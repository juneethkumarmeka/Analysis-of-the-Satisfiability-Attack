module basic_3000_30000_3500_6_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1120,In_2324);
nand U1 (N_1,In_993,In_2168);
nor U2 (N_2,In_2101,In_321);
nor U3 (N_3,In_2974,In_1556);
xnor U4 (N_4,In_2734,In_419);
xnor U5 (N_5,In_1196,In_2180);
nand U6 (N_6,In_402,In_1422);
or U7 (N_7,In_731,In_1642);
or U8 (N_8,In_2183,In_1036);
nand U9 (N_9,In_2259,In_1447);
nand U10 (N_10,In_34,In_2562);
nor U11 (N_11,In_2380,In_713);
nand U12 (N_12,In_172,In_791);
and U13 (N_13,In_1480,In_1550);
and U14 (N_14,In_2181,In_480);
or U15 (N_15,In_2772,In_716);
and U16 (N_16,In_1518,In_1271);
nand U17 (N_17,In_1652,In_35);
nor U18 (N_18,In_2241,In_96);
xor U19 (N_19,In_793,In_2938);
nand U20 (N_20,In_548,In_675);
and U21 (N_21,In_796,In_2091);
nand U22 (N_22,In_265,In_1640);
nand U23 (N_23,In_505,In_558);
or U24 (N_24,In_2114,In_2052);
or U25 (N_25,In_446,In_2461);
and U26 (N_26,In_515,In_2113);
xor U27 (N_27,In_1499,In_1723);
and U28 (N_28,In_1003,In_959);
nor U29 (N_29,In_928,In_2387);
nor U30 (N_30,In_1477,In_190);
or U31 (N_31,In_790,In_988);
nand U32 (N_32,In_563,In_2897);
nand U33 (N_33,In_2988,In_2149);
nand U34 (N_34,In_1688,In_2834);
and U35 (N_35,In_2264,In_32);
nand U36 (N_36,In_2673,In_2127);
and U37 (N_37,In_1472,In_2773);
and U38 (N_38,In_782,In_1620);
nand U39 (N_39,In_1114,In_207);
nand U40 (N_40,In_1337,In_593);
nand U41 (N_41,In_1947,In_2510);
nor U42 (N_42,In_1258,In_1430);
or U43 (N_43,In_1650,In_929);
nor U44 (N_44,In_1485,In_2458);
nand U45 (N_45,In_2158,In_1956);
or U46 (N_46,In_2295,In_2558);
nor U47 (N_47,In_2390,In_1040);
and U48 (N_48,In_2790,In_2551);
and U49 (N_49,In_651,In_483);
nor U50 (N_50,In_608,In_589);
or U51 (N_51,In_2234,In_1735);
nor U52 (N_52,In_1749,In_2396);
nor U53 (N_53,In_2316,In_2495);
xnor U54 (N_54,In_2742,In_2499);
and U55 (N_55,In_1884,In_654);
nand U56 (N_56,In_1299,In_1974);
or U57 (N_57,In_1561,In_2954);
nor U58 (N_58,In_1709,In_287);
nor U59 (N_59,In_1686,In_1403);
and U60 (N_60,In_1806,In_147);
and U61 (N_61,In_48,In_994);
nand U62 (N_62,In_2859,In_570);
nor U63 (N_63,In_1352,In_1641);
and U64 (N_64,In_2064,In_2015);
nor U65 (N_65,In_2927,In_2788);
or U66 (N_66,In_1533,In_1803);
nor U67 (N_67,In_1300,In_2069);
and U68 (N_68,In_77,In_2663);
xnor U69 (N_69,In_1910,In_1698);
and U70 (N_70,In_2167,In_1102);
or U71 (N_71,In_566,In_2642);
and U72 (N_72,In_1183,In_2753);
and U73 (N_73,In_1827,In_1629);
nor U74 (N_74,In_323,In_1333);
or U75 (N_75,In_161,In_1180);
nor U76 (N_76,In_2774,In_2508);
and U77 (N_77,In_1470,In_236);
nor U78 (N_78,In_191,In_2040);
nand U79 (N_79,In_1814,In_186);
nand U80 (N_80,In_441,In_359);
nand U81 (N_81,In_1763,In_657);
nor U82 (N_82,In_1232,In_1681);
nor U83 (N_83,In_243,In_1144);
nor U84 (N_84,In_387,In_1815);
or U85 (N_85,In_1573,In_2915);
nand U86 (N_86,In_58,In_322);
nand U87 (N_87,In_1809,In_2142);
or U88 (N_88,In_79,In_2115);
or U89 (N_89,In_653,In_1417);
or U90 (N_90,In_835,In_1607);
xnor U91 (N_91,In_1310,In_981);
nand U92 (N_92,In_2202,In_1972);
nor U93 (N_93,In_304,In_2802);
nor U94 (N_94,In_178,In_1828);
or U95 (N_95,In_2282,In_1553);
nor U96 (N_96,In_2146,In_2143);
and U97 (N_97,In_9,In_509);
nor U98 (N_98,In_57,In_478);
or U99 (N_99,In_2557,In_2166);
and U100 (N_100,In_2028,In_2949);
and U101 (N_101,In_2477,In_129);
nand U102 (N_102,In_2805,In_2366);
or U103 (N_103,In_760,In_2664);
or U104 (N_104,In_2189,In_2395);
or U105 (N_105,In_2197,In_299);
or U106 (N_106,In_1469,In_750);
nand U107 (N_107,In_1693,In_1013);
or U108 (N_108,In_842,In_1263);
nand U109 (N_109,In_1628,In_2615);
nor U110 (N_110,In_1708,In_1091);
and U111 (N_111,In_2036,In_954);
nor U112 (N_112,In_2945,In_2160);
xor U113 (N_113,In_904,In_808);
or U114 (N_114,In_1916,In_2090);
and U115 (N_115,In_2228,In_1960);
nor U116 (N_116,In_1172,In_1303);
and U117 (N_117,In_2951,In_720);
or U118 (N_118,In_2905,In_1181);
and U119 (N_119,In_702,In_2979);
nor U120 (N_120,In_1408,In_1928);
and U121 (N_121,In_893,In_156);
nor U122 (N_122,In_2864,In_683);
or U123 (N_123,In_2153,In_2590);
and U124 (N_124,In_2518,In_1679);
nor U125 (N_125,In_2850,In_1354);
and U126 (N_126,In_2039,In_2191);
nand U127 (N_127,In_1046,In_2381);
or U128 (N_128,In_2434,In_936);
nor U129 (N_129,In_2235,In_2047);
or U130 (N_130,In_409,In_1010);
xor U131 (N_131,In_1907,In_2330);
and U132 (N_132,In_2266,In_2061);
or U133 (N_133,In_137,In_405);
nor U134 (N_134,In_1311,In_229);
or U135 (N_135,In_2470,In_2074);
nand U136 (N_136,In_1504,In_396);
nand U137 (N_137,In_1820,In_1359);
nor U138 (N_138,In_1151,In_2471);
nor U139 (N_139,In_2591,In_1726);
nand U140 (N_140,In_1609,In_203);
nor U141 (N_141,In_2299,In_475);
nand U142 (N_142,In_1063,In_2781);
or U143 (N_143,In_1547,In_1881);
and U144 (N_144,In_1016,In_15);
and U145 (N_145,In_2710,In_2386);
nor U146 (N_146,In_1494,In_68);
or U147 (N_147,In_2797,In_2301);
nor U148 (N_148,In_1328,In_2870);
nand U149 (N_149,In_2447,In_457);
and U150 (N_150,In_195,In_2818);
nor U151 (N_151,In_1959,In_1022);
and U152 (N_152,In_1664,In_1478);
nor U153 (N_153,In_2478,In_2762);
nand U154 (N_154,In_2795,In_2020);
nand U155 (N_155,In_1836,In_920);
nand U156 (N_156,In_1255,In_2497);
nor U157 (N_157,In_635,In_1810);
nor U158 (N_158,In_1893,In_382);
nand U159 (N_159,In_2220,In_522);
or U160 (N_160,In_1946,In_2955);
or U161 (N_161,In_664,In_830);
and U162 (N_162,In_31,In_943);
and U163 (N_163,In_2904,In_426);
nand U164 (N_164,In_2021,In_1792);
nand U165 (N_165,In_2365,In_1692);
nor U166 (N_166,In_1505,In_2575);
and U167 (N_167,In_1855,In_2216);
and U168 (N_168,In_2674,In_818);
or U169 (N_169,In_1632,In_1018);
or U170 (N_170,In_392,In_184);
nor U171 (N_171,In_1211,In_365);
or U172 (N_172,In_1734,In_381);
nand U173 (N_173,In_792,In_1426);
or U174 (N_174,In_2851,In_2501);
or U175 (N_175,In_2319,In_2874);
and U176 (N_176,In_1848,In_541);
nor U177 (N_177,In_146,In_1621);
xor U178 (N_178,In_2082,In_757);
nor U179 (N_179,In_623,In_1130);
or U180 (N_180,In_1931,In_1405);
nor U181 (N_181,In_188,In_2637);
nor U182 (N_182,In_2199,In_1355);
xor U183 (N_183,In_756,In_170);
or U184 (N_184,In_2714,In_122);
nand U185 (N_185,In_1552,In_1966);
nand U186 (N_186,In_2880,In_6);
nand U187 (N_187,In_493,In_878);
xor U188 (N_188,In_55,In_2968);
and U189 (N_189,In_594,In_423);
nor U190 (N_190,In_1089,In_2875);
nand U191 (N_191,In_1161,In_843);
nand U192 (N_192,In_545,In_30);
and U193 (N_193,In_973,In_2981);
or U194 (N_194,In_1230,In_861);
nor U195 (N_195,In_1922,In_1979);
nor U196 (N_196,In_1812,In_1706);
xor U197 (N_197,In_228,In_1276);
xor U198 (N_198,In_99,In_105);
xnor U199 (N_199,In_733,In_2245);
and U200 (N_200,In_1218,In_1042);
and U201 (N_201,In_1381,In_2885);
or U202 (N_202,In_2249,In_741);
and U203 (N_203,In_931,In_2229);
or U204 (N_204,In_298,In_2690);
nand U205 (N_205,In_1746,In_2121);
or U206 (N_206,In_1983,In_2211);
nor U207 (N_207,In_2792,In_1982);
nand U208 (N_208,In_717,In_588);
and U209 (N_209,In_1944,In_2721);
or U210 (N_210,In_746,In_590);
nand U211 (N_211,In_992,In_1434);
or U212 (N_212,In_634,In_2572);
nand U213 (N_213,In_633,In_1326);
and U214 (N_214,In_1701,In_1203);
and U215 (N_215,In_347,In_2438);
or U216 (N_216,In_192,In_11);
and U217 (N_217,In_1129,In_1054);
and U218 (N_218,In_1794,In_2866);
and U219 (N_219,In_902,In_49);
xor U220 (N_220,In_544,In_2895);
nand U221 (N_221,In_1529,In_2007);
xnor U222 (N_222,In_2409,In_358);
and U223 (N_223,In_1158,In_513);
nand U224 (N_224,In_1514,In_1449);
and U225 (N_225,In_2527,In_2184);
nor U226 (N_226,In_425,In_1074);
and U227 (N_227,In_2588,In_1512);
nor U228 (N_228,In_2732,In_1256);
nor U229 (N_229,In_1630,In_2232);
nor U230 (N_230,In_1254,In_2983);
nand U231 (N_231,In_2129,In_1383);
nor U232 (N_232,In_831,In_1558);
and U233 (N_233,In_1275,In_2601);
and U234 (N_234,In_2822,In_2053);
xor U235 (N_235,In_766,In_2910);
xor U236 (N_236,In_1997,In_816);
and U237 (N_237,In_2454,In_985);
or U238 (N_238,In_1608,In_1797);
or U239 (N_239,In_2509,In_2860);
nand U240 (N_240,In_562,In_2374);
or U241 (N_241,In_1511,In_553);
and U242 (N_242,In_2190,In_2394);
nor U243 (N_243,In_2307,In_1007);
or U244 (N_244,In_2803,In_371);
and U245 (N_245,In_1740,In_277);
xor U246 (N_246,In_1564,In_2824);
or U247 (N_247,In_1549,In_1038);
nor U248 (N_248,In_519,In_2986);
or U249 (N_249,In_453,In_1534);
or U250 (N_250,In_2536,In_949);
nor U251 (N_251,In_526,In_957);
nand U252 (N_252,In_789,In_2956);
and U253 (N_253,In_1521,In_7);
xor U254 (N_254,In_2890,In_1577);
and U255 (N_255,In_727,In_967);
or U256 (N_256,In_571,In_2691);
and U257 (N_257,In_648,In_2088);
nand U258 (N_258,In_2760,In_1539);
and U259 (N_259,In_2472,In_596);
or U260 (N_260,In_1157,In_404);
xor U261 (N_261,In_1791,In_1567);
xnor U262 (N_262,In_303,In_1173);
and U263 (N_263,In_1115,In_1670);
nor U264 (N_264,In_1442,In_2619);
or U265 (N_265,In_1551,In_1135);
nand U266 (N_266,In_1327,In_771);
nor U267 (N_267,In_1025,In_1236);
nor U268 (N_268,In_2370,In_261);
and U269 (N_269,In_307,In_2273);
nand U270 (N_270,In_1186,In_1227);
or U271 (N_271,In_876,In_2672);
or U272 (N_272,In_1875,In_1546);
and U273 (N_273,In_24,In_1365);
nand U274 (N_274,In_2907,In_1741);
and U275 (N_275,In_865,In_242);
nor U276 (N_276,In_844,In_305);
or U277 (N_277,In_2328,In_338);
or U278 (N_278,In_2072,In_874);
and U279 (N_279,In_781,In_1479);
nand U280 (N_280,In_2119,In_2765);
and U281 (N_281,In_735,In_941);
nand U282 (N_282,In_1680,In_1147);
nand U283 (N_283,In_2679,In_2610);
nand U284 (N_284,In_529,In_1389);
nand U285 (N_285,In_2445,In_1523);
or U286 (N_286,In_1288,In_2185);
and U287 (N_287,In_2706,In_2489);
nor U288 (N_288,In_2013,In_1305);
and U289 (N_289,In_784,In_1773);
nor U290 (N_290,In_641,In_2027);
or U291 (N_291,In_2722,In_2128);
nor U292 (N_292,In_1660,In_1860);
nor U293 (N_293,In_336,In_1845);
nor U294 (N_294,In_2560,In_467);
and U295 (N_295,In_501,In_1164);
nor U296 (N_296,In_60,In_1678);
xor U297 (N_297,In_1039,In_987);
and U298 (N_298,In_2087,In_556);
nor U299 (N_299,In_2843,In_1729);
nand U300 (N_300,In_1919,In_1045);
and U301 (N_301,In_2656,In_1753);
nor U302 (N_302,In_1413,In_2215);
xor U303 (N_303,In_25,In_1483);
nor U304 (N_304,In_1341,In_2026);
or U305 (N_305,In_2066,In_5);
xnor U306 (N_306,In_2205,In_181);
nand U307 (N_307,In_944,In_2854);
and U308 (N_308,In_110,In_2737);
nor U309 (N_309,In_724,In_546);
nand U310 (N_310,In_1525,In_2704);
nor U311 (N_311,In_2046,In_1061);
nor U312 (N_312,In_1229,In_1962);
nand U313 (N_313,In_1099,In_1882);
nand U314 (N_314,In_921,In_132);
nand U315 (N_315,In_427,In_109);
nor U316 (N_316,In_1876,In_1116);
or U317 (N_317,In_1544,In_1414);
xnor U318 (N_318,In_1224,In_705);
or U319 (N_319,In_762,In_765);
and U320 (N_320,In_1588,In_2934);
nor U321 (N_321,In_1883,In_2868);
and U322 (N_322,In_2745,In_2561);
and U323 (N_323,In_1807,In_337);
nand U324 (N_324,In_348,In_451);
or U325 (N_325,In_1286,In_306);
nor U326 (N_326,In_385,In_1526);
nor U327 (N_327,In_1859,In_1323);
or U328 (N_328,In_2323,In_2349);
and U329 (N_329,In_1210,In_2775);
or U330 (N_330,In_1118,In_2353);
or U331 (N_331,In_330,In_1466);
nor U332 (N_332,In_268,In_2748);
nand U333 (N_333,In_1796,In_1360);
nand U334 (N_334,In_1293,In_1747);
nor U335 (N_335,In_899,In_1213);
xor U336 (N_336,In_209,In_690);
nor U337 (N_337,In_2586,In_897);
or U338 (N_338,In_1911,In_1362);
xnor U339 (N_339,In_880,In_1154);
xor U340 (N_340,In_1374,In_205);
and U341 (N_341,In_2102,In_1212);
and U342 (N_342,In_2278,In_2148);
nor U343 (N_343,In_1644,In_1395);
nor U344 (N_344,In_826,In_2195);
and U345 (N_345,In_492,In_1597);
or U346 (N_346,In_1216,In_2660);
and U347 (N_347,In_2720,In_1805);
nor U348 (N_348,In_1073,In_2545);
or U349 (N_349,In_2443,In_1586);
nand U350 (N_350,In_998,In_2914);
and U351 (N_351,In_2223,In_2923);
nor U352 (N_352,In_1481,In_176);
and U353 (N_353,In_532,In_2578);
nand U354 (N_354,In_269,In_92);
nor U355 (N_355,In_1456,In_617);
xor U356 (N_356,In_2118,In_1178);
or U357 (N_357,In_1937,In_1050);
nor U358 (N_358,In_230,In_130);
xnor U359 (N_359,In_2274,In_1611);
or U360 (N_360,In_1745,In_812);
nor U361 (N_361,In_964,In_1131);
nand U362 (N_362,In_2832,In_753);
and U363 (N_363,In_1078,In_1721);
or U364 (N_364,In_1712,In_136);
or U365 (N_365,In_2867,In_1268);
nor U366 (N_366,In_1606,In_1589);
and U367 (N_367,In_2780,In_471);
or U368 (N_368,In_700,In_2653);
nor U369 (N_369,In_389,In_2735);
nand U370 (N_370,In_2908,In_1965);
and U371 (N_371,In_1673,In_54);
or U372 (N_372,In_1339,In_2112);
nand U373 (N_373,In_615,In_1536);
nor U374 (N_374,In_1176,In_286);
and U375 (N_375,In_2889,In_1633);
xnor U376 (N_376,In_1555,In_461);
or U377 (N_377,In_583,In_1185);
or U378 (N_378,In_246,In_999);
and U379 (N_379,In_1237,In_552);
and U380 (N_380,In_2512,In_1361);
and U381 (N_381,In_1404,In_267);
nor U382 (N_382,In_2331,In_2516);
nand U383 (N_383,In_1108,In_1517);
nor U384 (N_384,In_460,In_890);
or U385 (N_385,In_512,In_1401);
nand U386 (N_386,In_1055,In_2617);
nor U387 (N_387,In_2188,In_142);
xnor U388 (N_388,In_2997,In_2280);
or U389 (N_389,In_1127,In_1927);
nor U390 (N_390,In_2863,In_2920);
nor U391 (N_391,In_2236,In_2618);
nor U392 (N_392,In_1064,In_2812);
nand U393 (N_393,In_2654,In_1731);
xor U394 (N_394,In_113,In_89);
and U395 (N_395,In_2446,In_915);
nand U396 (N_396,In_1051,In_46);
nand U397 (N_397,In_1319,In_1140);
or U398 (N_398,In_1802,In_2939);
and U399 (N_399,In_1231,In_759);
nor U400 (N_400,In_2755,In_1683);
nand U401 (N_401,In_1666,In_2621);
or U402 (N_402,In_1950,In_452);
nand U403 (N_403,In_2952,In_2784);
nand U404 (N_404,In_2998,In_914);
nand U405 (N_405,In_386,In_2203);
or U406 (N_406,In_1834,In_2507);
or U407 (N_407,In_1717,In_2752);
and U408 (N_408,In_2269,In_1122);
and U409 (N_409,In_1279,In_845);
and U410 (N_410,In_432,In_2369);
nand U411 (N_411,In_1580,In_665);
nand U412 (N_412,In_2918,In_282);
nand U413 (N_413,In_625,In_1508);
and U414 (N_414,In_2542,In_1832);
nand U415 (N_415,In_1134,In_279);
or U416 (N_416,In_2043,In_2255);
or U417 (N_417,In_496,In_1843);
nor U418 (N_418,In_1155,In_114);
nand U419 (N_419,In_828,In_2182);
nand U420 (N_420,In_2268,In_150);
nor U421 (N_421,In_2347,In_1424);
nor U422 (N_422,In_2999,In_106);
or U423 (N_423,In_2627,In_2756);
and U424 (N_424,In_2703,In_506);
nand U425 (N_425,In_104,In_1385);
nand U426 (N_426,In_316,In_2547);
xnor U427 (N_427,In_2921,In_732);
and U428 (N_428,In_855,In_2849);
or U429 (N_429,In_2935,In_2670);
or U430 (N_430,In_1639,In_1380);
or U431 (N_431,In_1696,In_619);
nor U432 (N_432,In_573,In_2420);
nor U433 (N_433,In_885,In_174);
or U434 (N_434,In_1861,In_1418);
nand U435 (N_435,In_1065,In_2503);
or U436 (N_436,In_1266,In_2916);
or U437 (N_437,In_2777,In_2985);
nor U438 (N_438,In_1363,In_543);
nand U439 (N_439,In_807,In_1128);
nand U440 (N_440,In_429,In_2894);
and U441 (N_441,In_701,In_1261);
xnor U442 (N_442,In_1874,In_2452);
xor U443 (N_443,In_829,In_525);
and U444 (N_444,In_308,In_2389);
nand U445 (N_445,In_1234,In_1501);
nand U446 (N_446,In_1917,In_1044);
nand U447 (N_447,In_2522,In_281);
nor U448 (N_448,In_997,In_1159);
or U449 (N_449,In_1566,In_2544);
and U450 (N_450,In_250,In_313);
xor U451 (N_451,In_1304,In_591);
and U452 (N_452,In_155,In_661);
or U453 (N_453,In_1011,In_817);
or U454 (N_454,In_2429,In_2716);
nor U455 (N_455,In_1087,In_88);
or U456 (N_456,In_1357,In_827);
or U457 (N_457,In_2624,In_1601);
or U458 (N_458,In_800,In_2929);
nor U459 (N_459,In_925,In_2511);
and U460 (N_460,In_1223,In_1842);
or U461 (N_461,In_946,In_1795);
xnor U462 (N_462,In_1668,In_2661);
nor U463 (N_463,In_2622,In_620);
nand U464 (N_464,In_231,In_52);
nand U465 (N_465,In_442,In_798);
nor U466 (N_466,In_1220,In_204);
nand U467 (N_467,In_1622,In_2367);
nand U468 (N_468,In_1789,In_1379);
xor U469 (N_469,In_1866,In_1557);
and U470 (N_470,In_1503,In_390);
nor U471 (N_471,In_2899,In_1110);
xor U472 (N_472,In_1728,In_2521);
nor U473 (N_473,In_2530,In_2778);
nand U474 (N_474,In_578,In_325);
nand U475 (N_475,In_2933,In_2265);
and U476 (N_476,In_1737,In_710);
and U477 (N_477,In_709,In_2094);
nand U478 (N_478,In_2540,In_2906);
nand U479 (N_479,In_399,In_226);
nand U480 (N_480,In_561,In_863);
and U481 (N_481,In_1345,In_1992);
or U482 (N_482,In_1847,In_63);
nand U483 (N_483,In_1800,In_1015);
nor U484 (N_484,In_2599,In_2702);
nor U485 (N_485,In_1782,In_1491);
nand U486 (N_486,In_847,In_2873);
and U487 (N_487,In_2635,In_454);
nand U488 (N_488,In_1986,In_802);
and U489 (N_489,In_2277,In_1459);
and U490 (N_490,In_485,In_430);
nor U491 (N_491,In_82,In_2807);
and U492 (N_492,In_2333,In_2965);
or U493 (N_493,In_2694,In_1583);
nand U494 (N_494,In_2827,In_1954);
and U495 (N_495,In_695,In_1098);
nor U496 (N_496,In_832,In_2723);
xor U497 (N_497,In_1160,In_990);
or U498 (N_498,In_1192,In_1700);
nor U499 (N_499,In_1468,In_1507);
nand U500 (N_500,In_2804,In_1985);
or U501 (N_501,In_1069,In_1981);
and U502 (N_502,In_1891,In_747);
nand U503 (N_503,In_2413,In_916);
nor U504 (N_504,In_2354,In_90);
or U505 (N_505,In_484,In_734);
and U506 (N_506,In_2237,In_463);
nor U507 (N_507,In_610,In_1971);
nand U508 (N_508,In_2491,In_860);
nor U509 (N_509,In_2246,In_627);
nand U510 (N_510,In_2383,In_241);
xnor U511 (N_511,In_489,In_2371);
and U512 (N_512,In_47,In_975);
and U513 (N_513,In_1209,In_1493);
and U514 (N_514,In_349,In_822);
nand U515 (N_515,In_586,In_712);
nor U516 (N_516,In_1190,In_2825);
nor U517 (N_517,In_2037,In_912);
nand U518 (N_518,In_1888,In_29);
or U519 (N_519,In_1301,In_2541);
nand U520 (N_520,In_2857,In_1646);
or U521 (N_521,In_41,In_2171);
or U522 (N_522,In_887,In_2937);
nor U523 (N_523,In_194,In_1579);
xor U524 (N_524,In_94,In_723);
nor U525 (N_525,In_1532,In_1427);
or U526 (N_526,In_1121,In_183);
or U527 (N_527,In_1153,In_1373);
or U528 (N_528,In_2029,In_1314);
nand U529 (N_529,In_2976,In_788);
and U530 (N_530,In_2571,In_768);
and U531 (N_531,In_50,In_2267);
or U532 (N_532,In_1587,In_2602);
and U533 (N_533,In_1667,In_1744);
nand U534 (N_534,In_1980,In_2177);
nand U535 (N_535,In_2163,In_2816);
or U536 (N_536,In_2798,In_1243);
or U537 (N_537,In_1315,In_2482);
nand U538 (N_538,In_115,In_602);
nor U539 (N_539,In_2936,In_838);
nand U540 (N_540,In_2150,In_2977);
or U541 (N_541,In_2724,In_646);
and U542 (N_542,In_1068,In_1446);
xnor U543 (N_543,In_1008,In_2698);
xor U544 (N_544,In_2201,In_1382);
or U545 (N_545,In_456,In_2829);
or U546 (N_546,In_2179,In_1535);
nor U547 (N_547,In_1189,In_368);
and U548 (N_548,In_445,In_811);
nand U549 (N_549,In_1017,In_256);
and U550 (N_550,In_2479,In_196);
nor U551 (N_551,In_2071,In_1562);
or U552 (N_552,In_1021,In_2140);
xnor U553 (N_553,In_2480,In_1793);
or U554 (N_554,In_1242,In_383);
or U555 (N_555,In_1977,In_1248);
and U556 (N_556,In_2131,In_1287);
and U557 (N_557,In_2884,In_2809);
or U558 (N_558,In_1614,In_1428);
xor U559 (N_559,In_2343,In_1733);
and U560 (N_560,In_27,In_864);
nor U561 (N_561,In_523,In_849);
nand U562 (N_562,In_1384,In_2808);
or U563 (N_563,In_1005,In_783);
nand U564 (N_564,In_225,In_437);
and U565 (N_565,In_13,In_2687);
and U566 (N_566,In_2651,In_2835);
nor U567 (N_567,In_2948,In_879);
nand U568 (N_568,In_687,In_1591);
or U569 (N_569,In_251,In_33);
or U570 (N_570,In_479,In_2891);
or U571 (N_571,In_2041,In_2194);
and U572 (N_572,In_2625,In_119);
and U573 (N_573,In_2432,In_36);
nand U574 (N_574,In_502,In_1704);
or U575 (N_575,In_2842,In_1902);
xnor U576 (N_576,In_2644,In_393);
nor U577 (N_577,In_1391,In_821);
or U578 (N_578,In_1169,In_909);
nand U579 (N_579,In_889,In_318);
xor U580 (N_580,In_1062,In_1171);
or U581 (N_581,In_1085,In_416);
and U582 (N_582,In_1431,In_2418);
and U583 (N_583,In_2392,In_2972);
and U584 (N_584,In_1879,In_1057);
xor U585 (N_585,In_1510,In_19);
nor U586 (N_586,In_640,In_2603);
nand U587 (N_587,In_1892,In_1351);
and U588 (N_588,In_528,In_2213);
xnor U589 (N_589,In_1020,In_2490);
nand U590 (N_590,In_1163,In_2248);
nand U591 (N_591,In_1071,In_953);
and U592 (N_592,In_1463,In_1425);
or U593 (N_593,In_854,In_962);
nor U594 (N_594,In_1941,In_2145);
or U595 (N_595,In_1784,In_2730);
nand U596 (N_596,In_2526,In_1296);
xor U597 (N_597,In_825,In_1249);
nor U598 (N_598,In_103,In_806);
nand U599 (N_599,In_2327,In_1410);
or U600 (N_600,In_1592,In_2065);
nor U601 (N_601,In_1623,In_794);
nor U602 (N_602,In_1838,In_1756);
and U603 (N_603,In_872,In_840);
nor U604 (N_604,In_2304,In_1291);
nor U605 (N_605,In_2993,In_2626);
or U606 (N_606,In_2106,In_2964);
or U607 (N_607,In_947,In_2961);
or U608 (N_608,In_1336,In_1766);
nand U609 (N_609,In_2671,In_2514);
or U610 (N_610,In_1610,In_2441);
and U611 (N_611,In_2982,In_1940);
xor U612 (N_612,In_1676,In_477);
nand U613 (N_613,In_1772,In_770);
and U614 (N_614,In_1202,In_1318);
and U615 (N_615,In_1295,In_2636);
nor U616 (N_616,In_1002,In_1790);
and U617 (N_617,In_2098,In_351);
nand U618 (N_618,In_850,In_2533);
or U619 (N_619,In_632,In_2502);
nor U620 (N_620,In_44,In_2309);
xor U621 (N_621,In_1294,In_1376);
or U622 (N_622,In_2840,In_152);
and U623 (N_623,In_1872,In_2204);
xnor U624 (N_624,In_551,In_2285);
nand U625 (N_625,In_1719,In_2589);
xor U626 (N_626,In_2493,In_630);
and U627 (N_627,In_1975,In_2574);
nor U628 (N_628,In_2110,In_1083);
nand U629 (N_629,In_1387,In_2097);
or U630 (N_630,In_2310,In_108);
nor U631 (N_631,In_2957,In_2813);
and U632 (N_632,In_595,In_1056);
or U633 (N_633,In_1452,In_2791);
xor U634 (N_634,In_1125,In_2496);
and U635 (N_635,In_2608,In_2684);
nor U636 (N_636,In_1049,In_2892);
and U637 (N_637,In_2911,In_984);
nand U638 (N_638,In_682,In_1043);
nand U639 (N_639,In_1167,In_2308);
and U640 (N_640,In_1104,In_2500);
and U641 (N_641,In_1409,In_331);
and U642 (N_642,In_857,In_379);
nor U643 (N_643,In_737,In_2862);
nor U644 (N_644,In_934,In_1331);
nor U645 (N_645,In_1575,In_1306);
nand U646 (N_646,In_2523,In_728);
or U647 (N_647,In_1335,In_1545);
nor U648 (N_648,In_584,In_1075);
xnor U649 (N_649,In_232,In_2073);
and U650 (N_650,In_1509,In_2594);
nor U651 (N_651,In_2172,In_2959);
and U652 (N_652,In_2341,In_2322);
or U653 (N_653,In_290,In_752);
or U654 (N_654,In_1097,In_2398);
nor U655 (N_655,In_868,In_1933);
nand U656 (N_656,In_2431,In_1101);
and U657 (N_657,In_1031,In_2067);
or U658 (N_658,In_913,In_1554);
and U659 (N_659,In_898,In_326);
nand U660 (N_660,In_1563,In_197);
nand U661 (N_661,In_2379,In_873);
nand U662 (N_662,In_924,In_2973);
nor U663 (N_663,In_1458,In_210);
or U664 (N_664,In_2406,In_23);
and U665 (N_665,In_126,In_102);
xnor U666 (N_666,In_2411,In_310);
nand U667 (N_667,In_2002,In_1613);
or U668 (N_668,In_1117,In_1433);
xor U669 (N_669,In_2117,In_2726);
nand U670 (N_670,In_1369,In_123);
or U671 (N_671,In_1060,In_2096);
or U672 (N_672,In_542,In_2225);
nand U673 (N_673,In_1201,In_2693);
nand U674 (N_674,In_2290,In_2796);
or U675 (N_675,In_2946,In_361);
nand U676 (N_676,In_2176,In_244);
nand U677 (N_677,In_1035,In_2334);
nor U678 (N_678,In_2050,In_1605);
nor U679 (N_679,In_2686,In_375);
and U680 (N_680,In_2404,In_2980);
nor U681 (N_681,In_2524,In_1877);
nor U682 (N_682,In_580,In_71);
and U683 (N_683,In_1991,In_373);
or U684 (N_684,In_2633,In_2419);
and U685 (N_685,In_2093,In_2917);
nor U686 (N_686,In_1471,In_1730);
or U687 (N_687,In_117,In_2567);
and U688 (N_688,In_2083,In_659);
or U689 (N_689,In_481,In_1262);
xnor U690 (N_690,In_2134,In_2666);
nand U691 (N_691,In_2990,In_2350);
and U692 (N_692,In_332,In_2095);
nor U693 (N_693,In_447,In_2212);
and U694 (N_694,In_1636,In_2318);
and U695 (N_695,In_688,In_1070);
xnor U696 (N_696,In_1393,In_293);
xnor U697 (N_697,In_1844,In_574);
xnor U698 (N_698,In_2358,In_1833);
nand U699 (N_699,In_814,In_2793);
and U700 (N_700,In_748,In_1949);
and U701 (N_701,In_3,In_886);
or U702 (N_702,In_521,In_1894);
nand U703 (N_703,In_958,In_1253);
nor U704 (N_704,In_2159,In_1252);
nor U705 (N_705,In_2450,In_1869);
or U706 (N_706,In_2057,In_328);
and U707 (N_707,In_2484,In_2062);
nand U708 (N_708,In_1152,In_531);
xor U709 (N_709,In_2227,In_61);
and U710 (N_710,In_1206,In_2833);
nand U711 (N_711,In_364,In_974);
xor U712 (N_712,In_2869,In_2435);
or U713 (N_713,In_1710,In_2410);
nor U714 (N_714,In_1955,In_488);
nand U715 (N_715,In_926,In_1217);
nand U716 (N_716,In_1625,In_407);
xor U717 (N_717,In_118,In_2239);
nand U718 (N_718,In_2244,In_2);
and U719 (N_719,In_1969,In_1811);
or U720 (N_720,In_2531,In_869);
or U721 (N_721,In_1758,In_841);
nor U722 (N_722,In_761,In_862);
and U723 (N_723,In_2931,In_2133);
and U724 (N_724,In_922,In_951);
and U725 (N_725,In_249,In_2359);
nor U726 (N_726,In_2132,In_2405);
nor U727 (N_727,In_2439,In_1432);
nor U728 (N_728,In_51,In_292);
nor U729 (N_729,In_2733,In_670);
nand U730 (N_730,In_2942,In_177);
nor U731 (N_731,In_1267,In_1476);
or U732 (N_732,In_1334,In_2763);
and U733 (N_733,In_1032,In_813);
nor U734 (N_734,In_1394,In_2563);
nor U735 (N_735,In_227,In_2596);
nand U736 (N_736,In_1088,In_2397);
or U737 (N_737,In_961,In_2958);
nand U738 (N_738,In_1958,In_1245);
or U739 (N_739,In_2221,In_1325);
nand U740 (N_740,In_1761,In_538);
nor U741 (N_741,In_237,In_918);
and U742 (N_742,In_1615,In_1119);
nor U743 (N_743,In_2006,In_17);
or U744 (N_744,In_1901,In_1771);
xnor U745 (N_745,In_2224,In_697);
or U746 (N_746,In_671,In_2462);
xnor U747 (N_747,In_1873,In_1265);
or U748 (N_748,In_910,In_662);
and U749 (N_749,In_2423,In_1578);
nand U750 (N_750,In_2576,In_1093);
or U751 (N_751,In_2054,In_1221);
nand U752 (N_752,In_749,In_21);
and U753 (N_753,In_2534,In_976);
and U754 (N_754,In_1297,In_202);
nand U755 (N_755,In_2616,In_1461);
or U756 (N_756,In_148,In_258);
or U757 (N_757,In_1465,In_819);
and U758 (N_758,In_2293,In_1783);
nor U759 (N_759,In_2436,In_266);
nor U760 (N_760,In_1926,In_2077);
and U761 (N_761,In_472,In_2697);
nand U762 (N_762,In_464,In_2841);
nor U763 (N_763,In_1849,In_1978);
nand U764 (N_764,In_2055,In_93);
nand U765 (N_765,In_575,In_1429);
nor U766 (N_766,In_1411,In_1938);
and U767 (N_767,In_2539,In_2887);
nor U768 (N_768,In_2284,In_0);
and U769 (N_769,In_1250,In_1490);
or U770 (N_770,In_2103,In_1024);
xor U771 (N_771,In_587,In_39);
nor U772 (N_772,In_415,In_626);
nand U773 (N_773,In_271,In_2058);
nand U774 (N_774,In_2712,In_1527);
nor U775 (N_775,In_1825,In_2583);
or U776 (N_776,In_2107,In_2975);
and U777 (N_777,In_2893,In_1531);
or U778 (N_778,In_1840,In_1829);
nand U779 (N_779,In_1624,In_2056);
nand U780 (N_780,In_1498,In_459);
or U781 (N_781,In_1457,In_40);
nand U782 (N_782,In_1662,In_2402);
nand U783 (N_783,In_568,In_1694);
or U784 (N_784,In_1388,In_377);
nand U785 (N_785,In_721,In_411);
or U786 (N_786,In_940,In_763);
or U787 (N_787,In_2296,In_80);
or U788 (N_788,In_421,In_2584);
or U789 (N_789,In_2217,In_2108);
and U790 (N_790,In_2984,In_883);
and U791 (N_791,In_2313,In_1885);
xor U792 (N_792,In_2453,In_866);
nand U793 (N_793,In_1289,In_2692);
nand U794 (N_794,In_2794,In_2678);
and U795 (N_795,In_2700,In_498);
or U796 (N_796,In_607,In_2747);
and U797 (N_797,In_2815,In_892);
and U798 (N_798,In_212,In_16);
nor U799 (N_799,In_621,In_1090);
and U800 (N_800,In_2782,In_2414);
and U801 (N_801,In_1308,In_2338);
and U802 (N_802,In_2799,In_1542);
and U803 (N_803,In_1540,In_354);
nand U804 (N_804,In_2378,In_2909);
and U805 (N_805,In_1748,In_647);
or U806 (N_806,In_2659,In_56);
or U807 (N_807,In_280,In_2048);
or U808 (N_808,In_1900,In_534);
or U809 (N_809,In_2900,In_668);
or U810 (N_810,In_1661,In_932);
and U811 (N_811,In_1538,In_1780);
nor U812 (N_812,In_1852,In_2085);
or U813 (N_813,In_2260,In_666);
nor U814 (N_814,In_2978,In_1939);
xor U815 (N_815,In_222,In_1909);
or U816 (N_816,In_1895,In_2068);
nor U817 (N_817,In_206,In_2016);
or U818 (N_818,In_1572,In_1081);
and U819 (N_819,In_1718,In_1139);
or U820 (N_820,In_637,In_1215);
nor U821 (N_821,In_1441,In_158);
nand U822 (N_822,In_660,In_1397);
nor U823 (N_823,In_554,In_439);
and U824 (N_824,In_1801,In_2675);
and U825 (N_825,In_1626,In_1407);
nor U826 (N_826,In_772,In_1651);
or U827 (N_827,In_1506,In_956);
nand U828 (N_828,In_2342,In_2162);
nand U829 (N_829,In_612,In_1942);
and U830 (N_830,In_240,In_1175);
xnor U831 (N_831,In_1496,In_1858);
and U832 (N_832,In_1779,In_2628);
or U833 (N_833,In_288,In_1482);
and U834 (N_834,In_2779,In_1821);
and U835 (N_835,In_614,In_1371);
nor U836 (N_836,In_2126,In_1200);
or U837 (N_837,In_1019,In_2151);
nor U838 (N_838,In_1000,In_674);
and U839 (N_839,In_1241,In_2593);
nand U840 (N_840,In_1813,In_2665);
xnor U841 (N_841,In_2078,In_164);
and U842 (N_842,In_785,In_2846);
nor U843 (N_843,In_517,In_2196);
nor U844 (N_844,In_1631,In_714);
or U845 (N_845,In_1390,In_642);
nor U846 (N_846,In_567,In_1896);
nand U847 (N_847,In_2385,In_1837);
and U848 (N_848,In_858,In_2360);
nor U849 (N_849,In_725,In_1439);
and U850 (N_850,In_2377,In_745);
or U851 (N_851,In_2130,In_1251);
nor U852 (N_852,In_1774,In_1246);
nand U853 (N_853,In_1785,In_4);
or U854 (N_854,In_965,In_1649);
or U855 (N_855,In_2218,In_900);
xnor U856 (N_856,In_458,In_329);
nand U857 (N_857,In_680,In_1460);
nor U858 (N_858,In_1402,In_2681);
nand U859 (N_859,In_2883,In_140);
or U860 (N_860,In_1489,In_2597);
nor U861 (N_861,In_622,In_618);
and U862 (N_862,In_2161,In_2853);
and U863 (N_863,In_2049,In_257);
nor U864 (N_864,In_719,In_2744);
or U865 (N_865,In_66,In_144);
or U866 (N_866,In_1370,In_773);
and U867 (N_867,In_1324,In_2012);
xor U868 (N_868,In_1332,In_2532);
nand U869 (N_869,In_417,In_1166);
and U870 (N_870,In_2550,In_2481);
and U871 (N_871,In_2519,In_1925);
or U872 (N_872,In_134,In_1145);
or U873 (N_873,In_2643,In_1675);
nor U874 (N_874,In_499,In_1034);
and U875 (N_875,In_2932,In_795);
nand U876 (N_876,In_903,In_2766);
nor U877 (N_877,In_1770,In_1219);
and U878 (N_878,In_1313,In_438);
and U879 (N_879,In_1871,In_969);
and U880 (N_880,In_278,In_1776);
nand U881 (N_881,In_422,In_420);
nand U882 (N_882,In_1228,In_1618);
nor U883 (N_883,In_1781,In_138);
nand U884 (N_884,In_376,In_1951);
nor U885 (N_885,In_233,In_2831);
nor U886 (N_886,In_2170,In_245);
nor U887 (N_887,In_2709,In_1270);
and U888 (N_888,In_2314,In_2966);
and U889 (N_889,In_2751,In_1707);
or U890 (N_890,In_1619,In_2018);
or U891 (N_891,In_2579,In_145);
nand U892 (N_892,In_2287,In_2876);
xor U893 (N_893,In_952,In_218);
or U894 (N_894,In_2005,In_2346);
nor U895 (N_895,In_291,In_2252);
and U896 (N_896,In_960,In_363);
nor U897 (N_897,In_972,In_2657);
nand U898 (N_898,In_613,In_950);
or U899 (N_899,In_905,In_1519);
nor U900 (N_900,In_1353,In_1897);
and U901 (N_901,In_1863,In_1999);
and U902 (N_902,In_684,In_1415);
nor U903 (N_903,In_302,In_1934);
nor U904 (N_904,In_743,In_497);
nand U905 (N_905,In_516,In_2620);
or U906 (N_906,In_945,In_2024);
and U907 (N_907,In_1027,In_2944);
or U908 (N_908,In_2922,In_2157);
or U909 (N_909,In_600,In_83);
nand U910 (N_910,In_2467,In_2124);
and U911 (N_911,In_214,In_1092);
nand U912 (N_912,In_2294,In_2960);
nand U913 (N_913,In_2577,In_1349);
or U914 (N_914,In_65,In_933);
nor U915 (N_915,In_579,In_1112);
or U916 (N_916,In_1560,In_1124);
nand U917 (N_917,In_1445,In_8);
or U918 (N_918,In_2950,In_2311);
nor U919 (N_919,In_2164,In_1474);
nor U920 (N_920,In_1816,In_180);
nand U921 (N_921,In_2600,In_73);
or U922 (N_922,In_1455,In_1416);
or U923 (N_923,In_1240,In_669);
xor U924 (N_924,In_317,In_601);
or U925 (N_925,In_638,In_2075);
and U926 (N_926,In_1994,In_2032);
nor U927 (N_927,In_1137,In_1993);
and U928 (N_928,In_1687,In_955);
nor U929 (N_929,In_2941,In_1870);
nand U930 (N_930,In_2553,In_1146);
xnor U931 (N_931,In_2076,In_2451);
and U932 (N_932,In_2427,In_2676);
or U933 (N_933,In_2559,In_1149);
and U934 (N_934,In_1138,In_1819);
and U935 (N_935,In_1136,In_2487);
or U936 (N_936,In_97,In_1344);
nor U937 (N_937,In_1193,In_2830);
nand U938 (N_938,In_1274,In_2852);
or U939 (N_939,In_1823,In_1086);
and U940 (N_940,In_1760,In_2104);
nand U941 (N_941,In_1697,In_2344);
and U942 (N_942,In_1759,In_1317);
nand U943 (N_943,In_2492,In_2038);
or U944 (N_944,In_2464,In_2222);
and U945 (N_945,In_143,In_888);
or U946 (N_946,In_2200,In_2630);
nand U947 (N_947,In_1400,In_1648);
nor U948 (N_948,In_343,In_804);
and U949 (N_949,In_1932,In_938);
xnor U950 (N_950,In_2345,In_2844);
nand U951 (N_951,In_2727,In_2658);
nand U952 (N_952,In_2498,In_2460);
nand U953 (N_953,In_2109,In_1364);
or U954 (N_954,In_2483,In_2810);
nor U955 (N_955,In_2306,In_1596);
and U956 (N_956,In_2468,In_547);
nor U957 (N_957,In_1348,In_1235);
or U958 (N_958,In_78,In_64);
xnor U959 (N_959,In_424,In_1616);
nor U960 (N_960,In_1132,In_663);
nand U961 (N_961,In_1346,In_200);
and U962 (N_962,In_2302,In_2401);
or U963 (N_963,In_2611,In_980);
or U964 (N_964,In_576,In_673);
and U965 (N_965,In_2995,In_2415);
nor U966 (N_966,In_2060,In_2486);
or U967 (N_967,In_2595,In_2819);
nor U968 (N_968,In_1585,In_1582);
nor U969 (N_969,In_2384,In_2254);
nor U970 (N_970,In_2786,In_718);
nor U971 (N_971,In_1905,In_1853);
nand U972 (N_972,In_2582,In_440);
or U973 (N_973,In_815,In_189);
or U974 (N_974,In_162,In_98);
nor U975 (N_975,In_2155,In_1123);
nand U976 (N_976,In_2647,In_1113);
nand U977 (N_977,In_2634,In_2357);
nor U978 (N_978,In_2994,In_2023);
and U979 (N_979,In_1943,In_2240);
xnor U980 (N_980,In_2736,In_2506);
or U981 (N_981,In_1156,In_2382);
xnor U982 (N_982,In_518,In_2650);
nand U983 (N_983,In_2407,In_1581);
nor U984 (N_984,In_1690,In_428);
nand U985 (N_985,In_474,In_2930);
and U986 (N_986,In_272,In_252);
nand U987 (N_987,In_1864,In_585);
nor U988 (N_988,In_1281,In_139);
nor U989 (N_989,In_38,In_179);
or U990 (N_990,In_2283,In_2474);
nor U991 (N_991,In_2456,In_1953);
nor U992 (N_992,In_315,In_1674);
xor U993 (N_993,In_650,In_1576);
nor U994 (N_994,In_539,In_12);
and U995 (N_995,In_2351,In_1787);
or U996 (N_996,In_201,In_769);
nor U997 (N_997,In_1665,In_1537);
nor U998 (N_998,In_2136,In_208);
or U999 (N_999,In_1967,In_1998);
nor U1000 (N_1000,In_678,In_45);
xnor U1001 (N_1001,In_2238,In_636);
nor U1002 (N_1002,In_977,In_2352);
or U1003 (N_1003,In_691,In_1435);
or U1004 (N_1004,In_2001,In_1148);
nand U1005 (N_1005,In_1280,In_1058);
nor U1006 (N_1006,In_520,In_2640);
xor U1007 (N_1007,In_100,In_1908);
or U1008 (N_1008,In_2198,In_894);
or U1009 (N_1009,In_2421,In_1654);
or U1010 (N_1010,In_1272,In_221);
or U1011 (N_1011,In_1316,In_645);
nand U1012 (N_1012,In_2174,In_408);
nor U1013 (N_1013,In_1444,In_1913);
and U1014 (N_1014,In_1617,In_1225);
nor U1015 (N_1015,In_69,In_2465);
nor U1016 (N_1016,In_2044,In_848);
and U1017 (N_1017,In_2789,In_2100);
nor U1018 (N_1018,In_2475,In_1358);
nand U1019 (N_1019,In_1298,In_1565);
and U1020 (N_1020,In_10,In_1107);
and U1021 (N_1021,In_2123,In_1851);
nand U1022 (N_1022,In_2122,In_2592);
nor U1023 (N_1023,In_353,In_1467);
and U1024 (N_1024,In_739,In_2321);
or U1025 (N_1025,In_2326,In_470);
or U1026 (N_1026,In_141,In_616);
xnor U1027 (N_1027,In_1672,In_1808);
or U1028 (N_1028,In_1473,In_2715);
nor U1029 (N_1029,In_2286,In_211);
or U1030 (N_1030,In_1222,In_157);
or U1031 (N_1031,In_2886,In_2317);
nor U1032 (N_1032,In_1804,In_859);
and U1033 (N_1033,In_942,In_1584);
nand U1034 (N_1034,In_834,In_1322);
nor U1035 (N_1035,In_223,In_906);
nand U1036 (N_1036,In_297,In_1725);
xnor U1037 (N_1037,In_1961,In_418);
nor U1038 (N_1038,In_199,In_163);
nand U1039 (N_1039,In_986,In_1590);
nor U1040 (N_1040,In_1769,In_264);
nand U1041 (N_1041,In_639,In_937);
or U1042 (N_1042,In_2556,In_309);
or U1043 (N_1043,In_2251,In_2645);
and U1044 (N_1044,In_882,In_2449);
nand U1045 (N_1045,In_2925,In_2362);
nand U1046 (N_1046,In_270,In_2505);
and U1047 (N_1047,In_1936,In_643);
nand U1048 (N_1048,In_1484,In_527);
nor U1049 (N_1049,In_219,In_1420);
or U1050 (N_1050,In_403,In_1682);
and U1051 (N_1051,In_2568,In_1386);
xor U1052 (N_1052,In_296,In_2783);
and U1053 (N_1053,In_871,In_1320);
and U1054 (N_1054,In_187,In_1283);
xnor U1055 (N_1055,In_2165,In_1052);
or U1056 (N_1056,In_1205,In_1378);
nor U1057 (N_1057,In_1399,In_1865);
nor U1058 (N_1058,In_597,In_1750);
nor U1059 (N_1059,In_2086,In_2272);
or U1060 (N_1060,In_2303,In_2139);
and U1061 (N_1061,In_2708,In_535);
nand U1062 (N_1062,In_1976,In_2070);
or U1063 (N_1063,In_1290,In_740);
nor U1064 (N_1064,In_1996,In_220);
nand U1065 (N_1065,In_706,In_1368);
nand U1066 (N_1066,In_1691,In_1657);
xor U1067 (N_1067,In_2837,In_1973);
and U1068 (N_1068,In_2652,In_466);
nor U1069 (N_1069,In_2872,In_234);
nor U1070 (N_1070,In_1645,In_435);
or U1071 (N_1071,In_2000,In_2648);
nand U1072 (N_1072,In_1889,In_1030);
nand U1073 (N_1073,In_2156,In_1059);
and U1074 (N_1074,In_1239,In_2888);
and U1075 (N_1075,In_2520,In_301);
or U1076 (N_1076,In_2817,In_510);
and U1077 (N_1077,In_62,In_372);
or U1078 (N_1078,In_312,In_1722);
or U1079 (N_1079,In_2417,In_1195);
nand U1080 (N_1080,In_2356,In_1685);
nand U1081 (N_1081,In_681,In_160);
nand U1082 (N_1082,In_694,In_2543);
and U1083 (N_1083,In_2080,In_2913);
or U1084 (N_1084,In_1856,In_799);
nand U1085 (N_1085,In_2416,In_1257);
nor U1086 (N_1086,In_1593,In_1912);
or U1087 (N_1087,In_604,In_1817);
xnor U1088 (N_1088,In_557,In_494);
or U1089 (N_1089,In_1464,In_1486);
nor U1090 (N_1090,In_2448,In_2811);
nand U1091 (N_1091,In_1495,In_107);
nor U1092 (N_1092,In_2175,In_1072);
nand U1093 (N_1093,In_1903,In_2668);
and U1094 (N_1094,In_1492,In_274);
nand U1095 (N_1095,In_1755,In_1440);
and U1096 (N_1096,In_2738,In_1739);
and U1097 (N_1097,In_1259,In_1421);
nand U1098 (N_1098,In_2528,In_1497);
nand U1099 (N_1099,In_1292,In_1775);
nand U1100 (N_1100,In_2529,In_1450);
and U1101 (N_1101,In_891,In_2288);
nor U1102 (N_1102,In_1500,In_2403);
nand U1103 (N_1103,In_2963,In_1406);
nand U1104 (N_1104,In_1026,In_111);
or U1105 (N_1105,In_1990,In_1207);
nand U1106 (N_1106,In_1366,In_84);
nand U1107 (N_1107,In_1935,In_1029);
xnor U1108 (N_1108,In_2667,In_2473);
or U1109 (N_1109,In_1177,In_2879);
nand U1110 (N_1110,In_2746,In_1702);
and U1111 (N_1111,In_852,In_982);
or U1112 (N_1112,In_692,In_1915);
or U1113 (N_1113,In_394,In_1392);
and U1114 (N_1114,In_2685,In_628);
nor U1115 (N_1115,In_1278,In_2771);
xor U1116 (N_1116,In_2555,In_2372);
and U1117 (N_1117,In_1930,In_2928);
xnor U1118 (N_1118,In_1133,In_1594);
and U1119 (N_1119,In_2565,In_2566);
nand U1120 (N_1120,In_168,In_2247);
or U1121 (N_1121,In_2739,In_2646);
nand U1122 (N_1122,In_2787,In_1187);
and U1123 (N_1123,In_742,In_1350);
nor U1124 (N_1124,In_851,In_1264);
nand U1125 (N_1125,In_1720,In_185);
nand U1126 (N_1126,In_1878,In_253);
or U1127 (N_1127,In_2242,In_473);
xnor U1128 (N_1128,In_2081,In_1970);
nand U1129 (N_1129,In_919,In_991);
or U1130 (N_1130,In_685,In_2270);
nand U1131 (N_1131,In_1699,In_1174);
and U1132 (N_1132,In_2008,In_1663);
or U1133 (N_1133,In_1079,In_514);
nor U1134 (N_1134,In_2424,In_2612);
nand U1135 (N_1135,In_979,In_476);
xnor U1136 (N_1136,In_870,In_1824);
or U1137 (N_1137,In_153,In_1448);
nor U1138 (N_1138,In_2943,In_2488);
xor U1139 (N_1139,In_1451,In_2253);
nor U1140 (N_1140,In_215,In_2535);
nor U1141 (N_1141,In_2169,In_1443);
or U1142 (N_1142,In_2466,In_2120);
nor U1143 (N_1143,In_2437,In_511);
or U1144 (N_1144,In_462,In_805);
nand U1145 (N_1145,In_803,In_1066);
or U1146 (N_1146,In_2312,In_1713);
nand U1147 (N_1147,In_1111,In_2877);
xnor U1148 (N_1148,In_2902,In_2587);
nor U1149 (N_1149,In_966,In_2340);
nor U1150 (N_1150,In_1338,In_1047);
nand U1151 (N_1151,In_2991,In_779);
xor U1152 (N_1152,In_2031,In_1968);
nor U1153 (N_1153,In_1453,In_1184);
or U1154 (N_1154,In_2701,In_2430);
and U1155 (N_1155,In_2632,In_2003);
or U1156 (N_1156,In_1396,In_127);
xnor U1157 (N_1157,In_2329,In_2336);
nand U1158 (N_1158,In_524,In_2719);
nor U1159 (N_1159,In_1012,In_2208);
or U1160 (N_1160,In_2231,In_2291);
nand U1161 (N_1161,In_1142,In_1574);
nand U1162 (N_1162,In_1198,In_2030);
and U1163 (N_1163,In_711,In_2649);
and U1164 (N_1164,In_362,In_824);
nand U1165 (N_1165,In_2856,In_1168);
and U1166 (N_1166,In_1899,In_1643);
nor U1167 (N_1167,In_91,In_907);
nand U1168 (N_1168,In_2769,In_2728);
nand U1169 (N_1169,In_2758,In_1604);
or U1170 (N_1170,In_1247,In_1603);
or U1171 (N_1171,In_884,In_2855);
nor U1172 (N_1172,In_2770,In_707);
xor U1173 (N_1173,In_2662,In_198);
nor U1174 (N_1174,In_1398,In_370);
nand U1175 (N_1175,In_333,In_1724);
and U1176 (N_1176,In_703,In_2711);
and U1177 (N_1177,In_2537,In_2258);
nand U1178 (N_1178,In_1170,In_1818);
nor U1179 (N_1179,In_2689,In_895);
nor U1180 (N_1180,In_836,In_2017);
xor U1181 (N_1181,In_708,In_930);
nor U1182 (N_1182,In_1887,In_262);
or U1183 (N_1183,In_1048,In_1282);
nand U1184 (N_1184,In_2713,In_2695);
nor U1185 (N_1185,In_2355,In_131);
nand U1186 (N_1186,In_2814,In_2806);
nand U1187 (N_1187,In_1321,In_2836);
or U1188 (N_1188,In_1528,In_1199);
nand U1189 (N_1189,In_2580,In_2729);
xnor U1190 (N_1190,In_996,In_369);
nand U1191 (N_1191,In_1736,In_2725);
or U1192 (N_1192,In_2987,In_2820);
or U1193 (N_1193,In_2214,In_2839);
xor U1194 (N_1194,In_1762,In_2871);
nand U1195 (N_1195,In_2717,In_74);
or U1196 (N_1196,In_1948,In_294);
or U1197 (N_1197,In_2609,In_2332);
nor U1198 (N_1198,In_1600,In_344);
or U1199 (N_1199,In_995,In_1284);
and U1200 (N_1200,In_624,In_2111);
nand U1201 (N_1201,In_968,In_1715);
xnor U1202 (N_1202,In_1367,In_649);
and U1203 (N_1203,In_289,In_1778);
nor U1204 (N_1204,In_2554,In_1165);
or U1205 (N_1205,In_412,In_14);
and U1206 (N_1206,In_533,In_2210);
and U1207 (N_1207,In_248,In_2549);
nand U1208 (N_1208,In_1377,In_777);
and U1209 (N_1209,In_1627,In_2552);
nand U1210 (N_1210,In_2428,In_2207);
or U1211 (N_1211,In_388,In_413);
or U1212 (N_1212,In_572,In_605);
nor U1213 (N_1213,In_1952,In_971);
nor U1214 (N_1214,In_2256,In_18);
nor U1215 (N_1215,In_2051,In_689);
nor U1216 (N_1216,In_1659,In_2569);
or U1217 (N_1217,In_983,In_1285);
or U1218 (N_1218,In_2373,In_837);
or U1219 (N_1219,In_1684,In_2821);
nor U1220 (N_1220,In_2517,In_2865);
nor U1221 (N_1221,In_2761,In_2996);
nor U1222 (N_1222,In_406,In_1906);
or U1223 (N_1223,In_125,In_559);
nor U1224 (N_1224,In_327,In_1343);
or U1225 (N_1225,In_948,In_465);
nand U1226 (N_1226,In_698,In_2173);
nand U1227 (N_1227,In_2878,In_341);
nand U1228 (N_1228,In_2219,In_565);
and U1229 (N_1229,In_1677,In_2463);
or U1230 (N_1230,In_1653,In_908);
nor U1231 (N_1231,In_1309,In_1743);
nand U1232 (N_1232,In_1522,In_901);
nor U1233 (N_1233,In_751,In_1423);
xnor U1234 (N_1234,In_787,In_2953);
nand U1235 (N_1235,In_2919,In_1541);
nor U1236 (N_1236,In_1084,In_2838);
and U1237 (N_1237,In_112,In_340);
nand U1238 (N_1238,In_2494,In_360);
and U1239 (N_1239,In_2677,In_2548);
nand U1240 (N_1240,In_1571,In_255);
and U1241 (N_1241,In_1987,In_755);
nand U1242 (N_1242,In_450,In_2320);
nand U1243 (N_1243,In_1695,In_2604);
and U1244 (N_1244,In_486,In_239);
and U1245 (N_1245,In_896,In_927);
nand U1246 (N_1246,In_2152,In_2947);
nand U1247 (N_1247,In_1053,In_1637);
nand U1248 (N_1248,In_1143,In_2233);
and U1249 (N_1249,In_366,In_401);
or U1250 (N_1250,In_2059,In_1356);
and U1251 (N_1251,In_677,In_507);
nand U1252 (N_1252,In_2276,In_2025);
and U1253 (N_1253,In_391,In_1106);
or U1254 (N_1254,In_963,In_319);
nand U1255 (N_1255,In_2861,In_2707);
nand U1256 (N_1256,In_726,In_2731);
and U1257 (N_1257,In_1188,In_560);
nor U1258 (N_1258,In_128,In_2801);
nor U1259 (N_1259,In_1103,In_550);
nor U1260 (N_1260,In_655,In_658);
or U1261 (N_1261,In_2606,In_1904);
or U1262 (N_1262,In_1826,In_356);
or U1263 (N_1263,In_2193,In_2099);
nand U1264 (N_1264,In_2376,In_2767);
nor U1265 (N_1265,In_2845,In_324);
and U1266 (N_1266,In_1233,In_193);
xnor U1267 (N_1267,In_577,In_722);
or U1268 (N_1268,In_1689,In_151);
nor U1269 (N_1269,In_1890,In_1634);
or U1270 (N_1270,In_2669,In_159);
or U1271 (N_1271,In_1822,In_867);
and U1272 (N_1272,In_395,In_37);
nand U1273 (N_1273,In_87,In_357);
or U1274 (N_1274,In_1767,In_433);
or U1275 (N_1275,In_1372,In_444);
xnor U1276 (N_1276,In_1612,In_247);
xnor U1277 (N_1277,In_2696,In_2154);
and U1278 (N_1278,In_350,In_2364);
and U1279 (N_1279,In_2971,In_696);
nand U1280 (N_1280,In_1543,In_2035);
nand U1281 (N_1281,In_1436,In_2325);
or U1282 (N_1282,In_2391,In_346);
nor U1283 (N_1283,In_881,In_2759);
nor U1284 (N_1284,In_320,In_2581);
xor U1285 (N_1285,In_2375,In_1831);
nand U1286 (N_1286,In_380,In_367);
nor U1287 (N_1287,In_213,In_2631);
or U1288 (N_1288,In_704,In_2967);
nor U1289 (N_1289,In_1703,In_2105);
nand U1290 (N_1290,In_283,In_1868);
or U1291 (N_1291,In_776,In_764);
or U1292 (N_1292,In_2848,In_2515);
and U1293 (N_1293,In_2442,In_686);
or U1294 (N_1294,In_1732,In_598);
or U1295 (N_1295,In_1041,In_76);
nand U1296 (N_1296,In_530,In_120);
nand U1297 (N_1297,In_1515,In_935);
xnor U1298 (N_1298,In_2641,In_2363);
and U1299 (N_1299,In_2614,In_431);
nand U1300 (N_1300,In_1602,In_2743);
and U1301 (N_1301,In_2138,In_1764);
and U1302 (N_1302,In_1924,In_2444);
xnor U1303 (N_1303,In_2962,In_1475);
nor U1304 (N_1304,In_1244,In_693);
xor U1305 (N_1305,In_2144,In_809);
and U1306 (N_1306,In_67,In_2513);
nand U1307 (N_1307,In_2629,In_2022);
nor U1308 (N_1308,In_2339,In_1839);
or U1309 (N_1309,In_1226,In_978);
xor U1310 (N_1310,In_679,In_2292);
and U1311 (N_1311,In_1340,In_1197);
nand U1312 (N_1312,In_1598,In_482);
nor U1313 (N_1313,In_2192,In_1105);
nor U1314 (N_1314,In_1711,In_1599);
or U1315 (N_1315,In_400,In_275);
and U1316 (N_1316,In_1412,In_1914);
xor U1317 (N_1317,In_1738,In_2348);
nor U1318 (N_1318,In_1179,In_1520);
nand U1319 (N_1319,In_2485,In_738);
and U1320 (N_1320,In_43,In_582);
or U1321 (N_1321,In_1754,In_414);
and U1322 (N_1322,In_167,In_1260);
and U1323 (N_1323,In_744,In_1705);
nand U1324 (N_1324,In_2969,In_154);
and U1325 (N_1325,In_536,In_352);
or U1326 (N_1326,In_652,In_149);
or U1327 (N_1327,In_2042,In_2422);
xnor U1328 (N_1328,In_1752,In_314);
nor U1329 (N_1329,In_335,In_1191);
and U1330 (N_1330,In_2147,In_1273);
nor U1331 (N_1331,In_1635,In_1023);
or U1332 (N_1332,In_1182,In_216);
and U1333 (N_1333,In_1454,In_1854);
nand U1334 (N_1334,In_2084,In_2764);
or U1335 (N_1335,In_2250,In_28);
nand U1336 (N_1336,In_2399,In_2092);
or U1337 (N_1337,In_923,In_22);
nor U1338 (N_1338,In_53,In_2682);
and U1339 (N_1339,In_1569,In_2800);
or U1340 (N_1340,In_2585,In_1001);
or U1341 (N_1341,In_2847,In_1194);
or U1342 (N_1342,In_801,In_2882);
nor U1343 (N_1343,In_2004,In_311);
nor U1344 (N_1344,In_1830,In_1329);
xnor U1345 (N_1345,In_374,In_1076);
xor U1346 (N_1346,In_2718,In_1);
nand U1347 (N_1347,In_1502,In_2504);
nand U1348 (N_1348,In_1037,In_672);
nor U1349 (N_1349,In_2924,In_1963);
nand U1350 (N_1350,In_2063,In_1751);
nor U1351 (N_1351,In_1638,In_2926);
or U1352 (N_1352,In_629,In_555);
nor U1353 (N_1353,In_2754,In_1656);
nor U1354 (N_1354,In_1786,In_2187);
nor U1355 (N_1355,In_1009,In_2033);
nand U1356 (N_1356,In_503,In_75);
nand U1357 (N_1357,In_124,In_2623);
nand U1358 (N_1358,In_2750,In_2546);
or U1359 (N_1359,In_2898,In_1559);
nand U1360 (N_1360,In_569,In_2741);
or U1361 (N_1361,In_1918,In_95);
nand U1362 (N_1362,In_2141,In_667);
or U1363 (N_1363,In_1347,In_182);
xnor U1364 (N_1364,In_273,In_2823);
or U1365 (N_1365,In_2683,In_2271);
nor U1366 (N_1366,In_2989,In_699);
nor U1367 (N_1367,In_1487,In_500);
nor U1368 (N_1368,In_1898,In_2828);
and U1369 (N_1369,In_345,In_166);
nand U1370 (N_1370,In_1984,In_2034);
and U1371 (N_1371,In_970,In_455);
and U1372 (N_1372,In_2116,In_611);
and U1373 (N_1373,In_2613,In_1141);
nand U1374 (N_1374,In_2912,In_599);
or U1375 (N_1375,In_1162,In_2045);
and U1376 (N_1376,In_355,In_1880);
or U1377 (N_1377,In_2940,In_1488);
or U1378 (N_1378,In_1841,In_1462);
nor U1379 (N_1379,In_656,In_2226);
nand U1380 (N_1380,In_2740,In_2279);
nor U1381 (N_1381,In_2564,In_410);
xor U1382 (N_1382,In_1867,In_606);
and U1383 (N_1383,In_259,In_2455);
or U1384 (N_1384,In_495,In_1765);
or U1385 (N_1385,In_797,In_2335);
xor U1386 (N_1386,In_285,In_2209);
nor U1387 (N_1387,In_2598,In_2261);
nor U1388 (N_1388,In_2426,In_676);
nand U1389 (N_1389,In_1923,In_1342);
and U1390 (N_1390,In_254,In_490);
and U1391 (N_1391,In_86,In_1850);
nor U1392 (N_1392,In_1929,In_2014);
or U1393 (N_1393,In_2605,In_101);
nor U1394 (N_1394,In_284,In_2476);
nand U1395 (N_1395,In_1082,In_1516);
or U1396 (N_1396,In_1438,In_2243);
or U1397 (N_1397,In_59,In_491);
or U1398 (N_1398,In_2992,In_1799);
or U1399 (N_1399,In_2655,In_1658);
and U1400 (N_1400,In_853,In_508);
nand U1401 (N_1401,In_1096,In_300);
nor U1402 (N_1402,In_1957,In_786);
nor U1403 (N_1403,In_839,In_2688);
nor U1404 (N_1404,In_775,In_1214);
nor U1405 (N_1405,In_609,In_592);
nor U1406 (N_1406,In_1570,In_1312);
nand U1407 (N_1407,In_2639,In_2785);
or U1408 (N_1408,In_729,In_235);
nand U1409 (N_1409,In_1595,In_2281);
xnor U1410 (N_1410,In_730,In_224);
nand U1411 (N_1411,In_85,In_1080);
nand U1412 (N_1412,In_2680,In_1862);
or U1413 (N_1413,In_1768,In_939);
and U1414 (N_1414,In_1714,In_1437);
nor U1415 (N_1415,In_2178,In_2573);
nand U1416 (N_1416,In_398,In_2337);
nand U1417 (N_1417,In_603,In_1727);
nor U1418 (N_1418,In_581,In_1568);
nor U1419 (N_1419,In_2412,In_81);
or U1420 (N_1420,In_436,In_469);
nor U1421 (N_1421,In_537,In_1530);
or U1422 (N_1422,In_1028,In_2125);
or U1423 (N_1423,In_1989,In_2408);
xor U1424 (N_1424,In_856,In_468);
xnor U1425 (N_1425,In_1419,In_42);
and U1426 (N_1426,In_1208,In_1964);
nor U1427 (N_1427,In_121,In_504);
or U1428 (N_1428,In_2525,In_2263);
and U1429 (N_1429,In_1277,In_1067);
or U1430 (N_1430,In_989,In_2289);
or U1431 (N_1431,In_1757,In_1742);
nor U1432 (N_1432,In_1945,In_2300);
or U1433 (N_1433,In_1655,In_1095);
and U1434 (N_1434,In_1204,In_2137);
or U1435 (N_1435,In_2896,In_2705);
nand U1436 (N_1436,In_175,In_823);
or U1437 (N_1437,In_2388,In_1846);
nor U1438 (N_1438,In_260,In_2881);
or U1439 (N_1439,In_631,In_820);
nand U1440 (N_1440,In_2186,In_2903);
nand U1441 (N_1441,In_2368,In_1307);
nor U1442 (N_1442,In_2433,In_1671);
nor U1443 (N_1443,In_1988,In_263);
nand U1444 (N_1444,In_1716,In_736);
and U1445 (N_1445,In_1788,In_1375);
nand U1446 (N_1446,In_1077,In_2206);
or U1447 (N_1447,In_833,In_2607);
nand U1448 (N_1448,In_2230,In_1269);
or U1449 (N_1449,In_1920,In_1033);
nand U1450 (N_1450,In_2858,In_715);
or U1451 (N_1451,In_2135,In_1302);
or U1452 (N_1452,In_2400,In_384);
nand U1453 (N_1453,In_1524,In_1006);
or U1454 (N_1454,In_339,In_1330);
xor U1455 (N_1455,In_1109,In_875);
nand U1456 (N_1456,In_116,In_1150);
or U1457 (N_1457,In_2009,In_1513);
or U1458 (N_1458,In_758,In_1798);
nor U1459 (N_1459,In_1777,In_2440);
nand U1460 (N_1460,In_448,In_2970);
and U1461 (N_1461,In_2393,In_173);
nor U1462 (N_1462,In_1094,In_20);
xnor U1463 (N_1463,In_1126,In_1669);
or U1464 (N_1464,In_2776,In_2538);
or U1465 (N_1465,In_2826,In_810);
nand U1466 (N_1466,In_2469,In_449);
nand U1467 (N_1467,In_1921,In_2297);
and U1468 (N_1468,In_780,In_2010);
nor U1469 (N_1469,In_1647,In_2768);
and U1470 (N_1470,In_644,In_1886);
nor U1471 (N_1471,In_70,In_2901);
nor U1472 (N_1472,In_334,In_342);
and U1473 (N_1473,In_2019,In_564);
nand U1474 (N_1474,In_135,In_434);
or U1475 (N_1475,In_754,In_1835);
xnor U1476 (N_1476,In_2757,In_397);
nor U1477 (N_1477,In_877,In_2315);
xor U1478 (N_1478,In_2459,In_1100);
and U1479 (N_1479,In_295,In_133);
or U1480 (N_1480,In_378,In_2298);
nand U1481 (N_1481,In_2089,In_171);
nor U1482 (N_1482,In_2257,In_165);
or U1483 (N_1483,In_917,In_846);
nand U1484 (N_1484,In_2011,In_2275);
xnor U1485 (N_1485,In_2638,In_2749);
nand U1486 (N_1486,In_238,In_72);
nor U1487 (N_1487,In_487,In_217);
nor U1488 (N_1488,In_2305,In_540);
nand U1489 (N_1489,In_2079,In_276);
and U1490 (N_1490,In_2262,In_2425);
and U1491 (N_1491,In_443,In_2699);
xor U1492 (N_1492,In_1995,In_1014);
nand U1493 (N_1493,In_774,In_2361);
nand U1494 (N_1494,In_2570,In_767);
or U1495 (N_1495,In_1548,In_26);
and U1496 (N_1496,In_911,In_1004);
or U1497 (N_1497,In_1238,In_169);
or U1498 (N_1498,In_1857,In_2457);
or U1499 (N_1499,In_778,In_549);
nor U1500 (N_1500,In_1690,In_364);
or U1501 (N_1501,In_640,In_754);
or U1502 (N_1502,In_1700,In_2409);
nor U1503 (N_1503,In_1300,In_33);
or U1504 (N_1504,In_1125,In_2065);
nor U1505 (N_1505,In_1754,In_2590);
nand U1506 (N_1506,In_1378,In_2449);
and U1507 (N_1507,In_2635,In_595);
nand U1508 (N_1508,In_1074,In_2847);
nor U1509 (N_1509,In_2508,In_2837);
or U1510 (N_1510,In_416,In_2764);
or U1511 (N_1511,In_2218,In_2087);
or U1512 (N_1512,In_1524,In_998);
nand U1513 (N_1513,In_588,In_1224);
xor U1514 (N_1514,In_2344,In_587);
and U1515 (N_1515,In_658,In_593);
nand U1516 (N_1516,In_2119,In_130);
nor U1517 (N_1517,In_1367,In_1692);
or U1518 (N_1518,In_2434,In_1216);
and U1519 (N_1519,In_2241,In_2192);
and U1520 (N_1520,In_2156,In_252);
nand U1521 (N_1521,In_2257,In_446);
nand U1522 (N_1522,In_758,In_2701);
nor U1523 (N_1523,In_89,In_2738);
or U1524 (N_1524,In_2102,In_1826);
nand U1525 (N_1525,In_237,In_2716);
nand U1526 (N_1526,In_1995,In_1299);
or U1527 (N_1527,In_2042,In_2019);
and U1528 (N_1528,In_247,In_2206);
and U1529 (N_1529,In_647,In_2652);
or U1530 (N_1530,In_74,In_1131);
nor U1531 (N_1531,In_1130,In_2107);
and U1532 (N_1532,In_2756,In_891);
and U1533 (N_1533,In_808,In_1107);
nor U1534 (N_1534,In_2330,In_324);
or U1535 (N_1535,In_2597,In_410);
and U1536 (N_1536,In_1670,In_921);
and U1537 (N_1537,In_418,In_1256);
xnor U1538 (N_1538,In_465,In_2267);
nor U1539 (N_1539,In_2583,In_692);
nor U1540 (N_1540,In_1387,In_2472);
or U1541 (N_1541,In_1392,In_1245);
or U1542 (N_1542,In_1187,In_2687);
and U1543 (N_1543,In_2983,In_1543);
nor U1544 (N_1544,In_1733,In_2996);
or U1545 (N_1545,In_555,In_2173);
and U1546 (N_1546,In_1813,In_894);
or U1547 (N_1547,In_2605,In_2604);
or U1548 (N_1548,In_1353,In_726);
xor U1549 (N_1549,In_1804,In_1961);
and U1550 (N_1550,In_1795,In_2382);
and U1551 (N_1551,In_2593,In_342);
nor U1552 (N_1552,In_2315,In_1373);
nor U1553 (N_1553,In_267,In_2494);
nand U1554 (N_1554,In_1584,In_1446);
nor U1555 (N_1555,In_2424,In_1512);
nor U1556 (N_1556,In_1421,In_978);
nand U1557 (N_1557,In_692,In_740);
nand U1558 (N_1558,In_965,In_669);
nand U1559 (N_1559,In_1595,In_2832);
or U1560 (N_1560,In_2646,In_2308);
nand U1561 (N_1561,In_372,In_2627);
and U1562 (N_1562,In_1051,In_825);
xnor U1563 (N_1563,In_2323,In_64);
xnor U1564 (N_1564,In_958,In_466);
and U1565 (N_1565,In_173,In_2083);
or U1566 (N_1566,In_1807,In_18);
nand U1567 (N_1567,In_968,In_2302);
nand U1568 (N_1568,In_2236,In_2184);
and U1569 (N_1569,In_2537,In_912);
and U1570 (N_1570,In_2439,In_2559);
xor U1571 (N_1571,In_1713,In_1003);
nand U1572 (N_1572,In_496,In_1134);
or U1573 (N_1573,In_1606,In_1412);
nor U1574 (N_1574,In_2801,In_2852);
or U1575 (N_1575,In_1786,In_2864);
nand U1576 (N_1576,In_2920,In_2665);
xor U1577 (N_1577,In_1035,In_2718);
xnor U1578 (N_1578,In_1167,In_657);
xnor U1579 (N_1579,In_1232,In_2901);
nand U1580 (N_1580,In_1354,In_777);
and U1581 (N_1581,In_2073,In_307);
or U1582 (N_1582,In_502,In_603);
nand U1583 (N_1583,In_1013,In_805);
and U1584 (N_1584,In_114,In_1089);
and U1585 (N_1585,In_2325,In_852);
xnor U1586 (N_1586,In_283,In_2201);
and U1587 (N_1587,In_1371,In_2030);
or U1588 (N_1588,In_1146,In_1858);
and U1589 (N_1589,In_161,In_299);
nand U1590 (N_1590,In_322,In_2149);
nor U1591 (N_1591,In_27,In_1834);
nand U1592 (N_1592,In_161,In_363);
and U1593 (N_1593,In_1422,In_1940);
or U1594 (N_1594,In_2927,In_879);
nand U1595 (N_1595,In_1649,In_1391);
nand U1596 (N_1596,In_1685,In_2644);
nor U1597 (N_1597,In_922,In_1017);
or U1598 (N_1598,In_1106,In_828);
nand U1599 (N_1599,In_2386,In_2199);
and U1600 (N_1600,In_1966,In_1720);
and U1601 (N_1601,In_1394,In_1740);
xnor U1602 (N_1602,In_1883,In_612);
nor U1603 (N_1603,In_2778,In_1422);
or U1604 (N_1604,In_1291,In_685);
nor U1605 (N_1605,In_2666,In_676);
nor U1606 (N_1606,In_1083,In_199);
nand U1607 (N_1607,In_2874,In_2728);
and U1608 (N_1608,In_1839,In_2076);
nand U1609 (N_1609,In_79,In_2544);
or U1610 (N_1610,In_2673,In_1132);
nor U1611 (N_1611,In_357,In_2181);
nand U1612 (N_1612,In_836,In_1675);
and U1613 (N_1613,In_63,In_77);
xor U1614 (N_1614,In_2727,In_731);
and U1615 (N_1615,In_1256,In_2515);
nand U1616 (N_1616,In_458,In_2517);
nor U1617 (N_1617,In_1710,In_2973);
or U1618 (N_1618,In_2102,In_2520);
nand U1619 (N_1619,In_345,In_1244);
or U1620 (N_1620,In_2262,In_2869);
nand U1621 (N_1621,In_340,In_2208);
or U1622 (N_1622,In_712,In_2649);
nand U1623 (N_1623,In_2166,In_296);
or U1624 (N_1624,In_2497,In_2324);
nor U1625 (N_1625,In_2821,In_1394);
xnor U1626 (N_1626,In_2170,In_374);
nand U1627 (N_1627,In_1870,In_343);
nor U1628 (N_1628,In_685,In_405);
nand U1629 (N_1629,In_2032,In_951);
and U1630 (N_1630,In_73,In_2160);
and U1631 (N_1631,In_2445,In_25);
or U1632 (N_1632,In_804,In_1785);
nor U1633 (N_1633,In_1939,In_1212);
xnor U1634 (N_1634,In_1976,In_2198);
and U1635 (N_1635,In_1262,In_1453);
nor U1636 (N_1636,In_444,In_2867);
nor U1637 (N_1637,In_461,In_143);
and U1638 (N_1638,In_2133,In_1884);
or U1639 (N_1639,In_251,In_1258);
nor U1640 (N_1640,In_211,In_2724);
and U1641 (N_1641,In_853,In_1034);
nand U1642 (N_1642,In_1804,In_2672);
nand U1643 (N_1643,In_32,In_828);
and U1644 (N_1644,In_702,In_1918);
nor U1645 (N_1645,In_42,In_1460);
or U1646 (N_1646,In_1618,In_2515);
or U1647 (N_1647,In_2948,In_1267);
nor U1648 (N_1648,In_1948,In_57);
or U1649 (N_1649,In_1675,In_2889);
nand U1650 (N_1650,In_1686,In_2943);
and U1651 (N_1651,In_1461,In_2015);
and U1652 (N_1652,In_2313,In_1416);
nor U1653 (N_1653,In_2378,In_312);
nor U1654 (N_1654,In_2507,In_223);
or U1655 (N_1655,In_2654,In_1414);
nand U1656 (N_1656,In_1750,In_1662);
and U1657 (N_1657,In_413,In_2151);
or U1658 (N_1658,In_915,In_2712);
xnor U1659 (N_1659,In_1311,In_1676);
and U1660 (N_1660,In_1923,In_2546);
and U1661 (N_1661,In_1732,In_2521);
nand U1662 (N_1662,In_1968,In_2473);
nand U1663 (N_1663,In_2969,In_2325);
nand U1664 (N_1664,In_531,In_1817);
or U1665 (N_1665,In_1203,In_1081);
nand U1666 (N_1666,In_287,In_1242);
or U1667 (N_1667,In_1264,In_1254);
or U1668 (N_1668,In_587,In_1720);
nand U1669 (N_1669,In_656,In_2703);
xnor U1670 (N_1670,In_970,In_1701);
xor U1671 (N_1671,In_2482,In_837);
and U1672 (N_1672,In_2956,In_689);
and U1673 (N_1673,In_2663,In_278);
xnor U1674 (N_1674,In_1612,In_1686);
nand U1675 (N_1675,In_102,In_1427);
nand U1676 (N_1676,In_2668,In_167);
xor U1677 (N_1677,In_1478,In_287);
and U1678 (N_1678,In_832,In_1830);
and U1679 (N_1679,In_2654,In_1959);
nor U1680 (N_1680,In_1398,In_2957);
nand U1681 (N_1681,In_2247,In_2206);
xor U1682 (N_1682,In_1619,In_1454);
nand U1683 (N_1683,In_1265,In_1966);
nor U1684 (N_1684,In_945,In_1303);
nor U1685 (N_1685,In_2991,In_1229);
nand U1686 (N_1686,In_2085,In_2749);
and U1687 (N_1687,In_2342,In_1983);
nand U1688 (N_1688,In_2002,In_2617);
nand U1689 (N_1689,In_1433,In_626);
and U1690 (N_1690,In_2310,In_122);
nand U1691 (N_1691,In_832,In_2072);
nand U1692 (N_1692,In_2642,In_263);
nor U1693 (N_1693,In_81,In_429);
or U1694 (N_1694,In_2082,In_2614);
xnor U1695 (N_1695,In_2978,In_841);
or U1696 (N_1696,In_2487,In_2615);
or U1697 (N_1697,In_606,In_1214);
nor U1698 (N_1698,In_548,In_1906);
nand U1699 (N_1699,In_2827,In_1865);
nand U1700 (N_1700,In_2243,In_1818);
nor U1701 (N_1701,In_2422,In_2760);
nand U1702 (N_1702,In_101,In_463);
and U1703 (N_1703,In_1861,In_342);
nand U1704 (N_1704,In_691,In_1020);
and U1705 (N_1705,In_560,In_1648);
nor U1706 (N_1706,In_1496,In_397);
or U1707 (N_1707,In_2364,In_2138);
nand U1708 (N_1708,In_1190,In_2285);
and U1709 (N_1709,In_726,In_924);
or U1710 (N_1710,In_520,In_1448);
and U1711 (N_1711,In_2713,In_565);
xor U1712 (N_1712,In_2718,In_570);
xor U1713 (N_1713,In_1785,In_1230);
xor U1714 (N_1714,In_379,In_2450);
nand U1715 (N_1715,In_1087,In_1884);
nor U1716 (N_1716,In_1172,In_1685);
and U1717 (N_1717,In_346,In_2056);
nor U1718 (N_1718,In_2263,In_2194);
and U1719 (N_1719,In_845,In_1222);
and U1720 (N_1720,In_2574,In_701);
and U1721 (N_1721,In_1460,In_1178);
nor U1722 (N_1722,In_1587,In_2796);
nand U1723 (N_1723,In_1073,In_2999);
nand U1724 (N_1724,In_695,In_2553);
nor U1725 (N_1725,In_1372,In_2188);
nor U1726 (N_1726,In_919,In_2293);
and U1727 (N_1727,In_1295,In_1392);
and U1728 (N_1728,In_2334,In_1874);
nand U1729 (N_1729,In_945,In_52);
nor U1730 (N_1730,In_393,In_2942);
nor U1731 (N_1731,In_1624,In_2115);
nor U1732 (N_1732,In_1809,In_2756);
nand U1733 (N_1733,In_2021,In_792);
nor U1734 (N_1734,In_1736,In_1155);
and U1735 (N_1735,In_169,In_1968);
nor U1736 (N_1736,In_1990,In_2634);
nand U1737 (N_1737,In_1649,In_1699);
or U1738 (N_1738,In_1114,In_196);
nand U1739 (N_1739,In_2080,In_940);
nor U1740 (N_1740,In_1971,In_1988);
nand U1741 (N_1741,In_649,In_1253);
or U1742 (N_1742,In_1841,In_1086);
and U1743 (N_1743,In_1099,In_1483);
and U1744 (N_1744,In_445,In_1429);
nand U1745 (N_1745,In_768,In_2958);
and U1746 (N_1746,In_2779,In_994);
and U1747 (N_1747,In_1390,In_1397);
or U1748 (N_1748,In_1065,In_2703);
and U1749 (N_1749,In_2407,In_781);
and U1750 (N_1750,In_1552,In_2792);
and U1751 (N_1751,In_2899,In_1651);
nor U1752 (N_1752,In_2958,In_382);
and U1753 (N_1753,In_431,In_2672);
or U1754 (N_1754,In_729,In_2311);
or U1755 (N_1755,In_2500,In_187);
nand U1756 (N_1756,In_409,In_1227);
nand U1757 (N_1757,In_2770,In_2625);
or U1758 (N_1758,In_572,In_2146);
nor U1759 (N_1759,In_622,In_2417);
or U1760 (N_1760,In_831,In_76);
nor U1761 (N_1761,In_1642,In_1919);
or U1762 (N_1762,In_1609,In_589);
nand U1763 (N_1763,In_1210,In_1448);
or U1764 (N_1764,In_1880,In_2823);
or U1765 (N_1765,In_61,In_1485);
nand U1766 (N_1766,In_2402,In_1489);
xor U1767 (N_1767,In_970,In_598);
nor U1768 (N_1768,In_397,In_2277);
nor U1769 (N_1769,In_2859,In_2688);
or U1770 (N_1770,In_673,In_1961);
nand U1771 (N_1771,In_219,In_117);
or U1772 (N_1772,In_556,In_1305);
and U1773 (N_1773,In_1272,In_189);
xnor U1774 (N_1774,In_1411,In_2060);
and U1775 (N_1775,In_2898,In_1760);
nor U1776 (N_1776,In_2031,In_1155);
nand U1777 (N_1777,In_1614,In_1890);
and U1778 (N_1778,In_1067,In_1648);
nor U1779 (N_1779,In_838,In_57);
nor U1780 (N_1780,In_1615,In_1665);
nor U1781 (N_1781,In_1859,In_1428);
nand U1782 (N_1782,In_2992,In_1043);
and U1783 (N_1783,In_1293,In_2517);
nor U1784 (N_1784,In_932,In_804);
xnor U1785 (N_1785,In_993,In_843);
xnor U1786 (N_1786,In_2009,In_2463);
or U1787 (N_1787,In_1289,In_204);
and U1788 (N_1788,In_1263,In_308);
and U1789 (N_1789,In_1671,In_1894);
or U1790 (N_1790,In_623,In_2576);
nor U1791 (N_1791,In_2132,In_102);
nand U1792 (N_1792,In_2319,In_1878);
and U1793 (N_1793,In_645,In_1320);
nand U1794 (N_1794,In_1692,In_858);
nor U1795 (N_1795,In_1966,In_2376);
or U1796 (N_1796,In_2580,In_974);
or U1797 (N_1797,In_1455,In_1673);
nor U1798 (N_1798,In_212,In_2186);
or U1799 (N_1799,In_1944,In_1841);
nand U1800 (N_1800,In_2186,In_1397);
nand U1801 (N_1801,In_353,In_719);
nand U1802 (N_1802,In_1392,In_2638);
nor U1803 (N_1803,In_1196,In_2913);
nand U1804 (N_1804,In_2178,In_2723);
or U1805 (N_1805,In_2405,In_827);
nor U1806 (N_1806,In_428,In_362);
nand U1807 (N_1807,In_522,In_2477);
and U1808 (N_1808,In_177,In_2581);
xnor U1809 (N_1809,In_2386,In_1950);
or U1810 (N_1810,In_609,In_393);
and U1811 (N_1811,In_758,In_306);
xor U1812 (N_1812,In_2295,In_2346);
nand U1813 (N_1813,In_2079,In_2741);
xor U1814 (N_1814,In_788,In_579);
nor U1815 (N_1815,In_2502,In_1924);
nand U1816 (N_1816,In_270,In_1279);
or U1817 (N_1817,In_2560,In_1286);
nand U1818 (N_1818,In_615,In_1657);
or U1819 (N_1819,In_902,In_2552);
xor U1820 (N_1820,In_1332,In_2752);
xnor U1821 (N_1821,In_1976,In_712);
or U1822 (N_1822,In_1906,In_1586);
nor U1823 (N_1823,In_679,In_1996);
nand U1824 (N_1824,In_911,In_1667);
nand U1825 (N_1825,In_2883,In_1035);
nand U1826 (N_1826,In_1239,In_2944);
nor U1827 (N_1827,In_1905,In_484);
or U1828 (N_1828,In_2204,In_2164);
or U1829 (N_1829,In_2771,In_432);
nand U1830 (N_1830,In_2600,In_2016);
or U1831 (N_1831,In_925,In_1353);
nor U1832 (N_1832,In_1900,In_1485);
nor U1833 (N_1833,In_694,In_514);
nor U1834 (N_1834,In_1624,In_2881);
or U1835 (N_1835,In_1065,In_2527);
xor U1836 (N_1836,In_2987,In_695);
nand U1837 (N_1837,In_1273,In_2694);
nand U1838 (N_1838,In_2973,In_415);
nand U1839 (N_1839,In_2496,In_2095);
and U1840 (N_1840,In_2965,In_725);
or U1841 (N_1841,In_365,In_1438);
nor U1842 (N_1842,In_58,In_829);
or U1843 (N_1843,In_300,In_936);
nand U1844 (N_1844,In_443,In_2879);
and U1845 (N_1845,In_1446,In_518);
or U1846 (N_1846,In_774,In_2777);
nor U1847 (N_1847,In_2736,In_228);
nor U1848 (N_1848,In_1769,In_807);
xor U1849 (N_1849,In_1706,In_1822);
and U1850 (N_1850,In_252,In_2287);
nor U1851 (N_1851,In_404,In_2442);
nand U1852 (N_1852,In_993,In_2720);
xor U1853 (N_1853,In_2478,In_2852);
or U1854 (N_1854,In_2794,In_943);
or U1855 (N_1855,In_116,In_2060);
or U1856 (N_1856,In_1081,In_1753);
nor U1857 (N_1857,In_778,In_345);
and U1858 (N_1858,In_581,In_1395);
nor U1859 (N_1859,In_1402,In_2589);
and U1860 (N_1860,In_1341,In_2029);
nor U1861 (N_1861,In_1117,In_2539);
and U1862 (N_1862,In_2820,In_1606);
nor U1863 (N_1863,In_2510,In_2803);
or U1864 (N_1864,In_2012,In_2604);
or U1865 (N_1865,In_1712,In_789);
xnor U1866 (N_1866,In_2272,In_1610);
nor U1867 (N_1867,In_1026,In_2539);
xnor U1868 (N_1868,In_2290,In_2913);
nor U1869 (N_1869,In_2375,In_2781);
xnor U1870 (N_1870,In_1023,In_1318);
or U1871 (N_1871,In_2350,In_2201);
nand U1872 (N_1872,In_1327,In_313);
or U1873 (N_1873,In_1066,In_649);
nor U1874 (N_1874,In_1105,In_1687);
and U1875 (N_1875,In_2033,In_1080);
nor U1876 (N_1876,In_989,In_520);
nand U1877 (N_1877,In_1205,In_2384);
nor U1878 (N_1878,In_337,In_2272);
xnor U1879 (N_1879,In_204,In_411);
or U1880 (N_1880,In_1719,In_464);
nor U1881 (N_1881,In_1223,In_802);
and U1882 (N_1882,In_1441,In_1052);
nor U1883 (N_1883,In_1045,In_127);
and U1884 (N_1884,In_549,In_2758);
nand U1885 (N_1885,In_1642,In_1848);
and U1886 (N_1886,In_1649,In_12);
or U1887 (N_1887,In_942,In_1455);
xnor U1888 (N_1888,In_2904,In_2565);
nand U1889 (N_1889,In_1767,In_733);
nor U1890 (N_1890,In_1467,In_1072);
nand U1891 (N_1891,In_2337,In_2566);
nand U1892 (N_1892,In_712,In_938);
nor U1893 (N_1893,In_2459,In_575);
nand U1894 (N_1894,In_2601,In_2551);
or U1895 (N_1895,In_377,In_1505);
or U1896 (N_1896,In_1550,In_259);
nor U1897 (N_1897,In_1067,In_335);
nor U1898 (N_1898,In_1558,In_1469);
and U1899 (N_1899,In_1180,In_2087);
and U1900 (N_1900,In_2860,In_1301);
nand U1901 (N_1901,In_1251,In_2887);
and U1902 (N_1902,In_2304,In_2237);
nor U1903 (N_1903,In_2903,In_1168);
xnor U1904 (N_1904,In_1869,In_720);
or U1905 (N_1905,In_760,In_1930);
nand U1906 (N_1906,In_1063,In_2406);
xnor U1907 (N_1907,In_2922,In_2210);
or U1908 (N_1908,In_1467,In_2019);
xor U1909 (N_1909,In_344,In_2259);
nor U1910 (N_1910,In_596,In_2959);
or U1911 (N_1911,In_357,In_973);
nor U1912 (N_1912,In_1429,In_490);
nand U1913 (N_1913,In_2379,In_2756);
nor U1914 (N_1914,In_1631,In_1749);
and U1915 (N_1915,In_2626,In_1506);
nand U1916 (N_1916,In_2597,In_1313);
or U1917 (N_1917,In_2002,In_1522);
and U1918 (N_1918,In_2561,In_2766);
nand U1919 (N_1919,In_2835,In_128);
xnor U1920 (N_1920,In_1790,In_1501);
xnor U1921 (N_1921,In_1210,In_2238);
and U1922 (N_1922,In_2133,In_67);
nand U1923 (N_1923,In_570,In_1427);
or U1924 (N_1924,In_241,In_1976);
or U1925 (N_1925,In_809,In_994);
and U1926 (N_1926,In_2905,In_1889);
xor U1927 (N_1927,In_161,In_1825);
and U1928 (N_1928,In_746,In_933);
or U1929 (N_1929,In_1283,In_2772);
nand U1930 (N_1930,In_681,In_2630);
and U1931 (N_1931,In_1162,In_2713);
nor U1932 (N_1932,In_1802,In_2940);
and U1933 (N_1933,In_378,In_44);
and U1934 (N_1934,In_2378,In_1402);
and U1935 (N_1935,In_1089,In_2153);
or U1936 (N_1936,In_2633,In_298);
nor U1937 (N_1937,In_2885,In_2979);
and U1938 (N_1938,In_1914,In_373);
or U1939 (N_1939,In_1396,In_1286);
and U1940 (N_1940,In_1301,In_2380);
or U1941 (N_1941,In_676,In_652);
nor U1942 (N_1942,In_313,In_41);
or U1943 (N_1943,In_346,In_62);
nor U1944 (N_1944,In_907,In_601);
or U1945 (N_1945,In_2682,In_871);
nor U1946 (N_1946,In_655,In_1815);
and U1947 (N_1947,In_1086,In_858);
nor U1948 (N_1948,In_28,In_1615);
and U1949 (N_1949,In_2179,In_2371);
or U1950 (N_1950,In_1643,In_545);
or U1951 (N_1951,In_2542,In_2121);
xnor U1952 (N_1952,In_1312,In_2999);
and U1953 (N_1953,In_1761,In_2716);
or U1954 (N_1954,In_591,In_2465);
nand U1955 (N_1955,In_1591,In_1143);
xor U1956 (N_1956,In_2771,In_787);
or U1957 (N_1957,In_2148,In_763);
or U1958 (N_1958,In_673,In_1648);
and U1959 (N_1959,In_2588,In_648);
xnor U1960 (N_1960,In_2605,In_1813);
and U1961 (N_1961,In_97,In_1468);
and U1962 (N_1962,In_421,In_1797);
or U1963 (N_1963,In_2040,In_2902);
and U1964 (N_1964,In_2402,In_953);
or U1965 (N_1965,In_1205,In_365);
nand U1966 (N_1966,In_2612,In_2968);
and U1967 (N_1967,In_1879,In_2541);
nand U1968 (N_1968,In_1978,In_170);
or U1969 (N_1969,In_1719,In_2568);
xnor U1970 (N_1970,In_2219,In_2341);
and U1971 (N_1971,In_1152,In_180);
or U1972 (N_1972,In_2941,In_601);
or U1973 (N_1973,In_1450,In_1498);
nor U1974 (N_1974,In_1893,In_2888);
nand U1975 (N_1975,In_1737,In_2347);
or U1976 (N_1976,In_229,In_1868);
nand U1977 (N_1977,In_2231,In_1359);
or U1978 (N_1978,In_1109,In_1412);
and U1979 (N_1979,In_1089,In_2181);
and U1980 (N_1980,In_1699,In_603);
nand U1981 (N_1981,In_378,In_2598);
nand U1982 (N_1982,In_2187,In_2422);
xnor U1983 (N_1983,In_367,In_1399);
or U1984 (N_1984,In_2518,In_2899);
and U1985 (N_1985,In_1957,In_442);
nand U1986 (N_1986,In_682,In_848);
and U1987 (N_1987,In_2202,In_2966);
or U1988 (N_1988,In_1717,In_229);
or U1989 (N_1989,In_1967,In_2997);
and U1990 (N_1990,In_1981,In_2568);
or U1991 (N_1991,In_2217,In_1421);
nor U1992 (N_1992,In_2231,In_1089);
nor U1993 (N_1993,In_668,In_1515);
nor U1994 (N_1994,In_1656,In_722);
xor U1995 (N_1995,In_1155,In_2668);
nor U1996 (N_1996,In_13,In_1999);
and U1997 (N_1997,In_1866,In_2755);
nand U1998 (N_1998,In_2900,In_619);
or U1999 (N_1999,In_2513,In_1609);
nand U2000 (N_2000,In_1003,In_779);
and U2001 (N_2001,In_917,In_2538);
nand U2002 (N_2002,In_2201,In_590);
xor U2003 (N_2003,In_2995,In_1832);
nor U2004 (N_2004,In_2325,In_1017);
and U2005 (N_2005,In_24,In_297);
nor U2006 (N_2006,In_399,In_1844);
or U2007 (N_2007,In_2033,In_717);
nor U2008 (N_2008,In_627,In_2623);
xnor U2009 (N_2009,In_808,In_2090);
nor U2010 (N_2010,In_283,In_2571);
and U2011 (N_2011,In_43,In_2782);
or U2012 (N_2012,In_111,In_2089);
nand U2013 (N_2013,In_2362,In_1871);
and U2014 (N_2014,In_36,In_1612);
nand U2015 (N_2015,In_896,In_2414);
and U2016 (N_2016,In_2607,In_2148);
or U2017 (N_2017,In_2808,In_345);
and U2018 (N_2018,In_758,In_2907);
nor U2019 (N_2019,In_632,In_776);
or U2020 (N_2020,In_2917,In_2606);
or U2021 (N_2021,In_2752,In_1197);
nor U2022 (N_2022,In_2600,In_1613);
nand U2023 (N_2023,In_112,In_1925);
nand U2024 (N_2024,In_2837,In_2666);
or U2025 (N_2025,In_2230,In_971);
nor U2026 (N_2026,In_368,In_2521);
nand U2027 (N_2027,In_913,In_1403);
or U2028 (N_2028,In_2277,In_1628);
and U2029 (N_2029,In_2743,In_390);
nor U2030 (N_2030,In_1299,In_453);
nor U2031 (N_2031,In_1353,In_467);
or U2032 (N_2032,In_2002,In_970);
nor U2033 (N_2033,In_1856,In_948);
nand U2034 (N_2034,In_2582,In_808);
or U2035 (N_2035,In_1117,In_1993);
nor U2036 (N_2036,In_1447,In_1344);
nor U2037 (N_2037,In_90,In_1835);
nor U2038 (N_2038,In_1354,In_2762);
and U2039 (N_2039,In_1885,In_58);
xor U2040 (N_2040,In_225,In_2301);
or U2041 (N_2041,In_2323,In_2475);
nand U2042 (N_2042,In_210,In_1918);
and U2043 (N_2043,In_2036,In_1001);
nor U2044 (N_2044,In_2473,In_2727);
and U2045 (N_2045,In_1599,In_623);
or U2046 (N_2046,In_1914,In_1527);
nand U2047 (N_2047,In_1459,In_1515);
or U2048 (N_2048,In_2726,In_800);
nand U2049 (N_2049,In_2568,In_206);
or U2050 (N_2050,In_2387,In_452);
xnor U2051 (N_2051,In_570,In_1771);
or U2052 (N_2052,In_1245,In_1173);
or U2053 (N_2053,In_1001,In_1621);
nand U2054 (N_2054,In_1870,In_737);
nand U2055 (N_2055,In_545,In_1852);
nand U2056 (N_2056,In_2955,In_1824);
and U2057 (N_2057,In_2036,In_937);
and U2058 (N_2058,In_1455,In_818);
and U2059 (N_2059,In_855,In_691);
xnor U2060 (N_2060,In_497,In_55);
nor U2061 (N_2061,In_2280,In_1351);
and U2062 (N_2062,In_862,In_122);
nand U2063 (N_2063,In_1309,In_245);
xnor U2064 (N_2064,In_1424,In_817);
nor U2065 (N_2065,In_2039,In_589);
and U2066 (N_2066,In_1666,In_16);
nand U2067 (N_2067,In_2046,In_773);
nand U2068 (N_2068,In_2216,In_409);
or U2069 (N_2069,In_2674,In_274);
xnor U2070 (N_2070,In_2304,In_1853);
or U2071 (N_2071,In_2464,In_1307);
nand U2072 (N_2072,In_2989,In_1134);
nand U2073 (N_2073,In_611,In_383);
xor U2074 (N_2074,In_2013,In_1846);
nor U2075 (N_2075,In_1608,In_293);
nand U2076 (N_2076,In_2710,In_899);
nand U2077 (N_2077,In_2394,In_2810);
nand U2078 (N_2078,In_159,In_288);
nand U2079 (N_2079,In_1775,In_2409);
and U2080 (N_2080,In_1952,In_1608);
and U2081 (N_2081,In_675,In_2626);
nor U2082 (N_2082,In_964,In_313);
nand U2083 (N_2083,In_187,In_2823);
or U2084 (N_2084,In_2795,In_2080);
nor U2085 (N_2085,In_1667,In_567);
nor U2086 (N_2086,In_12,In_2037);
nor U2087 (N_2087,In_2047,In_1466);
nor U2088 (N_2088,In_1045,In_2727);
and U2089 (N_2089,In_1070,In_604);
nand U2090 (N_2090,In_826,In_1206);
nand U2091 (N_2091,In_211,In_2641);
xnor U2092 (N_2092,In_758,In_1392);
nor U2093 (N_2093,In_251,In_2389);
and U2094 (N_2094,In_512,In_935);
nand U2095 (N_2095,In_2547,In_455);
nor U2096 (N_2096,In_355,In_2869);
or U2097 (N_2097,In_551,In_1098);
nand U2098 (N_2098,In_2031,In_1272);
nor U2099 (N_2099,In_1535,In_903);
and U2100 (N_2100,In_877,In_2888);
xor U2101 (N_2101,In_2104,In_1388);
xor U2102 (N_2102,In_422,In_1794);
or U2103 (N_2103,In_1432,In_1623);
and U2104 (N_2104,In_586,In_484);
xnor U2105 (N_2105,In_146,In_2678);
or U2106 (N_2106,In_1202,In_2556);
or U2107 (N_2107,In_263,In_1481);
nor U2108 (N_2108,In_2639,In_1740);
and U2109 (N_2109,In_1150,In_2488);
and U2110 (N_2110,In_363,In_953);
and U2111 (N_2111,In_2002,In_2954);
or U2112 (N_2112,In_1381,In_1443);
nor U2113 (N_2113,In_2885,In_1702);
and U2114 (N_2114,In_1151,In_1986);
xnor U2115 (N_2115,In_2350,In_2213);
and U2116 (N_2116,In_438,In_2539);
nand U2117 (N_2117,In_2041,In_2119);
or U2118 (N_2118,In_1052,In_1364);
nor U2119 (N_2119,In_2925,In_450);
nor U2120 (N_2120,In_1443,In_2230);
xnor U2121 (N_2121,In_1454,In_824);
nor U2122 (N_2122,In_709,In_829);
and U2123 (N_2123,In_601,In_786);
nand U2124 (N_2124,In_1505,In_2226);
nand U2125 (N_2125,In_81,In_2761);
nand U2126 (N_2126,In_1802,In_1379);
nand U2127 (N_2127,In_1246,In_2900);
nor U2128 (N_2128,In_1334,In_564);
or U2129 (N_2129,In_1893,In_242);
nor U2130 (N_2130,In_1937,In_1233);
nand U2131 (N_2131,In_2136,In_695);
nand U2132 (N_2132,In_2548,In_1873);
xor U2133 (N_2133,In_2271,In_1006);
nor U2134 (N_2134,In_926,In_1258);
and U2135 (N_2135,In_2777,In_157);
nor U2136 (N_2136,In_465,In_534);
nor U2137 (N_2137,In_586,In_2639);
or U2138 (N_2138,In_869,In_2110);
and U2139 (N_2139,In_1736,In_198);
nand U2140 (N_2140,In_2106,In_2774);
or U2141 (N_2141,In_1706,In_571);
nand U2142 (N_2142,In_1891,In_623);
xor U2143 (N_2143,In_1719,In_1437);
xnor U2144 (N_2144,In_1888,In_1300);
nor U2145 (N_2145,In_1799,In_2146);
nand U2146 (N_2146,In_51,In_2802);
nand U2147 (N_2147,In_2408,In_2932);
nor U2148 (N_2148,In_280,In_2267);
nor U2149 (N_2149,In_504,In_1883);
nor U2150 (N_2150,In_352,In_2193);
nor U2151 (N_2151,In_762,In_1749);
xnor U2152 (N_2152,In_2315,In_2219);
and U2153 (N_2153,In_1931,In_504);
and U2154 (N_2154,In_1537,In_1445);
nand U2155 (N_2155,In_933,In_1677);
nand U2156 (N_2156,In_663,In_916);
nor U2157 (N_2157,In_108,In_2664);
xnor U2158 (N_2158,In_1369,In_1055);
or U2159 (N_2159,In_1605,In_7);
and U2160 (N_2160,In_1420,In_1605);
nand U2161 (N_2161,In_1495,In_45);
and U2162 (N_2162,In_2344,In_2476);
or U2163 (N_2163,In_2676,In_323);
nor U2164 (N_2164,In_69,In_654);
or U2165 (N_2165,In_64,In_2694);
nand U2166 (N_2166,In_2984,In_2576);
and U2167 (N_2167,In_2766,In_2518);
nor U2168 (N_2168,In_2537,In_603);
nor U2169 (N_2169,In_2837,In_2623);
nor U2170 (N_2170,In_2944,In_2170);
nor U2171 (N_2171,In_1529,In_2354);
nand U2172 (N_2172,In_1597,In_499);
and U2173 (N_2173,In_2999,In_439);
nand U2174 (N_2174,In_2427,In_2820);
nor U2175 (N_2175,In_1946,In_944);
nor U2176 (N_2176,In_99,In_70);
xor U2177 (N_2177,In_1780,In_1950);
or U2178 (N_2178,In_2329,In_1412);
nor U2179 (N_2179,In_1108,In_1330);
nand U2180 (N_2180,In_1914,In_2904);
xor U2181 (N_2181,In_947,In_2375);
nor U2182 (N_2182,In_2285,In_1827);
nor U2183 (N_2183,In_1422,In_1578);
nand U2184 (N_2184,In_696,In_211);
xor U2185 (N_2185,In_2091,In_2728);
nor U2186 (N_2186,In_438,In_1870);
and U2187 (N_2187,In_2531,In_2037);
and U2188 (N_2188,In_2427,In_1502);
nor U2189 (N_2189,In_2051,In_208);
xor U2190 (N_2190,In_2516,In_2145);
nor U2191 (N_2191,In_1622,In_11);
or U2192 (N_2192,In_1870,In_2297);
and U2193 (N_2193,In_2318,In_956);
or U2194 (N_2194,In_545,In_2115);
nand U2195 (N_2195,In_685,In_1203);
nor U2196 (N_2196,In_2335,In_1895);
nor U2197 (N_2197,In_2525,In_954);
nand U2198 (N_2198,In_1192,In_1790);
nor U2199 (N_2199,In_2159,In_2288);
nand U2200 (N_2200,In_1776,In_2758);
xnor U2201 (N_2201,In_1739,In_1635);
or U2202 (N_2202,In_2268,In_142);
nor U2203 (N_2203,In_1636,In_2424);
and U2204 (N_2204,In_2669,In_2787);
or U2205 (N_2205,In_2775,In_2254);
or U2206 (N_2206,In_1229,In_469);
or U2207 (N_2207,In_2769,In_91);
nor U2208 (N_2208,In_597,In_1007);
xnor U2209 (N_2209,In_489,In_999);
xnor U2210 (N_2210,In_583,In_1008);
or U2211 (N_2211,In_424,In_1643);
and U2212 (N_2212,In_22,In_2968);
or U2213 (N_2213,In_2018,In_1711);
nand U2214 (N_2214,In_2674,In_1659);
xnor U2215 (N_2215,In_640,In_2133);
or U2216 (N_2216,In_2952,In_550);
nor U2217 (N_2217,In_187,In_754);
nor U2218 (N_2218,In_2304,In_1343);
nand U2219 (N_2219,In_2136,In_532);
nor U2220 (N_2220,In_1259,In_1340);
nor U2221 (N_2221,In_885,In_1185);
or U2222 (N_2222,In_555,In_234);
or U2223 (N_2223,In_253,In_1577);
or U2224 (N_2224,In_2641,In_2360);
nand U2225 (N_2225,In_2419,In_2130);
or U2226 (N_2226,In_1863,In_339);
nor U2227 (N_2227,In_2838,In_1413);
nor U2228 (N_2228,In_2870,In_2615);
nand U2229 (N_2229,In_1917,In_758);
or U2230 (N_2230,In_1150,In_2212);
xnor U2231 (N_2231,In_927,In_262);
nor U2232 (N_2232,In_959,In_1677);
nor U2233 (N_2233,In_1356,In_1045);
xnor U2234 (N_2234,In_1470,In_2891);
nand U2235 (N_2235,In_2268,In_2131);
and U2236 (N_2236,In_2835,In_708);
xor U2237 (N_2237,In_1607,In_1086);
nor U2238 (N_2238,In_611,In_1495);
nor U2239 (N_2239,In_713,In_636);
and U2240 (N_2240,In_2816,In_681);
nand U2241 (N_2241,In_347,In_2180);
or U2242 (N_2242,In_1263,In_1811);
and U2243 (N_2243,In_1527,In_393);
nand U2244 (N_2244,In_1538,In_2663);
and U2245 (N_2245,In_2041,In_278);
and U2246 (N_2246,In_905,In_1031);
nor U2247 (N_2247,In_1358,In_1064);
nor U2248 (N_2248,In_1425,In_2049);
or U2249 (N_2249,In_1932,In_2046);
xor U2250 (N_2250,In_2368,In_377);
and U2251 (N_2251,In_2635,In_2810);
or U2252 (N_2252,In_1338,In_1765);
and U2253 (N_2253,In_1851,In_153);
xnor U2254 (N_2254,In_1421,In_2741);
or U2255 (N_2255,In_1204,In_1506);
and U2256 (N_2256,In_934,In_994);
xnor U2257 (N_2257,In_2361,In_1679);
or U2258 (N_2258,In_1384,In_2388);
or U2259 (N_2259,In_2158,In_2514);
nor U2260 (N_2260,In_1341,In_457);
xnor U2261 (N_2261,In_2814,In_1733);
nand U2262 (N_2262,In_1304,In_1865);
or U2263 (N_2263,In_2838,In_833);
nor U2264 (N_2264,In_1859,In_1608);
or U2265 (N_2265,In_110,In_2350);
nor U2266 (N_2266,In_513,In_1469);
and U2267 (N_2267,In_1625,In_1608);
nor U2268 (N_2268,In_1151,In_69);
xnor U2269 (N_2269,In_1430,In_1727);
nor U2270 (N_2270,In_351,In_1735);
and U2271 (N_2271,In_1343,In_1392);
nand U2272 (N_2272,In_1752,In_1781);
and U2273 (N_2273,In_1801,In_999);
or U2274 (N_2274,In_1062,In_1813);
nand U2275 (N_2275,In_1738,In_2506);
or U2276 (N_2276,In_2192,In_1396);
or U2277 (N_2277,In_398,In_1240);
xnor U2278 (N_2278,In_2378,In_1288);
xor U2279 (N_2279,In_2624,In_2618);
nor U2280 (N_2280,In_1508,In_2136);
nand U2281 (N_2281,In_701,In_157);
and U2282 (N_2282,In_48,In_722);
or U2283 (N_2283,In_2155,In_1559);
and U2284 (N_2284,In_1310,In_2840);
xor U2285 (N_2285,In_2097,In_2601);
and U2286 (N_2286,In_1655,In_409);
nand U2287 (N_2287,In_476,In_1901);
or U2288 (N_2288,In_2027,In_1426);
nand U2289 (N_2289,In_514,In_48);
nor U2290 (N_2290,In_2468,In_1762);
xnor U2291 (N_2291,In_545,In_2962);
nor U2292 (N_2292,In_1356,In_2730);
or U2293 (N_2293,In_2472,In_1591);
nor U2294 (N_2294,In_1779,In_2769);
or U2295 (N_2295,In_460,In_1671);
nor U2296 (N_2296,In_2240,In_633);
nand U2297 (N_2297,In_847,In_2468);
or U2298 (N_2298,In_1007,In_1657);
nor U2299 (N_2299,In_1676,In_185);
or U2300 (N_2300,In_297,In_2913);
nand U2301 (N_2301,In_2232,In_1837);
nor U2302 (N_2302,In_2906,In_1360);
xnor U2303 (N_2303,In_1712,In_115);
and U2304 (N_2304,In_586,In_1057);
nor U2305 (N_2305,In_50,In_998);
nand U2306 (N_2306,In_1815,In_424);
or U2307 (N_2307,In_1255,In_2963);
and U2308 (N_2308,In_1220,In_979);
or U2309 (N_2309,In_2726,In_212);
or U2310 (N_2310,In_1590,In_254);
nor U2311 (N_2311,In_2503,In_471);
nand U2312 (N_2312,In_2630,In_452);
and U2313 (N_2313,In_2484,In_1515);
xnor U2314 (N_2314,In_2615,In_2308);
nor U2315 (N_2315,In_563,In_1356);
nand U2316 (N_2316,In_1346,In_2488);
nor U2317 (N_2317,In_1767,In_268);
xnor U2318 (N_2318,In_751,In_682);
or U2319 (N_2319,In_1619,In_1174);
and U2320 (N_2320,In_107,In_1535);
nand U2321 (N_2321,In_2298,In_16);
and U2322 (N_2322,In_427,In_2014);
or U2323 (N_2323,In_1946,In_2593);
nor U2324 (N_2324,In_2706,In_835);
or U2325 (N_2325,In_2668,In_223);
or U2326 (N_2326,In_2091,In_2510);
nor U2327 (N_2327,In_2565,In_1411);
nor U2328 (N_2328,In_2237,In_2056);
or U2329 (N_2329,In_678,In_605);
or U2330 (N_2330,In_257,In_2895);
nor U2331 (N_2331,In_967,In_1988);
or U2332 (N_2332,In_1341,In_523);
nor U2333 (N_2333,In_1084,In_558);
nand U2334 (N_2334,In_2366,In_514);
or U2335 (N_2335,In_392,In_985);
and U2336 (N_2336,In_2069,In_2301);
nand U2337 (N_2337,In_101,In_2820);
nand U2338 (N_2338,In_2804,In_1629);
nor U2339 (N_2339,In_2786,In_1363);
nor U2340 (N_2340,In_2682,In_682);
nor U2341 (N_2341,In_279,In_2606);
nand U2342 (N_2342,In_1674,In_2430);
nor U2343 (N_2343,In_2404,In_1379);
nor U2344 (N_2344,In_2724,In_870);
or U2345 (N_2345,In_863,In_2407);
nor U2346 (N_2346,In_2989,In_400);
nand U2347 (N_2347,In_1953,In_1605);
and U2348 (N_2348,In_2901,In_916);
or U2349 (N_2349,In_2690,In_1110);
nor U2350 (N_2350,In_2919,In_2067);
or U2351 (N_2351,In_1089,In_46);
nand U2352 (N_2352,In_2056,In_338);
and U2353 (N_2353,In_2539,In_1407);
or U2354 (N_2354,In_791,In_554);
and U2355 (N_2355,In_1462,In_1304);
and U2356 (N_2356,In_1556,In_834);
nor U2357 (N_2357,In_1830,In_1608);
and U2358 (N_2358,In_174,In_2722);
or U2359 (N_2359,In_377,In_2698);
xor U2360 (N_2360,In_1825,In_1076);
and U2361 (N_2361,In_1529,In_1725);
or U2362 (N_2362,In_2846,In_1286);
or U2363 (N_2363,In_1136,In_2440);
nor U2364 (N_2364,In_2039,In_1496);
nand U2365 (N_2365,In_1997,In_2989);
nand U2366 (N_2366,In_2841,In_1266);
or U2367 (N_2367,In_20,In_1399);
or U2368 (N_2368,In_2532,In_2310);
and U2369 (N_2369,In_1546,In_1313);
or U2370 (N_2370,In_1711,In_2785);
or U2371 (N_2371,In_2195,In_1499);
and U2372 (N_2372,In_2113,In_195);
and U2373 (N_2373,In_734,In_2679);
nand U2374 (N_2374,In_598,In_1683);
nand U2375 (N_2375,In_1349,In_1860);
nand U2376 (N_2376,In_912,In_1379);
or U2377 (N_2377,In_578,In_1381);
nand U2378 (N_2378,In_1666,In_1817);
and U2379 (N_2379,In_2650,In_2635);
nor U2380 (N_2380,In_2291,In_46);
and U2381 (N_2381,In_633,In_1102);
nand U2382 (N_2382,In_417,In_390);
and U2383 (N_2383,In_2736,In_1707);
xnor U2384 (N_2384,In_314,In_727);
nand U2385 (N_2385,In_1349,In_2969);
and U2386 (N_2386,In_431,In_1483);
xor U2387 (N_2387,In_1687,In_2355);
nand U2388 (N_2388,In_1649,In_2381);
nor U2389 (N_2389,In_2555,In_765);
or U2390 (N_2390,In_460,In_246);
or U2391 (N_2391,In_2752,In_731);
and U2392 (N_2392,In_1576,In_2606);
nor U2393 (N_2393,In_2917,In_1362);
or U2394 (N_2394,In_2967,In_1728);
or U2395 (N_2395,In_2135,In_1066);
or U2396 (N_2396,In_1560,In_2433);
or U2397 (N_2397,In_2355,In_2187);
or U2398 (N_2398,In_771,In_774);
and U2399 (N_2399,In_1262,In_2109);
or U2400 (N_2400,In_1326,In_2139);
nand U2401 (N_2401,In_1923,In_2044);
or U2402 (N_2402,In_594,In_2154);
or U2403 (N_2403,In_198,In_772);
or U2404 (N_2404,In_447,In_351);
nor U2405 (N_2405,In_2511,In_2294);
or U2406 (N_2406,In_377,In_1714);
or U2407 (N_2407,In_276,In_1184);
xor U2408 (N_2408,In_1068,In_914);
and U2409 (N_2409,In_1957,In_68);
and U2410 (N_2410,In_2472,In_2378);
nand U2411 (N_2411,In_2251,In_1168);
nor U2412 (N_2412,In_2662,In_1179);
and U2413 (N_2413,In_1024,In_562);
and U2414 (N_2414,In_1389,In_2214);
nand U2415 (N_2415,In_1723,In_695);
nor U2416 (N_2416,In_1286,In_951);
and U2417 (N_2417,In_285,In_1890);
and U2418 (N_2418,In_224,In_277);
and U2419 (N_2419,In_492,In_2870);
nor U2420 (N_2420,In_2989,In_1996);
nor U2421 (N_2421,In_1579,In_1434);
or U2422 (N_2422,In_2952,In_1310);
or U2423 (N_2423,In_2499,In_2100);
nor U2424 (N_2424,In_187,In_748);
and U2425 (N_2425,In_2487,In_2676);
nand U2426 (N_2426,In_1526,In_935);
nand U2427 (N_2427,In_2525,In_1106);
nor U2428 (N_2428,In_2597,In_429);
and U2429 (N_2429,In_1143,In_1626);
nor U2430 (N_2430,In_2483,In_1645);
or U2431 (N_2431,In_1914,In_110);
or U2432 (N_2432,In_2786,In_1588);
nand U2433 (N_2433,In_793,In_2898);
and U2434 (N_2434,In_1499,In_2134);
nor U2435 (N_2435,In_2602,In_480);
or U2436 (N_2436,In_274,In_1162);
and U2437 (N_2437,In_2299,In_1042);
nand U2438 (N_2438,In_92,In_1563);
or U2439 (N_2439,In_1099,In_1689);
nor U2440 (N_2440,In_785,In_2202);
nor U2441 (N_2441,In_392,In_2896);
and U2442 (N_2442,In_1911,In_432);
or U2443 (N_2443,In_2774,In_207);
and U2444 (N_2444,In_1225,In_2266);
or U2445 (N_2445,In_1292,In_2435);
or U2446 (N_2446,In_1143,In_2021);
nand U2447 (N_2447,In_1161,In_2768);
or U2448 (N_2448,In_1237,In_1213);
nand U2449 (N_2449,In_661,In_1084);
or U2450 (N_2450,In_2148,In_2007);
nand U2451 (N_2451,In_368,In_1555);
and U2452 (N_2452,In_2323,In_296);
xor U2453 (N_2453,In_445,In_924);
or U2454 (N_2454,In_1608,In_2812);
and U2455 (N_2455,In_2258,In_315);
xnor U2456 (N_2456,In_2290,In_1992);
and U2457 (N_2457,In_374,In_796);
or U2458 (N_2458,In_2157,In_2044);
or U2459 (N_2459,In_1098,In_2115);
or U2460 (N_2460,In_630,In_2375);
and U2461 (N_2461,In_2908,In_359);
nand U2462 (N_2462,In_1742,In_2726);
xnor U2463 (N_2463,In_669,In_2451);
and U2464 (N_2464,In_417,In_44);
and U2465 (N_2465,In_244,In_2155);
nor U2466 (N_2466,In_1718,In_2196);
and U2467 (N_2467,In_2165,In_1884);
nand U2468 (N_2468,In_175,In_747);
or U2469 (N_2469,In_2512,In_498);
xnor U2470 (N_2470,In_805,In_208);
and U2471 (N_2471,In_269,In_1115);
nand U2472 (N_2472,In_197,In_2125);
and U2473 (N_2473,In_2258,In_125);
nor U2474 (N_2474,In_2772,In_226);
and U2475 (N_2475,In_365,In_1504);
nand U2476 (N_2476,In_1953,In_1478);
and U2477 (N_2477,In_953,In_419);
xor U2478 (N_2478,In_770,In_2312);
and U2479 (N_2479,In_216,In_2851);
and U2480 (N_2480,In_2033,In_2394);
and U2481 (N_2481,In_338,In_980);
or U2482 (N_2482,In_39,In_611);
and U2483 (N_2483,In_465,In_2209);
nand U2484 (N_2484,In_487,In_2901);
nor U2485 (N_2485,In_57,In_2005);
xnor U2486 (N_2486,In_2395,In_881);
nand U2487 (N_2487,In_2278,In_1614);
nor U2488 (N_2488,In_569,In_2136);
nor U2489 (N_2489,In_430,In_2369);
xor U2490 (N_2490,In_1133,In_1096);
nand U2491 (N_2491,In_185,In_2001);
nor U2492 (N_2492,In_2937,In_1765);
xor U2493 (N_2493,In_2109,In_612);
or U2494 (N_2494,In_1905,In_1658);
or U2495 (N_2495,In_621,In_710);
nor U2496 (N_2496,In_1889,In_1505);
or U2497 (N_2497,In_842,In_2313);
and U2498 (N_2498,In_491,In_1702);
nand U2499 (N_2499,In_2260,In_2280);
and U2500 (N_2500,In_664,In_2364);
nor U2501 (N_2501,In_717,In_1152);
nand U2502 (N_2502,In_2112,In_140);
or U2503 (N_2503,In_1111,In_2792);
or U2504 (N_2504,In_806,In_535);
and U2505 (N_2505,In_2347,In_1539);
nand U2506 (N_2506,In_213,In_1719);
or U2507 (N_2507,In_2519,In_1200);
or U2508 (N_2508,In_256,In_2891);
xor U2509 (N_2509,In_1659,In_1866);
or U2510 (N_2510,In_1187,In_595);
xor U2511 (N_2511,In_986,In_460);
nor U2512 (N_2512,In_99,In_1574);
nand U2513 (N_2513,In_2727,In_2045);
nand U2514 (N_2514,In_1446,In_464);
and U2515 (N_2515,In_408,In_2979);
and U2516 (N_2516,In_1955,In_1030);
nand U2517 (N_2517,In_1407,In_1987);
or U2518 (N_2518,In_2799,In_2703);
and U2519 (N_2519,In_365,In_1384);
nand U2520 (N_2520,In_455,In_100);
nand U2521 (N_2521,In_2718,In_2375);
or U2522 (N_2522,In_1956,In_2906);
nor U2523 (N_2523,In_1155,In_976);
nor U2524 (N_2524,In_970,In_1112);
and U2525 (N_2525,In_473,In_306);
nor U2526 (N_2526,In_1411,In_264);
xor U2527 (N_2527,In_2831,In_2574);
nor U2528 (N_2528,In_2377,In_794);
nand U2529 (N_2529,In_253,In_2441);
nand U2530 (N_2530,In_430,In_2353);
nand U2531 (N_2531,In_2588,In_295);
nor U2532 (N_2532,In_1659,In_1718);
nand U2533 (N_2533,In_1001,In_934);
nor U2534 (N_2534,In_1609,In_2679);
or U2535 (N_2535,In_2719,In_2563);
and U2536 (N_2536,In_2700,In_1854);
nand U2537 (N_2537,In_449,In_644);
or U2538 (N_2538,In_2053,In_2204);
and U2539 (N_2539,In_1582,In_2395);
or U2540 (N_2540,In_1867,In_1761);
nor U2541 (N_2541,In_676,In_1363);
nor U2542 (N_2542,In_2209,In_936);
and U2543 (N_2543,In_1271,In_1631);
or U2544 (N_2544,In_2116,In_2993);
or U2545 (N_2545,In_1326,In_953);
nor U2546 (N_2546,In_471,In_2427);
and U2547 (N_2547,In_945,In_905);
nand U2548 (N_2548,In_2195,In_125);
and U2549 (N_2549,In_700,In_1847);
xor U2550 (N_2550,In_2049,In_941);
nor U2551 (N_2551,In_2364,In_2698);
or U2552 (N_2552,In_644,In_2211);
or U2553 (N_2553,In_744,In_2215);
nor U2554 (N_2554,In_1723,In_651);
and U2555 (N_2555,In_1279,In_2893);
xor U2556 (N_2556,In_713,In_1678);
nand U2557 (N_2557,In_586,In_761);
xnor U2558 (N_2558,In_1588,In_2367);
and U2559 (N_2559,In_370,In_821);
and U2560 (N_2560,In_2572,In_1216);
nor U2561 (N_2561,In_1352,In_488);
and U2562 (N_2562,In_194,In_73);
nor U2563 (N_2563,In_1,In_1787);
nand U2564 (N_2564,In_1826,In_1666);
or U2565 (N_2565,In_149,In_471);
nor U2566 (N_2566,In_1687,In_1454);
and U2567 (N_2567,In_1187,In_719);
xnor U2568 (N_2568,In_1633,In_216);
nand U2569 (N_2569,In_1869,In_1596);
or U2570 (N_2570,In_956,In_1565);
and U2571 (N_2571,In_2284,In_1909);
or U2572 (N_2572,In_2787,In_109);
nor U2573 (N_2573,In_1248,In_123);
xor U2574 (N_2574,In_268,In_1962);
nor U2575 (N_2575,In_988,In_812);
nand U2576 (N_2576,In_2174,In_2239);
nand U2577 (N_2577,In_2311,In_2027);
and U2578 (N_2578,In_2342,In_1134);
nand U2579 (N_2579,In_111,In_1347);
and U2580 (N_2580,In_1090,In_1395);
nor U2581 (N_2581,In_860,In_310);
nand U2582 (N_2582,In_562,In_1484);
and U2583 (N_2583,In_2926,In_183);
xor U2584 (N_2584,In_2818,In_2361);
or U2585 (N_2585,In_1512,In_2414);
nor U2586 (N_2586,In_2129,In_2385);
xnor U2587 (N_2587,In_2034,In_377);
and U2588 (N_2588,In_157,In_2837);
or U2589 (N_2589,In_2831,In_188);
xor U2590 (N_2590,In_2211,In_916);
or U2591 (N_2591,In_1407,In_67);
nand U2592 (N_2592,In_2525,In_2576);
or U2593 (N_2593,In_192,In_2594);
nor U2594 (N_2594,In_183,In_460);
or U2595 (N_2595,In_2840,In_1934);
nand U2596 (N_2596,In_367,In_728);
and U2597 (N_2597,In_1118,In_249);
nor U2598 (N_2598,In_755,In_1151);
and U2599 (N_2599,In_2604,In_1755);
xnor U2600 (N_2600,In_1769,In_2217);
nor U2601 (N_2601,In_2023,In_479);
nor U2602 (N_2602,In_1455,In_176);
nand U2603 (N_2603,In_2360,In_2135);
and U2604 (N_2604,In_933,In_1709);
and U2605 (N_2605,In_1796,In_2856);
nor U2606 (N_2606,In_667,In_1316);
nor U2607 (N_2607,In_2324,In_85);
xnor U2608 (N_2608,In_2520,In_2385);
and U2609 (N_2609,In_328,In_709);
or U2610 (N_2610,In_843,In_1789);
nand U2611 (N_2611,In_1756,In_504);
nand U2612 (N_2612,In_70,In_2526);
and U2613 (N_2613,In_2049,In_2315);
nand U2614 (N_2614,In_2875,In_1048);
or U2615 (N_2615,In_1268,In_2158);
nor U2616 (N_2616,In_312,In_733);
nor U2617 (N_2617,In_1649,In_646);
or U2618 (N_2618,In_341,In_1687);
and U2619 (N_2619,In_46,In_2895);
and U2620 (N_2620,In_2643,In_175);
nand U2621 (N_2621,In_1864,In_235);
and U2622 (N_2622,In_2755,In_570);
or U2623 (N_2623,In_1139,In_656);
or U2624 (N_2624,In_285,In_715);
xnor U2625 (N_2625,In_1383,In_2772);
nor U2626 (N_2626,In_10,In_2069);
or U2627 (N_2627,In_1430,In_1607);
and U2628 (N_2628,In_940,In_504);
nor U2629 (N_2629,In_1798,In_2653);
nor U2630 (N_2630,In_219,In_1331);
nand U2631 (N_2631,In_227,In_831);
xnor U2632 (N_2632,In_2377,In_2698);
and U2633 (N_2633,In_435,In_2414);
and U2634 (N_2634,In_613,In_727);
nor U2635 (N_2635,In_2540,In_2954);
or U2636 (N_2636,In_2089,In_1360);
nand U2637 (N_2637,In_2546,In_2020);
and U2638 (N_2638,In_2961,In_1229);
nor U2639 (N_2639,In_254,In_1614);
or U2640 (N_2640,In_1382,In_898);
nand U2641 (N_2641,In_2419,In_763);
nand U2642 (N_2642,In_2470,In_2278);
nor U2643 (N_2643,In_1535,In_1578);
nor U2644 (N_2644,In_418,In_948);
or U2645 (N_2645,In_273,In_1943);
nor U2646 (N_2646,In_932,In_2050);
nand U2647 (N_2647,In_476,In_2404);
xnor U2648 (N_2648,In_1343,In_857);
xnor U2649 (N_2649,In_959,In_2316);
nand U2650 (N_2650,In_1165,In_1916);
nand U2651 (N_2651,In_2219,In_95);
nand U2652 (N_2652,In_153,In_1750);
nor U2653 (N_2653,In_1123,In_670);
nor U2654 (N_2654,In_2344,In_496);
nand U2655 (N_2655,In_2447,In_2795);
nand U2656 (N_2656,In_2322,In_2515);
and U2657 (N_2657,In_2043,In_249);
and U2658 (N_2658,In_1354,In_310);
and U2659 (N_2659,In_2863,In_242);
nor U2660 (N_2660,In_490,In_709);
or U2661 (N_2661,In_2718,In_226);
nor U2662 (N_2662,In_687,In_2684);
nor U2663 (N_2663,In_1565,In_226);
nor U2664 (N_2664,In_2097,In_322);
or U2665 (N_2665,In_2763,In_167);
or U2666 (N_2666,In_806,In_673);
or U2667 (N_2667,In_1167,In_771);
nor U2668 (N_2668,In_2187,In_62);
or U2669 (N_2669,In_2487,In_2793);
or U2670 (N_2670,In_626,In_695);
and U2671 (N_2671,In_1576,In_933);
nor U2672 (N_2672,In_2196,In_1550);
xor U2673 (N_2673,In_1340,In_816);
nand U2674 (N_2674,In_2547,In_64);
xor U2675 (N_2675,In_1938,In_1217);
and U2676 (N_2676,In_2661,In_1769);
xnor U2677 (N_2677,In_177,In_644);
or U2678 (N_2678,In_2030,In_484);
xnor U2679 (N_2679,In_2571,In_1375);
or U2680 (N_2680,In_1527,In_1376);
nand U2681 (N_2681,In_395,In_1974);
or U2682 (N_2682,In_1324,In_205);
or U2683 (N_2683,In_654,In_855);
and U2684 (N_2684,In_814,In_78);
and U2685 (N_2685,In_1801,In_1709);
nor U2686 (N_2686,In_1960,In_1495);
xnor U2687 (N_2687,In_617,In_937);
or U2688 (N_2688,In_1438,In_1331);
nor U2689 (N_2689,In_1093,In_682);
nand U2690 (N_2690,In_2021,In_2072);
nor U2691 (N_2691,In_1104,In_2379);
or U2692 (N_2692,In_1567,In_2881);
and U2693 (N_2693,In_1487,In_2163);
nor U2694 (N_2694,In_188,In_1276);
nand U2695 (N_2695,In_1462,In_1536);
xnor U2696 (N_2696,In_2157,In_922);
or U2697 (N_2697,In_2119,In_1108);
nor U2698 (N_2698,In_2087,In_2191);
xnor U2699 (N_2699,In_2660,In_1249);
or U2700 (N_2700,In_371,In_1071);
nand U2701 (N_2701,In_1787,In_389);
or U2702 (N_2702,In_1080,In_1945);
xnor U2703 (N_2703,In_2403,In_2571);
or U2704 (N_2704,In_676,In_973);
and U2705 (N_2705,In_2446,In_1447);
or U2706 (N_2706,In_2625,In_2077);
or U2707 (N_2707,In_1394,In_1059);
nand U2708 (N_2708,In_2504,In_1201);
nor U2709 (N_2709,In_1959,In_1760);
nor U2710 (N_2710,In_548,In_1996);
nor U2711 (N_2711,In_1790,In_956);
and U2712 (N_2712,In_1272,In_2241);
nand U2713 (N_2713,In_623,In_860);
and U2714 (N_2714,In_1451,In_2407);
nand U2715 (N_2715,In_1582,In_1748);
nor U2716 (N_2716,In_2903,In_456);
nand U2717 (N_2717,In_2143,In_698);
nand U2718 (N_2718,In_1313,In_234);
nor U2719 (N_2719,In_1483,In_1998);
nor U2720 (N_2720,In_1539,In_2251);
and U2721 (N_2721,In_589,In_2802);
xnor U2722 (N_2722,In_1867,In_435);
and U2723 (N_2723,In_1271,In_98);
and U2724 (N_2724,In_2501,In_1178);
and U2725 (N_2725,In_309,In_773);
nor U2726 (N_2726,In_2728,In_2194);
nand U2727 (N_2727,In_213,In_2460);
and U2728 (N_2728,In_1938,In_2039);
nor U2729 (N_2729,In_151,In_993);
or U2730 (N_2730,In_1309,In_520);
and U2731 (N_2731,In_706,In_1279);
nand U2732 (N_2732,In_2666,In_574);
nand U2733 (N_2733,In_1762,In_677);
xor U2734 (N_2734,In_1534,In_1260);
nor U2735 (N_2735,In_1551,In_1595);
nand U2736 (N_2736,In_834,In_2260);
nor U2737 (N_2737,In_770,In_2492);
and U2738 (N_2738,In_24,In_1951);
nand U2739 (N_2739,In_534,In_2745);
nand U2740 (N_2740,In_2091,In_1113);
xor U2741 (N_2741,In_2645,In_1053);
or U2742 (N_2742,In_2733,In_142);
nand U2743 (N_2743,In_352,In_1368);
nor U2744 (N_2744,In_611,In_1789);
xnor U2745 (N_2745,In_2889,In_330);
nand U2746 (N_2746,In_1531,In_1465);
or U2747 (N_2747,In_2399,In_1337);
or U2748 (N_2748,In_2764,In_1518);
nor U2749 (N_2749,In_867,In_319);
nand U2750 (N_2750,In_2328,In_570);
nor U2751 (N_2751,In_2841,In_264);
or U2752 (N_2752,In_1587,In_2130);
or U2753 (N_2753,In_1637,In_2859);
xor U2754 (N_2754,In_465,In_1034);
and U2755 (N_2755,In_1780,In_1069);
and U2756 (N_2756,In_26,In_120);
nor U2757 (N_2757,In_636,In_1950);
nor U2758 (N_2758,In_1540,In_2013);
nand U2759 (N_2759,In_1081,In_1681);
and U2760 (N_2760,In_2637,In_1199);
or U2761 (N_2761,In_1084,In_847);
nor U2762 (N_2762,In_1119,In_1198);
or U2763 (N_2763,In_1338,In_245);
nand U2764 (N_2764,In_1941,In_469);
nand U2765 (N_2765,In_1573,In_2689);
or U2766 (N_2766,In_230,In_1041);
nor U2767 (N_2767,In_789,In_2033);
nand U2768 (N_2768,In_1688,In_2891);
nor U2769 (N_2769,In_1852,In_1002);
or U2770 (N_2770,In_2531,In_2307);
nand U2771 (N_2771,In_403,In_2152);
nand U2772 (N_2772,In_1452,In_65);
nand U2773 (N_2773,In_126,In_1167);
and U2774 (N_2774,In_2423,In_531);
xnor U2775 (N_2775,In_2040,In_2797);
or U2776 (N_2776,In_578,In_2203);
or U2777 (N_2777,In_1584,In_2500);
and U2778 (N_2778,In_1960,In_1256);
nor U2779 (N_2779,In_2498,In_2542);
nor U2780 (N_2780,In_353,In_2373);
or U2781 (N_2781,In_2881,In_191);
nor U2782 (N_2782,In_349,In_2066);
nand U2783 (N_2783,In_2799,In_632);
nand U2784 (N_2784,In_600,In_70);
nand U2785 (N_2785,In_138,In_2367);
or U2786 (N_2786,In_2071,In_650);
nor U2787 (N_2787,In_1526,In_1709);
or U2788 (N_2788,In_1888,In_1291);
nor U2789 (N_2789,In_1690,In_2410);
or U2790 (N_2790,In_560,In_2674);
and U2791 (N_2791,In_2308,In_128);
nor U2792 (N_2792,In_435,In_2487);
and U2793 (N_2793,In_2045,In_2774);
or U2794 (N_2794,In_474,In_1285);
or U2795 (N_2795,In_1424,In_1920);
or U2796 (N_2796,In_2924,In_2479);
nand U2797 (N_2797,In_2408,In_1562);
nand U2798 (N_2798,In_26,In_655);
and U2799 (N_2799,In_189,In_1973);
and U2800 (N_2800,In_2684,In_1277);
or U2801 (N_2801,In_426,In_347);
and U2802 (N_2802,In_335,In_1601);
xor U2803 (N_2803,In_2540,In_2643);
nand U2804 (N_2804,In_2109,In_1263);
or U2805 (N_2805,In_1637,In_2207);
and U2806 (N_2806,In_1257,In_4);
and U2807 (N_2807,In_2183,In_75);
xor U2808 (N_2808,In_2625,In_308);
nor U2809 (N_2809,In_2173,In_1994);
nor U2810 (N_2810,In_1125,In_537);
nor U2811 (N_2811,In_1704,In_1581);
nand U2812 (N_2812,In_2948,In_2840);
or U2813 (N_2813,In_2142,In_2758);
or U2814 (N_2814,In_851,In_2473);
or U2815 (N_2815,In_826,In_45);
nand U2816 (N_2816,In_102,In_1460);
nand U2817 (N_2817,In_2696,In_1650);
nor U2818 (N_2818,In_1803,In_2538);
or U2819 (N_2819,In_2937,In_1325);
and U2820 (N_2820,In_1669,In_1320);
or U2821 (N_2821,In_1584,In_2917);
nand U2822 (N_2822,In_1882,In_2532);
nor U2823 (N_2823,In_1067,In_971);
nand U2824 (N_2824,In_1438,In_1285);
xor U2825 (N_2825,In_671,In_1485);
or U2826 (N_2826,In_1355,In_236);
and U2827 (N_2827,In_1218,In_2733);
or U2828 (N_2828,In_1602,In_2486);
and U2829 (N_2829,In_1543,In_2761);
xor U2830 (N_2830,In_319,In_2676);
and U2831 (N_2831,In_2167,In_493);
or U2832 (N_2832,In_1009,In_44);
nor U2833 (N_2833,In_167,In_2199);
nor U2834 (N_2834,In_1864,In_231);
nand U2835 (N_2835,In_1505,In_2708);
or U2836 (N_2836,In_1628,In_1501);
nor U2837 (N_2837,In_2245,In_2614);
and U2838 (N_2838,In_96,In_2758);
nor U2839 (N_2839,In_318,In_1014);
and U2840 (N_2840,In_2542,In_2890);
nand U2841 (N_2841,In_612,In_543);
or U2842 (N_2842,In_1015,In_908);
nand U2843 (N_2843,In_2927,In_2482);
nor U2844 (N_2844,In_2789,In_828);
xnor U2845 (N_2845,In_1075,In_390);
and U2846 (N_2846,In_419,In_1869);
or U2847 (N_2847,In_2426,In_2138);
and U2848 (N_2848,In_1994,In_2090);
or U2849 (N_2849,In_2580,In_877);
nor U2850 (N_2850,In_1617,In_1370);
or U2851 (N_2851,In_496,In_2113);
xor U2852 (N_2852,In_1569,In_1506);
xor U2853 (N_2853,In_2643,In_2078);
nand U2854 (N_2854,In_2126,In_2082);
xnor U2855 (N_2855,In_259,In_2260);
nor U2856 (N_2856,In_121,In_626);
or U2857 (N_2857,In_2481,In_427);
or U2858 (N_2858,In_753,In_1122);
nor U2859 (N_2859,In_2099,In_970);
nand U2860 (N_2860,In_2480,In_2462);
xor U2861 (N_2861,In_2219,In_1518);
nor U2862 (N_2862,In_1255,In_2259);
xnor U2863 (N_2863,In_1272,In_2302);
or U2864 (N_2864,In_2235,In_2018);
or U2865 (N_2865,In_678,In_1969);
nand U2866 (N_2866,In_2769,In_1765);
or U2867 (N_2867,In_1648,In_1649);
nand U2868 (N_2868,In_2608,In_857);
nor U2869 (N_2869,In_2486,In_2247);
xor U2870 (N_2870,In_2949,In_2049);
nand U2871 (N_2871,In_1609,In_1012);
nand U2872 (N_2872,In_2833,In_2821);
or U2873 (N_2873,In_1097,In_1106);
or U2874 (N_2874,In_2118,In_2138);
xnor U2875 (N_2875,In_1477,In_966);
or U2876 (N_2876,In_2907,In_47);
nand U2877 (N_2877,In_2912,In_272);
or U2878 (N_2878,In_737,In_542);
or U2879 (N_2879,In_2274,In_660);
or U2880 (N_2880,In_354,In_2004);
and U2881 (N_2881,In_1683,In_646);
and U2882 (N_2882,In_2436,In_1737);
or U2883 (N_2883,In_246,In_1851);
nor U2884 (N_2884,In_1598,In_1833);
nand U2885 (N_2885,In_136,In_1652);
or U2886 (N_2886,In_2579,In_761);
nand U2887 (N_2887,In_444,In_2437);
and U2888 (N_2888,In_743,In_419);
or U2889 (N_2889,In_2527,In_2220);
or U2890 (N_2890,In_2966,In_849);
or U2891 (N_2891,In_2978,In_1582);
xor U2892 (N_2892,In_2906,In_896);
nand U2893 (N_2893,In_2410,In_1361);
and U2894 (N_2894,In_777,In_1719);
nand U2895 (N_2895,In_1467,In_2639);
nor U2896 (N_2896,In_303,In_1374);
nor U2897 (N_2897,In_150,In_2915);
or U2898 (N_2898,In_554,In_1541);
or U2899 (N_2899,In_2767,In_2840);
nor U2900 (N_2900,In_458,In_1470);
or U2901 (N_2901,In_2819,In_1616);
nor U2902 (N_2902,In_681,In_2340);
nor U2903 (N_2903,In_2446,In_1565);
xnor U2904 (N_2904,In_1288,In_1996);
nand U2905 (N_2905,In_3,In_363);
and U2906 (N_2906,In_2730,In_792);
or U2907 (N_2907,In_1855,In_2334);
xnor U2908 (N_2908,In_927,In_58);
and U2909 (N_2909,In_2214,In_270);
nor U2910 (N_2910,In_781,In_471);
nand U2911 (N_2911,In_694,In_2626);
nand U2912 (N_2912,In_359,In_2302);
nor U2913 (N_2913,In_2103,In_2833);
and U2914 (N_2914,In_730,In_302);
nor U2915 (N_2915,In_1945,In_2058);
nand U2916 (N_2916,In_13,In_1674);
xnor U2917 (N_2917,In_1805,In_2187);
nand U2918 (N_2918,In_133,In_488);
nand U2919 (N_2919,In_1083,In_91);
nor U2920 (N_2920,In_242,In_1903);
nand U2921 (N_2921,In_1772,In_1326);
or U2922 (N_2922,In_643,In_2174);
and U2923 (N_2923,In_1827,In_1281);
and U2924 (N_2924,In_1243,In_1469);
and U2925 (N_2925,In_2494,In_2914);
and U2926 (N_2926,In_267,In_1527);
nand U2927 (N_2927,In_1824,In_2518);
and U2928 (N_2928,In_58,In_1887);
or U2929 (N_2929,In_2041,In_634);
nor U2930 (N_2930,In_173,In_2108);
or U2931 (N_2931,In_446,In_374);
and U2932 (N_2932,In_1862,In_569);
xnor U2933 (N_2933,In_891,In_2176);
nand U2934 (N_2934,In_2964,In_2459);
nor U2935 (N_2935,In_2275,In_1426);
or U2936 (N_2936,In_1751,In_2644);
or U2937 (N_2937,In_815,In_242);
and U2938 (N_2938,In_1569,In_2001);
nand U2939 (N_2939,In_2202,In_2572);
or U2940 (N_2940,In_1273,In_1451);
nor U2941 (N_2941,In_1906,In_553);
nor U2942 (N_2942,In_2038,In_2780);
and U2943 (N_2943,In_1592,In_1551);
nand U2944 (N_2944,In_2249,In_2535);
or U2945 (N_2945,In_937,In_160);
nand U2946 (N_2946,In_383,In_598);
or U2947 (N_2947,In_2024,In_2706);
nand U2948 (N_2948,In_2097,In_2350);
nor U2949 (N_2949,In_2227,In_1090);
nor U2950 (N_2950,In_921,In_2951);
nand U2951 (N_2951,In_164,In_255);
nor U2952 (N_2952,In_1592,In_905);
and U2953 (N_2953,In_2571,In_1661);
and U2954 (N_2954,In_526,In_1066);
nor U2955 (N_2955,In_2283,In_798);
and U2956 (N_2956,In_2294,In_1514);
xor U2957 (N_2957,In_1550,In_1533);
and U2958 (N_2958,In_2142,In_1058);
xnor U2959 (N_2959,In_2471,In_495);
xor U2960 (N_2960,In_1169,In_2949);
or U2961 (N_2961,In_2552,In_272);
xor U2962 (N_2962,In_2989,In_2850);
nand U2963 (N_2963,In_451,In_2480);
nand U2964 (N_2964,In_1092,In_1139);
and U2965 (N_2965,In_159,In_67);
nor U2966 (N_2966,In_801,In_1161);
nor U2967 (N_2967,In_857,In_2290);
nor U2968 (N_2968,In_1568,In_493);
and U2969 (N_2969,In_1990,In_2112);
nand U2970 (N_2970,In_680,In_2553);
and U2971 (N_2971,In_1386,In_2234);
and U2972 (N_2972,In_1558,In_880);
nand U2973 (N_2973,In_1874,In_440);
nor U2974 (N_2974,In_335,In_2192);
or U2975 (N_2975,In_1854,In_1568);
or U2976 (N_2976,In_2133,In_2353);
or U2977 (N_2977,In_2237,In_457);
nand U2978 (N_2978,In_72,In_1291);
nand U2979 (N_2979,In_1295,In_176);
nand U2980 (N_2980,In_2875,In_1570);
nor U2981 (N_2981,In_1497,In_1217);
or U2982 (N_2982,In_364,In_583);
or U2983 (N_2983,In_2172,In_1604);
xnor U2984 (N_2984,In_142,In_162);
nor U2985 (N_2985,In_692,In_797);
and U2986 (N_2986,In_2927,In_1917);
or U2987 (N_2987,In_2156,In_891);
or U2988 (N_2988,In_672,In_939);
nor U2989 (N_2989,In_2390,In_1726);
or U2990 (N_2990,In_1468,In_210);
nand U2991 (N_2991,In_1030,In_699);
xnor U2992 (N_2992,In_644,In_915);
nor U2993 (N_2993,In_442,In_2525);
nand U2994 (N_2994,In_584,In_1065);
and U2995 (N_2995,In_1886,In_1659);
nand U2996 (N_2996,In_1560,In_876);
nor U2997 (N_2997,In_2347,In_363);
and U2998 (N_2998,In_474,In_393);
nor U2999 (N_2999,In_692,In_359);
nor U3000 (N_3000,In_1824,In_74);
and U3001 (N_3001,In_716,In_843);
nor U3002 (N_3002,In_905,In_2336);
xnor U3003 (N_3003,In_2187,In_2304);
nor U3004 (N_3004,In_1430,In_1100);
nand U3005 (N_3005,In_2281,In_2437);
nand U3006 (N_3006,In_2726,In_1906);
nand U3007 (N_3007,In_1835,In_2858);
nor U3008 (N_3008,In_2713,In_1790);
xor U3009 (N_3009,In_565,In_170);
xnor U3010 (N_3010,In_304,In_997);
nand U3011 (N_3011,In_480,In_524);
and U3012 (N_3012,In_397,In_2743);
or U3013 (N_3013,In_2770,In_201);
or U3014 (N_3014,In_1026,In_1593);
or U3015 (N_3015,In_1905,In_2591);
nor U3016 (N_3016,In_345,In_631);
nor U3017 (N_3017,In_37,In_632);
nor U3018 (N_3018,In_2727,In_2521);
nor U3019 (N_3019,In_2515,In_1405);
or U3020 (N_3020,In_292,In_855);
nand U3021 (N_3021,In_918,In_2139);
nor U3022 (N_3022,In_1474,In_1392);
and U3023 (N_3023,In_2528,In_589);
nor U3024 (N_3024,In_533,In_1100);
or U3025 (N_3025,In_1241,In_2007);
or U3026 (N_3026,In_2864,In_1385);
nor U3027 (N_3027,In_2643,In_2004);
nor U3028 (N_3028,In_2266,In_506);
nand U3029 (N_3029,In_1542,In_2090);
nor U3030 (N_3030,In_1955,In_2251);
and U3031 (N_3031,In_639,In_2492);
nor U3032 (N_3032,In_215,In_2315);
or U3033 (N_3033,In_1055,In_1214);
nor U3034 (N_3034,In_1799,In_2858);
xor U3035 (N_3035,In_2603,In_2675);
nor U3036 (N_3036,In_286,In_236);
nor U3037 (N_3037,In_1762,In_2331);
nor U3038 (N_3038,In_1303,In_919);
nor U3039 (N_3039,In_2803,In_1043);
nor U3040 (N_3040,In_1741,In_1198);
nand U3041 (N_3041,In_589,In_2301);
and U3042 (N_3042,In_582,In_1907);
nand U3043 (N_3043,In_21,In_2712);
and U3044 (N_3044,In_1498,In_2314);
nor U3045 (N_3045,In_1795,In_2675);
nand U3046 (N_3046,In_2857,In_2354);
nor U3047 (N_3047,In_724,In_947);
or U3048 (N_3048,In_1095,In_2698);
nor U3049 (N_3049,In_2612,In_311);
nor U3050 (N_3050,In_2802,In_2573);
nor U3051 (N_3051,In_1775,In_226);
and U3052 (N_3052,In_799,In_1934);
or U3053 (N_3053,In_1335,In_1264);
or U3054 (N_3054,In_2986,In_275);
xor U3055 (N_3055,In_2940,In_357);
nand U3056 (N_3056,In_95,In_414);
nor U3057 (N_3057,In_2963,In_1554);
or U3058 (N_3058,In_276,In_2762);
and U3059 (N_3059,In_2815,In_2850);
or U3060 (N_3060,In_537,In_1919);
or U3061 (N_3061,In_1115,In_403);
nand U3062 (N_3062,In_1166,In_2370);
nor U3063 (N_3063,In_755,In_2178);
nor U3064 (N_3064,In_583,In_2763);
nor U3065 (N_3065,In_1930,In_194);
and U3066 (N_3066,In_561,In_781);
and U3067 (N_3067,In_1736,In_61);
or U3068 (N_3068,In_1262,In_684);
nor U3069 (N_3069,In_1703,In_2229);
and U3070 (N_3070,In_253,In_1116);
xor U3071 (N_3071,In_2337,In_462);
and U3072 (N_3072,In_2072,In_1433);
or U3073 (N_3073,In_51,In_149);
and U3074 (N_3074,In_1064,In_2403);
and U3075 (N_3075,In_2035,In_2937);
nor U3076 (N_3076,In_1657,In_2236);
nand U3077 (N_3077,In_1790,In_2416);
nor U3078 (N_3078,In_872,In_587);
or U3079 (N_3079,In_1125,In_1781);
nor U3080 (N_3080,In_386,In_145);
or U3081 (N_3081,In_2422,In_365);
or U3082 (N_3082,In_2751,In_2561);
nand U3083 (N_3083,In_2909,In_1278);
nor U3084 (N_3084,In_764,In_103);
or U3085 (N_3085,In_1885,In_2241);
xor U3086 (N_3086,In_2233,In_2146);
nand U3087 (N_3087,In_12,In_1437);
nand U3088 (N_3088,In_624,In_2673);
nand U3089 (N_3089,In_914,In_2432);
xor U3090 (N_3090,In_1876,In_962);
or U3091 (N_3091,In_45,In_687);
or U3092 (N_3092,In_1533,In_677);
nor U3093 (N_3093,In_2430,In_917);
nand U3094 (N_3094,In_1187,In_259);
nand U3095 (N_3095,In_255,In_1075);
or U3096 (N_3096,In_1039,In_273);
nand U3097 (N_3097,In_1642,In_1683);
nand U3098 (N_3098,In_2184,In_384);
xor U3099 (N_3099,In_836,In_1891);
or U3100 (N_3100,In_2986,In_2991);
and U3101 (N_3101,In_611,In_1024);
or U3102 (N_3102,In_2363,In_469);
nand U3103 (N_3103,In_2485,In_1464);
or U3104 (N_3104,In_1066,In_421);
or U3105 (N_3105,In_2024,In_2612);
nor U3106 (N_3106,In_2752,In_692);
and U3107 (N_3107,In_693,In_1448);
nor U3108 (N_3108,In_126,In_2146);
nand U3109 (N_3109,In_1340,In_840);
and U3110 (N_3110,In_1041,In_1241);
nand U3111 (N_3111,In_1412,In_2832);
nor U3112 (N_3112,In_2731,In_2280);
nor U3113 (N_3113,In_2246,In_2977);
nor U3114 (N_3114,In_1911,In_75);
nor U3115 (N_3115,In_142,In_450);
xnor U3116 (N_3116,In_909,In_1751);
and U3117 (N_3117,In_999,In_144);
or U3118 (N_3118,In_2789,In_495);
nor U3119 (N_3119,In_1426,In_986);
and U3120 (N_3120,In_784,In_2411);
or U3121 (N_3121,In_1691,In_464);
nor U3122 (N_3122,In_350,In_2112);
or U3123 (N_3123,In_364,In_2806);
nand U3124 (N_3124,In_1266,In_2413);
nand U3125 (N_3125,In_1639,In_1012);
and U3126 (N_3126,In_228,In_748);
nor U3127 (N_3127,In_498,In_2752);
nand U3128 (N_3128,In_818,In_2818);
and U3129 (N_3129,In_2020,In_2584);
and U3130 (N_3130,In_1705,In_1139);
xor U3131 (N_3131,In_1550,In_2748);
or U3132 (N_3132,In_811,In_1353);
nor U3133 (N_3133,In_1633,In_2042);
or U3134 (N_3134,In_385,In_144);
nor U3135 (N_3135,In_2803,In_1623);
nor U3136 (N_3136,In_2433,In_1104);
nand U3137 (N_3137,In_2772,In_1627);
xor U3138 (N_3138,In_536,In_2712);
or U3139 (N_3139,In_1346,In_720);
or U3140 (N_3140,In_788,In_798);
and U3141 (N_3141,In_947,In_825);
nor U3142 (N_3142,In_2387,In_1660);
nor U3143 (N_3143,In_688,In_465);
xnor U3144 (N_3144,In_2151,In_2959);
nor U3145 (N_3145,In_1533,In_1045);
nand U3146 (N_3146,In_556,In_142);
nor U3147 (N_3147,In_550,In_930);
nor U3148 (N_3148,In_1244,In_2899);
or U3149 (N_3149,In_1171,In_2017);
or U3150 (N_3150,In_2266,In_402);
or U3151 (N_3151,In_1917,In_1603);
nor U3152 (N_3152,In_1718,In_1551);
and U3153 (N_3153,In_2729,In_1955);
xnor U3154 (N_3154,In_165,In_12);
or U3155 (N_3155,In_672,In_1123);
nor U3156 (N_3156,In_1178,In_1574);
nand U3157 (N_3157,In_788,In_2600);
nand U3158 (N_3158,In_811,In_1984);
and U3159 (N_3159,In_382,In_2465);
nor U3160 (N_3160,In_2361,In_972);
nand U3161 (N_3161,In_308,In_2544);
nor U3162 (N_3162,In_1612,In_2533);
nand U3163 (N_3163,In_1074,In_738);
nor U3164 (N_3164,In_488,In_236);
or U3165 (N_3165,In_1719,In_2954);
or U3166 (N_3166,In_941,In_761);
nor U3167 (N_3167,In_2495,In_2827);
and U3168 (N_3168,In_1535,In_2831);
or U3169 (N_3169,In_2384,In_1400);
or U3170 (N_3170,In_2984,In_1523);
or U3171 (N_3171,In_2156,In_875);
nand U3172 (N_3172,In_1722,In_1364);
nand U3173 (N_3173,In_984,In_2356);
nand U3174 (N_3174,In_1470,In_1783);
and U3175 (N_3175,In_2178,In_1198);
and U3176 (N_3176,In_2520,In_970);
and U3177 (N_3177,In_723,In_446);
nor U3178 (N_3178,In_2599,In_2182);
or U3179 (N_3179,In_2068,In_346);
nand U3180 (N_3180,In_561,In_2227);
nand U3181 (N_3181,In_110,In_2547);
or U3182 (N_3182,In_824,In_2409);
and U3183 (N_3183,In_2955,In_2017);
or U3184 (N_3184,In_1127,In_521);
xnor U3185 (N_3185,In_1468,In_864);
or U3186 (N_3186,In_1323,In_1904);
and U3187 (N_3187,In_1913,In_1069);
and U3188 (N_3188,In_506,In_2782);
nor U3189 (N_3189,In_1171,In_2894);
and U3190 (N_3190,In_2516,In_2156);
nor U3191 (N_3191,In_1388,In_181);
or U3192 (N_3192,In_2787,In_857);
or U3193 (N_3193,In_225,In_2967);
nor U3194 (N_3194,In_1820,In_2206);
or U3195 (N_3195,In_52,In_2001);
and U3196 (N_3196,In_1554,In_1114);
nand U3197 (N_3197,In_1496,In_616);
and U3198 (N_3198,In_1927,In_171);
nand U3199 (N_3199,In_488,In_554);
or U3200 (N_3200,In_1588,In_126);
nand U3201 (N_3201,In_672,In_1967);
and U3202 (N_3202,In_2508,In_1440);
xnor U3203 (N_3203,In_1003,In_749);
and U3204 (N_3204,In_1391,In_2263);
nand U3205 (N_3205,In_2984,In_1591);
nand U3206 (N_3206,In_1848,In_1856);
and U3207 (N_3207,In_701,In_1894);
nand U3208 (N_3208,In_2841,In_1790);
nand U3209 (N_3209,In_2416,In_561);
nand U3210 (N_3210,In_769,In_2305);
nand U3211 (N_3211,In_1654,In_1894);
or U3212 (N_3212,In_2333,In_2936);
xor U3213 (N_3213,In_1700,In_925);
and U3214 (N_3214,In_303,In_141);
or U3215 (N_3215,In_80,In_46);
nor U3216 (N_3216,In_1544,In_30);
nand U3217 (N_3217,In_2502,In_1051);
nor U3218 (N_3218,In_36,In_914);
nor U3219 (N_3219,In_697,In_2866);
nand U3220 (N_3220,In_2054,In_1452);
nor U3221 (N_3221,In_2602,In_921);
nand U3222 (N_3222,In_1812,In_218);
or U3223 (N_3223,In_681,In_615);
xor U3224 (N_3224,In_1004,In_1454);
or U3225 (N_3225,In_2855,In_2182);
or U3226 (N_3226,In_2797,In_349);
and U3227 (N_3227,In_86,In_869);
nor U3228 (N_3228,In_286,In_2495);
xnor U3229 (N_3229,In_2344,In_640);
nand U3230 (N_3230,In_2360,In_421);
or U3231 (N_3231,In_1251,In_395);
nand U3232 (N_3232,In_123,In_1291);
or U3233 (N_3233,In_1539,In_2615);
nor U3234 (N_3234,In_2579,In_2865);
and U3235 (N_3235,In_193,In_2600);
xor U3236 (N_3236,In_833,In_559);
or U3237 (N_3237,In_2799,In_2570);
xnor U3238 (N_3238,In_747,In_1455);
nor U3239 (N_3239,In_699,In_567);
nand U3240 (N_3240,In_2562,In_1837);
and U3241 (N_3241,In_807,In_247);
or U3242 (N_3242,In_1271,In_1703);
and U3243 (N_3243,In_1849,In_1478);
nor U3244 (N_3244,In_155,In_469);
nor U3245 (N_3245,In_717,In_823);
or U3246 (N_3246,In_1742,In_174);
and U3247 (N_3247,In_1591,In_83);
and U3248 (N_3248,In_2094,In_1513);
nand U3249 (N_3249,In_1314,In_2636);
and U3250 (N_3250,In_898,In_449);
or U3251 (N_3251,In_860,In_97);
nor U3252 (N_3252,In_1588,In_50);
or U3253 (N_3253,In_1063,In_2686);
or U3254 (N_3254,In_2437,In_2718);
and U3255 (N_3255,In_1231,In_879);
and U3256 (N_3256,In_2660,In_1688);
nand U3257 (N_3257,In_721,In_1989);
nor U3258 (N_3258,In_1223,In_73);
nand U3259 (N_3259,In_2092,In_1998);
nor U3260 (N_3260,In_545,In_2958);
nor U3261 (N_3261,In_450,In_2126);
or U3262 (N_3262,In_484,In_678);
and U3263 (N_3263,In_2789,In_2561);
or U3264 (N_3264,In_128,In_1041);
nand U3265 (N_3265,In_2550,In_782);
or U3266 (N_3266,In_2237,In_1017);
nand U3267 (N_3267,In_2605,In_1165);
or U3268 (N_3268,In_2245,In_335);
nor U3269 (N_3269,In_1938,In_2081);
nor U3270 (N_3270,In_138,In_1741);
nand U3271 (N_3271,In_2340,In_2888);
nor U3272 (N_3272,In_1127,In_247);
or U3273 (N_3273,In_2684,In_1184);
and U3274 (N_3274,In_885,In_1606);
xor U3275 (N_3275,In_1341,In_2064);
or U3276 (N_3276,In_1573,In_86);
and U3277 (N_3277,In_2130,In_1927);
nand U3278 (N_3278,In_700,In_2525);
nand U3279 (N_3279,In_373,In_1519);
or U3280 (N_3280,In_946,In_1528);
xnor U3281 (N_3281,In_1160,In_1032);
and U3282 (N_3282,In_1422,In_1976);
xnor U3283 (N_3283,In_2474,In_2692);
nand U3284 (N_3284,In_2559,In_443);
xnor U3285 (N_3285,In_1050,In_1134);
nand U3286 (N_3286,In_687,In_1571);
nand U3287 (N_3287,In_1400,In_2633);
and U3288 (N_3288,In_1234,In_2165);
and U3289 (N_3289,In_1373,In_100);
nor U3290 (N_3290,In_2527,In_771);
or U3291 (N_3291,In_866,In_2866);
and U3292 (N_3292,In_1091,In_1505);
nor U3293 (N_3293,In_2059,In_1272);
or U3294 (N_3294,In_1306,In_765);
and U3295 (N_3295,In_1521,In_2905);
nand U3296 (N_3296,In_1711,In_2254);
and U3297 (N_3297,In_1695,In_525);
and U3298 (N_3298,In_690,In_1059);
nand U3299 (N_3299,In_118,In_1534);
and U3300 (N_3300,In_1500,In_2359);
or U3301 (N_3301,In_2686,In_882);
or U3302 (N_3302,In_2667,In_1667);
or U3303 (N_3303,In_1054,In_2220);
nor U3304 (N_3304,In_2004,In_1033);
and U3305 (N_3305,In_2188,In_1728);
or U3306 (N_3306,In_2756,In_177);
nand U3307 (N_3307,In_2771,In_189);
nor U3308 (N_3308,In_2767,In_2506);
or U3309 (N_3309,In_2333,In_2989);
or U3310 (N_3310,In_1127,In_939);
xnor U3311 (N_3311,In_2126,In_879);
nand U3312 (N_3312,In_768,In_2329);
nor U3313 (N_3313,In_2777,In_2605);
nand U3314 (N_3314,In_1989,In_2447);
nor U3315 (N_3315,In_1203,In_1435);
nor U3316 (N_3316,In_1382,In_753);
nor U3317 (N_3317,In_1985,In_331);
and U3318 (N_3318,In_2568,In_2958);
and U3319 (N_3319,In_1833,In_2934);
or U3320 (N_3320,In_1136,In_1295);
xor U3321 (N_3321,In_518,In_250);
and U3322 (N_3322,In_1526,In_1570);
and U3323 (N_3323,In_2651,In_951);
or U3324 (N_3324,In_2895,In_2344);
and U3325 (N_3325,In_544,In_489);
nor U3326 (N_3326,In_2966,In_2002);
or U3327 (N_3327,In_1437,In_555);
and U3328 (N_3328,In_2018,In_205);
or U3329 (N_3329,In_677,In_853);
nor U3330 (N_3330,In_2771,In_1035);
and U3331 (N_3331,In_2312,In_415);
nand U3332 (N_3332,In_1976,In_749);
and U3333 (N_3333,In_1262,In_2138);
and U3334 (N_3334,In_352,In_525);
or U3335 (N_3335,In_127,In_1165);
nand U3336 (N_3336,In_306,In_871);
or U3337 (N_3337,In_2567,In_2505);
nor U3338 (N_3338,In_582,In_577);
or U3339 (N_3339,In_2654,In_2462);
nand U3340 (N_3340,In_1493,In_700);
nand U3341 (N_3341,In_1420,In_2626);
or U3342 (N_3342,In_1020,In_1521);
nor U3343 (N_3343,In_1382,In_1121);
or U3344 (N_3344,In_63,In_2543);
and U3345 (N_3345,In_2165,In_1875);
and U3346 (N_3346,In_2112,In_23);
xnor U3347 (N_3347,In_1858,In_180);
nand U3348 (N_3348,In_233,In_2777);
nand U3349 (N_3349,In_1587,In_1156);
and U3350 (N_3350,In_666,In_1655);
and U3351 (N_3351,In_1106,In_2904);
nand U3352 (N_3352,In_1039,In_2191);
nand U3353 (N_3353,In_1735,In_4);
nor U3354 (N_3354,In_1158,In_741);
and U3355 (N_3355,In_1298,In_620);
or U3356 (N_3356,In_904,In_1005);
or U3357 (N_3357,In_2108,In_268);
or U3358 (N_3358,In_1722,In_878);
nor U3359 (N_3359,In_2786,In_245);
or U3360 (N_3360,In_2143,In_1598);
nand U3361 (N_3361,In_1696,In_1923);
nand U3362 (N_3362,In_182,In_1545);
nand U3363 (N_3363,In_1646,In_1549);
xnor U3364 (N_3364,In_240,In_2302);
nand U3365 (N_3365,In_24,In_792);
nand U3366 (N_3366,In_2093,In_633);
nand U3367 (N_3367,In_2503,In_207);
or U3368 (N_3368,In_614,In_1865);
nor U3369 (N_3369,In_322,In_1215);
and U3370 (N_3370,In_2379,In_223);
xor U3371 (N_3371,In_2095,In_2461);
and U3372 (N_3372,In_2697,In_2583);
and U3373 (N_3373,In_2968,In_817);
nor U3374 (N_3374,In_1525,In_2455);
nor U3375 (N_3375,In_1985,In_1617);
nand U3376 (N_3376,In_87,In_1578);
or U3377 (N_3377,In_2676,In_648);
xor U3378 (N_3378,In_2344,In_1908);
and U3379 (N_3379,In_2333,In_2301);
or U3380 (N_3380,In_2940,In_2176);
and U3381 (N_3381,In_2571,In_2275);
nor U3382 (N_3382,In_2574,In_435);
or U3383 (N_3383,In_1253,In_87);
and U3384 (N_3384,In_2115,In_122);
and U3385 (N_3385,In_2039,In_2900);
xnor U3386 (N_3386,In_297,In_2053);
nor U3387 (N_3387,In_2109,In_115);
nand U3388 (N_3388,In_984,In_1283);
nand U3389 (N_3389,In_2709,In_576);
and U3390 (N_3390,In_2337,In_1966);
or U3391 (N_3391,In_2707,In_1545);
xnor U3392 (N_3392,In_1779,In_521);
or U3393 (N_3393,In_980,In_1904);
nand U3394 (N_3394,In_1090,In_1233);
nor U3395 (N_3395,In_1881,In_2547);
nand U3396 (N_3396,In_319,In_837);
or U3397 (N_3397,In_1968,In_1565);
nand U3398 (N_3398,In_2778,In_966);
nor U3399 (N_3399,In_2076,In_90);
or U3400 (N_3400,In_1027,In_2322);
nor U3401 (N_3401,In_1658,In_1683);
nand U3402 (N_3402,In_693,In_1433);
nand U3403 (N_3403,In_749,In_1143);
or U3404 (N_3404,In_1097,In_1580);
nor U3405 (N_3405,In_1707,In_1750);
nand U3406 (N_3406,In_1278,In_1303);
nor U3407 (N_3407,In_141,In_2151);
or U3408 (N_3408,In_706,In_2155);
nor U3409 (N_3409,In_2077,In_2622);
xnor U3410 (N_3410,In_2284,In_1565);
nand U3411 (N_3411,In_2042,In_242);
nand U3412 (N_3412,In_2428,In_1104);
or U3413 (N_3413,In_800,In_2346);
nor U3414 (N_3414,In_257,In_1670);
xor U3415 (N_3415,In_94,In_2643);
or U3416 (N_3416,In_2498,In_390);
nand U3417 (N_3417,In_230,In_1908);
or U3418 (N_3418,In_8,In_858);
xor U3419 (N_3419,In_2356,In_29);
xnor U3420 (N_3420,In_2922,In_2405);
or U3421 (N_3421,In_1047,In_2192);
or U3422 (N_3422,In_844,In_334);
nand U3423 (N_3423,In_482,In_864);
nand U3424 (N_3424,In_428,In_2382);
or U3425 (N_3425,In_1774,In_63);
nor U3426 (N_3426,In_2478,In_1191);
nor U3427 (N_3427,In_116,In_818);
nor U3428 (N_3428,In_945,In_703);
or U3429 (N_3429,In_558,In_249);
xor U3430 (N_3430,In_2960,In_2943);
and U3431 (N_3431,In_1948,In_2171);
and U3432 (N_3432,In_1483,In_1265);
nand U3433 (N_3433,In_889,In_1311);
and U3434 (N_3434,In_1798,In_2236);
or U3435 (N_3435,In_1488,In_1290);
and U3436 (N_3436,In_981,In_2846);
nor U3437 (N_3437,In_265,In_1493);
nor U3438 (N_3438,In_123,In_856);
nand U3439 (N_3439,In_1008,In_2351);
and U3440 (N_3440,In_1980,In_916);
and U3441 (N_3441,In_871,In_641);
nand U3442 (N_3442,In_2267,In_1325);
and U3443 (N_3443,In_1449,In_239);
or U3444 (N_3444,In_1202,In_1783);
xor U3445 (N_3445,In_2192,In_2885);
and U3446 (N_3446,In_1238,In_1493);
xor U3447 (N_3447,In_1759,In_217);
nor U3448 (N_3448,In_1951,In_1792);
xor U3449 (N_3449,In_1250,In_1564);
nor U3450 (N_3450,In_886,In_1775);
or U3451 (N_3451,In_1505,In_2745);
nor U3452 (N_3452,In_285,In_740);
and U3453 (N_3453,In_651,In_329);
and U3454 (N_3454,In_107,In_1136);
nor U3455 (N_3455,In_1877,In_338);
nor U3456 (N_3456,In_1301,In_1598);
nand U3457 (N_3457,In_1259,In_1616);
and U3458 (N_3458,In_1116,In_753);
nand U3459 (N_3459,In_1607,In_1352);
and U3460 (N_3460,In_488,In_1117);
nor U3461 (N_3461,In_1841,In_832);
or U3462 (N_3462,In_1483,In_2417);
nor U3463 (N_3463,In_117,In_158);
nand U3464 (N_3464,In_1737,In_1559);
nand U3465 (N_3465,In_1872,In_663);
or U3466 (N_3466,In_1552,In_2726);
or U3467 (N_3467,In_1534,In_840);
and U3468 (N_3468,In_1906,In_2610);
xor U3469 (N_3469,In_2148,In_2023);
and U3470 (N_3470,In_188,In_917);
nor U3471 (N_3471,In_2012,In_2611);
and U3472 (N_3472,In_2207,In_1232);
nor U3473 (N_3473,In_290,In_1085);
nor U3474 (N_3474,In_2182,In_1393);
nor U3475 (N_3475,In_1923,In_314);
or U3476 (N_3476,In_1382,In_1334);
and U3477 (N_3477,In_2329,In_715);
and U3478 (N_3478,In_1701,In_1394);
nand U3479 (N_3479,In_162,In_130);
nor U3480 (N_3480,In_863,In_1948);
and U3481 (N_3481,In_1022,In_718);
and U3482 (N_3482,In_1873,In_643);
or U3483 (N_3483,In_125,In_1430);
and U3484 (N_3484,In_2236,In_2696);
and U3485 (N_3485,In_2080,In_169);
or U3486 (N_3486,In_1644,In_726);
xnor U3487 (N_3487,In_183,In_462);
or U3488 (N_3488,In_2983,In_1250);
nand U3489 (N_3489,In_613,In_1533);
or U3490 (N_3490,In_829,In_821);
nand U3491 (N_3491,In_2735,In_1004);
xnor U3492 (N_3492,In_238,In_535);
and U3493 (N_3493,In_167,In_2397);
and U3494 (N_3494,In_1167,In_1733);
and U3495 (N_3495,In_2026,In_563);
nor U3496 (N_3496,In_1568,In_2606);
and U3497 (N_3497,In_2380,In_2788);
nand U3498 (N_3498,In_1352,In_1609);
or U3499 (N_3499,In_2774,In_1689);
and U3500 (N_3500,In_2191,In_2829);
or U3501 (N_3501,In_1009,In_2227);
nor U3502 (N_3502,In_26,In_2661);
xor U3503 (N_3503,In_2914,In_2772);
xnor U3504 (N_3504,In_1609,In_2077);
xnor U3505 (N_3505,In_583,In_912);
nand U3506 (N_3506,In_26,In_2818);
or U3507 (N_3507,In_1028,In_2670);
nand U3508 (N_3508,In_1165,In_1402);
nand U3509 (N_3509,In_1657,In_1313);
and U3510 (N_3510,In_1757,In_525);
nand U3511 (N_3511,In_1791,In_2824);
nor U3512 (N_3512,In_185,In_2380);
nand U3513 (N_3513,In_1647,In_1184);
nand U3514 (N_3514,In_317,In_2689);
or U3515 (N_3515,In_2410,In_125);
or U3516 (N_3516,In_1106,In_1195);
or U3517 (N_3517,In_2019,In_1600);
nand U3518 (N_3518,In_1387,In_2524);
nor U3519 (N_3519,In_2983,In_193);
nand U3520 (N_3520,In_141,In_137);
and U3521 (N_3521,In_2668,In_1739);
and U3522 (N_3522,In_2514,In_1877);
nor U3523 (N_3523,In_1106,In_2922);
or U3524 (N_3524,In_1134,In_1397);
nor U3525 (N_3525,In_1685,In_915);
xnor U3526 (N_3526,In_2733,In_2842);
nor U3527 (N_3527,In_187,In_2739);
nand U3528 (N_3528,In_279,In_389);
nor U3529 (N_3529,In_841,In_1662);
and U3530 (N_3530,In_2610,In_1917);
or U3531 (N_3531,In_2799,In_2148);
and U3532 (N_3532,In_243,In_641);
nor U3533 (N_3533,In_1534,In_326);
nand U3534 (N_3534,In_1339,In_1819);
or U3535 (N_3535,In_1777,In_2590);
or U3536 (N_3536,In_636,In_2939);
and U3537 (N_3537,In_2473,In_2848);
or U3538 (N_3538,In_99,In_1849);
nor U3539 (N_3539,In_2760,In_10);
nand U3540 (N_3540,In_153,In_1552);
or U3541 (N_3541,In_2336,In_2762);
and U3542 (N_3542,In_1269,In_2870);
nand U3543 (N_3543,In_1116,In_1277);
and U3544 (N_3544,In_2489,In_60);
nand U3545 (N_3545,In_2922,In_1579);
and U3546 (N_3546,In_1152,In_72);
and U3547 (N_3547,In_577,In_1520);
or U3548 (N_3548,In_2390,In_2914);
or U3549 (N_3549,In_1121,In_2417);
nor U3550 (N_3550,In_2905,In_42);
nand U3551 (N_3551,In_2989,In_1850);
nand U3552 (N_3552,In_1799,In_211);
or U3553 (N_3553,In_1903,In_1464);
xnor U3554 (N_3554,In_503,In_804);
nor U3555 (N_3555,In_1917,In_1868);
nand U3556 (N_3556,In_859,In_1377);
nor U3557 (N_3557,In_1573,In_402);
nand U3558 (N_3558,In_2072,In_919);
and U3559 (N_3559,In_2518,In_2244);
xnor U3560 (N_3560,In_1439,In_18);
nand U3561 (N_3561,In_574,In_2525);
nand U3562 (N_3562,In_2566,In_268);
and U3563 (N_3563,In_910,In_1167);
or U3564 (N_3564,In_1619,In_2019);
and U3565 (N_3565,In_262,In_984);
or U3566 (N_3566,In_1520,In_614);
and U3567 (N_3567,In_2382,In_617);
and U3568 (N_3568,In_2841,In_542);
nand U3569 (N_3569,In_597,In_558);
or U3570 (N_3570,In_2756,In_463);
and U3571 (N_3571,In_38,In_1108);
xnor U3572 (N_3572,In_548,In_929);
and U3573 (N_3573,In_1651,In_383);
nand U3574 (N_3574,In_2395,In_103);
xnor U3575 (N_3575,In_748,In_1065);
and U3576 (N_3576,In_597,In_1815);
or U3577 (N_3577,In_149,In_2466);
or U3578 (N_3578,In_1998,In_885);
nor U3579 (N_3579,In_753,In_1813);
or U3580 (N_3580,In_607,In_518);
and U3581 (N_3581,In_918,In_1344);
and U3582 (N_3582,In_2890,In_922);
xor U3583 (N_3583,In_1203,In_946);
or U3584 (N_3584,In_1185,In_2708);
or U3585 (N_3585,In_273,In_538);
xor U3586 (N_3586,In_348,In_2621);
nor U3587 (N_3587,In_954,In_1908);
nor U3588 (N_3588,In_2845,In_2763);
nor U3589 (N_3589,In_2849,In_242);
nand U3590 (N_3590,In_56,In_1321);
nand U3591 (N_3591,In_1350,In_382);
or U3592 (N_3592,In_966,In_2507);
xnor U3593 (N_3593,In_1193,In_819);
or U3594 (N_3594,In_462,In_626);
nand U3595 (N_3595,In_887,In_2551);
or U3596 (N_3596,In_473,In_766);
nor U3597 (N_3597,In_1239,In_2677);
nand U3598 (N_3598,In_304,In_1998);
xor U3599 (N_3599,In_2374,In_941);
or U3600 (N_3600,In_2958,In_365);
nor U3601 (N_3601,In_680,In_1897);
nand U3602 (N_3602,In_2392,In_534);
xor U3603 (N_3603,In_1785,In_2495);
nand U3604 (N_3604,In_2171,In_434);
or U3605 (N_3605,In_227,In_926);
or U3606 (N_3606,In_1994,In_592);
nand U3607 (N_3607,In_2386,In_1714);
and U3608 (N_3608,In_1661,In_1525);
xnor U3609 (N_3609,In_82,In_290);
and U3610 (N_3610,In_95,In_2597);
or U3611 (N_3611,In_1492,In_456);
and U3612 (N_3612,In_782,In_2114);
nand U3613 (N_3613,In_255,In_2166);
and U3614 (N_3614,In_726,In_1843);
or U3615 (N_3615,In_734,In_2181);
xnor U3616 (N_3616,In_876,In_558);
nor U3617 (N_3617,In_128,In_1231);
and U3618 (N_3618,In_979,In_1312);
and U3619 (N_3619,In_1177,In_1175);
nor U3620 (N_3620,In_1687,In_1359);
nand U3621 (N_3621,In_748,In_675);
and U3622 (N_3622,In_640,In_1526);
xnor U3623 (N_3623,In_1426,In_1397);
and U3624 (N_3624,In_2949,In_1513);
or U3625 (N_3625,In_894,In_1730);
nor U3626 (N_3626,In_1802,In_541);
nand U3627 (N_3627,In_948,In_2046);
or U3628 (N_3628,In_1849,In_1898);
and U3629 (N_3629,In_16,In_1895);
or U3630 (N_3630,In_1482,In_1896);
nand U3631 (N_3631,In_698,In_377);
nor U3632 (N_3632,In_1570,In_1380);
nand U3633 (N_3633,In_1336,In_2375);
nor U3634 (N_3634,In_1175,In_422);
nor U3635 (N_3635,In_2958,In_1839);
nor U3636 (N_3636,In_785,In_2019);
nand U3637 (N_3637,In_1405,In_2857);
nand U3638 (N_3638,In_2336,In_1280);
xor U3639 (N_3639,In_1238,In_1438);
or U3640 (N_3640,In_997,In_1489);
and U3641 (N_3641,In_1769,In_2330);
nor U3642 (N_3642,In_785,In_1606);
or U3643 (N_3643,In_2762,In_2311);
or U3644 (N_3644,In_2760,In_742);
xnor U3645 (N_3645,In_1123,In_2282);
xnor U3646 (N_3646,In_2852,In_1769);
nor U3647 (N_3647,In_1145,In_2198);
or U3648 (N_3648,In_920,In_2596);
nor U3649 (N_3649,In_1841,In_398);
nor U3650 (N_3650,In_303,In_2764);
xor U3651 (N_3651,In_833,In_2694);
nor U3652 (N_3652,In_2394,In_2835);
or U3653 (N_3653,In_2713,In_693);
nand U3654 (N_3654,In_2294,In_411);
nand U3655 (N_3655,In_201,In_1073);
and U3656 (N_3656,In_1853,In_1780);
or U3657 (N_3657,In_2828,In_884);
xor U3658 (N_3658,In_2444,In_866);
nand U3659 (N_3659,In_153,In_2394);
and U3660 (N_3660,In_2445,In_2479);
nand U3661 (N_3661,In_936,In_2161);
nand U3662 (N_3662,In_665,In_2366);
and U3663 (N_3663,In_782,In_1066);
nand U3664 (N_3664,In_59,In_512);
and U3665 (N_3665,In_2121,In_1429);
and U3666 (N_3666,In_390,In_2830);
or U3667 (N_3667,In_1270,In_2195);
or U3668 (N_3668,In_1197,In_1281);
nor U3669 (N_3669,In_22,In_310);
xor U3670 (N_3670,In_1995,In_1090);
nor U3671 (N_3671,In_662,In_2979);
and U3672 (N_3672,In_1467,In_1480);
nor U3673 (N_3673,In_2970,In_1878);
xor U3674 (N_3674,In_885,In_1302);
and U3675 (N_3675,In_804,In_1892);
or U3676 (N_3676,In_1301,In_2107);
and U3677 (N_3677,In_2544,In_800);
nand U3678 (N_3678,In_2281,In_2647);
or U3679 (N_3679,In_2902,In_1624);
nand U3680 (N_3680,In_1582,In_1304);
and U3681 (N_3681,In_1515,In_450);
and U3682 (N_3682,In_597,In_2431);
nor U3683 (N_3683,In_2972,In_2715);
nor U3684 (N_3684,In_296,In_1450);
nand U3685 (N_3685,In_65,In_1747);
or U3686 (N_3686,In_1566,In_19);
nand U3687 (N_3687,In_75,In_553);
and U3688 (N_3688,In_287,In_1793);
nor U3689 (N_3689,In_935,In_1134);
or U3690 (N_3690,In_1460,In_1179);
nand U3691 (N_3691,In_975,In_614);
xnor U3692 (N_3692,In_371,In_1347);
or U3693 (N_3693,In_2012,In_587);
nor U3694 (N_3694,In_1517,In_1395);
or U3695 (N_3695,In_739,In_1566);
or U3696 (N_3696,In_112,In_2116);
or U3697 (N_3697,In_1074,In_1517);
nor U3698 (N_3698,In_2391,In_1482);
or U3699 (N_3699,In_2278,In_951);
and U3700 (N_3700,In_2764,In_627);
nand U3701 (N_3701,In_588,In_762);
xor U3702 (N_3702,In_19,In_192);
xnor U3703 (N_3703,In_2072,In_2591);
nand U3704 (N_3704,In_1773,In_74);
nand U3705 (N_3705,In_2138,In_314);
and U3706 (N_3706,In_1501,In_849);
xnor U3707 (N_3707,In_976,In_1354);
xor U3708 (N_3708,In_434,In_1930);
nor U3709 (N_3709,In_1408,In_541);
nand U3710 (N_3710,In_1810,In_736);
nor U3711 (N_3711,In_1460,In_2657);
nand U3712 (N_3712,In_2931,In_427);
or U3713 (N_3713,In_2835,In_387);
nor U3714 (N_3714,In_2576,In_80);
nand U3715 (N_3715,In_2962,In_2987);
nand U3716 (N_3716,In_2105,In_827);
and U3717 (N_3717,In_2898,In_1941);
or U3718 (N_3718,In_610,In_1847);
or U3719 (N_3719,In_2575,In_2021);
nor U3720 (N_3720,In_986,In_942);
nand U3721 (N_3721,In_490,In_1545);
or U3722 (N_3722,In_1951,In_1005);
xnor U3723 (N_3723,In_1550,In_1169);
xor U3724 (N_3724,In_539,In_491);
or U3725 (N_3725,In_2013,In_674);
nand U3726 (N_3726,In_2120,In_2512);
and U3727 (N_3727,In_2541,In_1502);
and U3728 (N_3728,In_1003,In_2075);
nor U3729 (N_3729,In_2875,In_273);
or U3730 (N_3730,In_1380,In_2914);
nand U3731 (N_3731,In_826,In_2244);
nor U3732 (N_3732,In_325,In_1578);
or U3733 (N_3733,In_525,In_581);
or U3734 (N_3734,In_1810,In_2552);
nand U3735 (N_3735,In_682,In_1675);
and U3736 (N_3736,In_1928,In_2578);
and U3737 (N_3737,In_2527,In_695);
or U3738 (N_3738,In_1466,In_1549);
and U3739 (N_3739,In_1136,In_2309);
xor U3740 (N_3740,In_2096,In_2103);
or U3741 (N_3741,In_989,In_1196);
and U3742 (N_3742,In_372,In_644);
nand U3743 (N_3743,In_1187,In_879);
nand U3744 (N_3744,In_1572,In_306);
nor U3745 (N_3745,In_2788,In_313);
nor U3746 (N_3746,In_1750,In_257);
nand U3747 (N_3747,In_1082,In_1624);
and U3748 (N_3748,In_253,In_2986);
and U3749 (N_3749,In_323,In_2684);
or U3750 (N_3750,In_321,In_908);
and U3751 (N_3751,In_1360,In_1945);
xnor U3752 (N_3752,In_1012,In_782);
nand U3753 (N_3753,In_1863,In_2156);
nand U3754 (N_3754,In_2939,In_1910);
nor U3755 (N_3755,In_2829,In_1450);
xor U3756 (N_3756,In_1055,In_2390);
and U3757 (N_3757,In_2258,In_2436);
nand U3758 (N_3758,In_402,In_2949);
and U3759 (N_3759,In_1569,In_1730);
or U3760 (N_3760,In_2418,In_1550);
or U3761 (N_3761,In_1195,In_522);
and U3762 (N_3762,In_2082,In_1150);
nand U3763 (N_3763,In_2973,In_2741);
and U3764 (N_3764,In_1515,In_2755);
or U3765 (N_3765,In_1458,In_317);
or U3766 (N_3766,In_89,In_2304);
xnor U3767 (N_3767,In_759,In_500);
nand U3768 (N_3768,In_149,In_1041);
or U3769 (N_3769,In_1466,In_453);
xor U3770 (N_3770,In_1365,In_2643);
nand U3771 (N_3771,In_968,In_1022);
nand U3772 (N_3772,In_2327,In_605);
and U3773 (N_3773,In_284,In_2256);
or U3774 (N_3774,In_1642,In_2755);
nand U3775 (N_3775,In_1465,In_1204);
nand U3776 (N_3776,In_2103,In_2082);
or U3777 (N_3777,In_1981,In_2573);
and U3778 (N_3778,In_555,In_1090);
and U3779 (N_3779,In_2910,In_792);
nor U3780 (N_3780,In_2282,In_999);
nor U3781 (N_3781,In_2205,In_2106);
nand U3782 (N_3782,In_1005,In_710);
xnor U3783 (N_3783,In_2704,In_2999);
nand U3784 (N_3784,In_2003,In_1235);
nor U3785 (N_3785,In_559,In_2019);
nand U3786 (N_3786,In_1839,In_2980);
nor U3787 (N_3787,In_1803,In_1728);
nor U3788 (N_3788,In_1003,In_1448);
nor U3789 (N_3789,In_2027,In_125);
nand U3790 (N_3790,In_2595,In_682);
nor U3791 (N_3791,In_698,In_2119);
or U3792 (N_3792,In_77,In_2044);
xnor U3793 (N_3793,In_1348,In_1354);
and U3794 (N_3794,In_95,In_2496);
and U3795 (N_3795,In_221,In_2207);
and U3796 (N_3796,In_2543,In_605);
or U3797 (N_3797,In_1380,In_2318);
and U3798 (N_3798,In_2780,In_2579);
nand U3799 (N_3799,In_1250,In_2006);
or U3800 (N_3800,In_651,In_2636);
nand U3801 (N_3801,In_2509,In_2224);
nor U3802 (N_3802,In_2837,In_2560);
nand U3803 (N_3803,In_274,In_1949);
nand U3804 (N_3804,In_1807,In_1799);
nand U3805 (N_3805,In_2778,In_2303);
and U3806 (N_3806,In_173,In_1210);
nand U3807 (N_3807,In_2554,In_2747);
or U3808 (N_3808,In_1082,In_2463);
and U3809 (N_3809,In_1536,In_859);
nor U3810 (N_3810,In_72,In_897);
or U3811 (N_3811,In_18,In_2444);
nor U3812 (N_3812,In_1351,In_226);
nor U3813 (N_3813,In_2942,In_2703);
or U3814 (N_3814,In_2561,In_2640);
nor U3815 (N_3815,In_219,In_2355);
nor U3816 (N_3816,In_2428,In_1113);
and U3817 (N_3817,In_132,In_2394);
or U3818 (N_3818,In_749,In_1866);
or U3819 (N_3819,In_2192,In_1126);
xor U3820 (N_3820,In_2872,In_1446);
nor U3821 (N_3821,In_1683,In_78);
nand U3822 (N_3822,In_1516,In_2316);
nand U3823 (N_3823,In_642,In_1290);
nand U3824 (N_3824,In_1002,In_2298);
nor U3825 (N_3825,In_2769,In_2892);
nor U3826 (N_3826,In_2582,In_1409);
nand U3827 (N_3827,In_1115,In_2691);
nand U3828 (N_3828,In_11,In_2727);
or U3829 (N_3829,In_1156,In_1880);
or U3830 (N_3830,In_2584,In_673);
and U3831 (N_3831,In_275,In_536);
or U3832 (N_3832,In_2338,In_1148);
nor U3833 (N_3833,In_1571,In_2064);
and U3834 (N_3834,In_498,In_661);
nand U3835 (N_3835,In_1325,In_2105);
xnor U3836 (N_3836,In_2329,In_381);
and U3837 (N_3837,In_2179,In_1297);
or U3838 (N_3838,In_2785,In_1468);
and U3839 (N_3839,In_489,In_372);
or U3840 (N_3840,In_2863,In_1633);
and U3841 (N_3841,In_1772,In_457);
or U3842 (N_3842,In_485,In_932);
and U3843 (N_3843,In_1963,In_2987);
nor U3844 (N_3844,In_2336,In_238);
nand U3845 (N_3845,In_408,In_1313);
nand U3846 (N_3846,In_763,In_2081);
nand U3847 (N_3847,In_2549,In_1385);
nor U3848 (N_3848,In_634,In_2706);
and U3849 (N_3849,In_2112,In_2609);
xnor U3850 (N_3850,In_2468,In_1725);
or U3851 (N_3851,In_1346,In_1222);
nor U3852 (N_3852,In_1573,In_2521);
nand U3853 (N_3853,In_2399,In_347);
xor U3854 (N_3854,In_1491,In_792);
or U3855 (N_3855,In_471,In_2989);
nand U3856 (N_3856,In_373,In_1294);
nand U3857 (N_3857,In_1337,In_358);
nor U3858 (N_3858,In_144,In_2197);
nor U3859 (N_3859,In_2144,In_2136);
nor U3860 (N_3860,In_1350,In_2464);
or U3861 (N_3861,In_748,In_199);
and U3862 (N_3862,In_2169,In_1494);
and U3863 (N_3863,In_1573,In_2367);
nand U3864 (N_3864,In_981,In_193);
xnor U3865 (N_3865,In_1359,In_1269);
nor U3866 (N_3866,In_393,In_570);
nor U3867 (N_3867,In_2466,In_680);
nor U3868 (N_3868,In_902,In_25);
nor U3869 (N_3869,In_1226,In_1416);
and U3870 (N_3870,In_710,In_1389);
or U3871 (N_3871,In_2388,In_923);
xnor U3872 (N_3872,In_2967,In_2082);
and U3873 (N_3873,In_203,In_1722);
nand U3874 (N_3874,In_2571,In_1446);
and U3875 (N_3875,In_1398,In_1137);
nand U3876 (N_3876,In_878,In_1666);
and U3877 (N_3877,In_932,In_166);
nor U3878 (N_3878,In_241,In_527);
nand U3879 (N_3879,In_1444,In_2694);
nand U3880 (N_3880,In_1252,In_83);
or U3881 (N_3881,In_238,In_389);
and U3882 (N_3882,In_1470,In_956);
nand U3883 (N_3883,In_2895,In_2699);
nor U3884 (N_3884,In_312,In_2081);
xor U3885 (N_3885,In_2266,In_1741);
nor U3886 (N_3886,In_522,In_2664);
nor U3887 (N_3887,In_273,In_2681);
or U3888 (N_3888,In_623,In_2759);
nor U3889 (N_3889,In_2663,In_2024);
or U3890 (N_3890,In_1179,In_2576);
and U3891 (N_3891,In_213,In_1088);
and U3892 (N_3892,In_17,In_202);
xnor U3893 (N_3893,In_384,In_2415);
or U3894 (N_3894,In_1201,In_1125);
nand U3895 (N_3895,In_44,In_429);
and U3896 (N_3896,In_1008,In_1857);
nor U3897 (N_3897,In_982,In_1045);
and U3898 (N_3898,In_2963,In_108);
and U3899 (N_3899,In_2127,In_392);
or U3900 (N_3900,In_1039,In_376);
or U3901 (N_3901,In_2109,In_2320);
and U3902 (N_3902,In_302,In_2937);
nand U3903 (N_3903,In_2302,In_796);
nor U3904 (N_3904,In_432,In_865);
or U3905 (N_3905,In_726,In_2558);
or U3906 (N_3906,In_662,In_2191);
or U3907 (N_3907,In_1835,In_1096);
and U3908 (N_3908,In_1406,In_803);
nand U3909 (N_3909,In_2711,In_954);
and U3910 (N_3910,In_898,In_2388);
nor U3911 (N_3911,In_2724,In_2765);
or U3912 (N_3912,In_131,In_2677);
nand U3913 (N_3913,In_2725,In_120);
and U3914 (N_3914,In_1450,In_2567);
and U3915 (N_3915,In_1559,In_2742);
nand U3916 (N_3916,In_1403,In_1482);
xnor U3917 (N_3917,In_1446,In_1069);
xor U3918 (N_3918,In_371,In_2506);
nor U3919 (N_3919,In_1967,In_2908);
nand U3920 (N_3920,In_1317,In_894);
nor U3921 (N_3921,In_2624,In_458);
and U3922 (N_3922,In_1367,In_865);
nand U3923 (N_3923,In_2478,In_2716);
nand U3924 (N_3924,In_2478,In_1884);
nor U3925 (N_3925,In_30,In_2793);
or U3926 (N_3926,In_2614,In_1199);
nor U3927 (N_3927,In_959,In_2995);
xnor U3928 (N_3928,In_2636,In_951);
nand U3929 (N_3929,In_1313,In_1169);
and U3930 (N_3930,In_11,In_1532);
nand U3931 (N_3931,In_2199,In_2865);
and U3932 (N_3932,In_1301,In_346);
nand U3933 (N_3933,In_68,In_255);
xnor U3934 (N_3934,In_1949,In_1997);
and U3935 (N_3935,In_1455,In_1582);
nor U3936 (N_3936,In_2884,In_2788);
nor U3937 (N_3937,In_1913,In_2562);
nand U3938 (N_3938,In_2601,In_922);
nand U3939 (N_3939,In_2955,In_1412);
nand U3940 (N_3940,In_2245,In_863);
nand U3941 (N_3941,In_2874,In_1264);
or U3942 (N_3942,In_1896,In_1871);
or U3943 (N_3943,In_1493,In_1872);
or U3944 (N_3944,In_280,In_2464);
xor U3945 (N_3945,In_2415,In_2890);
nand U3946 (N_3946,In_2059,In_512);
and U3947 (N_3947,In_1279,In_2054);
nor U3948 (N_3948,In_1515,In_2839);
nand U3949 (N_3949,In_1116,In_1571);
and U3950 (N_3950,In_1365,In_721);
nor U3951 (N_3951,In_1619,In_1197);
or U3952 (N_3952,In_1722,In_1637);
and U3953 (N_3953,In_387,In_1204);
nor U3954 (N_3954,In_2371,In_199);
and U3955 (N_3955,In_2617,In_2779);
or U3956 (N_3956,In_1388,In_2887);
or U3957 (N_3957,In_2606,In_423);
nand U3958 (N_3958,In_1345,In_816);
nand U3959 (N_3959,In_1516,In_147);
nand U3960 (N_3960,In_444,In_2845);
or U3961 (N_3961,In_1353,In_86);
nand U3962 (N_3962,In_399,In_2453);
or U3963 (N_3963,In_518,In_2012);
xor U3964 (N_3964,In_1912,In_1259);
and U3965 (N_3965,In_1699,In_2278);
xnor U3966 (N_3966,In_1613,In_926);
and U3967 (N_3967,In_548,In_849);
xnor U3968 (N_3968,In_58,In_1029);
nor U3969 (N_3969,In_2919,In_2724);
or U3970 (N_3970,In_517,In_133);
and U3971 (N_3971,In_596,In_1694);
or U3972 (N_3972,In_658,In_2717);
nand U3973 (N_3973,In_991,In_1518);
and U3974 (N_3974,In_2045,In_79);
or U3975 (N_3975,In_1243,In_2588);
and U3976 (N_3976,In_2111,In_2090);
or U3977 (N_3977,In_894,In_1879);
and U3978 (N_3978,In_2613,In_2490);
or U3979 (N_3979,In_2769,In_1665);
xor U3980 (N_3980,In_424,In_2690);
xnor U3981 (N_3981,In_35,In_2311);
xor U3982 (N_3982,In_675,In_742);
and U3983 (N_3983,In_2810,In_2890);
and U3984 (N_3984,In_854,In_874);
nor U3985 (N_3985,In_1818,In_731);
or U3986 (N_3986,In_2952,In_2791);
and U3987 (N_3987,In_2461,In_2584);
or U3988 (N_3988,In_104,In_503);
or U3989 (N_3989,In_2744,In_1060);
nand U3990 (N_3990,In_2893,In_2109);
nor U3991 (N_3991,In_526,In_2168);
or U3992 (N_3992,In_1541,In_2484);
nor U3993 (N_3993,In_143,In_666);
nor U3994 (N_3994,In_2818,In_2954);
nand U3995 (N_3995,In_1587,In_1909);
and U3996 (N_3996,In_2517,In_923);
nor U3997 (N_3997,In_1602,In_135);
nor U3998 (N_3998,In_1732,In_2193);
and U3999 (N_3999,In_2608,In_2865);
nand U4000 (N_4000,In_106,In_1629);
and U4001 (N_4001,In_2536,In_1006);
and U4002 (N_4002,In_353,In_1813);
nor U4003 (N_4003,In_2736,In_355);
nand U4004 (N_4004,In_251,In_2996);
and U4005 (N_4005,In_2153,In_2509);
nor U4006 (N_4006,In_1213,In_1246);
nand U4007 (N_4007,In_1655,In_923);
xnor U4008 (N_4008,In_451,In_1016);
or U4009 (N_4009,In_2711,In_1154);
nor U4010 (N_4010,In_565,In_1291);
nor U4011 (N_4011,In_2868,In_478);
and U4012 (N_4012,In_409,In_918);
nand U4013 (N_4013,In_1389,In_922);
xor U4014 (N_4014,In_125,In_1019);
xnor U4015 (N_4015,In_693,In_1670);
xnor U4016 (N_4016,In_2287,In_2405);
or U4017 (N_4017,In_1601,In_2598);
xor U4018 (N_4018,In_1492,In_2409);
nand U4019 (N_4019,In_221,In_2997);
xor U4020 (N_4020,In_436,In_1489);
nand U4021 (N_4021,In_1308,In_1652);
nand U4022 (N_4022,In_286,In_1180);
and U4023 (N_4023,In_1969,In_477);
nor U4024 (N_4024,In_2342,In_2523);
or U4025 (N_4025,In_1788,In_2202);
and U4026 (N_4026,In_628,In_2137);
and U4027 (N_4027,In_1666,In_2196);
nor U4028 (N_4028,In_942,In_2805);
or U4029 (N_4029,In_517,In_915);
or U4030 (N_4030,In_2375,In_1618);
or U4031 (N_4031,In_166,In_1591);
xnor U4032 (N_4032,In_2003,In_1055);
and U4033 (N_4033,In_1948,In_994);
and U4034 (N_4034,In_1303,In_323);
nor U4035 (N_4035,In_155,In_577);
or U4036 (N_4036,In_480,In_795);
xor U4037 (N_4037,In_814,In_2836);
nor U4038 (N_4038,In_389,In_1426);
and U4039 (N_4039,In_45,In_2051);
nand U4040 (N_4040,In_484,In_326);
nand U4041 (N_4041,In_1119,In_1498);
and U4042 (N_4042,In_453,In_296);
nor U4043 (N_4043,In_36,In_1965);
nor U4044 (N_4044,In_1214,In_268);
and U4045 (N_4045,In_1769,In_1654);
nand U4046 (N_4046,In_595,In_1218);
and U4047 (N_4047,In_2797,In_1892);
and U4048 (N_4048,In_2072,In_2684);
and U4049 (N_4049,In_2983,In_1943);
and U4050 (N_4050,In_1276,In_415);
or U4051 (N_4051,In_233,In_745);
or U4052 (N_4052,In_1683,In_826);
nor U4053 (N_4053,In_2545,In_2586);
xor U4054 (N_4054,In_1756,In_2441);
or U4055 (N_4055,In_207,In_1559);
nand U4056 (N_4056,In_1768,In_1841);
and U4057 (N_4057,In_1049,In_1406);
xnor U4058 (N_4058,In_264,In_1175);
nand U4059 (N_4059,In_1578,In_1956);
nand U4060 (N_4060,In_2002,In_2936);
nand U4061 (N_4061,In_1642,In_1803);
nor U4062 (N_4062,In_704,In_1216);
nand U4063 (N_4063,In_1924,In_1059);
nand U4064 (N_4064,In_2492,In_568);
or U4065 (N_4065,In_320,In_1479);
and U4066 (N_4066,In_2335,In_2763);
nor U4067 (N_4067,In_398,In_1445);
nor U4068 (N_4068,In_1926,In_2382);
or U4069 (N_4069,In_801,In_2010);
xor U4070 (N_4070,In_1151,In_2186);
nor U4071 (N_4071,In_2731,In_2895);
nand U4072 (N_4072,In_801,In_1970);
or U4073 (N_4073,In_23,In_1704);
nor U4074 (N_4074,In_341,In_1526);
nand U4075 (N_4075,In_1029,In_2618);
nand U4076 (N_4076,In_2089,In_2843);
nand U4077 (N_4077,In_2486,In_331);
or U4078 (N_4078,In_2851,In_1331);
or U4079 (N_4079,In_1319,In_2545);
nor U4080 (N_4080,In_2759,In_2893);
xnor U4081 (N_4081,In_2142,In_1131);
nor U4082 (N_4082,In_1553,In_671);
nand U4083 (N_4083,In_742,In_2330);
and U4084 (N_4084,In_2885,In_897);
nand U4085 (N_4085,In_2551,In_399);
and U4086 (N_4086,In_1263,In_2551);
nand U4087 (N_4087,In_2496,In_1045);
nand U4088 (N_4088,In_2943,In_2918);
nor U4089 (N_4089,In_2248,In_2083);
nor U4090 (N_4090,In_2262,In_263);
nand U4091 (N_4091,In_2276,In_841);
nor U4092 (N_4092,In_2080,In_2840);
nand U4093 (N_4093,In_731,In_47);
and U4094 (N_4094,In_1471,In_1557);
xor U4095 (N_4095,In_1268,In_0);
nand U4096 (N_4096,In_417,In_23);
xnor U4097 (N_4097,In_808,In_2819);
nor U4098 (N_4098,In_1734,In_1264);
and U4099 (N_4099,In_309,In_53);
nand U4100 (N_4100,In_2902,In_980);
nor U4101 (N_4101,In_1168,In_1031);
and U4102 (N_4102,In_2075,In_709);
or U4103 (N_4103,In_569,In_738);
nor U4104 (N_4104,In_2365,In_1087);
nor U4105 (N_4105,In_1573,In_153);
nand U4106 (N_4106,In_2549,In_1831);
nand U4107 (N_4107,In_1268,In_1104);
xor U4108 (N_4108,In_772,In_2484);
nor U4109 (N_4109,In_1576,In_145);
and U4110 (N_4110,In_2990,In_364);
nor U4111 (N_4111,In_670,In_2223);
or U4112 (N_4112,In_356,In_2150);
nor U4113 (N_4113,In_734,In_2367);
and U4114 (N_4114,In_564,In_2962);
nand U4115 (N_4115,In_2461,In_2048);
and U4116 (N_4116,In_2478,In_216);
nand U4117 (N_4117,In_840,In_1059);
nand U4118 (N_4118,In_2815,In_806);
or U4119 (N_4119,In_311,In_2854);
or U4120 (N_4120,In_2591,In_698);
or U4121 (N_4121,In_1676,In_1417);
nand U4122 (N_4122,In_5,In_511);
nand U4123 (N_4123,In_2953,In_1146);
nor U4124 (N_4124,In_2644,In_1659);
or U4125 (N_4125,In_2947,In_2060);
nor U4126 (N_4126,In_80,In_2379);
or U4127 (N_4127,In_2985,In_2511);
or U4128 (N_4128,In_1819,In_2837);
nor U4129 (N_4129,In_2860,In_1881);
nand U4130 (N_4130,In_1687,In_2458);
nand U4131 (N_4131,In_323,In_782);
and U4132 (N_4132,In_379,In_632);
nor U4133 (N_4133,In_749,In_732);
and U4134 (N_4134,In_2330,In_2342);
xor U4135 (N_4135,In_856,In_834);
xor U4136 (N_4136,In_1458,In_1414);
and U4137 (N_4137,In_1020,In_2798);
or U4138 (N_4138,In_451,In_2052);
nand U4139 (N_4139,In_579,In_77);
nor U4140 (N_4140,In_984,In_2286);
and U4141 (N_4141,In_2636,In_497);
or U4142 (N_4142,In_64,In_142);
nor U4143 (N_4143,In_1832,In_2511);
and U4144 (N_4144,In_1784,In_1507);
and U4145 (N_4145,In_1343,In_1487);
nor U4146 (N_4146,In_2481,In_2810);
and U4147 (N_4147,In_603,In_2289);
xor U4148 (N_4148,In_2389,In_1873);
nor U4149 (N_4149,In_1031,In_1638);
nand U4150 (N_4150,In_2077,In_1229);
nand U4151 (N_4151,In_455,In_2645);
and U4152 (N_4152,In_631,In_638);
xnor U4153 (N_4153,In_589,In_1704);
or U4154 (N_4154,In_74,In_875);
nand U4155 (N_4155,In_602,In_1939);
and U4156 (N_4156,In_2145,In_2348);
nand U4157 (N_4157,In_779,In_1532);
nand U4158 (N_4158,In_2187,In_107);
or U4159 (N_4159,In_1581,In_754);
nand U4160 (N_4160,In_2087,In_412);
nor U4161 (N_4161,In_1003,In_920);
nor U4162 (N_4162,In_1275,In_1477);
and U4163 (N_4163,In_2641,In_2830);
and U4164 (N_4164,In_495,In_1116);
or U4165 (N_4165,In_2405,In_131);
or U4166 (N_4166,In_2612,In_218);
nand U4167 (N_4167,In_985,In_389);
nand U4168 (N_4168,In_1739,In_373);
nor U4169 (N_4169,In_1024,In_1698);
nand U4170 (N_4170,In_2768,In_2936);
nor U4171 (N_4171,In_2368,In_2819);
nand U4172 (N_4172,In_1923,In_1288);
and U4173 (N_4173,In_1190,In_2134);
or U4174 (N_4174,In_349,In_1864);
and U4175 (N_4175,In_1905,In_2899);
nor U4176 (N_4176,In_1108,In_2407);
nor U4177 (N_4177,In_638,In_2988);
nand U4178 (N_4178,In_2024,In_1290);
nand U4179 (N_4179,In_1646,In_1245);
nand U4180 (N_4180,In_205,In_42);
nor U4181 (N_4181,In_2948,In_1547);
nand U4182 (N_4182,In_543,In_2108);
nor U4183 (N_4183,In_1774,In_24);
nand U4184 (N_4184,In_291,In_892);
and U4185 (N_4185,In_2065,In_2445);
and U4186 (N_4186,In_375,In_2091);
nand U4187 (N_4187,In_199,In_2099);
nand U4188 (N_4188,In_616,In_517);
nand U4189 (N_4189,In_1199,In_686);
xnor U4190 (N_4190,In_2304,In_2175);
nor U4191 (N_4191,In_1594,In_1589);
or U4192 (N_4192,In_663,In_2981);
nor U4193 (N_4193,In_1763,In_402);
nand U4194 (N_4194,In_1642,In_1936);
nand U4195 (N_4195,In_572,In_985);
and U4196 (N_4196,In_2118,In_470);
and U4197 (N_4197,In_2007,In_1336);
nor U4198 (N_4198,In_2004,In_2840);
nand U4199 (N_4199,In_1350,In_1341);
nor U4200 (N_4200,In_1322,In_2194);
nand U4201 (N_4201,In_732,In_1980);
or U4202 (N_4202,In_2673,In_1906);
nor U4203 (N_4203,In_2273,In_930);
nor U4204 (N_4204,In_5,In_1526);
nor U4205 (N_4205,In_768,In_910);
and U4206 (N_4206,In_1688,In_2908);
and U4207 (N_4207,In_1175,In_456);
or U4208 (N_4208,In_2138,In_1462);
or U4209 (N_4209,In_2194,In_152);
nand U4210 (N_4210,In_2826,In_2849);
xnor U4211 (N_4211,In_687,In_1227);
nand U4212 (N_4212,In_1890,In_929);
xnor U4213 (N_4213,In_2527,In_423);
or U4214 (N_4214,In_122,In_1556);
nand U4215 (N_4215,In_1134,In_2250);
nor U4216 (N_4216,In_2814,In_449);
or U4217 (N_4217,In_735,In_2981);
nor U4218 (N_4218,In_2470,In_2795);
and U4219 (N_4219,In_1323,In_2076);
nand U4220 (N_4220,In_937,In_2394);
nand U4221 (N_4221,In_1905,In_703);
nor U4222 (N_4222,In_2937,In_1178);
or U4223 (N_4223,In_372,In_539);
or U4224 (N_4224,In_1391,In_1328);
xor U4225 (N_4225,In_664,In_2928);
or U4226 (N_4226,In_1921,In_377);
nor U4227 (N_4227,In_2710,In_140);
xor U4228 (N_4228,In_278,In_1603);
xor U4229 (N_4229,In_1534,In_1157);
xor U4230 (N_4230,In_2253,In_849);
or U4231 (N_4231,In_2237,In_1);
or U4232 (N_4232,In_2836,In_1234);
and U4233 (N_4233,In_2851,In_1212);
or U4234 (N_4234,In_2841,In_1570);
or U4235 (N_4235,In_651,In_738);
xor U4236 (N_4236,In_810,In_2137);
or U4237 (N_4237,In_2532,In_2464);
nor U4238 (N_4238,In_1556,In_1744);
or U4239 (N_4239,In_2360,In_2010);
nand U4240 (N_4240,In_1636,In_257);
nand U4241 (N_4241,In_1701,In_279);
nor U4242 (N_4242,In_330,In_1679);
and U4243 (N_4243,In_625,In_2569);
nand U4244 (N_4244,In_833,In_965);
nand U4245 (N_4245,In_165,In_1502);
and U4246 (N_4246,In_2425,In_1008);
nor U4247 (N_4247,In_2894,In_2662);
and U4248 (N_4248,In_709,In_2578);
or U4249 (N_4249,In_841,In_597);
and U4250 (N_4250,In_1172,In_6);
xnor U4251 (N_4251,In_1805,In_1724);
and U4252 (N_4252,In_853,In_2012);
and U4253 (N_4253,In_1650,In_1814);
or U4254 (N_4254,In_514,In_332);
nor U4255 (N_4255,In_1014,In_1557);
xor U4256 (N_4256,In_2247,In_2654);
nor U4257 (N_4257,In_1636,In_1747);
xor U4258 (N_4258,In_765,In_688);
and U4259 (N_4259,In_2828,In_593);
or U4260 (N_4260,In_965,In_1389);
or U4261 (N_4261,In_28,In_455);
or U4262 (N_4262,In_1575,In_1697);
and U4263 (N_4263,In_2561,In_1836);
and U4264 (N_4264,In_2222,In_408);
or U4265 (N_4265,In_2114,In_809);
or U4266 (N_4266,In_1543,In_2919);
nand U4267 (N_4267,In_33,In_226);
nand U4268 (N_4268,In_2126,In_2766);
nand U4269 (N_4269,In_1904,In_949);
or U4270 (N_4270,In_1109,In_317);
nand U4271 (N_4271,In_2396,In_2152);
nand U4272 (N_4272,In_639,In_780);
nor U4273 (N_4273,In_9,In_553);
or U4274 (N_4274,In_290,In_1017);
nand U4275 (N_4275,In_2518,In_1747);
nor U4276 (N_4276,In_376,In_1671);
nand U4277 (N_4277,In_280,In_2010);
nor U4278 (N_4278,In_1297,In_921);
nor U4279 (N_4279,In_44,In_1397);
or U4280 (N_4280,In_108,In_1250);
nor U4281 (N_4281,In_845,In_542);
nand U4282 (N_4282,In_888,In_432);
xnor U4283 (N_4283,In_1841,In_555);
nor U4284 (N_4284,In_2587,In_695);
nand U4285 (N_4285,In_756,In_2648);
nor U4286 (N_4286,In_289,In_2411);
and U4287 (N_4287,In_1142,In_1627);
or U4288 (N_4288,In_2974,In_1112);
and U4289 (N_4289,In_2095,In_2409);
or U4290 (N_4290,In_97,In_2581);
nand U4291 (N_4291,In_601,In_281);
nor U4292 (N_4292,In_271,In_373);
or U4293 (N_4293,In_2515,In_2273);
nand U4294 (N_4294,In_541,In_152);
nor U4295 (N_4295,In_1115,In_945);
or U4296 (N_4296,In_2664,In_1758);
and U4297 (N_4297,In_1815,In_411);
or U4298 (N_4298,In_2621,In_2180);
and U4299 (N_4299,In_1553,In_1987);
nor U4300 (N_4300,In_1130,In_260);
nand U4301 (N_4301,In_1406,In_1436);
nand U4302 (N_4302,In_2933,In_1270);
nand U4303 (N_4303,In_2490,In_2192);
or U4304 (N_4304,In_2021,In_2558);
nor U4305 (N_4305,In_2937,In_2245);
nor U4306 (N_4306,In_1474,In_2638);
nor U4307 (N_4307,In_1970,In_2797);
or U4308 (N_4308,In_2835,In_1029);
nor U4309 (N_4309,In_2712,In_2561);
or U4310 (N_4310,In_556,In_1671);
or U4311 (N_4311,In_400,In_568);
nand U4312 (N_4312,In_1325,In_499);
nor U4313 (N_4313,In_1601,In_2950);
nand U4314 (N_4314,In_592,In_1201);
or U4315 (N_4315,In_2426,In_1322);
and U4316 (N_4316,In_226,In_2493);
and U4317 (N_4317,In_803,In_1521);
nor U4318 (N_4318,In_2941,In_1685);
and U4319 (N_4319,In_1474,In_855);
nand U4320 (N_4320,In_179,In_1152);
nor U4321 (N_4321,In_2837,In_174);
nor U4322 (N_4322,In_2625,In_354);
nor U4323 (N_4323,In_832,In_1009);
and U4324 (N_4324,In_1650,In_842);
nand U4325 (N_4325,In_2744,In_2908);
or U4326 (N_4326,In_1292,In_1628);
nor U4327 (N_4327,In_2208,In_754);
and U4328 (N_4328,In_2696,In_2861);
nor U4329 (N_4329,In_1644,In_1892);
nand U4330 (N_4330,In_716,In_344);
nor U4331 (N_4331,In_71,In_1168);
nand U4332 (N_4332,In_2748,In_513);
and U4333 (N_4333,In_963,In_193);
nor U4334 (N_4334,In_1441,In_792);
nor U4335 (N_4335,In_1894,In_205);
nor U4336 (N_4336,In_34,In_468);
nor U4337 (N_4337,In_2874,In_2782);
nand U4338 (N_4338,In_1005,In_275);
and U4339 (N_4339,In_2290,In_1948);
nor U4340 (N_4340,In_801,In_2059);
nand U4341 (N_4341,In_518,In_2551);
or U4342 (N_4342,In_227,In_759);
nand U4343 (N_4343,In_702,In_2733);
nor U4344 (N_4344,In_699,In_138);
nor U4345 (N_4345,In_1672,In_1662);
nor U4346 (N_4346,In_650,In_1607);
nand U4347 (N_4347,In_798,In_1916);
xor U4348 (N_4348,In_2250,In_953);
or U4349 (N_4349,In_1612,In_2658);
and U4350 (N_4350,In_2501,In_2152);
or U4351 (N_4351,In_808,In_611);
and U4352 (N_4352,In_1358,In_756);
and U4353 (N_4353,In_915,In_1874);
xor U4354 (N_4354,In_1395,In_1276);
or U4355 (N_4355,In_218,In_2864);
or U4356 (N_4356,In_2117,In_2706);
nor U4357 (N_4357,In_730,In_1607);
xor U4358 (N_4358,In_1249,In_133);
and U4359 (N_4359,In_2602,In_1056);
nor U4360 (N_4360,In_789,In_2084);
xnor U4361 (N_4361,In_216,In_419);
xnor U4362 (N_4362,In_2416,In_757);
and U4363 (N_4363,In_1301,In_303);
or U4364 (N_4364,In_605,In_1820);
or U4365 (N_4365,In_1150,In_1764);
nand U4366 (N_4366,In_2986,In_65);
xor U4367 (N_4367,In_792,In_2835);
xnor U4368 (N_4368,In_1384,In_87);
or U4369 (N_4369,In_1119,In_2002);
or U4370 (N_4370,In_683,In_685);
and U4371 (N_4371,In_2935,In_1714);
or U4372 (N_4372,In_369,In_2839);
or U4373 (N_4373,In_813,In_1166);
nand U4374 (N_4374,In_1232,In_233);
xor U4375 (N_4375,In_2665,In_2993);
and U4376 (N_4376,In_2345,In_1956);
and U4377 (N_4377,In_1146,In_2193);
nor U4378 (N_4378,In_2025,In_2469);
or U4379 (N_4379,In_206,In_1638);
nor U4380 (N_4380,In_198,In_2427);
nand U4381 (N_4381,In_167,In_769);
nor U4382 (N_4382,In_153,In_2917);
and U4383 (N_4383,In_2181,In_2245);
nor U4384 (N_4384,In_2591,In_647);
and U4385 (N_4385,In_1030,In_2701);
nor U4386 (N_4386,In_2424,In_215);
nor U4387 (N_4387,In_2946,In_1603);
nand U4388 (N_4388,In_1939,In_1135);
and U4389 (N_4389,In_606,In_2130);
or U4390 (N_4390,In_1463,In_2269);
and U4391 (N_4391,In_1199,In_948);
nand U4392 (N_4392,In_1392,In_930);
nor U4393 (N_4393,In_546,In_454);
nor U4394 (N_4394,In_2146,In_2516);
xor U4395 (N_4395,In_2520,In_218);
nor U4396 (N_4396,In_1932,In_2478);
nand U4397 (N_4397,In_62,In_1335);
and U4398 (N_4398,In_435,In_2031);
nand U4399 (N_4399,In_2425,In_2992);
nand U4400 (N_4400,In_2802,In_476);
and U4401 (N_4401,In_886,In_2460);
or U4402 (N_4402,In_379,In_372);
or U4403 (N_4403,In_1501,In_1030);
and U4404 (N_4404,In_2433,In_2383);
or U4405 (N_4405,In_1915,In_183);
nand U4406 (N_4406,In_291,In_2260);
xnor U4407 (N_4407,In_2808,In_1789);
or U4408 (N_4408,In_231,In_801);
nor U4409 (N_4409,In_101,In_496);
nand U4410 (N_4410,In_1604,In_639);
xnor U4411 (N_4411,In_986,In_1096);
and U4412 (N_4412,In_2386,In_41);
or U4413 (N_4413,In_2061,In_603);
nor U4414 (N_4414,In_568,In_897);
and U4415 (N_4415,In_1490,In_727);
nor U4416 (N_4416,In_2779,In_476);
and U4417 (N_4417,In_1647,In_676);
or U4418 (N_4418,In_1767,In_246);
and U4419 (N_4419,In_1985,In_1377);
and U4420 (N_4420,In_1541,In_1094);
and U4421 (N_4421,In_2039,In_2793);
and U4422 (N_4422,In_918,In_2393);
nand U4423 (N_4423,In_1813,In_1357);
or U4424 (N_4424,In_1080,In_2945);
xnor U4425 (N_4425,In_604,In_227);
nor U4426 (N_4426,In_2627,In_866);
xnor U4427 (N_4427,In_375,In_1027);
or U4428 (N_4428,In_29,In_1870);
or U4429 (N_4429,In_2407,In_2641);
or U4430 (N_4430,In_1927,In_2686);
nand U4431 (N_4431,In_2993,In_1887);
xnor U4432 (N_4432,In_752,In_2070);
xnor U4433 (N_4433,In_1808,In_1293);
xnor U4434 (N_4434,In_1914,In_2893);
nor U4435 (N_4435,In_1754,In_2139);
nand U4436 (N_4436,In_1489,In_783);
nand U4437 (N_4437,In_1376,In_2012);
and U4438 (N_4438,In_1802,In_2720);
or U4439 (N_4439,In_2183,In_1553);
or U4440 (N_4440,In_884,In_2298);
nor U4441 (N_4441,In_452,In_539);
and U4442 (N_4442,In_2566,In_2529);
and U4443 (N_4443,In_1149,In_923);
nand U4444 (N_4444,In_2496,In_706);
and U4445 (N_4445,In_634,In_2461);
and U4446 (N_4446,In_67,In_1056);
and U4447 (N_4447,In_2340,In_45);
and U4448 (N_4448,In_2643,In_1709);
and U4449 (N_4449,In_1020,In_1181);
and U4450 (N_4450,In_746,In_105);
xor U4451 (N_4451,In_878,In_1592);
and U4452 (N_4452,In_404,In_2070);
xor U4453 (N_4453,In_406,In_2342);
and U4454 (N_4454,In_2049,In_2670);
nor U4455 (N_4455,In_2933,In_840);
xor U4456 (N_4456,In_2757,In_1508);
nand U4457 (N_4457,In_2347,In_845);
nand U4458 (N_4458,In_2683,In_1864);
or U4459 (N_4459,In_778,In_1561);
nand U4460 (N_4460,In_1809,In_2474);
and U4461 (N_4461,In_2697,In_517);
or U4462 (N_4462,In_259,In_1572);
or U4463 (N_4463,In_307,In_1720);
nand U4464 (N_4464,In_2303,In_611);
nand U4465 (N_4465,In_2122,In_367);
nand U4466 (N_4466,In_2352,In_956);
and U4467 (N_4467,In_1598,In_194);
xor U4468 (N_4468,In_1233,In_1092);
nor U4469 (N_4469,In_823,In_2668);
or U4470 (N_4470,In_1127,In_460);
and U4471 (N_4471,In_1478,In_1028);
nor U4472 (N_4472,In_2532,In_2911);
nand U4473 (N_4473,In_1593,In_2969);
nor U4474 (N_4474,In_2671,In_2261);
and U4475 (N_4475,In_681,In_1358);
nand U4476 (N_4476,In_94,In_2303);
or U4477 (N_4477,In_2882,In_1172);
and U4478 (N_4478,In_1072,In_2795);
nor U4479 (N_4479,In_131,In_723);
nand U4480 (N_4480,In_2842,In_2709);
nor U4481 (N_4481,In_2933,In_274);
and U4482 (N_4482,In_1138,In_2998);
and U4483 (N_4483,In_1776,In_1759);
or U4484 (N_4484,In_2731,In_2669);
nor U4485 (N_4485,In_1688,In_1110);
nor U4486 (N_4486,In_1644,In_1846);
nor U4487 (N_4487,In_1868,In_2780);
and U4488 (N_4488,In_1519,In_1261);
xor U4489 (N_4489,In_595,In_2051);
nand U4490 (N_4490,In_2680,In_774);
or U4491 (N_4491,In_2801,In_2758);
or U4492 (N_4492,In_229,In_1840);
or U4493 (N_4493,In_1522,In_831);
nand U4494 (N_4494,In_2594,In_2313);
nor U4495 (N_4495,In_666,In_1705);
or U4496 (N_4496,In_1934,In_118);
nand U4497 (N_4497,In_708,In_964);
and U4498 (N_4498,In_1902,In_2577);
or U4499 (N_4499,In_851,In_1350);
nand U4500 (N_4500,In_751,In_385);
and U4501 (N_4501,In_2613,In_1158);
nor U4502 (N_4502,In_731,In_1513);
or U4503 (N_4503,In_2451,In_1585);
nor U4504 (N_4504,In_995,In_921);
or U4505 (N_4505,In_1298,In_2767);
nand U4506 (N_4506,In_2969,In_2861);
nor U4507 (N_4507,In_663,In_841);
xor U4508 (N_4508,In_792,In_2359);
and U4509 (N_4509,In_2236,In_2924);
and U4510 (N_4510,In_1719,In_2407);
and U4511 (N_4511,In_2511,In_1756);
nor U4512 (N_4512,In_1446,In_1369);
nor U4513 (N_4513,In_572,In_1278);
nor U4514 (N_4514,In_188,In_2622);
and U4515 (N_4515,In_2350,In_2510);
nor U4516 (N_4516,In_2017,In_2229);
nor U4517 (N_4517,In_2417,In_2128);
nor U4518 (N_4518,In_1007,In_1235);
nor U4519 (N_4519,In_398,In_1355);
xor U4520 (N_4520,In_792,In_1060);
and U4521 (N_4521,In_590,In_2659);
and U4522 (N_4522,In_1975,In_2895);
or U4523 (N_4523,In_1680,In_2257);
nor U4524 (N_4524,In_1362,In_1777);
xor U4525 (N_4525,In_898,In_2603);
nand U4526 (N_4526,In_1855,In_1590);
or U4527 (N_4527,In_1988,In_442);
nor U4528 (N_4528,In_1245,In_2402);
or U4529 (N_4529,In_2125,In_1990);
nand U4530 (N_4530,In_1073,In_642);
nor U4531 (N_4531,In_1143,In_2616);
nor U4532 (N_4532,In_2585,In_2881);
nand U4533 (N_4533,In_2035,In_1483);
or U4534 (N_4534,In_1912,In_2288);
and U4535 (N_4535,In_2271,In_772);
nor U4536 (N_4536,In_2416,In_713);
xor U4537 (N_4537,In_1516,In_2277);
and U4538 (N_4538,In_95,In_2868);
nor U4539 (N_4539,In_1496,In_1353);
or U4540 (N_4540,In_253,In_2708);
nand U4541 (N_4541,In_187,In_2111);
xor U4542 (N_4542,In_1312,In_1552);
nand U4543 (N_4543,In_2624,In_1552);
and U4544 (N_4544,In_286,In_1282);
nand U4545 (N_4545,In_2596,In_947);
or U4546 (N_4546,In_2015,In_2839);
or U4547 (N_4547,In_1739,In_2684);
nor U4548 (N_4548,In_1395,In_1537);
nor U4549 (N_4549,In_120,In_2045);
nor U4550 (N_4550,In_1136,In_858);
or U4551 (N_4551,In_1629,In_2599);
nand U4552 (N_4552,In_685,In_883);
nor U4553 (N_4553,In_510,In_137);
or U4554 (N_4554,In_2328,In_2660);
nor U4555 (N_4555,In_1575,In_2746);
nor U4556 (N_4556,In_286,In_1803);
nor U4557 (N_4557,In_2087,In_372);
xor U4558 (N_4558,In_1359,In_105);
and U4559 (N_4559,In_384,In_166);
nand U4560 (N_4560,In_840,In_592);
nor U4561 (N_4561,In_2906,In_1162);
or U4562 (N_4562,In_1219,In_483);
or U4563 (N_4563,In_331,In_2004);
or U4564 (N_4564,In_1637,In_1519);
nor U4565 (N_4565,In_1420,In_37);
and U4566 (N_4566,In_1286,In_2135);
or U4567 (N_4567,In_1015,In_2647);
or U4568 (N_4568,In_1377,In_461);
nor U4569 (N_4569,In_102,In_1202);
nor U4570 (N_4570,In_710,In_729);
nand U4571 (N_4571,In_1964,In_1644);
nand U4572 (N_4572,In_2986,In_1317);
xor U4573 (N_4573,In_2580,In_1544);
nor U4574 (N_4574,In_2022,In_1336);
xnor U4575 (N_4575,In_2734,In_2468);
or U4576 (N_4576,In_1665,In_898);
nand U4577 (N_4577,In_536,In_1573);
nor U4578 (N_4578,In_802,In_2440);
or U4579 (N_4579,In_30,In_1709);
or U4580 (N_4580,In_2455,In_903);
or U4581 (N_4581,In_2658,In_2525);
or U4582 (N_4582,In_894,In_2746);
and U4583 (N_4583,In_24,In_1485);
or U4584 (N_4584,In_745,In_569);
nand U4585 (N_4585,In_1539,In_302);
nand U4586 (N_4586,In_160,In_2293);
and U4587 (N_4587,In_1516,In_2484);
or U4588 (N_4588,In_1157,In_2364);
nor U4589 (N_4589,In_284,In_2060);
xor U4590 (N_4590,In_2417,In_1094);
and U4591 (N_4591,In_67,In_2841);
nor U4592 (N_4592,In_2824,In_569);
nand U4593 (N_4593,In_2757,In_727);
xnor U4594 (N_4594,In_365,In_752);
and U4595 (N_4595,In_576,In_864);
nor U4596 (N_4596,In_1918,In_2593);
nor U4597 (N_4597,In_1901,In_1484);
and U4598 (N_4598,In_2344,In_2756);
xnor U4599 (N_4599,In_972,In_2471);
and U4600 (N_4600,In_966,In_1122);
and U4601 (N_4601,In_1450,In_2801);
nand U4602 (N_4602,In_1345,In_2804);
nand U4603 (N_4603,In_1094,In_2545);
nand U4604 (N_4604,In_938,In_1982);
nand U4605 (N_4605,In_467,In_2070);
or U4606 (N_4606,In_138,In_770);
and U4607 (N_4607,In_444,In_1957);
nor U4608 (N_4608,In_1917,In_1309);
or U4609 (N_4609,In_1068,In_21);
nand U4610 (N_4610,In_491,In_1832);
nor U4611 (N_4611,In_1934,In_189);
xor U4612 (N_4612,In_1781,In_1702);
or U4613 (N_4613,In_2475,In_185);
xor U4614 (N_4614,In_1713,In_1515);
or U4615 (N_4615,In_1017,In_950);
or U4616 (N_4616,In_1971,In_1868);
and U4617 (N_4617,In_1904,In_1729);
nor U4618 (N_4618,In_1429,In_745);
or U4619 (N_4619,In_1802,In_2709);
and U4620 (N_4620,In_1844,In_386);
or U4621 (N_4621,In_1404,In_1742);
and U4622 (N_4622,In_2214,In_2225);
and U4623 (N_4623,In_2391,In_279);
nand U4624 (N_4624,In_2171,In_1031);
nand U4625 (N_4625,In_1542,In_1639);
nand U4626 (N_4626,In_1682,In_15);
nand U4627 (N_4627,In_2773,In_2893);
nor U4628 (N_4628,In_388,In_471);
nor U4629 (N_4629,In_1866,In_1687);
xnor U4630 (N_4630,In_1327,In_716);
nand U4631 (N_4631,In_2765,In_2379);
nor U4632 (N_4632,In_1366,In_1127);
nor U4633 (N_4633,In_2197,In_2526);
nor U4634 (N_4634,In_2952,In_1949);
and U4635 (N_4635,In_1987,In_2994);
xor U4636 (N_4636,In_1707,In_1459);
nor U4637 (N_4637,In_1375,In_1371);
and U4638 (N_4638,In_322,In_756);
nand U4639 (N_4639,In_1568,In_1561);
nor U4640 (N_4640,In_1252,In_926);
or U4641 (N_4641,In_878,In_242);
nand U4642 (N_4642,In_1151,In_1487);
nor U4643 (N_4643,In_1255,In_2008);
or U4644 (N_4644,In_2714,In_218);
and U4645 (N_4645,In_2558,In_2);
or U4646 (N_4646,In_1420,In_1663);
nor U4647 (N_4647,In_2755,In_1826);
and U4648 (N_4648,In_2535,In_2554);
and U4649 (N_4649,In_1319,In_891);
nand U4650 (N_4650,In_1571,In_2414);
nand U4651 (N_4651,In_1657,In_515);
nand U4652 (N_4652,In_409,In_2361);
nor U4653 (N_4653,In_296,In_2865);
nor U4654 (N_4654,In_2515,In_1919);
nor U4655 (N_4655,In_1998,In_2166);
nand U4656 (N_4656,In_1241,In_2270);
nor U4657 (N_4657,In_2750,In_584);
xnor U4658 (N_4658,In_2065,In_1090);
or U4659 (N_4659,In_403,In_1200);
nand U4660 (N_4660,In_2489,In_1601);
nor U4661 (N_4661,In_555,In_2141);
nor U4662 (N_4662,In_2084,In_1732);
xor U4663 (N_4663,In_788,In_1349);
nand U4664 (N_4664,In_2733,In_527);
nor U4665 (N_4665,In_1852,In_2787);
nand U4666 (N_4666,In_994,In_1982);
or U4667 (N_4667,In_2485,In_1128);
and U4668 (N_4668,In_1388,In_1009);
nor U4669 (N_4669,In_1130,In_1354);
and U4670 (N_4670,In_1208,In_1476);
and U4671 (N_4671,In_2651,In_2477);
or U4672 (N_4672,In_640,In_1235);
or U4673 (N_4673,In_1062,In_2591);
and U4674 (N_4674,In_1047,In_1186);
nor U4675 (N_4675,In_451,In_758);
nand U4676 (N_4676,In_1642,In_588);
nand U4677 (N_4677,In_2127,In_465);
nand U4678 (N_4678,In_1458,In_2375);
and U4679 (N_4679,In_2509,In_2551);
and U4680 (N_4680,In_2107,In_1297);
nor U4681 (N_4681,In_566,In_1490);
or U4682 (N_4682,In_496,In_1285);
or U4683 (N_4683,In_1867,In_1999);
or U4684 (N_4684,In_1028,In_2704);
nand U4685 (N_4685,In_2616,In_616);
nand U4686 (N_4686,In_915,In_1304);
or U4687 (N_4687,In_2263,In_517);
and U4688 (N_4688,In_1238,In_814);
nand U4689 (N_4689,In_1676,In_1603);
and U4690 (N_4690,In_190,In_1163);
xor U4691 (N_4691,In_1871,In_225);
or U4692 (N_4692,In_1890,In_1064);
nand U4693 (N_4693,In_351,In_2506);
and U4694 (N_4694,In_1709,In_1604);
or U4695 (N_4695,In_2599,In_688);
nand U4696 (N_4696,In_1520,In_2721);
nor U4697 (N_4697,In_1662,In_1700);
nand U4698 (N_4698,In_49,In_2308);
and U4699 (N_4699,In_87,In_151);
nor U4700 (N_4700,In_1418,In_850);
nor U4701 (N_4701,In_1232,In_1076);
xor U4702 (N_4702,In_987,In_381);
nand U4703 (N_4703,In_2492,In_1340);
and U4704 (N_4704,In_530,In_1901);
nand U4705 (N_4705,In_1400,In_1356);
xor U4706 (N_4706,In_499,In_1894);
nand U4707 (N_4707,In_574,In_1037);
or U4708 (N_4708,In_1460,In_763);
or U4709 (N_4709,In_2132,In_963);
and U4710 (N_4710,In_435,In_440);
and U4711 (N_4711,In_1751,In_464);
and U4712 (N_4712,In_1968,In_1284);
xor U4713 (N_4713,In_790,In_2285);
or U4714 (N_4714,In_1114,In_2321);
and U4715 (N_4715,In_249,In_241);
or U4716 (N_4716,In_83,In_444);
or U4717 (N_4717,In_2602,In_2336);
and U4718 (N_4718,In_2673,In_53);
and U4719 (N_4719,In_2807,In_2099);
and U4720 (N_4720,In_2047,In_1089);
or U4721 (N_4721,In_2862,In_2702);
nor U4722 (N_4722,In_785,In_40);
nand U4723 (N_4723,In_1985,In_39);
and U4724 (N_4724,In_2614,In_44);
xnor U4725 (N_4725,In_995,In_2289);
nor U4726 (N_4726,In_704,In_1180);
nand U4727 (N_4727,In_668,In_2375);
nand U4728 (N_4728,In_1222,In_1450);
nand U4729 (N_4729,In_344,In_2123);
and U4730 (N_4730,In_554,In_715);
and U4731 (N_4731,In_1841,In_1699);
or U4732 (N_4732,In_1597,In_793);
nor U4733 (N_4733,In_167,In_815);
and U4734 (N_4734,In_719,In_2356);
nor U4735 (N_4735,In_2399,In_1650);
xor U4736 (N_4736,In_2621,In_1668);
or U4737 (N_4737,In_2062,In_726);
xor U4738 (N_4738,In_1666,In_2058);
xnor U4739 (N_4739,In_1842,In_912);
nor U4740 (N_4740,In_894,In_1722);
nor U4741 (N_4741,In_2653,In_1154);
nor U4742 (N_4742,In_2872,In_2231);
or U4743 (N_4743,In_2121,In_1334);
and U4744 (N_4744,In_1146,In_912);
and U4745 (N_4745,In_1734,In_2192);
nor U4746 (N_4746,In_1148,In_2722);
or U4747 (N_4747,In_2787,In_2092);
or U4748 (N_4748,In_659,In_2794);
nor U4749 (N_4749,In_2285,In_151);
or U4750 (N_4750,In_2172,In_1138);
or U4751 (N_4751,In_2050,In_833);
nand U4752 (N_4752,In_2962,In_2346);
and U4753 (N_4753,In_2310,In_881);
nand U4754 (N_4754,In_2323,In_2501);
and U4755 (N_4755,In_2137,In_2464);
nor U4756 (N_4756,In_493,In_1669);
xor U4757 (N_4757,In_1122,In_66);
xor U4758 (N_4758,In_48,In_1924);
nor U4759 (N_4759,In_1716,In_2503);
or U4760 (N_4760,In_326,In_1004);
nor U4761 (N_4761,In_743,In_1519);
xor U4762 (N_4762,In_1928,In_2650);
or U4763 (N_4763,In_622,In_2611);
nand U4764 (N_4764,In_2384,In_1788);
or U4765 (N_4765,In_1543,In_1882);
and U4766 (N_4766,In_505,In_2142);
nand U4767 (N_4767,In_1746,In_2958);
or U4768 (N_4768,In_354,In_1395);
nand U4769 (N_4769,In_1587,In_2306);
nand U4770 (N_4770,In_1020,In_573);
nor U4771 (N_4771,In_1517,In_2726);
nand U4772 (N_4772,In_827,In_2482);
nor U4773 (N_4773,In_2294,In_1114);
and U4774 (N_4774,In_2021,In_2780);
nand U4775 (N_4775,In_837,In_2413);
and U4776 (N_4776,In_1587,In_2848);
or U4777 (N_4777,In_439,In_1458);
xnor U4778 (N_4778,In_2826,In_2451);
nand U4779 (N_4779,In_996,In_609);
nor U4780 (N_4780,In_2894,In_1800);
nor U4781 (N_4781,In_722,In_755);
nand U4782 (N_4782,In_672,In_2377);
and U4783 (N_4783,In_544,In_790);
nand U4784 (N_4784,In_1885,In_859);
or U4785 (N_4785,In_2718,In_2370);
nand U4786 (N_4786,In_1690,In_195);
or U4787 (N_4787,In_762,In_928);
nor U4788 (N_4788,In_1792,In_2482);
and U4789 (N_4789,In_2515,In_879);
nor U4790 (N_4790,In_275,In_2982);
nand U4791 (N_4791,In_1415,In_718);
nor U4792 (N_4792,In_1161,In_2910);
nor U4793 (N_4793,In_145,In_2008);
or U4794 (N_4794,In_1089,In_471);
and U4795 (N_4795,In_1504,In_530);
nand U4796 (N_4796,In_543,In_404);
and U4797 (N_4797,In_1538,In_809);
or U4798 (N_4798,In_1982,In_2834);
nand U4799 (N_4799,In_262,In_2999);
nand U4800 (N_4800,In_1020,In_1051);
and U4801 (N_4801,In_1611,In_510);
or U4802 (N_4802,In_0,In_2467);
and U4803 (N_4803,In_1685,In_1544);
and U4804 (N_4804,In_2444,In_1398);
xor U4805 (N_4805,In_569,In_2639);
and U4806 (N_4806,In_2002,In_97);
nor U4807 (N_4807,In_1094,In_2889);
nand U4808 (N_4808,In_16,In_2210);
or U4809 (N_4809,In_2930,In_183);
nor U4810 (N_4810,In_1291,In_1325);
nand U4811 (N_4811,In_595,In_2306);
nand U4812 (N_4812,In_2848,In_1369);
nor U4813 (N_4813,In_2345,In_2171);
nor U4814 (N_4814,In_2654,In_1911);
or U4815 (N_4815,In_2569,In_1883);
or U4816 (N_4816,In_1174,In_285);
nor U4817 (N_4817,In_1149,In_615);
nor U4818 (N_4818,In_1194,In_2066);
and U4819 (N_4819,In_2622,In_1191);
nand U4820 (N_4820,In_797,In_2606);
nor U4821 (N_4821,In_2062,In_2335);
nor U4822 (N_4822,In_485,In_1378);
or U4823 (N_4823,In_1556,In_1683);
nand U4824 (N_4824,In_2539,In_391);
nand U4825 (N_4825,In_446,In_2656);
xnor U4826 (N_4826,In_543,In_1586);
nor U4827 (N_4827,In_909,In_1240);
and U4828 (N_4828,In_1939,In_906);
or U4829 (N_4829,In_2293,In_2595);
nor U4830 (N_4830,In_1762,In_1325);
nand U4831 (N_4831,In_1328,In_2079);
xor U4832 (N_4832,In_751,In_979);
xor U4833 (N_4833,In_2225,In_1415);
nand U4834 (N_4834,In_1708,In_2217);
nand U4835 (N_4835,In_1532,In_1602);
nand U4836 (N_4836,In_2944,In_1789);
or U4837 (N_4837,In_1029,In_118);
and U4838 (N_4838,In_2408,In_1003);
nor U4839 (N_4839,In_1285,In_1768);
xor U4840 (N_4840,In_2136,In_608);
xor U4841 (N_4841,In_1811,In_1000);
xor U4842 (N_4842,In_2350,In_2189);
or U4843 (N_4843,In_55,In_1227);
and U4844 (N_4844,In_1599,In_1268);
nand U4845 (N_4845,In_591,In_1890);
or U4846 (N_4846,In_498,In_1530);
nor U4847 (N_4847,In_300,In_1988);
or U4848 (N_4848,In_1917,In_1769);
nor U4849 (N_4849,In_147,In_2161);
or U4850 (N_4850,In_2270,In_1902);
and U4851 (N_4851,In_2000,In_338);
xor U4852 (N_4852,In_765,In_222);
or U4853 (N_4853,In_2530,In_2341);
or U4854 (N_4854,In_1185,In_1950);
and U4855 (N_4855,In_901,In_2061);
or U4856 (N_4856,In_1492,In_1730);
and U4857 (N_4857,In_2649,In_1740);
or U4858 (N_4858,In_892,In_629);
xnor U4859 (N_4859,In_1187,In_1018);
xnor U4860 (N_4860,In_1144,In_2747);
nand U4861 (N_4861,In_444,In_855);
nor U4862 (N_4862,In_1703,In_1431);
and U4863 (N_4863,In_1235,In_2175);
nand U4864 (N_4864,In_1095,In_2871);
and U4865 (N_4865,In_2455,In_2725);
or U4866 (N_4866,In_284,In_139);
and U4867 (N_4867,In_2847,In_1711);
nor U4868 (N_4868,In_2279,In_591);
nand U4869 (N_4869,In_1317,In_337);
and U4870 (N_4870,In_375,In_2792);
or U4871 (N_4871,In_1976,In_897);
nand U4872 (N_4872,In_1555,In_1914);
and U4873 (N_4873,In_1349,In_2587);
nor U4874 (N_4874,In_2132,In_987);
nand U4875 (N_4875,In_1186,In_951);
and U4876 (N_4876,In_1638,In_368);
nor U4877 (N_4877,In_1146,In_462);
and U4878 (N_4878,In_2962,In_1209);
nand U4879 (N_4879,In_762,In_238);
or U4880 (N_4880,In_935,In_1482);
nand U4881 (N_4881,In_1184,In_1956);
and U4882 (N_4882,In_1540,In_37);
or U4883 (N_4883,In_645,In_1626);
and U4884 (N_4884,In_1592,In_1657);
nor U4885 (N_4885,In_152,In_999);
or U4886 (N_4886,In_2045,In_121);
nand U4887 (N_4887,In_1989,In_2716);
or U4888 (N_4888,In_2580,In_680);
nor U4889 (N_4889,In_79,In_26);
or U4890 (N_4890,In_808,In_1924);
nor U4891 (N_4891,In_2785,In_558);
xor U4892 (N_4892,In_1076,In_85);
or U4893 (N_4893,In_1464,In_725);
nor U4894 (N_4894,In_2010,In_2610);
and U4895 (N_4895,In_1626,In_1910);
nor U4896 (N_4896,In_654,In_2281);
and U4897 (N_4897,In_2908,In_2953);
and U4898 (N_4898,In_2330,In_827);
nand U4899 (N_4899,In_2861,In_1775);
or U4900 (N_4900,In_2354,In_1148);
and U4901 (N_4901,In_874,In_777);
and U4902 (N_4902,In_418,In_137);
nand U4903 (N_4903,In_443,In_2119);
nand U4904 (N_4904,In_753,In_1008);
nand U4905 (N_4905,In_2895,In_1050);
nand U4906 (N_4906,In_61,In_2926);
and U4907 (N_4907,In_1471,In_1164);
nand U4908 (N_4908,In_2050,In_1354);
nand U4909 (N_4909,In_929,In_323);
nand U4910 (N_4910,In_2802,In_2158);
or U4911 (N_4911,In_1373,In_1279);
nand U4912 (N_4912,In_2547,In_1592);
nand U4913 (N_4913,In_780,In_497);
or U4914 (N_4914,In_2145,In_1479);
nand U4915 (N_4915,In_2129,In_2572);
nand U4916 (N_4916,In_2142,In_2936);
nand U4917 (N_4917,In_334,In_996);
nand U4918 (N_4918,In_1207,In_927);
or U4919 (N_4919,In_2482,In_1347);
nand U4920 (N_4920,In_1157,In_1188);
nor U4921 (N_4921,In_1877,In_2119);
and U4922 (N_4922,In_2631,In_2435);
nor U4923 (N_4923,In_1240,In_902);
and U4924 (N_4924,In_504,In_648);
xnor U4925 (N_4925,In_2501,In_2170);
or U4926 (N_4926,In_1161,In_258);
or U4927 (N_4927,In_1353,In_559);
and U4928 (N_4928,In_1537,In_1064);
and U4929 (N_4929,In_548,In_1101);
nor U4930 (N_4930,In_2766,In_945);
xnor U4931 (N_4931,In_1604,In_665);
nor U4932 (N_4932,In_1364,In_1746);
or U4933 (N_4933,In_2005,In_955);
nor U4934 (N_4934,In_882,In_2715);
nor U4935 (N_4935,In_1671,In_1784);
xor U4936 (N_4936,In_949,In_1722);
nor U4937 (N_4937,In_747,In_2760);
nand U4938 (N_4938,In_166,In_2614);
nand U4939 (N_4939,In_2837,In_1627);
or U4940 (N_4940,In_2178,In_2764);
nor U4941 (N_4941,In_523,In_2613);
xor U4942 (N_4942,In_2935,In_2214);
and U4943 (N_4943,In_1061,In_2540);
nand U4944 (N_4944,In_1851,In_457);
nand U4945 (N_4945,In_2573,In_787);
nand U4946 (N_4946,In_2111,In_2499);
nand U4947 (N_4947,In_2661,In_1350);
or U4948 (N_4948,In_726,In_1316);
nor U4949 (N_4949,In_903,In_831);
nor U4950 (N_4950,In_773,In_149);
or U4951 (N_4951,In_1759,In_1069);
nand U4952 (N_4952,In_1638,In_2082);
xnor U4953 (N_4953,In_2053,In_2707);
nand U4954 (N_4954,In_591,In_2719);
nor U4955 (N_4955,In_1489,In_2111);
or U4956 (N_4956,In_1243,In_2070);
nor U4957 (N_4957,In_2583,In_1548);
nand U4958 (N_4958,In_1368,In_1940);
xnor U4959 (N_4959,In_928,In_2899);
nor U4960 (N_4960,In_2117,In_2441);
and U4961 (N_4961,In_1713,In_237);
nand U4962 (N_4962,In_1023,In_1690);
nor U4963 (N_4963,In_671,In_2521);
and U4964 (N_4964,In_2804,In_2642);
and U4965 (N_4965,In_343,In_2452);
and U4966 (N_4966,In_1732,In_2101);
or U4967 (N_4967,In_2199,In_995);
xnor U4968 (N_4968,In_2237,In_874);
nor U4969 (N_4969,In_2888,In_31);
nor U4970 (N_4970,In_2183,In_2581);
nand U4971 (N_4971,In_1912,In_1610);
and U4972 (N_4972,In_2551,In_1023);
and U4973 (N_4973,In_1884,In_1489);
nand U4974 (N_4974,In_2557,In_447);
nand U4975 (N_4975,In_2877,In_740);
or U4976 (N_4976,In_507,In_2970);
or U4977 (N_4977,In_2542,In_1933);
nand U4978 (N_4978,In_2888,In_1599);
nor U4979 (N_4979,In_2908,In_1911);
nand U4980 (N_4980,In_2795,In_1934);
nand U4981 (N_4981,In_1845,In_1797);
nor U4982 (N_4982,In_1808,In_2427);
nor U4983 (N_4983,In_786,In_7);
or U4984 (N_4984,In_527,In_1450);
nor U4985 (N_4985,In_98,In_857);
nor U4986 (N_4986,In_450,In_22);
nor U4987 (N_4987,In_2622,In_2493);
or U4988 (N_4988,In_2120,In_2416);
nor U4989 (N_4989,In_686,In_445);
and U4990 (N_4990,In_825,In_2263);
and U4991 (N_4991,In_529,In_2955);
nand U4992 (N_4992,In_890,In_1061);
or U4993 (N_4993,In_747,In_2009);
nand U4994 (N_4994,In_681,In_316);
and U4995 (N_4995,In_171,In_2290);
nor U4996 (N_4996,In_1275,In_1488);
nor U4997 (N_4997,In_412,In_2941);
and U4998 (N_4998,In_1900,In_971);
or U4999 (N_4999,In_2324,In_1918);
xnor U5000 (N_5000,N_3797,N_2889);
nor U5001 (N_5001,N_654,N_2542);
nand U5002 (N_5002,N_3034,N_4325);
xor U5003 (N_5003,N_4260,N_922);
nor U5004 (N_5004,N_2840,N_3958);
nand U5005 (N_5005,N_883,N_2795);
nand U5006 (N_5006,N_3032,N_827);
xnor U5007 (N_5007,N_2733,N_768);
xnor U5008 (N_5008,N_1248,N_4447);
or U5009 (N_5009,N_2377,N_926);
nand U5010 (N_5010,N_4720,N_1417);
and U5011 (N_5011,N_317,N_755);
or U5012 (N_5012,N_2720,N_630);
nor U5013 (N_5013,N_3196,N_2585);
or U5014 (N_5014,N_1434,N_2679);
nand U5015 (N_5015,N_3777,N_3081);
or U5016 (N_5016,N_2212,N_3367);
xor U5017 (N_5017,N_2459,N_2645);
or U5018 (N_5018,N_2895,N_4555);
nand U5019 (N_5019,N_85,N_3174);
and U5020 (N_5020,N_4273,N_4449);
xor U5021 (N_5021,N_2649,N_4588);
and U5022 (N_5022,N_267,N_946);
and U5023 (N_5023,N_324,N_588);
nand U5024 (N_5024,N_2503,N_2379);
xor U5025 (N_5025,N_1017,N_1358);
nor U5026 (N_5026,N_984,N_4545);
and U5027 (N_5027,N_950,N_362);
and U5028 (N_5028,N_2093,N_4840);
nand U5029 (N_5029,N_3271,N_3823);
or U5030 (N_5030,N_2696,N_1567);
nand U5031 (N_5031,N_260,N_374);
or U5032 (N_5032,N_3928,N_2851);
xor U5033 (N_5033,N_742,N_1009);
and U5034 (N_5034,N_2873,N_1829);
or U5035 (N_5035,N_4266,N_3488);
nand U5036 (N_5036,N_3811,N_4208);
nand U5037 (N_5037,N_3495,N_4426);
and U5038 (N_5038,N_1984,N_2406);
nand U5039 (N_5039,N_3046,N_3068);
and U5040 (N_5040,N_2258,N_461);
and U5041 (N_5041,N_4275,N_1587);
nand U5042 (N_5042,N_3275,N_746);
nand U5043 (N_5043,N_3048,N_162);
nand U5044 (N_5044,N_2178,N_2639);
or U5045 (N_5045,N_1909,N_3339);
and U5046 (N_5046,N_1910,N_3840);
and U5047 (N_5047,N_2755,N_2552);
and U5048 (N_5048,N_918,N_2063);
or U5049 (N_5049,N_998,N_686);
and U5050 (N_5050,N_210,N_3424);
or U5051 (N_5051,N_1806,N_1274);
nor U5052 (N_5052,N_2702,N_4929);
nor U5053 (N_5053,N_3294,N_614);
and U5054 (N_5054,N_2670,N_4042);
nand U5055 (N_5055,N_3085,N_3964);
or U5056 (N_5056,N_3129,N_1459);
nor U5057 (N_5057,N_1246,N_5);
nor U5058 (N_5058,N_3882,N_3996);
and U5059 (N_5059,N_1818,N_3901);
and U5060 (N_5060,N_4284,N_452);
and U5061 (N_5061,N_3915,N_3494);
nor U5062 (N_5062,N_3920,N_1714);
or U5063 (N_5063,N_3062,N_3031);
or U5064 (N_5064,N_4335,N_1219);
nand U5065 (N_5065,N_497,N_1528);
nor U5066 (N_5066,N_2899,N_3900);
nor U5067 (N_5067,N_189,N_877);
or U5068 (N_5068,N_4951,N_4727);
nor U5069 (N_5069,N_951,N_985);
and U5070 (N_5070,N_3107,N_1223);
xor U5071 (N_5071,N_2605,N_257);
nand U5072 (N_5072,N_3155,N_2399);
nor U5073 (N_5073,N_3423,N_3320);
nor U5074 (N_5074,N_4666,N_1476);
and U5075 (N_5075,N_2501,N_4881);
or U5076 (N_5076,N_2532,N_3388);
nand U5077 (N_5077,N_4893,N_1841);
and U5078 (N_5078,N_4764,N_545);
or U5079 (N_5079,N_4674,N_3186);
or U5080 (N_5080,N_2419,N_4114);
or U5081 (N_5081,N_3855,N_2353);
nor U5082 (N_5082,N_3661,N_2727);
and U5083 (N_5083,N_1923,N_3607);
nand U5084 (N_5084,N_2615,N_541);
nor U5085 (N_5085,N_2666,N_1642);
nor U5086 (N_5086,N_4097,N_2913);
and U5087 (N_5087,N_4504,N_529);
and U5088 (N_5088,N_2978,N_2031);
nand U5089 (N_5089,N_2216,N_4531);
nor U5090 (N_5090,N_4312,N_1065);
and U5091 (N_5091,N_4597,N_3864);
and U5092 (N_5092,N_1804,N_695);
or U5093 (N_5093,N_592,N_2085);
or U5094 (N_5094,N_2121,N_1141);
nand U5095 (N_5095,N_1641,N_4548);
nand U5096 (N_5096,N_4746,N_516);
nand U5097 (N_5097,N_3534,N_2732);
and U5098 (N_5098,N_3714,N_2543);
or U5099 (N_5099,N_4985,N_2464);
and U5100 (N_5100,N_1530,N_4927);
and U5101 (N_5101,N_1364,N_2315);
and U5102 (N_5102,N_3878,N_35);
or U5103 (N_5103,N_2064,N_1666);
or U5104 (N_5104,N_2157,N_3002);
xnor U5105 (N_5105,N_4904,N_2407);
nor U5106 (N_5106,N_3839,N_2265);
and U5107 (N_5107,N_1594,N_3649);
or U5108 (N_5108,N_4387,N_3590);
nand U5109 (N_5109,N_2502,N_3166);
nand U5110 (N_5110,N_797,N_2741);
nor U5111 (N_5111,N_3470,N_3153);
or U5112 (N_5112,N_3486,N_942);
nor U5113 (N_5113,N_3184,N_1902);
or U5114 (N_5114,N_2324,N_1016);
nand U5115 (N_5115,N_3563,N_2841);
nor U5116 (N_5116,N_2907,N_4236);
nand U5117 (N_5117,N_4759,N_597);
nand U5118 (N_5118,N_2188,N_2109);
nor U5119 (N_5119,N_2317,N_2508);
xnor U5120 (N_5120,N_4380,N_416);
and U5121 (N_5121,N_4579,N_2438);
or U5122 (N_5122,N_1264,N_782);
or U5123 (N_5123,N_2183,N_1133);
and U5124 (N_5124,N_2677,N_4346);
and U5125 (N_5125,N_668,N_730);
and U5126 (N_5126,N_2263,N_641);
xnor U5127 (N_5127,N_816,N_1028);
or U5128 (N_5128,N_2339,N_1496);
nand U5129 (N_5129,N_2675,N_3451);
or U5130 (N_5130,N_3899,N_850);
and U5131 (N_5131,N_2245,N_2614);
nor U5132 (N_5132,N_1455,N_4090);
or U5133 (N_5133,N_3983,N_4280);
and U5134 (N_5134,N_2864,N_186);
nand U5135 (N_5135,N_206,N_3306);
nor U5136 (N_5136,N_4762,N_4327);
and U5137 (N_5137,N_4175,N_4660);
xnor U5138 (N_5138,N_975,N_3981);
xnor U5139 (N_5139,N_1071,N_43);
nor U5140 (N_5140,N_2955,N_1793);
and U5141 (N_5141,N_2777,N_4183);
or U5142 (N_5142,N_3654,N_1132);
and U5143 (N_5143,N_2549,N_4702);
xor U5144 (N_5144,N_143,N_4887);
nand U5145 (N_5145,N_2954,N_1032);
or U5146 (N_5146,N_4077,N_4729);
and U5147 (N_5147,N_1200,N_4288);
and U5148 (N_5148,N_460,N_3553);
or U5149 (N_5149,N_1457,N_1033);
nand U5150 (N_5150,N_4373,N_3157);
nor U5151 (N_5151,N_943,N_4664);
or U5152 (N_5152,N_860,N_2500);
or U5153 (N_5153,N_1247,N_1772);
nor U5154 (N_5154,N_3243,N_4388);
nor U5155 (N_5155,N_925,N_4832);
or U5156 (N_5156,N_1099,N_3954);
nor U5157 (N_5157,N_667,N_145);
nor U5158 (N_5158,N_4937,N_747);
or U5159 (N_5159,N_4263,N_3735);
nor U5160 (N_5160,N_219,N_4414);
and U5161 (N_5161,N_4146,N_2189);
and U5162 (N_5162,N_3611,N_2718);
nand U5163 (N_5163,N_2968,N_4307);
nor U5164 (N_5164,N_770,N_2694);
nor U5165 (N_5165,N_2253,N_4405);
or U5166 (N_5166,N_1925,N_3439);
and U5167 (N_5167,N_1573,N_4713);
and U5168 (N_5168,N_4022,N_3403);
nand U5169 (N_5169,N_1849,N_3598);
or U5170 (N_5170,N_4876,N_3577);
nand U5171 (N_5171,N_2411,N_3741);
nand U5172 (N_5172,N_4210,N_2294);
nand U5173 (N_5173,N_3302,N_930);
nand U5174 (N_5174,N_3137,N_181);
or U5175 (N_5175,N_4132,N_4317);
and U5176 (N_5176,N_2660,N_2710);
nand U5177 (N_5177,N_2689,N_203);
and U5178 (N_5178,N_3509,N_1342);
nor U5179 (N_5179,N_3724,N_1609);
nand U5180 (N_5180,N_2081,N_2652);
nand U5181 (N_5181,N_655,N_1324);
xnor U5182 (N_5182,N_1504,N_620);
and U5183 (N_5183,N_272,N_454);
nand U5184 (N_5184,N_37,N_2477);
xor U5185 (N_5185,N_2115,N_2402);
nor U5186 (N_5186,N_3987,N_4193);
nor U5187 (N_5187,N_2517,N_3799);
nand U5188 (N_5188,N_4877,N_3982);
nand U5189 (N_5189,N_2867,N_617);
or U5190 (N_5190,N_1025,N_3018);
and U5191 (N_5191,N_999,N_3537);
and U5192 (N_5192,N_4639,N_2229);
and U5193 (N_5193,N_3217,N_4155);
nor U5194 (N_5194,N_2586,N_2240);
nor U5195 (N_5195,N_3482,N_785);
nand U5196 (N_5196,N_1490,N_3730);
nand U5197 (N_5197,N_1908,N_2105);
xor U5198 (N_5198,N_3356,N_1869);
nor U5199 (N_5199,N_2273,N_550);
nor U5200 (N_5200,N_508,N_1506);
and U5201 (N_5201,N_1037,N_3206);
or U5202 (N_5202,N_3664,N_3195);
and U5203 (N_5203,N_2318,N_3407);
nand U5204 (N_5204,N_2142,N_448);
nor U5205 (N_5205,N_3487,N_1877);
nor U5206 (N_5206,N_2557,N_1309);
nand U5207 (N_5207,N_237,N_4040);
xor U5208 (N_5208,N_4247,N_3736);
or U5209 (N_5209,N_3962,N_3);
and U5210 (N_5210,N_428,N_3063);
nor U5211 (N_5211,N_4835,N_3581);
or U5212 (N_5212,N_456,N_1307);
or U5213 (N_5213,N_2998,N_3700);
xor U5214 (N_5214,N_1393,N_1172);
or U5215 (N_5215,N_1083,N_3222);
nor U5216 (N_5216,N_4763,N_2098);
nand U5217 (N_5217,N_3550,N_2092);
and U5218 (N_5218,N_4956,N_3197);
nor U5219 (N_5219,N_1548,N_1366);
and U5220 (N_5220,N_1701,N_706);
and U5221 (N_5221,N_4464,N_3112);
nand U5222 (N_5222,N_2228,N_3746);
xnor U5223 (N_5223,N_3385,N_1078);
or U5224 (N_5224,N_749,N_1308);
nand U5225 (N_5225,N_766,N_316);
and U5226 (N_5226,N_4196,N_632);
and U5227 (N_5227,N_4493,N_295);
nand U5228 (N_5228,N_3304,N_1379);
and U5229 (N_5229,N_1492,N_119);
nand U5230 (N_5230,N_1605,N_2144);
and U5231 (N_5231,N_3476,N_2219);
nor U5232 (N_5232,N_3378,N_4445);
and U5233 (N_5233,N_4103,N_18);
nor U5234 (N_5234,N_1543,N_1040);
and U5235 (N_5235,N_2089,N_2492);
and U5236 (N_5236,N_1993,N_4502);
and U5237 (N_5237,N_4629,N_4988);
nor U5238 (N_5238,N_4778,N_3663);
nand U5239 (N_5239,N_801,N_4558);
and U5240 (N_5240,N_2844,N_1374);
xor U5241 (N_5241,N_2535,N_3414);
or U5242 (N_5242,N_4153,N_1508);
and U5243 (N_5243,N_4882,N_2281);
nand U5244 (N_5244,N_1166,N_2007);
or U5245 (N_5245,N_4890,N_1552);
and U5246 (N_5246,N_1255,N_1621);
and U5247 (N_5247,N_4051,N_2238);
nand U5248 (N_5248,N_1004,N_2724);
and U5249 (N_5249,N_1768,N_3462);
and U5250 (N_5250,N_1432,N_3859);
nand U5251 (N_5251,N_4495,N_2322);
nor U5252 (N_5252,N_2202,N_1420);
nor U5253 (N_5253,N_2361,N_4747);
nor U5254 (N_5254,N_1940,N_2388);
and U5255 (N_5255,N_4136,N_1137);
and U5256 (N_5256,N_4370,N_4158);
nand U5257 (N_5257,N_4848,N_1510);
xnor U5258 (N_5258,N_3390,N_700);
and U5259 (N_5259,N_3043,N_3483);
nor U5260 (N_5260,N_1310,N_1178);
nor U5261 (N_5261,N_4024,N_1222);
xnor U5262 (N_5262,N_2824,N_4374);
or U5263 (N_5263,N_2765,N_862);
nor U5264 (N_5264,N_2529,N_1936);
or U5265 (N_5265,N_697,N_4698);
and U5266 (N_5266,N_638,N_335);
nand U5267 (N_5267,N_1332,N_2173);
nor U5268 (N_5268,N_78,N_1328);
or U5269 (N_5269,N_376,N_3150);
nor U5270 (N_5270,N_822,N_4138);
nand U5271 (N_5271,N_4498,N_222);
or U5272 (N_5272,N_2846,N_512);
and U5273 (N_5273,N_1898,N_4168);
and U5274 (N_5274,N_2625,N_2078);
and U5275 (N_5275,N_1146,N_4487);
nor U5276 (N_5276,N_4688,N_3169);
nor U5277 (N_5277,N_745,N_2553);
nor U5278 (N_5278,N_3175,N_202);
or U5279 (N_5279,N_2896,N_3616);
nor U5280 (N_5280,N_1553,N_1035);
nand U5281 (N_5281,N_927,N_4396);
or U5282 (N_5282,N_1343,N_2480);
nor U5283 (N_5283,N_634,N_750);
nand U5284 (N_5284,N_304,N_4306);
and U5285 (N_5285,N_666,N_205);
and U5286 (N_5286,N_1148,N_2497);
nand U5287 (N_5287,N_2974,N_1655);
and U5288 (N_5288,N_3065,N_3203);
and U5289 (N_5289,N_2785,N_3202);
and U5290 (N_5290,N_197,N_3528);
nor U5291 (N_5291,N_4482,N_4126);
and U5292 (N_5292,N_2369,N_1746);
nor U5293 (N_5293,N_2367,N_4105);
xor U5294 (N_5294,N_1495,N_4272);
nor U5295 (N_5295,N_1081,N_2374);
nor U5296 (N_5296,N_2192,N_3473);
nor U5297 (N_5297,N_4406,N_2383);
nand U5298 (N_5298,N_1335,N_4412);
xor U5299 (N_5299,N_3051,N_772);
and U5300 (N_5300,N_212,N_2310);
nand U5301 (N_5301,N_3884,N_3541);
and U5302 (N_5302,N_4584,N_4140);
and U5303 (N_5303,N_3352,N_1363);
or U5304 (N_5304,N_4943,N_1987);
or U5305 (N_5305,N_4323,N_4625);
nand U5306 (N_5306,N_2776,N_3665);
xnor U5307 (N_5307,N_2137,N_277);
and U5308 (N_5308,N_1302,N_4806);
nand U5309 (N_5309,N_4753,N_3709);
or U5310 (N_5310,N_4532,N_378);
nor U5311 (N_5311,N_4811,N_1879);
or U5312 (N_5312,N_4656,N_1722);
nand U5313 (N_5313,N_841,N_4041);
nor U5314 (N_5314,N_221,N_216);
and U5315 (N_5315,N_1547,N_546);
and U5316 (N_5316,N_180,N_2862);
nand U5317 (N_5317,N_294,N_217);
and U5318 (N_5318,N_1619,N_1242);
and U5319 (N_5319,N_3837,N_3231);
nand U5320 (N_5320,N_3959,N_1845);
xnor U5321 (N_5321,N_4712,N_902);
and U5322 (N_5322,N_1852,N_1618);
or U5323 (N_5323,N_1723,N_4993);
nand U5324 (N_5324,N_532,N_2457);
and U5325 (N_5325,N_3160,N_3705);
and U5326 (N_5326,N_3848,N_3397);
and U5327 (N_5327,N_2226,N_282);
or U5328 (N_5328,N_330,N_981);
nand U5329 (N_5329,N_4045,N_1600);
and U5330 (N_5330,N_2218,N_3193);
nor U5331 (N_5331,N_3118,N_3931);
nor U5332 (N_5332,N_4220,N_4783);
nand U5333 (N_5333,N_3697,N_4711);
nand U5334 (N_5334,N_891,N_4311);
and U5335 (N_5335,N_776,N_3545);
nand U5336 (N_5336,N_2661,N_325);
and U5337 (N_5337,N_2537,N_1256);
nand U5338 (N_5338,N_2260,N_3718);
and U5339 (N_5339,N_3047,N_825);
and U5340 (N_5340,N_184,N_4462);
nand U5341 (N_5341,N_1238,N_4612);
nand U5342 (N_5342,N_4213,N_4089);
nand U5343 (N_5343,N_236,N_3381);
nand U5344 (N_5344,N_1176,N_3694);
nand U5345 (N_5345,N_1582,N_284);
nand U5346 (N_5346,N_1224,N_3543);
nor U5347 (N_5347,N_230,N_4431);
nor U5348 (N_5348,N_3961,N_601);
nand U5349 (N_5349,N_3805,N_658);
xnor U5350 (N_5350,N_1931,N_3090);
nand U5351 (N_5351,N_2789,N_814);
and U5352 (N_5352,N_3591,N_1912);
or U5353 (N_5353,N_4790,N_1045);
nand U5354 (N_5354,N_3621,N_983);
and U5355 (N_5355,N_4807,N_227);
or U5356 (N_5356,N_1177,N_3605);
nor U5357 (N_5357,N_4507,N_959);
nor U5358 (N_5358,N_4074,N_2580);
and U5359 (N_5359,N_3000,N_3919);
and U5360 (N_5360,N_3387,N_4366);
nand U5361 (N_5361,N_1418,N_684);
nand U5362 (N_5362,N_1481,N_1182);
and U5363 (N_5363,N_4433,N_1314);
and U5364 (N_5364,N_4537,N_3923);
or U5365 (N_5365,N_1846,N_4015);
nor U5366 (N_5366,N_266,N_3921);
nor U5367 (N_5367,N_2003,N_331);
nor U5368 (N_5368,N_1697,N_4219);
nand U5369 (N_5369,N_4745,N_3104);
or U5370 (N_5370,N_2717,N_4377);
and U5371 (N_5371,N_1225,N_1779);
nor U5372 (N_5372,N_2009,N_1950);
nand U5373 (N_5373,N_2279,N_151);
nand U5374 (N_5374,N_1327,N_661);
or U5375 (N_5375,N_394,N_2651);
and U5376 (N_5376,N_3588,N_63);
nor U5377 (N_5377,N_1419,N_4722);
nor U5378 (N_5378,N_900,N_1960);
or U5379 (N_5379,N_4635,N_681);
or U5380 (N_5380,N_3761,N_979);
and U5381 (N_5381,N_2721,N_2931);
and U5382 (N_5382,N_4064,N_2210);
xor U5383 (N_5383,N_4486,N_2575);
nor U5384 (N_5384,N_3846,N_4160);
xor U5385 (N_5385,N_3087,N_2693);
or U5386 (N_5386,N_1676,N_4996);
or U5387 (N_5387,N_3830,N_4009);
nand U5388 (N_5388,N_4048,N_1799);
nand U5389 (N_5389,N_4873,N_4922);
nand U5390 (N_5390,N_2608,N_4365);
nand U5391 (N_5391,N_74,N_3073);
and U5392 (N_5392,N_849,N_1730);
and U5393 (N_5393,N_2635,N_2187);
and U5394 (N_5394,N_6,N_520);
xnor U5395 (N_5395,N_4233,N_3986);
nand U5396 (N_5396,N_949,N_4888);
nand U5397 (N_5397,N_1380,N_1997);
xor U5398 (N_5398,N_1991,N_3484);
nand U5399 (N_5399,N_3747,N_561);
xnor U5400 (N_5400,N_2338,N_1020);
and U5401 (N_5401,N_4821,N_4734);
or U5402 (N_5402,N_253,N_4100);
nand U5403 (N_5403,N_990,N_3334);
nor U5404 (N_5404,N_2044,N_2619);
and U5405 (N_5405,N_4201,N_13);
and U5406 (N_5406,N_829,N_1947);
xor U5407 (N_5407,N_723,N_2072);
nor U5408 (N_5408,N_2012,N_4669);
and U5409 (N_5409,N_558,N_726);
and U5410 (N_5410,N_4239,N_2282);
and U5411 (N_5411,N_3906,N_1161);
xnor U5412 (N_5412,N_4680,N_3755);
nand U5413 (N_5413,N_4419,N_157);
or U5414 (N_5414,N_3831,N_4889);
xnor U5415 (N_5415,N_3491,N_573);
nand U5416 (N_5416,N_2803,N_4653);
and U5417 (N_5417,N_1979,N_312);
or U5418 (N_5418,N_2792,N_232);
nand U5419 (N_5419,N_2359,N_646);
nor U5420 (N_5420,N_223,N_4065);
and U5421 (N_5421,N_3270,N_1531);
or U5422 (N_5422,N_2432,N_4257);
nand U5423 (N_5423,N_446,N_2819);
nor U5424 (N_5424,N_842,N_773);
nand U5425 (N_5425,N_36,N_1544);
or U5426 (N_5426,N_388,N_142);
nor U5427 (N_5427,N_4497,N_2321);
or U5428 (N_5428,N_3932,N_4321);
nand U5429 (N_5429,N_1890,N_2050);
and U5430 (N_5430,N_3519,N_3187);
nand U5431 (N_5431,N_2516,N_2155);
and U5432 (N_5432,N_1,N_4586);
nor U5433 (N_5433,N_3521,N_451);
nor U5434 (N_5434,N_3583,N_3331);
nor U5435 (N_5435,N_2865,N_117);
nor U5436 (N_5436,N_1549,N_3907);
nand U5437 (N_5437,N_3386,N_2977);
nor U5438 (N_5438,N_2588,N_1319);
nand U5439 (N_5439,N_3013,N_3529);
xnor U5440 (N_5440,N_4006,N_1217);
nand U5441 (N_5441,N_1817,N_4809);
or U5442 (N_5442,N_4204,N_4242);
or U5443 (N_5443,N_759,N_420);
and U5444 (N_5444,N_4071,N_738);
or U5445 (N_5445,N_2022,N_3402);
nor U5446 (N_5446,N_194,N_4084);
xnor U5447 (N_5447,N_4453,N_4187);
or U5448 (N_5448,N_720,N_761);
xor U5449 (N_5449,N_3659,N_50);
nor U5450 (N_5450,N_1199,N_4027);
xor U5451 (N_5451,N_1140,N_4375);
and U5452 (N_5452,N_4983,N_4390);
xor U5453 (N_5453,N_3345,N_3952);
or U5454 (N_5454,N_2932,N_1372);
and U5455 (N_5455,N_540,N_2804);
nor U5456 (N_5456,N_910,N_3007);
nand U5457 (N_5457,N_4329,N_141);
nand U5458 (N_5458,N_3219,N_2331);
xnor U5459 (N_5459,N_4144,N_3096);
and U5460 (N_5460,N_1976,N_3891);
or U5461 (N_5461,N_3168,N_1637);
xnor U5462 (N_5462,N_2740,N_2002);
nor U5463 (N_5463,N_762,N_1063);
or U5464 (N_5464,N_3673,N_2962);
nand U5465 (N_5465,N_441,N_226);
nand U5466 (N_5466,N_3852,N_255);
nand U5467 (N_5467,N_2515,N_4189);
and U5468 (N_5468,N_3875,N_1982);
nand U5469 (N_5469,N_1597,N_719);
xor U5470 (N_5470,N_4202,N_3369);
nor U5471 (N_5471,N_3795,N_4017);
and U5472 (N_5472,N_1783,N_1102);
nor U5473 (N_5473,N_938,N_359);
or U5474 (N_5474,N_3950,N_1764);
nor U5475 (N_5475,N_4954,N_4611);
or U5476 (N_5476,N_4276,N_2570);
and U5477 (N_5477,N_3426,N_2133);
nand U5478 (N_5478,N_3238,N_894);
nor U5479 (N_5479,N_4650,N_4206);
xor U5480 (N_5480,N_3310,N_3430);
and U5481 (N_5481,N_2082,N_2108);
xnor U5482 (N_5482,N_758,N_1651);
and U5483 (N_5483,N_3936,N_3978);
or U5484 (N_5484,N_4372,N_2903);
nor U5485 (N_5485,N_4787,N_4351);
and U5486 (N_5486,N_246,N_3708);
nand U5487 (N_5487,N_1671,N_3834);
and U5488 (N_5488,N_4032,N_563);
and U5489 (N_5489,N_3028,N_3968);
nor U5490 (N_5490,N_935,N_4358);
and U5491 (N_5491,N_3643,N_4198);
nand U5492 (N_5492,N_1175,N_1123);
or U5493 (N_5493,N_1911,N_1679);
nor U5494 (N_5494,N_1320,N_4770);
nand U5495 (N_5495,N_1945,N_1860);
nand U5496 (N_5496,N_3867,N_1079);
or U5497 (N_5497,N_3030,N_1514);
nand U5498 (N_5498,N_3699,N_298);
or U5499 (N_5499,N_4647,N_3566);
nand U5500 (N_5500,N_305,N_3512);
nor U5501 (N_5501,N_1124,N_4569);
nand U5502 (N_5502,N_4483,N_4613);
and U5503 (N_5503,N_4805,N_2988);
or U5504 (N_5504,N_3468,N_1561);
or U5505 (N_5505,N_3399,N_1026);
xor U5506 (N_5506,N_4489,N_2019);
nor U5507 (N_5507,N_3069,N_3567);
or U5508 (N_5508,N_2332,N_1499);
nor U5509 (N_5509,N_1832,N_1630);
and U5510 (N_5510,N_2150,N_1542);
nand U5511 (N_5511,N_3518,N_1788);
nor U5512 (N_5512,N_2211,N_796);
nand U5513 (N_5513,N_948,N_969);
xor U5514 (N_5514,N_496,N_2598);
xnor U5515 (N_5515,N_3911,N_249);
nand U5516 (N_5516,N_1271,N_4853);
nand U5517 (N_5517,N_3721,N_1244);
nand U5518 (N_5518,N_149,N_537);
nand U5519 (N_5519,N_3719,N_2644);
nor U5520 (N_5520,N_4268,N_478);
nor U5521 (N_5521,N_321,N_4820);
nand U5522 (N_5522,N_731,N_1387);
and U5523 (N_5523,N_1464,N_3435);
and U5524 (N_5524,N_100,N_4353);
and U5525 (N_5525,N_21,N_4892);
nand U5526 (N_5526,N_2312,N_1725);
or U5527 (N_5527,N_865,N_1656);
nor U5528 (N_5528,N_3319,N_2395);
nor U5529 (N_5529,N_4651,N_483);
nor U5530 (N_5530,N_108,N_377);
or U5531 (N_5531,N_4417,N_4057);
nand U5532 (N_5532,N_3560,N_4076);
or U5533 (N_5533,N_3237,N_4630);
and U5534 (N_5534,N_3948,N_1185);
nor U5535 (N_5535,N_2746,N_4383);
nor U5536 (N_5536,N_1661,N_673);
nand U5537 (N_5537,N_1294,N_3743);
nand U5538 (N_5538,N_433,N_4691);
or U5539 (N_5539,N_4053,N_553);
nand U5540 (N_5540,N_2214,N_778);
xnor U5541 (N_5541,N_4440,N_309);
or U5542 (N_5542,N_1710,N_4468);
nand U5543 (N_5543,N_2191,N_3038);
and U5544 (N_5544,N_3114,N_4511);
nor U5545 (N_5545,N_413,N_3888);
xor U5546 (N_5546,N_3542,N_1477);
or U5547 (N_5547,N_2306,N_1915);
nor U5548 (N_5548,N_1355,N_2878);
nor U5549 (N_5549,N_1472,N_2827);
and U5550 (N_5550,N_4178,N_715);
and U5551 (N_5551,N_4207,N_2094);
and U5552 (N_5552,N_2859,N_1626);
nor U5553 (N_5553,N_32,N_1488);
nand U5554 (N_5554,N_707,N_2832);
nand U5555 (N_5555,N_3636,N_3841);
or U5556 (N_5556,N_2354,N_468);
or U5557 (N_5557,N_3335,N_4092);
nor U5558 (N_5558,N_4928,N_919);
nor U5559 (N_5559,N_1765,N_3625);
and U5560 (N_5560,N_2623,N_3922);
and U5561 (N_5561,N_4768,N_600);
or U5562 (N_5562,N_873,N_3210);
nand U5563 (N_5563,N_310,N_466);
nor U5564 (N_5564,N_1522,N_2633);
and U5565 (N_5565,N_2224,N_1330);
and U5566 (N_5566,N_4452,N_358);
and U5567 (N_5567,N_4392,N_4895);
or U5568 (N_5568,N_2530,N_815);
nand U5569 (N_5569,N_3433,N_286);
and U5570 (N_5570,N_4561,N_1165);
nor U5571 (N_5571,N_2242,N_4850);
nor U5572 (N_5572,N_4244,N_3253);
nand U5573 (N_5573,N_4641,N_3740);
and U5574 (N_5574,N_1763,N_907);
nor U5575 (N_5575,N_830,N_1965);
nor U5576 (N_5576,N_275,N_3493);
nand U5577 (N_5577,N_1889,N_714);
nand U5578 (N_5578,N_1670,N_1321);
nor U5579 (N_5579,N_4499,N_4860);
or U5580 (N_5580,N_4553,N_4423);
or U5581 (N_5581,N_2786,N_2106);
or U5582 (N_5582,N_1828,N_4190);
or U5583 (N_5583,N_1050,N_3300);
and U5584 (N_5584,N_3977,N_3620);
or U5585 (N_5585,N_2509,N_127);
nand U5586 (N_5586,N_261,N_2385);
nand U5587 (N_5587,N_920,N_931);
nor U5588 (N_5588,N_3301,N_1389);
nor U5589 (N_5589,N_193,N_1311);
nand U5590 (N_5590,N_251,N_1385);
nand U5591 (N_5591,N_439,N_4829);
or U5592 (N_5592,N_2771,N_1589);
xor U5593 (N_5593,N_610,N_1534);
nand U5594 (N_5594,N_3255,N_4450);
nor U5595 (N_5595,N_4792,N_4229);
nor U5596 (N_5596,N_2449,N_4725);
or U5597 (N_5597,N_2482,N_1090);
nand U5598 (N_5598,N_4991,N_4580);
nand U5599 (N_5599,N_4294,N_4872);
nand U5600 (N_5600,N_2636,N_3535);
or U5601 (N_5601,N_3316,N_436);
or U5602 (N_5602,N_4348,N_1570);
or U5603 (N_5603,N_1583,N_380);
xnor U5604 (N_5604,N_4708,N_4339);
and U5605 (N_5605,N_2234,N_4384);
xnor U5606 (N_5606,N_3815,N_552);
and U5607 (N_5607,N_2384,N_4142);
xor U5608 (N_5608,N_4769,N_3147);
nand U5609 (N_5609,N_28,N_2448);
nor U5610 (N_5610,N_415,N_4836);
and U5611 (N_5611,N_3053,N_4139);
and U5612 (N_5612,N_2117,N_1273);
nor U5613 (N_5613,N_3416,N_3817);
or U5614 (N_5614,N_3707,N_1628);
and U5615 (N_5615,N_1507,N_1635);
or U5616 (N_5616,N_4283,N_4551);
and U5617 (N_5617,N_1526,N_2695);
or U5618 (N_5618,N_2734,N_2944);
and U5619 (N_5619,N_2316,N_2275);
nor U5620 (N_5620,N_647,N_1649);
nor U5621 (N_5621,N_2952,N_4199);
nor U5622 (N_5622,N_914,N_3292);
or U5623 (N_5623,N_4672,N_2861);
xnor U5624 (N_5624,N_3376,N_3312);
nor U5625 (N_5625,N_2830,N_4723);
nand U5626 (N_5626,N_105,N_2601);
and U5627 (N_5627,N_3240,N_31);
nand U5628 (N_5628,N_4901,N_3248);
nand U5629 (N_5629,N_54,N_1100);
nor U5630 (N_5630,N_4049,N_4604);
and U5631 (N_5631,N_2166,N_3821);
or U5632 (N_5632,N_1952,N_2882);
or U5633 (N_5633,N_1266,N_4174);
and U5634 (N_5634,N_3380,N_435);
and U5635 (N_5635,N_1116,N_3772);
nor U5636 (N_5636,N_2203,N_2730);
and U5637 (N_5637,N_2141,N_3009);
or U5638 (N_5638,N_3516,N_3615);
and U5639 (N_5639,N_4170,N_4638);
and U5640 (N_5640,N_1059,N_3973);
or U5641 (N_5641,N_1031,N_821);
nor U5642 (N_5642,N_3568,N_2838);
or U5643 (N_5643,N_1824,N_1443);
and U5644 (N_5644,N_4589,N_125);
and U5645 (N_5645,N_3097,N_1648);
and U5646 (N_5646,N_2688,N_527);
and U5647 (N_5647,N_2505,N_419);
or U5648 (N_5648,N_2493,N_4813);
nor U5649 (N_5649,N_1155,N_4616);
nor U5650 (N_5650,N_328,N_405);
nor U5651 (N_5651,N_4252,N_2393);
nor U5652 (N_5652,N_1608,N_1181);
or U5653 (N_5653,N_2966,N_3067);
xnor U5654 (N_5654,N_370,N_2650);
and U5655 (N_5655,N_4133,N_4743);
or U5656 (N_5656,N_1770,N_4182);
and U5657 (N_5657,N_905,N_1288);
nand U5658 (N_5658,N_1475,N_175);
or U5659 (N_5659,N_4432,N_3448);
nor U5660 (N_5660,N_2563,N_72);
nand U5661 (N_5661,N_4303,N_642);
nand U5662 (N_5662,N_280,N_4437);
nor U5663 (N_5663,N_3666,N_3070);
or U5664 (N_5664,N_640,N_3832);
and U5665 (N_5665,N_4262,N_3162);
nor U5666 (N_5666,N_4345,N_4844);
xnor U5667 (N_5667,N_4330,N_1080);
or U5668 (N_5668,N_4917,N_3720);
nor U5669 (N_5669,N_4606,N_2398);
nor U5670 (N_5670,N_1740,N_1985);
or U5671 (N_5671,N_297,N_4167);
or U5672 (N_5672,N_3422,N_2034);
nand U5673 (N_5673,N_3517,N_1489);
nand U5674 (N_5674,N_3116,N_4458);
or U5675 (N_5675,N_2074,N_2016);
nor U5676 (N_5676,N_1511,N_1186);
nand U5677 (N_5677,N_2000,N_2524);
nand U5678 (N_5678,N_2848,N_3612);
or U5679 (N_5679,N_1298,N_2934);
and U5680 (N_5680,N_2458,N_4484);
xnor U5681 (N_5681,N_4070,N_1093);
nor U5682 (N_5682,N_2368,N_2251);
and U5683 (N_5683,N_677,N_1907);
and U5684 (N_5684,N_565,N_687);
nand U5685 (N_5685,N_909,N_3533);
nor U5686 (N_5686,N_1955,N_2521);
or U5687 (N_5687,N_3600,N_107);
and U5688 (N_5688,N_4563,N_870);
xnor U5689 (N_5689,N_1706,N_2087);
and U5690 (N_5690,N_4851,N_341);
or U5691 (N_5691,N_3119,N_3679);
nor U5692 (N_5692,N_1195,N_4395);
nor U5693 (N_5693,N_3077,N_4855);
and U5694 (N_5694,N_582,N_2372);
nor U5695 (N_5695,N_1060,N_3624);
nand U5696 (N_5696,N_3646,N_3064);
and U5697 (N_5697,N_4724,N_2607);
xnor U5698 (N_5698,N_4066,N_3770);
xor U5699 (N_5699,N_4610,N_3765);
nand U5700 (N_5700,N_3918,N_3870);
xor U5701 (N_5701,N_2025,N_2573);
and U5702 (N_5702,N_2829,N_3489);
nand U5703 (N_5703,N_994,N_1170);
xor U5704 (N_5704,N_1197,N_4299);
or U5705 (N_5705,N_4602,N_4852);
nor U5706 (N_5706,N_437,N_2463);
nand U5707 (N_5707,N_4857,N_3861);
nand U5708 (N_5708,N_1354,N_2208);
and U5709 (N_5709,N_4817,N_4240);
nand U5710 (N_5710,N_3185,N_2264);
xnor U5711 (N_5711,N_3400,N_4854);
nand U5712 (N_5712,N_3886,N_128);
or U5713 (N_5713,N_3602,N_2336);
or U5714 (N_5714,N_2184,N_191);
nor U5715 (N_5715,N_741,N_4350);
nand U5716 (N_5716,N_4773,N_670);
nand U5717 (N_5717,N_2423,N_1516);
nand U5718 (N_5718,N_1616,N_4342);
and U5719 (N_5719,N_2980,N_4381);
and U5720 (N_5720,N_1044,N_76);
nand U5721 (N_5721,N_3934,N_2930);
or U5722 (N_5722,N_3794,N_980);
and U5723 (N_5723,N_4808,N_3232);
nor U5724 (N_5724,N_4494,N_2005);
xnor U5725 (N_5725,N_3330,N_4116);
nor U5726 (N_5726,N_586,N_3671);
and U5727 (N_5727,N_422,N_4034);
and U5728 (N_5728,N_431,N_2778);
or U5729 (N_5729,N_2572,N_2412);
or U5730 (N_5730,N_3684,N_4535);
nor U5731 (N_5731,N_4915,N_3825);
nand U5732 (N_5732,N_302,N_4309);
and U5733 (N_5733,N_2090,N_4442);
nor U5734 (N_5734,N_2043,N_327);
nor U5735 (N_5735,N_886,N_3288);
nor U5736 (N_5736,N_1500,N_3604);
nor U5737 (N_5737,N_4012,N_3223);
nand U5738 (N_5738,N_2863,N_1326);
or U5739 (N_5739,N_3371,N_1891);
xnor U5740 (N_5740,N_788,N_1375);
or U5741 (N_5741,N_106,N_2409);
nor U5742 (N_5742,N_2006,N_944);
and U5743 (N_5743,N_3974,N_165);
nand U5744 (N_5744,N_1453,N_3789);
nor U5745 (N_5745,N_3723,N_4068);
nand U5746 (N_5746,N_4846,N_1193);
nor U5747 (N_5747,N_133,N_1313);
nor U5748 (N_5748,N_2146,N_3054);
nand U5749 (N_5749,N_1074,N_4195);
nor U5750 (N_5750,N_1174,N_1316);
or U5751 (N_5751,N_4101,N_751);
nor U5752 (N_5752,N_2262,N_2613);
nand U5753 (N_5753,N_2852,N_4749);
or U5754 (N_5754,N_4241,N_3016);
nand U5755 (N_5755,N_2991,N_3750);
or U5756 (N_5756,N_4930,N_1049);
or U5757 (N_5757,N_3045,N_1913);
nand U5758 (N_5758,N_490,N_2637);
and U5759 (N_5759,N_1833,N_2571);
xor U5760 (N_5760,N_575,N_807);
and U5761 (N_5761,N_99,N_2943);
or U5762 (N_5762,N_55,N_2344);
and U5763 (N_5763,N_2431,N_3633);
and U5764 (N_5764,N_3254,N_70);
xor U5765 (N_5765,N_2937,N_674);
or U5766 (N_5766,N_4441,N_607);
xnor U5767 (N_5767,N_4083,N_953);
or U5768 (N_5768,N_1992,N_1057);
and U5769 (N_5769,N_4127,N_1103);
nor U5770 (N_5770,N_2697,N_340);
and U5771 (N_5771,N_542,N_2849);
and U5772 (N_5772,N_2065,N_965);
nor U5773 (N_5773,N_2255,N_1663);
and U5774 (N_5774,N_1468,N_3258);
nor U5775 (N_5775,N_3716,N_2925);
and U5776 (N_5776,N_4750,N_572);
xor U5777 (N_5777,N_812,N_228);
or U5778 (N_5778,N_2070,N_140);
or U5779 (N_5779,N_3296,N_2949);
nand U5780 (N_5780,N_1231,N_445);
nand U5781 (N_5781,N_9,N_2686);
nor U5782 (N_5782,N_1204,N_1937);
or U5783 (N_5783,N_49,N_3963);
nand U5784 (N_5784,N_2165,N_473);
nand U5785 (N_5785,N_4935,N_3146);
nor U5786 (N_5786,N_1834,N_1973);
or U5787 (N_5787,N_1023,N_1269);
nand U5788 (N_5788,N_3551,N_3917);
nor U5789 (N_5789,N_3477,N_1645);
and U5790 (N_5790,N_3309,N_937);
and U5791 (N_5791,N_4179,N_913);
or U5792 (N_5792,N_120,N_2668);
nand U5793 (N_5793,N_4289,N_2351);
nand U5794 (N_5794,N_220,N_214);
or U5795 (N_5795,N_3142,N_3843);
or U5796 (N_5796,N_4824,N_2559);
xor U5797 (N_5797,N_1565,N_3003);
nor U5798 (N_5798,N_4005,N_1771);
and U5799 (N_5799,N_2806,N_4169);
nor U5800 (N_5800,N_4751,N_4677);
and U5801 (N_5801,N_475,N_3585);
and U5802 (N_5802,N_1021,N_611);
nor U5803 (N_5803,N_2814,N_4668);
nand U5804 (N_5804,N_3781,N_2886);
and U5805 (N_5805,N_535,N_888);
nand U5806 (N_5806,N_3953,N_2021);
xor U5807 (N_5807,N_1953,N_1362);
or U5808 (N_5808,N_4640,N_3990);
nand U5809 (N_5809,N_1287,N_3163);
and U5810 (N_5810,N_3569,N_1899);
or U5811 (N_5811,N_2346,N_472);
or U5812 (N_5812,N_2454,N_4970);
nor U5813 (N_5813,N_1220,N_2347);
nor U5814 (N_5814,N_4721,N_2565);
and U5815 (N_5815,N_1785,N_3303);
or U5816 (N_5816,N_2893,N_392);
nor U5817 (N_5817,N_1586,N_692);
or U5818 (N_5818,N_3445,N_3252);
nand U5819 (N_5819,N_101,N_3364);
and U5820 (N_5820,N_3868,N_1240);
or U5821 (N_5821,N_1603,N_2941);
xor U5822 (N_5822,N_4293,N_4422);
nor U5823 (N_5823,N_1560,N_4546);
nand U5824 (N_5824,N_718,N_3608);
and U5825 (N_5825,N_989,N_4972);
nor U5826 (N_5826,N_4981,N_1892);
nor U5827 (N_5827,N_1694,N_2345);
or U5828 (N_5828,N_3594,N_729);
xnor U5829 (N_5829,N_2970,N_3572);
and U5830 (N_5830,N_570,N_2909);
or U5831 (N_5831,N_3141,N_4591);
and U5832 (N_5832,N_903,N_615);
nor U5833 (N_5833,N_3241,N_1317);
nand U5834 (N_5834,N_1471,N_3744);
and U5835 (N_5835,N_4512,N_1878);
xor U5836 (N_5836,N_1721,N_2705);
nand U5837 (N_5837,N_1386,N_656);
nor U5838 (N_5838,N_241,N_3949);
or U5839 (N_5839,N_3485,N_2206);
or U5840 (N_5840,N_604,N_956);
or U5841 (N_5841,N_4491,N_3152);
and U5842 (N_5842,N_2634,N_1980);
nor U5843 (N_5843,N_721,N_1755);
nor U5844 (N_5844,N_3703,N_2111);
nand U5845 (N_5845,N_176,N_1719);
and U5846 (N_5846,N_3546,N_649);
nand U5847 (N_5847,N_1485,N_486);
and U5848 (N_5848,N_121,N_2638);
nand U5849 (N_5849,N_3327,N_2513);
nand U5850 (N_5850,N_2918,N_928);
nor U5851 (N_5851,N_137,N_4028);
and U5852 (N_5852,N_4044,N_373);
nand U5853 (N_5853,N_2340,N_4628);
and U5854 (N_5854,N_4469,N_1280);
and U5855 (N_5855,N_1988,N_1118);
and U5856 (N_5856,N_2723,N_1875);
or U5857 (N_5857,N_813,N_2185);
and U5858 (N_5858,N_1820,N_2576);
nand U5859 (N_5859,N_346,N_2236);
nor U5860 (N_5860,N_2314,N_3463);
or U5861 (N_5861,N_3346,N_831);
or U5862 (N_5862,N_4963,N_2127);
and U5863 (N_5863,N_4363,N_1776);
or U5864 (N_5864,N_1233,N_3229);
nand U5865 (N_5865,N_2452,N_4258);
and U5866 (N_5866,N_1689,N_4568);
nor U5867 (N_5867,N_3458,N_4662);
nor U5868 (N_5868,N_2837,N_498);
or U5869 (N_5869,N_2061,N_2629);
nand U5870 (N_5870,N_3041,N_1267);
or U5871 (N_5871,N_4570,N_2136);
nand U5872 (N_5872,N_300,N_3504);
and U5873 (N_5873,N_2773,N_3638);
nor U5874 (N_5874,N_854,N_2667);
nor U5875 (N_5875,N_4194,N_940);
and U5876 (N_5876,N_1433,N_1819);
nor U5877 (N_5877,N_1962,N_135);
nand U5878 (N_5878,N_569,N_467);
and U5879 (N_5879,N_2525,N_177);
and U5880 (N_5880,N_798,N_3291);
nand U5881 (N_5881,N_2039,N_2261);
or U5882 (N_5882,N_971,N_2397);
or U5883 (N_5883,N_3357,N_576);
nor U5884 (N_5884,N_613,N_3540);
nand U5885 (N_5885,N_4822,N_4079);
or U5886 (N_5886,N_3619,N_4757);
nand U5887 (N_5887,N_2742,N_2898);
nand U5888 (N_5888,N_285,N_4154);
or U5889 (N_5889,N_1700,N_872);
nor U5890 (N_5890,N_3592,N_263);
or U5891 (N_5891,N_491,N_4223);
and U5892 (N_5892,N_402,N_1720);
or U5893 (N_5893,N_4795,N_2427);
nor U5894 (N_5894,N_2788,N_66);
or U5895 (N_5895,N_1752,N_1470);
nor U5896 (N_5896,N_1136,N_4400);
and U5897 (N_5897,N_740,N_2462);
nand U5898 (N_5898,N_1876,N_273);
or U5899 (N_5899,N_3020,N_2597);
and U5900 (N_5900,N_834,N_4761);
xnor U5901 (N_5901,N_2951,N_1290);
or U5902 (N_5902,N_4,N_4355);
or U5903 (N_5903,N_4000,N_3108);
nor U5904 (N_5904,N_3775,N_4205);
nand U5905 (N_5905,N_1707,N_2278);
xor U5906 (N_5906,N_3370,N_1253);
nor U5907 (N_5907,N_4990,N_2434);
or U5908 (N_5908,N_4599,N_4878);
and U5909 (N_5909,N_131,N_4137);
nand U5910 (N_5910,N_1444,N_4300);
or U5911 (N_5911,N_711,N_2768);
nor U5912 (N_5912,N_1932,N_2241);
and U5913 (N_5913,N_4617,N_3273);
or U5914 (N_5914,N_4522,N_2479);
and U5915 (N_5915,N_423,N_4953);
and U5916 (N_5916,N_4619,N_3937);
nand U5917 (N_5917,N_2975,N_997);
and U5918 (N_5918,N_4324,N_3767);
or U5919 (N_5919,N_2747,N_182);
nand U5920 (N_5920,N_4115,N_3001);
and U5921 (N_5921,N_213,N_411);
and U5922 (N_5922,N_4378,N_735);
and U5923 (N_5923,N_4585,N_3657);
nand U5924 (N_5924,N_3093,N_80);
and U5925 (N_5925,N_465,N_4758);
xor U5926 (N_5926,N_4534,N_3234);
nor U5927 (N_5927,N_307,N_1801);
or U5928 (N_5928,N_3148,N_2728);
nor U5929 (N_5929,N_4564,N_676);
or U5930 (N_5930,N_845,N_1011);
nor U5931 (N_5931,N_3199,N_506);
nand U5932 (N_5932,N_716,N_494);
nand U5933 (N_5933,N_1502,N_3353);
and U5934 (N_5934,N_2578,N_781);
nor U5935 (N_5935,N_4004,N_581);
xnor U5936 (N_5936,N_3216,N_1285);
nand U5937 (N_5937,N_360,N_1821);
and U5938 (N_5938,N_4217,N_4485);
nor U5939 (N_5939,N_4292,N_3558);
or U5940 (N_5940,N_2286,N_2780);
nand U5941 (N_5941,N_1966,N_4601);
nor U5942 (N_5942,N_2443,N_166);
or U5943 (N_5943,N_2564,N_1376);
and U5944 (N_5944,N_351,N_4859);
or U5945 (N_5945,N_2271,N_1933);
xnor U5946 (N_5946,N_3872,N_3984);
or U5947 (N_5947,N_1906,N_1569);
xor U5948 (N_5948,N_2946,N_4754);
and U5949 (N_5949,N_3536,N_4106);
or U5950 (N_5950,N_1207,N_1634);
and U5951 (N_5951,N_2872,N_1034);
and U5952 (N_5952,N_3228,N_2160);
xor U5953 (N_5953,N_602,N_1494);
and U5954 (N_5954,N_2049,N_2906);
nor U5955 (N_5955,N_458,N_1449);
nand U5956 (N_5956,N_1110,N_68);
and U5957 (N_5957,N_1322,N_4402);
nor U5958 (N_5958,N_4117,N_2982);
nand U5959 (N_5959,N_4026,N_1239);
or U5960 (N_5960,N_1480,N_2069);
nand U5961 (N_5961,N_4430,N_262);
nor U5962 (N_5962,N_2124,N_2646);
nand U5963 (N_5963,N_1058,N_2868);
and U5964 (N_5964,N_4819,N_4338);
nand U5965 (N_5965,N_2073,N_3967);
nand U5966 (N_5966,N_1134,N_190);
and U5967 (N_5967,N_3896,N_1830);
xor U5968 (N_5968,N_3729,N_3272);
nor U5969 (N_5969,N_208,N_4416);
nand U5970 (N_5970,N_4434,N_19);
nand U5971 (N_5971,N_3871,N_3008);
nor U5972 (N_5972,N_3075,N_479);
xor U5973 (N_5973,N_2033,N_239);
nand U5974 (N_5974,N_530,N_2600);
xor U5975 (N_5975,N_1087,N_4163);
nor U5976 (N_5976,N_3404,N_2990);
nor U5977 (N_5977,N_3084,N_1250);
and U5978 (N_5978,N_574,N_148);
nand U5979 (N_5979,N_2328,N_2526);
nor U5980 (N_5980,N_789,N_2839);
and U5981 (N_5981,N_4389,N_2313);
nand U5982 (N_5982,N_2114,N_2101);
nand U5983 (N_5983,N_4062,N_240);
or U5984 (N_5984,N_1668,N_1210);
nand U5985 (N_5985,N_2523,N_2560);
or U5986 (N_5986,N_704,N_1211);
xnor U5987 (N_5987,N_4731,N_1243);
nor U5988 (N_5988,N_4960,N_933);
nor U5989 (N_5989,N_438,N_484);
nor U5990 (N_5990,N_2584,N_4784);
nor U5991 (N_5991,N_525,N_4478);
and U5992 (N_5992,N_383,N_833);
and U5993 (N_5993,N_2833,N_4397);
nor U5994 (N_5994,N_2784,N_2041);
or U5995 (N_5995,N_4479,N_748);
nor U5996 (N_5996,N_2182,N_3224);
nor U5997 (N_5997,N_4515,N_3980);
or U5998 (N_5998,N_3110,N_1926);
nand U5999 (N_5999,N_4130,N_2495);
or U6000 (N_6000,N_1096,N_584);
and U6001 (N_6001,N_3154,N_1888);
xnor U6002 (N_6002,N_3758,N_4875);
nor U6003 (N_6003,N_3164,N_2831);
or U6004 (N_6004,N_4235,N_116);
nor U6005 (N_6005,N_3279,N_1517);
or U6006 (N_6006,N_2963,N_2616);
or U6007 (N_6007,N_2739,N_4227);
xor U6008 (N_6008,N_2797,N_2091);
and U6009 (N_6009,N_4679,N_2325);
nand U6010 (N_6010,N_1261,N_2680);
or U6011 (N_6011,N_1082,N_4533);
nand U6012 (N_6012,N_2343,N_3637);
and U6013 (N_6013,N_4596,N_3844);
and U6014 (N_6014,N_1711,N_4243);
xor U6015 (N_6015,N_2444,N_112);
nand U6016 (N_6016,N_1138,N_2179);
nand U6017 (N_6017,N_2762,N_881);
nand U6018 (N_6018,N_1766,N_3791);
nand U6019 (N_6019,N_91,N_1447);
nor U6020 (N_6020,N_2957,N_60);
and U6021 (N_6021,N_348,N_1941);
nor U6022 (N_6022,N_3641,N_4667);
nor U6023 (N_6023,N_103,N_1347);
or U6024 (N_6024,N_387,N_3698);
or U6025 (N_6025,N_1008,N_1467);
xor U6026 (N_6026,N_2483,N_2993);
or U6027 (N_6027,N_1463,N_832);
or U6028 (N_6028,N_924,N_4980);
nor U6029 (N_6029,N_17,N_1109);
nor U6030 (N_6030,N_2938,N_1042);
or U6031 (N_6031,N_982,N_4418);
or U6032 (N_6032,N_4544,N_4145);
and U6033 (N_6033,N_4023,N_8);
xor U6034 (N_6034,N_3393,N_3375);
and U6035 (N_6035,N_1221,N_804);
xnor U6036 (N_6036,N_3342,N_3773);
nor U6037 (N_6037,N_1241,N_1345);
nor U6038 (N_6038,N_4697,N_1678);
nand U6039 (N_6039,N_469,N_2413);
or U6040 (N_6040,N_3425,N_2707);
nor U6041 (N_6041,N_2186,N_1227);
and U6042 (N_6042,N_3282,N_3822);
nor U6043 (N_6043,N_4007,N_2879);
nand U6044 (N_6044,N_3383,N_4782);
and U6045 (N_6045,N_4823,N_2394);
or U6046 (N_6046,N_2729,N_2669);
or U6047 (N_6047,N_765,N_1777);
or U6048 (N_6048,N_1963,N_274);
nor U6049 (N_6049,N_3173,N_1512);
nor U6050 (N_6050,N_339,N_3130);
and U6051 (N_6051,N_2664,N_1781);
nand U6052 (N_6052,N_4095,N_3208);
or U6053 (N_6053,N_2916,N_596);
or U6054 (N_6054,N_3836,N_4391);
or U6055 (N_6055,N_775,N_3971);
nand U6056 (N_6056,N_502,N_4510);
nor U6057 (N_6057,N_1213,N_2088);
nor U6058 (N_6058,N_1505,N_1396);
xnor U6059 (N_6059,N_3410,N_1585);
nor U6060 (N_6060,N_3678,N_2257);
or U6061 (N_6061,N_2825,N_3055);
and U6062 (N_6062,N_3609,N_590);
or U6063 (N_6063,N_4529,N_4689);
and U6064 (N_6064,N_2731,N_4950);
xor U6065 (N_6065,N_185,N_440);
nor U6066 (N_6066,N_3685,N_3165);
and U6067 (N_6067,N_4637,N_4932);
and U6068 (N_6068,N_510,N_624);
nor U6069 (N_6069,N_4909,N_1095);
xor U6070 (N_6070,N_4245,N_4815);
or U6071 (N_6071,N_4197,N_1163);
and U6072 (N_6072,N_218,N_2381);
and U6073 (N_6073,N_3318,N_1279);
nand U6074 (N_6074,N_3192,N_1717);
nand U6075 (N_6075,N_4752,N_395);
nand U6076 (N_6076,N_2217,N_1305);
nor U6077 (N_6077,N_3338,N_4232);
nor U6078 (N_6078,N_2620,N_514);
and U6079 (N_6079,N_3230,N_2823);
or U6080 (N_6080,N_608,N_696);
nand U6081 (N_6081,N_3737,N_1053);
xnor U6082 (N_6082,N_996,N_2812);
and U6083 (N_6083,N_2299,N_1084);
nor U6084 (N_6084,N_869,N_3539);
nand U6085 (N_6085,N_1572,N_369);
or U6086 (N_6086,N_4939,N_523);
nor U6087 (N_6087,N_1437,N_528);
nand U6088 (N_6088,N_3688,N_3820);
xor U6089 (N_6089,N_4073,N_3348);
and U6090 (N_6090,N_4575,N_4856);
or U6091 (N_6091,N_3431,N_4538);
and U6092 (N_6092,N_3874,N_1786);
nor U6093 (N_6093,N_2756,N_1414);
nand U6094 (N_6094,N_1130,N_3490);
and U6095 (N_6095,N_3847,N_2148);
xor U6096 (N_6096,N_4192,N_2456);
nor U6097 (N_6097,N_1930,N_733);
or U6098 (N_6098,N_2297,N_671);
or U6099 (N_6099,N_291,N_2011);
or U6100 (N_6100,N_1022,N_4562);
nand U6101 (N_6101,N_3059,N_4831);
or U6102 (N_6102,N_1885,N_618);
nand U6103 (N_6103,N_4765,N_880);
or U6104 (N_6104,N_345,N_3499);
and U6105 (N_6105,N_1152,N_3212);
and U6106 (N_6106,N_4237,N_4052);
nor U6107 (N_6107,N_3575,N_4735);
nand U6108 (N_6108,N_4914,N_2370);
and U6109 (N_6109,N_3889,N_1451);
nor U6110 (N_6110,N_1257,N_338);
and U6111 (N_6111,N_86,N_4156);
or U6112 (N_6112,N_1939,N_4772);
and U6113 (N_6113,N_2225,N_4238);
or U6114 (N_6114,N_852,N_3428);
or U6115 (N_6115,N_3337,N_3547);
or U6116 (N_6116,N_1329,N_1425);
nand U6117 (N_6117,N_4622,N_4259);
nand U6118 (N_6118,N_1584,N_211);
nor U6119 (N_6119,N_1758,N_1893);
or U6120 (N_6120,N_4578,N_1334);
and U6121 (N_6121,N_1683,N_2591);
nor U6122 (N_6122,N_3739,N_1357);
and U6123 (N_6123,N_3017,N_896);
or U6124 (N_6124,N_477,N_1690);
nand U6125 (N_6125,N_2252,N_2430);
and U6126 (N_6126,N_67,N_504);
nor U6127 (N_6127,N_1999,N_4916);
nor U6128 (N_6128,N_1660,N_1318);
nand U6129 (N_6129,N_4659,N_1904);
nor U6130 (N_6130,N_2612,N_3599);
nor U6131 (N_6131,N_2555,N_515);
or U6132 (N_6132,N_2914,N_2135);
and U6133 (N_6133,N_3102,N_299);
nand U6134 (N_6134,N_4715,N_1070);
or U6135 (N_6135,N_3204,N_3818);
xnor U6136 (N_6136,N_2858,N_366);
or U6137 (N_6137,N_818,N_4060);
or U6138 (N_6138,N_4124,N_4285);
nand U6139 (N_6139,N_2953,N_2881);
and U6140 (N_6140,N_2169,N_4096);
and U6141 (N_6141,N_808,N_2239);
nor U6142 (N_6142,N_3573,N_3019);
and U6143 (N_6143,N_1918,N_3266);
nand U6144 (N_6144,N_1052,N_867);
and U6145 (N_6145,N_4796,N_1698);
and U6146 (N_6146,N_2030,N_4265);
nor U6147 (N_6147,N_1183,N_2700);
and U6148 (N_6148,N_4279,N_3835);
nand U6149 (N_6149,N_1959,N_3544);
nor U6150 (N_6150,N_4393,N_1555);
xnor U6151 (N_6151,N_4086,N_846);
nand U6152 (N_6152,N_2749,N_4577);
and U6153 (N_6153,N_679,N_1413);
and U6154 (N_6154,N_970,N_2196);
nor U6155 (N_6155,N_4767,N_4075);
and U6156 (N_6156,N_1391,N_567);
or U6157 (N_6157,N_1206,N_2536);
nand U6158 (N_6158,N_2854,N_2813);
xor U6159 (N_6159,N_4739,N_3105);
or U6160 (N_6160,N_2964,N_1708);
and U6161 (N_6161,N_4678,N_46);
nand U6162 (N_6162,N_1927,N_1537);
nor U6163 (N_6163,N_4087,N_2471);
nand U6164 (N_6164,N_2075,N_1214);
nand U6165 (N_6165,N_2860,N_3574);
nand U6166 (N_6166,N_1805,N_3475);
nand U6167 (N_6167,N_3171,N_3358);
and U6168 (N_6168,N_2470,N_59);
and U6169 (N_6169,N_4595,N_2274);
nor U6170 (N_6170,N_2905,N_178);
nand U6171 (N_6171,N_3256,N_2);
and U6172 (N_6172,N_4999,N_173);
and U6173 (N_6173,N_603,N_2309);
nand U6174 (N_6174,N_1536,N_4368);
nand U6175 (N_6175,N_557,N_3461);
and U6176 (N_6176,N_287,N_4298);
or U6177 (N_6177,N_599,N_1406);
nand U6178 (N_6178,N_3853,N_252);
nand U6179 (N_6179,N_1840,N_3308);
nand U6180 (N_6180,N_2231,N_407);
xnor U6181 (N_6181,N_1515,N_3221);
nor U6182 (N_6182,N_4919,N_764);
or U6183 (N_6183,N_1886,N_794);
nor U6184 (N_6184,N_1858,N_2562);
or U6185 (N_6185,N_4029,N_4180);
nor U6186 (N_6186,N_3326,N_3502);
xor U6187 (N_6187,N_2489,N_4891);
or U6188 (N_6188,N_3128,N_820);
nor U6189 (N_6189,N_4203,N_4924);
and U6190 (N_6190,N_2790,N_2942);
and U6191 (N_6191,N_2999,N_1297);
nor U6192 (N_6192,N_4261,N_2223);
nor U6193 (N_6193,N_2752,N_4655);
nand U6194 (N_6194,N_3454,N_3525);
nor U6195 (N_6195,N_1981,N_4744);
and U6196 (N_6196,N_4337,N_242);
and U6197 (N_6197,N_1412,N_3183);
or U6198 (N_6198,N_2935,N_1125);
nand U6199 (N_6199,N_957,N_1203);
or U6200 (N_6200,N_2469,N_1815);
or U6201 (N_6201,N_64,N_2304);
nor U6202 (N_6202,N_1144,N_3549);
or U6203 (N_6203,N_3505,N_4941);
nor U6204 (N_6204,N_2857,N_2227);
nand U6205 (N_6205,N_2029,N_779);
or U6206 (N_6206,N_1596,N_1782);
and U6207 (N_6207,N_3438,N_2062);
nor U6208 (N_6208,N_4966,N_2390);
or U6209 (N_6209,N_40,N_4949);
nand U6210 (N_6210,N_3813,N_2981);
and U6211 (N_6211,N_56,N_2683);
and U6212 (N_6212,N_389,N_1862);
nor U6213 (N_6213,N_3732,N_1623);
nor U6214 (N_6214,N_1088,N_1392);
nand U6215 (N_6215,N_858,N_1662);
nor U6216 (N_6216,N_3712,N_311);
nor U6217 (N_6217,N_3395,N_2908);
and U6218 (N_6218,N_1127,N_2038);
nand U6219 (N_6219,N_2967,N_4446);
nand U6220 (N_6220,N_2417,N_2972);
and U6221 (N_6221,N_1229,N_3913);
nand U6222 (N_6222,N_408,N_583);
nand U6223 (N_6223,N_1558,N_2047);
nand U6224 (N_6224,N_114,N_4528);
nor U6225 (N_6225,N_3050,N_4899);
nor U6226 (N_6226,N_1226,N_1838);
or U6227 (N_6227,N_505,N_703);
nor U6228 (N_6228,N_4554,N_1769);
nor U6229 (N_6229,N_705,N_1048);
or U6230 (N_6230,N_2791,N_4652);
and U6231 (N_6231,N_1695,N_1704);
nand U6232 (N_6232,N_1484,N_4812);
nand U6233 (N_6233,N_2948,N_4134);
nand U6234 (N_6234,N_156,N_4884);
or U6235 (N_6235,N_2996,N_2194);
nor U6236 (N_6236,N_3869,N_1633);
nand U6237 (N_6237,N_1062,N_278);
nor U6238 (N_6238,N_4113,N_4775);
xnor U6239 (N_6239,N_4861,N_3925);
xor U6240 (N_6240,N_1972,N_4683);
nor U6241 (N_6241,N_4291,N_3742);
xnor U6242 (N_6242,N_1880,N_4186);
xor U6243 (N_6243,N_3456,N_4098);
nor U6244 (N_6244,N_2647,N_3161);
and U6245 (N_6245,N_3289,N_3895);
nor U6246 (N_6246,N_2648,N_4352);
and U6247 (N_6247,N_353,N_4847);
nand U6248 (N_6248,N_2176,N_4843);
and U6249 (N_6249,N_1559,N_1967);
xnor U6250 (N_6250,N_3564,N_3727);
nand U6251 (N_6251,N_756,N_2066);
and U6252 (N_6252,N_4868,N_4143);
or U6253 (N_6253,N_4310,N_921);
or U6254 (N_6254,N_2375,N_2193);
and U6255 (N_6255,N_1800,N_4900);
nor U6256 (N_6256,N_201,N_2352);
and U6257 (N_6257,N_1112,N_2556);
nor U6258 (N_6258,N_2541,N_2414);
nand U6259 (N_6259,N_3138,N_4593);
and U6260 (N_6260,N_2904,N_4908);
nor U6261 (N_6261,N_2885,N_1881);
nor U6262 (N_6262,N_4255,N_1790);
or U6263 (N_6263,N_3283,N_3373);
and U6264 (N_6264,N_664,N_1498);
or U6265 (N_6265,N_4415,N_1732);
and U6266 (N_6266,N_3613,N_1557);
and U6267 (N_6267,N_4188,N_1283);
nand U6268 (N_6268,N_4732,N_1787);
and U6269 (N_6269,N_4620,N_2594);
nand U6270 (N_6270,N_568,N_1245);
nand U6271 (N_6271,N_450,N_4465);
or U6272 (N_6272,N_449,N_4047);
and U6273 (N_6273,N_4379,N_1868);
nor U6274 (N_6274,N_4598,N_4925);
or U6275 (N_6275,N_2376,N_1101);
nand U6276 (N_6276,N_2811,N_2821);
and U6277 (N_6277,N_2174,N_1729);
nand U6278 (N_6278,N_1296,N_1113);
nand U6279 (N_6279,N_2604,N_3151);
xnor U6280 (N_6280,N_4118,N_728);
and U6281 (N_6281,N_1384,N_2847);
nand U6282 (N_6282,N_235,N_2876);
nor U6283 (N_6283,N_2845,N_1168);
nor U6284 (N_6284,N_124,N_3449);
or U6285 (N_6285,N_4176,N_4738);
xor U6286 (N_6286,N_289,N_639);
nor U6287 (N_6287,N_960,N_2622);
or U6288 (N_6288,N_1039,N_2716);
nand U6289 (N_6289,N_1029,N_3181);
nand U6290 (N_6290,N_2665,N_3798);
and U6291 (N_6291,N_4278,N_2681);
and U6292 (N_6292,N_3006,N_1974);
xnor U6293 (N_6293,N_1822,N_2940);
or U6294 (N_6294,N_3455,N_4439);
and U6295 (N_6295,N_3500,N_1540);
and U6296 (N_6296,N_2396,N_868);
or U6297 (N_6297,N_4649,N_1680);
and U6298 (N_6298,N_4061,N_2363);
nand U6299 (N_6299,N_354,N_3215);
or U6300 (N_6300,N_4694,N_2719);
and U6301 (N_6301,N_1150,N_4256);
nand U6302 (N_6302,N_3783,N_3955);
and U6303 (N_6303,N_1620,N_308);
nand U6304 (N_6304,N_487,N_1871);
nand U6305 (N_6305,N_2547,N_1802);
and U6306 (N_6306,N_3653,N_4228);
nand U6307 (N_6307,N_2528,N_2131);
and U6308 (N_6308,N_146,N_1686);
nor U6309 (N_6309,N_4707,N_4952);
nand U6310 (N_6310,N_3086,N_3244);
nand U6311 (N_6311,N_3172,N_3322);
nor U6312 (N_6312,N_2950,N_2794);
nand U6313 (N_6313,N_2329,N_3603);
nor U6314 (N_6314,N_3827,N_2138);
nand U6315 (N_6315,N_318,N_839);
nand U6316 (N_6316,N_4643,N_61);
nand U6317 (N_6317,N_2035,N_3269);
or U6318 (N_6318,N_1089,N_3779);
nand U6319 (N_6319,N_2167,N_3960);
nand U6320 (N_6320,N_1590,N_4451);
or U6321 (N_6321,N_605,N_1702);
and U6322 (N_6322,N_1237,N_2915);
nor U6323 (N_6323,N_3610,N_2190);
nand U6324 (N_6324,N_3194,N_4177);
xor U6325 (N_6325,N_3176,N_4547);
or U6326 (N_6326,N_593,N_1395);
or U6327 (N_6327,N_1454,N_2641);
nand U6328 (N_6328,N_171,N_4360);
nor U6329 (N_6329,N_2162,N_799);
nor U6330 (N_6330,N_1014,N_2514);
nand U6331 (N_6331,N_1159,N_4514);
and U6332 (N_6332,N_4942,N_1595);
nand U6333 (N_6333,N_2510,N_2161);
nand U6334 (N_6334,N_1187,N_609);
nor U6335 (N_6335,N_4107,N_1126);
nand U6336 (N_6336,N_4055,N_1390);
or U6337 (N_6337,N_4099,N_3412);
or U6338 (N_6338,N_2057,N_2611);
and U6339 (N_6339,N_4885,N_3078);
nor U6340 (N_6340,N_4693,N_1416);
xnor U6341 (N_6341,N_1825,N_4385);
nor U6342 (N_6342,N_701,N_4603);
or U6343 (N_6343,N_3998,N_3328);
or U6344 (N_6344,N_77,N_3026);
or U6345 (N_6345,N_1692,N_3926);
nand U6346 (N_6346,N_356,N_144);
or U6347 (N_6347,N_4173,N_3384);
or U6348 (N_6348,N_3995,N_3025);
and U6349 (N_6349,N_3728,N_2947);
and U6350 (N_6350,N_1289,N_513);
nor U6351 (N_6351,N_626,N_1131);
or U6352 (N_6352,N_4281,N_3515);
or U6353 (N_6353,N_1440,N_1184);
xor U6354 (N_6354,N_322,N_2097);
or U6355 (N_6355,N_3877,N_4121);
nor U6356 (N_6356,N_2153,N_2205);
and U6357 (N_6357,N_73,N_3763);
or U6358 (N_6358,N_1986,N_2642);
nand U6359 (N_6359,N_2292,N_1969);
xnor U6360 (N_6360,N_934,N_962);
and U6361 (N_6361,N_4828,N_680);
nor U6362 (N_6362,N_2805,N_352);
and U6363 (N_6363,N_4567,N_693);
nand U6364 (N_6364,N_118,N_349);
and U6365 (N_6365,N_270,N_1847);
nor U6366 (N_6366,N_1688,N_4356);
and U6367 (N_6367,N_739,N_2958);
xnor U6368 (N_6368,N_4021,N_1848);
nand U6369 (N_6369,N_4148,N_2386);
or U6370 (N_6370,N_4172,N_2305);
nor U6371 (N_6371,N_2168,N_524);
and U6372 (N_6372,N_3508,N_4420);
or U6373 (N_6373,N_1580,N_167);
nand U6374 (N_6374,N_2270,N_4833);
or U6375 (N_6375,N_4933,N_1520);
nand U6376 (N_6376,N_1350,N_698);
nand U6377 (N_6377,N_3492,N_4685);
nor U6378 (N_6378,N_4797,N_3095);
or U6379 (N_6379,N_3632,N_350);
xnor U6380 (N_6380,N_1465,N_3557);
or U6381 (N_6381,N_4120,N_836);
xnor U6382 (N_6382,N_2566,N_2096);
and U6383 (N_6383,N_878,N_4014);
nand U6384 (N_6384,N_2453,N_824);
nor U6385 (N_6385,N_963,N_2473);
xor U6386 (N_6386,N_2761,N_2726);
nand U6387 (N_6387,N_4527,N_1436);
or U6388 (N_6388,N_1809,N_1916);
xnor U6389 (N_6389,N_1106,N_3702);
xor U6390 (N_6390,N_3552,N_464);
xor U6391 (N_6391,N_3774,N_265);
nand U6392 (N_6392,N_3951,N_3554);
nand U6393 (N_6393,N_2235,N_3651);
nor U6394 (N_6394,N_3405,N_1839);
and U6395 (N_6395,N_192,N_2326);
or U6396 (N_6396,N_3060,N_964);
nor U6397 (N_6397,N_1277,N_3989);
or U6398 (N_6398,N_1971,N_2079);
nand U6399 (N_6399,N_1228,N_3284);
or U6400 (N_6400,N_3368,N_3211);
and U6401 (N_6401,N_2424,N_2583);
and U6402 (N_6402,N_481,N_2280);
nand U6403 (N_6403,N_790,N_3733);
nor U6404 (N_6404,N_3074,N_4463);
or U6405 (N_6405,N_397,N_2945);
xor U6406 (N_6406,N_4800,N_2610);
or U6407 (N_6407,N_1452,N_3099);
xor U6408 (N_6408,N_4524,N_3942);
nor U6409 (N_6409,N_866,N_2001);
nand U6410 (N_6410,N_2071,N_3738);
and U6411 (N_6411,N_1735,N_3092);
nand U6412 (N_6412,N_2995,N_1883);
or U6413 (N_6413,N_3682,N_3752);
nand U6414 (N_6414,N_4036,N_2095);
nor U6415 (N_6415,N_2441,N_3548);
and U6416 (N_6416,N_2295,N_3012);
and U6417 (N_6417,N_343,N_254);
nand U6418 (N_6418,N_2589,N_2285);
xor U6419 (N_6419,N_4091,N_3904);
or U6420 (N_6420,N_336,N_2027);
or U6421 (N_6421,N_4995,N_1995);
nor U6422 (N_6422,N_4403,N_2128);
nand U6423 (N_6423,N_1796,N_1019);
or U6424 (N_6424,N_4871,N_1361);
nor U6425 (N_6425,N_2711,N_2828);
nor U6426 (N_6426,N_2621,N_2308);
nand U6427 (N_6427,N_2737,N_4215);
and U6428 (N_6428,N_1162,N_233);
nand U6429 (N_6429,N_3630,N_1696);
or U6430 (N_6430,N_442,N_4394);
and U6431 (N_6431,N_4523,N_3704);
or U6432 (N_6432,N_384,N_871);
or U6433 (N_6433,N_4067,N_1968);
and U6434 (N_6434,N_2067,N_519);
and U6435 (N_6435,N_1736,N_1775);
and U6436 (N_6436,N_1814,N_3044);
nand U6437 (N_6437,N_3908,N_2199);
xnor U6438 (N_6438,N_4896,N_2774);
nand U6439 (N_6439,N_1382,N_760);
and U6440 (N_6440,N_1996,N_3695);
nand U6441 (N_6441,N_492,N_4913);
and U6442 (N_6442,N_4975,N_3856);
and U6443 (N_6443,N_160,N_4825);
nand U6444 (N_6444,N_2894,N_3459);
nand U6445 (N_6445,N_2793,N_2715);
nor U6446 (N_6446,N_3131,N_2897);
or U6447 (N_6447,N_1438,N_3409);
and U6448 (N_6448,N_386,N_1823);
nor U6449 (N_6449,N_4359,N_3824);
and U6450 (N_6450,N_3819,N_493);
xnor U6451 (N_6451,N_517,N_709);
or U6452 (N_6452,N_1061,N_2024);
nand U6453 (N_6453,N_754,N_1518);
xnor U6454 (N_6454,N_292,N_4102);
nand U6455 (N_6455,N_4671,N_897);
nand U6456 (N_6456,N_2519,N_4838);
and U6457 (N_6457,N_1935,N_4501);
nor U6458 (N_6458,N_3011,N_4477);
nor U6459 (N_6459,N_3033,N_2926);
or U6460 (N_6460,N_2222,N_4957);
nor U6461 (N_6461,N_3506,N_29);
nand U6462 (N_6462,N_4305,N_1751);
nor U6463 (N_6463,N_459,N_594);
and U6464 (N_6464,N_4264,N_4277);
or U6465 (N_6465,N_4271,N_917);
nor U6466 (N_6466,N_1258,N_1728);
or U6467 (N_6467,N_3394,N_1180);
nor U6468 (N_6468,N_323,N_2476);
or U6469 (N_6469,N_333,N_848);
and U6470 (N_6470,N_534,N_4583);
and U6471 (N_6471,N_2348,N_4157);
and U6472 (N_6472,N_1612,N_2320);
or U6473 (N_6473,N_651,N_3251);
or U6474 (N_6474,N_4516,N_1756);
or U6475 (N_6475,N_1733,N_3885);
xnor U6476 (N_6476,N_2451,N_2436);
and U6477 (N_6477,N_4043,N_4862);
nand U6478 (N_6478,N_3498,N_579);
and U6479 (N_6479,N_2401,N_3631);
or U6480 (N_6480,N_3443,N_511);
nor U6481 (N_6481,N_4398,N_780);
nand U6482 (N_6482,N_2422,N_368);
nand U6483 (N_6483,N_507,N_3305);
nand U6484 (N_6484,N_1336,N_1551);
and U6485 (N_6485,N_616,N_4506);
xor U6486 (N_6486,N_4513,N_2548);
nand U6487 (N_6487,N_1368,N_1359);
nor U6488 (N_6488,N_1625,N_4645);
or U6489 (N_6489,N_2130,N_2826);
nand U6490 (N_6490,N_3377,N_2818);
xnor U6491 (N_6491,N_4994,N_3670);
or U6492 (N_6492,N_1188,N_2113);
and U6493 (N_6493,N_1739,N_2687);
and U6494 (N_6494,N_2051,N_2499);
or U6495 (N_6495,N_4517,N_911);
nand U6496 (N_6496,N_843,N_4287);
nand U6497 (N_6497,N_4556,N_4304);
nor U6498 (N_6498,N_1151,N_7);
and U6499 (N_6499,N_1333,N_1450);
xor U6500 (N_6500,N_4509,N_3866);
nand U6501 (N_6501,N_4673,N_1003);
and U6502 (N_6502,N_3298,N_3189);
nor U6503 (N_6503,N_1954,N_4774);
nand U6504 (N_6504,N_3814,N_4407);
nor U6505 (N_6505,N_26,N_4119);
and U6506 (N_6506,N_147,N_659);
nand U6507 (N_6507,N_3576,N_4290);
nor U6508 (N_6508,N_4454,N_1346);
nor U6509 (N_6509,N_810,N_110);
nor U6510 (N_6510,N_4742,N_1249);
or U6511 (N_6511,N_1900,N_470);
or U6512 (N_6512,N_4830,N_3863);
nand U6513 (N_6513,N_4129,N_3768);
and U6514 (N_6514,N_3640,N_915);
or U6515 (N_6515,N_195,N_3669);
nand U6516 (N_6516,N_1232,N_736);
nor U6517 (N_6517,N_1644,N_3800);
and U6518 (N_6518,N_2973,N_4863);
and U6519 (N_6519,N_4401,N_895);
or U6520 (N_6520,N_3472,N_1421);
nor U6521 (N_6521,N_521,N_2159);
xnor U6522 (N_6522,N_1602,N_3214);
xor U6523 (N_6523,N_4560,N_4013);
nand U6524 (N_6524,N_1286,N_2323);
nand U6525 (N_6525,N_3522,N_4123);
or U6526 (N_6526,N_499,N_1677);
and U6527 (N_6527,N_3526,N_4151);
or U6528 (N_6528,N_89,N_859);
or U6529 (N_6529,N_2129,N_3293);
and U6530 (N_6530,N_1120,N_3947);
and U6531 (N_6531,N_1291,N_2880);
nor U6532 (N_6532,N_1030,N_3122);
or U6533 (N_6533,N_3693,N_1943);
or U6534 (N_6534,N_3333,N_3801);
nand U6535 (N_6535,N_1190,N_2053);
or U6536 (N_6536,N_3809,N_977);
xor U6537 (N_6537,N_2484,N_1377);
xor U6538 (N_6538,N_1795,N_2927);
or U6539 (N_6539,N_3845,N_3280);
and U6540 (N_6540,N_744,N_2341);
xnor U6541 (N_6541,N_4642,N_3880);
and U6542 (N_6542,N_3816,N_2461);
nor U6543 (N_6543,N_2609,N_887);
nor U6544 (N_6544,N_2373,N_3726);
and U6545 (N_6545,N_1424,N_314);
and U6546 (N_6546,N_1235,N_3793);
and U6547 (N_6547,N_122,N_2447);
nand U6548 (N_6548,N_4644,N_1265);
xnor U6549 (N_6549,N_1613,N_4253);
nor U6550 (N_6550,N_3123,N_391);
xor U6551 (N_6551,N_1353,N_1325);
or U6552 (N_6552,N_1792,N_3497);
nand U6553 (N_6553,N_4152,N_3004);
and U6554 (N_6554,N_4703,N_3235);
or U6555 (N_6555,N_3263,N_2760);
nand U6556 (N_6556,N_3556,N_3313);
nand U6557 (N_6557,N_33,N_3167);
xnor U6558 (N_6558,N_1143,N_4841);
and U6559 (N_6559,N_1399,N_2327);
and U6560 (N_6560,N_4609,N_2084);
nand U6561 (N_6561,N_418,N_2366);
nand U6562 (N_6562,N_4926,N_1111);
nand U6563 (N_6563,N_1007,N_2890);
nand U6564 (N_6564,N_4968,N_1921);
and U6565 (N_6565,N_4505,N_1870);
nand U6566 (N_6566,N_3101,N_1873);
and U6567 (N_6567,N_4326,N_163);
nand U6568 (N_6568,N_234,N_1653);
xor U6569 (N_6569,N_1942,N_4866);
or U6570 (N_6570,N_306,N_1791);
xor U6571 (N_6571,N_771,N_912);
nor U6572 (N_6572,N_1409,N_1149);
and U6573 (N_6573,N_4566,N_3513);
nor U6574 (N_6574,N_2692,N_2437);
or U6575 (N_6575,N_1378,N_24);
xor U6576 (N_6576,N_2653,N_1142);
and U6577 (N_6577,N_2171,N_279);
or U6578 (N_6578,N_1073,N_2595);
nand U6579 (N_6579,N_2869,N_653);
nor U6580 (N_6580,N_4592,N_1066);
or U6581 (N_6581,N_4755,N_3109);
nor U6582 (N_6582,N_1901,N_3143);
and U6583 (N_6583,N_2698,N_4675);
xor U6584 (N_6584,N_432,N_4467);
and U6585 (N_6585,N_3938,N_2059);
nor U6586 (N_6586,N_2596,N_1574);
xor U6587 (N_6587,N_4002,N_1550);
and U6588 (N_6588,N_96,N_1811);
and U6589 (N_6589,N_2997,N_3247);
nor U6590 (N_6590,N_111,N_2266);
nor U6591 (N_6591,N_4965,N_365);
nor U6592 (N_6592,N_2956,N_4460);
nand U6593 (N_6593,N_3940,N_319);
xor U6594 (N_6594,N_4382,N_3239);
and U6595 (N_6595,N_3366,N_1807);
and U6596 (N_6596,N_961,N_786);
and U6597 (N_6597,N_811,N_1054);
nand U6598 (N_6598,N_1851,N_4408);
or U6599 (N_6599,N_1349,N_4605);
xnor U6600 (N_6600,N_4466,N_769);
and U6601 (N_6601,N_1929,N_2520);
and U6602 (N_6602,N_1842,N_757);
and U6603 (N_6603,N_4165,N_4756);
or U6604 (N_6604,N_4072,N_1348);
nor U6605 (N_6605,N_4992,N_4867);
and U6606 (N_6606,N_4222,N_2685);
nor U6607 (N_6607,N_2139,N_2358);
and U6608 (N_6608,N_4946,N_2145);
and U6609 (N_6609,N_3261,N_1360);
nor U6610 (N_6610,N_2531,N_2877);
and U6611 (N_6611,N_3580,N_2272);
nand U6612 (N_6612,N_536,N_531);
or U6613 (N_6613,N_52,N_4020);
nand U6614 (N_6614,N_4766,N_1975);
nand U6615 (N_6615,N_3985,N_3117);
and U6616 (N_6616,N_3876,N_2708);
nor U6617 (N_6617,N_3341,N_2020);
nand U6618 (N_6618,N_158,N_489);
nor U6619 (N_6619,N_2593,N_1784);
nor U6620 (N_6620,N_3250,N_3323);
nor U6621 (N_6621,N_2799,N_4413);
nand U6622 (N_6622,N_2017,N_4308);
nand U6623 (N_6623,N_4448,N_4500);
nand U6624 (N_6624,N_2118,N_4503);
and U6625 (N_6625,N_3975,N_1734);
or U6626 (N_6626,N_724,N_4984);
and U6627 (N_6627,N_1473,N_2086);
nand U6628 (N_6628,N_1164,N_2928);
and U6629 (N_6629,N_2013,N_4185);
and U6630 (N_6630,N_904,N_4033);
nand U6631 (N_6631,N_3259,N_3873);
or U6632 (N_6632,N_2400,N_434);
or U6633 (N_6633,N_2816,N_3057);
nand U6634 (N_6634,N_4912,N_2911);
xor U6635 (N_6635,N_3311,N_1863);
and U6636 (N_6636,N_2291,N_2758);
xnor U6637 (N_6637,N_363,N_2450);
nand U6638 (N_6638,N_966,N_1351);
xor U6639 (N_6639,N_699,N_4001);
and U6640 (N_6640,N_3532,N_3749);
nand U6641 (N_6641,N_3127,N_3559);
nand U6642 (N_6642,N_2037,N_4897);
nand U6643 (N_6643,N_4147,N_38);
and U6644 (N_6644,N_4549,N_2077);
and U6645 (N_6645,N_2311,N_4367);
or U6646 (N_6646,N_717,N_3645);
and U6647 (N_6647,N_1300,N_1038);
or U6648 (N_6648,N_3040,N_1077);
and U6649 (N_6649,N_2654,N_3514);
nor U6650 (N_6650,N_3691,N_1056);
nor U6651 (N_6651,N_207,N_2663);
or U6652 (N_6652,N_2511,N_2307);
nand U6653 (N_6653,N_4519,N_4600);
and U6654 (N_6654,N_2763,N_3290);
xor U6655 (N_6655,N_4539,N_1615);
nand U6656 (N_6656,N_885,N_1491);
or U6657 (N_6657,N_4741,N_2800);
nor U6658 (N_6658,N_4771,N_4633);
and U6659 (N_6659,N_3851,N_3227);
and U6660 (N_6660,N_4661,N_1826);
nor U6661 (N_6661,N_3941,N_1441);
or U6662 (N_6662,N_2293,N_4131);
nand U6663 (N_6663,N_4166,N_2582);
and U6664 (N_6664,N_2382,N_1610);
nor U6665 (N_6665,N_225,N_159);
or U6666 (N_6666,N_1299,N_403);
nand U6667 (N_6667,N_2933,N_258);
and U6668 (N_6668,N_2699,N_929);
xor U6669 (N_6669,N_3113,N_1398);
and U6670 (N_6670,N_2054,N_1407);
nor U6671 (N_6671,N_4921,N_2391);
nand U6672 (N_6672,N_3453,N_1482);
nand U6673 (N_6673,N_3391,N_3924);
and U6674 (N_6674,N_1114,N_2874);
nand U6675 (N_6675,N_179,N_4998);
or U6676 (N_6676,N_2468,N_1005);
nand U6677 (N_6677,N_4940,N_488);
and U6678 (N_6678,N_939,N_1724);
and U6679 (N_6679,N_215,N_2177);
nor U6680 (N_6680,N_4438,N_4969);
or U6681 (N_6681,N_589,N_549);
nand U6682 (N_6682,N_889,N_1107);
nor U6683 (N_6683,N_4814,N_1252);
and U6684 (N_6684,N_2770,N_4695);
and U6685 (N_6685,N_2820,N_978);
and U6686 (N_6686,N_2917,N_4221);
or U6687 (N_6687,N_1895,N_2269);
nor U6688 (N_6688,N_1292,N_2691);
or U6689 (N_6689,N_3437,N_3850);
or U6690 (N_6690,N_2250,N_1647);
nand U6691 (N_6691,N_2783,N_1753);
and U6692 (N_6692,N_1145,N_169);
or U6693 (N_6693,N_3623,N_2276);
xor U6694 (N_6694,N_3207,N_3833);
nand U6695 (N_6695,N_82,N_3220);
xnor U6696 (N_6696,N_1119,N_840);
and U6697 (N_6697,N_908,N_4934);
nand U6698 (N_6698,N_1230,N_390);
and U6699 (N_6699,N_566,N_1158);
xnor U6700 (N_6700,N_4181,N_3351);
nand U6701 (N_6701,N_509,N_4801);
nor U6702 (N_6702,N_2058,N_1315);
nor U6703 (N_6703,N_3969,N_853);
or U6704 (N_6704,N_2112,N_2357);
nor U6705 (N_6705,N_1672,N_4429);
or U6706 (N_6706,N_1803,N_1884);
and U6707 (N_6707,N_3363,N_3570);
and U6708 (N_6708,N_3759,N_4025);
or U6709 (N_6709,N_2989,N_2655);
nor U6710 (N_6710,N_4018,N_3480);
and U6711 (N_6711,N_2076,N_1894);
xor U6712 (N_6712,N_3771,N_139);
xor U6713 (N_6713,N_2538,N_3935);
or U6714 (N_6714,N_3389,N_3415);
and U6715 (N_6715,N_3365,N_4818);
and U6716 (N_6716,N_1571,N_2207);
and U6717 (N_6717,N_281,N_1479);
nand U6718 (N_6718,N_4737,N_1738);
nand U6719 (N_6719,N_3350,N_2040);
xor U6720 (N_6720,N_4902,N_247);
nand U6721 (N_6721,N_4058,N_2140);
nand U6722 (N_6722,N_399,N_1024);
nor U6723 (N_6723,N_3132,N_1160);
or U6724 (N_6724,N_2640,N_3692);
or U6725 (N_6725,N_4149,N_538);
nor U6726 (N_6726,N_3711,N_51);
nor U6727 (N_6727,N_2850,N_3281);
nand U6728 (N_6728,N_129,N_2428);
xor U6729 (N_6729,N_1554,N_3893);
nand U6730 (N_6730,N_1121,N_1439);
nand U6731 (N_6731,N_4557,N_2080);
or U6732 (N_6732,N_2855,N_2550);
nand U6733 (N_6733,N_1874,N_4424);
or U6734 (N_6734,N_1429,N_2632);
and U6735 (N_6735,N_2764,N_4125);
nand U6736 (N_6736,N_2319,N_2350);
nand U6737 (N_6737,N_3343,N_787);
and U6738 (N_6738,N_1627,N_1681);
and U6739 (N_6739,N_1503,N_2403);
or U6740 (N_6740,N_1532,N_3587);
and U6741 (N_6741,N_4443,N_2672);
and U6742 (N_6742,N_1262,N_1403);
xnor U6743 (N_6743,N_2808,N_1713);
and U6744 (N_6744,N_1780,N_4705);
nand U6745 (N_6745,N_3392,N_3321);
and U6746 (N_6746,N_1592,N_3965);
or U6747 (N_6747,N_2154,N_3879);
nor U6748 (N_6748,N_2151,N_3810);
and U6749 (N_6749,N_986,N_3910);
or U6750 (N_6750,N_2283,N_48);
nor U6751 (N_6751,N_4550,N_425);
and U6752 (N_6752,N_644,N_544);
and U6753 (N_6753,N_4267,N_932);
nor U6754 (N_6754,N_83,N_1944);
and U6755 (N_6755,N_3325,N_1816);
nor U6756 (N_6756,N_153,N_2103);
and U6757 (N_6757,N_802,N_2152);
nor U6758 (N_6758,N_1928,N_4111);
nand U6759 (N_6759,N_3285,N_4435);
or U6760 (N_6760,N_2268,N_4135);
nor U6761 (N_6761,N_629,N_2775);
nand U6762 (N_6762,N_2888,N_3268);
or U6763 (N_6763,N_3336,N_3467);
nor U6764 (N_6764,N_3894,N_4318);
and U6765 (N_6765,N_2671,N_1778);
and U6766 (N_6766,N_2561,N_712);
or U6767 (N_6767,N_1404,N_4776);
and U6768 (N_6768,N_4627,N_650);
xnor U6769 (N_6769,N_1405,N_1201);
and U6770 (N_6770,N_2590,N_767);
xor U6771 (N_6771,N_2512,N_4684);
nor U6772 (N_6772,N_3027,N_3881);
nand U6773 (N_6773,N_2772,N_4411);
and U6774 (N_6774,N_2533,N_4344);
and U6775 (N_6775,N_1857,N_1281);
nand U6776 (N_6776,N_4212,N_329);
and U6777 (N_6777,N_4962,N_1854);
nand U6778 (N_6778,N_3979,N_2175);
and U6779 (N_6779,N_3471,N_2301);
nand U6780 (N_6780,N_2581,N_1275);
nand U6781 (N_6781,N_2690,N_2195);
and U6782 (N_6782,N_1401,N_4918);
nor U6783 (N_6783,N_3675,N_4214);
or U6784 (N_6784,N_974,N_1046);
nor U6785 (N_6785,N_2288,N_501);
nor U6786 (N_6786,N_4037,N_856);
or U6787 (N_6787,N_3260,N_1946);
nor U6788 (N_6788,N_2883,N_4362);
nor U6789 (N_6789,N_1427,N_12);
and U6790 (N_6790,N_3465,N_3734);
nand U6791 (N_6791,N_2365,N_1097);
or U6792 (N_6792,N_3474,N_1426);
and U6793 (N_6793,N_3538,N_4607);
nor U6794 (N_6794,N_161,N_3421);
or U6795 (N_6795,N_3398,N_2674);
or U6796 (N_6796,N_3317,N_4093);
or U6797 (N_6797,N_898,N_3748);
nand U6798 (N_6798,N_4386,N_4967);
nor U6799 (N_6799,N_3715,N_1394);
nor U6800 (N_6800,N_3627,N_3717);
xor U6801 (N_6801,N_3807,N_3056);
or U6802 (N_6802,N_1194,N_1588);
or U6803 (N_6803,N_1047,N_268);
and U6804 (N_6804,N_3106,N_690);
nor U6805 (N_6805,N_1036,N_90);
xor U6806 (N_6806,N_2435,N_3957);
nand U6807 (N_6807,N_2330,N_1855);
or U6808 (N_6808,N_94,N_1657);
and U6809 (N_6809,N_2656,N_1339);
or U6810 (N_6810,N_1850,N_3854);
xor U6811 (N_6811,N_1301,N_864);
and U6812 (N_6812,N_4670,N_75);
xnor U6813 (N_6813,N_847,N_2244);
and U6814 (N_6814,N_1445,N_857);
nor U6815 (N_6815,N_4657,N_4760);
or U6816 (N_6816,N_4250,N_2467);
and U6817 (N_6817,N_2902,N_2659);
nand U6818 (N_6818,N_1196,N_4615);
nor U6819 (N_6819,N_1041,N_1268);
nor U6820 (N_6820,N_3629,N_1442);
and U6821 (N_6821,N_2751,N_2606);
or U6822 (N_6822,N_198,N_2254);
xnor U6823 (N_6823,N_4314,N_3562);
xnor U6824 (N_6824,N_2599,N_337);
or U6825 (N_6825,N_1064,N_4050);
or U6826 (N_6826,N_2920,N_1607);
xor U6827 (N_6827,N_4874,N_1757);
or U6828 (N_6828,N_1388,N_2754);
nor U6829 (N_6829,N_1276,N_4781);
or U6830 (N_6830,N_884,N_3803);
nor U6831 (N_6831,N_1831,N_1747);
or U6832 (N_6832,N_4349,N_1674);
nand U6833 (N_6833,N_1856,N_4826);
nand U6834 (N_6834,N_1446,N_1415);
nand U6835 (N_6835,N_2901,N_3072);
or U6836 (N_6836,N_2256,N_3145);
or U6837 (N_6837,N_4476,N_3757);
and U6838 (N_6838,N_4376,N_725);
or U6839 (N_6839,N_2042,N_4251);
nand U6840 (N_6840,N_3401,N_1234);
nor U6841 (N_6841,N_1864,N_2701);
nor U6842 (N_6842,N_2221,N_3658);
xnor U6843 (N_6843,N_1687,N_3804);
and U6844 (N_6844,N_3660,N_3005);
or U6845 (N_6845,N_1664,N_1566);
and U6846 (N_6846,N_2290,N_1295);
and U6847 (N_6847,N_1270,N_1611);
nand U6848 (N_6848,N_3039,N_264);
and U6849 (N_6849,N_3121,N_577);
nor U6850 (N_6850,N_256,N_3992);
or U6851 (N_6851,N_1705,N_4690);
nand U6852 (N_6852,N_1914,N_3408);
nor U6853 (N_6853,N_3429,N_4246);
xnor U6854 (N_6854,N_14,N_1665);
or U6855 (N_6855,N_1749,N_882);
xnor U6856 (N_6856,N_1422,N_4804);
nand U6857 (N_6857,N_22,N_92);
or U6858 (N_6858,N_3672,N_1684);
nor U6859 (N_6859,N_3769,N_1167);
nand U6860 (N_6860,N_4837,N_2429);
nor U6861 (N_6861,N_1523,N_3427);
and U6862 (N_6862,N_2158,N_4191);
and U6863 (N_6863,N_3680,N_4654);
or U6864 (N_6864,N_2643,N_1837);
nand U6865 (N_6865,N_2534,N_3379);
nand U6866 (N_6866,N_1905,N_4056);
and U6867 (N_6867,N_2163,N_2782);
or U6868 (N_6868,N_1606,N_3565);
and U6869 (N_6869,N_4456,N_4802);
or U6870 (N_6870,N_4726,N_1726);
or U6871 (N_6871,N_2682,N_2164);
nand U6872 (N_6872,N_3035,N_3469);
nor U6873 (N_6873,N_727,N_3213);
xnor U6874 (N_6874,N_3022,N_1658);
or U6875 (N_6875,N_4869,N_2298);
nor U6876 (N_6876,N_2246,N_2507);
xor U6877 (N_6877,N_1659,N_1556);
or U6878 (N_6878,N_4842,N_482);
nor U6879 (N_6879,N_2442,N_835);
nor U6880 (N_6880,N_4122,N_3683);
nor U6881 (N_6881,N_10,N_3170);
and U6882 (N_6882,N_3792,N_710);
nand U6883 (N_6883,N_2684,N_1098);
nor U6884 (N_6884,N_4110,N_1581);
and U6885 (N_6885,N_3674,N_3897);
or U6886 (N_6886,N_838,N_2243);
and U6887 (N_6887,N_1767,N_1709);
nand U6888 (N_6888,N_2965,N_1529);
and U6889 (N_6889,N_3246,N_1774);
and U6890 (N_6890,N_4297,N_1091);
nand U6891 (N_6891,N_1456,N_1461);
and U6892 (N_6892,N_2984,N_3578);
nand U6893 (N_6893,N_1737,N_1638);
nand U6894 (N_6894,N_2418,N_3299);
nor U6895 (N_6895,N_2102,N_2249);
nand U6896 (N_6896,N_1075,N_4104);
or U6897 (N_6897,N_637,N_2891);
or U6898 (N_6898,N_4574,N_3527);
nand U6899 (N_6899,N_4898,N_4789);
and U6900 (N_6900,N_3778,N_4496);
or U6901 (N_6901,N_3037,N_3745);
nor U6902 (N_6902,N_625,N_371);
and U6903 (N_6903,N_2725,N_4786);
or U6904 (N_6904,N_1189,N_4938);
nand U6905 (N_6905,N_443,N_805);
nor U6906 (N_6906,N_4164,N_3042);
nor U6907 (N_6907,N_2961,N_1139);
or U6908 (N_6908,N_2979,N_694);
nand U6909 (N_6909,N_941,N_4552);
nand U6910 (N_6910,N_622,N_4526);
xor U6911 (N_6911,N_2518,N_421);
and U6912 (N_6912,N_4472,N_4162);
or U6913 (N_6913,N_861,N_174);
nand U6914 (N_6914,N_429,N_2842);
and U6915 (N_6915,N_4540,N_2355);
nand U6916 (N_6916,N_4410,N_3589);
xor U6917 (N_6917,N_4328,N_4109);
and U6918 (N_6918,N_1383,N_4019);
or U6919 (N_6919,N_4958,N_109);
nor U6920 (N_6920,N_4976,N_417);
and U6921 (N_6921,N_1872,N_3264);
nand U6922 (N_6922,N_3776,N_3460);
nor U6923 (N_6923,N_412,N_2181);
and U6924 (N_6924,N_3159,N_2439);
nand U6925 (N_6925,N_2032,N_1352);
xor U6926 (N_6926,N_2237,N_2486);
and U6927 (N_6927,N_2119,N_3523);
nand U6928 (N_6928,N_3571,N_3584);
and U6929 (N_6929,N_288,N_4989);
nor U6930 (N_6930,N_1251,N_4225);
nor U6931 (N_6931,N_164,N_4269);
and U6932 (N_6932,N_1497,N_1808);
nand U6933 (N_6933,N_2490,N_1501);
and U6934 (N_6934,N_1513,N_4319);
and U6935 (N_6935,N_2360,N_457);
and U6936 (N_6936,N_1731,N_1961);
nand U6937 (N_6937,N_1012,N_1156);
xnor U6938 (N_6938,N_84,N_3124);
nand U6939 (N_6939,N_559,N_1509);
or U6940 (N_6940,N_2807,N_732);
nand U6941 (N_6941,N_200,N_3354);
nor U6942 (N_6942,N_2123,N_901);
xor U6943 (N_6943,N_4333,N_3411);
or U6944 (N_6944,N_4834,N_3676);
or U6945 (N_6945,N_4286,N_4428);
nand U6946 (N_6946,N_1754,N_2781);
nand U6947 (N_6947,N_619,N_3115);
and U6948 (N_6948,N_763,N_526);
or U6949 (N_6949,N_4883,N_3806);
nor U6950 (N_6950,N_2284,N_4159);
and U6951 (N_6951,N_4254,N_4404);
nand U6952 (N_6952,N_4209,N_3796);
xnor U6953 (N_6953,N_4112,N_876);
nor U6954 (N_6954,N_3079,N_4490);
nand U6955 (N_6955,N_410,N_4565);
or U6956 (N_6956,N_474,N_57);
nor U6957 (N_6957,N_2046,N_2045);
nand U6958 (N_6958,N_132,N_4923);
nand U6959 (N_6959,N_3784,N_398);
nor U6960 (N_6960,N_784,N_2587);
and U6961 (N_6961,N_4911,N_1191);
and U6962 (N_6962,N_1105,N_683);
nor U6963 (N_6963,N_1067,N_3178);
and U6964 (N_6964,N_1015,N_1576);
and U6965 (N_6965,N_1887,N_4571);
and U6966 (N_6966,N_1922,N_2884);
or U6967 (N_6967,N_3903,N_1810);
nand U6968 (N_6968,N_4587,N_2801);
and U6969 (N_6969,N_115,N_2522);
nand U6970 (N_6970,N_4736,N_3956);
nand U6971 (N_6971,N_1323,N_2472);
xnor U6972 (N_6972,N_1254,N_2455);
and U6973 (N_6973,N_1727,N_4648);
xor U6974 (N_6974,N_992,N_3314);
nor U6975 (N_6975,N_2969,N_4827);
nand U6976 (N_6976,N_3066,N_2267);
nand U6977 (N_6977,N_4982,N_4296);
nand U6978 (N_6978,N_826,N_1639);
or U6979 (N_6979,N_2204,N_1598);
xnor U6980 (N_6980,N_2617,N_972);
and U6981 (N_6981,N_3858,N_2630);
xnor U6982 (N_6982,N_2415,N_4336);
nor U6983 (N_6983,N_662,N_3945);
or U6984 (N_6984,N_444,N_1284);
nand U6985 (N_6985,N_4788,N_4480);
and U6986 (N_6986,N_1293,N_3686);
and U6987 (N_6987,N_2420,N_547);
nand U6988 (N_6988,N_453,N_993);
or U6989 (N_6989,N_3826,N_2378);
and U6990 (N_6990,N_248,N_3614);
nor U6991 (N_6991,N_2494,N_1636);
nand U6992 (N_6992,N_3883,N_2603);
and U6993 (N_6993,N_2389,N_1430);
or U6994 (N_6994,N_2209,N_4582);
or U6995 (N_6995,N_238,N_2478);
nand U6996 (N_6996,N_1964,N_4920);
and U6997 (N_6997,N_476,N_3083);
and U6998 (N_6998,N_3177,N_564);
and U6999 (N_6999,N_4704,N_3149);
nand U7000 (N_7000,N_2574,N_3842);
and U7001 (N_7001,N_3689,N_1272);
nand U7002 (N_7002,N_2544,N_916);
nand U7003 (N_7003,N_1760,N_290);
and U7004 (N_7004,N_3464,N_4031);
nor U7005 (N_7005,N_4481,N_1631);
nand U7006 (N_7006,N_2971,N_427);
nor U7007 (N_7007,N_2678,N_3681);
nand U7008 (N_7008,N_4716,N_3307);
nand U7009 (N_7009,N_4987,N_1198);
nand U7010 (N_7010,N_463,N_3344);
xor U7011 (N_7011,N_2673,N_4085);
nand U7012 (N_7012,N_2986,N_3479);
nor U7013 (N_7013,N_4315,N_713);
and U7014 (N_7014,N_3061,N_3764);
nand U7015 (N_7015,N_1006,N_2985);
or U7016 (N_7016,N_4184,N_3849);
nand U7017 (N_7017,N_4475,N_3329);
or U7018 (N_7018,N_792,N_1169);
nor U7019 (N_7019,N_4849,N_3933);
nor U7020 (N_7020,N_522,N_783);
xor U7021 (N_7021,N_2099,N_1743);
nor U7022 (N_7022,N_1682,N_2704);
nor U7023 (N_7023,N_168,N_551);
nand U7024 (N_7024,N_4624,N_2334);
nor U7025 (N_7025,N_41,N_4302);
nor U7026 (N_7026,N_2172,N_1593);
nor U7027 (N_7027,N_2052,N_4361);
or U7028 (N_7028,N_3182,N_837);
and U7029 (N_7029,N_2779,N_1654);
and U7030 (N_7030,N_691,N_2618);
xnor U7031 (N_7031,N_2068,N_3786);
nand U7032 (N_7032,N_2602,N_2922);
nand U7033 (N_7033,N_1989,N_2048);
and U7034 (N_7034,N_555,N_2866);
or U7035 (N_7035,N_3766,N_4231);
xnor U7036 (N_7036,N_806,N_2744);
nor U7037 (N_7037,N_988,N_1699);
or U7038 (N_7038,N_4520,N_3135);
nor U7039 (N_7039,N_4997,N_2247);
nand U7040 (N_7040,N_2936,N_828);
nor U7041 (N_7041,N_3927,N_2706);
nand U7042 (N_7042,N_3652,N_1312);
xnor U7043 (N_7043,N_3233,N_3785);
or U7044 (N_7044,N_3295,N_3790);
or U7045 (N_7045,N_809,N_2387);
nand U7046 (N_7046,N_3788,N_1998);
xor U7047 (N_7047,N_4341,N_612);
nand U7048 (N_7048,N_3909,N_3265);
xnor U7049 (N_7049,N_495,N_1896);
nand U7050 (N_7050,N_462,N_4799);
or U7051 (N_7051,N_2787,N_2676);
and U7052 (N_7052,N_4696,N_4886);
nand U7053 (N_7053,N_4907,N_722);
and U7054 (N_7054,N_606,N_3103);
nor U7055 (N_7055,N_702,N_3555);
and U7056 (N_7056,N_4030,N_3722);
nand U7057 (N_7057,N_4728,N_172);
nand U7058 (N_7058,N_320,N_2545);
nor U7059 (N_7059,N_3249,N_1216);
nor U7060 (N_7060,N_1147,N_4094);
xor U7061 (N_7061,N_2853,N_4525);
and U7062 (N_7062,N_1055,N_4080);
or U7063 (N_7063,N_4955,N_3593);
nor U7064 (N_7064,N_4903,N_4594);
nand U7065 (N_7065,N_3994,N_4977);
or U7066 (N_7066,N_4530,N_3315);
xor U7067 (N_7067,N_3731,N_1469);
or U7068 (N_7068,N_1742,N_2992);
nand U7069 (N_7069,N_342,N_3058);
nor U7070 (N_7070,N_2083,N_2149);
nor U7071 (N_7071,N_3360,N_1994);
or U7072 (N_7072,N_4492,N_250);
nor U7073 (N_7073,N_1622,N_2539);
or U7074 (N_7074,N_244,N_1675);
nor U7075 (N_7075,N_2815,N_2259);
nor U7076 (N_7076,N_4218,N_4572);
nand U7077 (N_7077,N_1750,N_3667);
nand U7078 (N_7078,N_1460,N_2569);
and U7079 (N_7079,N_3361,N_3015);
nand U7080 (N_7080,N_2929,N_669);
nor U7081 (N_7081,N_1624,N_4332);
xor U7082 (N_7082,N_3892,N_1092);
nor U7083 (N_7083,N_1010,N_3267);
and U7084 (N_7084,N_3180,N_1741);
nand U7085 (N_7085,N_2287,N_2126);
and U7086 (N_7086,N_817,N_2147);
xor U7087 (N_7087,N_2657,N_3225);
and U7088 (N_7088,N_3278,N_1086);
and U7089 (N_7089,N_3860,N_27);
nand U7090 (N_7090,N_1978,N_4141);
or U7091 (N_7091,N_4016,N_2714);
nor U7092 (N_7092,N_3126,N_4608);
nand U7093 (N_7093,N_3156,N_3939);
nand U7094 (N_7094,N_1304,N_1431);
nor U7095 (N_7095,N_1632,N_1650);
and U7096 (N_7096,N_155,N_3076);
xnor U7097 (N_7097,N_2289,N_364);
or U7098 (N_7098,N_2546,N_2750);
or U7099 (N_7099,N_1794,N_1179);
nor U7100 (N_7100,N_3902,N_2371);
nor U7101 (N_7101,N_1260,N_4845);
nand U7102 (N_7102,N_3628,N_20);
nand U7103 (N_7103,N_2628,N_623);
or U7104 (N_7104,N_4791,N_2506);
or U7105 (N_7105,N_3436,N_1072);
and U7106 (N_7106,N_621,N_2362);
and U7107 (N_7107,N_2939,N_3324);
nor U7108 (N_7108,N_1068,N_2488);
nor U7109 (N_7109,N_3418,N_3887);
or U7110 (N_7110,N_2296,N_2405);
xnor U7111 (N_7111,N_1917,N_1411);
and U7112 (N_7112,N_2568,N_3049);
and U7113 (N_7113,N_1990,N_2474);
xnor U7114 (N_7114,N_2738,N_1340);
or U7115 (N_7115,N_3690,N_79);
nand U7116 (N_7116,N_1745,N_3158);
or U7117 (N_7117,N_2627,N_2624);
or U7118 (N_7118,N_3374,N_2122);
and U7119 (N_7119,N_3190,N_2421);
nor U7120 (N_7120,N_791,N_1835);
nor U7121 (N_7121,N_4295,N_973);
xor U7122 (N_7122,N_2809,N_1076);
or U7123 (N_7123,N_892,N_4211);
nand U7124 (N_7124,N_3417,N_1001);
nand U7125 (N_7125,N_3993,N_2722);
nand U7126 (N_7126,N_2100,N_1208);
or U7127 (N_7127,N_4706,N_2567);
and U7128 (N_7128,N_800,N_154);
nor U7129 (N_7129,N_3656,N_400);
or U7130 (N_7130,N_3446,N_1535);
and U7131 (N_7131,N_1812,N_4436);
nor U7132 (N_7132,N_4559,N_503);
or U7133 (N_7133,N_855,N_1466);
nand U7134 (N_7134,N_4035,N_3601);
xor U7135 (N_7135,N_3972,N_4128);
nor U7136 (N_7136,N_245,N_2132);
and U7137 (N_7137,N_4334,N_2658);
nor U7138 (N_7138,N_3530,N_752);
xor U7139 (N_7139,N_102,N_645);
or U7140 (N_7140,N_393,N_556);
nor U7141 (N_7141,N_3218,N_591);
nor U7142 (N_7142,N_4894,N_4320);
or U7143 (N_7143,N_2356,N_3286);
or U7144 (N_7144,N_3052,N_682);
and U7145 (N_7145,N_4879,N_803);
nand U7146 (N_7146,N_1546,N_3828);
and U7147 (N_7147,N_2180,N_1956);
and U7148 (N_7148,N_4200,N_598);
and U7149 (N_7149,N_4331,N_2425);
or U7150 (N_7150,N_4249,N_3029);
nor U7151 (N_7151,N_2015,N_2233);
nor U7152 (N_7152,N_1356,N_1866);
and U7153 (N_7153,N_1202,N_899);
and U7154 (N_7154,N_3242,N_3701);
nand U7155 (N_7155,N_3297,N_3133);
nand U7156 (N_7156,N_2703,N_3347);
or U7157 (N_7157,N_1773,N_2487);
nor U7158 (N_7158,N_4621,N_3274);
and U7159 (N_7159,N_1577,N_4216);
or U7160 (N_7160,N_737,N_409);
or U7161 (N_7161,N_1085,N_3930);
and U7162 (N_7162,N_628,N_3857);
or U7163 (N_7163,N_893,N_3595);
and U7164 (N_7164,N_4364,N_3245);
and U7165 (N_7165,N_283,N_2796);
and U7166 (N_7166,N_4931,N_2125);
or U7167 (N_7167,N_1474,N_3420);
nor U7168 (N_7168,N_4108,N_4681);
nand U7169 (N_7169,N_4864,N_595);
nand U7170 (N_7170,N_2592,N_580);
and U7171 (N_7171,N_4718,N_1949);
nor U7172 (N_7172,N_2766,N_3442);
nor U7173 (N_7173,N_1370,N_4794);
nor U7174 (N_7174,N_3139,N_560);
nor U7175 (N_7175,N_3668,N_313);
and U7176 (N_7176,N_4399,N_3751);
or U7177 (N_7177,N_4508,N_3520);
nor U7178 (N_7178,N_3662,N_414);
nand U7179 (N_7179,N_4371,N_936);
or U7180 (N_7180,N_3946,N_3760);
or U7181 (N_7181,N_406,N_1209);
xnor U7182 (N_7182,N_2364,N_1527);
nor U7183 (N_7183,N_3100,N_1115);
and U7184 (N_7184,N_1400,N_2527);
or U7185 (N_7185,N_2709,N_4536);
and U7186 (N_7186,N_4971,N_3125);
nand U7187 (N_7187,N_2921,N_4171);
xor U7188 (N_7188,N_382,N_1919);
nor U7189 (N_7189,N_3970,N_4905);
nor U7190 (N_7190,N_3466,N_3457);
nand U7191 (N_7191,N_2230,N_3452);
xnor U7192 (N_7192,N_98,N_890);
and U7193 (N_7193,N_4686,N_2856);
or U7194 (N_7194,N_30,N_2213);
nand U7195 (N_7195,N_3635,N_2014);
and U7196 (N_7196,N_3639,N_1337);
nor U7197 (N_7197,N_430,N_1331);
nor U7198 (N_7198,N_4581,N_2843);
and U7199 (N_7199,N_1669,N_2875);
nand U7200 (N_7200,N_1762,N_875);
nand U7201 (N_7201,N_34,N_3419);
xor U7202 (N_7202,N_991,N_3648);
nor U7203 (N_7203,N_471,N_2416);
nor U7204 (N_7204,N_4011,N_562);
or U7205 (N_7205,N_2745,N_4974);
nand U7206 (N_7206,N_3812,N_4234);
nand U7207 (N_7207,N_4936,N_1652);
nand U7208 (N_7208,N_276,N_1813);
or U7209 (N_7209,N_150,N_4088);
and U7210 (N_7210,N_1397,N_53);
nand U7211 (N_7211,N_518,N_2460);
nor U7212 (N_7212,N_2107,N_4947);
or U7213 (N_7213,N_455,N_1629);
nor U7214 (N_7214,N_4542,N_500);
xor U7215 (N_7215,N_1718,N_3991);
nor U7216 (N_7216,N_665,N_3413);
or U7217 (N_7217,N_2498,N_4369);
nand U7218 (N_7218,N_548,N_2836);
or U7219 (N_7219,N_1341,N_1575);
nor U7220 (N_7220,N_4226,N_3226);
or U7221 (N_7221,N_4701,N_3140);
and U7222 (N_7222,N_688,N_187);
nor U7223 (N_7223,N_4161,N_657);
nor U7224 (N_7224,N_1882,N_1000);
nor U7225 (N_7225,N_88,N_4046);
or U7226 (N_7226,N_2445,N_1129);
nor U7227 (N_7227,N_152,N_1408);
nand U7228 (N_7228,N_1410,N_2735);
xnor U7229 (N_7229,N_113,N_4343);
and U7230 (N_7230,N_1951,N_3023);
nor U7231 (N_7231,N_3898,N_259);
or U7232 (N_7232,N_3080,N_1614);
nor U7233 (N_7233,N_2277,N_3441);
nand U7234 (N_7234,N_183,N_344);
or U7235 (N_7235,N_955,N_385);
nand U7236 (N_7236,N_4322,N_2170);
and U7237 (N_7237,N_3262,N_3205);
nor U7238 (N_7238,N_1259,N_271);
or U7239 (N_7239,N_367,N_2736);
or U7240 (N_7240,N_1579,N_4944);
or U7241 (N_7241,N_4081,N_44);
xor U7242 (N_7242,N_967,N_3082);
nand U7243 (N_7243,N_1748,N_4518);
or U7244 (N_7244,N_3622,N_3098);
and U7245 (N_7245,N_2056,N_2008);
and U7246 (N_7246,N_404,N_69);
or U7247 (N_7247,N_3372,N_4003);
and U7248 (N_7248,N_1483,N_4865);
and U7249 (N_7249,N_4665,N_2466);
xnor U7250 (N_7250,N_1667,N_16);
and U7251 (N_7251,N_15,N_753);
and U7252 (N_7252,N_1402,N_87);
and U7253 (N_7253,N_1865,N_2036);
nand U7254 (N_7254,N_1069,N_326);
xnor U7255 (N_7255,N_4961,N_1646);
and U7256 (N_7256,N_4488,N_4870);
or U7257 (N_7257,N_3644,N_315);
or U7258 (N_7258,N_3094,N_1538);
nor U7259 (N_7259,N_2023,N_4986);
nor U7260 (N_7260,N_3626,N_3406);
and U7261 (N_7261,N_3447,N_293);
nand U7262 (N_7262,N_4626,N_1263);
nand U7263 (N_7263,N_4461,N_2446);
nand U7264 (N_7264,N_947,N_4054);
or U7265 (N_7265,N_4457,N_4777);
or U7266 (N_7266,N_1478,N_1601);
or U7267 (N_7267,N_2134,N_224);
or U7268 (N_7268,N_1617,N_303);
nor U7269 (N_7269,N_3198,N_1744);
or U7270 (N_7270,N_2900,N_1303);
and U7271 (N_7271,N_3618,N_1493);
nand U7272 (N_7272,N_1797,N_663);
nor U7273 (N_7273,N_361,N_1897);
nand U7274 (N_7274,N_3916,N_3802);
nor U7275 (N_7275,N_2554,N_2197);
xor U7276 (N_7276,N_2976,N_42);
nand U7277 (N_7277,N_652,N_3531);
nand U7278 (N_7278,N_2631,N_426);
nand U7279 (N_7279,N_3713,N_1591);
nand U7280 (N_7280,N_196,N_4421);
and U7281 (N_7281,N_2440,N_675);
or U7282 (N_7282,N_2662,N_4347);
nor U7283 (N_7283,N_1853,N_823);
nand U7284 (N_7284,N_4632,N_381);
or U7285 (N_7285,N_2713,N_533);
and U7286 (N_7286,N_2408,N_4816);
nand U7287 (N_7287,N_4313,N_1002);
and U7288 (N_7288,N_1218,N_4709);
nor U7289 (N_7289,N_3579,N_3332);
or U7290 (N_7290,N_170,N_93);
nor U7291 (N_7291,N_123,N_3501);
xor U7292 (N_7292,N_2959,N_11);
and U7293 (N_7293,N_2028,N_1525);
or U7294 (N_7294,N_357,N_4636);
or U7295 (N_7295,N_4979,N_4063);
nor U7296 (N_7296,N_4717,N_1171);
and U7297 (N_7297,N_2817,N_4700);
and U7298 (N_7298,N_2496,N_874);
nand U7299 (N_7299,N_1128,N_1381);
or U7300 (N_7300,N_4409,N_2798);
xor U7301 (N_7301,N_2987,N_585);
or U7302 (N_7302,N_375,N_3236);
nor U7303 (N_7303,N_1365,N_1215);
nand U7304 (N_7304,N_968,N_71);
nand U7305 (N_7305,N_0,N_2748);
or U7306 (N_7306,N_4224,N_3340);
nand U7307 (N_7307,N_3905,N_958);
xor U7308 (N_7308,N_4780,N_3710);
and U7309 (N_7309,N_2577,N_2120);
nand U7310 (N_7310,N_209,N_4748);
xor U7311 (N_7311,N_1524,N_3355);
nand U7312 (N_7312,N_4964,N_447);
nor U7313 (N_7313,N_2143,N_4658);
nor U7314 (N_7314,N_2481,N_2871);
and U7315 (N_7315,N_1970,N_4710);
and U7316 (N_7316,N_1716,N_1712);
nand U7317 (N_7317,N_301,N_1948);
xnor U7318 (N_7318,N_4316,N_774);
or U7319 (N_7319,N_2769,N_4282);
nand U7320 (N_7320,N_3089,N_3382);
xor U7321 (N_7321,N_1924,N_1117);
xnor U7322 (N_7322,N_2551,N_3696);
nor U7323 (N_7323,N_3753,N_3606);
nor U7324 (N_7324,N_1371,N_643);
nor U7325 (N_7325,N_3091,N_4614);
nand U7326 (N_7326,N_4740,N_1691);
or U7327 (N_7327,N_396,N_1153);
nor U7328 (N_7328,N_379,N_2912);
and U7329 (N_7329,N_3111,N_3478);
nor U7330 (N_7330,N_1192,N_2924);
xnor U7331 (N_7331,N_3134,N_4682);
nand U7332 (N_7332,N_2433,N_3524);
nor U7333 (N_7333,N_3432,N_1369);
nand U7334 (N_7334,N_954,N_3287);
and U7335 (N_7335,N_134,N_4714);
nand U7336 (N_7336,N_923,N_3943);
nand U7337 (N_7337,N_2579,N_636);
or U7338 (N_7338,N_851,N_4301);
xor U7339 (N_7339,N_734,N_3597);
xnor U7340 (N_7340,N_1563,N_3725);
or U7341 (N_7341,N_58,N_4444);
xnor U7342 (N_7342,N_1789,N_2200);
and U7343 (N_7343,N_793,N_4590);
nand U7344 (N_7344,N_1568,N_4543);
or U7345 (N_7345,N_3349,N_3582);
nand U7346 (N_7346,N_3617,N_3188);
xor U7347 (N_7347,N_1903,N_777);
or U7348 (N_7348,N_3191,N_689);
and U7349 (N_7349,N_2834,N_3677);
nor U7350 (N_7350,N_3561,N_1154);
xor U7351 (N_7351,N_1519,N_3450);
and U7352 (N_7352,N_3444,N_1423);
or U7353 (N_7353,N_4521,N_3586);
and U7354 (N_7354,N_976,N_3010);
nor U7355 (N_7355,N_45,N_3036);
and U7356 (N_7356,N_3179,N_1761);
or U7357 (N_7357,N_2198,N_1759);
and U7358 (N_7358,N_995,N_1693);
nand U7359 (N_7359,N_4687,N_3988);
nand U7360 (N_7360,N_660,N_4038);
and U7361 (N_7361,N_4573,N_1487);
xnor U7362 (N_7362,N_1957,N_2104);
or U7363 (N_7363,N_819,N_2337);
and U7364 (N_7364,N_2335,N_3277);
and U7365 (N_7365,N_3510,N_3650);
or U7366 (N_7366,N_2540,N_1458);
nand U7367 (N_7367,N_4910,N_2892);
nor U7368 (N_7368,N_3976,N_2626);
nor U7369 (N_7369,N_3136,N_1278);
or U7370 (N_7370,N_1604,N_1958);
xor U7371 (N_7371,N_1715,N_1643);
nor U7372 (N_7372,N_2743,N_3209);
nand U7373 (N_7373,N_332,N_3756);
nor U7374 (N_7374,N_3434,N_863);
and U7375 (N_7375,N_3655,N_1934);
and U7376 (N_7376,N_229,N_3071);
or U7377 (N_7377,N_4357,N_1205);
nand U7378 (N_7378,N_62,N_4973);
nand U7379 (N_7379,N_678,N_1843);
or U7380 (N_7380,N_130,N_1043);
and U7381 (N_7381,N_138,N_2303);
nand U7382 (N_7382,N_3144,N_3929);
nor U7383 (N_7383,N_3362,N_4948);
nor U7384 (N_7384,N_1640,N_2802);
nor U7385 (N_7385,N_4248,N_347);
or U7386 (N_7386,N_631,N_424);
nand U7387 (N_7387,N_1173,N_2349);
or U7388 (N_7388,N_4474,N_4978);
or U7389 (N_7389,N_1533,N_65);
nor U7390 (N_7390,N_4858,N_1094);
nand U7391 (N_7391,N_3829,N_1104);
or U7392 (N_7392,N_2919,N_3088);
and U7393 (N_7393,N_3276,N_4274);
nand U7394 (N_7394,N_3997,N_3496);
or U7395 (N_7395,N_126,N_554);
nand U7396 (N_7396,N_743,N_1051);
and U7397 (N_7397,N_3687,N_136);
nor U7398 (N_7398,N_2810,N_3966);
or U7399 (N_7399,N_2300,N_1578);
or U7400 (N_7400,N_2983,N_4082);
nor U7401 (N_7401,N_1836,N_2116);
or U7402 (N_7402,N_3754,N_1859);
or U7403 (N_7403,N_4646,N_2822);
nand U7404 (N_7404,N_3201,N_104);
or U7405 (N_7405,N_188,N_3890);
nand U7406 (N_7406,N_2060,N_571);
nor U7407 (N_7407,N_480,N_3706);
or U7408 (N_7408,N_2004,N_3999);
or U7409 (N_7409,N_4793,N_1983);
nand U7410 (N_7410,N_4541,N_269);
xnor U7411 (N_7411,N_648,N_4618);
nor U7412 (N_7412,N_4906,N_2465);
and U7413 (N_7413,N_1013,N_3912);
and U7414 (N_7414,N_4959,N_3862);
or U7415 (N_7415,N_4078,N_952);
and U7416 (N_7416,N_1541,N_4354);
and U7417 (N_7417,N_2910,N_4676);
and U7418 (N_7418,N_95,N_2712);
or U7419 (N_7419,N_3511,N_1462);
nand U7420 (N_7420,N_3021,N_1564);
and U7421 (N_7421,N_543,N_987);
nand U7422 (N_7422,N_3865,N_1703);
or U7423 (N_7423,N_4719,N_2018);
nor U7424 (N_7424,N_1373,N_795);
nand U7425 (N_7425,N_685,N_1135);
nor U7426 (N_7426,N_2342,N_3647);
nor U7427 (N_7427,N_1212,N_633);
or U7428 (N_7428,N_372,N_2485);
nand U7429 (N_7429,N_3120,N_4730);
nand U7430 (N_7430,N_4634,N_4150);
or U7431 (N_7431,N_204,N_1486);
xor U7432 (N_7432,N_4623,N_1867);
xnor U7433 (N_7433,N_2010,N_3944);
xor U7434 (N_7434,N_23,N_47);
or U7435 (N_7435,N_1844,N_3634);
nor U7436 (N_7436,N_3808,N_1236);
nor U7437 (N_7437,N_2026,N_1673);
and U7438 (N_7438,N_945,N_578);
nor U7439 (N_7439,N_3780,N_4810);
nor U7440 (N_7440,N_3503,N_2753);
xor U7441 (N_7441,N_4039,N_25);
nand U7442 (N_7442,N_2426,N_2055);
nor U7443 (N_7443,N_4692,N_672);
or U7444 (N_7444,N_4069,N_3782);
nor U7445 (N_7445,N_2215,N_3481);
nand U7446 (N_7446,N_4798,N_4473);
nand U7447 (N_7447,N_4779,N_2759);
xor U7448 (N_7448,N_4470,N_2410);
nor U7449 (N_7449,N_2156,N_1539);
nor U7450 (N_7450,N_1018,N_243);
xor U7451 (N_7451,N_2491,N_4803);
and U7452 (N_7452,N_3596,N_879);
nor U7453 (N_7453,N_1977,N_3642);
xor U7454 (N_7454,N_39,N_4631);
or U7455 (N_7455,N_635,N_2404);
xnor U7456 (N_7456,N_97,N_1448);
nand U7457 (N_7457,N_231,N_4059);
nor U7458 (N_7458,N_1027,N_4459);
nor U7459 (N_7459,N_2110,N_485);
xor U7460 (N_7460,N_1122,N_627);
or U7461 (N_7461,N_1157,N_4576);
and U7462 (N_7462,N_1282,N_2475);
nor U7463 (N_7463,N_1562,N_844);
or U7464 (N_7464,N_2504,N_2248);
nor U7465 (N_7465,N_296,N_2870);
nor U7466 (N_7466,N_4425,N_1344);
nand U7467 (N_7467,N_2767,N_1435);
nand U7468 (N_7468,N_539,N_708);
or U7469 (N_7469,N_3257,N_4471);
nand U7470 (N_7470,N_1338,N_2201);
nand U7471 (N_7471,N_4270,N_1367);
and U7472 (N_7472,N_2923,N_2220);
and U7473 (N_7473,N_1798,N_1685);
or U7474 (N_7474,N_3396,N_2380);
nor U7475 (N_7475,N_4663,N_3359);
or U7476 (N_7476,N_1545,N_1938);
and U7477 (N_7477,N_1108,N_4455);
or U7478 (N_7478,N_3200,N_4785);
or U7479 (N_7479,N_4427,N_4699);
xnor U7480 (N_7480,N_4839,N_1521);
nand U7481 (N_7481,N_1920,N_2302);
nand U7482 (N_7482,N_1861,N_4340);
or U7483 (N_7483,N_199,N_1428);
or U7484 (N_7484,N_4010,N_1306);
and U7485 (N_7485,N_4945,N_2835);
or U7486 (N_7486,N_1827,N_81);
and U7487 (N_7487,N_334,N_3014);
xor U7488 (N_7488,N_906,N_355);
nand U7489 (N_7489,N_2392,N_2558);
nand U7490 (N_7490,N_4008,N_401);
or U7491 (N_7491,N_2887,N_2333);
or U7492 (N_7492,N_2757,N_3024);
or U7493 (N_7493,N_587,N_2232);
xnor U7494 (N_7494,N_4230,N_3838);
and U7495 (N_7495,N_3914,N_4733);
or U7496 (N_7496,N_1599,N_3762);
or U7497 (N_7497,N_3507,N_3787);
xnor U7498 (N_7498,N_2960,N_4880);
xor U7499 (N_7499,N_2994,N_3440);
nor U7500 (N_7500,N_3609,N_1828);
nand U7501 (N_7501,N_300,N_3221);
nor U7502 (N_7502,N_306,N_1465);
and U7503 (N_7503,N_1166,N_813);
xor U7504 (N_7504,N_1883,N_686);
nor U7505 (N_7505,N_1133,N_2162);
and U7506 (N_7506,N_3503,N_3009);
nor U7507 (N_7507,N_518,N_1111);
or U7508 (N_7508,N_1236,N_538);
nor U7509 (N_7509,N_87,N_4692);
nor U7510 (N_7510,N_4044,N_2668);
nand U7511 (N_7511,N_2875,N_1826);
xnor U7512 (N_7512,N_4497,N_2330);
and U7513 (N_7513,N_332,N_1161);
xor U7514 (N_7514,N_2383,N_3379);
or U7515 (N_7515,N_1251,N_4914);
xnor U7516 (N_7516,N_87,N_4191);
and U7517 (N_7517,N_1136,N_1559);
xnor U7518 (N_7518,N_4889,N_4528);
and U7519 (N_7519,N_1527,N_3840);
nand U7520 (N_7520,N_499,N_2627);
nand U7521 (N_7521,N_4255,N_1669);
and U7522 (N_7522,N_4005,N_394);
nand U7523 (N_7523,N_2340,N_3007);
nor U7524 (N_7524,N_841,N_4781);
or U7525 (N_7525,N_77,N_2933);
or U7526 (N_7526,N_4132,N_2485);
and U7527 (N_7527,N_1915,N_3173);
and U7528 (N_7528,N_4438,N_4109);
xnor U7529 (N_7529,N_1920,N_2509);
and U7530 (N_7530,N_72,N_916);
nor U7531 (N_7531,N_4336,N_382);
and U7532 (N_7532,N_1288,N_1348);
nand U7533 (N_7533,N_3905,N_2855);
nor U7534 (N_7534,N_3152,N_3430);
nor U7535 (N_7535,N_2087,N_1067);
and U7536 (N_7536,N_2435,N_2552);
nand U7537 (N_7537,N_4095,N_3005);
nor U7538 (N_7538,N_3793,N_1190);
nand U7539 (N_7539,N_398,N_4932);
and U7540 (N_7540,N_4153,N_3372);
xnor U7541 (N_7541,N_568,N_4540);
and U7542 (N_7542,N_2961,N_921);
nand U7543 (N_7543,N_4943,N_3066);
nor U7544 (N_7544,N_1919,N_3643);
nand U7545 (N_7545,N_3897,N_547);
and U7546 (N_7546,N_3818,N_4265);
or U7547 (N_7547,N_4469,N_763);
or U7548 (N_7548,N_3542,N_2355);
nand U7549 (N_7549,N_4731,N_4498);
nand U7550 (N_7550,N_2950,N_2845);
nor U7551 (N_7551,N_704,N_1240);
or U7552 (N_7552,N_2449,N_469);
nor U7553 (N_7553,N_1013,N_2217);
nand U7554 (N_7554,N_3004,N_2837);
nor U7555 (N_7555,N_2424,N_3642);
and U7556 (N_7556,N_1510,N_4161);
xor U7557 (N_7557,N_2099,N_2356);
and U7558 (N_7558,N_2178,N_4200);
xor U7559 (N_7559,N_23,N_3321);
xor U7560 (N_7560,N_2611,N_1407);
or U7561 (N_7561,N_1920,N_3720);
xor U7562 (N_7562,N_3054,N_1975);
nand U7563 (N_7563,N_525,N_2769);
or U7564 (N_7564,N_2061,N_273);
and U7565 (N_7565,N_551,N_811);
or U7566 (N_7566,N_4703,N_1384);
or U7567 (N_7567,N_4472,N_1999);
and U7568 (N_7568,N_1386,N_1136);
nor U7569 (N_7569,N_2501,N_525);
nand U7570 (N_7570,N_2179,N_3604);
nor U7571 (N_7571,N_4289,N_668);
or U7572 (N_7572,N_2435,N_1845);
nor U7573 (N_7573,N_3170,N_1573);
or U7574 (N_7574,N_1270,N_3415);
nor U7575 (N_7575,N_2938,N_4666);
xnor U7576 (N_7576,N_2700,N_760);
xor U7577 (N_7577,N_4497,N_1929);
or U7578 (N_7578,N_3758,N_2617);
nand U7579 (N_7579,N_1984,N_3673);
nand U7580 (N_7580,N_693,N_2866);
and U7581 (N_7581,N_3068,N_4340);
nor U7582 (N_7582,N_4042,N_3919);
nor U7583 (N_7583,N_3016,N_1775);
xor U7584 (N_7584,N_4526,N_1920);
xnor U7585 (N_7585,N_2497,N_1072);
nand U7586 (N_7586,N_76,N_2552);
or U7587 (N_7587,N_4358,N_3870);
nor U7588 (N_7588,N_366,N_1775);
nor U7589 (N_7589,N_1350,N_4401);
or U7590 (N_7590,N_2037,N_3384);
and U7591 (N_7591,N_4177,N_1582);
nand U7592 (N_7592,N_2648,N_4664);
and U7593 (N_7593,N_2764,N_4599);
and U7594 (N_7594,N_1347,N_3014);
nor U7595 (N_7595,N_799,N_1613);
nand U7596 (N_7596,N_4330,N_3850);
and U7597 (N_7597,N_3524,N_2378);
nor U7598 (N_7598,N_1056,N_2385);
nand U7599 (N_7599,N_2340,N_2910);
nand U7600 (N_7600,N_4732,N_1359);
nor U7601 (N_7601,N_109,N_3213);
or U7602 (N_7602,N_3782,N_1689);
or U7603 (N_7603,N_817,N_3823);
and U7604 (N_7604,N_3266,N_1023);
nand U7605 (N_7605,N_330,N_3628);
nor U7606 (N_7606,N_4761,N_3245);
and U7607 (N_7607,N_2800,N_2805);
and U7608 (N_7608,N_4257,N_2877);
and U7609 (N_7609,N_2444,N_3065);
nand U7610 (N_7610,N_3123,N_217);
or U7611 (N_7611,N_2198,N_2922);
nor U7612 (N_7612,N_584,N_1083);
nor U7613 (N_7613,N_58,N_861);
xnor U7614 (N_7614,N_3230,N_3816);
nor U7615 (N_7615,N_4672,N_1254);
nor U7616 (N_7616,N_3050,N_2383);
or U7617 (N_7617,N_1946,N_3525);
nand U7618 (N_7618,N_1003,N_4789);
nand U7619 (N_7619,N_58,N_2814);
nand U7620 (N_7620,N_4293,N_3252);
nand U7621 (N_7621,N_4778,N_3383);
nor U7622 (N_7622,N_735,N_4085);
nand U7623 (N_7623,N_4320,N_4880);
or U7624 (N_7624,N_2086,N_300);
or U7625 (N_7625,N_2283,N_822);
or U7626 (N_7626,N_3811,N_3004);
nor U7627 (N_7627,N_560,N_1329);
or U7628 (N_7628,N_496,N_4388);
nand U7629 (N_7629,N_2289,N_4922);
or U7630 (N_7630,N_1498,N_1779);
nor U7631 (N_7631,N_2879,N_4053);
nor U7632 (N_7632,N_700,N_4872);
and U7633 (N_7633,N_3284,N_212);
or U7634 (N_7634,N_3325,N_2913);
nand U7635 (N_7635,N_3717,N_3644);
nor U7636 (N_7636,N_1137,N_4040);
xor U7637 (N_7637,N_105,N_3524);
nand U7638 (N_7638,N_282,N_4092);
nand U7639 (N_7639,N_1018,N_146);
nand U7640 (N_7640,N_207,N_922);
or U7641 (N_7641,N_3114,N_4157);
nand U7642 (N_7642,N_776,N_1258);
and U7643 (N_7643,N_2178,N_631);
nor U7644 (N_7644,N_3770,N_1379);
xnor U7645 (N_7645,N_480,N_1919);
nand U7646 (N_7646,N_1910,N_114);
and U7647 (N_7647,N_3840,N_38);
or U7648 (N_7648,N_638,N_4332);
or U7649 (N_7649,N_4705,N_2018);
or U7650 (N_7650,N_182,N_3383);
nor U7651 (N_7651,N_79,N_2175);
or U7652 (N_7652,N_97,N_2654);
nor U7653 (N_7653,N_2783,N_1289);
nand U7654 (N_7654,N_1064,N_1509);
or U7655 (N_7655,N_2186,N_535);
and U7656 (N_7656,N_3812,N_2376);
and U7657 (N_7657,N_2606,N_3955);
and U7658 (N_7658,N_2421,N_4426);
nand U7659 (N_7659,N_1804,N_4059);
and U7660 (N_7660,N_4331,N_2309);
nor U7661 (N_7661,N_3613,N_3591);
and U7662 (N_7662,N_279,N_2838);
nor U7663 (N_7663,N_2293,N_1740);
or U7664 (N_7664,N_1535,N_409);
and U7665 (N_7665,N_1613,N_1175);
and U7666 (N_7666,N_2928,N_4204);
nor U7667 (N_7667,N_846,N_612);
nor U7668 (N_7668,N_4170,N_2485);
or U7669 (N_7669,N_2081,N_2876);
nand U7670 (N_7670,N_2464,N_997);
or U7671 (N_7671,N_1023,N_3306);
or U7672 (N_7672,N_1743,N_2956);
or U7673 (N_7673,N_907,N_3327);
nand U7674 (N_7674,N_197,N_3763);
or U7675 (N_7675,N_2954,N_733);
nand U7676 (N_7676,N_4483,N_1617);
nor U7677 (N_7677,N_3304,N_2363);
or U7678 (N_7678,N_1660,N_2125);
nor U7679 (N_7679,N_4419,N_2260);
xor U7680 (N_7680,N_2646,N_210);
or U7681 (N_7681,N_4579,N_420);
and U7682 (N_7682,N_1974,N_960);
or U7683 (N_7683,N_899,N_1037);
nor U7684 (N_7684,N_4273,N_173);
or U7685 (N_7685,N_3811,N_3501);
nand U7686 (N_7686,N_4083,N_4988);
or U7687 (N_7687,N_2194,N_3920);
or U7688 (N_7688,N_766,N_148);
nor U7689 (N_7689,N_117,N_2806);
nand U7690 (N_7690,N_3084,N_2739);
nor U7691 (N_7691,N_1453,N_2471);
nor U7692 (N_7692,N_3559,N_1005);
and U7693 (N_7693,N_4628,N_4685);
nor U7694 (N_7694,N_3859,N_3273);
or U7695 (N_7695,N_2263,N_1330);
or U7696 (N_7696,N_2892,N_518);
nand U7697 (N_7697,N_4042,N_840);
or U7698 (N_7698,N_866,N_1705);
and U7699 (N_7699,N_3636,N_1724);
or U7700 (N_7700,N_2389,N_828);
nand U7701 (N_7701,N_2723,N_1793);
nor U7702 (N_7702,N_2921,N_3305);
nand U7703 (N_7703,N_2865,N_3210);
nand U7704 (N_7704,N_3531,N_2263);
nor U7705 (N_7705,N_3088,N_120);
nor U7706 (N_7706,N_1721,N_669);
nand U7707 (N_7707,N_3763,N_2768);
or U7708 (N_7708,N_750,N_2889);
and U7709 (N_7709,N_697,N_983);
and U7710 (N_7710,N_1984,N_788);
nor U7711 (N_7711,N_2747,N_2640);
nand U7712 (N_7712,N_4128,N_2138);
and U7713 (N_7713,N_1711,N_468);
nor U7714 (N_7714,N_3954,N_4381);
nand U7715 (N_7715,N_3716,N_1748);
or U7716 (N_7716,N_165,N_1833);
xnor U7717 (N_7717,N_42,N_218);
nor U7718 (N_7718,N_3425,N_914);
nand U7719 (N_7719,N_3389,N_2055);
and U7720 (N_7720,N_4385,N_2187);
and U7721 (N_7721,N_4056,N_3039);
nand U7722 (N_7722,N_960,N_4213);
and U7723 (N_7723,N_2278,N_120);
and U7724 (N_7724,N_3495,N_3033);
xnor U7725 (N_7725,N_2885,N_3617);
and U7726 (N_7726,N_2826,N_3649);
and U7727 (N_7727,N_1783,N_2993);
nor U7728 (N_7728,N_4951,N_334);
nor U7729 (N_7729,N_49,N_1950);
or U7730 (N_7730,N_3916,N_4645);
xnor U7731 (N_7731,N_2558,N_4752);
or U7732 (N_7732,N_2597,N_4870);
and U7733 (N_7733,N_4910,N_1461);
nor U7734 (N_7734,N_857,N_26);
and U7735 (N_7735,N_1961,N_3814);
nor U7736 (N_7736,N_3517,N_1398);
xnor U7737 (N_7737,N_4343,N_1617);
nor U7738 (N_7738,N_1026,N_3126);
or U7739 (N_7739,N_3760,N_2561);
nand U7740 (N_7740,N_1992,N_3050);
nand U7741 (N_7741,N_4504,N_1952);
nand U7742 (N_7742,N_3367,N_3448);
or U7743 (N_7743,N_4794,N_956);
and U7744 (N_7744,N_3275,N_3568);
or U7745 (N_7745,N_3478,N_378);
nand U7746 (N_7746,N_3523,N_4316);
nand U7747 (N_7747,N_1794,N_126);
and U7748 (N_7748,N_4697,N_1227);
or U7749 (N_7749,N_3532,N_3129);
nand U7750 (N_7750,N_4894,N_3615);
or U7751 (N_7751,N_2973,N_4450);
nor U7752 (N_7752,N_2551,N_1167);
or U7753 (N_7753,N_837,N_1100);
and U7754 (N_7754,N_4763,N_3465);
or U7755 (N_7755,N_2219,N_1863);
nor U7756 (N_7756,N_1100,N_3822);
or U7757 (N_7757,N_3044,N_1535);
or U7758 (N_7758,N_2885,N_1624);
nand U7759 (N_7759,N_3298,N_2630);
nor U7760 (N_7760,N_3471,N_3427);
nor U7761 (N_7761,N_1282,N_2975);
xor U7762 (N_7762,N_3391,N_4873);
nand U7763 (N_7763,N_2761,N_4793);
nor U7764 (N_7764,N_706,N_226);
and U7765 (N_7765,N_4847,N_2118);
or U7766 (N_7766,N_2501,N_2871);
nor U7767 (N_7767,N_3771,N_3379);
nand U7768 (N_7768,N_1970,N_4600);
or U7769 (N_7769,N_766,N_1007);
nor U7770 (N_7770,N_2421,N_1025);
nand U7771 (N_7771,N_3080,N_4126);
or U7772 (N_7772,N_3162,N_1307);
or U7773 (N_7773,N_3983,N_2214);
or U7774 (N_7774,N_4959,N_1108);
nor U7775 (N_7775,N_4280,N_325);
nor U7776 (N_7776,N_4563,N_2711);
and U7777 (N_7777,N_250,N_4273);
nand U7778 (N_7778,N_612,N_2493);
or U7779 (N_7779,N_2824,N_2151);
and U7780 (N_7780,N_1989,N_4077);
and U7781 (N_7781,N_2975,N_2177);
and U7782 (N_7782,N_4032,N_1095);
and U7783 (N_7783,N_3171,N_1861);
nand U7784 (N_7784,N_2836,N_4027);
nand U7785 (N_7785,N_2350,N_3052);
xor U7786 (N_7786,N_4130,N_800);
or U7787 (N_7787,N_341,N_4468);
or U7788 (N_7788,N_3589,N_35);
or U7789 (N_7789,N_2962,N_1335);
nand U7790 (N_7790,N_4461,N_3676);
and U7791 (N_7791,N_4126,N_380);
and U7792 (N_7792,N_506,N_524);
and U7793 (N_7793,N_3000,N_3390);
nand U7794 (N_7794,N_4691,N_3313);
or U7795 (N_7795,N_4930,N_1023);
or U7796 (N_7796,N_2933,N_4101);
or U7797 (N_7797,N_3324,N_2793);
nor U7798 (N_7798,N_4840,N_1506);
or U7799 (N_7799,N_1538,N_1223);
nor U7800 (N_7800,N_600,N_1986);
or U7801 (N_7801,N_1612,N_1551);
or U7802 (N_7802,N_1436,N_1374);
nand U7803 (N_7803,N_2483,N_3465);
nor U7804 (N_7804,N_2829,N_1262);
or U7805 (N_7805,N_2211,N_3793);
xor U7806 (N_7806,N_139,N_1610);
or U7807 (N_7807,N_3106,N_4617);
xor U7808 (N_7808,N_3317,N_316);
nand U7809 (N_7809,N_2304,N_1132);
or U7810 (N_7810,N_3357,N_3320);
and U7811 (N_7811,N_2523,N_2600);
nor U7812 (N_7812,N_1830,N_4760);
nor U7813 (N_7813,N_2695,N_2759);
nand U7814 (N_7814,N_4545,N_1004);
nor U7815 (N_7815,N_3047,N_947);
or U7816 (N_7816,N_3356,N_44);
nor U7817 (N_7817,N_3197,N_4882);
xnor U7818 (N_7818,N_1721,N_4878);
nand U7819 (N_7819,N_1702,N_4234);
nand U7820 (N_7820,N_4038,N_4514);
nor U7821 (N_7821,N_1383,N_2075);
and U7822 (N_7822,N_4215,N_2324);
and U7823 (N_7823,N_2718,N_732);
xnor U7824 (N_7824,N_1273,N_3037);
xor U7825 (N_7825,N_169,N_1590);
xnor U7826 (N_7826,N_2368,N_4766);
nand U7827 (N_7827,N_4238,N_1986);
nand U7828 (N_7828,N_4594,N_4327);
nand U7829 (N_7829,N_167,N_3772);
xor U7830 (N_7830,N_2449,N_4082);
nand U7831 (N_7831,N_2823,N_2875);
and U7832 (N_7832,N_4232,N_3347);
and U7833 (N_7833,N_4407,N_3032);
nand U7834 (N_7834,N_2634,N_3888);
and U7835 (N_7835,N_1146,N_1211);
or U7836 (N_7836,N_491,N_2864);
or U7837 (N_7837,N_3379,N_1614);
and U7838 (N_7838,N_4544,N_795);
nand U7839 (N_7839,N_2571,N_2534);
nand U7840 (N_7840,N_1513,N_321);
and U7841 (N_7841,N_900,N_906);
xor U7842 (N_7842,N_1593,N_617);
nand U7843 (N_7843,N_4382,N_4098);
or U7844 (N_7844,N_4037,N_4671);
nand U7845 (N_7845,N_4574,N_3862);
nor U7846 (N_7846,N_803,N_793);
nor U7847 (N_7847,N_1215,N_2536);
nor U7848 (N_7848,N_1096,N_4582);
or U7849 (N_7849,N_2552,N_4079);
and U7850 (N_7850,N_4890,N_1228);
or U7851 (N_7851,N_4951,N_4022);
nor U7852 (N_7852,N_1551,N_851);
xnor U7853 (N_7853,N_2378,N_3566);
and U7854 (N_7854,N_413,N_2230);
nand U7855 (N_7855,N_2637,N_589);
nor U7856 (N_7856,N_4403,N_3578);
xnor U7857 (N_7857,N_3299,N_1166);
xnor U7858 (N_7858,N_365,N_256);
and U7859 (N_7859,N_280,N_3793);
nand U7860 (N_7860,N_3853,N_3676);
nand U7861 (N_7861,N_360,N_3631);
or U7862 (N_7862,N_909,N_2060);
or U7863 (N_7863,N_515,N_4551);
xnor U7864 (N_7864,N_4910,N_1197);
or U7865 (N_7865,N_431,N_1097);
xnor U7866 (N_7866,N_1757,N_4734);
nor U7867 (N_7867,N_4051,N_2749);
and U7868 (N_7868,N_4967,N_1976);
nand U7869 (N_7869,N_3994,N_3740);
xor U7870 (N_7870,N_3516,N_2318);
nor U7871 (N_7871,N_4351,N_3523);
nand U7872 (N_7872,N_894,N_2194);
or U7873 (N_7873,N_4923,N_380);
nor U7874 (N_7874,N_2522,N_208);
xor U7875 (N_7875,N_4836,N_3745);
nand U7876 (N_7876,N_3235,N_1075);
nor U7877 (N_7877,N_3990,N_1567);
and U7878 (N_7878,N_3844,N_467);
nand U7879 (N_7879,N_4145,N_4716);
nand U7880 (N_7880,N_3600,N_2544);
or U7881 (N_7881,N_834,N_2931);
and U7882 (N_7882,N_376,N_2036);
nand U7883 (N_7883,N_1775,N_3581);
nor U7884 (N_7884,N_2629,N_4420);
nor U7885 (N_7885,N_1133,N_4527);
nor U7886 (N_7886,N_2366,N_4397);
or U7887 (N_7887,N_4834,N_1942);
or U7888 (N_7888,N_256,N_3447);
nand U7889 (N_7889,N_2074,N_2054);
nor U7890 (N_7890,N_3,N_4351);
nor U7891 (N_7891,N_2696,N_886);
nand U7892 (N_7892,N_4068,N_2405);
nor U7893 (N_7893,N_4511,N_3621);
and U7894 (N_7894,N_2933,N_176);
or U7895 (N_7895,N_2073,N_4356);
or U7896 (N_7896,N_4745,N_2453);
or U7897 (N_7897,N_1096,N_4913);
nand U7898 (N_7898,N_2883,N_342);
or U7899 (N_7899,N_1288,N_3896);
nand U7900 (N_7900,N_1877,N_1816);
nand U7901 (N_7901,N_2697,N_1001);
or U7902 (N_7902,N_2886,N_175);
nand U7903 (N_7903,N_4029,N_2977);
and U7904 (N_7904,N_4137,N_4059);
nand U7905 (N_7905,N_4467,N_3359);
or U7906 (N_7906,N_951,N_1982);
nand U7907 (N_7907,N_2939,N_1346);
nor U7908 (N_7908,N_3232,N_485);
nand U7909 (N_7909,N_4260,N_4183);
nand U7910 (N_7910,N_4004,N_3343);
xor U7911 (N_7911,N_2083,N_281);
or U7912 (N_7912,N_2619,N_2141);
and U7913 (N_7913,N_3222,N_2283);
nand U7914 (N_7914,N_2521,N_95);
nor U7915 (N_7915,N_2575,N_176);
or U7916 (N_7916,N_2922,N_607);
nor U7917 (N_7917,N_3695,N_910);
xnor U7918 (N_7918,N_390,N_276);
nand U7919 (N_7919,N_173,N_3353);
and U7920 (N_7920,N_3997,N_697);
and U7921 (N_7921,N_2909,N_3896);
or U7922 (N_7922,N_2201,N_1596);
nor U7923 (N_7923,N_3039,N_809);
nand U7924 (N_7924,N_3998,N_2609);
xor U7925 (N_7925,N_294,N_3136);
and U7926 (N_7926,N_3944,N_830);
and U7927 (N_7927,N_4653,N_203);
or U7928 (N_7928,N_1543,N_1429);
or U7929 (N_7929,N_2525,N_3790);
nor U7930 (N_7930,N_2850,N_3195);
nor U7931 (N_7931,N_1928,N_4284);
xor U7932 (N_7932,N_2297,N_1637);
or U7933 (N_7933,N_539,N_3571);
or U7934 (N_7934,N_486,N_2462);
nand U7935 (N_7935,N_2729,N_1653);
and U7936 (N_7936,N_2624,N_3834);
xor U7937 (N_7937,N_886,N_1118);
nand U7938 (N_7938,N_199,N_1783);
xnor U7939 (N_7939,N_3946,N_534);
nand U7940 (N_7940,N_3074,N_2262);
nand U7941 (N_7941,N_3987,N_479);
or U7942 (N_7942,N_740,N_1354);
and U7943 (N_7943,N_3204,N_2927);
or U7944 (N_7944,N_943,N_3280);
xnor U7945 (N_7945,N_380,N_974);
or U7946 (N_7946,N_766,N_1093);
or U7947 (N_7947,N_2408,N_3356);
nand U7948 (N_7948,N_531,N_1401);
xor U7949 (N_7949,N_891,N_4419);
or U7950 (N_7950,N_1885,N_1588);
and U7951 (N_7951,N_2928,N_4090);
nand U7952 (N_7952,N_1922,N_4162);
and U7953 (N_7953,N_2436,N_1383);
and U7954 (N_7954,N_147,N_4475);
and U7955 (N_7955,N_4469,N_3547);
xor U7956 (N_7956,N_4885,N_195);
nor U7957 (N_7957,N_4576,N_2900);
nor U7958 (N_7958,N_1356,N_1472);
nand U7959 (N_7959,N_177,N_3189);
nor U7960 (N_7960,N_3730,N_793);
nand U7961 (N_7961,N_4881,N_36);
and U7962 (N_7962,N_744,N_999);
or U7963 (N_7963,N_2673,N_1489);
or U7964 (N_7964,N_709,N_2687);
nand U7965 (N_7965,N_3432,N_676);
nor U7966 (N_7966,N_3592,N_658);
nand U7967 (N_7967,N_3354,N_10);
nand U7968 (N_7968,N_906,N_4666);
or U7969 (N_7969,N_4852,N_4943);
nor U7970 (N_7970,N_1135,N_1148);
nor U7971 (N_7971,N_663,N_3232);
xnor U7972 (N_7972,N_4752,N_3130);
xor U7973 (N_7973,N_4013,N_695);
or U7974 (N_7974,N_1626,N_833);
nand U7975 (N_7975,N_3536,N_1962);
nand U7976 (N_7976,N_2318,N_1828);
and U7977 (N_7977,N_171,N_1442);
nor U7978 (N_7978,N_1986,N_2533);
or U7979 (N_7979,N_38,N_1310);
and U7980 (N_7980,N_3132,N_411);
or U7981 (N_7981,N_4788,N_2417);
and U7982 (N_7982,N_2105,N_3422);
and U7983 (N_7983,N_1198,N_3027);
nor U7984 (N_7984,N_1214,N_1893);
nand U7985 (N_7985,N_3579,N_2413);
nand U7986 (N_7986,N_3972,N_248);
and U7987 (N_7987,N_2364,N_3918);
nor U7988 (N_7988,N_4025,N_4628);
xor U7989 (N_7989,N_1735,N_3039);
and U7990 (N_7990,N_4119,N_381);
or U7991 (N_7991,N_7,N_2760);
or U7992 (N_7992,N_4820,N_3187);
nor U7993 (N_7993,N_3841,N_4078);
nor U7994 (N_7994,N_3596,N_986);
nor U7995 (N_7995,N_716,N_190);
nor U7996 (N_7996,N_4062,N_1022);
nor U7997 (N_7997,N_2413,N_2863);
xor U7998 (N_7998,N_2450,N_2423);
nand U7999 (N_7999,N_4589,N_3839);
or U8000 (N_8000,N_4303,N_98);
nand U8001 (N_8001,N_608,N_4112);
and U8002 (N_8002,N_3510,N_758);
and U8003 (N_8003,N_2824,N_4560);
and U8004 (N_8004,N_2511,N_3936);
nor U8005 (N_8005,N_461,N_2254);
or U8006 (N_8006,N_106,N_1892);
and U8007 (N_8007,N_4681,N_1699);
or U8008 (N_8008,N_3799,N_477);
nand U8009 (N_8009,N_3204,N_2004);
or U8010 (N_8010,N_1709,N_2290);
and U8011 (N_8011,N_1254,N_614);
nand U8012 (N_8012,N_1182,N_166);
or U8013 (N_8013,N_2546,N_2910);
or U8014 (N_8014,N_2433,N_3031);
or U8015 (N_8015,N_4491,N_3128);
xor U8016 (N_8016,N_2380,N_1121);
or U8017 (N_8017,N_2840,N_3003);
and U8018 (N_8018,N_1354,N_1992);
and U8019 (N_8019,N_1397,N_32);
nand U8020 (N_8020,N_1106,N_2112);
xnor U8021 (N_8021,N_1133,N_2660);
nor U8022 (N_8022,N_2924,N_4777);
nor U8023 (N_8023,N_3019,N_3544);
and U8024 (N_8024,N_2487,N_1202);
and U8025 (N_8025,N_2294,N_94);
and U8026 (N_8026,N_1253,N_279);
or U8027 (N_8027,N_824,N_77);
or U8028 (N_8028,N_1410,N_1061);
nand U8029 (N_8029,N_3259,N_601);
and U8030 (N_8030,N_1780,N_613);
nor U8031 (N_8031,N_3397,N_2905);
xnor U8032 (N_8032,N_604,N_1901);
or U8033 (N_8033,N_2542,N_467);
or U8034 (N_8034,N_3631,N_4112);
and U8035 (N_8035,N_4581,N_4542);
and U8036 (N_8036,N_1876,N_1172);
nand U8037 (N_8037,N_1813,N_4209);
nand U8038 (N_8038,N_2268,N_4690);
and U8039 (N_8039,N_3433,N_1298);
or U8040 (N_8040,N_232,N_1143);
and U8041 (N_8041,N_3877,N_4103);
xnor U8042 (N_8042,N_3065,N_4986);
nor U8043 (N_8043,N_4930,N_2468);
or U8044 (N_8044,N_2440,N_2188);
nor U8045 (N_8045,N_3986,N_1000);
nor U8046 (N_8046,N_2245,N_1284);
and U8047 (N_8047,N_2678,N_4180);
or U8048 (N_8048,N_880,N_547);
nor U8049 (N_8049,N_2549,N_936);
nor U8050 (N_8050,N_4611,N_2518);
and U8051 (N_8051,N_4359,N_3030);
nor U8052 (N_8052,N_3059,N_4385);
or U8053 (N_8053,N_3987,N_1702);
nand U8054 (N_8054,N_2259,N_1732);
and U8055 (N_8055,N_4235,N_3758);
nand U8056 (N_8056,N_1158,N_1751);
or U8057 (N_8057,N_1347,N_3483);
nor U8058 (N_8058,N_3145,N_4105);
or U8059 (N_8059,N_2101,N_237);
and U8060 (N_8060,N_435,N_1887);
nor U8061 (N_8061,N_2781,N_961);
and U8062 (N_8062,N_3556,N_3938);
or U8063 (N_8063,N_4486,N_3137);
and U8064 (N_8064,N_600,N_3427);
and U8065 (N_8065,N_1219,N_1214);
nand U8066 (N_8066,N_3870,N_2136);
and U8067 (N_8067,N_1584,N_448);
or U8068 (N_8068,N_2121,N_2783);
nor U8069 (N_8069,N_1593,N_257);
or U8070 (N_8070,N_4285,N_3094);
nand U8071 (N_8071,N_37,N_3631);
and U8072 (N_8072,N_974,N_3267);
nor U8073 (N_8073,N_3998,N_1907);
nand U8074 (N_8074,N_3980,N_3297);
nor U8075 (N_8075,N_2959,N_3513);
and U8076 (N_8076,N_3522,N_2047);
or U8077 (N_8077,N_3267,N_1713);
nor U8078 (N_8078,N_2566,N_3745);
nand U8079 (N_8079,N_4044,N_2230);
nor U8080 (N_8080,N_4003,N_1120);
nand U8081 (N_8081,N_57,N_3040);
and U8082 (N_8082,N_275,N_2315);
xnor U8083 (N_8083,N_150,N_335);
nand U8084 (N_8084,N_1402,N_2061);
xor U8085 (N_8085,N_2788,N_4266);
or U8086 (N_8086,N_3025,N_2119);
nor U8087 (N_8087,N_2049,N_136);
and U8088 (N_8088,N_4168,N_3965);
nor U8089 (N_8089,N_3120,N_1109);
nor U8090 (N_8090,N_2132,N_1281);
nand U8091 (N_8091,N_4856,N_268);
or U8092 (N_8092,N_1681,N_351);
and U8093 (N_8093,N_2672,N_3198);
nand U8094 (N_8094,N_2578,N_1708);
and U8095 (N_8095,N_3415,N_882);
nand U8096 (N_8096,N_510,N_2016);
and U8097 (N_8097,N_1076,N_1328);
or U8098 (N_8098,N_374,N_2224);
or U8099 (N_8099,N_3252,N_235);
nor U8100 (N_8100,N_659,N_1858);
nand U8101 (N_8101,N_4093,N_3881);
xor U8102 (N_8102,N_610,N_2929);
nor U8103 (N_8103,N_4427,N_3938);
and U8104 (N_8104,N_1953,N_3569);
or U8105 (N_8105,N_3810,N_3731);
nand U8106 (N_8106,N_1792,N_2068);
nand U8107 (N_8107,N_1728,N_4863);
and U8108 (N_8108,N_3612,N_3649);
or U8109 (N_8109,N_4797,N_4784);
or U8110 (N_8110,N_3456,N_4059);
and U8111 (N_8111,N_4405,N_3993);
nor U8112 (N_8112,N_4238,N_170);
and U8113 (N_8113,N_4621,N_1309);
and U8114 (N_8114,N_2603,N_1786);
nand U8115 (N_8115,N_3612,N_3838);
or U8116 (N_8116,N_4006,N_366);
nand U8117 (N_8117,N_4545,N_1611);
and U8118 (N_8118,N_351,N_2541);
and U8119 (N_8119,N_2052,N_960);
nand U8120 (N_8120,N_1490,N_4405);
and U8121 (N_8121,N_2424,N_4759);
nor U8122 (N_8122,N_4022,N_909);
nand U8123 (N_8123,N_643,N_1538);
or U8124 (N_8124,N_3511,N_1595);
and U8125 (N_8125,N_624,N_1249);
and U8126 (N_8126,N_4702,N_4635);
nor U8127 (N_8127,N_3620,N_1582);
or U8128 (N_8128,N_569,N_238);
nor U8129 (N_8129,N_2177,N_2598);
or U8130 (N_8130,N_651,N_1429);
nand U8131 (N_8131,N_2361,N_3526);
or U8132 (N_8132,N_1598,N_284);
nor U8133 (N_8133,N_1613,N_4616);
xor U8134 (N_8134,N_4312,N_1676);
and U8135 (N_8135,N_3199,N_1462);
nor U8136 (N_8136,N_1497,N_2218);
nor U8137 (N_8137,N_1801,N_1056);
or U8138 (N_8138,N_4649,N_3189);
and U8139 (N_8139,N_4061,N_2251);
and U8140 (N_8140,N_1903,N_4177);
and U8141 (N_8141,N_1571,N_2117);
xor U8142 (N_8142,N_3488,N_3684);
nand U8143 (N_8143,N_246,N_3345);
or U8144 (N_8144,N_4837,N_3828);
or U8145 (N_8145,N_4265,N_1182);
and U8146 (N_8146,N_1327,N_2189);
nand U8147 (N_8147,N_1496,N_3417);
and U8148 (N_8148,N_3777,N_105);
nand U8149 (N_8149,N_2851,N_244);
nand U8150 (N_8150,N_1252,N_3169);
nor U8151 (N_8151,N_2426,N_2182);
and U8152 (N_8152,N_805,N_2430);
or U8153 (N_8153,N_4987,N_356);
nor U8154 (N_8154,N_3665,N_2006);
nor U8155 (N_8155,N_2704,N_1822);
or U8156 (N_8156,N_4616,N_1212);
xor U8157 (N_8157,N_1136,N_2107);
and U8158 (N_8158,N_368,N_211);
or U8159 (N_8159,N_544,N_506);
xor U8160 (N_8160,N_622,N_1378);
nand U8161 (N_8161,N_1375,N_3669);
nand U8162 (N_8162,N_4717,N_497);
nand U8163 (N_8163,N_4165,N_2598);
nor U8164 (N_8164,N_2585,N_3416);
and U8165 (N_8165,N_3660,N_1477);
or U8166 (N_8166,N_1112,N_2860);
and U8167 (N_8167,N_210,N_4129);
or U8168 (N_8168,N_4773,N_4124);
nand U8169 (N_8169,N_4842,N_3183);
and U8170 (N_8170,N_939,N_172);
and U8171 (N_8171,N_461,N_3992);
nor U8172 (N_8172,N_4972,N_950);
nand U8173 (N_8173,N_3217,N_2105);
nand U8174 (N_8174,N_4505,N_3169);
or U8175 (N_8175,N_112,N_2352);
nor U8176 (N_8176,N_4844,N_1462);
or U8177 (N_8177,N_3488,N_3964);
nand U8178 (N_8178,N_3452,N_1111);
and U8179 (N_8179,N_127,N_2858);
nor U8180 (N_8180,N_2244,N_1436);
or U8181 (N_8181,N_2654,N_4171);
xnor U8182 (N_8182,N_3489,N_3526);
nor U8183 (N_8183,N_4720,N_2648);
or U8184 (N_8184,N_3053,N_4415);
nor U8185 (N_8185,N_13,N_3692);
or U8186 (N_8186,N_596,N_1269);
and U8187 (N_8187,N_2366,N_4852);
xnor U8188 (N_8188,N_2062,N_4167);
and U8189 (N_8189,N_154,N_4049);
nor U8190 (N_8190,N_2596,N_2550);
xor U8191 (N_8191,N_4000,N_1977);
xor U8192 (N_8192,N_2013,N_2908);
nor U8193 (N_8193,N_154,N_2796);
nand U8194 (N_8194,N_2930,N_4090);
or U8195 (N_8195,N_4735,N_3297);
nor U8196 (N_8196,N_869,N_3039);
nor U8197 (N_8197,N_4906,N_4970);
nand U8198 (N_8198,N_2378,N_3197);
nor U8199 (N_8199,N_721,N_1926);
or U8200 (N_8200,N_1350,N_3000);
nand U8201 (N_8201,N_2710,N_1664);
or U8202 (N_8202,N_4192,N_4068);
or U8203 (N_8203,N_2431,N_1742);
nor U8204 (N_8204,N_2204,N_207);
and U8205 (N_8205,N_1893,N_1586);
and U8206 (N_8206,N_2615,N_3916);
and U8207 (N_8207,N_892,N_1585);
and U8208 (N_8208,N_2616,N_2713);
or U8209 (N_8209,N_3928,N_2030);
and U8210 (N_8210,N_3337,N_2752);
and U8211 (N_8211,N_1222,N_1433);
and U8212 (N_8212,N_3418,N_1249);
or U8213 (N_8213,N_2742,N_267);
and U8214 (N_8214,N_1600,N_4223);
and U8215 (N_8215,N_969,N_1527);
nand U8216 (N_8216,N_3259,N_4315);
and U8217 (N_8217,N_4804,N_3650);
and U8218 (N_8218,N_3473,N_1132);
nor U8219 (N_8219,N_1710,N_4385);
nor U8220 (N_8220,N_2248,N_1433);
and U8221 (N_8221,N_2117,N_631);
nor U8222 (N_8222,N_3391,N_2439);
nand U8223 (N_8223,N_816,N_3233);
nor U8224 (N_8224,N_4934,N_1951);
nand U8225 (N_8225,N_1734,N_1832);
nor U8226 (N_8226,N_3293,N_1378);
nor U8227 (N_8227,N_1040,N_898);
or U8228 (N_8228,N_1960,N_4361);
nor U8229 (N_8229,N_4679,N_4369);
nand U8230 (N_8230,N_3430,N_3270);
nor U8231 (N_8231,N_2205,N_4412);
xnor U8232 (N_8232,N_4660,N_871);
or U8233 (N_8233,N_668,N_1722);
nand U8234 (N_8234,N_2038,N_321);
nor U8235 (N_8235,N_1908,N_4344);
nand U8236 (N_8236,N_710,N_3416);
or U8237 (N_8237,N_2037,N_208);
nor U8238 (N_8238,N_4731,N_3712);
nor U8239 (N_8239,N_4529,N_3023);
and U8240 (N_8240,N_4221,N_3137);
and U8241 (N_8241,N_1731,N_3536);
nor U8242 (N_8242,N_2460,N_2456);
nor U8243 (N_8243,N_2108,N_2488);
nor U8244 (N_8244,N_2919,N_1848);
or U8245 (N_8245,N_2919,N_914);
or U8246 (N_8246,N_3825,N_3334);
xnor U8247 (N_8247,N_416,N_2561);
nand U8248 (N_8248,N_1740,N_4292);
or U8249 (N_8249,N_3600,N_1354);
or U8250 (N_8250,N_2396,N_4296);
nor U8251 (N_8251,N_2261,N_1188);
or U8252 (N_8252,N_3623,N_2640);
nor U8253 (N_8253,N_3627,N_4361);
nor U8254 (N_8254,N_2504,N_3174);
or U8255 (N_8255,N_2326,N_2568);
nor U8256 (N_8256,N_1195,N_3022);
and U8257 (N_8257,N_1059,N_2316);
xnor U8258 (N_8258,N_1999,N_3094);
or U8259 (N_8259,N_1159,N_1461);
and U8260 (N_8260,N_1672,N_2998);
and U8261 (N_8261,N_1016,N_1690);
nor U8262 (N_8262,N_204,N_3306);
nand U8263 (N_8263,N_910,N_3703);
nor U8264 (N_8264,N_3157,N_511);
nor U8265 (N_8265,N_1503,N_2648);
and U8266 (N_8266,N_999,N_1346);
or U8267 (N_8267,N_2645,N_3772);
or U8268 (N_8268,N_4139,N_2906);
or U8269 (N_8269,N_1636,N_1847);
or U8270 (N_8270,N_4567,N_3695);
or U8271 (N_8271,N_4274,N_398);
nor U8272 (N_8272,N_87,N_839);
or U8273 (N_8273,N_1584,N_3337);
nor U8274 (N_8274,N_1230,N_1724);
xor U8275 (N_8275,N_2464,N_3173);
or U8276 (N_8276,N_4952,N_3638);
nor U8277 (N_8277,N_1241,N_1220);
nand U8278 (N_8278,N_1226,N_1018);
nor U8279 (N_8279,N_4847,N_742);
or U8280 (N_8280,N_1810,N_3843);
nand U8281 (N_8281,N_3605,N_3190);
nor U8282 (N_8282,N_1660,N_2351);
nor U8283 (N_8283,N_4268,N_751);
nor U8284 (N_8284,N_741,N_4679);
or U8285 (N_8285,N_3464,N_3355);
nor U8286 (N_8286,N_4886,N_2399);
nor U8287 (N_8287,N_2528,N_1985);
nor U8288 (N_8288,N_2647,N_471);
or U8289 (N_8289,N_1309,N_3866);
or U8290 (N_8290,N_3014,N_2702);
or U8291 (N_8291,N_560,N_4608);
or U8292 (N_8292,N_4220,N_4699);
nor U8293 (N_8293,N_521,N_712);
and U8294 (N_8294,N_232,N_2961);
and U8295 (N_8295,N_3976,N_2979);
nor U8296 (N_8296,N_21,N_1445);
nand U8297 (N_8297,N_3459,N_3721);
nand U8298 (N_8298,N_4882,N_655);
nand U8299 (N_8299,N_4145,N_4413);
or U8300 (N_8300,N_1845,N_2570);
nor U8301 (N_8301,N_1574,N_389);
nand U8302 (N_8302,N_2516,N_426);
and U8303 (N_8303,N_4886,N_1161);
or U8304 (N_8304,N_1745,N_1921);
or U8305 (N_8305,N_3939,N_737);
nand U8306 (N_8306,N_209,N_1832);
and U8307 (N_8307,N_1205,N_2413);
or U8308 (N_8308,N_2147,N_1985);
and U8309 (N_8309,N_2648,N_401);
nand U8310 (N_8310,N_2079,N_2864);
and U8311 (N_8311,N_4111,N_2862);
nand U8312 (N_8312,N_2391,N_1428);
or U8313 (N_8313,N_4056,N_4832);
nand U8314 (N_8314,N_913,N_2360);
nor U8315 (N_8315,N_493,N_4967);
and U8316 (N_8316,N_4740,N_2286);
and U8317 (N_8317,N_1113,N_575);
or U8318 (N_8318,N_4632,N_333);
xnor U8319 (N_8319,N_4721,N_3033);
and U8320 (N_8320,N_4102,N_2568);
or U8321 (N_8321,N_943,N_2733);
and U8322 (N_8322,N_2586,N_1907);
and U8323 (N_8323,N_603,N_2999);
and U8324 (N_8324,N_4133,N_3476);
or U8325 (N_8325,N_4279,N_1707);
nand U8326 (N_8326,N_1361,N_2334);
nor U8327 (N_8327,N_1515,N_2763);
or U8328 (N_8328,N_3189,N_4392);
nand U8329 (N_8329,N_166,N_2591);
or U8330 (N_8330,N_4549,N_1404);
or U8331 (N_8331,N_2283,N_832);
and U8332 (N_8332,N_3220,N_84);
and U8333 (N_8333,N_3411,N_2742);
and U8334 (N_8334,N_4464,N_1525);
nor U8335 (N_8335,N_2319,N_4266);
and U8336 (N_8336,N_4919,N_1868);
or U8337 (N_8337,N_877,N_4621);
nor U8338 (N_8338,N_1274,N_3897);
and U8339 (N_8339,N_4865,N_26);
nor U8340 (N_8340,N_2304,N_3104);
or U8341 (N_8341,N_606,N_1626);
or U8342 (N_8342,N_2870,N_4957);
nand U8343 (N_8343,N_3662,N_4141);
or U8344 (N_8344,N_1300,N_349);
nor U8345 (N_8345,N_4874,N_3817);
and U8346 (N_8346,N_3977,N_893);
nand U8347 (N_8347,N_2601,N_1735);
and U8348 (N_8348,N_4433,N_802);
or U8349 (N_8349,N_1026,N_3647);
nor U8350 (N_8350,N_4438,N_3037);
nand U8351 (N_8351,N_28,N_1426);
or U8352 (N_8352,N_2382,N_190);
nor U8353 (N_8353,N_1445,N_1927);
and U8354 (N_8354,N_188,N_2399);
and U8355 (N_8355,N_3953,N_2296);
xnor U8356 (N_8356,N_2654,N_3694);
and U8357 (N_8357,N_4193,N_3332);
xor U8358 (N_8358,N_3083,N_2775);
nand U8359 (N_8359,N_276,N_707);
or U8360 (N_8360,N_3776,N_2084);
nor U8361 (N_8361,N_2263,N_3009);
nand U8362 (N_8362,N_4833,N_747);
and U8363 (N_8363,N_2825,N_4915);
and U8364 (N_8364,N_485,N_1591);
xor U8365 (N_8365,N_1535,N_4631);
nand U8366 (N_8366,N_1856,N_2853);
and U8367 (N_8367,N_357,N_208);
nand U8368 (N_8368,N_251,N_615);
nor U8369 (N_8369,N_2068,N_3704);
and U8370 (N_8370,N_2185,N_2719);
xnor U8371 (N_8371,N_4311,N_1703);
nand U8372 (N_8372,N_2797,N_3455);
nand U8373 (N_8373,N_1997,N_549);
or U8374 (N_8374,N_3225,N_1985);
or U8375 (N_8375,N_2464,N_1548);
xor U8376 (N_8376,N_3530,N_1338);
and U8377 (N_8377,N_2987,N_3426);
and U8378 (N_8378,N_218,N_1749);
or U8379 (N_8379,N_2286,N_3476);
nor U8380 (N_8380,N_2366,N_867);
or U8381 (N_8381,N_344,N_3931);
and U8382 (N_8382,N_3423,N_3032);
or U8383 (N_8383,N_251,N_2672);
or U8384 (N_8384,N_1930,N_4490);
nand U8385 (N_8385,N_847,N_1180);
nor U8386 (N_8386,N_2847,N_4920);
and U8387 (N_8387,N_203,N_4804);
and U8388 (N_8388,N_4925,N_3591);
xor U8389 (N_8389,N_2202,N_4277);
and U8390 (N_8390,N_3603,N_205);
or U8391 (N_8391,N_2302,N_1492);
or U8392 (N_8392,N_2119,N_37);
nand U8393 (N_8393,N_1428,N_449);
or U8394 (N_8394,N_1389,N_263);
and U8395 (N_8395,N_3425,N_20);
and U8396 (N_8396,N_4603,N_3364);
and U8397 (N_8397,N_3154,N_2770);
nand U8398 (N_8398,N_1583,N_4907);
nor U8399 (N_8399,N_2846,N_711);
or U8400 (N_8400,N_2945,N_2002);
or U8401 (N_8401,N_4672,N_4630);
nand U8402 (N_8402,N_2391,N_4558);
nand U8403 (N_8403,N_1573,N_3213);
nor U8404 (N_8404,N_1608,N_3904);
nor U8405 (N_8405,N_545,N_3686);
and U8406 (N_8406,N_42,N_88);
or U8407 (N_8407,N_1547,N_4354);
xor U8408 (N_8408,N_3834,N_1126);
nand U8409 (N_8409,N_1978,N_268);
xor U8410 (N_8410,N_4694,N_3757);
xnor U8411 (N_8411,N_2884,N_3712);
nor U8412 (N_8412,N_1806,N_2660);
or U8413 (N_8413,N_629,N_500);
or U8414 (N_8414,N_3618,N_2730);
nor U8415 (N_8415,N_1068,N_329);
nand U8416 (N_8416,N_4545,N_1704);
xor U8417 (N_8417,N_1305,N_1788);
and U8418 (N_8418,N_4334,N_1350);
nor U8419 (N_8419,N_2323,N_3318);
nor U8420 (N_8420,N_453,N_583);
nor U8421 (N_8421,N_471,N_1834);
and U8422 (N_8422,N_1018,N_4135);
or U8423 (N_8423,N_3620,N_3556);
nor U8424 (N_8424,N_3676,N_1142);
and U8425 (N_8425,N_1152,N_3259);
or U8426 (N_8426,N_914,N_770);
nand U8427 (N_8427,N_3300,N_3984);
and U8428 (N_8428,N_1376,N_175);
nor U8429 (N_8429,N_1929,N_4192);
and U8430 (N_8430,N_4391,N_971);
or U8431 (N_8431,N_2240,N_2861);
nor U8432 (N_8432,N_3878,N_1053);
and U8433 (N_8433,N_2679,N_3744);
or U8434 (N_8434,N_4924,N_2069);
nor U8435 (N_8435,N_4624,N_2375);
nor U8436 (N_8436,N_4975,N_1571);
nand U8437 (N_8437,N_2857,N_1965);
nor U8438 (N_8438,N_2644,N_2280);
nand U8439 (N_8439,N_3237,N_4035);
nor U8440 (N_8440,N_464,N_2216);
or U8441 (N_8441,N_2948,N_1129);
or U8442 (N_8442,N_972,N_1587);
nor U8443 (N_8443,N_4609,N_2100);
or U8444 (N_8444,N_297,N_3484);
and U8445 (N_8445,N_3166,N_2765);
or U8446 (N_8446,N_1334,N_4770);
or U8447 (N_8447,N_2965,N_3044);
and U8448 (N_8448,N_3555,N_147);
nand U8449 (N_8449,N_555,N_1447);
and U8450 (N_8450,N_3663,N_4636);
nand U8451 (N_8451,N_4494,N_1333);
xor U8452 (N_8452,N_1152,N_539);
and U8453 (N_8453,N_3617,N_1425);
or U8454 (N_8454,N_2402,N_3603);
nor U8455 (N_8455,N_2933,N_3134);
and U8456 (N_8456,N_442,N_4030);
nor U8457 (N_8457,N_1485,N_1198);
and U8458 (N_8458,N_3474,N_2350);
nor U8459 (N_8459,N_1808,N_3493);
and U8460 (N_8460,N_408,N_3262);
nor U8461 (N_8461,N_4662,N_1620);
nand U8462 (N_8462,N_92,N_3899);
or U8463 (N_8463,N_3141,N_4574);
or U8464 (N_8464,N_3408,N_2998);
or U8465 (N_8465,N_1371,N_1211);
nand U8466 (N_8466,N_273,N_1913);
and U8467 (N_8467,N_1589,N_3410);
and U8468 (N_8468,N_35,N_4894);
nor U8469 (N_8469,N_2890,N_2755);
nand U8470 (N_8470,N_1736,N_1676);
nor U8471 (N_8471,N_2821,N_3745);
nor U8472 (N_8472,N_4156,N_33);
nand U8473 (N_8473,N_3719,N_631);
xor U8474 (N_8474,N_95,N_2297);
xnor U8475 (N_8475,N_265,N_462);
or U8476 (N_8476,N_1140,N_1263);
xnor U8477 (N_8477,N_3534,N_2031);
nor U8478 (N_8478,N_291,N_2377);
nor U8479 (N_8479,N_2732,N_4729);
and U8480 (N_8480,N_2166,N_4302);
or U8481 (N_8481,N_1528,N_504);
or U8482 (N_8482,N_3711,N_1673);
nor U8483 (N_8483,N_2533,N_1604);
and U8484 (N_8484,N_2963,N_1826);
or U8485 (N_8485,N_3794,N_4322);
nor U8486 (N_8486,N_3315,N_243);
nand U8487 (N_8487,N_27,N_234);
xnor U8488 (N_8488,N_2811,N_4643);
xor U8489 (N_8489,N_469,N_4450);
and U8490 (N_8490,N_104,N_2076);
xor U8491 (N_8491,N_2718,N_2354);
nand U8492 (N_8492,N_1808,N_4821);
or U8493 (N_8493,N_549,N_4744);
nand U8494 (N_8494,N_2074,N_2087);
and U8495 (N_8495,N_16,N_4033);
xor U8496 (N_8496,N_3759,N_1477);
and U8497 (N_8497,N_498,N_4832);
nand U8498 (N_8498,N_3553,N_4601);
nand U8499 (N_8499,N_523,N_4862);
nor U8500 (N_8500,N_2418,N_4697);
and U8501 (N_8501,N_3315,N_150);
nor U8502 (N_8502,N_3863,N_2973);
nand U8503 (N_8503,N_992,N_419);
nor U8504 (N_8504,N_2308,N_2158);
nor U8505 (N_8505,N_2607,N_2179);
or U8506 (N_8506,N_1864,N_1638);
or U8507 (N_8507,N_2291,N_3660);
nor U8508 (N_8508,N_3251,N_3017);
nand U8509 (N_8509,N_4313,N_4471);
xnor U8510 (N_8510,N_2554,N_1853);
xor U8511 (N_8511,N_3935,N_1072);
and U8512 (N_8512,N_490,N_2961);
nand U8513 (N_8513,N_4695,N_3369);
and U8514 (N_8514,N_1067,N_926);
nor U8515 (N_8515,N_2402,N_1783);
and U8516 (N_8516,N_1595,N_2042);
nand U8517 (N_8517,N_268,N_1019);
or U8518 (N_8518,N_4610,N_2156);
nor U8519 (N_8519,N_1283,N_1869);
or U8520 (N_8520,N_1970,N_574);
or U8521 (N_8521,N_2427,N_914);
or U8522 (N_8522,N_3264,N_1251);
nand U8523 (N_8523,N_4802,N_4886);
nor U8524 (N_8524,N_4740,N_2683);
nand U8525 (N_8525,N_19,N_630);
and U8526 (N_8526,N_1143,N_1087);
or U8527 (N_8527,N_2025,N_3186);
nor U8528 (N_8528,N_4127,N_1699);
or U8529 (N_8529,N_3555,N_3776);
nor U8530 (N_8530,N_3502,N_4789);
nor U8531 (N_8531,N_4463,N_1194);
or U8532 (N_8532,N_627,N_1520);
nor U8533 (N_8533,N_3351,N_270);
or U8534 (N_8534,N_329,N_3605);
nor U8535 (N_8535,N_3838,N_3900);
nor U8536 (N_8536,N_4077,N_4559);
nor U8537 (N_8537,N_1345,N_852);
nand U8538 (N_8538,N_1294,N_4677);
and U8539 (N_8539,N_3551,N_1075);
nand U8540 (N_8540,N_77,N_1682);
nand U8541 (N_8541,N_155,N_1026);
and U8542 (N_8542,N_1363,N_4184);
nand U8543 (N_8543,N_876,N_4395);
nor U8544 (N_8544,N_1867,N_3059);
nor U8545 (N_8545,N_1288,N_3240);
nor U8546 (N_8546,N_848,N_3079);
nor U8547 (N_8547,N_4889,N_1707);
xnor U8548 (N_8548,N_3769,N_359);
nor U8549 (N_8549,N_1458,N_2773);
nand U8550 (N_8550,N_4935,N_4096);
nand U8551 (N_8551,N_500,N_3259);
nor U8552 (N_8552,N_3007,N_948);
nor U8553 (N_8553,N_3174,N_4924);
or U8554 (N_8554,N_2840,N_4276);
or U8555 (N_8555,N_3568,N_2118);
or U8556 (N_8556,N_5,N_1632);
nand U8557 (N_8557,N_4574,N_2525);
nand U8558 (N_8558,N_3146,N_274);
nand U8559 (N_8559,N_532,N_2371);
nor U8560 (N_8560,N_1367,N_952);
nand U8561 (N_8561,N_3602,N_3038);
xnor U8562 (N_8562,N_4414,N_1203);
and U8563 (N_8563,N_2349,N_1351);
nand U8564 (N_8564,N_1414,N_1355);
nor U8565 (N_8565,N_2979,N_1784);
and U8566 (N_8566,N_3173,N_3415);
xnor U8567 (N_8567,N_463,N_3924);
or U8568 (N_8568,N_3202,N_4298);
and U8569 (N_8569,N_2056,N_4826);
and U8570 (N_8570,N_1884,N_647);
nor U8571 (N_8571,N_3608,N_4245);
nor U8572 (N_8572,N_3105,N_3503);
and U8573 (N_8573,N_2821,N_2566);
nand U8574 (N_8574,N_1729,N_4868);
nand U8575 (N_8575,N_3700,N_4281);
xnor U8576 (N_8576,N_662,N_3359);
nor U8577 (N_8577,N_4994,N_1806);
xnor U8578 (N_8578,N_2855,N_1965);
nand U8579 (N_8579,N_4196,N_70);
or U8580 (N_8580,N_4479,N_4756);
and U8581 (N_8581,N_3685,N_2569);
and U8582 (N_8582,N_959,N_3740);
xor U8583 (N_8583,N_1035,N_138);
or U8584 (N_8584,N_355,N_1915);
nor U8585 (N_8585,N_792,N_4316);
or U8586 (N_8586,N_3113,N_253);
and U8587 (N_8587,N_409,N_2584);
nand U8588 (N_8588,N_1296,N_1637);
nand U8589 (N_8589,N_4688,N_2370);
xor U8590 (N_8590,N_1262,N_3191);
or U8591 (N_8591,N_2286,N_2784);
nand U8592 (N_8592,N_3875,N_2494);
nand U8593 (N_8593,N_3170,N_3991);
nor U8594 (N_8594,N_2126,N_4542);
nand U8595 (N_8595,N_1264,N_4884);
nand U8596 (N_8596,N_4943,N_3674);
nand U8597 (N_8597,N_3930,N_1883);
or U8598 (N_8598,N_1062,N_821);
xor U8599 (N_8599,N_4857,N_2960);
nor U8600 (N_8600,N_3516,N_1939);
or U8601 (N_8601,N_3449,N_4101);
nand U8602 (N_8602,N_3610,N_2490);
xor U8603 (N_8603,N_2576,N_3165);
nand U8604 (N_8604,N_4880,N_4271);
nand U8605 (N_8605,N_4315,N_1478);
xor U8606 (N_8606,N_2565,N_1439);
or U8607 (N_8607,N_2382,N_2450);
and U8608 (N_8608,N_2444,N_2802);
or U8609 (N_8609,N_2244,N_928);
or U8610 (N_8610,N_4887,N_2127);
nand U8611 (N_8611,N_934,N_648);
nor U8612 (N_8612,N_2004,N_1196);
nor U8613 (N_8613,N_2647,N_2695);
and U8614 (N_8614,N_4122,N_537);
or U8615 (N_8615,N_4672,N_3916);
or U8616 (N_8616,N_1485,N_4902);
nor U8617 (N_8617,N_3315,N_2717);
and U8618 (N_8618,N_606,N_3875);
nand U8619 (N_8619,N_523,N_545);
nand U8620 (N_8620,N_4380,N_4200);
and U8621 (N_8621,N_4188,N_722);
nor U8622 (N_8622,N_3166,N_1030);
and U8623 (N_8623,N_2066,N_1691);
and U8624 (N_8624,N_237,N_4548);
nand U8625 (N_8625,N_3347,N_2917);
nor U8626 (N_8626,N_2709,N_3617);
nand U8627 (N_8627,N_262,N_507);
or U8628 (N_8628,N_4322,N_2888);
nand U8629 (N_8629,N_435,N_2689);
nand U8630 (N_8630,N_2762,N_579);
xor U8631 (N_8631,N_4425,N_2234);
xor U8632 (N_8632,N_4802,N_2037);
or U8633 (N_8633,N_1695,N_1624);
xor U8634 (N_8634,N_4454,N_2922);
nand U8635 (N_8635,N_449,N_1919);
and U8636 (N_8636,N_2987,N_3629);
and U8637 (N_8637,N_4687,N_3141);
or U8638 (N_8638,N_3841,N_256);
xor U8639 (N_8639,N_2620,N_3340);
or U8640 (N_8640,N_832,N_3219);
or U8641 (N_8641,N_3161,N_2243);
nor U8642 (N_8642,N_175,N_2872);
or U8643 (N_8643,N_4040,N_3536);
or U8644 (N_8644,N_4609,N_338);
and U8645 (N_8645,N_2619,N_1182);
or U8646 (N_8646,N_3823,N_4871);
nor U8647 (N_8647,N_3230,N_2577);
nand U8648 (N_8648,N_1222,N_1160);
or U8649 (N_8649,N_2255,N_2135);
and U8650 (N_8650,N_4751,N_1217);
or U8651 (N_8651,N_1721,N_3433);
nor U8652 (N_8652,N_2987,N_4885);
or U8653 (N_8653,N_1803,N_4081);
and U8654 (N_8654,N_1805,N_1246);
nand U8655 (N_8655,N_2753,N_1369);
and U8656 (N_8656,N_495,N_4284);
and U8657 (N_8657,N_403,N_4097);
xor U8658 (N_8658,N_3763,N_3355);
nand U8659 (N_8659,N_2246,N_1657);
nor U8660 (N_8660,N_1404,N_4205);
and U8661 (N_8661,N_626,N_1552);
or U8662 (N_8662,N_4117,N_2985);
or U8663 (N_8663,N_3420,N_3886);
and U8664 (N_8664,N_1071,N_1154);
and U8665 (N_8665,N_4486,N_1874);
nand U8666 (N_8666,N_1780,N_339);
and U8667 (N_8667,N_3121,N_4724);
or U8668 (N_8668,N_4585,N_1915);
or U8669 (N_8669,N_3807,N_3015);
and U8670 (N_8670,N_4196,N_80);
nand U8671 (N_8671,N_4743,N_3972);
xnor U8672 (N_8672,N_371,N_1855);
nor U8673 (N_8673,N_3045,N_2000);
or U8674 (N_8674,N_3253,N_1979);
nor U8675 (N_8675,N_4168,N_519);
nand U8676 (N_8676,N_2954,N_68);
or U8677 (N_8677,N_805,N_3952);
or U8678 (N_8678,N_4810,N_1697);
or U8679 (N_8679,N_1,N_3827);
nand U8680 (N_8680,N_1088,N_4308);
or U8681 (N_8681,N_4009,N_287);
nand U8682 (N_8682,N_870,N_2092);
xor U8683 (N_8683,N_4418,N_2111);
nor U8684 (N_8684,N_783,N_603);
and U8685 (N_8685,N_785,N_3854);
nor U8686 (N_8686,N_345,N_4015);
xnor U8687 (N_8687,N_3026,N_2166);
nor U8688 (N_8688,N_1131,N_4674);
or U8689 (N_8689,N_1085,N_1333);
and U8690 (N_8690,N_3133,N_2757);
xnor U8691 (N_8691,N_1443,N_2956);
nand U8692 (N_8692,N_1567,N_4272);
nor U8693 (N_8693,N_1635,N_1001);
and U8694 (N_8694,N_364,N_2962);
and U8695 (N_8695,N_2898,N_743);
nand U8696 (N_8696,N_3028,N_1654);
nor U8697 (N_8697,N_834,N_2280);
xnor U8698 (N_8698,N_4427,N_3962);
or U8699 (N_8699,N_3343,N_1309);
nor U8700 (N_8700,N_2035,N_959);
and U8701 (N_8701,N_1748,N_1668);
or U8702 (N_8702,N_1635,N_2504);
nand U8703 (N_8703,N_1171,N_3645);
and U8704 (N_8704,N_4102,N_4581);
nand U8705 (N_8705,N_694,N_3262);
or U8706 (N_8706,N_842,N_3804);
or U8707 (N_8707,N_234,N_2099);
xnor U8708 (N_8708,N_392,N_187);
nor U8709 (N_8709,N_490,N_3063);
nor U8710 (N_8710,N_134,N_2747);
xnor U8711 (N_8711,N_1485,N_1982);
and U8712 (N_8712,N_1096,N_4307);
xor U8713 (N_8713,N_3489,N_2117);
or U8714 (N_8714,N_4238,N_4078);
or U8715 (N_8715,N_1763,N_3730);
or U8716 (N_8716,N_4816,N_936);
or U8717 (N_8717,N_2970,N_2801);
or U8718 (N_8718,N_297,N_472);
and U8719 (N_8719,N_2524,N_3933);
or U8720 (N_8720,N_603,N_3672);
nand U8721 (N_8721,N_1488,N_3095);
nand U8722 (N_8722,N_464,N_1582);
nor U8723 (N_8723,N_1626,N_167);
nand U8724 (N_8724,N_1860,N_4663);
or U8725 (N_8725,N_3626,N_249);
or U8726 (N_8726,N_808,N_455);
or U8727 (N_8727,N_3394,N_2997);
and U8728 (N_8728,N_600,N_2222);
nand U8729 (N_8729,N_852,N_3756);
or U8730 (N_8730,N_2286,N_4379);
nor U8731 (N_8731,N_1053,N_1045);
and U8732 (N_8732,N_3283,N_2226);
and U8733 (N_8733,N_881,N_4514);
nand U8734 (N_8734,N_365,N_3109);
and U8735 (N_8735,N_3070,N_2705);
or U8736 (N_8736,N_4437,N_394);
nand U8737 (N_8737,N_4327,N_2574);
and U8738 (N_8738,N_2721,N_403);
or U8739 (N_8739,N_4227,N_2138);
xor U8740 (N_8740,N_3836,N_2653);
xnor U8741 (N_8741,N_2843,N_1024);
nand U8742 (N_8742,N_1679,N_4966);
and U8743 (N_8743,N_1362,N_4214);
and U8744 (N_8744,N_1665,N_4743);
and U8745 (N_8745,N_988,N_3505);
xor U8746 (N_8746,N_4624,N_2710);
or U8747 (N_8747,N_1393,N_3312);
nand U8748 (N_8748,N_1956,N_1178);
and U8749 (N_8749,N_3086,N_4114);
nor U8750 (N_8750,N_2210,N_2346);
or U8751 (N_8751,N_3069,N_1591);
nand U8752 (N_8752,N_748,N_2595);
nand U8753 (N_8753,N_3870,N_4205);
or U8754 (N_8754,N_4731,N_4162);
nor U8755 (N_8755,N_3483,N_2906);
xnor U8756 (N_8756,N_4860,N_2451);
or U8757 (N_8757,N_1762,N_4830);
and U8758 (N_8758,N_664,N_3244);
nor U8759 (N_8759,N_3715,N_1716);
or U8760 (N_8760,N_481,N_4342);
or U8761 (N_8761,N_1417,N_2781);
or U8762 (N_8762,N_3107,N_2204);
and U8763 (N_8763,N_856,N_629);
or U8764 (N_8764,N_2873,N_1948);
and U8765 (N_8765,N_1047,N_1259);
nor U8766 (N_8766,N_4150,N_1591);
nand U8767 (N_8767,N_2339,N_4257);
or U8768 (N_8768,N_3872,N_747);
nor U8769 (N_8769,N_595,N_1203);
nor U8770 (N_8770,N_1814,N_970);
nand U8771 (N_8771,N_601,N_1848);
or U8772 (N_8772,N_2137,N_3165);
xor U8773 (N_8773,N_2160,N_4126);
nand U8774 (N_8774,N_173,N_313);
nand U8775 (N_8775,N_1929,N_3835);
nor U8776 (N_8776,N_3518,N_818);
nor U8777 (N_8777,N_1355,N_3250);
and U8778 (N_8778,N_1162,N_908);
and U8779 (N_8779,N_1953,N_3067);
nor U8780 (N_8780,N_1676,N_196);
nor U8781 (N_8781,N_2777,N_3611);
nand U8782 (N_8782,N_4604,N_1676);
nor U8783 (N_8783,N_3537,N_9);
nand U8784 (N_8784,N_716,N_3884);
nand U8785 (N_8785,N_3765,N_282);
nor U8786 (N_8786,N_3150,N_2003);
and U8787 (N_8787,N_3977,N_616);
xnor U8788 (N_8788,N_2855,N_2561);
nor U8789 (N_8789,N_1386,N_1154);
or U8790 (N_8790,N_3089,N_3969);
xor U8791 (N_8791,N_2699,N_2706);
or U8792 (N_8792,N_4734,N_2004);
nand U8793 (N_8793,N_1929,N_851);
xnor U8794 (N_8794,N_4987,N_4605);
and U8795 (N_8795,N_277,N_1286);
xnor U8796 (N_8796,N_2734,N_4976);
xor U8797 (N_8797,N_3658,N_1471);
nor U8798 (N_8798,N_1629,N_4235);
and U8799 (N_8799,N_1336,N_4013);
nand U8800 (N_8800,N_1202,N_4589);
and U8801 (N_8801,N_3529,N_4174);
or U8802 (N_8802,N_443,N_4316);
and U8803 (N_8803,N_431,N_577);
or U8804 (N_8804,N_2928,N_261);
xor U8805 (N_8805,N_96,N_607);
and U8806 (N_8806,N_2637,N_4937);
nor U8807 (N_8807,N_2850,N_2251);
nand U8808 (N_8808,N_4611,N_297);
nand U8809 (N_8809,N_1550,N_3442);
xor U8810 (N_8810,N_4135,N_3066);
and U8811 (N_8811,N_3611,N_3786);
nor U8812 (N_8812,N_4791,N_4571);
or U8813 (N_8813,N_3400,N_2270);
and U8814 (N_8814,N_3727,N_802);
and U8815 (N_8815,N_4214,N_1690);
nand U8816 (N_8816,N_4306,N_2350);
or U8817 (N_8817,N_4834,N_2547);
nor U8818 (N_8818,N_105,N_1222);
or U8819 (N_8819,N_2724,N_3836);
xnor U8820 (N_8820,N_434,N_3747);
xnor U8821 (N_8821,N_2355,N_709);
nand U8822 (N_8822,N_1186,N_22);
nor U8823 (N_8823,N_1612,N_1078);
nand U8824 (N_8824,N_3970,N_4734);
xnor U8825 (N_8825,N_3987,N_4458);
nor U8826 (N_8826,N_1552,N_1640);
or U8827 (N_8827,N_3066,N_1214);
xnor U8828 (N_8828,N_226,N_55);
and U8829 (N_8829,N_1677,N_2088);
xor U8830 (N_8830,N_609,N_4636);
nand U8831 (N_8831,N_4710,N_4688);
or U8832 (N_8832,N_4126,N_3180);
nor U8833 (N_8833,N_1059,N_4746);
and U8834 (N_8834,N_1701,N_3738);
and U8835 (N_8835,N_596,N_3963);
nor U8836 (N_8836,N_797,N_4079);
and U8837 (N_8837,N_3625,N_3693);
or U8838 (N_8838,N_3007,N_1831);
nor U8839 (N_8839,N_3986,N_3418);
and U8840 (N_8840,N_1758,N_2464);
nand U8841 (N_8841,N_4424,N_2879);
xnor U8842 (N_8842,N_468,N_253);
and U8843 (N_8843,N_717,N_3879);
nand U8844 (N_8844,N_188,N_4656);
nor U8845 (N_8845,N_4653,N_3695);
xor U8846 (N_8846,N_2627,N_680);
or U8847 (N_8847,N_1346,N_3740);
nand U8848 (N_8848,N_4285,N_1759);
and U8849 (N_8849,N_3197,N_678);
nor U8850 (N_8850,N_187,N_4875);
nand U8851 (N_8851,N_4224,N_2844);
or U8852 (N_8852,N_1997,N_4458);
nor U8853 (N_8853,N_10,N_1255);
and U8854 (N_8854,N_2828,N_3915);
nor U8855 (N_8855,N_3946,N_2363);
nand U8856 (N_8856,N_3992,N_3347);
and U8857 (N_8857,N_3868,N_276);
or U8858 (N_8858,N_3035,N_2772);
and U8859 (N_8859,N_3105,N_4821);
and U8860 (N_8860,N_1681,N_2542);
nor U8861 (N_8861,N_2517,N_420);
and U8862 (N_8862,N_4952,N_36);
or U8863 (N_8863,N_1691,N_190);
and U8864 (N_8864,N_2625,N_2929);
or U8865 (N_8865,N_4673,N_4142);
and U8866 (N_8866,N_4017,N_1384);
and U8867 (N_8867,N_1974,N_4164);
nand U8868 (N_8868,N_2929,N_322);
xnor U8869 (N_8869,N_2098,N_3018);
nor U8870 (N_8870,N_1900,N_3111);
nor U8871 (N_8871,N_3460,N_2197);
and U8872 (N_8872,N_1825,N_1498);
and U8873 (N_8873,N_40,N_2367);
nor U8874 (N_8874,N_1991,N_2339);
nand U8875 (N_8875,N_8,N_4587);
nand U8876 (N_8876,N_3825,N_957);
and U8877 (N_8877,N_2313,N_993);
nor U8878 (N_8878,N_3243,N_4415);
and U8879 (N_8879,N_688,N_4058);
xnor U8880 (N_8880,N_4962,N_281);
nor U8881 (N_8881,N_2464,N_1452);
or U8882 (N_8882,N_1611,N_1466);
nand U8883 (N_8883,N_2037,N_4971);
and U8884 (N_8884,N_3345,N_3228);
nor U8885 (N_8885,N_2509,N_482);
or U8886 (N_8886,N_3230,N_3934);
nand U8887 (N_8887,N_1567,N_4982);
and U8888 (N_8888,N_310,N_323);
xnor U8889 (N_8889,N_2301,N_1778);
nor U8890 (N_8890,N_3824,N_1270);
or U8891 (N_8891,N_3884,N_2763);
nand U8892 (N_8892,N_2634,N_4793);
or U8893 (N_8893,N_210,N_3070);
nor U8894 (N_8894,N_2419,N_3362);
nand U8895 (N_8895,N_3815,N_4086);
nand U8896 (N_8896,N_2508,N_4994);
and U8897 (N_8897,N_1092,N_1872);
and U8898 (N_8898,N_4574,N_1666);
nand U8899 (N_8899,N_480,N_4591);
nand U8900 (N_8900,N_1465,N_1534);
or U8901 (N_8901,N_2156,N_3586);
nand U8902 (N_8902,N_3987,N_1665);
or U8903 (N_8903,N_1646,N_4161);
nand U8904 (N_8904,N_2567,N_535);
nor U8905 (N_8905,N_3552,N_2466);
nand U8906 (N_8906,N_2616,N_1613);
and U8907 (N_8907,N_1257,N_1379);
and U8908 (N_8908,N_1493,N_4109);
or U8909 (N_8909,N_665,N_2479);
nor U8910 (N_8910,N_2546,N_3956);
nor U8911 (N_8911,N_698,N_79);
or U8912 (N_8912,N_3155,N_1549);
nor U8913 (N_8913,N_405,N_4446);
xor U8914 (N_8914,N_1718,N_2569);
nand U8915 (N_8915,N_657,N_4022);
or U8916 (N_8916,N_3774,N_247);
nand U8917 (N_8917,N_1571,N_4519);
nor U8918 (N_8918,N_109,N_2753);
xor U8919 (N_8919,N_3901,N_1833);
and U8920 (N_8920,N_2137,N_4853);
nand U8921 (N_8921,N_963,N_4772);
nor U8922 (N_8922,N_4007,N_257);
or U8923 (N_8923,N_4072,N_913);
and U8924 (N_8924,N_2078,N_2892);
nor U8925 (N_8925,N_496,N_2810);
or U8926 (N_8926,N_2875,N_1972);
or U8927 (N_8927,N_1257,N_2797);
or U8928 (N_8928,N_3131,N_2070);
or U8929 (N_8929,N_3160,N_677);
nand U8930 (N_8930,N_3179,N_4197);
or U8931 (N_8931,N_774,N_4125);
and U8932 (N_8932,N_502,N_4861);
or U8933 (N_8933,N_4537,N_4137);
nor U8934 (N_8934,N_866,N_3660);
nand U8935 (N_8935,N_2902,N_1262);
nor U8936 (N_8936,N_3133,N_3685);
or U8937 (N_8937,N_1883,N_825);
nor U8938 (N_8938,N_1323,N_4222);
or U8939 (N_8939,N_4495,N_3021);
nand U8940 (N_8940,N_1708,N_488);
nor U8941 (N_8941,N_528,N_1759);
and U8942 (N_8942,N_288,N_1440);
or U8943 (N_8943,N_4113,N_2874);
xnor U8944 (N_8944,N_2604,N_4587);
or U8945 (N_8945,N_3733,N_601);
nor U8946 (N_8946,N_4572,N_2886);
xor U8947 (N_8947,N_3263,N_1686);
nand U8948 (N_8948,N_4716,N_2421);
and U8949 (N_8949,N_2420,N_2685);
and U8950 (N_8950,N_4042,N_4649);
and U8951 (N_8951,N_1812,N_478);
or U8952 (N_8952,N_3466,N_1848);
xnor U8953 (N_8953,N_2270,N_2478);
and U8954 (N_8954,N_3361,N_4621);
and U8955 (N_8955,N_3895,N_1229);
nor U8956 (N_8956,N_945,N_1021);
nor U8957 (N_8957,N_810,N_2645);
nor U8958 (N_8958,N_560,N_4998);
and U8959 (N_8959,N_3703,N_4014);
nor U8960 (N_8960,N_4025,N_783);
or U8961 (N_8961,N_1609,N_250);
and U8962 (N_8962,N_2036,N_4361);
and U8963 (N_8963,N_19,N_733);
nor U8964 (N_8964,N_674,N_3957);
and U8965 (N_8965,N_393,N_1766);
nand U8966 (N_8966,N_1564,N_3879);
nand U8967 (N_8967,N_3072,N_3464);
nand U8968 (N_8968,N_1115,N_1813);
and U8969 (N_8969,N_1504,N_3200);
or U8970 (N_8970,N_736,N_4204);
or U8971 (N_8971,N_4796,N_4871);
xor U8972 (N_8972,N_4038,N_3267);
nand U8973 (N_8973,N_843,N_1153);
xor U8974 (N_8974,N_4501,N_2338);
and U8975 (N_8975,N_3218,N_1238);
xnor U8976 (N_8976,N_1272,N_4539);
nor U8977 (N_8977,N_2659,N_318);
nor U8978 (N_8978,N_3904,N_557);
and U8979 (N_8979,N_822,N_1231);
or U8980 (N_8980,N_2567,N_3465);
nand U8981 (N_8981,N_4951,N_4469);
nand U8982 (N_8982,N_3055,N_2331);
or U8983 (N_8983,N_724,N_1194);
nand U8984 (N_8984,N_1081,N_39);
xor U8985 (N_8985,N_80,N_1395);
nand U8986 (N_8986,N_1721,N_2344);
nor U8987 (N_8987,N_1142,N_726);
and U8988 (N_8988,N_2131,N_4011);
xor U8989 (N_8989,N_1866,N_1776);
or U8990 (N_8990,N_2446,N_665);
xnor U8991 (N_8991,N_985,N_3648);
or U8992 (N_8992,N_729,N_2994);
nand U8993 (N_8993,N_298,N_4828);
or U8994 (N_8994,N_2534,N_3277);
and U8995 (N_8995,N_4330,N_2371);
nand U8996 (N_8996,N_4688,N_1884);
nor U8997 (N_8997,N_4188,N_1078);
and U8998 (N_8998,N_3601,N_2666);
or U8999 (N_8999,N_1380,N_1073);
or U9000 (N_9000,N_1701,N_2892);
nand U9001 (N_9001,N_3011,N_1237);
or U9002 (N_9002,N_2782,N_2301);
xor U9003 (N_9003,N_1127,N_372);
and U9004 (N_9004,N_3538,N_356);
or U9005 (N_9005,N_4701,N_2429);
nand U9006 (N_9006,N_2028,N_3517);
and U9007 (N_9007,N_3895,N_3170);
xor U9008 (N_9008,N_2774,N_2586);
nand U9009 (N_9009,N_4810,N_62);
and U9010 (N_9010,N_4933,N_1502);
nor U9011 (N_9011,N_1089,N_4377);
and U9012 (N_9012,N_3875,N_439);
nor U9013 (N_9013,N_1869,N_2211);
or U9014 (N_9014,N_2954,N_2915);
and U9015 (N_9015,N_3334,N_4110);
nand U9016 (N_9016,N_4600,N_963);
xor U9017 (N_9017,N_1553,N_2735);
and U9018 (N_9018,N_3001,N_2693);
nand U9019 (N_9019,N_1609,N_2569);
nor U9020 (N_9020,N_2404,N_4995);
nor U9021 (N_9021,N_4454,N_4650);
nand U9022 (N_9022,N_2639,N_2567);
nand U9023 (N_9023,N_1656,N_4757);
or U9024 (N_9024,N_2513,N_380);
nor U9025 (N_9025,N_4892,N_4317);
and U9026 (N_9026,N_2083,N_1595);
nor U9027 (N_9027,N_4373,N_2327);
nor U9028 (N_9028,N_4298,N_4424);
or U9029 (N_9029,N_1485,N_3987);
nand U9030 (N_9030,N_4571,N_3715);
nand U9031 (N_9031,N_3435,N_535);
or U9032 (N_9032,N_399,N_657);
nor U9033 (N_9033,N_2960,N_4876);
or U9034 (N_9034,N_4624,N_1281);
or U9035 (N_9035,N_191,N_540);
and U9036 (N_9036,N_3219,N_3509);
and U9037 (N_9037,N_1540,N_1738);
or U9038 (N_9038,N_3989,N_1025);
xnor U9039 (N_9039,N_3204,N_1300);
or U9040 (N_9040,N_3543,N_2678);
nor U9041 (N_9041,N_2637,N_3161);
nor U9042 (N_9042,N_2350,N_1984);
nor U9043 (N_9043,N_4391,N_2330);
and U9044 (N_9044,N_481,N_476);
and U9045 (N_9045,N_4404,N_1754);
nor U9046 (N_9046,N_4652,N_4388);
nand U9047 (N_9047,N_1927,N_4708);
and U9048 (N_9048,N_131,N_3280);
nor U9049 (N_9049,N_3974,N_2645);
and U9050 (N_9050,N_4443,N_1812);
nand U9051 (N_9051,N_4913,N_1789);
or U9052 (N_9052,N_4361,N_1478);
and U9053 (N_9053,N_4748,N_2833);
nand U9054 (N_9054,N_1759,N_1695);
and U9055 (N_9055,N_4662,N_3592);
xnor U9056 (N_9056,N_2810,N_1559);
nand U9057 (N_9057,N_1470,N_3203);
or U9058 (N_9058,N_908,N_1135);
and U9059 (N_9059,N_1505,N_886);
or U9060 (N_9060,N_2294,N_257);
xnor U9061 (N_9061,N_4607,N_1789);
or U9062 (N_9062,N_4689,N_914);
nand U9063 (N_9063,N_3629,N_4130);
nor U9064 (N_9064,N_4459,N_1558);
and U9065 (N_9065,N_4343,N_1293);
xor U9066 (N_9066,N_1262,N_239);
or U9067 (N_9067,N_1854,N_1235);
and U9068 (N_9068,N_823,N_3667);
nor U9069 (N_9069,N_353,N_4913);
nor U9070 (N_9070,N_640,N_276);
nand U9071 (N_9071,N_1703,N_3632);
or U9072 (N_9072,N_4036,N_1626);
and U9073 (N_9073,N_3258,N_920);
and U9074 (N_9074,N_2405,N_3767);
nor U9075 (N_9075,N_3023,N_1819);
nand U9076 (N_9076,N_4212,N_348);
or U9077 (N_9077,N_54,N_2157);
and U9078 (N_9078,N_2983,N_1398);
xnor U9079 (N_9079,N_689,N_2934);
nor U9080 (N_9080,N_589,N_393);
xor U9081 (N_9081,N_4453,N_657);
and U9082 (N_9082,N_3513,N_1741);
nand U9083 (N_9083,N_1918,N_3768);
nor U9084 (N_9084,N_2746,N_2431);
xor U9085 (N_9085,N_3399,N_1399);
xor U9086 (N_9086,N_1453,N_3957);
nand U9087 (N_9087,N_116,N_1980);
nor U9088 (N_9088,N_4731,N_4205);
or U9089 (N_9089,N_1330,N_2805);
or U9090 (N_9090,N_2791,N_2812);
nand U9091 (N_9091,N_88,N_4759);
nor U9092 (N_9092,N_3645,N_3087);
or U9093 (N_9093,N_866,N_4897);
nand U9094 (N_9094,N_2862,N_3400);
nand U9095 (N_9095,N_1654,N_407);
xor U9096 (N_9096,N_4694,N_1667);
nand U9097 (N_9097,N_3561,N_96);
nor U9098 (N_9098,N_3773,N_3815);
nor U9099 (N_9099,N_3409,N_1056);
nor U9100 (N_9100,N_3854,N_1823);
xor U9101 (N_9101,N_4832,N_4713);
or U9102 (N_9102,N_3157,N_2259);
nor U9103 (N_9103,N_1697,N_2282);
and U9104 (N_9104,N_654,N_4178);
and U9105 (N_9105,N_2146,N_4778);
or U9106 (N_9106,N_2327,N_29);
and U9107 (N_9107,N_4108,N_3082);
and U9108 (N_9108,N_1525,N_547);
nand U9109 (N_9109,N_3405,N_3784);
nand U9110 (N_9110,N_2003,N_3898);
and U9111 (N_9111,N_2757,N_3137);
or U9112 (N_9112,N_4892,N_3577);
or U9113 (N_9113,N_2491,N_2316);
nor U9114 (N_9114,N_556,N_1828);
nand U9115 (N_9115,N_3699,N_1173);
or U9116 (N_9116,N_316,N_2775);
nor U9117 (N_9117,N_4686,N_1825);
and U9118 (N_9118,N_4292,N_653);
and U9119 (N_9119,N_2678,N_1020);
and U9120 (N_9120,N_1218,N_4643);
or U9121 (N_9121,N_4278,N_4413);
nand U9122 (N_9122,N_4953,N_4289);
nor U9123 (N_9123,N_545,N_4376);
xnor U9124 (N_9124,N_2969,N_4472);
or U9125 (N_9125,N_1430,N_3528);
and U9126 (N_9126,N_4431,N_553);
nor U9127 (N_9127,N_267,N_3577);
and U9128 (N_9128,N_3411,N_615);
xnor U9129 (N_9129,N_180,N_716);
or U9130 (N_9130,N_4434,N_1839);
nand U9131 (N_9131,N_273,N_1152);
and U9132 (N_9132,N_3137,N_84);
and U9133 (N_9133,N_1852,N_4488);
nand U9134 (N_9134,N_208,N_2951);
xnor U9135 (N_9135,N_3405,N_509);
or U9136 (N_9136,N_4955,N_903);
nand U9137 (N_9137,N_2682,N_580);
or U9138 (N_9138,N_252,N_4726);
or U9139 (N_9139,N_539,N_4642);
nand U9140 (N_9140,N_1551,N_4176);
nor U9141 (N_9141,N_1327,N_3732);
and U9142 (N_9142,N_1278,N_958);
or U9143 (N_9143,N_2329,N_777);
or U9144 (N_9144,N_2877,N_4026);
nand U9145 (N_9145,N_402,N_3929);
nor U9146 (N_9146,N_4108,N_865);
nor U9147 (N_9147,N_2090,N_2246);
xnor U9148 (N_9148,N_550,N_284);
and U9149 (N_9149,N_1552,N_805);
xor U9150 (N_9150,N_3864,N_4360);
and U9151 (N_9151,N_3123,N_4913);
and U9152 (N_9152,N_4556,N_295);
or U9153 (N_9153,N_3020,N_3027);
nor U9154 (N_9154,N_968,N_1669);
nand U9155 (N_9155,N_2908,N_4338);
or U9156 (N_9156,N_2147,N_4717);
xnor U9157 (N_9157,N_2903,N_4400);
nand U9158 (N_9158,N_3719,N_4785);
or U9159 (N_9159,N_588,N_1521);
nor U9160 (N_9160,N_1185,N_3734);
nor U9161 (N_9161,N_3438,N_431);
xor U9162 (N_9162,N_895,N_4950);
xnor U9163 (N_9163,N_496,N_3637);
or U9164 (N_9164,N_3516,N_1142);
nand U9165 (N_9165,N_4968,N_2468);
nor U9166 (N_9166,N_2372,N_1446);
nor U9167 (N_9167,N_3755,N_4528);
nand U9168 (N_9168,N_2362,N_1257);
nand U9169 (N_9169,N_827,N_4450);
nor U9170 (N_9170,N_3078,N_99);
nor U9171 (N_9171,N_751,N_745);
and U9172 (N_9172,N_731,N_4519);
and U9173 (N_9173,N_856,N_1701);
nor U9174 (N_9174,N_1710,N_3468);
and U9175 (N_9175,N_2816,N_3999);
nor U9176 (N_9176,N_1767,N_4428);
and U9177 (N_9177,N_4939,N_3106);
nand U9178 (N_9178,N_4394,N_2544);
nand U9179 (N_9179,N_4217,N_788);
xor U9180 (N_9180,N_220,N_959);
xnor U9181 (N_9181,N_1620,N_3896);
and U9182 (N_9182,N_3495,N_912);
and U9183 (N_9183,N_4967,N_2717);
or U9184 (N_9184,N_1611,N_2948);
nor U9185 (N_9185,N_316,N_3329);
and U9186 (N_9186,N_2764,N_2248);
nor U9187 (N_9187,N_4808,N_1092);
and U9188 (N_9188,N_1464,N_3419);
or U9189 (N_9189,N_3707,N_1853);
xnor U9190 (N_9190,N_4252,N_4166);
nor U9191 (N_9191,N_2649,N_110);
nand U9192 (N_9192,N_721,N_3401);
nand U9193 (N_9193,N_1029,N_2494);
xor U9194 (N_9194,N_3925,N_3160);
and U9195 (N_9195,N_612,N_787);
nor U9196 (N_9196,N_3499,N_2686);
or U9197 (N_9197,N_4510,N_2499);
or U9198 (N_9198,N_1594,N_2003);
nand U9199 (N_9199,N_242,N_1329);
and U9200 (N_9200,N_3415,N_970);
and U9201 (N_9201,N_184,N_2605);
and U9202 (N_9202,N_3927,N_402);
nor U9203 (N_9203,N_2811,N_3663);
nand U9204 (N_9204,N_407,N_1066);
or U9205 (N_9205,N_2199,N_3567);
nand U9206 (N_9206,N_483,N_463);
and U9207 (N_9207,N_2110,N_2398);
nor U9208 (N_9208,N_926,N_3503);
xnor U9209 (N_9209,N_3048,N_1392);
nand U9210 (N_9210,N_1680,N_678);
nor U9211 (N_9211,N_208,N_1753);
nor U9212 (N_9212,N_3387,N_4707);
or U9213 (N_9213,N_2290,N_3965);
and U9214 (N_9214,N_2822,N_4214);
and U9215 (N_9215,N_1124,N_4615);
nand U9216 (N_9216,N_1767,N_4851);
nor U9217 (N_9217,N_2445,N_1442);
nor U9218 (N_9218,N_2459,N_1147);
nor U9219 (N_9219,N_4928,N_4522);
nor U9220 (N_9220,N_3207,N_415);
and U9221 (N_9221,N_3546,N_4418);
and U9222 (N_9222,N_4685,N_4568);
nor U9223 (N_9223,N_2467,N_2772);
nor U9224 (N_9224,N_973,N_82);
nand U9225 (N_9225,N_135,N_1432);
nor U9226 (N_9226,N_2052,N_4061);
nor U9227 (N_9227,N_2553,N_2802);
and U9228 (N_9228,N_1431,N_1606);
nor U9229 (N_9229,N_293,N_2321);
nor U9230 (N_9230,N_41,N_504);
nand U9231 (N_9231,N_4375,N_2812);
or U9232 (N_9232,N_3078,N_398);
nor U9233 (N_9233,N_2675,N_2393);
nor U9234 (N_9234,N_1580,N_4244);
nor U9235 (N_9235,N_4729,N_4208);
nand U9236 (N_9236,N_4525,N_3166);
or U9237 (N_9237,N_4743,N_4642);
and U9238 (N_9238,N_4889,N_3636);
and U9239 (N_9239,N_3600,N_2504);
or U9240 (N_9240,N_462,N_3816);
or U9241 (N_9241,N_2218,N_2970);
nor U9242 (N_9242,N_4333,N_3305);
and U9243 (N_9243,N_128,N_2772);
and U9244 (N_9244,N_3540,N_1760);
and U9245 (N_9245,N_3844,N_443);
xor U9246 (N_9246,N_3587,N_4121);
and U9247 (N_9247,N_3174,N_728);
nor U9248 (N_9248,N_2088,N_769);
nor U9249 (N_9249,N_4536,N_920);
xor U9250 (N_9250,N_2099,N_2744);
or U9251 (N_9251,N_10,N_343);
and U9252 (N_9252,N_1408,N_472);
nor U9253 (N_9253,N_2357,N_1318);
nor U9254 (N_9254,N_397,N_2638);
or U9255 (N_9255,N_4449,N_3246);
nor U9256 (N_9256,N_558,N_4181);
nand U9257 (N_9257,N_980,N_1126);
or U9258 (N_9258,N_3394,N_2946);
and U9259 (N_9259,N_2827,N_1314);
nor U9260 (N_9260,N_755,N_2355);
nor U9261 (N_9261,N_2278,N_4383);
and U9262 (N_9262,N_67,N_1786);
nor U9263 (N_9263,N_2923,N_44);
or U9264 (N_9264,N_450,N_1260);
nor U9265 (N_9265,N_1897,N_3307);
nor U9266 (N_9266,N_723,N_4438);
and U9267 (N_9267,N_3168,N_1062);
nand U9268 (N_9268,N_3823,N_455);
or U9269 (N_9269,N_2952,N_3036);
nor U9270 (N_9270,N_2189,N_4816);
nand U9271 (N_9271,N_2192,N_4569);
nand U9272 (N_9272,N_2302,N_4229);
nand U9273 (N_9273,N_871,N_1145);
nor U9274 (N_9274,N_921,N_2348);
nor U9275 (N_9275,N_4163,N_4323);
xor U9276 (N_9276,N_1090,N_832);
nand U9277 (N_9277,N_2789,N_2326);
nor U9278 (N_9278,N_3422,N_768);
and U9279 (N_9279,N_785,N_2478);
nor U9280 (N_9280,N_3471,N_4642);
nand U9281 (N_9281,N_808,N_3908);
xnor U9282 (N_9282,N_4562,N_2518);
or U9283 (N_9283,N_3080,N_534);
nand U9284 (N_9284,N_1506,N_4467);
nand U9285 (N_9285,N_236,N_4446);
nand U9286 (N_9286,N_1555,N_2621);
nor U9287 (N_9287,N_615,N_1104);
nand U9288 (N_9288,N_3174,N_4302);
nand U9289 (N_9289,N_173,N_437);
nor U9290 (N_9290,N_138,N_3393);
xor U9291 (N_9291,N_1599,N_4776);
and U9292 (N_9292,N_1103,N_3963);
or U9293 (N_9293,N_3336,N_4605);
nor U9294 (N_9294,N_3142,N_4020);
nand U9295 (N_9295,N_4201,N_994);
or U9296 (N_9296,N_1796,N_2644);
nand U9297 (N_9297,N_2698,N_4735);
nand U9298 (N_9298,N_4269,N_464);
nor U9299 (N_9299,N_2203,N_1474);
nor U9300 (N_9300,N_4703,N_4900);
or U9301 (N_9301,N_2041,N_1254);
or U9302 (N_9302,N_2230,N_3071);
xnor U9303 (N_9303,N_2866,N_3211);
nand U9304 (N_9304,N_1551,N_2684);
and U9305 (N_9305,N_310,N_758);
nand U9306 (N_9306,N_524,N_535);
nand U9307 (N_9307,N_3493,N_3051);
or U9308 (N_9308,N_3932,N_791);
nor U9309 (N_9309,N_1180,N_220);
or U9310 (N_9310,N_1635,N_3511);
and U9311 (N_9311,N_4174,N_1122);
nor U9312 (N_9312,N_2257,N_2232);
nand U9313 (N_9313,N_4082,N_2455);
and U9314 (N_9314,N_968,N_2383);
nor U9315 (N_9315,N_799,N_3623);
and U9316 (N_9316,N_4419,N_2790);
nor U9317 (N_9317,N_1466,N_1609);
and U9318 (N_9318,N_4383,N_4860);
nor U9319 (N_9319,N_274,N_3963);
and U9320 (N_9320,N_1313,N_4374);
nor U9321 (N_9321,N_1351,N_3695);
or U9322 (N_9322,N_2857,N_3732);
nor U9323 (N_9323,N_4619,N_1273);
nor U9324 (N_9324,N_4811,N_1637);
and U9325 (N_9325,N_3770,N_4947);
nand U9326 (N_9326,N_2515,N_3648);
or U9327 (N_9327,N_2648,N_360);
nor U9328 (N_9328,N_3827,N_2789);
and U9329 (N_9329,N_3755,N_2571);
nor U9330 (N_9330,N_3628,N_3048);
nor U9331 (N_9331,N_3230,N_3129);
nand U9332 (N_9332,N_3194,N_4840);
nor U9333 (N_9333,N_3113,N_3849);
or U9334 (N_9334,N_2259,N_1125);
and U9335 (N_9335,N_1222,N_672);
and U9336 (N_9336,N_4560,N_680);
nor U9337 (N_9337,N_4730,N_2455);
or U9338 (N_9338,N_995,N_161);
and U9339 (N_9339,N_4073,N_1980);
or U9340 (N_9340,N_2175,N_59);
nor U9341 (N_9341,N_247,N_4846);
nand U9342 (N_9342,N_2737,N_2682);
or U9343 (N_9343,N_1940,N_427);
and U9344 (N_9344,N_1438,N_1678);
nor U9345 (N_9345,N_2368,N_284);
nor U9346 (N_9346,N_1074,N_1631);
or U9347 (N_9347,N_4339,N_2215);
or U9348 (N_9348,N_1650,N_4902);
or U9349 (N_9349,N_1538,N_4396);
or U9350 (N_9350,N_4734,N_1803);
nand U9351 (N_9351,N_3814,N_3561);
nand U9352 (N_9352,N_1522,N_1595);
nor U9353 (N_9353,N_2071,N_2239);
or U9354 (N_9354,N_2112,N_216);
and U9355 (N_9355,N_3120,N_2974);
nor U9356 (N_9356,N_4512,N_1195);
and U9357 (N_9357,N_1151,N_1418);
and U9358 (N_9358,N_1197,N_3770);
and U9359 (N_9359,N_1747,N_3610);
or U9360 (N_9360,N_1746,N_4075);
or U9361 (N_9361,N_300,N_246);
nand U9362 (N_9362,N_2315,N_3236);
and U9363 (N_9363,N_4068,N_4929);
and U9364 (N_9364,N_3045,N_357);
xor U9365 (N_9365,N_738,N_1556);
nand U9366 (N_9366,N_2215,N_4876);
nor U9367 (N_9367,N_2396,N_4510);
nor U9368 (N_9368,N_343,N_4364);
and U9369 (N_9369,N_342,N_2966);
nand U9370 (N_9370,N_3895,N_3423);
nand U9371 (N_9371,N_2566,N_3498);
nor U9372 (N_9372,N_3969,N_4000);
and U9373 (N_9373,N_4438,N_3463);
or U9374 (N_9374,N_2366,N_163);
or U9375 (N_9375,N_899,N_3870);
and U9376 (N_9376,N_4233,N_3916);
or U9377 (N_9377,N_4214,N_2700);
nor U9378 (N_9378,N_2982,N_4522);
and U9379 (N_9379,N_2311,N_3092);
or U9380 (N_9380,N_66,N_3173);
xnor U9381 (N_9381,N_1032,N_552);
or U9382 (N_9382,N_1731,N_4481);
or U9383 (N_9383,N_3696,N_2552);
nor U9384 (N_9384,N_1196,N_1749);
nand U9385 (N_9385,N_1659,N_4830);
nand U9386 (N_9386,N_1550,N_3845);
or U9387 (N_9387,N_4447,N_1936);
nor U9388 (N_9388,N_4768,N_1112);
and U9389 (N_9389,N_4690,N_732);
or U9390 (N_9390,N_3675,N_4240);
nand U9391 (N_9391,N_604,N_4650);
nor U9392 (N_9392,N_4086,N_1928);
nor U9393 (N_9393,N_123,N_1555);
and U9394 (N_9394,N_1808,N_4722);
and U9395 (N_9395,N_111,N_4124);
and U9396 (N_9396,N_3426,N_2277);
xnor U9397 (N_9397,N_3821,N_4325);
or U9398 (N_9398,N_4855,N_1333);
nor U9399 (N_9399,N_4123,N_826);
and U9400 (N_9400,N_3365,N_542);
or U9401 (N_9401,N_634,N_2082);
nor U9402 (N_9402,N_2816,N_416);
nor U9403 (N_9403,N_1069,N_3398);
nor U9404 (N_9404,N_2416,N_2517);
nor U9405 (N_9405,N_3528,N_1469);
xnor U9406 (N_9406,N_2371,N_2893);
or U9407 (N_9407,N_4956,N_4202);
and U9408 (N_9408,N_504,N_2010);
and U9409 (N_9409,N_1357,N_325);
xor U9410 (N_9410,N_3265,N_2905);
and U9411 (N_9411,N_3051,N_3769);
nor U9412 (N_9412,N_3188,N_1857);
and U9413 (N_9413,N_3160,N_945);
nor U9414 (N_9414,N_1486,N_3365);
nor U9415 (N_9415,N_4260,N_4456);
xor U9416 (N_9416,N_1627,N_2431);
and U9417 (N_9417,N_3358,N_3722);
or U9418 (N_9418,N_3274,N_2313);
nor U9419 (N_9419,N_705,N_2942);
or U9420 (N_9420,N_813,N_2662);
nor U9421 (N_9421,N_1069,N_99);
or U9422 (N_9422,N_443,N_3911);
nor U9423 (N_9423,N_302,N_1144);
nor U9424 (N_9424,N_1130,N_4991);
nor U9425 (N_9425,N_2614,N_4900);
or U9426 (N_9426,N_4784,N_1109);
nand U9427 (N_9427,N_2963,N_4416);
and U9428 (N_9428,N_1569,N_547);
or U9429 (N_9429,N_1945,N_4067);
nand U9430 (N_9430,N_4599,N_2374);
nor U9431 (N_9431,N_3100,N_1122);
nand U9432 (N_9432,N_3074,N_2742);
nand U9433 (N_9433,N_1284,N_1745);
nor U9434 (N_9434,N_551,N_648);
nor U9435 (N_9435,N_53,N_4008);
nor U9436 (N_9436,N_4753,N_3295);
nand U9437 (N_9437,N_735,N_2780);
nand U9438 (N_9438,N_220,N_2984);
or U9439 (N_9439,N_1277,N_258);
or U9440 (N_9440,N_2178,N_1995);
nand U9441 (N_9441,N_4972,N_3746);
or U9442 (N_9442,N_3200,N_4884);
nor U9443 (N_9443,N_491,N_4609);
nand U9444 (N_9444,N_711,N_1346);
or U9445 (N_9445,N_318,N_2862);
or U9446 (N_9446,N_739,N_3419);
and U9447 (N_9447,N_3881,N_331);
nand U9448 (N_9448,N_2187,N_2660);
xnor U9449 (N_9449,N_4406,N_1991);
or U9450 (N_9450,N_4334,N_1213);
nand U9451 (N_9451,N_1313,N_3888);
or U9452 (N_9452,N_1341,N_240);
nor U9453 (N_9453,N_301,N_3456);
or U9454 (N_9454,N_905,N_1631);
xor U9455 (N_9455,N_4010,N_1636);
and U9456 (N_9456,N_4780,N_4434);
or U9457 (N_9457,N_3607,N_639);
or U9458 (N_9458,N_3490,N_942);
nor U9459 (N_9459,N_3511,N_3889);
and U9460 (N_9460,N_189,N_4287);
nand U9461 (N_9461,N_2413,N_4205);
nand U9462 (N_9462,N_3346,N_373);
or U9463 (N_9463,N_1645,N_2296);
or U9464 (N_9464,N_49,N_2991);
nand U9465 (N_9465,N_1056,N_3000);
or U9466 (N_9466,N_2625,N_1371);
nor U9467 (N_9467,N_730,N_2554);
and U9468 (N_9468,N_2130,N_791);
or U9469 (N_9469,N_3068,N_4321);
or U9470 (N_9470,N_3793,N_2637);
and U9471 (N_9471,N_4508,N_760);
or U9472 (N_9472,N_1770,N_2425);
nor U9473 (N_9473,N_3218,N_1578);
and U9474 (N_9474,N_810,N_3237);
nand U9475 (N_9475,N_4165,N_3162);
and U9476 (N_9476,N_4614,N_603);
nor U9477 (N_9477,N_1609,N_4323);
xor U9478 (N_9478,N_1351,N_3127);
and U9479 (N_9479,N_803,N_3725);
nor U9480 (N_9480,N_3234,N_4180);
nor U9481 (N_9481,N_802,N_1987);
and U9482 (N_9482,N_4436,N_2873);
nor U9483 (N_9483,N_3467,N_2097);
or U9484 (N_9484,N_352,N_4644);
nand U9485 (N_9485,N_686,N_1291);
nor U9486 (N_9486,N_1564,N_1835);
or U9487 (N_9487,N_1900,N_4627);
or U9488 (N_9488,N_68,N_2559);
nor U9489 (N_9489,N_47,N_2395);
xor U9490 (N_9490,N_3542,N_2212);
nor U9491 (N_9491,N_1458,N_1382);
nand U9492 (N_9492,N_2373,N_714);
or U9493 (N_9493,N_2477,N_4248);
nor U9494 (N_9494,N_4436,N_3005);
and U9495 (N_9495,N_2555,N_4632);
nand U9496 (N_9496,N_757,N_1837);
nor U9497 (N_9497,N_674,N_378);
xnor U9498 (N_9498,N_279,N_4579);
nand U9499 (N_9499,N_3433,N_2656);
nor U9500 (N_9500,N_3288,N_4560);
nand U9501 (N_9501,N_4266,N_3734);
or U9502 (N_9502,N_4710,N_4344);
or U9503 (N_9503,N_1089,N_214);
or U9504 (N_9504,N_1059,N_4455);
or U9505 (N_9505,N_4644,N_1780);
nor U9506 (N_9506,N_306,N_3475);
nand U9507 (N_9507,N_4900,N_2247);
nor U9508 (N_9508,N_4131,N_2017);
nand U9509 (N_9509,N_4473,N_533);
xnor U9510 (N_9510,N_4156,N_3678);
and U9511 (N_9511,N_3700,N_2471);
nor U9512 (N_9512,N_1767,N_3050);
and U9513 (N_9513,N_3420,N_2870);
nor U9514 (N_9514,N_4903,N_1499);
and U9515 (N_9515,N_1898,N_4846);
and U9516 (N_9516,N_3744,N_3105);
nand U9517 (N_9517,N_4772,N_4540);
and U9518 (N_9518,N_1802,N_4036);
or U9519 (N_9519,N_2045,N_3067);
and U9520 (N_9520,N_3522,N_490);
and U9521 (N_9521,N_3297,N_297);
and U9522 (N_9522,N_2772,N_1594);
nor U9523 (N_9523,N_1614,N_1649);
or U9524 (N_9524,N_138,N_169);
and U9525 (N_9525,N_2170,N_2553);
nor U9526 (N_9526,N_4092,N_482);
nand U9527 (N_9527,N_4287,N_4855);
nand U9528 (N_9528,N_802,N_1114);
nor U9529 (N_9529,N_1253,N_1605);
nand U9530 (N_9530,N_2928,N_1135);
nand U9531 (N_9531,N_2755,N_4206);
and U9532 (N_9532,N_1451,N_2295);
nand U9533 (N_9533,N_4723,N_3784);
or U9534 (N_9534,N_36,N_4500);
or U9535 (N_9535,N_2674,N_4630);
or U9536 (N_9536,N_3575,N_2610);
nor U9537 (N_9537,N_4692,N_3321);
nor U9538 (N_9538,N_1725,N_1987);
nor U9539 (N_9539,N_1337,N_4944);
nor U9540 (N_9540,N_4351,N_1172);
or U9541 (N_9541,N_4523,N_4229);
nand U9542 (N_9542,N_2005,N_3055);
and U9543 (N_9543,N_1306,N_798);
nand U9544 (N_9544,N_2830,N_573);
and U9545 (N_9545,N_1431,N_1654);
nor U9546 (N_9546,N_1509,N_501);
and U9547 (N_9547,N_3207,N_3394);
and U9548 (N_9548,N_1670,N_4015);
or U9549 (N_9549,N_1418,N_3056);
nand U9550 (N_9550,N_4015,N_2260);
xor U9551 (N_9551,N_2731,N_799);
or U9552 (N_9552,N_1565,N_4256);
or U9553 (N_9553,N_4224,N_4837);
nand U9554 (N_9554,N_3033,N_1537);
nand U9555 (N_9555,N_3191,N_4362);
nor U9556 (N_9556,N_677,N_1241);
nand U9557 (N_9557,N_4318,N_2341);
or U9558 (N_9558,N_4126,N_2211);
nand U9559 (N_9559,N_4703,N_516);
nor U9560 (N_9560,N_1540,N_2927);
nand U9561 (N_9561,N_3767,N_3151);
nand U9562 (N_9562,N_129,N_2354);
and U9563 (N_9563,N_2376,N_2653);
and U9564 (N_9564,N_4640,N_3579);
nand U9565 (N_9565,N_3202,N_3775);
or U9566 (N_9566,N_3876,N_1040);
or U9567 (N_9567,N_3178,N_4165);
nand U9568 (N_9568,N_3112,N_364);
or U9569 (N_9569,N_4204,N_3769);
or U9570 (N_9570,N_1158,N_548);
nor U9571 (N_9571,N_1014,N_2970);
nor U9572 (N_9572,N_4425,N_3248);
or U9573 (N_9573,N_1368,N_376);
and U9574 (N_9574,N_1802,N_2911);
and U9575 (N_9575,N_1314,N_3784);
or U9576 (N_9576,N_1918,N_905);
and U9577 (N_9577,N_4001,N_4074);
or U9578 (N_9578,N_610,N_12);
and U9579 (N_9579,N_1946,N_3481);
or U9580 (N_9580,N_1433,N_3230);
nand U9581 (N_9581,N_3887,N_373);
xnor U9582 (N_9582,N_4480,N_1123);
nand U9583 (N_9583,N_2494,N_4044);
or U9584 (N_9584,N_3576,N_1114);
or U9585 (N_9585,N_103,N_3341);
nor U9586 (N_9586,N_829,N_4143);
nand U9587 (N_9587,N_731,N_1727);
or U9588 (N_9588,N_4014,N_3336);
nand U9589 (N_9589,N_4348,N_4141);
and U9590 (N_9590,N_3532,N_2928);
or U9591 (N_9591,N_1172,N_430);
and U9592 (N_9592,N_1650,N_4552);
and U9593 (N_9593,N_1749,N_3952);
nor U9594 (N_9594,N_3250,N_2559);
xnor U9595 (N_9595,N_3292,N_4877);
and U9596 (N_9596,N_3319,N_4166);
and U9597 (N_9597,N_4402,N_3945);
nand U9598 (N_9598,N_1402,N_2522);
nor U9599 (N_9599,N_4591,N_2767);
nand U9600 (N_9600,N_1442,N_1713);
nand U9601 (N_9601,N_3093,N_3939);
xor U9602 (N_9602,N_205,N_4955);
nor U9603 (N_9603,N_4427,N_1921);
or U9604 (N_9604,N_480,N_3384);
and U9605 (N_9605,N_739,N_3647);
nor U9606 (N_9606,N_3512,N_3963);
nor U9607 (N_9607,N_1798,N_1117);
or U9608 (N_9608,N_4950,N_2730);
nand U9609 (N_9609,N_3589,N_4567);
or U9610 (N_9610,N_4021,N_3064);
and U9611 (N_9611,N_2853,N_3521);
nor U9612 (N_9612,N_1293,N_3851);
or U9613 (N_9613,N_1268,N_1536);
nor U9614 (N_9614,N_548,N_1163);
or U9615 (N_9615,N_1473,N_4061);
xor U9616 (N_9616,N_2762,N_3337);
or U9617 (N_9617,N_1553,N_2533);
nor U9618 (N_9618,N_4871,N_4741);
and U9619 (N_9619,N_4636,N_2922);
xnor U9620 (N_9620,N_469,N_2290);
xor U9621 (N_9621,N_2303,N_4552);
or U9622 (N_9622,N_4610,N_1896);
and U9623 (N_9623,N_2854,N_1623);
and U9624 (N_9624,N_4638,N_3076);
nor U9625 (N_9625,N_4234,N_3506);
or U9626 (N_9626,N_2280,N_4659);
nor U9627 (N_9627,N_3917,N_1016);
xor U9628 (N_9628,N_2083,N_417);
or U9629 (N_9629,N_4263,N_3146);
or U9630 (N_9630,N_2779,N_2825);
nand U9631 (N_9631,N_257,N_383);
and U9632 (N_9632,N_3878,N_1835);
or U9633 (N_9633,N_1105,N_4630);
or U9634 (N_9634,N_3017,N_782);
nand U9635 (N_9635,N_3617,N_3813);
and U9636 (N_9636,N_2209,N_253);
or U9637 (N_9637,N_1804,N_47);
and U9638 (N_9638,N_3425,N_3334);
nor U9639 (N_9639,N_4839,N_3988);
and U9640 (N_9640,N_2922,N_840);
and U9641 (N_9641,N_2687,N_4949);
or U9642 (N_9642,N_4263,N_963);
nor U9643 (N_9643,N_3054,N_254);
nor U9644 (N_9644,N_2103,N_4770);
and U9645 (N_9645,N_4280,N_4247);
nand U9646 (N_9646,N_1184,N_3811);
and U9647 (N_9647,N_3690,N_2918);
nand U9648 (N_9648,N_3442,N_2574);
nor U9649 (N_9649,N_3470,N_4519);
or U9650 (N_9650,N_3048,N_3058);
or U9651 (N_9651,N_453,N_801);
or U9652 (N_9652,N_1691,N_215);
and U9653 (N_9653,N_2646,N_1078);
nand U9654 (N_9654,N_1837,N_3980);
nor U9655 (N_9655,N_4371,N_1976);
nor U9656 (N_9656,N_1099,N_1504);
nand U9657 (N_9657,N_494,N_4612);
nor U9658 (N_9658,N_2439,N_1339);
and U9659 (N_9659,N_4773,N_2044);
nand U9660 (N_9660,N_1887,N_3340);
nor U9661 (N_9661,N_4451,N_903);
nand U9662 (N_9662,N_277,N_2156);
or U9663 (N_9663,N_2020,N_3221);
and U9664 (N_9664,N_1788,N_348);
nand U9665 (N_9665,N_1102,N_613);
and U9666 (N_9666,N_1491,N_1204);
and U9667 (N_9667,N_3165,N_1332);
or U9668 (N_9668,N_4828,N_3410);
and U9669 (N_9669,N_1398,N_2233);
or U9670 (N_9670,N_2274,N_937);
or U9671 (N_9671,N_839,N_2227);
and U9672 (N_9672,N_3163,N_4176);
nand U9673 (N_9673,N_4970,N_4220);
nor U9674 (N_9674,N_2759,N_3088);
nand U9675 (N_9675,N_691,N_90);
and U9676 (N_9676,N_4978,N_2501);
xnor U9677 (N_9677,N_1777,N_4411);
and U9678 (N_9678,N_3345,N_100);
nand U9679 (N_9679,N_2433,N_3115);
xor U9680 (N_9680,N_2590,N_178);
nand U9681 (N_9681,N_2406,N_2338);
nor U9682 (N_9682,N_2007,N_940);
and U9683 (N_9683,N_3801,N_2511);
nor U9684 (N_9684,N_3823,N_3485);
nor U9685 (N_9685,N_1806,N_1129);
nor U9686 (N_9686,N_2516,N_4594);
xnor U9687 (N_9687,N_4136,N_763);
xnor U9688 (N_9688,N_4605,N_77);
nor U9689 (N_9689,N_2069,N_186);
and U9690 (N_9690,N_4354,N_2870);
nand U9691 (N_9691,N_2018,N_1919);
and U9692 (N_9692,N_1138,N_4304);
and U9693 (N_9693,N_3341,N_3310);
or U9694 (N_9694,N_4184,N_4088);
nor U9695 (N_9695,N_4506,N_4866);
and U9696 (N_9696,N_830,N_3249);
nand U9697 (N_9697,N_3488,N_1752);
nor U9698 (N_9698,N_2600,N_157);
nand U9699 (N_9699,N_1121,N_2501);
or U9700 (N_9700,N_1032,N_953);
or U9701 (N_9701,N_3671,N_688);
or U9702 (N_9702,N_816,N_1217);
and U9703 (N_9703,N_766,N_1458);
nand U9704 (N_9704,N_1517,N_4254);
nand U9705 (N_9705,N_432,N_1422);
or U9706 (N_9706,N_4410,N_1538);
nor U9707 (N_9707,N_4322,N_468);
nand U9708 (N_9708,N_53,N_2604);
or U9709 (N_9709,N_2317,N_1998);
nand U9710 (N_9710,N_1590,N_3536);
or U9711 (N_9711,N_2531,N_3571);
nor U9712 (N_9712,N_957,N_7);
and U9713 (N_9713,N_1137,N_1530);
nand U9714 (N_9714,N_4036,N_669);
xor U9715 (N_9715,N_3030,N_3803);
nand U9716 (N_9716,N_1095,N_4440);
nor U9717 (N_9717,N_3122,N_4129);
or U9718 (N_9718,N_424,N_2529);
nand U9719 (N_9719,N_226,N_4856);
xnor U9720 (N_9720,N_3859,N_2224);
and U9721 (N_9721,N_117,N_3198);
nand U9722 (N_9722,N_4742,N_984);
or U9723 (N_9723,N_669,N_4424);
and U9724 (N_9724,N_2941,N_2966);
and U9725 (N_9725,N_3323,N_2904);
or U9726 (N_9726,N_4924,N_4066);
and U9727 (N_9727,N_3590,N_1178);
nand U9728 (N_9728,N_534,N_1294);
and U9729 (N_9729,N_4439,N_1108);
xor U9730 (N_9730,N_2742,N_2126);
or U9731 (N_9731,N_4343,N_4097);
and U9732 (N_9732,N_2600,N_4005);
and U9733 (N_9733,N_3527,N_2483);
and U9734 (N_9734,N_4375,N_2150);
or U9735 (N_9735,N_4496,N_182);
nand U9736 (N_9736,N_1016,N_4854);
nor U9737 (N_9737,N_3602,N_4670);
or U9738 (N_9738,N_4634,N_3739);
nor U9739 (N_9739,N_1160,N_3642);
and U9740 (N_9740,N_476,N_3841);
nor U9741 (N_9741,N_1442,N_4352);
or U9742 (N_9742,N_4035,N_4271);
or U9743 (N_9743,N_570,N_1181);
or U9744 (N_9744,N_4917,N_2574);
and U9745 (N_9745,N_1192,N_2122);
and U9746 (N_9746,N_799,N_3460);
xor U9747 (N_9747,N_1460,N_4706);
and U9748 (N_9748,N_2679,N_3607);
or U9749 (N_9749,N_3609,N_4693);
or U9750 (N_9750,N_3869,N_2957);
nand U9751 (N_9751,N_2314,N_570);
or U9752 (N_9752,N_3893,N_706);
xor U9753 (N_9753,N_1407,N_1770);
or U9754 (N_9754,N_4780,N_4896);
and U9755 (N_9755,N_446,N_241);
nand U9756 (N_9756,N_2943,N_436);
nand U9757 (N_9757,N_2548,N_4440);
nand U9758 (N_9758,N_3846,N_1937);
nor U9759 (N_9759,N_2352,N_3565);
and U9760 (N_9760,N_2954,N_3668);
and U9761 (N_9761,N_4416,N_4611);
xor U9762 (N_9762,N_1405,N_1071);
or U9763 (N_9763,N_518,N_1532);
nand U9764 (N_9764,N_100,N_2340);
and U9765 (N_9765,N_4686,N_4294);
and U9766 (N_9766,N_3253,N_2549);
xnor U9767 (N_9767,N_4958,N_3567);
nand U9768 (N_9768,N_4153,N_2260);
xor U9769 (N_9769,N_78,N_2646);
nand U9770 (N_9770,N_4067,N_4478);
or U9771 (N_9771,N_1216,N_3987);
nand U9772 (N_9772,N_4836,N_4866);
nand U9773 (N_9773,N_3195,N_1085);
nor U9774 (N_9774,N_2108,N_664);
nor U9775 (N_9775,N_1732,N_4517);
or U9776 (N_9776,N_1568,N_1808);
nor U9777 (N_9777,N_4463,N_4983);
or U9778 (N_9778,N_1191,N_3571);
and U9779 (N_9779,N_285,N_1872);
nor U9780 (N_9780,N_1832,N_109);
and U9781 (N_9781,N_3175,N_4280);
or U9782 (N_9782,N_3890,N_1178);
nand U9783 (N_9783,N_1606,N_2413);
or U9784 (N_9784,N_1376,N_3023);
nor U9785 (N_9785,N_4630,N_455);
or U9786 (N_9786,N_2794,N_4532);
nor U9787 (N_9787,N_4128,N_664);
and U9788 (N_9788,N_2757,N_1709);
nand U9789 (N_9789,N_2593,N_2380);
nand U9790 (N_9790,N_256,N_3414);
nand U9791 (N_9791,N_2692,N_1633);
xnor U9792 (N_9792,N_1542,N_3888);
nand U9793 (N_9793,N_4029,N_3163);
nand U9794 (N_9794,N_1706,N_3635);
and U9795 (N_9795,N_701,N_241);
or U9796 (N_9796,N_4391,N_4517);
xor U9797 (N_9797,N_1125,N_4327);
or U9798 (N_9798,N_4834,N_2325);
nor U9799 (N_9799,N_1865,N_1903);
and U9800 (N_9800,N_3717,N_799);
and U9801 (N_9801,N_1178,N_2172);
nor U9802 (N_9802,N_4582,N_3311);
and U9803 (N_9803,N_1165,N_2419);
or U9804 (N_9804,N_950,N_3767);
or U9805 (N_9805,N_4492,N_802);
or U9806 (N_9806,N_1276,N_3947);
xnor U9807 (N_9807,N_1938,N_2160);
and U9808 (N_9808,N_2276,N_4388);
and U9809 (N_9809,N_4235,N_2483);
and U9810 (N_9810,N_1358,N_3575);
and U9811 (N_9811,N_4741,N_4184);
nand U9812 (N_9812,N_1537,N_3146);
nand U9813 (N_9813,N_731,N_4259);
xnor U9814 (N_9814,N_2784,N_325);
nor U9815 (N_9815,N_3072,N_3020);
and U9816 (N_9816,N_1290,N_945);
nor U9817 (N_9817,N_3878,N_407);
and U9818 (N_9818,N_3417,N_2982);
or U9819 (N_9819,N_1797,N_179);
nor U9820 (N_9820,N_4852,N_3003);
nor U9821 (N_9821,N_2972,N_1706);
xor U9822 (N_9822,N_2938,N_2648);
nand U9823 (N_9823,N_3427,N_1449);
nand U9824 (N_9824,N_4805,N_4402);
nand U9825 (N_9825,N_1756,N_2235);
or U9826 (N_9826,N_2388,N_1429);
nor U9827 (N_9827,N_4777,N_2152);
xnor U9828 (N_9828,N_3018,N_2459);
nor U9829 (N_9829,N_4355,N_1129);
nor U9830 (N_9830,N_3170,N_3278);
or U9831 (N_9831,N_4917,N_1458);
xnor U9832 (N_9832,N_511,N_445);
and U9833 (N_9833,N_4004,N_3955);
nand U9834 (N_9834,N_3381,N_1837);
nand U9835 (N_9835,N_369,N_1873);
or U9836 (N_9836,N_2813,N_4326);
and U9837 (N_9837,N_4512,N_4723);
and U9838 (N_9838,N_1945,N_1219);
or U9839 (N_9839,N_3036,N_3996);
xor U9840 (N_9840,N_2959,N_3320);
or U9841 (N_9841,N_4131,N_3166);
nor U9842 (N_9842,N_1838,N_3768);
and U9843 (N_9843,N_2836,N_2308);
nor U9844 (N_9844,N_2354,N_849);
nor U9845 (N_9845,N_3903,N_3284);
nand U9846 (N_9846,N_1148,N_2224);
and U9847 (N_9847,N_713,N_4854);
nand U9848 (N_9848,N_3116,N_4832);
nor U9849 (N_9849,N_3355,N_735);
or U9850 (N_9850,N_2110,N_3122);
nor U9851 (N_9851,N_4341,N_4980);
nand U9852 (N_9852,N_1625,N_4700);
and U9853 (N_9853,N_1011,N_2641);
or U9854 (N_9854,N_2151,N_4247);
or U9855 (N_9855,N_845,N_1191);
xor U9856 (N_9856,N_1814,N_4606);
or U9857 (N_9857,N_3387,N_3239);
or U9858 (N_9858,N_1003,N_3718);
nand U9859 (N_9859,N_4254,N_1393);
or U9860 (N_9860,N_4272,N_4021);
nand U9861 (N_9861,N_126,N_4986);
and U9862 (N_9862,N_4234,N_764);
nand U9863 (N_9863,N_4865,N_4578);
and U9864 (N_9864,N_3133,N_350);
or U9865 (N_9865,N_1264,N_310);
nand U9866 (N_9866,N_4873,N_1707);
xor U9867 (N_9867,N_3771,N_1684);
or U9868 (N_9868,N_2618,N_3580);
nand U9869 (N_9869,N_3502,N_760);
and U9870 (N_9870,N_459,N_4049);
and U9871 (N_9871,N_3658,N_1742);
nor U9872 (N_9872,N_2722,N_2458);
nand U9873 (N_9873,N_2904,N_1151);
nor U9874 (N_9874,N_3591,N_792);
xnor U9875 (N_9875,N_4290,N_3509);
or U9876 (N_9876,N_1297,N_2843);
nor U9877 (N_9877,N_4950,N_2878);
or U9878 (N_9878,N_3132,N_2077);
xnor U9879 (N_9879,N_1827,N_3691);
nand U9880 (N_9880,N_1520,N_4494);
nor U9881 (N_9881,N_1052,N_3974);
nor U9882 (N_9882,N_4369,N_2786);
nand U9883 (N_9883,N_1824,N_2006);
or U9884 (N_9884,N_1214,N_2570);
nor U9885 (N_9885,N_4125,N_3206);
and U9886 (N_9886,N_1218,N_3665);
and U9887 (N_9887,N_4184,N_2000);
nand U9888 (N_9888,N_434,N_4734);
or U9889 (N_9889,N_2546,N_944);
or U9890 (N_9890,N_2217,N_3786);
or U9891 (N_9891,N_612,N_3829);
nor U9892 (N_9892,N_3102,N_1329);
xor U9893 (N_9893,N_330,N_2333);
nor U9894 (N_9894,N_2191,N_2534);
and U9895 (N_9895,N_413,N_728);
xnor U9896 (N_9896,N_4079,N_3419);
or U9897 (N_9897,N_2556,N_2012);
or U9898 (N_9898,N_1841,N_4119);
nand U9899 (N_9899,N_4834,N_2990);
nand U9900 (N_9900,N_3783,N_104);
nor U9901 (N_9901,N_3341,N_3866);
or U9902 (N_9902,N_4603,N_4936);
and U9903 (N_9903,N_532,N_2134);
or U9904 (N_9904,N_1232,N_2928);
or U9905 (N_9905,N_260,N_2090);
nand U9906 (N_9906,N_4124,N_3989);
or U9907 (N_9907,N_3063,N_2361);
nor U9908 (N_9908,N_4031,N_4133);
and U9909 (N_9909,N_134,N_4733);
or U9910 (N_9910,N_1087,N_1844);
nor U9911 (N_9911,N_4362,N_4946);
or U9912 (N_9912,N_868,N_1674);
or U9913 (N_9913,N_4832,N_803);
nand U9914 (N_9914,N_4733,N_634);
xnor U9915 (N_9915,N_3919,N_1100);
or U9916 (N_9916,N_234,N_1289);
xor U9917 (N_9917,N_711,N_3413);
or U9918 (N_9918,N_391,N_1028);
or U9919 (N_9919,N_2572,N_4245);
and U9920 (N_9920,N_3784,N_865);
and U9921 (N_9921,N_933,N_954);
or U9922 (N_9922,N_4594,N_3376);
nor U9923 (N_9923,N_4712,N_4842);
and U9924 (N_9924,N_52,N_1435);
and U9925 (N_9925,N_2789,N_1362);
and U9926 (N_9926,N_2389,N_4935);
nor U9927 (N_9927,N_926,N_3074);
or U9928 (N_9928,N_1839,N_4729);
nand U9929 (N_9929,N_1531,N_347);
and U9930 (N_9930,N_1649,N_968);
nand U9931 (N_9931,N_4061,N_3242);
or U9932 (N_9932,N_870,N_4812);
nor U9933 (N_9933,N_1508,N_1007);
nor U9934 (N_9934,N_1757,N_515);
and U9935 (N_9935,N_963,N_3286);
nand U9936 (N_9936,N_2375,N_4140);
nand U9937 (N_9937,N_741,N_3648);
nor U9938 (N_9938,N_1167,N_3624);
and U9939 (N_9939,N_1016,N_2126);
nor U9940 (N_9940,N_1565,N_3253);
and U9941 (N_9941,N_4961,N_1183);
nand U9942 (N_9942,N_1364,N_266);
nand U9943 (N_9943,N_4783,N_2449);
nor U9944 (N_9944,N_1334,N_4790);
nand U9945 (N_9945,N_2308,N_2330);
or U9946 (N_9946,N_4207,N_887);
nand U9947 (N_9947,N_4280,N_3211);
nand U9948 (N_9948,N_1959,N_76);
nand U9949 (N_9949,N_2027,N_2388);
and U9950 (N_9950,N_3445,N_3751);
xor U9951 (N_9951,N_1908,N_4180);
nor U9952 (N_9952,N_1643,N_2765);
nand U9953 (N_9953,N_468,N_541);
nor U9954 (N_9954,N_2976,N_3001);
or U9955 (N_9955,N_648,N_2202);
nor U9956 (N_9956,N_2106,N_4251);
or U9957 (N_9957,N_4355,N_4182);
or U9958 (N_9958,N_4140,N_3529);
and U9959 (N_9959,N_3877,N_2260);
nor U9960 (N_9960,N_2088,N_4135);
xor U9961 (N_9961,N_1159,N_4617);
or U9962 (N_9962,N_4244,N_1635);
xnor U9963 (N_9963,N_2483,N_1812);
nand U9964 (N_9964,N_593,N_2528);
nand U9965 (N_9965,N_1990,N_2611);
and U9966 (N_9966,N_4781,N_1260);
and U9967 (N_9967,N_3472,N_2651);
xnor U9968 (N_9968,N_2605,N_4004);
nor U9969 (N_9969,N_3679,N_812);
or U9970 (N_9970,N_1161,N_2505);
nor U9971 (N_9971,N_1126,N_52);
and U9972 (N_9972,N_1164,N_2969);
xor U9973 (N_9973,N_27,N_3785);
nor U9974 (N_9974,N_4858,N_3484);
or U9975 (N_9975,N_1622,N_403);
or U9976 (N_9976,N_4810,N_4451);
nand U9977 (N_9977,N_66,N_37);
nand U9978 (N_9978,N_1454,N_2703);
nor U9979 (N_9979,N_847,N_1147);
nor U9980 (N_9980,N_840,N_4447);
nor U9981 (N_9981,N_1309,N_1183);
or U9982 (N_9982,N_3465,N_4390);
or U9983 (N_9983,N_4487,N_4927);
or U9984 (N_9984,N_2283,N_2091);
or U9985 (N_9985,N_905,N_3384);
nand U9986 (N_9986,N_3411,N_1282);
nand U9987 (N_9987,N_1110,N_3024);
nor U9988 (N_9988,N_2348,N_3529);
nor U9989 (N_9989,N_780,N_538);
or U9990 (N_9990,N_4009,N_4321);
nand U9991 (N_9991,N_1437,N_1837);
nor U9992 (N_9992,N_4319,N_1223);
xnor U9993 (N_9993,N_1557,N_74);
and U9994 (N_9994,N_4298,N_674);
and U9995 (N_9995,N_1422,N_4067);
nor U9996 (N_9996,N_3383,N_55);
nand U9997 (N_9997,N_3225,N_4103);
and U9998 (N_9998,N_1425,N_857);
and U9999 (N_9999,N_2326,N_1973);
nor U10000 (N_10000,N_5649,N_7876);
or U10001 (N_10001,N_7471,N_7198);
and U10002 (N_10002,N_7123,N_9036);
nor U10003 (N_10003,N_5194,N_5899);
nand U10004 (N_10004,N_6171,N_7040);
nand U10005 (N_10005,N_8929,N_6071);
or U10006 (N_10006,N_8940,N_5879);
or U10007 (N_10007,N_7808,N_9822);
nand U10008 (N_10008,N_9844,N_9725);
nor U10009 (N_10009,N_5225,N_5255);
or U10010 (N_10010,N_7813,N_9897);
nor U10011 (N_10011,N_9669,N_9419);
or U10012 (N_10012,N_6388,N_6989);
nor U10013 (N_10013,N_9227,N_7036);
nand U10014 (N_10014,N_7935,N_8764);
xnor U10015 (N_10015,N_5990,N_7320);
and U10016 (N_10016,N_7892,N_9717);
nand U10017 (N_10017,N_8139,N_7174);
xnor U10018 (N_10018,N_9362,N_6583);
and U10019 (N_10019,N_9743,N_5207);
or U10020 (N_10020,N_8721,N_7529);
xor U10021 (N_10021,N_9349,N_7060);
nor U10022 (N_10022,N_8798,N_6074);
nor U10023 (N_10023,N_7211,N_7694);
and U10024 (N_10024,N_8009,N_8039);
or U10025 (N_10025,N_5617,N_7362);
or U10026 (N_10026,N_7696,N_8274);
nor U10027 (N_10027,N_5790,N_8404);
or U10028 (N_10028,N_5144,N_6352);
or U10029 (N_10029,N_6220,N_9054);
or U10030 (N_10030,N_5286,N_7888);
nand U10031 (N_10031,N_9931,N_9788);
and U10032 (N_10032,N_8273,N_6005);
nand U10033 (N_10033,N_7941,N_8614);
and U10034 (N_10034,N_9285,N_9826);
nor U10035 (N_10035,N_5957,N_5741);
nor U10036 (N_10036,N_6937,N_7121);
nand U10037 (N_10037,N_8248,N_9742);
nand U10038 (N_10038,N_8724,N_9014);
nand U10039 (N_10039,N_6905,N_7252);
nor U10040 (N_10040,N_5665,N_5468);
nand U10041 (N_10041,N_7844,N_9495);
and U10042 (N_10042,N_9821,N_6666);
and U10043 (N_10043,N_8576,N_5680);
nor U10044 (N_10044,N_5750,N_5052);
or U10045 (N_10045,N_9368,N_5441);
or U10046 (N_10046,N_8328,N_9566);
and U10047 (N_10047,N_5925,N_8971);
xor U10048 (N_10048,N_6477,N_6415);
and U10049 (N_10049,N_7422,N_5009);
nand U10050 (N_10050,N_9574,N_6286);
or U10051 (N_10051,N_6073,N_9787);
nor U10052 (N_10052,N_9924,N_7641);
nor U10053 (N_10053,N_5094,N_9379);
and U10054 (N_10054,N_9217,N_5498);
and U10055 (N_10055,N_9012,N_8413);
nand U10056 (N_10056,N_6459,N_6120);
nand U10057 (N_10057,N_5252,N_9329);
nor U10058 (N_10058,N_6257,N_9492);
nand U10059 (N_10059,N_6068,N_9575);
nand U10060 (N_10060,N_6125,N_5438);
nor U10061 (N_10061,N_9613,N_7091);
xor U10062 (N_10062,N_7009,N_5206);
nand U10063 (N_10063,N_8398,N_9758);
nor U10064 (N_10064,N_7236,N_6264);
and U10065 (N_10065,N_5942,N_5014);
nand U10066 (N_10066,N_5743,N_8411);
or U10067 (N_10067,N_8160,N_5291);
nor U10068 (N_10068,N_8163,N_9837);
nor U10069 (N_10069,N_9972,N_6662);
nand U10070 (N_10070,N_6924,N_9569);
nand U10071 (N_10071,N_8106,N_7113);
and U10072 (N_10072,N_9614,N_8321);
nor U10073 (N_10073,N_9868,N_6488);
or U10074 (N_10074,N_6793,N_9775);
or U10075 (N_10075,N_8080,N_9366);
nand U10076 (N_10076,N_9702,N_5547);
or U10077 (N_10077,N_8640,N_8800);
nand U10078 (N_10078,N_5030,N_7991);
nor U10079 (N_10079,N_5857,N_6469);
and U10080 (N_10080,N_9802,N_5415);
nand U10081 (N_10081,N_7660,N_8966);
and U10082 (N_10082,N_5368,N_5417);
or U10083 (N_10083,N_8405,N_7470);
or U10084 (N_10084,N_8378,N_5082);
and U10085 (N_10085,N_9185,N_7788);
or U10086 (N_10086,N_9796,N_6768);
or U10087 (N_10087,N_6996,N_9245);
and U10088 (N_10088,N_6288,N_8133);
and U10089 (N_10089,N_9988,N_6334);
or U10090 (N_10090,N_9771,N_6077);
nand U10091 (N_10091,N_7648,N_5972);
xor U10092 (N_10092,N_5530,N_6336);
or U10093 (N_10093,N_8412,N_6133);
nand U10094 (N_10094,N_6997,N_5039);
nand U10095 (N_10095,N_9451,N_6833);
nor U10096 (N_10096,N_7084,N_7406);
and U10097 (N_10097,N_7322,N_9374);
and U10098 (N_10098,N_7718,N_5936);
nand U10099 (N_10099,N_7631,N_6323);
and U10100 (N_10100,N_8366,N_8192);
and U10101 (N_10101,N_6260,N_7834);
nor U10102 (N_10102,N_7617,N_9405);
and U10103 (N_10103,N_5639,N_8898);
and U10104 (N_10104,N_9096,N_7469);
nor U10105 (N_10105,N_7147,N_7081);
nor U10106 (N_10106,N_7150,N_6880);
or U10107 (N_10107,N_7549,N_6080);
nor U10108 (N_10108,N_5213,N_8842);
nand U10109 (N_10109,N_5200,N_6660);
nor U10110 (N_10110,N_8060,N_8058);
nor U10111 (N_10111,N_8628,N_7971);
nand U10112 (N_10112,N_5054,N_6229);
nor U10113 (N_10113,N_5120,N_7429);
nand U10114 (N_10114,N_7784,N_7143);
nand U10115 (N_10115,N_7608,N_8341);
nor U10116 (N_10116,N_8194,N_9387);
and U10117 (N_10117,N_9886,N_7911);
nand U10118 (N_10118,N_6308,N_8262);
nor U10119 (N_10119,N_8770,N_7160);
nor U10120 (N_10120,N_9101,N_7110);
and U10121 (N_10121,N_8708,N_8758);
nand U10122 (N_10122,N_7568,N_5823);
and U10123 (N_10123,N_8911,N_8023);
nand U10124 (N_10124,N_8678,N_7595);
nor U10125 (N_10125,N_7449,N_9081);
or U10126 (N_10126,N_5600,N_7933);
or U10127 (N_10127,N_9567,N_9730);
and U10128 (N_10128,N_6084,N_9425);
and U10129 (N_10129,N_8061,N_9734);
nand U10130 (N_10130,N_7129,N_6735);
or U10131 (N_10131,N_7651,N_6703);
or U10132 (N_10132,N_6566,N_6526);
nand U10133 (N_10133,N_6023,N_8070);
or U10134 (N_10134,N_8314,N_9146);
and U10135 (N_10135,N_6307,N_8443);
or U10136 (N_10136,N_6726,N_6127);
nand U10137 (N_10137,N_7779,N_9439);
nand U10138 (N_10138,N_5168,N_8199);
nor U10139 (N_10139,N_9556,N_6507);
and U10140 (N_10140,N_6092,N_5129);
or U10141 (N_10141,N_9793,N_9378);
nor U10142 (N_10142,N_6378,N_8693);
nor U10143 (N_10143,N_8822,N_5379);
or U10144 (N_10144,N_9183,N_7261);
and U10145 (N_10145,N_6917,N_5980);
or U10146 (N_10146,N_7321,N_9208);
and U10147 (N_10147,N_5926,N_5888);
and U10148 (N_10148,N_6647,N_9710);
or U10149 (N_10149,N_6346,N_7639);
nor U10150 (N_10150,N_6528,N_5138);
or U10151 (N_10151,N_7116,N_9021);
and U10152 (N_10152,N_8930,N_7524);
nor U10153 (N_10153,N_8004,N_7542);
or U10154 (N_10154,N_8575,N_7293);
and U10155 (N_10155,N_7890,N_6207);
nor U10156 (N_10156,N_9949,N_9141);
and U10157 (N_10157,N_6197,N_6659);
or U10158 (N_10158,N_7825,N_5999);
xor U10159 (N_10159,N_6813,N_6716);
or U10160 (N_10160,N_9635,N_7672);
nand U10161 (N_10161,N_8333,N_6501);
or U10162 (N_10162,N_6369,N_9709);
nor U10163 (N_10163,N_9565,N_7936);
nor U10164 (N_10164,N_6331,N_5018);
nor U10165 (N_10165,N_5278,N_7872);
nor U10166 (N_10166,N_6798,N_8242);
or U10167 (N_10167,N_7340,N_6912);
or U10168 (N_10168,N_8539,N_9713);
nor U10169 (N_10169,N_5623,N_8688);
or U10170 (N_10170,N_6474,N_6343);
nor U10171 (N_10171,N_9571,N_9319);
nor U10172 (N_10172,N_7454,N_5222);
nand U10173 (N_10173,N_9736,N_8292);
or U10174 (N_10174,N_8702,N_9213);
nor U10175 (N_10175,N_9699,N_8747);
and U10176 (N_10176,N_6616,N_8980);
or U10177 (N_10177,N_6141,N_5075);
nand U10178 (N_10178,N_7120,N_7783);
nor U10179 (N_10179,N_7804,N_8953);
and U10180 (N_10180,N_5552,N_9925);
nor U10181 (N_10181,N_5603,N_8277);
nand U10182 (N_10182,N_9573,N_8237);
nand U10183 (N_10183,N_8159,N_8261);
and U10184 (N_10184,N_6658,N_6100);
nand U10185 (N_10185,N_6419,N_9643);
nor U10186 (N_10186,N_9063,N_8045);
nor U10187 (N_10187,N_6743,N_7332);
nand U10188 (N_10188,N_8958,N_7386);
and U10189 (N_10189,N_5924,N_8959);
or U10190 (N_10190,N_6497,N_9662);
or U10191 (N_10191,N_6253,N_7433);
or U10192 (N_10192,N_9392,N_6039);
nor U10193 (N_10193,N_7766,N_6856);
and U10194 (N_10194,N_7959,N_7507);
nor U10195 (N_10195,N_5059,N_5243);
nor U10196 (N_10196,N_8742,N_6215);
and U10197 (N_10197,N_5845,N_9448);
xor U10198 (N_10198,N_8428,N_8505);
nor U10199 (N_10199,N_5581,N_7535);
or U10200 (N_10200,N_6262,N_8989);
xnor U10201 (N_10201,N_7823,N_5409);
or U10202 (N_10202,N_8228,N_6724);
nor U10203 (N_10203,N_7038,N_9267);
and U10204 (N_10204,N_6928,N_5986);
xnor U10205 (N_10205,N_5418,N_9422);
xnor U10206 (N_10206,N_9391,N_7791);
nand U10207 (N_10207,N_7680,N_5152);
nor U10208 (N_10208,N_9407,N_7064);
and U10209 (N_10209,N_7401,N_7917);
nor U10210 (N_10210,N_8063,N_6102);
or U10211 (N_10211,N_9884,N_9470);
and U10212 (N_10212,N_8586,N_9660);
nand U10213 (N_10213,N_8831,N_6000);
and U10214 (N_10214,N_8837,N_7200);
nand U10215 (N_10215,N_9905,N_8786);
nand U10216 (N_10216,N_5551,N_5556);
nor U10217 (N_10217,N_5852,N_7603);
or U10218 (N_10218,N_8543,N_7135);
xor U10219 (N_10219,N_5933,N_6546);
or U10220 (N_10220,N_5481,N_8790);
or U10221 (N_10221,N_9632,N_8182);
and U10222 (N_10222,N_6097,N_8105);
nand U10223 (N_10223,N_8801,N_9618);
and U10224 (N_10224,N_8491,N_7452);
xnor U10225 (N_10225,N_9863,N_8797);
or U10226 (N_10226,N_8089,N_9845);
or U10227 (N_10227,N_8281,N_6509);
or U10228 (N_10228,N_8014,N_7356);
nor U10229 (N_10229,N_9105,N_6302);
nor U10230 (N_10230,N_6978,N_9854);
nand U10231 (N_10231,N_6250,N_7707);
xor U10232 (N_10232,N_8901,N_6910);
xnor U10233 (N_10233,N_7606,N_5470);
nor U10234 (N_10234,N_9969,N_5906);
nor U10235 (N_10235,N_5602,N_6019);
and U10236 (N_10236,N_7013,N_7565);
or U10237 (N_10237,N_9927,N_5722);
nand U10238 (N_10238,N_8087,N_7809);
xor U10239 (N_10239,N_8463,N_9965);
or U10240 (N_10240,N_5491,N_8767);
nand U10241 (N_10241,N_5615,N_6188);
nand U10242 (N_10242,N_6840,N_7914);
nor U10243 (N_10243,N_5251,N_5087);
and U10244 (N_10244,N_7430,N_8353);
nor U10245 (N_10245,N_7836,N_7913);
and U10246 (N_10246,N_6961,N_5661);
and U10247 (N_10247,N_5482,N_5019);
nand U10248 (N_10248,N_9129,N_8417);
nand U10249 (N_10249,N_8263,N_8414);
and U10250 (N_10250,N_8541,N_8617);
or U10251 (N_10251,N_8251,N_5882);
or U10252 (N_10252,N_5620,N_5385);
nor U10253 (N_10253,N_7599,N_8932);
or U10254 (N_10254,N_8469,N_8477);
nand U10255 (N_10255,N_6060,N_7269);
nand U10256 (N_10256,N_9551,N_8457);
nand U10257 (N_10257,N_9441,N_9889);
nand U10258 (N_10258,N_6045,N_8871);
nor U10259 (N_10259,N_8476,N_9481);
nand U10260 (N_10260,N_7420,N_5586);
nand U10261 (N_10261,N_8458,N_5850);
and U10262 (N_10262,N_9322,N_9260);
nor U10263 (N_10263,N_5713,N_8426);
nand U10264 (N_10264,N_9918,N_5902);
and U10265 (N_10265,N_9221,N_6156);
nor U10266 (N_10266,N_7640,N_5275);
nand U10267 (N_10267,N_5821,N_6050);
or U10268 (N_10268,N_8354,N_8975);
or U10269 (N_10269,N_7233,N_8645);
nor U10270 (N_10270,N_6634,N_6822);
nand U10271 (N_10271,N_8915,N_5775);
nor U10272 (N_10272,N_9154,N_9489);
nor U10273 (N_10273,N_8503,N_8157);
and U10274 (N_10274,N_9747,N_8664);
or U10275 (N_10275,N_6399,N_9738);
nand U10276 (N_10276,N_8069,N_8172);
nor U10277 (N_10277,N_8140,N_7148);
nor U10278 (N_10278,N_5416,N_5812);
and U10279 (N_10279,N_6682,N_6210);
nor U10280 (N_10280,N_7659,N_9352);
nor U10281 (N_10281,N_8610,N_7188);
or U10282 (N_10282,N_9232,N_5118);
nor U10283 (N_10283,N_6228,N_9511);
or U10284 (N_10284,N_9610,N_8291);
nand U10285 (N_10285,N_8051,N_5110);
nor U10286 (N_10286,N_8917,N_7954);
nand U10287 (N_10287,N_7924,N_8399);
xor U10288 (N_10288,N_5351,N_6648);
nor U10289 (N_10289,N_9752,N_9576);
nor U10290 (N_10290,N_6931,N_8870);
nor U10291 (N_10291,N_7031,N_7965);
nor U10292 (N_10292,N_9740,N_5563);
nand U10293 (N_10293,N_9706,N_5521);
or U10294 (N_10294,N_6581,N_9288);
nand U10295 (N_10295,N_7860,N_5178);
nor U10296 (N_10296,N_5197,N_9193);
nand U10297 (N_10297,N_7214,N_6008);
nor U10298 (N_10298,N_6650,N_6107);
and U10299 (N_10299,N_5124,N_7627);
and U10300 (N_10300,N_6649,N_8092);
or U10301 (N_10301,N_9334,N_7828);
nor U10302 (N_10302,N_5513,N_8056);
nand U10303 (N_10303,N_7354,N_7282);
or U10304 (N_10304,N_5172,N_9472);
and U10305 (N_10305,N_5725,N_8000);
nor U10306 (N_10306,N_7105,N_9690);
and U10307 (N_10307,N_9432,N_7494);
nand U10308 (N_10308,N_7725,N_8694);
or U10309 (N_10309,N_5844,N_8789);
nor U10310 (N_10310,N_9795,N_8381);
nand U10311 (N_10311,N_7968,N_6478);
xor U10312 (N_10312,N_9843,N_6637);
xnor U10313 (N_10313,N_8619,N_6476);
xnor U10314 (N_10314,N_5909,N_6324);
xor U10315 (N_10315,N_5046,N_7534);
and U10316 (N_10316,N_8739,N_5645);
nor U10317 (N_10317,N_7816,N_9666);
nor U10318 (N_10318,N_7224,N_9981);
nor U10319 (N_10319,N_7763,N_6174);
nand U10320 (N_10320,N_8497,N_5627);
or U10321 (N_10321,N_6234,N_6609);
and U10322 (N_10322,N_9963,N_7794);
or U10323 (N_10323,N_7716,N_9537);
and U10324 (N_10324,N_9513,N_6527);
xor U10325 (N_10325,N_7140,N_6873);
or U10326 (N_10326,N_6004,N_7467);
nand U10327 (N_10327,N_8754,N_8266);
nor U10328 (N_10328,N_8712,N_8465);
nor U10329 (N_10329,N_6520,N_7159);
nor U10330 (N_10330,N_5634,N_9398);
nor U10331 (N_10331,N_6877,N_7062);
and U10332 (N_10332,N_6130,N_6926);
and U10333 (N_10333,N_5466,N_6773);
nand U10334 (N_10334,N_6145,N_5130);
xnor U10335 (N_10335,N_7088,N_5536);
and U10336 (N_10336,N_6495,N_7993);
and U10337 (N_10337,N_7096,N_7842);
nand U10338 (N_10338,N_6782,N_6279);
nor U10339 (N_10339,N_9825,N_8072);
nand U10340 (N_10340,N_7540,N_7000);
or U10341 (N_10341,N_7366,N_7518);
or U10342 (N_10342,N_7216,N_7682);
nand U10343 (N_10343,N_9282,N_6599);
nand U10344 (N_10344,N_9572,N_6487);
and U10345 (N_10345,N_6175,N_9568);
or U10346 (N_10346,N_6222,N_8081);
or U10347 (N_10347,N_8048,N_7799);
and U10348 (N_10348,N_8514,N_9350);
nand U10349 (N_10349,N_9406,N_5212);
or U10350 (N_10350,N_6452,N_7512);
or U10351 (N_10351,N_5260,N_9536);
nand U10352 (N_10352,N_9848,N_5234);
nand U10353 (N_10353,N_7417,N_8485);
or U10354 (N_10354,N_5073,N_9135);
or U10355 (N_10355,N_5204,N_6112);
or U10356 (N_10356,N_5831,N_8952);
and U10357 (N_10357,N_7803,N_7538);
or U10358 (N_10358,N_5992,N_8456);
or U10359 (N_10359,N_9806,N_5727);
and U10360 (N_10360,N_9830,N_7756);
or U10361 (N_10361,N_6031,N_6362);
nor U10362 (N_10362,N_8785,N_7026);
xor U10363 (N_10363,N_6680,N_9627);
or U10364 (N_10364,N_9371,N_9922);
nor U10365 (N_10365,N_9181,N_9040);
and U10366 (N_10366,N_9238,N_6412);
nand U10367 (N_10367,N_6236,N_6226);
and U10368 (N_10368,N_9418,N_8109);
nor U10369 (N_10369,N_5985,N_6765);
or U10370 (N_10370,N_5614,N_7436);
or U10371 (N_10371,N_6639,N_8379);
nor U10372 (N_10372,N_7598,N_8283);
xor U10373 (N_10373,N_6598,N_7781);
and U10374 (N_10374,N_9277,N_8918);
and U10375 (N_10375,N_8099,N_6786);
xor U10376 (N_10376,N_6217,N_5188);
and U10377 (N_10377,N_5300,N_5652);
nor U10378 (N_10378,N_8126,N_6020);
nor U10379 (N_10379,N_8779,N_6913);
nand U10380 (N_10380,N_8442,N_5191);
nor U10381 (N_10381,N_9957,N_8373);
nand U10382 (N_10382,N_5066,N_7531);
nor U10383 (N_10383,N_7744,N_9791);
nor U10384 (N_10384,N_7901,N_6778);
and U10385 (N_10385,N_5542,N_8067);
and U10386 (N_10386,N_7922,N_6098);
nor U10387 (N_10387,N_5241,N_9373);
and U10388 (N_10388,N_9296,N_6800);
or U10389 (N_10389,N_5607,N_9190);
and U10390 (N_10390,N_8974,N_7193);
or U10391 (N_10391,N_8096,N_6168);
or U10392 (N_10392,N_6705,N_8956);
and U10393 (N_10393,N_7112,N_5187);
and U10394 (N_10394,N_6759,N_7043);
and U10395 (N_10395,N_7620,N_5777);
xor U10396 (N_10396,N_7275,N_9681);
or U10397 (N_10397,N_8138,N_9546);
nand U10398 (N_10398,N_7453,N_5987);
nand U10399 (N_10399,N_6370,N_5742);
or U10400 (N_10400,N_5320,N_6240);
or U10401 (N_10401,N_5329,N_8627);
or U10402 (N_10402,N_9505,N_7445);
nor U10403 (N_10403,N_6295,N_6608);
and U10404 (N_10404,N_7299,N_6281);
or U10405 (N_10405,N_8210,N_7881);
nor U10406 (N_10406,N_5483,N_8490);
nand U10407 (N_10407,N_7495,N_7774);
or U10408 (N_10408,N_9257,N_8097);
nor U10409 (N_10409,N_5748,N_8348);
or U10410 (N_10410,N_5254,N_5084);
nor U10411 (N_10411,N_7448,N_9249);
or U10412 (N_10412,N_6561,N_8186);
nand U10413 (N_10413,N_5545,N_6310);
nand U10414 (N_10414,N_9941,N_7930);
or U10415 (N_10415,N_9695,N_5758);
nor U10416 (N_10416,N_9893,N_5383);
and U10417 (N_10417,N_5115,N_8219);
or U10418 (N_10418,N_7286,N_6938);
or U10419 (N_10419,N_5116,N_5892);
or U10420 (N_10420,N_7944,N_5451);
and U10421 (N_10421,N_9563,N_8362);
and U10422 (N_10422,N_5445,N_6933);
or U10423 (N_10423,N_8221,N_7374);
nand U10424 (N_10424,N_7578,N_9529);
or U10425 (N_10425,N_6468,N_8508);
nand U10426 (N_10426,N_7636,N_9920);
nand U10427 (N_10427,N_5668,N_5395);
and U10428 (N_10428,N_8162,N_7748);
nand U10429 (N_10429,N_5937,N_7894);
nor U10430 (N_10430,N_5905,N_9469);
or U10431 (N_10431,N_6923,N_5345);
nand U10432 (N_10432,N_8472,N_6285);
or U10433 (N_10433,N_8916,N_8833);
nor U10434 (N_10434,N_7812,N_9239);
nand U10435 (N_10435,N_5696,N_9256);
nor U10436 (N_10436,N_5272,N_8808);
xnor U10437 (N_10437,N_9330,N_7691);
nand U10438 (N_10438,N_6749,N_6342);
and U10439 (N_10439,N_8637,N_7848);
xor U10440 (N_10440,N_7325,N_9401);
or U10441 (N_10441,N_8933,N_7776);
nand U10442 (N_10442,N_8950,N_7411);
xnor U10443 (N_10443,N_9543,N_6594);
and U10444 (N_10444,N_9750,N_6988);
or U10445 (N_10445,N_9408,N_7482);
xnor U10446 (N_10446,N_7197,N_5421);
nor U10447 (N_10447,N_7007,N_6199);
and U10448 (N_10448,N_5891,N_8127);
and U10449 (N_10449,N_9134,N_9150);
or U10450 (N_10450,N_7029,N_5512);
and U10451 (N_10451,N_9411,N_5885);
and U10452 (N_10452,N_6806,N_5969);
nor U10453 (N_10453,N_9145,N_7442);
nand U10454 (N_10454,N_5447,N_6941);
or U10455 (N_10455,N_8095,N_6032);
nand U10456 (N_10456,N_7658,N_6667);
nor U10457 (N_10457,N_5145,N_5164);
and U10458 (N_10458,N_9746,N_8303);
nand U10459 (N_10459,N_7835,N_5315);
nand U10460 (N_10460,N_9852,N_6113);
and U10461 (N_10461,N_6805,N_5819);
nand U10462 (N_10462,N_8151,N_9119);
and U10463 (N_10463,N_9649,N_8707);
nand U10464 (N_10464,N_6436,N_9525);
xnor U10465 (N_10465,N_8315,N_9066);
nand U10466 (N_10466,N_5877,N_9633);
nor U10467 (N_10467,N_7050,N_5125);
and U10468 (N_10468,N_8977,N_7814);
and U10469 (N_10469,N_5367,N_8904);
and U10470 (N_10470,N_7479,N_5156);
and U10471 (N_10471,N_9586,N_5787);
nor U10472 (N_10472,N_9042,N_9314);
nand U10473 (N_10473,N_7859,N_5338);
nand U10474 (N_10474,N_6979,N_8703);
nor U10475 (N_10475,N_7223,N_7023);
nor U10476 (N_10476,N_8165,N_6652);
or U10477 (N_10477,N_7052,N_9850);
xnor U10478 (N_10478,N_5355,N_8715);
and U10479 (N_10479,N_5175,N_5822);
and U10480 (N_10480,N_5676,N_6027);
nor U10481 (N_10481,N_9044,N_9093);
or U10482 (N_10482,N_7301,N_9636);
nor U10483 (N_10483,N_9622,N_5883);
nor U10484 (N_10484,N_8632,N_7296);
xnor U10485 (N_10485,N_9015,N_8784);
and U10486 (N_10486,N_7372,N_5248);
nor U10487 (N_10487,N_9073,N_6431);
xor U10488 (N_10488,N_7095,N_6967);
nor U10489 (N_10489,N_8451,N_8108);
nor U10490 (N_10490,N_9547,N_7962);
or U10491 (N_10491,N_6698,N_7734);
nand U10492 (N_10492,N_5535,N_6335);
nor U10493 (N_10493,N_9026,N_9173);
nand U10494 (N_10494,N_5499,N_6319);
or U10495 (N_10495,N_6954,N_9253);
nand U10496 (N_10496,N_5051,N_5584);
nand U10497 (N_10497,N_6748,N_9443);
or U10498 (N_10498,N_7058,N_8749);
xnor U10499 (N_10499,N_6956,N_6983);
nand U10500 (N_10500,N_6492,N_9389);
or U10501 (N_10501,N_6225,N_8117);
nor U10502 (N_10502,N_7266,N_8187);
nor U10503 (N_10503,N_7369,N_6559);
nor U10504 (N_10504,N_9685,N_5550);
or U10505 (N_10505,N_5846,N_9088);
nor U10506 (N_10506,N_9022,N_8890);
nand U10507 (N_10507,N_9756,N_8846);
or U10508 (N_10508,N_8436,N_7612);
and U10509 (N_10509,N_8597,N_5043);
nor U10510 (N_10510,N_9766,N_5002);
nand U10511 (N_10511,N_5364,N_6920);
and U10512 (N_10512,N_5796,N_7483);
or U10513 (N_10513,N_7870,N_7946);
and U10514 (N_10514,N_8841,N_7068);
nand U10515 (N_10515,N_5838,N_9053);
xnor U10516 (N_10516,N_5836,N_9112);
xnor U10517 (N_10517,N_7869,N_6152);
nand U10518 (N_10518,N_6948,N_5113);
and U10519 (N_10519,N_7124,N_8836);
and U10520 (N_10520,N_6086,N_7335);
or U10521 (N_10521,N_6733,N_7942);
nor U10522 (N_10522,N_5808,N_5277);
or U10523 (N_10523,N_9030,N_8603);
and U10524 (N_10524,N_8606,N_7472);
and U10525 (N_10525,N_7185,N_8008);
nand U10526 (N_10526,N_9718,N_8775);
and U10527 (N_10527,N_5070,N_5310);
nand U10528 (N_10528,N_5702,N_9872);
xnor U10529 (N_10529,N_5765,N_6239);
nand U10530 (N_10530,N_7457,N_6897);
nor U10531 (N_10531,N_8111,N_7435);
nor U10532 (N_10532,N_5183,N_6407);
or U10533 (N_10533,N_8197,N_9544);
and U10534 (N_10534,N_6109,N_9209);
nand U10535 (N_10535,N_5694,N_7071);
or U10536 (N_10536,N_9315,N_5699);
nand U10537 (N_10537,N_5439,N_7852);
and U10538 (N_10538,N_9393,N_9989);
nor U10539 (N_10539,N_5538,N_6316);
or U10540 (N_10540,N_9211,N_7409);
or U10541 (N_10541,N_6246,N_6016);
and U10542 (N_10542,N_8188,N_9092);
and U10543 (N_10543,N_8049,N_8776);
or U10544 (N_10544,N_8230,N_9108);
or U10545 (N_10545,N_6939,N_8034);
and U10546 (N_10546,N_7378,N_6792);
and U10547 (N_10547,N_9477,N_7240);
and U10548 (N_10548,N_8207,N_7426);
nand U10549 (N_10549,N_9287,N_5406);
or U10550 (N_10550,N_9548,N_5829);
nor U10551 (N_10551,N_8036,N_5944);
and U10552 (N_10552,N_9560,N_8114);
nand U10553 (N_10553,N_8193,N_6816);
and U10554 (N_10554,N_7350,N_5497);
or U10555 (N_10555,N_8440,N_6015);
nand U10556 (N_10556,N_7826,N_5932);
nand U10557 (N_10557,N_9813,N_6424);
and U10558 (N_10558,N_6427,N_8286);
and U10559 (N_10559,N_7421,N_6219);
xnor U10560 (N_10560,N_6065,N_7796);
xor U10561 (N_10561,N_9975,N_6290);
and U10562 (N_10562,N_6182,N_6413);
and U10563 (N_10563,N_7441,N_5544);
nand U10564 (N_10564,N_9431,N_8488);
and U10565 (N_10565,N_5675,N_6908);
or U10566 (N_10566,N_7720,N_9733);
nor U10567 (N_10567,N_6361,N_5760);
xnor U10568 (N_10568,N_9117,N_5214);
or U10569 (N_10569,N_7403,N_6504);
or U10570 (N_10570,N_8448,N_8889);
and U10571 (N_10571,N_6591,N_7271);
or U10572 (N_10572,N_8175,N_9545);
nor U10573 (N_10573,N_8598,N_5967);
nor U10574 (N_10574,N_6013,N_7331);
or U10575 (N_10575,N_8329,N_5103);
and U10576 (N_10576,N_9087,N_6301);
and U10577 (N_10577,N_8983,N_9624);
and U10578 (N_10578,N_6916,N_6162);
nor U10579 (N_10579,N_9521,N_7678);
nor U10580 (N_10580,N_7918,N_8370);
xor U10581 (N_10581,N_6844,N_8256);
or U10582 (N_10582,N_5055,N_5163);
or U10583 (N_10583,N_8431,N_9413);
xnor U10584 (N_10584,N_5610,N_9799);
and U10585 (N_10585,N_6345,N_5721);
nand U10586 (N_10586,N_7017,N_5561);
or U10587 (N_10587,N_8960,N_7693);
or U10588 (N_10588,N_8681,N_9055);
and U10589 (N_10589,N_9344,N_7937);
nor U10590 (N_10590,N_5824,N_8103);
nand U10591 (N_10591,N_7294,N_5456);
nor U10592 (N_10592,N_7865,N_8146);
or U10593 (N_10593,N_8234,N_8912);
or U10594 (N_10594,N_8406,N_9671);
and U10595 (N_10595,N_9687,N_7570);
or U10596 (N_10596,N_9812,N_5624);
xnor U10597 (N_10597,N_5865,N_5250);
nor U10598 (N_10598,N_6915,N_8304);
or U10599 (N_10599,N_6590,N_5480);
nor U10600 (N_10600,N_8757,N_8729);
nand U10601 (N_10601,N_6975,N_9235);
nand U10602 (N_10602,N_6953,N_8564);
and U10603 (N_10603,N_8920,N_7897);
or U10604 (N_10604,N_8392,N_6853);
or U10605 (N_10605,N_5419,N_6397);
and U10606 (N_10606,N_8418,N_6091);
nand U10607 (N_10607,N_9721,N_8942);
nor U10608 (N_10608,N_9914,N_7175);
nor U10609 (N_10609,N_6356,N_8317);
nor U10610 (N_10610,N_6393,N_5446);
and U10611 (N_10611,N_9534,N_8859);
nand U10612 (N_10612,N_8604,N_5593);
nand U10613 (N_10613,N_5346,N_5626);
xor U10614 (N_10614,N_8809,N_5647);
xor U10615 (N_10615,N_8685,N_6218);
nor U10616 (N_10616,N_8131,N_5640);
nand U10617 (N_10617,N_7569,N_7559);
and U10618 (N_10618,N_6149,N_9735);
nor U10619 (N_10619,N_7502,N_7415);
nand U10620 (N_10620,N_6820,N_6535);
and U10621 (N_10621,N_9306,N_9065);
or U10622 (N_10622,N_8142,N_5598);
or U10623 (N_10623,N_9180,N_9785);
nor U10624 (N_10624,N_6318,N_5943);
or U10625 (N_10625,N_9264,N_7360);
or U10626 (N_10626,N_9767,N_9337);
nand U10627 (N_10627,N_7137,N_5653);
nor U10628 (N_10628,N_5531,N_9363);
nor U10629 (N_10629,N_7365,N_6284);
and U10630 (N_10630,N_5737,N_5734);
xnor U10631 (N_10631,N_9156,N_5484);
nand U10632 (N_10632,N_7487,N_6815);
xnor U10633 (N_10633,N_5566,N_6633);
nor U10634 (N_10634,N_5915,N_5236);
and U10635 (N_10635,N_6871,N_5599);
or U10636 (N_10636,N_9926,N_9212);
nand U10637 (N_10637,N_8523,N_7257);
nand U10638 (N_10638,N_5437,N_7202);
nand U10639 (N_10639,N_8492,N_6242);
and U10640 (N_10640,N_7926,N_7972);
and U10641 (N_10641,N_7357,N_9580);
or U10642 (N_10642,N_5712,N_5855);
nor U10643 (N_10643,N_8850,N_7134);
nand U10644 (N_10644,N_6885,N_9272);
nand U10645 (N_10645,N_8385,N_9585);
xnor U10646 (N_10646,N_8330,N_7337);
nand U10647 (N_10647,N_9298,N_9038);
nor U10648 (N_10648,N_6809,N_6902);
nand U10649 (N_10649,N_6213,N_6617);
or U10650 (N_10650,N_6110,N_5293);
nor U10651 (N_10651,N_8184,N_7769);
or U10652 (N_10652,N_8257,N_5528);
or U10653 (N_10653,N_9278,N_8085);
nor U10654 (N_10654,N_7652,N_6552);
and U10655 (N_10655,N_8802,N_9276);
and U10656 (N_10656,N_6325,N_7742);
and U10657 (N_10657,N_8946,N_7561);
or U10658 (N_10658,N_5710,N_8825);
nor U10659 (N_10659,N_5785,N_9762);
or U10660 (N_10660,N_6847,N_7144);
and U10661 (N_10661,N_7861,N_5641);
and U10662 (N_10662,N_5973,N_6973);
or U10663 (N_10663,N_7098,N_9930);
xnor U10664 (N_10664,N_7955,N_6303);
xor U10665 (N_10665,N_9050,N_8643);
nand U10666 (N_10666,N_8571,N_7949);
nor U10667 (N_10667,N_5674,N_8282);
or U10668 (N_10668,N_8579,N_6494);
nand U10669 (N_10669,N_7451,N_7862);
nor U10670 (N_10670,N_6408,N_6101);
xnor U10671 (N_10671,N_8427,N_9532);
nor U10672 (N_10672,N_5302,N_6959);
nor U10673 (N_10673,N_6305,N_6958);
nand U10674 (N_10674,N_7880,N_5866);
nand U10675 (N_10675,N_9381,N_8355);
or U10676 (N_10676,N_5011,N_9683);
and U10677 (N_10677,N_5928,N_6061);
or U10678 (N_10678,N_8813,N_5749);
nand U10679 (N_10679,N_8017,N_6982);
nand U10680 (N_10680,N_6542,N_7895);
xnor U10681 (N_10681,N_5035,N_9188);
nand U10682 (N_10682,N_5874,N_5815);
xor U10683 (N_10683,N_7992,N_6072);
nand U10684 (N_10684,N_8745,N_6111);
nor U10685 (N_10685,N_8424,N_6057);
or U10686 (N_10686,N_7733,N_7710);
nor U10687 (N_10687,N_9400,N_5273);
nor U10688 (N_10688,N_5403,N_7511);
nor U10689 (N_10689,N_8154,N_6510);
and U10690 (N_10690,N_6169,N_6878);
nand U10691 (N_10691,N_8387,N_8868);
and U10692 (N_10692,N_8409,N_5703);
and U10693 (N_10693,N_6433,N_5658);
and U10694 (N_10694,N_7241,N_7908);
nor U10695 (N_10695,N_5038,N_7999);
and U10696 (N_10696,N_6106,N_9320);
nand U10697 (N_10697,N_7751,N_5763);
or U10698 (N_10698,N_6313,N_7455);
nand U10699 (N_10699,N_8402,N_9510);
nor U10700 (N_10700,N_9895,N_8517);
nor U10701 (N_10701,N_8894,N_7705);
and U10702 (N_10702,N_7632,N_8677);
nand U10703 (N_10703,N_7093,N_6977);
or U10704 (N_10704,N_6692,N_7800);
and U10705 (N_10705,N_9814,N_6512);
nor U10706 (N_10706,N_5478,N_7295);
nor U10707 (N_10707,N_5148,N_6766);
nand U10708 (N_10708,N_9316,N_6819);
or U10709 (N_10709,N_6825,N_5223);
and U10710 (N_10710,N_9482,N_9996);
and U10711 (N_10711,N_8041,N_7513);
nand U10712 (N_10712,N_8687,N_6223);
xnor U10713 (N_10713,N_5618,N_9291);
or U10714 (N_10714,N_6767,N_8542);
nor U10715 (N_10715,N_6569,N_7832);
xor U10716 (N_10716,N_5102,N_9940);
nor U10717 (N_10717,N_5660,N_5380);
nand U10718 (N_10718,N_9429,N_6636);
and U10719 (N_10719,N_7581,N_7272);
and U10720 (N_10720,N_6723,N_5266);
nand U10721 (N_10721,N_5503,N_8396);
nand U10722 (N_10722,N_7264,N_9455);
nand U10723 (N_10723,N_8148,N_7522);
nor U10724 (N_10724,N_8196,N_9360);
or U10725 (N_10725,N_5424,N_9097);
nor U10726 (N_10726,N_6321,N_9052);
xnor U10727 (N_10727,N_7145,N_8909);
xor U10728 (N_10728,N_5683,N_9280);
nor U10729 (N_10729,N_5889,N_8130);
nand U10730 (N_10730,N_9621,N_9628);
and U10731 (N_10731,N_7960,N_5348);
and U10732 (N_10732,N_8861,N_7997);
or U10733 (N_10733,N_8887,N_9116);
nand U10734 (N_10734,N_6038,N_6482);
nor U10735 (N_10735,N_6205,N_9881);
and U10736 (N_10736,N_9883,N_8369);
xor U10737 (N_10737,N_7229,N_5311);
or U10738 (N_10738,N_9915,N_9967);
and U10739 (N_10739,N_8589,N_5012);
nand U10740 (N_10740,N_9458,N_6062);
and U10741 (N_10741,N_8957,N_8389);
nor U10742 (N_10742,N_8149,N_6570);
or U10743 (N_10743,N_6677,N_6126);
xnor U10744 (N_10744,N_7662,N_8420);
nor U10745 (N_10745,N_6862,N_8336);
nor U10746 (N_10746,N_9480,N_9686);
nor U10747 (N_10747,N_9680,N_9728);
and U10748 (N_10748,N_5568,N_7065);
nand U10749 (N_10749,N_7130,N_9255);
nand U10750 (N_10750,N_8124,N_9639);
nor U10751 (N_10751,N_9754,N_9017);
and U10752 (N_10752,N_5195,N_5041);
nand U10753 (N_10753,N_8218,N_9072);
nand U10754 (N_10754,N_9907,N_8863);
and U10755 (N_10755,N_9980,N_8482);
and U10756 (N_10756,N_8762,N_9057);
nor U10757 (N_10757,N_9910,N_8278);
or U10758 (N_10758,N_9974,N_6750);
nor U10759 (N_10759,N_7934,N_7136);
xnor U10760 (N_10760,N_8856,N_8596);
nor U10761 (N_10761,N_6893,N_5856);
nand U10762 (N_10762,N_7187,N_7126);
or U10763 (N_10763,N_7625,N_5114);
nand U10764 (N_10764,N_7873,N_7753);
and U10765 (N_10765,N_7558,N_8591);
nand U10766 (N_10766,N_5292,N_8308);
or U10767 (N_10767,N_9892,N_6186);
nor U10768 (N_10768,N_5034,N_7253);
nor U10769 (N_10769,N_8997,N_7437);
nand U10770 (N_10770,N_5628,N_7277);
xnor U10771 (N_10771,N_7317,N_8121);
xnor U10772 (N_10772,N_6999,N_5050);
nor U10773 (N_10773,N_6836,N_7080);
nor U10774 (N_10774,N_7545,N_8631);
xor U10775 (N_10775,N_7533,N_5518);
xnor U10776 (N_10776,N_7508,N_9001);
or U10777 (N_10777,N_6344,N_5644);
nor U10778 (N_10778,N_9332,N_5230);
and U10779 (N_10779,N_5826,N_7290);
nor U10780 (N_10780,N_6712,N_6037);
nand U10781 (N_10781,N_5585,N_5376);
nand U10782 (N_10782,N_5622,N_7027);
or U10783 (N_10783,N_5386,N_6589);
and U10784 (N_10784,N_8446,N_6464);
and U10785 (N_10785,N_7650,N_6661);
nand U10786 (N_10786,N_7276,N_8936);
or U10787 (N_10787,N_5520,N_6466);
nand U10788 (N_10788,N_8029,N_8119);
xor U10789 (N_10789,N_9908,N_8011);
nor U10790 (N_10790,N_8873,N_6483);
or U10791 (N_10791,N_9853,N_7963);
nor U10792 (N_10792,N_6780,N_5952);
and U10793 (N_10793,N_5401,N_5506);
nand U10794 (N_10794,N_6968,N_9415);
nand U10795 (N_10795,N_5921,N_8788);
nand U10796 (N_10796,N_8449,N_9928);
and U10797 (N_10797,N_7142,N_8882);
and U10798 (N_10798,N_5284,N_9076);
and U10799 (N_10799,N_5502,N_7478);
or U10800 (N_10800,N_6178,N_8268);
nor U10801 (N_10801,N_9579,N_5840);
or U10802 (N_10802,N_7076,N_9933);
or U10803 (N_10803,N_5695,N_6010);
or U10804 (N_10804,N_5739,N_7583);
or U10805 (N_10805,N_9761,N_5793);
nor U10806 (N_10806,N_6621,N_8147);
and U10807 (N_10807,N_8122,N_8710);
nor U10808 (N_10808,N_8515,N_7986);
nand U10809 (N_10809,N_9869,N_7864);
or U10810 (N_10810,N_5930,N_5807);
nor U10811 (N_10811,N_8239,N_6124);
and U10812 (N_10812,N_9358,N_9644);
nand U10813 (N_10813,N_8520,N_7094);
or U10814 (N_10814,N_6443,N_8258);
and U10815 (N_10815,N_8580,N_7623);
xnor U10816 (N_10816,N_5537,N_9008);
nor U10817 (N_10817,N_5228,N_8824);
and U10818 (N_10818,N_7067,N_7673);
nand U10819 (N_10819,N_8756,N_9661);
nor U10820 (N_10820,N_7586,N_5294);
nand U10821 (N_10821,N_5825,N_7576);
and U10822 (N_10822,N_8867,N_7447);
nand U10823 (N_10823,N_8507,N_5256);
and U10824 (N_10824,N_5895,N_8073);
nor U10825 (N_10825,N_7582,N_8214);
nor U10826 (N_10826,N_5473,N_5576);
nor U10827 (N_10827,N_9394,N_6752);
nor U10828 (N_10828,N_6409,N_7634);
or U10829 (N_10829,N_8419,N_6329);
nand U10830 (N_10830,N_5301,N_8650);
nor U10831 (N_10831,N_7305,N_5245);
nor U10832 (N_10832,N_5509,N_6818);
xor U10833 (N_10833,N_7444,N_5425);
or U10834 (N_10834,N_9873,N_7133);
nor U10835 (N_10835,N_7490,N_6935);
nor U10836 (N_10836,N_6103,N_6432);
or U10837 (N_10837,N_9798,N_6627);
nand U10838 (N_10838,N_7206,N_8141);
and U10839 (N_10839,N_5015,N_9345);
nor U10840 (N_10840,N_6644,N_8649);
xor U10841 (N_10841,N_8992,N_6663);
or U10842 (N_10842,N_7994,N_6914);
and U10843 (N_10843,N_9024,N_8031);
or U10844 (N_10844,N_7849,N_5574);
and U10845 (N_10845,N_9056,N_8896);
and U10846 (N_10846,N_7111,N_7303);
nand U10847 (N_10847,N_8053,N_8796);
nor U10848 (N_10848,N_8435,N_8374);
nor U10849 (N_10849,N_6009,N_6622);
or U10850 (N_10850,N_9899,N_8881);
nor U10851 (N_10851,N_9707,N_5373);
xnor U10852 (N_10852,N_8352,N_5396);
nor U10853 (N_10853,N_9998,N_6777);
and U10854 (N_10854,N_8322,N_9473);
or U10855 (N_10855,N_6568,N_8015);
or U10856 (N_10856,N_8013,N_8990);
nand U10857 (N_10857,N_7073,N_6866);
nor U10858 (N_10858,N_5601,N_8245);
nand U10859 (N_10859,N_6539,N_9230);
and U10860 (N_10860,N_8460,N_9279);
nand U10861 (N_10861,N_5279,N_8057);
and U10862 (N_10862,N_9939,N_5978);
xnor U10863 (N_10863,N_6689,N_5633);
nor U10864 (N_10864,N_7297,N_8176);
or U10865 (N_10865,N_9107,N_9748);
nand U10866 (N_10866,N_7425,N_8506);
nand U10867 (N_10867,N_7855,N_5475);
xnor U10868 (N_10868,N_6254,N_9715);
xnor U10869 (N_10869,N_5201,N_6401);
or U10870 (N_10870,N_5107,N_6580);
nand U10871 (N_10871,N_5917,N_7389);
and U10872 (N_10872,N_9629,N_5233);
or U10873 (N_10873,N_6267,N_8252);
nor U10874 (N_10874,N_9901,N_8624);
or U10875 (N_10875,N_8408,N_7030);
or U10876 (N_10876,N_7683,N_7450);
and U10877 (N_10877,N_6709,N_9711);
nand U10878 (N_10878,N_5625,N_6700);
and U10879 (N_10879,N_6554,N_9157);
and U10880 (N_10880,N_7011,N_5352);
or U10881 (N_10881,N_8213,N_5288);
and U10882 (N_10882,N_9719,N_5290);
nand U10883 (N_10883,N_5768,N_5109);
nand U10884 (N_10884,N_8875,N_7474);
and U10885 (N_10885,N_8864,N_9526);
or U10886 (N_10886,N_7764,N_8660);
and U10887 (N_10887,N_9166,N_6874);
nand U10888 (N_10888,N_9720,N_5693);
and U10889 (N_10889,N_5074,N_5328);
nand U10890 (N_10890,N_8862,N_9626);
or U10891 (N_10891,N_9089,N_8700);
and U10892 (N_10892,N_7746,N_7419);
nand U10893 (N_10893,N_9353,N_6787);
or U10894 (N_10894,N_8331,N_5604);
or U10895 (N_10895,N_6249,N_5122);
and U10896 (N_10896,N_8452,N_5871);
xor U10897 (N_10897,N_6251,N_6593);
or U10898 (N_10898,N_6421,N_8068);
and U10899 (N_10899,N_8616,N_7544);
and U10900 (N_10900,N_6934,N_8307);
nor U10901 (N_10901,N_8074,N_5166);
and U10902 (N_10902,N_8722,N_9946);
nand U10903 (N_10903,N_5339,N_6994);
or U10904 (N_10904,N_7370,N_9290);
nor U10905 (N_10905,N_7334,N_7856);
and U10906 (N_10906,N_5121,N_5654);
or U10907 (N_10907,N_9938,N_6270);
or U10908 (N_10908,N_8112,N_8538);
and U10909 (N_10909,N_7351,N_9109);
nand U10910 (N_10910,N_9607,N_7209);
nor U10911 (N_10911,N_7975,N_6348);
nor U10912 (N_10912,N_6276,N_6189);
and U10913 (N_10913,N_9772,N_8927);
nand U10914 (N_10914,N_5318,N_6696);
and U10915 (N_10915,N_9223,N_6006);
and U10916 (N_10916,N_8024,N_9460);
nor U10917 (N_10917,N_6144,N_6312);
nand U10918 (N_10918,N_8269,N_5716);
nor U10919 (N_10919,N_7243,N_7190);
and U10920 (N_10920,N_6503,N_8346);
or U10921 (N_10921,N_7898,N_8982);
or U10922 (N_10922,N_6585,N_8979);
nor U10923 (N_10923,N_9159,N_8390);
xnor U10924 (N_10924,N_7249,N_6950);
nor U10925 (N_10925,N_8075,N_9783);
nand U10926 (N_10926,N_5472,N_7567);
nand U10927 (N_10927,N_7407,N_7817);
nor U10928 (N_10928,N_8483,N_7740);
and U10929 (N_10929,N_6772,N_7427);
xor U10930 (N_10930,N_8470,N_9823);
nor U10931 (N_10931,N_6925,N_8748);
nor U10932 (N_10932,N_7767,N_6620);
nand U10933 (N_10933,N_5820,N_9491);
nor U10934 (N_10934,N_8852,N_5149);
and U10935 (N_10935,N_7853,N_9755);
nand U10936 (N_10936,N_5786,N_8403);
or U10937 (N_10937,N_6350,N_5024);
and U10938 (N_10938,N_8988,N_7438);
nor U10939 (N_10939,N_5705,N_8164);
nor U10940 (N_10940,N_6564,N_6085);
nor U10941 (N_10941,N_6525,N_6490);
nand U10942 (N_10942,N_5738,N_9171);
and U10943 (N_10943,N_5872,N_9642);
and U10944 (N_10944,N_9659,N_8574);
nor U10945 (N_10945,N_5929,N_8367);
nand U10946 (N_10946,N_7738,N_7863);
or U10947 (N_10947,N_8924,N_5258);
nand U10948 (N_10948,N_9247,N_5851);
or U10949 (N_10949,N_8201,N_8782);
or U10950 (N_10950,N_6012,N_9535);
and U10951 (N_10951,N_8377,N_8530);
and U10952 (N_10952,N_8495,N_5366);
nor U10953 (N_10953,N_9437,N_6522);
nor U10954 (N_10954,N_9148,N_9189);
nor U10955 (N_10955,N_7379,N_9452);
and U10956 (N_10956,N_5182,N_8937);
nor U10957 (N_10957,N_6596,N_7183);
and U10958 (N_10958,N_9541,N_9542);
or U10959 (N_10959,N_6952,N_6976);
nand U10960 (N_10960,N_9376,N_8962);
or U10961 (N_10961,N_6514,N_8609);
or U10962 (N_10962,N_5590,N_8641);
nand U10963 (N_10963,N_8265,N_9522);
xor U10964 (N_10964,N_6775,N_6224);
nand U10965 (N_10965,N_5308,N_9595);
or U10966 (N_10966,N_7726,N_5799);
or U10967 (N_10967,N_5570,N_6789);
and U10968 (N_10968,N_6030,N_7952);
nand U10969 (N_10969,N_9838,N_5539);
and U10970 (N_10970,N_8270,N_5975);
nand U10971 (N_10971,N_9465,N_6586);
nor U10972 (N_10972,N_7072,N_5219);
nor U10973 (N_10973,N_5261,N_7217);
nand U10974 (N_10974,N_8973,N_5578);
or U10975 (N_10975,N_8718,N_8584);
nor U10976 (N_10976,N_8587,N_7602);
or U10977 (N_10977,N_8338,N_7989);
and U10978 (N_10978,N_6460,N_5525);
nand U10979 (N_10979,N_9500,N_6894);
or U10980 (N_10980,N_7117,N_7815);
nor U10981 (N_10981,N_5504,N_8527);
or U10982 (N_10982,N_7923,N_7681);
and U10983 (N_10983,N_6209,N_9688);
xor U10984 (N_10984,N_9139,N_6383);
xor U10985 (N_10985,N_8395,N_5782);
xor U10986 (N_10986,N_8851,N_6491);
and U10987 (N_10987,N_6379,N_7684);
nor U10988 (N_10988,N_9999,N_8673);
or U10989 (N_10989,N_6364,N_5285);
or U10990 (N_10990,N_6674,N_6995);
or U10991 (N_10991,N_9790,N_5996);
xnor U10992 (N_10992,N_9297,N_9667);
or U10993 (N_10993,N_6887,N_8552);
xor U10994 (N_10994,N_9722,N_6769);
nor U10995 (N_10995,N_7891,N_8116);
and U10996 (N_10996,N_8804,N_6742);
and U10997 (N_10997,N_5977,N_5143);
or U10998 (N_10998,N_6007,N_6718);
and U10999 (N_10999,N_7408,N_5463);
xor U11000 (N_11000,N_8522,N_9768);
nand U11001 (N_11001,N_9078,N_6069);
nand U11002 (N_11002,N_6615,N_9149);
or U11003 (N_11003,N_8935,N_7182);
and U11004 (N_11004,N_9357,N_9777);
nor U11005 (N_11005,N_7951,N_5269);
and U11006 (N_11006,N_8335,N_7584);
nand U11007 (N_11007,N_6376,N_5778);
xnor U11008 (N_11008,N_6670,N_7822);
or U11009 (N_11009,N_8088,N_6732);
xnor U11010 (N_11010,N_6903,N_7128);
nor U11011 (N_11011,N_6830,N_9111);
or U11012 (N_11012,N_9835,N_5132);
and U11013 (N_11013,N_9829,N_7592);
and U11014 (N_11014,N_6089,N_9133);
nor U11015 (N_11015,N_5264,N_5448);
nor U11016 (N_11016,N_6823,N_9849);
and U11017 (N_11017,N_6841,N_7637);
or U11018 (N_11018,N_9792,N_8222);
or U11019 (N_11019,N_9549,N_6888);
and U11020 (N_11020,N_6457,N_5592);
and U11021 (N_11021,N_7056,N_8365);
and U11022 (N_11022,N_9479,N_9906);
and U11023 (N_11023,N_6861,N_6707);
nor U11024 (N_11024,N_5363,N_6115);
nand U11025 (N_11025,N_6040,N_7491);
and U11026 (N_11026,N_8978,N_9932);
xor U11027 (N_11027,N_7377,N_7324);
nor U11028 (N_11028,N_8670,N_7347);
and U11029 (N_11029,N_7336,N_5001);
nand U11030 (N_11030,N_8736,N_6839);
xor U11031 (N_11031,N_9739,N_9004);
nand U11032 (N_11032,N_6461,N_9828);
and U11033 (N_11033,N_6991,N_7996);
nor U11034 (N_11034,N_8101,N_8967);
nor U11035 (N_11035,N_7793,N_5211);
nor U11036 (N_11036,N_5630,N_7896);
nand U11037 (N_11037,N_9882,N_6351);
xnor U11038 (N_11038,N_6611,N_8858);
or U11039 (N_11039,N_5827,N_7866);
nor U11040 (N_11040,N_9421,N_7900);
or U11041 (N_11041,N_5956,N_9266);
and U11042 (N_11042,N_6971,N_5546);
nor U11043 (N_11043,N_9403,N_9144);
nor U11044 (N_11044,N_5764,N_9311);
and U11045 (N_11045,N_5690,N_6811);
nand U11046 (N_11046,N_8572,N_7613);
or U11047 (N_11047,N_7412,N_8086);
nor U11048 (N_11048,N_8500,N_7739);
nor U11049 (N_11049,N_6024,N_5108);
or U11050 (N_11050,N_5434,N_8473);
and U11051 (N_11051,N_8646,N_8227);
or U11052 (N_11052,N_6034,N_9951);
and U11053 (N_11053,N_6704,N_8753);
or U11054 (N_11054,N_5170,N_8595);
nand U11055 (N_11055,N_6258,N_5524);
or U11056 (N_11056,N_5274,N_9450);
or U11057 (N_11057,N_7687,N_8787);
or U11058 (N_11058,N_6567,N_6602);
nand U11059 (N_11059,N_5072,N_8380);
xor U11060 (N_11060,N_9888,N_6244);
and U11061 (N_11061,N_7476,N_7001);
nand U11062 (N_11062,N_8501,N_6694);
or U11063 (N_11063,N_9170,N_9486);
and U11064 (N_11064,N_9966,N_7646);
nand U11065 (N_11065,N_5839,N_8620);
or U11066 (N_11066,N_8394,N_9655);
or U11067 (N_11067,N_8512,N_8696);
nand U11068 (N_11068,N_6440,N_6282);
or U11069 (N_11069,N_5527,N_6428);
or U11070 (N_11070,N_5670,N_5876);
or U11071 (N_11071,N_7760,N_8038);
and U11072 (N_11072,N_5964,N_8719);
nor U11073 (N_11073,N_8888,N_5863);
and U11074 (N_11074,N_8177,N_7956);
nand U11075 (N_11075,N_8475,N_6268);
or U11076 (N_11076,N_5792,N_6889);
nand U11077 (N_11077,N_5237,N_9652);
and U11078 (N_11078,N_7025,N_8524);
xor U11079 (N_11079,N_8714,N_5920);
or U11080 (N_11080,N_5423,N_6087);
nand U11081 (N_11081,N_9726,N_5903);
or U11082 (N_11082,N_8908,N_5078);
nand U11083 (N_11083,N_8136,N_6932);
nor U11084 (N_11084,N_6484,N_9043);
nor U11085 (N_11085,N_6451,N_8683);
nor U11086 (N_11086,N_5854,N_7831);
nor U11087 (N_11087,N_8525,N_8318);
or U11088 (N_11088,N_8519,N_9234);
nand U11089 (N_11089,N_9242,N_5408);
and U11090 (N_11090,N_6505,N_6201);
nor U11091 (N_11091,N_5246,N_8450);
nand U11092 (N_11092,N_7893,N_5832);
or U11093 (N_11093,N_8020,N_8319);
and U11094 (N_11094,N_8016,N_6266);
nand U11095 (N_11095,N_7053,N_5493);
nand U11096 (N_11096,N_6048,N_5998);
xnor U11097 (N_11097,N_9840,N_7547);
or U11098 (N_11098,N_5065,N_5776);
nor U11099 (N_11099,N_5752,N_5136);
or U11100 (N_11100,N_7504,N_5534);
xnor U11101 (N_11101,N_8076,N_5714);
and U11102 (N_11102,N_6537,N_6341);
and U11103 (N_11103,N_7003,N_5006);
xor U11104 (N_11104,N_5887,N_6533);
or U11105 (N_11105,N_7615,N_6423);
or U11106 (N_11106,N_7122,N_5005);
nand U11107 (N_11107,N_8573,N_8298);
nand U11108 (N_11108,N_7843,N_9416);
and U11109 (N_11109,N_6797,N_5128);
nor U11110 (N_11110,N_9131,N_5818);
xor U11111 (N_11111,N_5723,N_6645);
or U11112 (N_11112,N_8383,N_6448);
or U11113 (N_11113,N_8012,N_8104);
or U11114 (N_11114,N_9202,N_7782);
nand U11115 (N_11115,N_8563,N_5802);
and U11116 (N_11116,N_7785,N_9776);
nor U11117 (N_11117,N_9196,N_9395);
or U11118 (N_11118,N_9731,N_6669);
and U11119 (N_11119,N_5719,N_5021);
or U11120 (N_11120,N_5789,N_9200);
nor U11121 (N_11121,N_5220,N_7819);
nand U11122 (N_11122,N_9122,N_6190);
and U11123 (N_11123,N_6990,N_7916);
and U11124 (N_11124,N_8855,N_8518);
or U11125 (N_11125,N_6758,N_6299);
nand U11126 (N_11126,N_7138,N_5185);
and U11127 (N_11127,N_8332,N_6386);
and U11128 (N_11128,N_5282,N_7605);
and U11129 (N_11129,N_9047,N_7218);
and U11130 (N_11130,N_8468,N_6890);
nor U11131 (N_11131,N_8544,N_7980);
xnor U11132 (N_11132,N_5461,N_5817);
or U11133 (N_11133,N_9318,N_8903);
or U11134 (N_11134,N_6578,N_5837);
nor U11135 (N_11135,N_6181,N_9435);
and U11136 (N_11136,N_8865,N_8158);
and U11137 (N_11137,N_7609,N_8951);
nor U11138 (N_11138,N_9302,N_7727);
xnor U11139 (N_11139,N_7899,N_9348);
or U11140 (N_11140,N_9531,N_8895);
nand U11141 (N_11141,N_5390,N_7787);
or U11142 (N_11142,N_7353,N_6702);
or U11143 (N_11143,N_7614,N_9404);
and U11144 (N_11144,N_5023,N_8433);
and U11145 (N_11145,N_8447,N_7012);
or U11146 (N_11146,N_7837,N_5988);
nand U11147 (N_11147,N_6055,N_7698);
and U11148 (N_11148,N_6355,N_7220);
and U11149 (N_11149,N_7367,N_7985);
or U11150 (N_11150,N_7798,N_9675);
nor U11151 (N_11151,N_8945,N_8287);
xnor U11152 (N_11152,N_6746,N_8893);
nand U11153 (N_11153,N_9466,N_6676);
xnor U11154 (N_11154,N_7840,N_9308);
and U11155 (N_11155,N_8582,N_6523);
and U11156 (N_11156,N_7821,N_7464);
xor U11157 (N_11157,N_8125,N_9059);
and U11158 (N_11158,N_9152,N_7530);
nand U11159 (N_11159,N_9917,N_9137);
or U11160 (N_11160,N_9818,N_5229);
nor U11161 (N_11161,N_5553,N_5514);
nor U11162 (N_11162,N_6136,N_9143);
and U11163 (N_11163,N_6296,N_7752);
or U11164 (N_11164,N_8778,N_5631);
or U11165 (N_11165,N_5770,N_7265);
and U11166 (N_11166,N_8549,N_7070);
and U11167 (N_11167,N_5435,N_5811);
nand U11168 (N_11168,N_7207,N_9051);
nor U11169 (N_11169,N_8658,N_7663);
xor U11170 (N_11170,N_8084,N_6259);
or U11171 (N_11171,N_5319,N_7373);
and U11172 (N_11172,N_9385,N_7797);
nand U11173 (N_11173,N_5359,N_9114);
nor U11174 (N_11174,N_5881,N_8551);
nand U11175 (N_11175,N_9589,N_8249);
and U11176 (N_11176,N_8260,N_9494);
nand U11177 (N_11177,N_8566,N_9617);
and U11178 (N_11178,N_5147,N_7416);
and U11179 (N_11179,N_9630,N_8055);
nor U11180 (N_11180,N_8625,N_8173);
xnor U11181 (N_11181,N_6003,N_9986);
nand U11182 (N_11182,N_7018,N_9968);
nor U11183 (N_11183,N_7889,N_5979);
nand U11184 (N_11184,N_7622,N_5176);
xnor U11185 (N_11185,N_5327,N_9034);
nand U11186 (N_11186,N_8554,N_6868);
and U11187 (N_11187,N_5587,N_6571);
or U11188 (N_11188,N_5045,N_8054);
and U11189 (N_11189,N_8963,N_8815);
or U11190 (N_11190,N_5389,N_8689);
nand U11191 (N_11191,N_8052,N_7180);
and U11192 (N_11192,N_9128,N_5086);
nand U11193 (N_11193,N_9265,N_5688);
xnor U11194 (N_11194,N_7695,N_6148);
xor U11195 (N_11195,N_5666,N_8397);
nand U11196 (N_11196,N_7368,N_6684);
nor U11197 (N_11197,N_7439,N_8623);
or U11198 (N_11198,N_7086,N_7905);
nand U11199 (N_11199,N_8926,N_6653);
nand U11200 (N_11200,N_5381,N_8832);
and U11201 (N_11201,N_7260,N_6159);
xnor U11202 (N_11202,N_6090,N_5180);
and U11203 (N_11203,N_6628,N_9365);
and U11204 (N_11204,N_6135,N_9424);
or U11205 (N_11205,N_8910,N_5347);
or U11206 (N_11206,N_7621,N_9786);
nand U11207 (N_11207,N_7259,N_7168);
and U11208 (N_11208,N_5961,N_8630);
nand U11209 (N_11209,N_8244,N_8079);
and U11210 (N_11210,N_7600,N_5784);
nor U11211 (N_11211,N_9590,N_7227);
nand U11212 (N_11212,N_6557,N_5867);
nor U11213 (N_11213,N_8285,N_6831);
nor U11214 (N_11214,N_6185,N_8356);
or U11215 (N_11215,N_5462,N_6619);
or U11216 (N_11216,N_9328,N_7035);
or U11217 (N_11217,N_9801,N_7315);
nor U11218 (N_11218,N_7730,N_9887);
and U11219 (N_11219,N_5697,N_7712);
or U11220 (N_11220,N_7885,N_9507);
or U11221 (N_11221,N_8536,N_7388);
or U11222 (N_11222,N_7928,N_6638);
nor U11223 (N_11223,N_5374,N_9760);
nor U11224 (N_11224,N_6366,N_9061);
or U11225 (N_11225,N_8772,N_9912);
nand U11226 (N_11226,N_7151,N_5217);
nand U11227 (N_11227,N_8969,N_8531);
and U11228 (N_11228,N_5646,N_9861);
nor U11229 (N_11229,N_8532,N_8793);
and U11230 (N_11230,N_6965,N_5361);
nand U11231 (N_11231,N_8546,N_8884);
nor U11232 (N_11232,N_6966,N_5360);
xnor U11233 (N_11233,N_7428,N_6420);
or U11234 (N_11234,N_6610,N_5126);
nor U11235 (N_11235,N_6835,N_9275);
nand U11236 (N_11236,N_5322,N_7221);
nand U11237 (N_11237,N_9070,N_8590);
and U11238 (N_11238,N_9729,N_9011);
nand U11239 (N_11239,N_5989,N_7109);
and U11240 (N_11240,N_9692,N_8027);
nor U11241 (N_11241,N_7957,N_9085);
or U11242 (N_11242,N_5029,N_7465);
and U11243 (N_11243,N_6444,N_6486);
xnor U11244 (N_11244,N_7208,N_5745);
and U11245 (N_11245,N_7163,N_5414);
or U11246 (N_11246,N_9647,N_8878);
nand U11247 (N_11247,N_5946,N_6721);
nand U11248 (N_11248,N_5870,N_7945);
nand U11249 (N_11249,N_5609,N_5762);
nor U11250 (N_11250,N_9442,N_8820);
and U11251 (N_11251,N_8897,N_5982);
nor U11252 (N_11252,N_5632,N_9779);
nor U11253 (N_11253,N_7496,N_6565);
or U11254 (N_11254,N_5548,N_5377);
nand U11255 (N_11255,N_9871,N_8602);
nand U11256 (N_11256,N_7556,N_5117);
nand U11257 (N_11257,N_7127,N_6449);
xor U11258 (N_11258,N_9982,N_9714);
nor U11259 (N_11259,N_7958,N_8665);
nand U11260 (N_11260,N_8098,N_5090);
or U11261 (N_11261,N_9241,N_5077);
or U11262 (N_11262,N_7611,N_9041);
or U11263 (N_11263,N_8999,N_7154);
or U11264 (N_11264,N_8902,N_5104);
nor U11265 (N_11265,N_8692,N_7874);
nand U11266 (N_11266,N_6340,N_8010);
nor U11267 (N_11267,N_8386,N_9944);
and U11268 (N_11268,N_8811,N_6673);
or U11269 (N_11269,N_8022,N_5684);
xnor U11270 (N_11270,N_8170,N_6385);
or U11271 (N_11271,N_9077,N_5910);
or U11272 (N_11272,N_9502,N_5963);
or U11273 (N_11273,N_5271,N_6472);
nand U11274 (N_11274,N_5567,N_9342);
xor U11275 (N_11275,N_9858,N_8046);
and U11276 (N_11276,N_8516,N_5140);
and U11277 (N_11277,N_7667,N_5287);
or U11278 (N_11278,N_6465,N_5735);
xnor U11279 (N_11279,N_6693,N_5270);
or U11280 (N_11280,N_9142,N_8238);
or U11281 (N_11281,N_9104,N_8919);
nor U11282 (N_11282,N_8528,N_7204);
nor U11283 (N_11283,N_6657,N_5247);
nand U11284 (N_11284,N_6900,N_6708);
xor U11285 (N_11285,N_7987,N_9118);
nand U11286 (N_11286,N_5759,N_5262);
nand U11287 (N_11287,N_7722,N_8504);
nor U11288 (N_11288,N_7157,N_8247);
or U11289 (N_11289,N_5794,N_7473);
or U11290 (N_11290,N_6398,N_6829);
nor U11291 (N_11291,N_6895,N_8830);
and U11292 (N_11292,N_8189,N_6064);
or U11293 (N_11293,N_6998,N_5464);
or U11294 (N_11294,N_5405,N_9898);
or U11295 (N_11295,N_5332,N_9964);
nand U11296 (N_11296,N_6458,N_6231);
xor U11297 (N_11297,N_8030,N_5677);
xor U11298 (N_11298,N_7685,N_9600);
and U11299 (N_11299,N_9155,N_7983);
nand U11300 (N_11300,N_9619,N_9773);
or U11301 (N_11301,N_5911,N_9457);
and U11302 (N_11302,N_8986,N_6516);
or U11303 (N_11303,N_7107,N_5133);
and U11304 (N_11304,N_5724,N_7594);
nor U11305 (N_11305,N_9172,N_5101);
nor U11306 (N_11306,N_9646,N_9090);
nand U11307 (N_11307,N_5398,N_9284);
and U11308 (N_11308,N_5884,N_6771);
nand U11309 (N_11309,N_7181,N_9555);
nor U11310 (N_11310,N_6794,N_5709);
xor U11311 (N_11311,N_6936,N_6722);
or U11312 (N_11312,N_6543,N_7686);
and U11313 (N_11313,N_9071,N_7131);
or U11314 (N_11314,N_7566,N_9664);
nor U11315 (N_11315,N_6717,N_8713);
or U11316 (N_11316,N_8548,N_7579);
nand U11317 (N_11317,N_7099,N_7714);
and U11318 (N_11318,N_9292,N_6202);
and U11319 (N_11319,N_8728,N_9679);
or U11320 (N_11320,N_9640,N_7046);
or U11321 (N_11321,N_6668,N_8777);
nand U11322 (N_11322,N_6579,N_6180);
nand U11323 (N_11323,N_5142,N_7488);
nand U11324 (N_11324,N_9222,N_5687);
nand U11325 (N_11325,N_8676,N_7323);
or U11326 (N_11326,N_7792,N_7256);
or U11327 (N_11327,N_9243,N_9916);
nand U11328 (N_11328,N_6243,N_7158);
nor U11329 (N_11329,N_6629,N_5100);
and U11330 (N_11330,N_8636,N_5099);
or U11331 (N_11331,N_7222,N_7239);
and U11332 (N_11332,N_5981,N_9902);
nand U11333 (N_11333,N_8276,N_9335);
and U11334 (N_11334,N_9514,N_9168);
or U11335 (N_11335,N_5112,N_9979);
nor U11336 (N_11336,N_7004,N_8019);
and U11337 (N_11337,N_6898,N_5061);
and U11338 (N_11338,N_8233,N_8032);
nand U11339 (N_11339,N_8513,N_8866);
nand U11340 (N_11340,N_6730,N_6943);
and U11341 (N_11341,N_8844,N_6395);
and U11342 (N_11342,N_9562,N_6517);
and U11343 (N_11343,N_8695,N_5436);
nor U11344 (N_11344,N_5529,N_7670);
and U11345 (N_11345,N_7348,N_7526);
or U11346 (N_11346,N_9832,N_6686);
nor U11347 (N_11347,N_7970,N_6606);
xor U11348 (N_11348,N_5841,N_9412);
nand U11349 (N_11349,N_8174,N_8204);
and U11350 (N_11350,N_5636,N_8090);
and U11351 (N_11351,N_9879,N_5235);
nand U11352 (N_11352,N_6560,N_6439);
and U11353 (N_11353,N_7085,N_5393);
and U11354 (N_11354,N_5340,N_9028);
or U11355 (N_11355,N_7344,N_7346);
nor U11356 (N_11356,N_5431,N_9177);
nor U11357 (N_11357,N_9765,N_9309);
nand U11358 (N_11358,N_5991,N_8494);
nor U11359 (N_11359,N_7314,N_5068);
and U11360 (N_11360,N_9367,N_6297);
xnor U11361 (N_11361,N_5391,N_9948);
or U11362 (N_11362,N_6618,N_6381);
nor U11363 (N_11363,N_9891,N_5215);
xor U11364 (N_11364,N_8553,N_8690);
or U11365 (N_11365,N_5289,N_6774);
and U11366 (N_11366,N_5500,N_7342);
nor U11367 (N_11367,N_9167,N_7083);
nor U11368 (N_11368,N_5621,N_7573);
or U11369 (N_11369,N_6053,N_9461);
nand U11370 (N_11370,N_8744,N_7690);
nor U11371 (N_11371,N_9701,N_6151);
and U11372 (N_11372,N_5177,N_9426);
nor U11373 (N_11373,N_7485,N_7736);
nor U11374 (N_11374,N_9517,N_7284);
and U11375 (N_11375,N_8003,N_5244);
nor U11376 (N_11376,N_7382,N_9997);
nor U11377 (N_11377,N_9520,N_6059);
or U11378 (N_11378,N_7978,N_7967);
or U11379 (N_11379,N_7775,N_9670);
nor U11380 (N_11380,N_7539,N_6720);
nor U11381 (N_11381,N_9165,N_8275);
xor U11382 (N_11382,N_5190,N_9269);
and U11383 (N_11383,N_8360,N_5443);
or U11384 (N_11384,N_6287,N_5828);
nand U11385 (N_11385,N_7647,N_9763);
nand U11386 (N_11386,N_6121,N_8225);
and U11387 (N_11387,N_8486,N_8680);
xor U11388 (N_11388,N_7604,N_7984);
and U11389 (N_11389,N_9397,N_8144);
nand U11390 (N_11390,N_7857,N_6322);
or U11391 (N_11391,N_9369,N_7171);
nor U11392 (N_11392,N_6167,N_7480);
nor U11393 (N_11393,N_9582,N_5399);
or U11394 (N_11394,N_6605,N_9361);
or U11395 (N_11395,N_8550,N_5769);
xor U11396 (N_11396,N_5161,N_5202);
nor U11397 (N_11397,N_5643,N_7616);
nand U11398 (N_11398,N_9286,N_9006);
and U11399 (N_11399,N_7162,N_7300);
or U11400 (N_11400,N_7475,N_6834);
xor U11401 (N_11401,N_5783,N_5210);
nor U11402 (N_11402,N_8943,N_5167);
or U11403 (N_11403,N_8611,N_8422);
xnor U11404 (N_11404,N_9956,N_8040);
or U11405 (N_11405,N_8781,N_7199);
and U11406 (N_11406,N_8416,N_5886);
or U11407 (N_11407,N_9983,N_8705);
xnor U11408 (N_11408,N_8388,N_8955);
nand U11409 (N_11409,N_9490,N_6980);
xor U11410 (N_11410,N_7298,N_9909);
or U11411 (N_11411,N_7638,N_6881);
or U11412 (N_11412,N_9125,N_9612);
nor U11413 (N_11413,N_5154,N_9620);
nor U11414 (N_11414,N_7486,N_8581);
and U11415 (N_11415,N_5095,N_8484);
and U11416 (N_11416,N_8618,N_6416);
nor U11417 (N_11417,N_6946,N_9809);
nor U11418 (N_11418,N_8615,N_7689);
xor U11419 (N_11419,N_6632,N_7724);
and U11420 (N_11420,N_6795,N_9370);
nor U11421 (N_11421,N_8359,N_8299);
or U11422 (N_11422,N_6993,N_6300);
or U11423 (N_11423,N_6864,N_7326);
nor U11424 (N_11424,N_8821,N_7505);
and U11425 (N_11425,N_6315,N_9351);
nor U11426 (N_11426,N_6757,N_6865);
xor U11427 (N_11427,N_8613,N_7339);
nand U11428 (N_11428,N_7194,N_8301);
xnor U11429 (N_11429,N_5341,N_5540);
nand U11430 (N_11430,N_5198,N_8350);
nand U11431 (N_11431,N_6921,N_5835);
nor U11432 (N_11432,N_5025,N_8814);
nor U11433 (N_11433,N_7665,N_6025);
xor U11434 (N_11434,N_6011,N_8340);
nor U11435 (N_11435,N_6575,N_8143);
nand U11436 (N_11436,N_7841,N_6513);
nand U11437 (N_11437,N_9390,N_6985);
or U11438 (N_11438,N_8883,N_8877);
or U11439 (N_11439,N_7248,N_7868);
nand U11440 (N_11440,N_8737,N_8393);
nor U11441 (N_11441,N_6671,N_7287);
or U11442 (N_11442,N_7699,N_8648);
nand U11443 (N_11443,N_5971,N_8511);
nand U11444 (N_11444,N_8622,N_8612);
nand U11445 (N_11445,N_9067,N_5356);
or U11446 (N_11446,N_6643,N_9194);
xor U11447 (N_11447,N_8570,N_6911);
or U11448 (N_11448,N_9528,N_8559);
nand U11449 (N_11449,N_9615,N_8661);
nor U11450 (N_11450,N_9084,N_9252);
nand U11451 (N_11451,N_7244,N_6269);
or U11452 (N_11452,N_6944,N_6601);
xnor U11453 (N_11453,N_6425,N_5938);
or U11454 (N_11454,N_8605,N_6096);
and U11455 (N_11455,N_9420,N_7352);
nand U11456 (N_11456,N_7291,N_5580);
xor U11457 (N_11457,N_8461,N_6161);
and U11458 (N_11458,N_6076,N_8880);
xor U11459 (N_11459,N_7089,N_5691);
nand U11460 (N_11460,N_8025,N_7311);
nand U11461 (N_11461,N_7886,N_6332);
and U11462 (N_11462,N_6846,N_6377);
xnor U11463 (N_11463,N_7773,N_7713);
nand U11464 (N_11464,N_6922,N_6445);
nor U11465 (N_11465,N_7528,N_5432);
and U11466 (N_11466,N_9603,N_7966);
nand U11467 (N_11467,N_5960,N_5196);
or U11468 (N_11468,N_8178,N_8259);
and U11469 (N_11469,N_6473,N_9326);
or U11470 (N_11470,N_8949,N_6330);
xor U11471 (N_11471,N_6681,N_5460);
nand U11472 (N_11472,N_6283,N_9199);
nand U11473 (N_11473,N_9598,N_6371);
and U11474 (N_11474,N_6863,N_8558);
and U11475 (N_11475,N_6711,N_9299);
and U11476 (N_11476,N_9029,N_6918);
xor U11477 (N_11477,N_8368,N_6070);
nand U11478 (N_11478,N_9339,N_7082);
xnor U11479 (N_11479,N_7503,N_6802);
nor U11480 (N_11480,N_8496,N_6374);
or U11481 (N_11481,N_7021,N_6737);
nand U11482 (N_11482,N_8535,N_8725);
xnor U11483 (N_11483,N_7061,N_8701);
nor U11484 (N_11484,N_8656,N_5429);
or U11485 (N_11485,N_5199,N_6614);
nor U11486 (N_11486,N_6697,N_9388);
nor U11487 (N_11487,N_7910,N_6827);
and U11488 (N_11488,N_9343,N_5814);
nand U11489 (N_11489,N_9697,N_7288);
nand U11490 (N_11490,N_9225,N_8459);
or U11491 (N_11491,N_6623,N_5993);
nor U11492 (N_11492,N_8310,N_9753);
or U11493 (N_11493,N_7443,N_5951);
nand U11494 (N_11494,N_7463,N_6761);
nand U11495 (N_11495,N_5974,N_8981);
nand U11496 (N_11496,N_9216,N_7008);
or U11497 (N_11497,N_7550,N_5044);
nand U11498 (N_11498,N_7002,N_9819);
and U11499 (N_11499,N_8726,N_8062);
nand U11500 (N_11500,N_7319,N_5711);
and U11501 (N_11501,N_7103,N_9955);
and U11502 (N_11502,N_7976,N_8639);
nor U11503 (N_11503,N_6170,N_8735);
nand U11504 (N_11504,N_7033,N_9684);
nor U11505 (N_11505,N_8415,N_5276);
nor U11506 (N_11506,N_5469,N_7459);
or U11507 (N_11507,N_9130,N_5131);
and U11508 (N_11508,N_9324,N_6791);
nor U11509 (N_11509,N_6529,N_9113);
and U11510 (N_11510,N_7226,N_7230);
and U11511 (N_11511,N_6886,N_6116);
and U11512 (N_11512,N_6745,N_8899);
nand U11513 (N_11513,N_5375,N_5809);
nand U11514 (N_11514,N_8401,N_8444);
and U11515 (N_11515,N_9516,N_7921);
nor U11516 (N_11516,N_5465,N_6817);
xnor U11517 (N_11517,N_9025,N_8699);
nand U11518 (N_11518,N_6261,N_5354);
nor U11519 (N_11519,N_5965,N_8599);
and U11520 (N_11520,N_8638,N_8668);
xnor U11521 (N_11521,N_7656,N_8502);
nand U11522 (N_11522,N_6403,N_9340);
nor U11523 (N_11523,N_6664,N_9584);
or U11524 (N_11524,N_6550,N_6592);
or U11525 (N_11525,N_8965,N_5492);
or U11526 (N_11526,N_6855,N_7912);
nand U11527 (N_11527,N_6751,N_5349);
xor U11528 (N_11528,N_5642,N_6776);
nor U11529 (N_11529,N_8035,N_7982);
nand U11530 (N_11530,N_9100,N_6556);
xnor U11531 (N_11531,N_9380,N_5036);
nor U11532 (N_11532,N_5155,N_7995);
or U11533 (N_11533,N_6265,N_6271);
nand U11534 (N_11534,N_9035,N_9158);
nand U11535 (N_11535,N_9303,N_8018);
nor U11536 (N_11536,N_8741,N_7700);
nor U11537 (N_11537,N_5913,N_5325);
or U11538 (N_11538,N_9312,N_5516);
and U11539 (N_11539,N_6277,N_6906);
nor U11540 (N_11540,N_8766,N_6804);
nand U11541 (N_11541,N_7761,N_8985);
nand U11542 (N_11542,N_5940,N_8711);
nand U11543 (N_11543,N_6095,N_7279);
or U11544 (N_11544,N_9625,N_6577);
nand U11545 (N_11545,N_9258,N_7575);
or U11546 (N_11546,N_8662,N_5655);
nor U11547 (N_11547,N_8759,N_9638);
or U11548 (N_11548,N_5698,N_7047);
nand U11549 (N_11549,N_7805,N_9518);
xor U11550 (N_11550,N_8874,N_9410);
and U11551 (N_11551,N_5283,N_5193);
xor U11552 (N_11552,N_9987,N_6176);
nand U11553 (N_11553,N_6678,N_5757);
nor U11554 (N_11554,N_5400,N_8297);
and U11555 (N_11555,N_5324,N_6518);
and U11556 (N_11556,N_6058,N_6043);
and U11557 (N_11557,N_6843,N_7668);
xnor U11558 (N_11558,N_9581,N_9124);
nor U11559 (N_11559,N_7977,N_5744);
or U11560 (N_11560,N_7795,N_5227);
or U11561 (N_11561,N_6128,N_9827);
or U11562 (N_11562,N_7051,N_5842);
and U11563 (N_11563,N_9977,N_5671);
nand U11564 (N_11564,N_8078,N_5020);
or U11565 (N_11565,N_6173,N_8970);
nand U11566 (N_11566,N_8794,N_7591);
nor U11567 (N_11567,N_8371,N_9224);
or U11568 (N_11568,N_9774,N_9608);
and U11569 (N_11569,N_5105,N_9176);
nand U11570 (N_11570,N_7854,N_6930);
nor U11571 (N_11571,N_5312,N_9086);
and U11572 (N_11572,N_9327,N_6238);
and U11573 (N_11573,N_6294,N_5554);
xnor U11574 (N_11574,N_8891,N_7543);
nand U11575 (N_11575,N_9865,N_8529);
and U11576 (N_11576,N_5515,N_7517);
and U11577 (N_11577,N_5387,N_8302);
or U11578 (N_11578,N_6604,N_7953);
or U11579 (N_11579,N_6392,N_5517);
nand U11580 (N_11580,N_9197,N_7418);
nand U11581 (N_11581,N_5249,N_6754);
nand U11582 (N_11582,N_6738,N_7732);
nand U11583 (N_11583,N_8364,N_9651);
nor U11584 (N_11584,N_5606,N_6626);
and U11585 (N_11585,N_9807,N_9973);
xnor U11586 (N_11586,N_5474,N_6400);
and U11587 (N_11587,N_7165,N_7327);
and U11588 (N_11588,N_7316,N_7555);
or U11589 (N_11589,N_7964,N_5455);
and U11590 (N_11590,N_8560,N_8755);
and U11591 (N_11591,N_5751,N_9855);
xor U11592 (N_11592,N_6940,N_7059);
nand U11593 (N_11593,N_9512,N_8246);
or U11594 (N_11594,N_6957,N_9399);
xor U11595 (N_11595,N_5523,N_6713);
nor U11596 (N_11596,N_6241,N_9781);
nor U11597 (N_11597,N_5267,N_6907);
or U11598 (N_11598,N_7210,N_8537);
or U11599 (N_11599,N_5532,N_6547);
or U11600 (N_11600,N_6154,N_8309);
or U11601 (N_11601,N_5588,N_9045);
nand U11602 (N_11602,N_8306,N_9031);
and U11603 (N_11603,N_9147,N_5321);
or U11604 (N_11604,N_7902,N_6292);
xnor U11605 (N_11605,N_7232,N_9300);
or U11606 (N_11606,N_5707,N_8325);
or U11607 (N_11607,N_9493,N_7754);
nand U11608 (N_11608,N_7057,N_5047);
or U11609 (N_11609,N_8006,N_7034);
and U11610 (N_11610,N_5032,N_6317);
or U11611 (N_11611,N_5667,N_8167);
nor U11612 (N_11612,N_5231,N_9060);
nor U11613 (N_11613,N_5306,N_7909);
or U11614 (N_11614,N_7410,N_6756);
xnor U11615 (N_11615,N_6755,N_7328);
and U11616 (N_11616,N_7624,N_7743);
and U11617 (N_11617,N_8751,N_7280);
xor U11618 (N_11618,N_6216,N_9601);
or U11619 (N_11619,N_6075,N_6785);
and U11620 (N_11620,N_7585,N_5313);
nand U11621 (N_11621,N_5560,N_6531);
and U11622 (N_11622,N_5659,N_7552);
or U11623 (N_11623,N_8914,N_7153);
nand U11624 (N_11624,N_9436,N_9058);
or U11625 (N_11625,N_6496,N_9094);
nand U11626 (N_11626,N_8432,N_5549);
or U11627 (N_11627,N_7998,N_6821);
xnor U11628 (N_11628,N_6824,N_6046);
nand U11629 (N_11629,N_6672,N_5878);
nand U11630 (N_11630,N_5813,N_6500);
nand U11631 (N_11631,N_7078,N_8100);
nand U11632 (N_11632,N_8626,N_9654);
nor U11633 (N_11633,N_8357,N_6081);
or U11634 (N_11634,N_7807,N_9016);
or U11635 (N_11635,N_9231,N_9831);
nor U11636 (N_11636,N_7498,N_9875);
or U11637 (N_11637,N_8761,N_7850);
xnor U11638 (N_11638,N_9007,N_7851);
nor U11639 (N_11639,N_9509,N_8993);
nand U11640 (N_11640,N_5510,N_8059);
or U11641 (N_11641,N_5378,N_5573);
nand U11642 (N_11642,N_5594,N_5795);
nand U11643 (N_11643,N_5489,N_7875);
nor U11644 (N_11644,N_9009,N_8083);
and U11645 (N_11645,N_7580,N_5611);
and U11646 (N_11646,N_7618,N_6082);
nand U11647 (N_11647,N_5372,N_6587);
nand U11648 (N_11648,N_9961,N_8400);
nand U11649 (N_11649,N_6347,N_9310);
nand U11650 (N_11650,N_5650,N_7247);
nand U11651 (N_11651,N_6339,N_6909);
nand U11652 (N_11652,N_9703,N_8730);
or U11653 (N_11653,N_8568,N_5803);
or U11654 (N_11654,N_5608,N_8421);
xor U11655 (N_11655,N_7456,N_5717);
nor U11656 (N_11656,N_8241,N_9164);
nor U11657 (N_11657,N_5362,N_9834);
or U11658 (N_11658,N_6155,N_9506);
nand U11659 (N_11659,N_5388,N_7554);
nand U11660 (N_11660,N_6942,N_9508);
and U11661 (N_11661,N_7268,N_6904);
or U11662 (N_11662,N_6410,N_8209);
nor U11663 (N_11663,N_6446,N_6063);
and U11664 (N_11664,N_8817,N_7546);
and U11665 (N_11665,N_8466,N_9971);
or U11666 (N_11666,N_9048,N_9524);
and U11667 (N_11667,N_8375,N_5949);
xnor U11668 (N_11668,N_7706,N_5402);
and U11669 (N_11669,N_8976,N_6122);
nor U11670 (N_11670,N_7731,N_8326);
or U11671 (N_11671,N_5353,N_5923);
or U11672 (N_11672,N_7735,N_9123);
nor U11673 (N_11673,N_6463,N_7635);
xor U11674 (N_11674,N_7041,N_9993);
or U11675 (N_11675,N_5898,N_7943);
and U11676 (N_11676,N_7778,N_6502);
xor U11677 (N_11677,N_5134,N_7877);
or U11678 (N_11678,N_8860,N_9485);
or U11679 (N_11679,N_8869,N_7042);
or U11680 (N_11680,N_8812,N_6422);
and U11681 (N_11681,N_6655,N_5413);
and U11682 (N_11682,N_7564,N_6545);
nand U11683 (N_11683,N_5605,N_7780);
and U11684 (N_11684,N_5092,N_8337);
and U11685 (N_11685,N_6417,N_8240);
nor U11686 (N_11686,N_8780,N_7981);
nand U11687 (N_11687,N_8727,N_7119);
xnor U11688 (N_11688,N_8913,N_8900);
or U11689 (N_11689,N_5384,N_7285);
nor U11690 (N_11690,N_5394,N_6022);
nand U11691 (N_11691,N_9616,N_6553);
or U11692 (N_11692,N_8629,N_9246);
or U11693 (N_11693,N_7460,N_5511);
nand U11694 (N_11694,N_9498,N_6640);
nor U11695 (N_11695,N_8474,N_9623);
nand U11696 (N_11696,N_9226,N_5577);
and U11697 (N_11697,N_9484,N_5151);
and U11698 (N_11698,N_7273,N_5454);
or U11699 (N_11699,N_8153,N_6047);
and U11700 (N_11700,N_6360,N_5422);
nor U11701 (N_11701,N_9248,N_5444);
nor U11702 (N_11702,N_8135,N_8806);
xor U11703 (N_11703,N_7717,N_9102);
and U11704 (N_11704,N_9414,N_6563);
nor U11705 (N_11705,N_5679,N_5057);
or U11706 (N_11706,N_8947,N_7838);
and U11707 (N_11707,N_6247,N_9737);
or U11708 (N_11708,N_7657,N_5397);
and U11709 (N_11709,N_6273,N_9010);
nand U11710 (N_11710,N_5708,N_5900);
xnor U11711 (N_11711,N_6851,N_6558);
and U11712 (N_11712,N_5559,N_9677);
and U11713 (N_11713,N_9250,N_5729);
xnor U11714 (N_11714,N_6326,N_8509);
nor U11715 (N_11715,N_6051,N_9789);
nor U11716 (N_11716,N_6828,N_8264);
nor U11717 (N_11717,N_7015,N_6949);
nor U11718 (N_11718,N_7179,N_8838);
or U11719 (N_11719,N_9846,N_7728);
and U11720 (N_11720,N_5771,N_5365);
or U11721 (N_11721,N_7669,N_9293);
or U11722 (N_11722,N_9936,N_9757);
and U11723 (N_11723,N_5656,N_8185);
and U11724 (N_11724,N_9120,N_9583);
nor U11725 (N_11725,N_8608,N_7802);
xnor U11726 (N_11726,N_5772,N_6544);
or U11727 (N_11727,N_7055,N_8968);
xor U11728 (N_11728,N_8621,N_5268);
xnor U11729 (N_11729,N_9262,N_9103);
nor U11730 (N_11730,N_7255,N_9527);
nand U11731 (N_11731,N_9240,N_6192);
xnor U11732 (N_11732,N_8774,N_7312);
and U11733 (N_11733,N_5950,N_9784);
nor U11734 (N_11734,N_8110,N_7423);
nor U11735 (N_11735,N_8441,N_5890);
nor U11736 (N_11736,N_7254,N_9770);
nor U11737 (N_11737,N_6747,N_7358);
nand U11738 (N_11738,N_8481,N_9658);
or U11739 (N_11739,N_5914,N_9593);
nor U11740 (N_11740,N_9878,N_6688);
or U11741 (N_11741,N_5088,N_8091);
or U11742 (N_11742,N_8107,N_9577);
and U11743 (N_11743,N_8467,N_6964);
and U11744 (N_11744,N_6026,N_6275);
nor U11745 (N_11745,N_5579,N_7884);
or U11746 (N_11746,N_8635,N_5616);
xor U11747 (N_11747,N_9446,N_8044);
and U11748 (N_11748,N_8961,N_7655);
or U11749 (N_11749,N_5582,N_5927);
or U11750 (N_11750,N_8849,N_9488);
nor U11751 (N_11751,N_9434,N_9000);
and U11752 (N_11752,N_7557,N_8115);
or U11753 (N_11753,N_6838,N_6138);
and U11754 (N_11754,N_9244,N_9402);
nor U11755 (N_11755,N_8007,N_9602);
and U11756 (N_11756,N_8885,N_7414);
xnor U11757 (N_11757,N_7553,N_6117);
or U11758 (N_11758,N_5488,N_7845);
or U11759 (N_11759,N_7010,N_6426);
and U11760 (N_11760,N_8305,N_9751);
and U11761 (N_11761,N_5205,N_6418);
or U11762 (N_11762,N_5337,N_8578);
and U11763 (N_11763,N_6123,N_6945);
or U11764 (N_11764,N_8533,N_5186);
and U11765 (N_11765,N_5471,N_8819);
nor U11766 (N_11766,N_6365,N_6211);
or U11767 (N_11767,N_6078,N_5880);
or U11768 (N_11768,N_9454,N_5062);
nand U11769 (N_11769,N_6524,N_6892);
xnor U11770 (N_11770,N_5096,N_8430);
or U11771 (N_11771,N_8996,N_9027);
nor U11772 (N_11772,N_6631,N_8829);
or U11773 (N_11773,N_9808,N_8478);
or U11774 (N_11774,N_7510,N_7231);
and U11775 (N_11775,N_7161,N_6675);
nor U11776 (N_11776,N_9372,N_7014);
nand U11777 (N_11777,N_7395,N_6129);
nor U11778 (N_11778,N_6506,N_7394);
or U11779 (N_11779,N_8050,N_9496);
or U11780 (N_11780,N_8684,N_6679);
nand U11781 (N_11781,N_9663,N_6471);
nand U11782 (N_11782,N_6508,N_8669);
nor U11783 (N_11783,N_9218,N_6710);
nand U11784 (N_11784,N_8232,N_5908);
or U11785 (N_11785,N_9186,N_8783);
and U11786 (N_11786,N_9347,N_5411);
nand U11787 (N_11787,N_7461,N_6992);
nor U11788 (N_11788,N_7664,N_6536);
or U11789 (N_11789,N_8434,N_9764);
nor U11790 (N_11790,N_5860,N_9317);
and U11791 (N_11791,N_6837,N_6562);
nor U11792 (N_11792,N_9236,N_7574);
and U11793 (N_11793,N_6165,N_5119);
or U11794 (N_11794,N_7988,N_9032);
nor U11795 (N_11795,N_5430,N_7309);
nor U11796 (N_11796,N_8498,N_8113);
xnor U11797 (N_11797,N_9794,N_5303);
xnor U11798 (N_11798,N_9153,N_9727);
and U11799 (N_11799,N_9237,N_8807);
nor U11800 (N_11800,N_7519,N_5779);
nor U11801 (N_11801,N_9184,N_7391);
nand U11802 (N_11802,N_6849,N_7969);
or U11803 (N_11803,N_9700,N_5037);
and U11804 (N_11804,N_5490,N_5663);
nor U11805 (N_11805,N_7432,N_9945);
or U11806 (N_11806,N_7114,N_7629);
and U11807 (N_11807,N_9355,N_6198);
nor U11808 (N_11808,N_5689,N_7228);
and U11809 (N_11809,N_6018,N_5053);
or U11810 (N_11810,N_6870,N_6358);
or U11811 (N_11811,N_7250,N_8540);
nand U11812 (N_11812,N_6233,N_8853);
or U11813 (N_11813,N_9198,N_9864);
xor U11814 (N_11814,N_5022,N_9476);
and U11815 (N_11815,N_7166,N_5382);
and U11816 (N_11816,N_5309,N_6739);
nand U11817 (N_11817,N_7100,N_5834);
or U11818 (N_11818,N_8391,N_8001);
nand U11819 (N_11819,N_9179,N_7610);
nand U11820 (N_11820,N_6986,N_6534);
xnor U11821 (N_11821,N_7468,N_8120);
xnor U11822 (N_11822,N_6984,N_8211);
or U11823 (N_11823,N_8534,N_9935);
xor U11824 (N_11824,N_6153,N_6656);
nor U11825 (N_11825,N_6919,N_7887);
or U11826 (N_11826,N_7176,N_5558);
nor U11827 (N_11827,N_8723,N_9215);
nand U11828 (N_11828,N_9570,N_6354);
and U11829 (N_11829,N_9797,N_6160);
nand U11830 (N_11830,N_9075,N_5323);
or U11831 (N_11831,N_8155,N_8243);
nor U11832 (N_11832,N_6455,N_8382);
nor U11833 (N_11833,N_7811,N_5931);
nor U11834 (N_11834,N_5919,N_7399);
nand U11835 (N_11835,N_5941,N_8805);
or U11836 (N_11836,N_8043,N_7141);
or U11837 (N_11837,N_5858,N_7092);
or U11838 (N_11838,N_9665,N_8939);
nor U11839 (N_11839,N_6184,N_7709);
nor U11840 (N_11840,N_6430,N_6595);
xor U11841 (N_11841,N_9515,N_5830);
and U11842 (N_11842,N_7155,N_9191);
nor U11843 (N_11843,N_5756,N_6142);
nor U11844 (N_11844,N_9921,N_7772);
and U11845 (N_11845,N_9195,N_6363);
or U11846 (N_11846,N_8033,N_9428);
and U11847 (N_11847,N_7310,N_9880);
and U11848 (N_11848,N_9885,N_6359);
nand U11849 (N_11849,N_9037,N_6114);
and U11850 (N_11850,N_7882,N_8746);
nor U11851 (N_11851,N_6699,N_8667);
or U11852 (N_11852,N_5296,N_8823);
or U11853 (N_11853,N_6411,N_6435);
nand U11854 (N_11854,N_5158,N_7499);
nand U11855 (N_11855,N_9540,N_8220);
nor U11856 (N_11856,N_7677,N_5171);
nand U11857 (N_11857,N_8454,N_6157);
nor U11858 (N_11858,N_5736,N_6770);
and U11859 (N_11859,N_6441,N_5067);
or U11860 (N_11860,N_7446,N_5049);
or U11861 (N_11861,N_7431,N_9182);
and U11862 (N_11862,N_7397,N_7262);
xor U11863 (N_11863,N_9068,N_5410);
xnor U11864 (N_11864,N_5619,N_5700);
and U11865 (N_11865,N_9668,N_6796);
and U11866 (N_11866,N_6033,N_6382);
nand U11867 (N_11867,N_5371,N_5596);
nor U11868 (N_11868,N_6685,N_5788);
xor U11869 (N_11869,N_9958,N_6867);
xnor U11870 (N_11870,N_6139,N_7715);
or U11871 (N_11871,N_5427,N_7497);
nor U11872 (N_11872,N_9782,N_9817);
nor U11873 (N_11873,N_7371,N_6612);
and U11874 (N_11874,N_9890,N_7186);
nor U11875 (N_11875,N_7536,N_7653);
nand U11876 (N_11876,N_6691,N_6104);
or U11877 (N_11877,N_6665,N_5780);
nand U11878 (N_11878,N_7115,N_6235);
nand U11879 (N_11879,N_5174,N_5028);
or U11880 (N_11880,N_5153,N_8342);
and U11881 (N_11881,N_7628,N_5181);
nand U11882 (N_11882,N_8583,N_8601);
nor U11883 (N_11883,N_6725,N_8743);
xor U11884 (N_11884,N_7589,N_9396);
and U11885 (N_11885,N_6947,N_5281);
nand U11886 (N_11886,N_8324,N_8137);
or U11887 (N_11887,N_6206,N_6654);
or U11888 (N_11888,N_7101,N_5467);
and U11889 (N_11889,N_8633,N_8706);
nand U11890 (N_11890,N_7619,N_6630);
or U11891 (N_11891,N_5165,N_7387);
nor U11892 (N_11892,N_6320,N_5333);
nor U11893 (N_11893,N_9857,N_8288);
nor U11894 (N_11894,N_9002,N_7688);
nand U11895 (N_11895,N_6017,N_6278);
nand U11896 (N_11896,N_5753,N_7173);
nor U11897 (N_11897,N_5810,N_7607);
or U11898 (N_11898,N_5007,N_6056);
nor U11899 (N_11899,N_7931,N_5428);
or U11900 (N_11900,N_9860,N_5918);
nor U11901 (N_11901,N_8202,N_6799);
or U11902 (N_11902,N_5426,N_6291);
nand U11903 (N_11903,N_6187,N_8312);
nand U11904 (N_11904,N_9696,N_7548);
and U11905 (N_11905,N_5543,N_8284);
xnor U11906 (N_11906,N_6108,N_6447);
nor U11907 (N_11907,N_8839,N_7940);
nor U11908 (N_11908,N_7630,N_7938);
nand U11909 (N_11909,N_5806,N_8964);
nand U11910 (N_11910,N_5613,N_6143);
and U11911 (N_11911,N_8195,N_7755);
nor U11912 (N_11912,N_9656,N_6036);
xor U11913 (N_11913,N_6353,N_6607);
and U11914 (N_11914,N_8892,N_9178);
or U11915 (N_11915,N_8250,N_5805);
or U11916 (N_11916,N_8835,N_5853);
and U11917 (N_11917,N_6083,N_5008);
or U11918 (N_11918,N_6049,N_8064);
nor U11919 (N_11919,N_7827,N_8002);
nor U11920 (N_11920,N_8845,N_5976);
nand U11921 (N_11921,N_5939,N_6333);
xnor U11922 (N_11922,N_8921,N_7562);
xor U11923 (N_11923,N_8686,N_9676);
and U11924 (N_11924,N_8763,N_5458);
and U11925 (N_11925,N_8334,N_7879);
nand U11926 (N_11926,N_9020,N_6044);
and U11927 (N_11927,N_6328,N_8720);
and U11928 (N_11928,N_7523,N_7597);
nand U11929 (N_11929,N_6054,N_6875);
or U11930 (N_11930,N_8425,N_5063);
nor U11931 (N_11931,N_6812,N_9475);
or U11932 (N_11932,N_5583,N_9161);
and U11933 (N_11933,N_9445,N_6784);
and U11934 (N_11934,N_8760,N_8437);
or U11935 (N_11935,N_7005,N_8445);
or U11936 (N_11936,N_6456,N_8799);
nor U11937 (N_11937,N_7307,N_6969);
and U11938 (N_11938,N_5953,N_7466);
nand U11939 (N_11939,N_7749,N_7203);
or U11940 (N_11940,N_7765,N_8077);
and U11941 (N_11941,N_8200,N_6002);
nor U11942 (N_11942,N_5849,N_9082);
xnor U11943 (N_11943,N_5263,N_8691);
nor U11944 (N_11944,N_9174,N_8588);
nor U11945 (N_11945,N_9321,N_6373);
nand U11946 (N_11946,N_9851,N_7489);
nand U11947 (N_11947,N_9558,N_6788);
nand U11948 (N_11948,N_6394,N_9637);
and U11949 (N_11949,N_6532,N_7948);
nor U11950 (N_11950,N_9483,N_9433);
nand U11951 (N_11951,N_8290,N_6901);
or U11952 (N_11952,N_8655,N_8487);
nand U11953 (N_11953,N_9960,N_7402);
and U11954 (N_11954,N_9187,N_9423);
nand U11955 (N_11955,N_9301,N_7481);
or U11956 (N_11956,N_7939,N_8499);
and U11957 (N_11957,N_8954,N_9091);
and U11958 (N_11958,N_7541,N_9841);
nand U11959 (N_11959,N_9169,N_6372);
or U11960 (N_11960,N_9138,N_7363);
nand U11961 (N_11961,N_8827,N_6442);
nand U11962 (N_11962,N_9984,N_9305);
or U11963 (N_11963,N_9554,N_6807);
and U11964 (N_11964,N_8272,N_6387);
nand U11965 (N_11965,N_8556,N_6067);
nor U11966 (N_11966,N_5081,N_6227);
xor U11967 (N_11967,N_6221,N_7393);
and U11968 (N_11968,N_5026,N_6252);
xor U11969 (N_11969,N_9769,N_9811);
or U11970 (N_11970,N_9023,N_7770);
or U11971 (N_11971,N_7801,N_9005);
nor U11972 (N_11972,N_8709,N_9530);
nand U11973 (N_11973,N_8679,N_9954);
or U11974 (N_11974,N_6538,N_9591);
nand U11975 (N_11975,N_7246,N_7195);
and U11976 (N_11976,N_6872,N_5307);
and U11977 (N_11977,N_6237,N_6810);
nor U11978 (N_11978,N_7818,N_5358);
nand U11979 (N_11979,N_7375,N_5798);
or U11980 (N_11980,N_7790,N_9694);
or U11981 (N_11981,N_8994,N_9205);
nor U11982 (N_11982,N_8294,N_5127);
nand U11983 (N_11983,N_8938,N_5295);
nor U11984 (N_11984,N_5773,N_6493);
nor U11985 (N_11985,N_5449,N_9594);
or U11986 (N_11986,N_8212,N_7177);
and U11987 (N_11987,N_7514,N_6163);
or U11988 (N_11988,N_6489,N_6597);
nor U11989 (N_11989,N_6762,N_7079);
and U11990 (N_11990,N_7645,N_5013);
nand U11991 (N_11991,N_9810,N_9033);
and U11992 (N_11992,N_7106,N_6434);
nor U11993 (N_11993,N_6404,N_5027);
xnor U11994 (N_11994,N_5253,N_6485);
nor U11995 (N_11995,N_8876,N_9354);
nor U11996 (N_11996,N_5612,N_7022);
xnor U11997 (N_11997,N_6832,N_9990);
and U11998 (N_11998,N_6814,N_5218);
or U11999 (N_11999,N_6293,N_6927);
nand U12000 (N_12000,N_8168,N_9539);
xnor U12001 (N_12001,N_6548,N_9336);
or U12002 (N_12002,N_9597,N_6744);
nand U12003 (N_12003,N_7527,N_5635);
and U12004 (N_12004,N_7758,N_6783);
or U12005 (N_12005,N_8547,N_5970);
nand U12006 (N_12006,N_6368,N_9804);
nand U12007 (N_12007,N_9341,N_6166);
nor U12008 (N_12008,N_5071,N_6191);
and U12009 (N_12009,N_7063,N_5916);
nor U12010 (N_12010,N_6195,N_7757);
and U12011 (N_12011,N_8293,N_7037);
nor U12012 (N_12012,N_9923,N_9192);
nor U12013 (N_12013,N_9550,N_6530);
nand U12014 (N_12014,N_5056,N_8480);
and U12015 (N_12015,N_5907,N_5966);
nand U12016 (N_12016,N_5316,N_8358);
nand U12017 (N_12017,N_7520,N_9121);
or U12018 (N_12018,N_9836,N_9210);
nor U12019 (N_12019,N_8254,N_7829);
or U12020 (N_12020,N_7947,N_7973);
xnor U12021 (N_12021,N_7927,N_9018);
and U12022 (N_12022,N_9338,N_7750);
nor U12023 (N_12023,N_5833,N_6779);
and U12024 (N_12024,N_7178,N_6338);
nor U12025 (N_12025,N_8907,N_7833);
and U12026 (N_12026,N_8489,N_7196);
and U12027 (N_12027,N_7172,N_6255);
nor U12028 (N_12028,N_5507,N_5000);
and U12029 (N_12029,N_9064,N_8423);
and U12030 (N_12030,N_5565,N_5335);
nand U12031 (N_12031,N_8593,N_8198);
or U12032 (N_12032,N_5896,N_9723);
nor U12033 (N_12033,N_9080,N_9325);
and U12034 (N_12034,N_8271,N_9127);
xnor U12035 (N_12035,N_8179,N_8215);
nand U12036 (N_12036,N_9693,N_9261);
xor U12037 (N_12037,N_9866,N_5209);
and U12038 (N_12038,N_7839,N_9942);
and U12039 (N_12039,N_7878,N_6790);
or U12040 (N_12040,N_5508,N_7506);
or U12041 (N_12041,N_5093,N_7170);
nand U12042 (N_12042,N_5331,N_8226);
xnor U12043 (N_12043,N_6499,N_5091);
and U12044 (N_12044,N_7146,N_8569);
nand U12045 (N_12045,N_6584,N_5184);
or U12046 (N_12046,N_9160,N_9386);
or U12047 (N_12047,N_5774,N_8343);
nor U12048 (N_12048,N_7024,N_8922);
or U12049 (N_12049,N_6879,N_9375);
nand U12050 (N_12050,N_8847,N_7643);
nor U12051 (N_12051,N_6146,N_9847);
or U12052 (N_12052,N_6857,N_6955);
xnor U12053 (N_12053,N_6119,N_9251);
nor U12054 (N_12054,N_9561,N_5934);
xor U12055 (N_12055,N_7404,N_9705);
xnor U12056 (N_12056,N_7729,N_8733);
xor U12057 (N_12057,N_9745,N_7213);
nand U12058 (N_12058,N_8738,N_9271);
or U12059 (N_12059,N_7274,N_9136);
or U12060 (N_12060,N_6850,N_6183);
and U12061 (N_12061,N_7205,N_6179);
xor U12062 (N_12062,N_6981,N_5571);
and U12063 (N_12063,N_9346,N_6521);
or U12064 (N_12064,N_9083,N_8231);
nand U12065 (N_12065,N_7267,N_6462);
nor U12066 (N_12066,N_9523,N_8351);
xor U12067 (N_12067,N_5369,N_9474);
nand U12068 (N_12068,N_7719,N_6635);
and U12069 (N_12069,N_5912,N_5629);
or U12070 (N_12070,N_6572,N_7919);
and U12071 (N_12071,N_6079,N_5486);
nand U12072 (N_12072,N_5040,N_5146);
nand U12073 (N_12073,N_5704,N_7020);
or U12074 (N_12074,N_9856,N_7509);
nor U12075 (N_12075,N_5305,N_8223);
nor U12076 (N_12076,N_9283,N_9274);
or U12077 (N_12077,N_6651,N_8732);
and U12078 (N_12078,N_5058,N_5342);
xor U12079 (N_12079,N_7676,N_7361);
nand U12080 (N_12080,N_9596,N_6118);
nand U12081 (N_12081,N_6540,N_8768);
xnor U12082 (N_12082,N_6248,N_9140);
nand U12083 (N_12083,N_9995,N_7304);
nand U12084 (N_12084,N_7191,N_6327);
nand U12085 (N_12085,N_9937,N_9219);
or U12086 (N_12086,N_8828,N_9464);
nor U12087 (N_12087,N_8697,N_7184);
nand U12088 (N_12088,N_5280,N_7049);
or U12089 (N_12089,N_7492,N_7028);
and U12090 (N_12090,N_7633,N_7278);
xnor U12091 (N_12091,N_6041,N_8666);
nor U12092 (N_12092,N_6263,N_7345);
nor U12093 (N_12093,N_9294,N_6480);
or U12094 (N_12094,N_7306,N_6289);
and U12095 (N_12095,N_8311,N_6402);
nor U12096 (N_12096,N_9833,N_6852);
nand U12097 (N_12097,N_9950,N_9691);
nor U12098 (N_12098,N_9049,N_8642);
and U12099 (N_12099,N_8600,N_9732);
or U12100 (N_12100,N_9013,N_5265);
nor U12101 (N_12101,N_6963,N_5097);
or U12102 (N_12102,N_6414,N_5730);
nand U12103 (N_12103,N_8521,N_7383);
nor U12104 (N_12104,N_7066,N_8065);
xor U12105 (N_12105,N_7847,N_5299);
nand U12106 (N_12106,N_6147,N_5685);
or U12107 (N_12107,N_7349,N_5945);
or U12108 (N_12108,N_5766,N_9456);
nand U12109 (N_12109,N_6467,N_7069);
nand U12110 (N_12110,N_7577,N_9504);
and U12111 (N_12111,N_6203,N_9499);
or U12112 (N_12112,N_7745,N_7118);
or U12113 (N_12113,N_9913,N_9503);
nor U12114 (N_12114,N_5076,N_9359);
nor U12115 (N_12115,N_7920,N_5591);
or U12116 (N_12116,N_5139,N_7516);
or U12117 (N_12117,N_6573,N_6208);
nor U12118 (N_12118,N_9254,N_8716);
xor U12119 (N_12119,N_5575,N_9440);
and U12120 (N_12120,N_9501,N_6574);
nor U12121 (N_12121,N_8594,N_8654);
and U12122 (N_12122,N_9689,N_7661);
or U12123 (N_12123,N_7329,N_8510);
or U12124 (N_12124,N_7741,N_9313);
nand U12125 (N_12125,N_9578,N_7039);
nand U12126 (N_12126,N_7215,N_6029);
nand U12127 (N_12127,N_5862,N_9904);
and U12128 (N_12128,N_6014,N_9903);
and U12129 (N_12129,N_5922,N_5479);
and U12130 (N_12130,N_8471,N_6970);
and U12131 (N_12131,N_8816,N_5761);
and U12132 (N_12132,N_7762,N_7458);
or U12133 (N_12133,N_9800,N_5672);
nor U12134 (N_12134,N_5079,N_9839);
and U12135 (N_12135,N_5179,N_6093);
and U12136 (N_12136,N_7593,N_9487);
or U12137 (N_12137,N_6511,N_5995);
nor U12138 (N_12138,N_9862,N_6131);
nor U12139 (N_12139,N_7588,N_7318);
nand U12140 (N_12140,N_9099,N_8429);
and U12141 (N_12141,N_5843,N_8224);
nor U12142 (N_12142,N_9867,N_7723);
nor U12143 (N_12143,N_8128,N_7903);
nor U12144 (N_12144,N_5060,N_9553);
nand U12145 (N_12145,N_7364,N_5968);
and U12146 (N_12146,N_9605,N_5728);
nand U12147 (N_12147,N_6028,N_5031);
and U12148 (N_12148,N_9564,N_6896);
nor U12149 (N_12149,N_8557,N_8675);
nand U12150 (N_12150,N_8810,N_7381);
nand U12151 (N_12151,N_6731,N_9220);
and U12152 (N_12152,N_7697,N_5997);
nor U12153 (N_12153,N_8236,N_9985);
or U12154 (N_12154,N_6551,N_7974);
nand U12155 (N_12155,N_8652,N_8647);
nand U12156 (N_12156,N_9323,N_5747);
or U12157 (N_12157,N_8545,N_6021);
nor U12158 (N_12158,N_8129,N_6826);
nand U12159 (N_12159,N_7302,N_9815);
nor U12160 (N_12160,N_6391,N_8150);
xnor U12161 (N_12161,N_7674,N_6475);
and U12162 (N_12162,N_5496,N_8704);
xor U12163 (N_12163,N_8279,N_8657);
nand U12164 (N_12164,N_6150,N_9449);
nand U12165 (N_12165,N_9201,N_5791);
and U12166 (N_12166,N_8565,N_8229);
or U12167 (N_12167,N_6481,N_7572);
and U12168 (N_12168,N_6298,N_9842);
xor U12169 (N_12169,N_9151,N_9463);
and U12170 (N_12170,N_9749,N_9270);
nand U12171 (N_12171,N_7560,N_8906);
xor U12172 (N_12172,N_6763,N_9214);
xnor U12173 (N_12173,N_8795,N_8455);
and U12174 (N_12174,N_8771,N_7405);
and U12175 (N_12175,N_7424,N_7759);
xor U12176 (N_12176,N_9384,N_6498);
or U12177 (N_12177,N_7087,N_7596);
or U12178 (N_12178,N_6588,N_8066);
nor U12179 (N_12179,N_9095,N_8363);
or U12180 (N_12180,N_7708,N_8323);
xnor U12181 (N_12181,N_7961,N_9673);
nor U12182 (N_12182,N_8854,N_7164);
nand U12183 (N_12183,N_9559,N_6001);
nand U12184 (N_12184,N_9994,N_5562);
nand U12185 (N_12185,N_8255,N_5242);
xor U12186 (N_12186,N_5208,N_9953);
xnor U12187 (N_12187,N_7532,N_8651);
nor U12188 (N_12188,N_5715,N_8923);
and U12189 (N_12189,N_7125,N_6960);
nand U12190 (N_12190,N_6642,N_8339);
or U12191 (N_12191,N_6860,N_9962);
or U12192 (N_12192,N_6715,N_6438);
and U12193 (N_12193,N_7737,N_7990);
and U12194 (N_12194,N_5800,N_9759);
nand U12195 (N_12195,N_9674,N_5754);
or U12196 (N_12196,N_6479,N_6736);
nand U12197 (N_12197,N_5984,N_8663);
nand U12198 (N_12198,N_6375,N_8752);
or U12199 (N_12199,N_8984,N_9698);
or U12200 (N_12200,N_8672,N_8118);
nand U12201 (N_12201,N_7045,N_6706);
and U12202 (N_12202,N_7054,N_9098);
nor U12203 (N_12203,N_8991,N_8773);
nor U12204 (N_12204,N_6137,N_6781);
and U12205 (N_12205,N_7626,N_5304);
or U12206 (N_12206,N_9430,N_8462);
nor U12207 (N_12207,N_5994,N_6848);
nor U12208 (N_12208,N_5726,N_7225);
and U12209 (N_12209,N_6099,N_7219);
or U12210 (N_12210,N_5433,N_5239);
nand U12211 (N_12211,N_8585,N_9307);
and U12212 (N_12212,N_5681,N_5533);
nand U12213 (N_12213,N_8653,N_5894);
nand U12214 (N_12214,N_9552,N_6603);
nor U12215 (N_12215,N_7904,N_5569);
nand U12216 (N_12216,N_6306,N_7654);
and U12217 (N_12217,N_5098,N_8145);
nand U12218 (N_12218,N_7330,N_9538);
or U12219 (N_12219,N_7283,N_9911);
or U12220 (N_12220,N_9648,N_6625);
nand U12221 (N_12221,N_5085,N_6734);
nor U12222 (N_12222,N_8717,N_9672);
xor U12223 (N_12223,N_5816,N_5495);
nor U12224 (N_12224,N_6140,N_8765);
xnor U12225 (N_12225,N_9588,N_7019);
and U12226 (N_12226,N_5216,N_5526);
and U12227 (N_12227,N_6854,N_6066);
nand U12228 (N_12228,N_7238,N_8123);
or U12229 (N_12229,N_7132,N_5224);
or U12230 (N_12230,N_7152,N_8644);
nand U12231 (N_12231,N_8803,N_9778);
or U12232 (N_12232,N_8313,N_7671);
or U12233 (N_12233,N_5869,N_5505);
or U12234 (N_12234,N_9383,N_7016);
nand U12235 (N_12235,N_7108,N_7359);
and U12236 (N_12236,N_6214,N_6641);
nor U12237 (N_12237,N_8349,N_8410);
or U12238 (N_12238,N_6304,N_5948);
and U12239 (N_12239,N_5767,N_5257);
xor U12240 (N_12240,N_7090,N_6582);
and U12241 (N_12241,N_7907,N_9115);
or U12242 (N_12242,N_9377,N_6367);
xnor U12243 (N_12243,N_9409,N_6987);
and U12244 (N_12244,N_7500,N_6245);
xnor U12245 (N_12245,N_5897,N_5959);
and U12246 (N_12246,N_8634,N_6274);
nor U12247 (N_12247,N_6929,N_8132);
or U12248 (N_12248,N_6624,N_9604);
and U12249 (N_12249,N_9132,N_5150);
and U12250 (N_12250,N_5106,N_6052);
or U12251 (N_12251,N_7484,N_5682);
or U12252 (N_12252,N_5701,N_8021);
nand U12253 (N_12253,N_8750,N_7702);
nand U12254 (N_12254,N_7237,N_7235);
xor U12255 (N_12255,N_6429,N_9894);
and U12256 (N_12256,N_6727,N_9364);
and U12257 (N_12257,N_5935,N_9724);
or U12258 (N_12258,N_9062,N_8464);
or U12259 (N_12259,N_6801,N_6453);
nor U12260 (N_12260,N_9970,N_7167);
xnor U12261 (N_12261,N_5522,N_6357);
or U12262 (N_12262,N_7721,N_8156);
and U12263 (N_12263,N_9259,N_8384);
nand U12264 (N_12264,N_5648,N_8134);
or U12265 (N_12265,N_5048,N_7355);
nor U12266 (N_12266,N_9333,N_9459);
and U12267 (N_12267,N_8592,N_8376);
and U12268 (N_12268,N_5519,N_8567);
xor U12269 (N_12269,N_6390,N_9611);
xnor U12270 (N_12270,N_7333,N_7515);
nand U12271 (N_12271,N_8042,N_8934);
nor U12272 (N_12272,N_7830,N_5221);
nand U12273 (N_12273,N_5746,N_5420);
or U12274 (N_12274,N_5589,N_6549);
nor U12275 (N_12275,N_8886,N_9331);
nand U12276 (N_12276,N_8093,N_9587);
xor U12277 (N_12277,N_5864,N_7915);
nand U12278 (N_12278,N_7587,N_6196);
nor U12279 (N_12279,N_8826,N_7551);
or U12280 (N_12280,N_7398,N_9805);
nor U12281 (N_12281,N_8191,N_5962);
nor U12282 (N_12282,N_7234,N_9978);
nor U12283 (N_12283,N_6232,N_8791);
and U12284 (N_12284,N_5442,N_5501);
nor U12285 (N_12285,N_7704,N_9206);
or U12286 (N_12286,N_8659,N_9468);
and U12287 (N_12287,N_9919,N_5947);
and U12288 (N_12288,N_8987,N_9991);
or U12289 (N_12289,N_7313,N_5638);
nor U12290 (N_12290,N_7858,N_5240);
and U12291 (N_12291,N_5083,N_6753);
or U12292 (N_12292,N_9959,N_5859);
and U12293 (N_12293,N_9106,N_6808);
nand U12294 (N_12294,N_5317,N_5016);
or U12295 (N_12295,N_7384,N_9744);
nand U12296 (N_12296,N_6646,N_5459);
and U12297 (N_12297,N_8998,N_8208);
nor U12298 (N_12298,N_5557,N_8555);
nor U12299 (N_12299,N_9870,N_8879);
nor U12300 (N_12300,N_8561,N_5875);
nor U12301 (N_12301,N_8361,N_7434);
nor U12302 (N_12302,N_7242,N_9046);
nand U12303 (N_12303,N_5954,N_8843);
or U12304 (N_12304,N_7675,N_5314);
or U12305 (N_12305,N_5692,N_9356);
and U12306 (N_12306,N_6194,N_6695);
nand U12307 (N_12307,N_9304,N_8217);
or U12308 (N_12308,N_5238,N_8253);
and U12309 (N_12309,N_9634,N_9896);
xnor U12310 (N_12310,N_6683,N_5111);
nor U12311 (N_12311,N_7077,N_6687);
nor U12312 (N_12312,N_5123,N_9289);
or U12313 (N_12313,N_6105,N_5004);
or U12314 (N_12314,N_9204,N_5412);
or U12315 (N_12315,N_6515,N_8280);
nor U12316 (N_12316,N_8296,N_5958);
and U12317 (N_12317,N_7768,N_9478);
xor U12318 (N_12318,N_6891,N_8320);
nor U12319 (N_12319,N_6519,N_9641);
nand U12320 (N_12320,N_8818,N_7006);
and U12321 (N_12321,N_9444,N_8698);
and U12322 (N_12322,N_6764,N_8493);
xnor U12323 (N_12323,N_8071,N_5343);
and U12324 (N_12324,N_7281,N_7376);
and U12325 (N_12325,N_6309,N_9820);
nor U12326 (N_12326,N_9816,N_9447);
nand U12327 (N_12327,N_9877,N_5893);
xnor U12328 (N_12328,N_5042,N_8205);
nor U12329 (N_12329,N_7571,N_7789);
nor U12330 (N_12330,N_7292,N_9557);
and U12331 (N_12331,N_9079,N_7493);
or U12332 (N_12332,N_6450,N_8372);
and U12333 (N_12333,N_8848,N_9281);
and U12334 (N_12334,N_5983,N_5651);
nand U12335 (N_12335,N_5564,N_5597);
nand U12336 (N_12336,N_5226,N_5162);
or U12337 (N_12337,N_8152,N_6158);
and U12338 (N_12338,N_6858,N_9471);
or U12339 (N_12339,N_8792,N_6701);
nand U12340 (N_12340,N_6349,N_9803);
or U12341 (N_12341,N_6728,N_5440);
nor U12342 (N_12342,N_7156,N_5450);
and U12343 (N_12343,N_8453,N_7846);
or U12344 (N_12344,N_7692,N_6132);
nor U12345 (N_12345,N_9126,N_7263);
nand U12346 (N_12346,N_6972,N_6714);
nand U12347 (N_12347,N_7390,N_5330);
nor U12348 (N_12348,N_5669,N_8407);
or U12349 (N_12349,N_8181,N_9203);
nor U12350 (N_12350,N_9947,N_5344);
nor U12351 (N_12351,N_6876,N_8928);
or U12352 (N_12352,N_5453,N_5901);
or U12353 (N_12353,N_6760,N_6337);
or U12354 (N_12354,N_9678,N_9657);
nand U12355 (N_12355,N_5657,N_7642);
or U12356 (N_12356,N_9943,N_7102);
or U12357 (N_12357,N_5010,N_8840);
and U12358 (N_12358,N_7537,N_7771);
and U12359 (N_12359,N_8183,N_7701);
nand U12360 (N_12360,N_6200,N_5733);
or U12361 (N_12361,N_6405,N_5069);
nand U12362 (N_12362,N_9273,N_7149);
and U12363 (N_12363,N_6845,N_8972);
and U12364 (N_12364,N_7400,N_9704);
and U12365 (N_12365,N_9653,N_6719);
nor U12366 (N_12366,N_8300,N_8671);
nor U12367 (N_12367,N_7044,N_7525);
nand U12368 (N_12368,N_7929,N_5404);
or U12369 (N_12369,N_6193,N_7590);
or U12370 (N_12370,N_6899,N_6094);
or U12371 (N_12371,N_8345,N_9650);
or U12372 (N_12372,N_8267,N_7392);
nor U12373 (N_12373,N_8526,N_7251);
nor U12374 (N_12374,N_5160,N_8925);
nand U12375 (N_12375,N_9497,N_9929);
and U12376 (N_12376,N_6212,N_9606);
nor U12377 (N_12377,N_7867,N_5706);
nand U12378 (N_12378,N_6741,N_9712);
or U12379 (N_12379,N_7212,N_9952);
and U12380 (N_12380,N_5336,N_5686);
and U12381 (N_12381,N_5664,N_9645);
or U12382 (N_12382,N_7270,N_6729);
nor U12383 (N_12383,N_9163,N_6384);
nor U12384 (N_12384,N_5350,N_6177);
xnor U12385 (N_12385,N_8995,N_5392);
or U12386 (N_12386,N_6884,N_8216);
nand U12387 (N_12387,N_8438,N_7777);
or U12388 (N_12388,N_5740,N_7139);
or U12389 (N_12389,N_6613,N_8180);
and U12390 (N_12390,N_5135,N_6088);
xnor U12391 (N_12391,N_7413,N_5137);
or U12392 (N_12392,N_8005,N_7338);
or U12393 (N_12393,N_9207,N_9780);
xor U12394 (N_12394,N_5847,N_6256);
or U12395 (N_12395,N_7820,N_6314);
or U12396 (N_12396,N_5370,N_9900);
nor U12397 (N_12397,N_6541,N_6974);
and U12398 (N_12398,N_9976,N_9003);
nand U12399 (N_12399,N_6454,N_5017);
or U12400 (N_12400,N_5801,N_7824);
nand U12401 (N_12401,N_9228,N_6437);
and U12402 (N_12402,N_6842,N_5033);
nor U12403 (N_12403,N_5003,N_9229);
nand U12404 (N_12404,N_9462,N_6470);
and U12405 (N_12405,N_7048,N_9716);
nand U12406 (N_12406,N_7563,N_5203);
nand U12407 (N_12407,N_9019,N_8171);
nand U12408 (N_12408,N_5637,N_5848);
nand U12409 (N_12409,N_8102,N_9438);
or U12410 (N_12410,N_6272,N_5720);
or U12411 (N_12411,N_6389,N_7810);
and U12412 (N_12412,N_5326,N_9162);
xor U12413 (N_12413,N_6172,N_5157);
nand U12414 (N_12414,N_8439,N_5868);
nand U12415 (N_12415,N_5297,N_5678);
nand U12416 (N_12416,N_9039,N_8479);
nor U12417 (N_12417,N_9268,N_5452);
nand U12418 (N_12418,N_9631,N_8037);
nand U12419 (N_12419,N_8948,N_5673);
or U12420 (N_12420,N_5080,N_6035);
xor U12421 (N_12421,N_7501,N_8872);
nand U12422 (N_12422,N_5755,N_6576);
nand U12423 (N_12423,N_5662,N_7308);
nor U12424 (N_12424,N_8203,N_7521);
nand U12425 (N_12425,N_6882,N_8190);
nand U12426 (N_12426,N_8562,N_8166);
or U12427 (N_12427,N_6600,N_7380);
and U12428 (N_12428,N_7666,N_7440);
or U12429 (N_12429,N_5173,N_7385);
xnor U12430 (N_12430,N_5407,N_7341);
or U12431 (N_12431,N_5781,N_8944);
xor U12432 (N_12432,N_5804,N_8344);
and U12433 (N_12433,N_9592,N_7258);
and U12434 (N_12434,N_7950,N_7925);
nor U12435 (N_12435,N_8905,N_5159);
nand U12436 (N_12436,N_6311,N_5334);
or U12437 (N_12437,N_5357,N_9519);
nor U12438 (N_12438,N_5731,N_8169);
and U12439 (N_12439,N_8931,N_8082);
xor U12440 (N_12440,N_8577,N_9599);
or U12441 (N_12441,N_8607,N_8740);
nand U12442 (N_12442,N_8235,N_7192);
nand U12443 (N_12443,N_7932,N_9175);
and U12444 (N_12444,N_5797,N_6204);
xor U12445 (N_12445,N_7032,N_5861);
and U12446 (N_12446,N_7189,N_8026);
xnor U12447 (N_12447,N_6803,N_6869);
or U12448 (N_12448,N_5064,N_7871);
and U12449 (N_12449,N_9110,N_7075);
nand U12450 (N_12450,N_8674,N_5541);
xor U12451 (N_12451,N_6380,N_5494);
and U12452 (N_12452,N_7679,N_7201);
or U12453 (N_12453,N_5572,N_8734);
or U12454 (N_12454,N_7786,N_7245);
nor U12455 (N_12455,N_5955,N_8047);
nor U12456 (N_12456,N_7883,N_9295);
nand U12457 (N_12457,N_6951,N_8206);
nor U12458 (N_12458,N_6740,N_7462);
nor U12459 (N_12459,N_9992,N_6042);
and U12460 (N_12460,N_5477,N_7747);
nor U12461 (N_12461,N_6164,N_9874);
or U12462 (N_12462,N_9427,N_7806);
or U12463 (N_12463,N_5089,N_8295);
nand U12464 (N_12464,N_8028,N_5169);
and U12465 (N_12465,N_7477,N_8941);
nor U12466 (N_12466,N_5232,N_7711);
nor U12467 (N_12467,N_7644,N_5555);
and U12468 (N_12468,N_8289,N_8769);
or U12469 (N_12469,N_7649,N_9382);
nor U12470 (N_12470,N_5873,N_9467);
and U12471 (N_12471,N_8316,N_6396);
or U12472 (N_12472,N_6690,N_9682);
nand U12473 (N_12473,N_5595,N_9417);
xor U12474 (N_12474,N_7703,N_9074);
nor U12475 (N_12475,N_7169,N_7097);
and U12476 (N_12476,N_7601,N_9859);
nand U12477 (N_12477,N_6134,N_7343);
nand U12478 (N_12478,N_9263,N_7396);
nor U12479 (N_12479,N_9453,N_6406);
xnor U12480 (N_12480,N_5189,N_5298);
nand U12481 (N_12481,N_6859,N_9069);
and U12482 (N_12482,N_9934,N_5141);
nor U12483 (N_12483,N_5192,N_6230);
and U12484 (N_12484,N_7979,N_8857);
or U12485 (N_12485,N_8094,N_7289);
nor U12486 (N_12486,N_8834,N_5259);
xnor U12487 (N_12487,N_6883,N_9233);
and U12488 (N_12488,N_6555,N_6280);
nand U12489 (N_12489,N_9876,N_8731);
or U12490 (N_12490,N_9741,N_7074);
and U12491 (N_12491,N_9824,N_5487);
xnor U12492 (N_12492,N_8327,N_5476);
nand U12493 (N_12493,N_6962,N_9609);
and U12494 (N_12494,N_9533,N_8161);
nand U12495 (N_12495,N_5718,N_8682);
nor U12496 (N_12496,N_7906,N_5732);
or U12497 (N_12497,N_5904,N_9708);
and U12498 (N_12498,N_7104,N_5485);
nand U12499 (N_12499,N_8347,N_5457);
xnor U12500 (N_12500,N_9813,N_8972);
nand U12501 (N_12501,N_5598,N_9767);
nand U12502 (N_12502,N_7391,N_8729);
nand U12503 (N_12503,N_9298,N_8001);
nand U12504 (N_12504,N_6025,N_6514);
and U12505 (N_12505,N_8748,N_8071);
xor U12506 (N_12506,N_6498,N_8400);
xor U12507 (N_12507,N_7391,N_7990);
and U12508 (N_12508,N_5411,N_5197);
nand U12509 (N_12509,N_7461,N_8725);
nor U12510 (N_12510,N_9209,N_7650);
or U12511 (N_12511,N_8999,N_6616);
and U12512 (N_12512,N_6339,N_9677);
nor U12513 (N_12513,N_8818,N_8793);
xor U12514 (N_12514,N_6827,N_9876);
nand U12515 (N_12515,N_5738,N_9200);
and U12516 (N_12516,N_7207,N_8744);
or U12517 (N_12517,N_6617,N_6670);
nor U12518 (N_12518,N_7732,N_7615);
nand U12519 (N_12519,N_5531,N_5989);
nand U12520 (N_12520,N_9672,N_5513);
and U12521 (N_12521,N_8958,N_7515);
nor U12522 (N_12522,N_7007,N_5874);
and U12523 (N_12523,N_7981,N_7671);
xnor U12524 (N_12524,N_5029,N_8910);
nand U12525 (N_12525,N_7038,N_8502);
or U12526 (N_12526,N_5248,N_5677);
nor U12527 (N_12527,N_7898,N_9509);
nor U12528 (N_12528,N_5351,N_8020);
or U12529 (N_12529,N_7157,N_8094);
nand U12530 (N_12530,N_9798,N_5414);
nor U12531 (N_12531,N_7327,N_8938);
xor U12532 (N_12532,N_8113,N_6141);
nand U12533 (N_12533,N_8033,N_5229);
and U12534 (N_12534,N_9188,N_5827);
and U12535 (N_12535,N_9138,N_8402);
or U12536 (N_12536,N_9710,N_8681);
or U12537 (N_12537,N_5836,N_5710);
nor U12538 (N_12538,N_7871,N_8771);
nand U12539 (N_12539,N_5384,N_5141);
xnor U12540 (N_12540,N_8387,N_6037);
nor U12541 (N_12541,N_5083,N_8511);
or U12542 (N_12542,N_9656,N_5999);
and U12543 (N_12543,N_6246,N_5305);
and U12544 (N_12544,N_5199,N_8876);
nand U12545 (N_12545,N_7134,N_7166);
or U12546 (N_12546,N_7544,N_7826);
nor U12547 (N_12547,N_7974,N_5296);
xor U12548 (N_12548,N_6286,N_7304);
or U12549 (N_12549,N_9542,N_5738);
and U12550 (N_12550,N_7125,N_7106);
or U12551 (N_12551,N_7227,N_9846);
or U12552 (N_12552,N_6966,N_7045);
and U12553 (N_12553,N_7823,N_8068);
nor U12554 (N_12554,N_7097,N_5723);
and U12555 (N_12555,N_9487,N_8703);
and U12556 (N_12556,N_5124,N_6052);
or U12557 (N_12557,N_7845,N_6764);
or U12558 (N_12558,N_5027,N_9345);
or U12559 (N_12559,N_5706,N_5123);
and U12560 (N_12560,N_8058,N_8113);
nor U12561 (N_12561,N_7616,N_9561);
and U12562 (N_12562,N_8323,N_8239);
nor U12563 (N_12563,N_6880,N_6689);
nor U12564 (N_12564,N_9272,N_5517);
xor U12565 (N_12565,N_7845,N_8036);
or U12566 (N_12566,N_9960,N_9324);
or U12567 (N_12567,N_9999,N_8790);
and U12568 (N_12568,N_9579,N_7724);
nor U12569 (N_12569,N_8336,N_8450);
nand U12570 (N_12570,N_6360,N_6132);
nor U12571 (N_12571,N_5114,N_7964);
nor U12572 (N_12572,N_7173,N_6502);
nor U12573 (N_12573,N_7991,N_7438);
nand U12574 (N_12574,N_8297,N_9663);
or U12575 (N_12575,N_6828,N_7436);
or U12576 (N_12576,N_6180,N_6383);
nor U12577 (N_12577,N_5153,N_9280);
and U12578 (N_12578,N_7505,N_8850);
nor U12579 (N_12579,N_5668,N_8788);
nand U12580 (N_12580,N_5973,N_7641);
nor U12581 (N_12581,N_9427,N_8452);
nand U12582 (N_12582,N_8993,N_9758);
nand U12583 (N_12583,N_9035,N_6041);
nor U12584 (N_12584,N_6449,N_9073);
and U12585 (N_12585,N_5843,N_5247);
nor U12586 (N_12586,N_8876,N_6382);
nand U12587 (N_12587,N_9221,N_7378);
xnor U12588 (N_12588,N_8446,N_7238);
xor U12589 (N_12589,N_8550,N_5501);
nand U12590 (N_12590,N_6087,N_5339);
or U12591 (N_12591,N_7970,N_6520);
or U12592 (N_12592,N_9724,N_6256);
nor U12593 (N_12593,N_6267,N_7162);
nor U12594 (N_12594,N_6193,N_9464);
nand U12595 (N_12595,N_5992,N_9124);
nor U12596 (N_12596,N_9305,N_8543);
and U12597 (N_12597,N_7594,N_6324);
and U12598 (N_12598,N_6793,N_5923);
or U12599 (N_12599,N_5384,N_5666);
nand U12600 (N_12600,N_8650,N_9804);
nor U12601 (N_12601,N_9908,N_8928);
or U12602 (N_12602,N_5552,N_6334);
nor U12603 (N_12603,N_9091,N_5871);
and U12604 (N_12604,N_7028,N_5650);
or U12605 (N_12605,N_9550,N_6902);
nand U12606 (N_12606,N_7043,N_6270);
nor U12607 (N_12607,N_7218,N_6245);
nor U12608 (N_12608,N_6312,N_7555);
or U12609 (N_12609,N_6622,N_6808);
nor U12610 (N_12610,N_9048,N_9017);
xnor U12611 (N_12611,N_5056,N_5523);
nand U12612 (N_12612,N_7224,N_5542);
and U12613 (N_12613,N_7216,N_9251);
nand U12614 (N_12614,N_5853,N_9405);
nand U12615 (N_12615,N_8123,N_8362);
nand U12616 (N_12616,N_8139,N_6039);
and U12617 (N_12617,N_5292,N_7580);
nand U12618 (N_12618,N_6522,N_7291);
nand U12619 (N_12619,N_5864,N_9070);
nor U12620 (N_12620,N_7382,N_9592);
or U12621 (N_12621,N_5593,N_5598);
and U12622 (N_12622,N_6570,N_8935);
and U12623 (N_12623,N_9497,N_5816);
and U12624 (N_12624,N_9355,N_9579);
and U12625 (N_12625,N_6368,N_7863);
nand U12626 (N_12626,N_5507,N_9417);
nand U12627 (N_12627,N_9452,N_7520);
xor U12628 (N_12628,N_6896,N_7203);
nand U12629 (N_12629,N_7702,N_7096);
or U12630 (N_12630,N_7800,N_6883);
xor U12631 (N_12631,N_8447,N_5353);
or U12632 (N_12632,N_8135,N_6881);
nand U12633 (N_12633,N_5787,N_8381);
nand U12634 (N_12634,N_8215,N_9907);
xnor U12635 (N_12635,N_6993,N_5316);
and U12636 (N_12636,N_5288,N_9934);
nand U12637 (N_12637,N_5713,N_7738);
nand U12638 (N_12638,N_7310,N_8144);
and U12639 (N_12639,N_5612,N_8194);
or U12640 (N_12640,N_5371,N_6476);
and U12641 (N_12641,N_9360,N_5800);
or U12642 (N_12642,N_7972,N_8028);
nor U12643 (N_12643,N_5298,N_8315);
nor U12644 (N_12644,N_5003,N_7497);
and U12645 (N_12645,N_7627,N_6955);
xor U12646 (N_12646,N_6064,N_5143);
xnor U12647 (N_12647,N_9866,N_7738);
xnor U12648 (N_12648,N_9385,N_9249);
or U12649 (N_12649,N_8260,N_5469);
xnor U12650 (N_12650,N_5301,N_5138);
and U12651 (N_12651,N_7201,N_7061);
and U12652 (N_12652,N_7144,N_7326);
nor U12653 (N_12653,N_8808,N_9044);
and U12654 (N_12654,N_5680,N_8937);
xor U12655 (N_12655,N_7665,N_7798);
and U12656 (N_12656,N_8022,N_5728);
or U12657 (N_12657,N_6711,N_8375);
or U12658 (N_12658,N_9878,N_5964);
nor U12659 (N_12659,N_5502,N_7956);
xnor U12660 (N_12660,N_8611,N_9652);
nand U12661 (N_12661,N_8623,N_7313);
or U12662 (N_12662,N_8490,N_5364);
nor U12663 (N_12663,N_9629,N_7968);
and U12664 (N_12664,N_5762,N_8906);
nor U12665 (N_12665,N_9239,N_7606);
nor U12666 (N_12666,N_7050,N_9880);
nand U12667 (N_12667,N_8064,N_9544);
and U12668 (N_12668,N_7651,N_5752);
and U12669 (N_12669,N_5105,N_7914);
xor U12670 (N_12670,N_6098,N_5172);
or U12671 (N_12671,N_5985,N_6050);
or U12672 (N_12672,N_9893,N_7352);
nand U12673 (N_12673,N_8905,N_7995);
and U12674 (N_12674,N_8617,N_5584);
nand U12675 (N_12675,N_6965,N_9320);
nand U12676 (N_12676,N_8927,N_6665);
and U12677 (N_12677,N_8175,N_6156);
and U12678 (N_12678,N_6508,N_8918);
and U12679 (N_12679,N_9817,N_9956);
xor U12680 (N_12680,N_7850,N_8328);
or U12681 (N_12681,N_9490,N_7844);
or U12682 (N_12682,N_6853,N_7351);
and U12683 (N_12683,N_5435,N_8179);
or U12684 (N_12684,N_9053,N_9113);
and U12685 (N_12685,N_9402,N_7379);
and U12686 (N_12686,N_8676,N_9274);
xnor U12687 (N_12687,N_5341,N_8890);
xnor U12688 (N_12688,N_8357,N_7210);
or U12689 (N_12689,N_6803,N_9952);
nor U12690 (N_12690,N_9386,N_7200);
and U12691 (N_12691,N_8349,N_6832);
and U12692 (N_12692,N_8191,N_5012);
nand U12693 (N_12693,N_7745,N_8599);
nand U12694 (N_12694,N_8520,N_9598);
and U12695 (N_12695,N_6645,N_5607);
nand U12696 (N_12696,N_5788,N_5414);
or U12697 (N_12697,N_7943,N_8947);
nand U12698 (N_12698,N_8925,N_5649);
nor U12699 (N_12699,N_5354,N_8343);
nor U12700 (N_12700,N_8297,N_6871);
and U12701 (N_12701,N_6888,N_7049);
and U12702 (N_12702,N_7222,N_8048);
or U12703 (N_12703,N_6817,N_6703);
nand U12704 (N_12704,N_9655,N_7769);
and U12705 (N_12705,N_5117,N_6227);
or U12706 (N_12706,N_8365,N_5327);
nand U12707 (N_12707,N_5123,N_6674);
nor U12708 (N_12708,N_9621,N_8767);
and U12709 (N_12709,N_8030,N_7909);
and U12710 (N_12710,N_5530,N_6707);
nor U12711 (N_12711,N_6420,N_8848);
nand U12712 (N_12712,N_9891,N_8675);
or U12713 (N_12713,N_5043,N_5113);
xnor U12714 (N_12714,N_9370,N_9393);
xnor U12715 (N_12715,N_6405,N_8271);
or U12716 (N_12716,N_9261,N_5189);
nand U12717 (N_12717,N_5163,N_8508);
and U12718 (N_12718,N_9281,N_5620);
nand U12719 (N_12719,N_5258,N_8295);
nor U12720 (N_12720,N_5551,N_7929);
and U12721 (N_12721,N_9599,N_7984);
or U12722 (N_12722,N_5323,N_5885);
nor U12723 (N_12723,N_9393,N_9968);
and U12724 (N_12724,N_5420,N_8706);
xnor U12725 (N_12725,N_9671,N_8421);
nor U12726 (N_12726,N_9664,N_6895);
xnor U12727 (N_12727,N_9111,N_6344);
and U12728 (N_12728,N_7797,N_9281);
nand U12729 (N_12729,N_6139,N_9494);
and U12730 (N_12730,N_8831,N_8794);
nor U12731 (N_12731,N_8362,N_8986);
xnor U12732 (N_12732,N_9956,N_7050);
nand U12733 (N_12733,N_7153,N_6257);
or U12734 (N_12734,N_8568,N_7202);
nand U12735 (N_12735,N_7601,N_5908);
or U12736 (N_12736,N_8044,N_5189);
or U12737 (N_12737,N_7792,N_5844);
nor U12738 (N_12738,N_8691,N_9290);
and U12739 (N_12739,N_5520,N_8518);
xor U12740 (N_12740,N_7059,N_7411);
and U12741 (N_12741,N_6663,N_9865);
xor U12742 (N_12742,N_8764,N_8463);
or U12743 (N_12743,N_7046,N_5646);
and U12744 (N_12744,N_8110,N_8132);
nand U12745 (N_12745,N_6712,N_6699);
or U12746 (N_12746,N_8217,N_7486);
and U12747 (N_12747,N_9546,N_9583);
and U12748 (N_12748,N_9449,N_8783);
or U12749 (N_12749,N_9749,N_7620);
nand U12750 (N_12750,N_5559,N_7918);
xor U12751 (N_12751,N_9848,N_9610);
nor U12752 (N_12752,N_6894,N_7561);
and U12753 (N_12753,N_8180,N_5108);
nand U12754 (N_12754,N_6433,N_7162);
and U12755 (N_12755,N_8054,N_5386);
xor U12756 (N_12756,N_7995,N_8660);
nor U12757 (N_12757,N_7877,N_5153);
and U12758 (N_12758,N_9557,N_7924);
or U12759 (N_12759,N_5604,N_7560);
or U12760 (N_12760,N_8445,N_7698);
or U12761 (N_12761,N_9253,N_9356);
and U12762 (N_12762,N_5425,N_5781);
nor U12763 (N_12763,N_9754,N_8535);
xor U12764 (N_12764,N_5877,N_5515);
nor U12765 (N_12765,N_8571,N_6834);
nor U12766 (N_12766,N_6421,N_9612);
and U12767 (N_12767,N_6910,N_9077);
xnor U12768 (N_12768,N_6565,N_5718);
and U12769 (N_12769,N_8643,N_8341);
and U12770 (N_12770,N_9611,N_9597);
or U12771 (N_12771,N_8116,N_6407);
nand U12772 (N_12772,N_5130,N_5375);
or U12773 (N_12773,N_7420,N_7325);
xnor U12774 (N_12774,N_8368,N_5011);
and U12775 (N_12775,N_5165,N_8811);
nand U12776 (N_12776,N_5815,N_8880);
xor U12777 (N_12777,N_5733,N_6220);
nand U12778 (N_12778,N_5608,N_9536);
or U12779 (N_12779,N_5069,N_7715);
nor U12780 (N_12780,N_9327,N_5414);
or U12781 (N_12781,N_7673,N_9558);
or U12782 (N_12782,N_6434,N_9205);
nand U12783 (N_12783,N_7104,N_6391);
and U12784 (N_12784,N_8676,N_5064);
nor U12785 (N_12785,N_9424,N_8851);
or U12786 (N_12786,N_9679,N_5565);
and U12787 (N_12787,N_6993,N_8774);
nand U12788 (N_12788,N_6761,N_9291);
nand U12789 (N_12789,N_9445,N_6773);
nand U12790 (N_12790,N_6877,N_9004);
nor U12791 (N_12791,N_6789,N_5246);
xnor U12792 (N_12792,N_9398,N_5210);
and U12793 (N_12793,N_6119,N_8490);
or U12794 (N_12794,N_8545,N_9278);
xor U12795 (N_12795,N_8401,N_8275);
or U12796 (N_12796,N_5362,N_7648);
nand U12797 (N_12797,N_9877,N_8483);
and U12798 (N_12798,N_9283,N_6185);
and U12799 (N_12799,N_7908,N_9115);
and U12800 (N_12800,N_6962,N_7023);
nand U12801 (N_12801,N_7318,N_6689);
or U12802 (N_12802,N_6648,N_9667);
or U12803 (N_12803,N_8732,N_6005);
and U12804 (N_12804,N_7799,N_6962);
or U12805 (N_12805,N_5711,N_7729);
or U12806 (N_12806,N_7359,N_9332);
and U12807 (N_12807,N_5079,N_8066);
nor U12808 (N_12808,N_6398,N_6861);
or U12809 (N_12809,N_9725,N_9568);
and U12810 (N_12810,N_8605,N_5662);
or U12811 (N_12811,N_5416,N_9872);
nor U12812 (N_12812,N_7633,N_5059);
or U12813 (N_12813,N_8734,N_5837);
or U12814 (N_12814,N_8743,N_6883);
or U12815 (N_12815,N_7737,N_7768);
or U12816 (N_12816,N_6210,N_8966);
and U12817 (N_12817,N_5992,N_6819);
or U12818 (N_12818,N_5864,N_8000);
nor U12819 (N_12819,N_7896,N_8632);
xor U12820 (N_12820,N_7212,N_9530);
or U12821 (N_12821,N_5727,N_9682);
xnor U12822 (N_12822,N_7879,N_8689);
nor U12823 (N_12823,N_5876,N_6633);
and U12824 (N_12824,N_8590,N_8629);
nor U12825 (N_12825,N_8356,N_7775);
or U12826 (N_12826,N_5377,N_9497);
and U12827 (N_12827,N_7240,N_6670);
nand U12828 (N_12828,N_5556,N_6177);
and U12829 (N_12829,N_7936,N_6890);
nor U12830 (N_12830,N_9962,N_7641);
and U12831 (N_12831,N_7466,N_5891);
or U12832 (N_12832,N_8839,N_8539);
nor U12833 (N_12833,N_9141,N_9003);
or U12834 (N_12834,N_8036,N_9059);
xor U12835 (N_12835,N_8861,N_7933);
or U12836 (N_12836,N_7463,N_5471);
and U12837 (N_12837,N_7619,N_5182);
or U12838 (N_12838,N_8063,N_7044);
nand U12839 (N_12839,N_7645,N_9119);
and U12840 (N_12840,N_8782,N_8592);
nor U12841 (N_12841,N_6013,N_9338);
xnor U12842 (N_12842,N_9958,N_6053);
or U12843 (N_12843,N_5960,N_6990);
and U12844 (N_12844,N_5276,N_8318);
and U12845 (N_12845,N_9073,N_7354);
and U12846 (N_12846,N_7543,N_8337);
nor U12847 (N_12847,N_5695,N_7882);
nor U12848 (N_12848,N_9800,N_5967);
and U12849 (N_12849,N_8868,N_6711);
and U12850 (N_12850,N_9040,N_6742);
and U12851 (N_12851,N_7373,N_5825);
or U12852 (N_12852,N_6193,N_6949);
and U12853 (N_12853,N_8776,N_6491);
or U12854 (N_12854,N_9634,N_9515);
and U12855 (N_12855,N_5745,N_5928);
or U12856 (N_12856,N_9876,N_8617);
nor U12857 (N_12857,N_6649,N_9632);
and U12858 (N_12858,N_8496,N_9156);
and U12859 (N_12859,N_9786,N_9764);
xnor U12860 (N_12860,N_5857,N_9495);
and U12861 (N_12861,N_6114,N_9490);
nor U12862 (N_12862,N_6412,N_9809);
and U12863 (N_12863,N_5600,N_7355);
nand U12864 (N_12864,N_7914,N_6810);
or U12865 (N_12865,N_9108,N_9510);
or U12866 (N_12866,N_8502,N_7522);
and U12867 (N_12867,N_9103,N_6292);
nor U12868 (N_12868,N_5212,N_9294);
nor U12869 (N_12869,N_9028,N_7411);
xnor U12870 (N_12870,N_7248,N_8191);
nand U12871 (N_12871,N_9836,N_6542);
or U12872 (N_12872,N_5259,N_5638);
or U12873 (N_12873,N_9984,N_5018);
nor U12874 (N_12874,N_6926,N_5406);
nor U12875 (N_12875,N_8137,N_5684);
nand U12876 (N_12876,N_5426,N_6890);
xnor U12877 (N_12877,N_9369,N_5934);
nand U12878 (N_12878,N_9388,N_7265);
nand U12879 (N_12879,N_5370,N_5845);
and U12880 (N_12880,N_6910,N_6922);
nand U12881 (N_12881,N_5978,N_9003);
nor U12882 (N_12882,N_5140,N_9427);
and U12883 (N_12883,N_9821,N_5729);
nand U12884 (N_12884,N_5896,N_9362);
and U12885 (N_12885,N_6055,N_8052);
xnor U12886 (N_12886,N_5191,N_6629);
nand U12887 (N_12887,N_6594,N_5242);
or U12888 (N_12888,N_8146,N_6697);
or U12889 (N_12889,N_8804,N_8985);
nand U12890 (N_12890,N_7704,N_5554);
and U12891 (N_12891,N_9713,N_9185);
or U12892 (N_12892,N_7650,N_5979);
or U12893 (N_12893,N_5388,N_6175);
xnor U12894 (N_12894,N_9837,N_8928);
or U12895 (N_12895,N_9382,N_7347);
xnor U12896 (N_12896,N_6349,N_8755);
or U12897 (N_12897,N_7568,N_9775);
nor U12898 (N_12898,N_9570,N_7077);
nand U12899 (N_12899,N_9220,N_9212);
or U12900 (N_12900,N_7848,N_9507);
nand U12901 (N_12901,N_8544,N_5407);
or U12902 (N_12902,N_9359,N_8532);
and U12903 (N_12903,N_6695,N_8978);
nand U12904 (N_12904,N_8913,N_9573);
nand U12905 (N_12905,N_7674,N_7251);
nor U12906 (N_12906,N_5416,N_7654);
nor U12907 (N_12907,N_9560,N_6357);
nor U12908 (N_12908,N_9582,N_9457);
nor U12909 (N_12909,N_8029,N_8469);
nand U12910 (N_12910,N_7497,N_7711);
nor U12911 (N_12911,N_8502,N_9384);
nand U12912 (N_12912,N_9236,N_5375);
nand U12913 (N_12913,N_7488,N_5750);
nor U12914 (N_12914,N_8299,N_6233);
or U12915 (N_12915,N_9940,N_8488);
nand U12916 (N_12916,N_7223,N_5006);
xor U12917 (N_12917,N_6827,N_5901);
or U12918 (N_12918,N_8681,N_8743);
nor U12919 (N_12919,N_5817,N_9563);
nand U12920 (N_12920,N_5006,N_8778);
and U12921 (N_12921,N_7088,N_5959);
or U12922 (N_12922,N_7075,N_6803);
or U12923 (N_12923,N_8355,N_7558);
xor U12924 (N_12924,N_8798,N_9956);
or U12925 (N_12925,N_8171,N_6273);
or U12926 (N_12926,N_9524,N_8457);
or U12927 (N_12927,N_7603,N_7540);
nand U12928 (N_12928,N_5271,N_5564);
nor U12929 (N_12929,N_8647,N_7193);
xor U12930 (N_12930,N_5596,N_5333);
nand U12931 (N_12931,N_9117,N_9518);
and U12932 (N_12932,N_5336,N_9875);
nand U12933 (N_12933,N_9456,N_6299);
xnor U12934 (N_12934,N_6943,N_9427);
or U12935 (N_12935,N_7083,N_8090);
and U12936 (N_12936,N_7002,N_8301);
and U12937 (N_12937,N_8446,N_5191);
or U12938 (N_12938,N_8170,N_6000);
or U12939 (N_12939,N_7436,N_9271);
nor U12940 (N_12940,N_8379,N_5555);
nand U12941 (N_12941,N_5016,N_5051);
or U12942 (N_12942,N_6063,N_9380);
xnor U12943 (N_12943,N_9829,N_6005);
or U12944 (N_12944,N_5727,N_6201);
or U12945 (N_12945,N_6520,N_7775);
nand U12946 (N_12946,N_7445,N_6048);
and U12947 (N_12947,N_6795,N_6914);
or U12948 (N_12948,N_9976,N_9200);
and U12949 (N_12949,N_7739,N_8268);
xnor U12950 (N_12950,N_7977,N_9917);
nor U12951 (N_12951,N_7046,N_8518);
and U12952 (N_12952,N_6152,N_6149);
nand U12953 (N_12953,N_9806,N_5561);
nand U12954 (N_12954,N_5654,N_5719);
and U12955 (N_12955,N_7421,N_6711);
or U12956 (N_12956,N_7103,N_9832);
nor U12957 (N_12957,N_6258,N_6684);
nand U12958 (N_12958,N_6119,N_7916);
or U12959 (N_12959,N_8613,N_8752);
and U12960 (N_12960,N_8298,N_8540);
and U12961 (N_12961,N_5636,N_9185);
and U12962 (N_12962,N_9863,N_5320);
nor U12963 (N_12963,N_5049,N_9983);
and U12964 (N_12964,N_6285,N_5276);
xnor U12965 (N_12965,N_5301,N_9654);
nand U12966 (N_12966,N_9455,N_8636);
or U12967 (N_12967,N_9591,N_8172);
nor U12968 (N_12968,N_8658,N_5095);
nand U12969 (N_12969,N_5234,N_8875);
and U12970 (N_12970,N_6395,N_6959);
and U12971 (N_12971,N_7420,N_6952);
and U12972 (N_12972,N_7915,N_6403);
and U12973 (N_12973,N_9317,N_5815);
nor U12974 (N_12974,N_7979,N_7268);
nand U12975 (N_12975,N_6265,N_6536);
nand U12976 (N_12976,N_7751,N_9396);
nand U12977 (N_12977,N_9620,N_6190);
and U12978 (N_12978,N_5908,N_7100);
xor U12979 (N_12979,N_8195,N_8662);
and U12980 (N_12980,N_9895,N_5225);
and U12981 (N_12981,N_7508,N_5167);
nand U12982 (N_12982,N_5658,N_5606);
or U12983 (N_12983,N_9503,N_5393);
nand U12984 (N_12984,N_7584,N_7860);
and U12985 (N_12985,N_8952,N_9593);
and U12986 (N_12986,N_5575,N_9309);
nor U12987 (N_12987,N_5571,N_5083);
or U12988 (N_12988,N_6769,N_6713);
nor U12989 (N_12989,N_9045,N_8803);
or U12990 (N_12990,N_6303,N_8520);
and U12991 (N_12991,N_7550,N_9372);
and U12992 (N_12992,N_6816,N_9395);
nand U12993 (N_12993,N_7719,N_5445);
and U12994 (N_12994,N_8828,N_6991);
or U12995 (N_12995,N_9554,N_9531);
or U12996 (N_12996,N_6118,N_8408);
or U12997 (N_12997,N_6592,N_9035);
or U12998 (N_12998,N_7162,N_7917);
or U12999 (N_12999,N_5045,N_9218);
xnor U13000 (N_13000,N_9110,N_5493);
xnor U13001 (N_13001,N_7215,N_9217);
xnor U13002 (N_13002,N_7046,N_5495);
or U13003 (N_13003,N_7127,N_8635);
nor U13004 (N_13004,N_6855,N_9035);
and U13005 (N_13005,N_8379,N_8782);
nand U13006 (N_13006,N_8367,N_6495);
xnor U13007 (N_13007,N_7095,N_5179);
nand U13008 (N_13008,N_5039,N_5120);
xnor U13009 (N_13009,N_5083,N_6509);
or U13010 (N_13010,N_7904,N_9902);
nand U13011 (N_13011,N_9920,N_8158);
nor U13012 (N_13012,N_6084,N_7031);
nor U13013 (N_13013,N_7413,N_7739);
or U13014 (N_13014,N_8897,N_6463);
nand U13015 (N_13015,N_6156,N_8631);
nor U13016 (N_13016,N_5833,N_7614);
nor U13017 (N_13017,N_9880,N_9349);
or U13018 (N_13018,N_9268,N_7842);
nand U13019 (N_13019,N_5674,N_9905);
or U13020 (N_13020,N_9505,N_6686);
and U13021 (N_13021,N_8147,N_8050);
nand U13022 (N_13022,N_9316,N_5447);
nand U13023 (N_13023,N_5965,N_7440);
and U13024 (N_13024,N_7441,N_6203);
or U13025 (N_13025,N_8275,N_5157);
nand U13026 (N_13026,N_6670,N_7289);
and U13027 (N_13027,N_9558,N_7354);
xor U13028 (N_13028,N_6408,N_8722);
nor U13029 (N_13029,N_5583,N_8652);
nand U13030 (N_13030,N_8316,N_7318);
and U13031 (N_13031,N_5332,N_9098);
or U13032 (N_13032,N_7488,N_9835);
or U13033 (N_13033,N_6256,N_9113);
xor U13034 (N_13034,N_5309,N_7677);
and U13035 (N_13035,N_7760,N_7238);
nor U13036 (N_13036,N_5212,N_5115);
nand U13037 (N_13037,N_9190,N_6568);
and U13038 (N_13038,N_7406,N_5743);
or U13039 (N_13039,N_9803,N_5495);
nor U13040 (N_13040,N_9018,N_6116);
nand U13041 (N_13041,N_7627,N_5806);
nand U13042 (N_13042,N_8202,N_8635);
and U13043 (N_13043,N_6333,N_9857);
or U13044 (N_13044,N_6539,N_9160);
nor U13045 (N_13045,N_5051,N_8172);
nand U13046 (N_13046,N_7132,N_5999);
or U13047 (N_13047,N_5058,N_7087);
xnor U13048 (N_13048,N_7908,N_7180);
nand U13049 (N_13049,N_9140,N_9755);
or U13050 (N_13050,N_8498,N_6497);
and U13051 (N_13051,N_9295,N_8287);
nand U13052 (N_13052,N_6754,N_6215);
or U13053 (N_13053,N_8318,N_7861);
or U13054 (N_13054,N_6402,N_6239);
and U13055 (N_13055,N_6424,N_9582);
nor U13056 (N_13056,N_6581,N_8720);
and U13057 (N_13057,N_5411,N_9097);
and U13058 (N_13058,N_8016,N_8765);
and U13059 (N_13059,N_9280,N_9152);
nand U13060 (N_13060,N_7333,N_7870);
or U13061 (N_13061,N_9891,N_5756);
and U13062 (N_13062,N_9010,N_7600);
xor U13063 (N_13063,N_7711,N_8978);
nand U13064 (N_13064,N_9454,N_7167);
and U13065 (N_13065,N_5066,N_8498);
nor U13066 (N_13066,N_7002,N_7861);
and U13067 (N_13067,N_6490,N_5802);
and U13068 (N_13068,N_6024,N_9987);
or U13069 (N_13069,N_8527,N_8404);
and U13070 (N_13070,N_8457,N_9334);
xor U13071 (N_13071,N_6704,N_9166);
nor U13072 (N_13072,N_9776,N_6879);
nand U13073 (N_13073,N_7896,N_5511);
and U13074 (N_13074,N_6724,N_8082);
nand U13075 (N_13075,N_6879,N_8350);
and U13076 (N_13076,N_9301,N_9530);
nor U13077 (N_13077,N_7688,N_9949);
nand U13078 (N_13078,N_7603,N_8624);
and U13079 (N_13079,N_8940,N_9360);
nor U13080 (N_13080,N_9042,N_9592);
nor U13081 (N_13081,N_6328,N_7621);
or U13082 (N_13082,N_5574,N_7634);
nor U13083 (N_13083,N_7591,N_7848);
nand U13084 (N_13084,N_6805,N_8001);
and U13085 (N_13085,N_7016,N_5063);
or U13086 (N_13086,N_5009,N_8005);
nor U13087 (N_13087,N_8118,N_7257);
or U13088 (N_13088,N_5617,N_8652);
nand U13089 (N_13089,N_7620,N_5243);
nand U13090 (N_13090,N_5871,N_9070);
nand U13091 (N_13091,N_7179,N_5610);
or U13092 (N_13092,N_5377,N_5278);
and U13093 (N_13093,N_6331,N_5971);
nand U13094 (N_13094,N_7478,N_8792);
nor U13095 (N_13095,N_7571,N_5619);
nor U13096 (N_13096,N_5490,N_7772);
nand U13097 (N_13097,N_7558,N_5945);
and U13098 (N_13098,N_6286,N_7756);
or U13099 (N_13099,N_7578,N_9301);
and U13100 (N_13100,N_9939,N_9340);
nor U13101 (N_13101,N_8896,N_9255);
nand U13102 (N_13102,N_8686,N_9348);
xor U13103 (N_13103,N_6679,N_9479);
and U13104 (N_13104,N_5891,N_8811);
nand U13105 (N_13105,N_7898,N_9092);
xor U13106 (N_13106,N_9556,N_7875);
nand U13107 (N_13107,N_9732,N_7387);
nand U13108 (N_13108,N_5655,N_9123);
or U13109 (N_13109,N_9695,N_9208);
nand U13110 (N_13110,N_6202,N_8582);
nand U13111 (N_13111,N_9379,N_5726);
nand U13112 (N_13112,N_6372,N_7716);
nor U13113 (N_13113,N_6910,N_5668);
nand U13114 (N_13114,N_8000,N_6426);
and U13115 (N_13115,N_9046,N_9819);
or U13116 (N_13116,N_7406,N_7087);
and U13117 (N_13117,N_7882,N_8857);
or U13118 (N_13118,N_5899,N_5264);
and U13119 (N_13119,N_7842,N_9280);
xor U13120 (N_13120,N_6382,N_9124);
nor U13121 (N_13121,N_8324,N_5825);
and U13122 (N_13122,N_6834,N_8939);
nor U13123 (N_13123,N_6075,N_6765);
or U13124 (N_13124,N_9556,N_7663);
xnor U13125 (N_13125,N_5142,N_7666);
or U13126 (N_13126,N_6697,N_7665);
or U13127 (N_13127,N_6963,N_8051);
and U13128 (N_13128,N_6569,N_5382);
nand U13129 (N_13129,N_9089,N_9645);
and U13130 (N_13130,N_8251,N_7325);
nor U13131 (N_13131,N_8413,N_6933);
nand U13132 (N_13132,N_7321,N_8633);
and U13133 (N_13133,N_8679,N_9338);
nor U13134 (N_13134,N_6449,N_5772);
or U13135 (N_13135,N_6513,N_9156);
or U13136 (N_13136,N_9319,N_6756);
nand U13137 (N_13137,N_8077,N_7793);
nor U13138 (N_13138,N_5314,N_8741);
and U13139 (N_13139,N_7609,N_7702);
nand U13140 (N_13140,N_8882,N_7251);
and U13141 (N_13141,N_6099,N_6117);
and U13142 (N_13142,N_9940,N_9435);
nand U13143 (N_13143,N_5778,N_7826);
xor U13144 (N_13144,N_8594,N_8570);
xnor U13145 (N_13145,N_9816,N_8901);
nand U13146 (N_13146,N_9460,N_6656);
nand U13147 (N_13147,N_7686,N_5817);
and U13148 (N_13148,N_5134,N_6855);
or U13149 (N_13149,N_7653,N_7046);
or U13150 (N_13150,N_6439,N_7925);
and U13151 (N_13151,N_9391,N_9502);
nor U13152 (N_13152,N_9183,N_6651);
nand U13153 (N_13153,N_5693,N_6856);
xor U13154 (N_13154,N_7367,N_6724);
nand U13155 (N_13155,N_6110,N_8996);
nand U13156 (N_13156,N_6528,N_9753);
nand U13157 (N_13157,N_6567,N_9471);
or U13158 (N_13158,N_9626,N_6892);
nand U13159 (N_13159,N_5729,N_7460);
or U13160 (N_13160,N_9366,N_9725);
nor U13161 (N_13161,N_7749,N_8135);
and U13162 (N_13162,N_9045,N_6665);
nand U13163 (N_13163,N_7324,N_9364);
and U13164 (N_13164,N_5687,N_9540);
nor U13165 (N_13165,N_5770,N_6912);
or U13166 (N_13166,N_6416,N_8288);
nand U13167 (N_13167,N_5071,N_5371);
xnor U13168 (N_13168,N_7543,N_8853);
nor U13169 (N_13169,N_6810,N_8537);
or U13170 (N_13170,N_7467,N_5617);
nand U13171 (N_13171,N_8880,N_9040);
nand U13172 (N_13172,N_6892,N_7665);
nand U13173 (N_13173,N_7987,N_7432);
or U13174 (N_13174,N_9980,N_7195);
and U13175 (N_13175,N_9446,N_8518);
nand U13176 (N_13176,N_9795,N_9812);
nor U13177 (N_13177,N_8628,N_7229);
or U13178 (N_13178,N_5516,N_6618);
nand U13179 (N_13179,N_8906,N_5342);
nand U13180 (N_13180,N_6873,N_6370);
nor U13181 (N_13181,N_8396,N_8758);
nor U13182 (N_13182,N_5298,N_8500);
nor U13183 (N_13183,N_9644,N_5141);
or U13184 (N_13184,N_5641,N_8126);
nor U13185 (N_13185,N_7290,N_6126);
nor U13186 (N_13186,N_7291,N_8888);
and U13187 (N_13187,N_6751,N_6724);
or U13188 (N_13188,N_9741,N_8084);
xor U13189 (N_13189,N_8076,N_7417);
nand U13190 (N_13190,N_8917,N_9016);
nor U13191 (N_13191,N_7508,N_9766);
or U13192 (N_13192,N_6366,N_5309);
and U13193 (N_13193,N_9014,N_8576);
xor U13194 (N_13194,N_8587,N_6457);
nor U13195 (N_13195,N_6735,N_7654);
nand U13196 (N_13196,N_5649,N_8426);
or U13197 (N_13197,N_7282,N_5076);
nand U13198 (N_13198,N_8782,N_9837);
xnor U13199 (N_13199,N_6101,N_6543);
nor U13200 (N_13200,N_6360,N_7022);
xnor U13201 (N_13201,N_5932,N_5364);
nand U13202 (N_13202,N_5153,N_5897);
nor U13203 (N_13203,N_8794,N_9139);
nor U13204 (N_13204,N_8985,N_8186);
or U13205 (N_13205,N_9234,N_7637);
nor U13206 (N_13206,N_5832,N_6393);
nand U13207 (N_13207,N_9690,N_5126);
nand U13208 (N_13208,N_9760,N_5216);
or U13209 (N_13209,N_9479,N_6746);
nand U13210 (N_13210,N_6948,N_6541);
xnor U13211 (N_13211,N_6447,N_6015);
and U13212 (N_13212,N_5962,N_5781);
or U13213 (N_13213,N_8796,N_9710);
or U13214 (N_13214,N_8649,N_5890);
nor U13215 (N_13215,N_7945,N_7720);
or U13216 (N_13216,N_7098,N_7577);
or U13217 (N_13217,N_6309,N_9728);
nand U13218 (N_13218,N_9933,N_6017);
and U13219 (N_13219,N_6541,N_6429);
or U13220 (N_13220,N_8877,N_6287);
nor U13221 (N_13221,N_6358,N_5168);
and U13222 (N_13222,N_7563,N_5775);
or U13223 (N_13223,N_9163,N_7394);
or U13224 (N_13224,N_7753,N_5319);
xor U13225 (N_13225,N_5356,N_5748);
or U13226 (N_13226,N_8651,N_9642);
nor U13227 (N_13227,N_8927,N_5040);
and U13228 (N_13228,N_9888,N_5847);
or U13229 (N_13229,N_9482,N_8778);
nor U13230 (N_13230,N_5504,N_7515);
or U13231 (N_13231,N_8460,N_7781);
or U13232 (N_13232,N_9115,N_8675);
nand U13233 (N_13233,N_7782,N_7623);
nor U13234 (N_13234,N_8111,N_6511);
and U13235 (N_13235,N_5096,N_5385);
nor U13236 (N_13236,N_8795,N_9840);
nand U13237 (N_13237,N_8483,N_9166);
or U13238 (N_13238,N_9198,N_7103);
or U13239 (N_13239,N_7883,N_6573);
and U13240 (N_13240,N_9355,N_6046);
nand U13241 (N_13241,N_8409,N_6123);
xor U13242 (N_13242,N_6930,N_9892);
or U13243 (N_13243,N_6780,N_9294);
nor U13244 (N_13244,N_5769,N_5553);
nand U13245 (N_13245,N_7389,N_5083);
nand U13246 (N_13246,N_7014,N_6004);
nand U13247 (N_13247,N_5297,N_8747);
nor U13248 (N_13248,N_6551,N_5119);
xor U13249 (N_13249,N_7649,N_5733);
and U13250 (N_13250,N_9109,N_6814);
or U13251 (N_13251,N_8343,N_7389);
nor U13252 (N_13252,N_8218,N_7940);
nor U13253 (N_13253,N_7037,N_5377);
or U13254 (N_13254,N_9803,N_5944);
or U13255 (N_13255,N_8025,N_9239);
and U13256 (N_13256,N_9306,N_5877);
xnor U13257 (N_13257,N_9886,N_5182);
or U13258 (N_13258,N_8283,N_7314);
nand U13259 (N_13259,N_8749,N_7571);
and U13260 (N_13260,N_5860,N_6034);
nor U13261 (N_13261,N_9124,N_8469);
or U13262 (N_13262,N_5252,N_5819);
nor U13263 (N_13263,N_5929,N_6250);
or U13264 (N_13264,N_9005,N_9990);
nand U13265 (N_13265,N_9948,N_7942);
nor U13266 (N_13266,N_9523,N_9285);
and U13267 (N_13267,N_5663,N_7095);
nor U13268 (N_13268,N_5315,N_7805);
nor U13269 (N_13269,N_5765,N_9340);
and U13270 (N_13270,N_8592,N_5253);
nand U13271 (N_13271,N_7956,N_8964);
nand U13272 (N_13272,N_7282,N_6783);
and U13273 (N_13273,N_7636,N_8446);
or U13274 (N_13274,N_7949,N_8029);
or U13275 (N_13275,N_7374,N_7325);
nand U13276 (N_13276,N_5855,N_8341);
or U13277 (N_13277,N_6443,N_5842);
or U13278 (N_13278,N_5884,N_9716);
or U13279 (N_13279,N_8053,N_8434);
nor U13280 (N_13280,N_6953,N_5740);
or U13281 (N_13281,N_6126,N_8886);
or U13282 (N_13282,N_7995,N_9775);
and U13283 (N_13283,N_8060,N_6757);
nor U13284 (N_13284,N_5285,N_8864);
xor U13285 (N_13285,N_8482,N_6530);
xnor U13286 (N_13286,N_5278,N_5000);
xor U13287 (N_13287,N_5084,N_8191);
or U13288 (N_13288,N_7021,N_7683);
and U13289 (N_13289,N_9577,N_8662);
or U13290 (N_13290,N_8301,N_9410);
or U13291 (N_13291,N_9971,N_5129);
or U13292 (N_13292,N_5767,N_8609);
nor U13293 (N_13293,N_9554,N_8438);
and U13294 (N_13294,N_8009,N_7305);
or U13295 (N_13295,N_8160,N_7131);
nand U13296 (N_13296,N_8982,N_7591);
nor U13297 (N_13297,N_9692,N_5980);
nand U13298 (N_13298,N_5613,N_8979);
or U13299 (N_13299,N_5705,N_8815);
or U13300 (N_13300,N_8234,N_9079);
nand U13301 (N_13301,N_5021,N_9287);
or U13302 (N_13302,N_9352,N_9815);
nor U13303 (N_13303,N_5341,N_7515);
nor U13304 (N_13304,N_8801,N_6949);
and U13305 (N_13305,N_5744,N_5584);
nor U13306 (N_13306,N_9866,N_9094);
and U13307 (N_13307,N_8495,N_7688);
and U13308 (N_13308,N_5246,N_5315);
xnor U13309 (N_13309,N_7539,N_9434);
xor U13310 (N_13310,N_9993,N_7080);
nor U13311 (N_13311,N_6788,N_5677);
nor U13312 (N_13312,N_6040,N_9364);
and U13313 (N_13313,N_9181,N_6700);
xnor U13314 (N_13314,N_6885,N_5947);
nand U13315 (N_13315,N_8515,N_9915);
nor U13316 (N_13316,N_9753,N_5535);
xnor U13317 (N_13317,N_9040,N_5902);
or U13318 (N_13318,N_5422,N_6182);
xnor U13319 (N_13319,N_7583,N_5557);
or U13320 (N_13320,N_7784,N_6777);
or U13321 (N_13321,N_5286,N_9803);
and U13322 (N_13322,N_5770,N_7880);
nand U13323 (N_13323,N_6837,N_7915);
nand U13324 (N_13324,N_9355,N_5663);
or U13325 (N_13325,N_5776,N_7939);
and U13326 (N_13326,N_7146,N_6994);
and U13327 (N_13327,N_6236,N_6882);
nor U13328 (N_13328,N_9664,N_8217);
or U13329 (N_13329,N_6666,N_5167);
xnor U13330 (N_13330,N_9663,N_9277);
nand U13331 (N_13331,N_7502,N_9142);
nor U13332 (N_13332,N_6364,N_7376);
or U13333 (N_13333,N_6428,N_7440);
xor U13334 (N_13334,N_6229,N_6142);
and U13335 (N_13335,N_6690,N_8454);
nor U13336 (N_13336,N_6882,N_5123);
or U13337 (N_13337,N_8251,N_9344);
nand U13338 (N_13338,N_7258,N_5227);
or U13339 (N_13339,N_8354,N_5604);
and U13340 (N_13340,N_9437,N_7773);
or U13341 (N_13341,N_5341,N_9960);
xor U13342 (N_13342,N_5117,N_5630);
nor U13343 (N_13343,N_9585,N_6286);
nor U13344 (N_13344,N_7599,N_8916);
nand U13345 (N_13345,N_8403,N_7413);
and U13346 (N_13346,N_7976,N_6624);
and U13347 (N_13347,N_7992,N_9943);
xor U13348 (N_13348,N_6696,N_8626);
and U13349 (N_13349,N_8892,N_8026);
nand U13350 (N_13350,N_5280,N_5282);
or U13351 (N_13351,N_6497,N_6405);
and U13352 (N_13352,N_6085,N_8689);
xor U13353 (N_13353,N_6672,N_6831);
nand U13354 (N_13354,N_9829,N_8961);
nor U13355 (N_13355,N_7977,N_6850);
nor U13356 (N_13356,N_5557,N_8588);
or U13357 (N_13357,N_9564,N_5486);
nor U13358 (N_13358,N_8286,N_9829);
or U13359 (N_13359,N_5823,N_9301);
or U13360 (N_13360,N_9598,N_9783);
xnor U13361 (N_13361,N_9550,N_5845);
or U13362 (N_13362,N_7754,N_6328);
nor U13363 (N_13363,N_7383,N_6554);
or U13364 (N_13364,N_6559,N_9412);
or U13365 (N_13365,N_6316,N_7862);
nor U13366 (N_13366,N_7839,N_7711);
nor U13367 (N_13367,N_6198,N_9413);
or U13368 (N_13368,N_9441,N_6258);
nor U13369 (N_13369,N_6236,N_6864);
and U13370 (N_13370,N_7280,N_9026);
and U13371 (N_13371,N_6609,N_7849);
or U13372 (N_13372,N_8909,N_5911);
and U13373 (N_13373,N_5556,N_9804);
or U13374 (N_13374,N_7577,N_5357);
nand U13375 (N_13375,N_6882,N_9317);
or U13376 (N_13376,N_8258,N_7593);
and U13377 (N_13377,N_5166,N_5890);
nor U13378 (N_13378,N_6483,N_7174);
or U13379 (N_13379,N_8592,N_6198);
nand U13380 (N_13380,N_5875,N_9987);
or U13381 (N_13381,N_5147,N_5705);
or U13382 (N_13382,N_5400,N_7148);
nor U13383 (N_13383,N_6348,N_7097);
nand U13384 (N_13384,N_7364,N_5980);
xnor U13385 (N_13385,N_9003,N_7090);
and U13386 (N_13386,N_9947,N_6435);
and U13387 (N_13387,N_8938,N_9418);
or U13388 (N_13388,N_5118,N_5060);
xor U13389 (N_13389,N_9975,N_6699);
nand U13390 (N_13390,N_5353,N_8000);
and U13391 (N_13391,N_5424,N_8514);
or U13392 (N_13392,N_8744,N_9136);
nor U13393 (N_13393,N_9707,N_5251);
nor U13394 (N_13394,N_6629,N_6093);
and U13395 (N_13395,N_9316,N_6390);
nand U13396 (N_13396,N_8353,N_6899);
and U13397 (N_13397,N_7954,N_7685);
nand U13398 (N_13398,N_8792,N_8536);
and U13399 (N_13399,N_9432,N_5382);
nand U13400 (N_13400,N_5707,N_8161);
or U13401 (N_13401,N_9436,N_9294);
nand U13402 (N_13402,N_8761,N_6717);
and U13403 (N_13403,N_9895,N_9671);
nand U13404 (N_13404,N_7797,N_5183);
xnor U13405 (N_13405,N_5241,N_9386);
nand U13406 (N_13406,N_5355,N_6646);
or U13407 (N_13407,N_9320,N_9710);
and U13408 (N_13408,N_9559,N_5879);
nand U13409 (N_13409,N_8597,N_9035);
and U13410 (N_13410,N_5042,N_8239);
and U13411 (N_13411,N_8325,N_7510);
nand U13412 (N_13412,N_5764,N_6987);
nor U13413 (N_13413,N_9924,N_6871);
nor U13414 (N_13414,N_7912,N_9995);
and U13415 (N_13415,N_6267,N_7363);
nor U13416 (N_13416,N_6541,N_7199);
and U13417 (N_13417,N_9603,N_7487);
nand U13418 (N_13418,N_9690,N_6213);
and U13419 (N_13419,N_8058,N_8208);
or U13420 (N_13420,N_9461,N_5618);
and U13421 (N_13421,N_7102,N_5063);
and U13422 (N_13422,N_5778,N_6502);
nor U13423 (N_13423,N_9237,N_7010);
xnor U13424 (N_13424,N_5118,N_5810);
or U13425 (N_13425,N_6533,N_6730);
or U13426 (N_13426,N_6110,N_6496);
xor U13427 (N_13427,N_5706,N_8967);
nand U13428 (N_13428,N_9930,N_6209);
nand U13429 (N_13429,N_7274,N_9175);
nor U13430 (N_13430,N_7695,N_8811);
nor U13431 (N_13431,N_8730,N_6410);
or U13432 (N_13432,N_5685,N_5176);
and U13433 (N_13433,N_5532,N_8284);
or U13434 (N_13434,N_7367,N_7603);
and U13435 (N_13435,N_9313,N_6363);
or U13436 (N_13436,N_8799,N_9043);
and U13437 (N_13437,N_6749,N_5786);
nand U13438 (N_13438,N_5023,N_9194);
nor U13439 (N_13439,N_6087,N_7909);
nor U13440 (N_13440,N_8797,N_8717);
and U13441 (N_13441,N_5106,N_6806);
and U13442 (N_13442,N_7034,N_9180);
nand U13443 (N_13443,N_7661,N_7415);
nor U13444 (N_13444,N_6567,N_5246);
or U13445 (N_13445,N_9826,N_7798);
or U13446 (N_13446,N_6968,N_8614);
or U13447 (N_13447,N_8152,N_7564);
nor U13448 (N_13448,N_8481,N_8524);
or U13449 (N_13449,N_9528,N_9622);
and U13450 (N_13450,N_7445,N_5190);
nor U13451 (N_13451,N_6810,N_7682);
and U13452 (N_13452,N_5027,N_8378);
and U13453 (N_13453,N_7859,N_5991);
nand U13454 (N_13454,N_9212,N_7750);
and U13455 (N_13455,N_6265,N_5871);
and U13456 (N_13456,N_8151,N_5296);
or U13457 (N_13457,N_5448,N_9611);
or U13458 (N_13458,N_7841,N_6581);
or U13459 (N_13459,N_5788,N_5545);
xnor U13460 (N_13460,N_9047,N_8027);
and U13461 (N_13461,N_9326,N_5973);
or U13462 (N_13462,N_5486,N_8177);
nand U13463 (N_13463,N_6666,N_6109);
or U13464 (N_13464,N_8915,N_5947);
xor U13465 (N_13465,N_8585,N_5410);
and U13466 (N_13466,N_8052,N_7995);
nand U13467 (N_13467,N_8423,N_8139);
nor U13468 (N_13468,N_9859,N_5703);
or U13469 (N_13469,N_8024,N_5831);
nand U13470 (N_13470,N_7243,N_7640);
nor U13471 (N_13471,N_7970,N_7269);
nor U13472 (N_13472,N_9139,N_8508);
nor U13473 (N_13473,N_9253,N_8134);
and U13474 (N_13474,N_5163,N_6877);
xnor U13475 (N_13475,N_7449,N_8228);
nor U13476 (N_13476,N_8492,N_7317);
nor U13477 (N_13477,N_7829,N_6924);
xor U13478 (N_13478,N_7906,N_9351);
or U13479 (N_13479,N_6456,N_5437);
nor U13480 (N_13480,N_7450,N_6955);
nor U13481 (N_13481,N_9485,N_7020);
and U13482 (N_13482,N_7880,N_9966);
xnor U13483 (N_13483,N_5047,N_7221);
nand U13484 (N_13484,N_5550,N_5213);
and U13485 (N_13485,N_5316,N_8317);
and U13486 (N_13486,N_7741,N_6418);
nor U13487 (N_13487,N_9867,N_8104);
xnor U13488 (N_13488,N_8018,N_8466);
xor U13489 (N_13489,N_8953,N_6015);
and U13490 (N_13490,N_6911,N_8037);
nand U13491 (N_13491,N_6919,N_8625);
or U13492 (N_13492,N_7605,N_9013);
xor U13493 (N_13493,N_8943,N_8900);
and U13494 (N_13494,N_6695,N_8473);
and U13495 (N_13495,N_5139,N_5006);
or U13496 (N_13496,N_7337,N_7004);
nor U13497 (N_13497,N_8809,N_8887);
or U13498 (N_13498,N_8689,N_8722);
nand U13499 (N_13499,N_6120,N_8138);
nor U13500 (N_13500,N_6543,N_5331);
nor U13501 (N_13501,N_8407,N_9681);
nor U13502 (N_13502,N_7297,N_7130);
or U13503 (N_13503,N_5676,N_5140);
xor U13504 (N_13504,N_8972,N_6949);
nand U13505 (N_13505,N_8622,N_6513);
xor U13506 (N_13506,N_6442,N_8858);
or U13507 (N_13507,N_8269,N_6182);
nor U13508 (N_13508,N_7518,N_8673);
nand U13509 (N_13509,N_9293,N_7179);
nand U13510 (N_13510,N_9532,N_8989);
and U13511 (N_13511,N_8791,N_8052);
or U13512 (N_13512,N_8737,N_6372);
xnor U13513 (N_13513,N_9396,N_6230);
nor U13514 (N_13514,N_8985,N_5122);
nor U13515 (N_13515,N_6781,N_9716);
nor U13516 (N_13516,N_7848,N_8689);
or U13517 (N_13517,N_5919,N_5181);
nor U13518 (N_13518,N_5844,N_5888);
or U13519 (N_13519,N_7834,N_6398);
xnor U13520 (N_13520,N_6977,N_6371);
and U13521 (N_13521,N_8292,N_6058);
or U13522 (N_13522,N_6698,N_8033);
nor U13523 (N_13523,N_5417,N_9524);
nor U13524 (N_13524,N_9630,N_9113);
or U13525 (N_13525,N_5387,N_6421);
nor U13526 (N_13526,N_5063,N_6511);
xnor U13527 (N_13527,N_8693,N_8654);
or U13528 (N_13528,N_9075,N_7586);
xnor U13529 (N_13529,N_8334,N_9350);
nor U13530 (N_13530,N_9809,N_5553);
nor U13531 (N_13531,N_7557,N_9468);
xor U13532 (N_13532,N_7113,N_7994);
and U13533 (N_13533,N_5870,N_5812);
and U13534 (N_13534,N_8943,N_8786);
nand U13535 (N_13535,N_6663,N_9108);
and U13536 (N_13536,N_5218,N_8734);
or U13537 (N_13537,N_7494,N_5083);
and U13538 (N_13538,N_7644,N_5055);
nor U13539 (N_13539,N_8014,N_6526);
nand U13540 (N_13540,N_7069,N_9079);
xnor U13541 (N_13541,N_7395,N_9406);
nand U13542 (N_13542,N_5495,N_8526);
nand U13543 (N_13543,N_5897,N_8839);
xnor U13544 (N_13544,N_6248,N_7717);
nor U13545 (N_13545,N_5661,N_5867);
or U13546 (N_13546,N_6162,N_8944);
nor U13547 (N_13547,N_9393,N_8324);
and U13548 (N_13548,N_9219,N_7001);
and U13549 (N_13549,N_5652,N_5048);
nand U13550 (N_13550,N_6534,N_7044);
nand U13551 (N_13551,N_5889,N_8155);
nor U13552 (N_13552,N_8973,N_8846);
nor U13553 (N_13553,N_5110,N_5745);
nand U13554 (N_13554,N_8461,N_6472);
and U13555 (N_13555,N_7250,N_7076);
nand U13556 (N_13556,N_8367,N_6806);
nand U13557 (N_13557,N_8899,N_9917);
or U13558 (N_13558,N_5480,N_7474);
nor U13559 (N_13559,N_6522,N_5915);
or U13560 (N_13560,N_6443,N_7738);
or U13561 (N_13561,N_7614,N_6840);
and U13562 (N_13562,N_7144,N_6299);
and U13563 (N_13563,N_5227,N_6644);
or U13564 (N_13564,N_7508,N_9917);
or U13565 (N_13565,N_6980,N_9853);
nor U13566 (N_13566,N_8391,N_9872);
or U13567 (N_13567,N_8031,N_7912);
or U13568 (N_13568,N_5985,N_5126);
or U13569 (N_13569,N_6280,N_7927);
and U13570 (N_13570,N_9733,N_7675);
nor U13571 (N_13571,N_6725,N_8516);
and U13572 (N_13572,N_8249,N_5376);
nor U13573 (N_13573,N_6180,N_9023);
or U13574 (N_13574,N_6908,N_7207);
or U13575 (N_13575,N_7979,N_8752);
nor U13576 (N_13576,N_7901,N_6670);
or U13577 (N_13577,N_6811,N_5234);
nor U13578 (N_13578,N_6547,N_9855);
and U13579 (N_13579,N_5239,N_7934);
nand U13580 (N_13580,N_5076,N_7049);
xor U13581 (N_13581,N_5743,N_9451);
xor U13582 (N_13582,N_7187,N_9313);
or U13583 (N_13583,N_7874,N_6612);
and U13584 (N_13584,N_6256,N_6936);
nand U13585 (N_13585,N_6540,N_8906);
and U13586 (N_13586,N_5911,N_8595);
or U13587 (N_13587,N_7582,N_5346);
and U13588 (N_13588,N_8411,N_9331);
nor U13589 (N_13589,N_5375,N_8014);
and U13590 (N_13590,N_8662,N_8745);
xor U13591 (N_13591,N_8313,N_8674);
nor U13592 (N_13592,N_9852,N_7896);
or U13593 (N_13593,N_7329,N_6002);
or U13594 (N_13594,N_8941,N_8763);
or U13595 (N_13595,N_8150,N_6536);
nor U13596 (N_13596,N_5346,N_6713);
and U13597 (N_13597,N_5513,N_5429);
nor U13598 (N_13598,N_5700,N_5814);
nor U13599 (N_13599,N_5370,N_7994);
nand U13600 (N_13600,N_7994,N_6020);
nor U13601 (N_13601,N_8284,N_6730);
nor U13602 (N_13602,N_6936,N_9734);
or U13603 (N_13603,N_9656,N_9537);
or U13604 (N_13604,N_7862,N_9072);
or U13605 (N_13605,N_5808,N_5665);
or U13606 (N_13606,N_8459,N_9537);
nor U13607 (N_13607,N_8040,N_6163);
xor U13608 (N_13608,N_7732,N_7824);
nor U13609 (N_13609,N_6222,N_8719);
nor U13610 (N_13610,N_9184,N_5230);
nand U13611 (N_13611,N_5307,N_6692);
nand U13612 (N_13612,N_8383,N_8008);
nor U13613 (N_13613,N_6165,N_7780);
nor U13614 (N_13614,N_6284,N_7054);
or U13615 (N_13615,N_9480,N_8160);
nor U13616 (N_13616,N_7683,N_5915);
nor U13617 (N_13617,N_9536,N_6976);
nor U13618 (N_13618,N_8817,N_8756);
and U13619 (N_13619,N_9484,N_9834);
and U13620 (N_13620,N_6258,N_7970);
and U13621 (N_13621,N_6346,N_6416);
nor U13622 (N_13622,N_6369,N_6311);
and U13623 (N_13623,N_8687,N_8356);
or U13624 (N_13624,N_7674,N_8361);
and U13625 (N_13625,N_6111,N_6639);
and U13626 (N_13626,N_8723,N_5713);
or U13627 (N_13627,N_8708,N_6717);
or U13628 (N_13628,N_9252,N_5063);
nor U13629 (N_13629,N_6662,N_6483);
or U13630 (N_13630,N_9584,N_6889);
and U13631 (N_13631,N_9523,N_8465);
nand U13632 (N_13632,N_7361,N_8773);
and U13633 (N_13633,N_5992,N_5087);
and U13634 (N_13634,N_8859,N_7428);
nand U13635 (N_13635,N_9014,N_9723);
nand U13636 (N_13636,N_9016,N_7215);
or U13637 (N_13637,N_5059,N_9986);
nor U13638 (N_13638,N_7920,N_9916);
nor U13639 (N_13639,N_5004,N_9524);
and U13640 (N_13640,N_9555,N_6883);
nand U13641 (N_13641,N_9972,N_6707);
nor U13642 (N_13642,N_8777,N_6563);
and U13643 (N_13643,N_5534,N_8538);
or U13644 (N_13644,N_7018,N_8924);
and U13645 (N_13645,N_6507,N_6418);
and U13646 (N_13646,N_8625,N_7186);
xnor U13647 (N_13647,N_7403,N_5144);
and U13648 (N_13648,N_5661,N_6061);
xnor U13649 (N_13649,N_7621,N_8735);
xor U13650 (N_13650,N_6308,N_5380);
nor U13651 (N_13651,N_5190,N_7506);
nand U13652 (N_13652,N_7805,N_6564);
nor U13653 (N_13653,N_6915,N_9984);
nor U13654 (N_13654,N_8901,N_6602);
xnor U13655 (N_13655,N_9403,N_8994);
nor U13656 (N_13656,N_5009,N_7633);
or U13657 (N_13657,N_5345,N_9869);
or U13658 (N_13658,N_7481,N_9793);
nor U13659 (N_13659,N_6488,N_5063);
or U13660 (N_13660,N_5955,N_6143);
nor U13661 (N_13661,N_6839,N_6051);
or U13662 (N_13662,N_8052,N_7699);
nand U13663 (N_13663,N_7312,N_8396);
and U13664 (N_13664,N_5035,N_5261);
nand U13665 (N_13665,N_6775,N_7266);
nand U13666 (N_13666,N_7866,N_7888);
and U13667 (N_13667,N_5152,N_6076);
xnor U13668 (N_13668,N_8615,N_7130);
or U13669 (N_13669,N_7758,N_5013);
nand U13670 (N_13670,N_8310,N_9198);
or U13671 (N_13671,N_7916,N_5607);
and U13672 (N_13672,N_9756,N_9646);
xor U13673 (N_13673,N_8273,N_9979);
nor U13674 (N_13674,N_7322,N_6309);
nand U13675 (N_13675,N_9596,N_8861);
and U13676 (N_13676,N_7998,N_7993);
nand U13677 (N_13677,N_7513,N_7627);
and U13678 (N_13678,N_8773,N_7368);
or U13679 (N_13679,N_8503,N_9441);
nand U13680 (N_13680,N_9296,N_6017);
nand U13681 (N_13681,N_7626,N_8272);
and U13682 (N_13682,N_6351,N_8464);
or U13683 (N_13683,N_9829,N_9110);
xnor U13684 (N_13684,N_6716,N_7285);
xor U13685 (N_13685,N_7247,N_8528);
or U13686 (N_13686,N_8678,N_5756);
and U13687 (N_13687,N_7881,N_8205);
nor U13688 (N_13688,N_8053,N_9948);
or U13689 (N_13689,N_6606,N_6078);
xnor U13690 (N_13690,N_9176,N_9386);
nand U13691 (N_13691,N_8260,N_7031);
and U13692 (N_13692,N_9476,N_8733);
or U13693 (N_13693,N_5708,N_7852);
and U13694 (N_13694,N_8502,N_5398);
nor U13695 (N_13695,N_9885,N_9780);
nor U13696 (N_13696,N_5169,N_5792);
nor U13697 (N_13697,N_5654,N_5224);
or U13698 (N_13698,N_9495,N_5030);
or U13699 (N_13699,N_8084,N_5826);
nor U13700 (N_13700,N_8795,N_7689);
nor U13701 (N_13701,N_6741,N_6951);
nor U13702 (N_13702,N_5239,N_7265);
and U13703 (N_13703,N_5082,N_6888);
nand U13704 (N_13704,N_7146,N_6648);
nor U13705 (N_13705,N_9239,N_9106);
nor U13706 (N_13706,N_7777,N_5809);
nand U13707 (N_13707,N_8929,N_7817);
xor U13708 (N_13708,N_8156,N_5244);
nand U13709 (N_13709,N_6557,N_8841);
or U13710 (N_13710,N_9692,N_5211);
or U13711 (N_13711,N_8534,N_5043);
nand U13712 (N_13712,N_5158,N_9444);
or U13713 (N_13713,N_8010,N_6604);
nand U13714 (N_13714,N_8292,N_7155);
nand U13715 (N_13715,N_5460,N_8983);
or U13716 (N_13716,N_9947,N_9811);
nor U13717 (N_13717,N_8924,N_6402);
xnor U13718 (N_13718,N_9714,N_8416);
nor U13719 (N_13719,N_5796,N_8991);
nand U13720 (N_13720,N_8426,N_6282);
nand U13721 (N_13721,N_7598,N_7987);
xor U13722 (N_13722,N_5202,N_5746);
nor U13723 (N_13723,N_6367,N_6804);
nand U13724 (N_13724,N_8282,N_6848);
xnor U13725 (N_13725,N_6318,N_8949);
and U13726 (N_13726,N_9381,N_9324);
nor U13727 (N_13727,N_9347,N_7699);
nand U13728 (N_13728,N_8492,N_7003);
nand U13729 (N_13729,N_5163,N_8255);
or U13730 (N_13730,N_8566,N_9910);
or U13731 (N_13731,N_8967,N_6567);
and U13732 (N_13732,N_6225,N_8436);
nand U13733 (N_13733,N_9369,N_5705);
nand U13734 (N_13734,N_5354,N_6006);
and U13735 (N_13735,N_5514,N_8350);
xor U13736 (N_13736,N_8519,N_5308);
nand U13737 (N_13737,N_5487,N_8896);
nand U13738 (N_13738,N_5098,N_6442);
nor U13739 (N_13739,N_6555,N_8132);
nand U13740 (N_13740,N_9011,N_6413);
and U13741 (N_13741,N_8977,N_5347);
nand U13742 (N_13742,N_7849,N_7005);
nand U13743 (N_13743,N_6087,N_9071);
and U13744 (N_13744,N_9532,N_6928);
nor U13745 (N_13745,N_8484,N_6555);
nand U13746 (N_13746,N_9183,N_7340);
nand U13747 (N_13747,N_9803,N_9031);
nand U13748 (N_13748,N_8857,N_8433);
and U13749 (N_13749,N_6941,N_7880);
and U13750 (N_13750,N_8224,N_7621);
nor U13751 (N_13751,N_6817,N_8569);
or U13752 (N_13752,N_9469,N_7719);
nor U13753 (N_13753,N_7484,N_8151);
nand U13754 (N_13754,N_6830,N_9813);
nor U13755 (N_13755,N_9090,N_8582);
and U13756 (N_13756,N_8646,N_8864);
or U13757 (N_13757,N_9572,N_9419);
or U13758 (N_13758,N_6525,N_5854);
or U13759 (N_13759,N_8820,N_6500);
nand U13760 (N_13760,N_6772,N_9591);
nor U13761 (N_13761,N_5126,N_9345);
xor U13762 (N_13762,N_5559,N_7971);
and U13763 (N_13763,N_6375,N_9994);
and U13764 (N_13764,N_7587,N_9121);
nand U13765 (N_13765,N_5290,N_5168);
or U13766 (N_13766,N_6965,N_9803);
nor U13767 (N_13767,N_8425,N_9575);
nand U13768 (N_13768,N_6065,N_5079);
xnor U13769 (N_13769,N_6190,N_9672);
nor U13770 (N_13770,N_8321,N_5886);
or U13771 (N_13771,N_8353,N_6469);
xnor U13772 (N_13772,N_6508,N_8107);
or U13773 (N_13773,N_8400,N_8175);
nand U13774 (N_13774,N_6636,N_6818);
and U13775 (N_13775,N_9488,N_9181);
nor U13776 (N_13776,N_9142,N_7209);
and U13777 (N_13777,N_5908,N_5569);
nor U13778 (N_13778,N_8233,N_9710);
nand U13779 (N_13779,N_6514,N_9330);
nor U13780 (N_13780,N_7054,N_8777);
xor U13781 (N_13781,N_9104,N_6541);
or U13782 (N_13782,N_5716,N_9170);
or U13783 (N_13783,N_6175,N_7034);
nand U13784 (N_13784,N_6704,N_5896);
xor U13785 (N_13785,N_8612,N_9799);
nand U13786 (N_13786,N_5614,N_7747);
xor U13787 (N_13787,N_5515,N_7928);
nand U13788 (N_13788,N_7722,N_5774);
or U13789 (N_13789,N_9603,N_5518);
nor U13790 (N_13790,N_9659,N_9035);
and U13791 (N_13791,N_6178,N_6722);
or U13792 (N_13792,N_7440,N_7725);
nor U13793 (N_13793,N_7778,N_5118);
nor U13794 (N_13794,N_5839,N_7422);
or U13795 (N_13795,N_6526,N_7562);
nand U13796 (N_13796,N_7502,N_6333);
nand U13797 (N_13797,N_9371,N_7206);
nand U13798 (N_13798,N_8402,N_8436);
nor U13799 (N_13799,N_9790,N_7699);
or U13800 (N_13800,N_7012,N_9199);
nor U13801 (N_13801,N_7818,N_5554);
or U13802 (N_13802,N_9285,N_7475);
nor U13803 (N_13803,N_5511,N_8003);
or U13804 (N_13804,N_8461,N_7497);
or U13805 (N_13805,N_5927,N_8936);
or U13806 (N_13806,N_9704,N_8693);
xor U13807 (N_13807,N_7888,N_5139);
and U13808 (N_13808,N_7883,N_9861);
and U13809 (N_13809,N_6226,N_7920);
and U13810 (N_13810,N_5111,N_7948);
nand U13811 (N_13811,N_5581,N_5337);
and U13812 (N_13812,N_5519,N_8032);
nand U13813 (N_13813,N_8872,N_7993);
nand U13814 (N_13814,N_7021,N_8397);
xor U13815 (N_13815,N_8823,N_8662);
and U13816 (N_13816,N_7336,N_5192);
and U13817 (N_13817,N_8265,N_6078);
nand U13818 (N_13818,N_6912,N_7853);
nand U13819 (N_13819,N_8589,N_7690);
nor U13820 (N_13820,N_6684,N_6822);
xor U13821 (N_13821,N_7158,N_8777);
or U13822 (N_13822,N_8795,N_9531);
and U13823 (N_13823,N_9677,N_5113);
nor U13824 (N_13824,N_6921,N_7982);
nor U13825 (N_13825,N_7763,N_7362);
nor U13826 (N_13826,N_6529,N_7824);
and U13827 (N_13827,N_8465,N_5705);
and U13828 (N_13828,N_8665,N_9037);
and U13829 (N_13829,N_8707,N_7498);
nor U13830 (N_13830,N_5627,N_8043);
xnor U13831 (N_13831,N_8167,N_7840);
nor U13832 (N_13832,N_5648,N_9919);
nand U13833 (N_13833,N_6083,N_9842);
nand U13834 (N_13834,N_5134,N_8038);
nor U13835 (N_13835,N_5560,N_7740);
or U13836 (N_13836,N_6853,N_9539);
nand U13837 (N_13837,N_8879,N_7617);
xor U13838 (N_13838,N_5082,N_9828);
nand U13839 (N_13839,N_9193,N_6616);
or U13840 (N_13840,N_7088,N_7063);
or U13841 (N_13841,N_7828,N_9964);
or U13842 (N_13842,N_6467,N_7210);
nor U13843 (N_13843,N_5471,N_6573);
xnor U13844 (N_13844,N_7053,N_6055);
or U13845 (N_13845,N_5176,N_9735);
and U13846 (N_13846,N_6407,N_7603);
or U13847 (N_13847,N_7055,N_7458);
nor U13848 (N_13848,N_5710,N_7405);
and U13849 (N_13849,N_7936,N_5070);
nand U13850 (N_13850,N_9910,N_6176);
nor U13851 (N_13851,N_5534,N_9865);
nand U13852 (N_13852,N_8366,N_9276);
and U13853 (N_13853,N_5011,N_6524);
or U13854 (N_13854,N_7852,N_5107);
and U13855 (N_13855,N_9565,N_9910);
nor U13856 (N_13856,N_7616,N_8184);
nand U13857 (N_13857,N_8358,N_5015);
nand U13858 (N_13858,N_8962,N_8813);
nor U13859 (N_13859,N_9421,N_7924);
and U13860 (N_13860,N_5790,N_5691);
or U13861 (N_13861,N_8724,N_5885);
nand U13862 (N_13862,N_8100,N_8158);
or U13863 (N_13863,N_6892,N_9256);
or U13864 (N_13864,N_9878,N_8047);
nand U13865 (N_13865,N_7853,N_9349);
nand U13866 (N_13866,N_9870,N_6659);
or U13867 (N_13867,N_9980,N_8490);
nor U13868 (N_13868,N_5699,N_9733);
nor U13869 (N_13869,N_5356,N_9257);
nand U13870 (N_13870,N_9176,N_8269);
or U13871 (N_13871,N_5678,N_8588);
nand U13872 (N_13872,N_9327,N_5556);
nand U13873 (N_13873,N_6503,N_6762);
and U13874 (N_13874,N_8693,N_5476);
nand U13875 (N_13875,N_7519,N_6970);
nor U13876 (N_13876,N_5460,N_9947);
or U13877 (N_13877,N_9886,N_6344);
or U13878 (N_13878,N_5628,N_7116);
nor U13879 (N_13879,N_5565,N_9435);
and U13880 (N_13880,N_5698,N_8418);
or U13881 (N_13881,N_8428,N_8574);
nor U13882 (N_13882,N_6462,N_9805);
nand U13883 (N_13883,N_6186,N_7898);
or U13884 (N_13884,N_6713,N_7197);
or U13885 (N_13885,N_6835,N_8288);
and U13886 (N_13886,N_9653,N_6193);
nor U13887 (N_13887,N_5453,N_8395);
and U13888 (N_13888,N_9800,N_7159);
and U13889 (N_13889,N_7218,N_6753);
nor U13890 (N_13890,N_5765,N_5970);
nand U13891 (N_13891,N_8649,N_6758);
and U13892 (N_13892,N_5195,N_8545);
nand U13893 (N_13893,N_8168,N_9409);
nand U13894 (N_13894,N_7954,N_8285);
or U13895 (N_13895,N_7488,N_9288);
xor U13896 (N_13896,N_7638,N_5588);
or U13897 (N_13897,N_5074,N_7587);
and U13898 (N_13898,N_6237,N_6161);
nand U13899 (N_13899,N_7923,N_9604);
xnor U13900 (N_13900,N_9446,N_7811);
or U13901 (N_13901,N_9182,N_7849);
or U13902 (N_13902,N_5121,N_5753);
or U13903 (N_13903,N_8436,N_8951);
or U13904 (N_13904,N_7949,N_8223);
nand U13905 (N_13905,N_6113,N_7920);
or U13906 (N_13906,N_8105,N_7713);
xor U13907 (N_13907,N_6021,N_6087);
nand U13908 (N_13908,N_6269,N_6085);
nor U13909 (N_13909,N_8409,N_6409);
or U13910 (N_13910,N_6271,N_6284);
and U13911 (N_13911,N_9740,N_8324);
and U13912 (N_13912,N_6802,N_5089);
and U13913 (N_13913,N_8046,N_5510);
nor U13914 (N_13914,N_6164,N_9904);
or U13915 (N_13915,N_8631,N_8510);
nor U13916 (N_13916,N_6546,N_8862);
nor U13917 (N_13917,N_7186,N_6070);
or U13918 (N_13918,N_9162,N_6676);
nor U13919 (N_13919,N_9357,N_6507);
or U13920 (N_13920,N_9734,N_8256);
or U13921 (N_13921,N_7308,N_7567);
nor U13922 (N_13922,N_5680,N_5993);
or U13923 (N_13923,N_8179,N_9178);
nand U13924 (N_13924,N_7272,N_9197);
and U13925 (N_13925,N_6871,N_6671);
or U13926 (N_13926,N_6367,N_8202);
or U13927 (N_13927,N_9000,N_5999);
and U13928 (N_13928,N_5533,N_6361);
nand U13929 (N_13929,N_9899,N_9091);
and U13930 (N_13930,N_9279,N_6753);
nor U13931 (N_13931,N_7924,N_5211);
nand U13932 (N_13932,N_8168,N_8640);
nand U13933 (N_13933,N_8373,N_9882);
nand U13934 (N_13934,N_9606,N_6193);
and U13935 (N_13935,N_5261,N_7066);
nand U13936 (N_13936,N_7944,N_8100);
nor U13937 (N_13937,N_6876,N_6860);
nor U13938 (N_13938,N_7205,N_6516);
nor U13939 (N_13939,N_7685,N_8985);
nor U13940 (N_13940,N_7831,N_7363);
nand U13941 (N_13941,N_5850,N_6139);
and U13942 (N_13942,N_7960,N_9442);
or U13943 (N_13943,N_6020,N_5131);
xor U13944 (N_13944,N_9480,N_6108);
nor U13945 (N_13945,N_6595,N_6206);
and U13946 (N_13946,N_8212,N_5520);
and U13947 (N_13947,N_7305,N_8408);
nand U13948 (N_13948,N_8184,N_9635);
nand U13949 (N_13949,N_8984,N_5930);
nand U13950 (N_13950,N_7461,N_9521);
and U13951 (N_13951,N_6305,N_9977);
nor U13952 (N_13952,N_6198,N_6341);
and U13953 (N_13953,N_9626,N_7391);
or U13954 (N_13954,N_8227,N_6011);
or U13955 (N_13955,N_8916,N_7546);
and U13956 (N_13956,N_9259,N_7409);
nand U13957 (N_13957,N_5069,N_9916);
nand U13958 (N_13958,N_6662,N_9065);
or U13959 (N_13959,N_6710,N_7405);
nor U13960 (N_13960,N_8096,N_8011);
or U13961 (N_13961,N_6303,N_8935);
or U13962 (N_13962,N_6332,N_5968);
and U13963 (N_13963,N_8268,N_7960);
and U13964 (N_13964,N_6752,N_5104);
and U13965 (N_13965,N_6766,N_6287);
or U13966 (N_13966,N_8245,N_9768);
and U13967 (N_13967,N_5542,N_5002);
or U13968 (N_13968,N_9540,N_9599);
or U13969 (N_13969,N_7227,N_5120);
nand U13970 (N_13970,N_6589,N_5272);
nand U13971 (N_13971,N_6961,N_5258);
nand U13972 (N_13972,N_6941,N_5668);
or U13973 (N_13973,N_7312,N_5309);
or U13974 (N_13974,N_5320,N_9982);
or U13975 (N_13975,N_6801,N_9141);
or U13976 (N_13976,N_6635,N_9879);
and U13977 (N_13977,N_6742,N_6356);
or U13978 (N_13978,N_6339,N_6366);
nor U13979 (N_13979,N_5857,N_8057);
nand U13980 (N_13980,N_6735,N_9987);
or U13981 (N_13981,N_5021,N_6189);
nand U13982 (N_13982,N_8089,N_8507);
or U13983 (N_13983,N_7062,N_7736);
nand U13984 (N_13984,N_5641,N_9596);
nand U13985 (N_13985,N_6567,N_7400);
and U13986 (N_13986,N_7918,N_6451);
and U13987 (N_13987,N_6924,N_5958);
nand U13988 (N_13988,N_7727,N_6205);
or U13989 (N_13989,N_7956,N_7635);
nand U13990 (N_13990,N_7997,N_9640);
nor U13991 (N_13991,N_7197,N_5370);
and U13992 (N_13992,N_5522,N_7284);
nand U13993 (N_13993,N_6544,N_6370);
or U13994 (N_13994,N_6822,N_5888);
nor U13995 (N_13995,N_5946,N_5598);
or U13996 (N_13996,N_8248,N_6249);
or U13997 (N_13997,N_9455,N_6641);
nand U13998 (N_13998,N_7628,N_8863);
nand U13999 (N_13999,N_5960,N_5491);
nor U14000 (N_14000,N_6693,N_6940);
or U14001 (N_14001,N_6528,N_7970);
or U14002 (N_14002,N_9953,N_6202);
nand U14003 (N_14003,N_6705,N_7220);
nor U14004 (N_14004,N_7246,N_8713);
xnor U14005 (N_14005,N_5387,N_5184);
xnor U14006 (N_14006,N_8912,N_8044);
or U14007 (N_14007,N_7700,N_9017);
xor U14008 (N_14008,N_6656,N_7101);
or U14009 (N_14009,N_7002,N_9645);
nor U14010 (N_14010,N_5589,N_6716);
nor U14011 (N_14011,N_6399,N_5672);
or U14012 (N_14012,N_9170,N_6427);
or U14013 (N_14013,N_6823,N_6178);
nor U14014 (N_14014,N_9173,N_8565);
nor U14015 (N_14015,N_5031,N_5223);
nor U14016 (N_14016,N_9069,N_5750);
and U14017 (N_14017,N_6938,N_8011);
nand U14018 (N_14018,N_5042,N_8078);
and U14019 (N_14019,N_5080,N_6415);
nand U14020 (N_14020,N_6019,N_9320);
xnor U14021 (N_14021,N_6215,N_9465);
nor U14022 (N_14022,N_5365,N_5560);
or U14023 (N_14023,N_9911,N_9595);
nand U14024 (N_14024,N_5355,N_5202);
and U14025 (N_14025,N_6885,N_9832);
nor U14026 (N_14026,N_8841,N_8390);
xnor U14027 (N_14027,N_5368,N_5334);
or U14028 (N_14028,N_6298,N_8610);
and U14029 (N_14029,N_8352,N_5632);
or U14030 (N_14030,N_8395,N_9103);
nor U14031 (N_14031,N_7961,N_7534);
or U14032 (N_14032,N_5055,N_8388);
and U14033 (N_14033,N_8833,N_7256);
nand U14034 (N_14034,N_9446,N_8754);
xor U14035 (N_14035,N_7718,N_7404);
or U14036 (N_14036,N_5358,N_9134);
nand U14037 (N_14037,N_5369,N_7000);
nor U14038 (N_14038,N_6387,N_7689);
nand U14039 (N_14039,N_5849,N_7703);
and U14040 (N_14040,N_9552,N_6641);
and U14041 (N_14041,N_8164,N_6733);
xor U14042 (N_14042,N_5865,N_7576);
nand U14043 (N_14043,N_7246,N_9701);
or U14044 (N_14044,N_5577,N_6668);
nand U14045 (N_14045,N_6797,N_5753);
or U14046 (N_14046,N_7986,N_7682);
nand U14047 (N_14047,N_8702,N_9990);
xor U14048 (N_14048,N_6854,N_9273);
or U14049 (N_14049,N_8116,N_9975);
nand U14050 (N_14050,N_8462,N_9742);
or U14051 (N_14051,N_6869,N_9370);
or U14052 (N_14052,N_7713,N_5292);
or U14053 (N_14053,N_6392,N_8667);
nor U14054 (N_14054,N_9872,N_7997);
or U14055 (N_14055,N_9429,N_8285);
nor U14056 (N_14056,N_5546,N_8669);
nand U14057 (N_14057,N_6758,N_7462);
and U14058 (N_14058,N_5718,N_6213);
nor U14059 (N_14059,N_6617,N_7528);
or U14060 (N_14060,N_8809,N_6888);
nand U14061 (N_14061,N_9301,N_8288);
nand U14062 (N_14062,N_8833,N_5872);
xnor U14063 (N_14063,N_7862,N_8944);
nor U14064 (N_14064,N_8683,N_7135);
xnor U14065 (N_14065,N_5993,N_6348);
and U14066 (N_14066,N_7397,N_5731);
xnor U14067 (N_14067,N_6764,N_9770);
nand U14068 (N_14068,N_5558,N_7979);
or U14069 (N_14069,N_7098,N_9294);
xor U14070 (N_14070,N_6786,N_7580);
or U14071 (N_14071,N_7426,N_7417);
nor U14072 (N_14072,N_5629,N_6538);
nor U14073 (N_14073,N_7891,N_5576);
nor U14074 (N_14074,N_6959,N_9654);
nand U14075 (N_14075,N_9027,N_8992);
and U14076 (N_14076,N_8892,N_7346);
nor U14077 (N_14077,N_8372,N_9794);
nor U14078 (N_14078,N_6033,N_8219);
and U14079 (N_14079,N_6436,N_6908);
or U14080 (N_14080,N_6417,N_8690);
or U14081 (N_14081,N_7370,N_9080);
or U14082 (N_14082,N_7776,N_8350);
and U14083 (N_14083,N_8007,N_5377);
and U14084 (N_14084,N_7285,N_9452);
and U14085 (N_14085,N_8896,N_9512);
nand U14086 (N_14086,N_6221,N_9295);
nand U14087 (N_14087,N_8750,N_8749);
or U14088 (N_14088,N_7415,N_8714);
nor U14089 (N_14089,N_7896,N_9620);
nor U14090 (N_14090,N_5864,N_8596);
xor U14091 (N_14091,N_8890,N_6530);
or U14092 (N_14092,N_6541,N_7783);
and U14093 (N_14093,N_8847,N_7213);
nor U14094 (N_14094,N_5837,N_8147);
nor U14095 (N_14095,N_8036,N_6603);
or U14096 (N_14096,N_8830,N_5717);
nand U14097 (N_14097,N_8958,N_9831);
nor U14098 (N_14098,N_8427,N_5726);
or U14099 (N_14099,N_5207,N_9169);
xor U14100 (N_14100,N_7453,N_6296);
nor U14101 (N_14101,N_8465,N_9500);
nor U14102 (N_14102,N_8562,N_8142);
nor U14103 (N_14103,N_9252,N_6863);
nand U14104 (N_14104,N_7505,N_7455);
or U14105 (N_14105,N_5695,N_7357);
nor U14106 (N_14106,N_8634,N_9207);
or U14107 (N_14107,N_8739,N_9626);
nand U14108 (N_14108,N_5297,N_8458);
or U14109 (N_14109,N_5661,N_7250);
nand U14110 (N_14110,N_9728,N_7062);
or U14111 (N_14111,N_6374,N_7947);
or U14112 (N_14112,N_9141,N_6494);
or U14113 (N_14113,N_8733,N_6888);
and U14114 (N_14114,N_9281,N_9206);
nor U14115 (N_14115,N_7632,N_7217);
xnor U14116 (N_14116,N_6405,N_5707);
and U14117 (N_14117,N_5993,N_8032);
or U14118 (N_14118,N_5409,N_7213);
nand U14119 (N_14119,N_5604,N_5550);
and U14120 (N_14120,N_5653,N_5679);
or U14121 (N_14121,N_9571,N_8067);
nand U14122 (N_14122,N_5253,N_5718);
or U14123 (N_14123,N_5206,N_7253);
nor U14124 (N_14124,N_9578,N_8514);
or U14125 (N_14125,N_9958,N_8441);
or U14126 (N_14126,N_6824,N_7472);
and U14127 (N_14127,N_8906,N_8516);
nor U14128 (N_14128,N_5348,N_7734);
nor U14129 (N_14129,N_5533,N_5782);
nand U14130 (N_14130,N_7244,N_6504);
and U14131 (N_14131,N_6036,N_8725);
and U14132 (N_14132,N_9036,N_5786);
nor U14133 (N_14133,N_6328,N_7755);
nor U14134 (N_14134,N_5784,N_9784);
nand U14135 (N_14135,N_7967,N_9589);
nand U14136 (N_14136,N_5480,N_8777);
nor U14137 (N_14137,N_7302,N_8608);
or U14138 (N_14138,N_8791,N_8364);
nor U14139 (N_14139,N_9499,N_9003);
or U14140 (N_14140,N_7964,N_5403);
nand U14141 (N_14141,N_8759,N_8089);
nor U14142 (N_14142,N_5944,N_9089);
or U14143 (N_14143,N_8951,N_9428);
or U14144 (N_14144,N_5229,N_7841);
or U14145 (N_14145,N_9307,N_5009);
nor U14146 (N_14146,N_7074,N_8984);
nand U14147 (N_14147,N_9688,N_6882);
or U14148 (N_14148,N_8087,N_6576);
or U14149 (N_14149,N_6587,N_9215);
nor U14150 (N_14150,N_9598,N_7430);
nand U14151 (N_14151,N_7613,N_5195);
nand U14152 (N_14152,N_6221,N_5165);
and U14153 (N_14153,N_6074,N_7724);
or U14154 (N_14154,N_7921,N_9694);
nor U14155 (N_14155,N_7886,N_9210);
nand U14156 (N_14156,N_5310,N_8075);
xor U14157 (N_14157,N_7297,N_9099);
nor U14158 (N_14158,N_7937,N_6127);
xor U14159 (N_14159,N_5616,N_8122);
and U14160 (N_14160,N_8382,N_5655);
nand U14161 (N_14161,N_6022,N_6811);
or U14162 (N_14162,N_6800,N_9973);
or U14163 (N_14163,N_6371,N_5035);
xor U14164 (N_14164,N_5655,N_9202);
and U14165 (N_14165,N_5634,N_8173);
and U14166 (N_14166,N_8620,N_9166);
or U14167 (N_14167,N_9904,N_7379);
and U14168 (N_14168,N_5053,N_6221);
or U14169 (N_14169,N_8438,N_5974);
nand U14170 (N_14170,N_7026,N_8557);
xor U14171 (N_14171,N_9869,N_7957);
or U14172 (N_14172,N_9610,N_7684);
or U14173 (N_14173,N_5784,N_8262);
and U14174 (N_14174,N_9141,N_8181);
nand U14175 (N_14175,N_8015,N_8436);
nand U14176 (N_14176,N_5845,N_7498);
nor U14177 (N_14177,N_8915,N_6331);
or U14178 (N_14178,N_7045,N_8449);
nor U14179 (N_14179,N_9444,N_9671);
nand U14180 (N_14180,N_5409,N_5888);
nand U14181 (N_14181,N_9566,N_8285);
nand U14182 (N_14182,N_5222,N_9458);
or U14183 (N_14183,N_6619,N_9010);
or U14184 (N_14184,N_8213,N_6897);
and U14185 (N_14185,N_9576,N_6217);
or U14186 (N_14186,N_5987,N_8335);
and U14187 (N_14187,N_5883,N_9379);
xnor U14188 (N_14188,N_5231,N_7865);
and U14189 (N_14189,N_8824,N_9837);
or U14190 (N_14190,N_7327,N_8411);
xor U14191 (N_14191,N_6125,N_6986);
and U14192 (N_14192,N_5475,N_8092);
and U14193 (N_14193,N_6727,N_7980);
xor U14194 (N_14194,N_5811,N_9759);
or U14195 (N_14195,N_6868,N_8248);
nand U14196 (N_14196,N_5573,N_8682);
nor U14197 (N_14197,N_7420,N_8478);
or U14198 (N_14198,N_8424,N_6536);
nand U14199 (N_14199,N_6300,N_9473);
nand U14200 (N_14200,N_8939,N_5474);
xor U14201 (N_14201,N_8474,N_6694);
or U14202 (N_14202,N_7454,N_6393);
or U14203 (N_14203,N_8853,N_5942);
or U14204 (N_14204,N_5084,N_7327);
and U14205 (N_14205,N_8204,N_8994);
or U14206 (N_14206,N_8305,N_5895);
nand U14207 (N_14207,N_6635,N_6074);
nand U14208 (N_14208,N_7092,N_6119);
and U14209 (N_14209,N_9673,N_7346);
nand U14210 (N_14210,N_9180,N_8863);
nand U14211 (N_14211,N_6909,N_6460);
and U14212 (N_14212,N_8532,N_8921);
nor U14213 (N_14213,N_6831,N_7342);
nor U14214 (N_14214,N_5787,N_5511);
nor U14215 (N_14215,N_8295,N_8267);
nand U14216 (N_14216,N_9890,N_8485);
nand U14217 (N_14217,N_9907,N_5871);
or U14218 (N_14218,N_6004,N_8060);
or U14219 (N_14219,N_5980,N_7376);
and U14220 (N_14220,N_8721,N_6640);
and U14221 (N_14221,N_8455,N_6444);
nor U14222 (N_14222,N_6056,N_5956);
nor U14223 (N_14223,N_5644,N_9084);
nor U14224 (N_14224,N_8708,N_8939);
xor U14225 (N_14225,N_5647,N_6170);
and U14226 (N_14226,N_5329,N_7012);
nand U14227 (N_14227,N_9195,N_5260);
xor U14228 (N_14228,N_8677,N_6326);
or U14229 (N_14229,N_7436,N_9341);
xor U14230 (N_14230,N_6308,N_5835);
nand U14231 (N_14231,N_8172,N_6185);
or U14232 (N_14232,N_8806,N_9406);
nand U14233 (N_14233,N_9654,N_8147);
nor U14234 (N_14234,N_7727,N_8485);
and U14235 (N_14235,N_5334,N_9816);
xor U14236 (N_14236,N_8813,N_7367);
nor U14237 (N_14237,N_7019,N_8994);
and U14238 (N_14238,N_6063,N_5162);
xor U14239 (N_14239,N_5638,N_7176);
xnor U14240 (N_14240,N_6232,N_6014);
nor U14241 (N_14241,N_9495,N_8217);
nand U14242 (N_14242,N_6860,N_6487);
nor U14243 (N_14243,N_8152,N_9055);
nor U14244 (N_14244,N_5735,N_9300);
nor U14245 (N_14245,N_8970,N_8862);
nand U14246 (N_14246,N_9006,N_5382);
or U14247 (N_14247,N_8004,N_8574);
or U14248 (N_14248,N_8858,N_6128);
nand U14249 (N_14249,N_8543,N_8127);
or U14250 (N_14250,N_9136,N_5560);
nor U14251 (N_14251,N_7194,N_7203);
nand U14252 (N_14252,N_6633,N_9849);
nand U14253 (N_14253,N_6311,N_8142);
nand U14254 (N_14254,N_9416,N_5054);
and U14255 (N_14255,N_6963,N_6853);
nand U14256 (N_14256,N_9954,N_7216);
and U14257 (N_14257,N_5962,N_5062);
and U14258 (N_14258,N_5985,N_7613);
nand U14259 (N_14259,N_5677,N_9813);
and U14260 (N_14260,N_9720,N_7038);
or U14261 (N_14261,N_6908,N_8099);
nor U14262 (N_14262,N_6756,N_6107);
xor U14263 (N_14263,N_6912,N_8240);
and U14264 (N_14264,N_5461,N_7776);
or U14265 (N_14265,N_8063,N_8874);
and U14266 (N_14266,N_8106,N_7796);
xnor U14267 (N_14267,N_8569,N_9990);
and U14268 (N_14268,N_9418,N_8061);
or U14269 (N_14269,N_5743,N_7354);
nor U14270 (N_14270,N_5573,N_7465);
and U14271 (N_14271,N_7001,N_8321);
nand U14272 (N_14272,N_9019,N_9383);
xnor U14273 (N_14273,N_6119,N_6405);
and U14274 (N_14274,N_8410,N_8753);
or U14275 (N_14275,N_6000,N_7167);
and U14276 (N_14276,N_7075,N_8689);
nand U14277 (N_14277,N_5883,N_6494);
nor U14278 (N_14278,N_6656,N_8963);
and U14279 (N_14279,N_7311,N_5286);
and U14280 (N_14280,N_8232,N_7846);
or U14281 (N_14281,N_7970,N_8232);
nand U14282 (N_14282,N_5488,N_9991);
nand U14283 (N_14283,N_6563,N_6520);
and U14284 (N_14284,N_8554,N_5239);
and U14285 (N_14285,N_6812,N_6709);
or U14286 (N_14286,N_9538,N_7009);
nor U14287 (N_14287,N_5529,N_5972);
and U14288 (N_14288,N_7330,N_6618);
and U14289 (N_14289,N_6647,N_8071);
nor U14290 (N_14290,N_7874,N_6030);
nand U14291 (N_14291,N_6844,N_8442);
nand U14292 (N_14292,N_7717,N_5053);
or U14293 (N_14293,N_5731,N_9127);
xnor U14294 (N_14294,N_7507,N_6441);
nand U14295 (N_14295,N_5681,N_7435);
nor U14296 (N_14296,N_9213,N_8131);
or U14297 (N_14297,N_7146,N_9924);
or U14298 (N_14298,N_6857,N_8140);
or U14299 (N_14299,N_7473,N_5532);
and U14300 (N_14300,N_8935,N_7672);
nor U14301 (N_14301,N_5992,N_6434);
or U14302 (N_14302,N_6338,N_6523);
and U14303 (N_14303,N_8973,N_7627);
or U14304 (N_14304,N_7339,N_6377);
nor U14305 (N_14305,N_6038,N_6131);
or U14306 (N_14306,N_6571,N_5891);
nor U14307 (N_14307,N_7482,N_8971);
or U14308 (N_14308,N_6364,N_9299);
nand U14309 (N_14309,N_7826,N_6432);
nand U14310 (N_14310,N_5938,N_8948);
nand U14311 (N_14311,N_5714,N_5937);
nor U14312 (N_14312,N_5895,N_8118);
nor U14313 (N_14313,N_8520,N_9408);
nor U14314 (N_14314,N_9010,N_7769);
and U14315 (N_14315,N_9373,N_8715);
nand U14316 (N_14316,N_9616,N_9107);
and U14317 (N_14317,N_6251,N_8371);
or U14318 (N_14318,N_9586,N_8131);
and U14319 (N_14319,N_8757,N_5992);
nor U14320 (N_14320,N_7483,N_7145);
and U14321 (N_14321,N_8468,N_6657);
nor U14322 (N_14322,N_7315,N_7905);
and U14323 (N_14323,N_8598,N_7730);
nand U14324 (N_14324,N_9929,N_6006);
nand U14325 (N_14325,N_8380,N_9110);
xor U14326 (N_14326,N_7271,N_6378);
or U14327 (N_14327,N_7795,N_6314);
and U14328 (N_14328,N_7510,N_8502);
and U14329 (N_14329,N_7481,N_8511);
nand U14330 (N_14330,N_6639,N_7769);
and U14331 (N_14331,N_6546,N_6596);
or U14332 (N_14332,N_6297,N_6361);
and U14333 (N_14333,N_6760,N_9765);
nor U14334 (N_14334,N_9539,N_7887);
nor U14335 (N_14335,N_9128,N_6223);
nor U14336 (N_14336,N_7495,N_8690);
or U14337 (N_14337,N_6902,N_9972);
or U14338 (N_14338,N_5581,N_9783);
nand U14339 (N_14339,N_8651,N_7199);
and U14340 (N_14340,N_5382,N_6335);
nor U14341 (N_14341,N_6588,N_8656);
and U14342 (N_14342,N_9925,N_9932);
nand U14343 (N_14343,N_5944,N_8137);
nor U14344 (N_14344,N_9470,N_8590);
nand U14345 (N_14345,N_9539,N_5825);
xnor U14346 (N_14346,N_6482,N_5907);
nor U14347 (N_14347,N_6637,N_5163);
or U14348 (N_14348,N_7230,N_5899);
nor U14349 (N_14349,N_5040,N_9065);
or U14350 (N_14350,N_9991,N_7328);
nor U14351 (N_14351,N_8021,N_7190);
nand U14352 (N_14352,N_8765,N_9198);
nand U14353 (N_14353,N_5308,N_9849);
nand U14354 (N_14354,N_7212,N_6724);
or U14355 (N_14355,N_9344,N_6626);
xor U14356 (N_14356,N_8084,N_6993);
and U14357 (N_14357,N_5797,N_6229);
or U14358 (N_14358,N_9390,N_8584);
or U14359 (N_14359,N_9866,N_6394);
or U14360 (N_14360,N_9686,N_8628);
nor U14361 (N_14361,N_7869,N_7128);
or U14362 (N_14362,N_9369,N_9727);
or U14363 (N_14363,N_5993,N_8426);
and U14364 (N_14364,N_5078,N_6795);
nand U14365 (N_14365,N_9279,N_8098);
nor U14366 (N_14366,N_7952,N_8733);
or U14367 (N_14367,N_9110,N_8064);
nand U14368 (N_14368,N_6971,N_9480);
or U14369 (N_14369,N_7585,N_5270);
xor U14370 (N_14370,N_6246,N_7040);
nand U14371 (N_14371,N_8086,N_9840);
nor U14372 (N_14372,N_8144,N_6391);
nand U14373 (N_14373,N_6129,N_5581);
nand U14374 (N_14374,N_8694,N_5211);
nand U14375 (N_14375,N_9538,N_6123);
or U14376 (N_14376,N_8793,N_7806);
nand U14377 (N_14377,N_5774,N_6879);
nor U14378 (N_14378,N_5886,N_9835);
nor U14379 (N_14379,N_8278,N_7917);
or U14380 (N_14380,N_7067,N_6421);
nor U14381 (N_14381,N_6068,N_8614);
or U14382 (N_14382,N_9089,N_7269);
nand U14383 (N_14383,N_5407,N_9493);
nor U14384 (N_14384,N_6579,N_9196);
and U14385 (N_14385,N_8393,N_6719);
nand U14386 (N_14386,N_6921,N_5337);
nand U14387 (N_14387,N_5662,N_9159);
nand U14388 (N_14388,N_8868,N_5860);
and U14389 (N_14389,N_9190,N_6041);
nand U14390 (N_14390,N_6830,N_6695);
nand U14391 (N_14391,N_8554,N_9553);
xnor U14392 (N_14392,N_5364,N_6290);
nor U14393 (N_14393,N_9559,N_6943);
and U14394 (N_14394,N_9562,N_5417);
xor U14395 (N_14395,N_8296,N_8631);
and U14396 (N_14396,N_7590,N_6404);
nand U14397 (N_14397,N_6492,N_9515);
and U14398 (N_14398,N_5521,N_8328);
nand U14399 (N_14399,N_9563,N_9731);
and U14400 (N_14400,N_7136,N_9633);
or U14401 (N_14401,N_7393,N_6090);
xnor U14402 (N_14402,N_7962,N_8837);
xnor U14403 (N_14403,N_5908,N_9997);
and U14404 (N_14404,N_9670,N_9100);
nand U14405 (N_14405,N_5217,N_9672);
nand U14406 (N_14406,N_7874,N_6689);
xor U14407 (N_14407,N_5528,N_9183);
or U14408 (N_14408,N_5149,N_5783);
and U14409 (N_14409,N_9452,N_6762);
xnor U14410 (N_14410,N_9312,N_9585);
or U14411 (N_14411,N_5490,N_9353);
and U14412 (N_14412,N_9468,N_8121);
nand U14413 (N_14413,N_6582,N_5809);
or U14414 (N_14414,N_8236,N_5833);
or U14415 (N_14415,N_6052,N_7869);
nand U14416 (N_14416,N_9211,N_9691);
and U14417 (N_14417,N_9852,N_9995);
nand U14418 (N_14418,N_8334,N_6857);
or U14419 (N_14419,N_9272,N_7986);
and U14420 (N_14420,N_7603,N_5235);
or U14421 (N_14421,N_7025,N_5199);
nor U14422 (N_14422,N_8502,N_8789);
and U14423 (N_14423,N_9129,N_8267);
or U14424 (N_14424,N_8529,N_7494);
or U14425 (N_14425,N_7869,N_6299);
nand U14426 (N_14426,N_9420,N_8636);
or U14427 (N_14427,N_9877,N_6837);
nand U14428 (N_14428,N_9644,N_5815);
xnor U14429 (N_14429,N_8961,N_8919);
nand U14430 (N_14430,N_9285,N_7623);
or U14431 (N_14431,N_7630,N_9263);
nor U14432 (N_14432,N_6833,N_9453);
nand U14433 (N_14433,N_5666,N_7487);
nand U14434 (N_14434,N_8240,N_7994);
or U14435 (N_14435,N_8628,N_8497);
nor U14436 (N_14436,N_6463,N_9120);
and U14437 (N_14437,N_7368,N_6457);
nand U14438 (N_14438,N_9976,N_7651);
nor U14439 (N_14439,N_9662,N_6255);
or U14440 (N_14440,N_5041,N_8875);
or U14441 (N_14441,N_5455,N_7257);
xor U14442 (N_14442,N_6843,N_9071);
nand U14443 (N_14443,N_8540,N_9754);
and U14444 (N_14444,N_7947,N_5656);
and U14445 (N_14445,N_8776,N_5385);
and U14446 (N_14446,N_8776,N_9948);
or U14447 (N_14447,N_5531,N_6349);
nor U14448 (N_14448,N_6671,N_5182);
xor U14449 (N_14449,N_8685,N_5465);
and U14450 (N_14450,N_5651,N_6438);
or U14451 (N_14451,N_6350,N_9404);
and U14452 (N_14452,N_9587,N_8547);
or U14453 (N_14453,N_9098,N_9603);
nor U14454 (N_14454,N_8965,N_9322);
nor U14455 (N_14455,N_5689,N_6099);
or U14456 (N_14456,N_8675,N_6832);
nor U14457 (N_14457,N_8718,N_8909);
xnor U14458 (N_14458,N_6090,N_6884);
nor U14459 (N_14459,N_5413,N_9738);
nand U14460 (N_14460,N_8119,N_8716);
nand U14461 (N_14461,N_8149,N_5474);
or U14462 (N_14462,N_5555,N_9570);
and U14463 (N_14463,N_6176,N_9617);
or U14464 (N_14464,N_9796,N_8882);
xor U14465 (N_14465,N_9680,N_8870);
nand U14466 (N_14466,N_6924,N_6121);
and U14467 (N_14467,N_5392,N_6754);
nand U14468 (N_14468,N_8003,N_9083);
nand U14469 (N_14469,N_8872,N_8446);
or U14470 (N_14470,N_5462,N_9686);
or U14471 (N_14471,N_6064,N_6453);
nor U14472 (N_14472,N_5453,N_6817);
or U14473 (N_14473,N_9016,N_7844);
or U14474 (N_14474,N_8558,N_6067);
and U14475 (N_14475,N_6542,N_7969);
nor U14476 (N_14476,N_6179,N_5290);
nor U14477 (N_14477,N_8266,N_8481);
nand U14478 (N_14478,N_6373,N_8084);
nand U14479 (N_14479,N_5185,N_6331);
nor U14480 (N_14480,N_7482,N_8555);
nand U14481 (N_14481,N_6343,N_6525);
nor U14482 (N_14482,N_5627,N_8854);
xor U14483 (N_14483,N_9700,N_7748);
nor U14484 (N_14484,N_9359,N_5490);
or U14485 (N_14485,N_9640,N_9976);
nor U14486 (N_14486,N_6906,N_7472);
or U14487 (N_14487,N_8748,N_6616);
or U14488 (N_14488,N_9465,N_5247);
or U14489 (N_14489,N_7168,N_8370);
nor U14490 (N_14490,N_8642,N_8957);
and U14491 (N_14491,N_9117,N_9962);
nor U14492 (N_14492,N_7342,N_9096);
or U14493 (N_14493,N_9591,N_8735);
nor U14494 (N_14494,N_8666,N_8401);
nand U14495 (N_14495,N_9341,N_9365);
or U14496 (N_14496,N_6331,N_9358);
nor U14497 (N_14497,N_9123,N_5396);
and U14498 (N_14498,N_8554,N_7781);
nand U14499 (N_14499,N_8598,N_7006);
or U14500 (N_14500,N_8373,N_6058);
or U14501 (N_14501,N_5925,N_9340);
or U14502 (N_14502,N_6518,N_7515);
or U14503 (N_14503,N_5289,N_6213);
and U14504 (N_14504,N_9191,N_7584);
xor U14505 (N_14505,N_5925,N_8146);
and U14506 (N_14506,N_7986,N_6472);
nand U14507 (N_14507,N_9012,N_5969);
or U14508 (N_14508,N_7584,N_5888);
or U14509 (N_14509,N_7655,N_5591);
and U14510 (N_14510,N_6173,N_9728);
nor U14511 (N_14511,N_8603,N_5793);
and U14512 (N_14512,N_8862,N_7087);
nand U14513 (N_14513,N_5856,N_8966);
or U14514 (N_14514,N_8637,N_8388);
nor U14515 (N_14515,N_5833,N_7854);
nand U14516 (N_14516,N_6624,N_8083);
nand U14517 (N_14517,N_5895,N_6449);
xnor U14518 (N_14518,N_8157,N_5202);
and U14519 (N_14519,N_7122,N_5116);
nor U14520 (N_14520,N_9342,N_5177);
and U14521 (N_14521,N_8821,N_6026);
xor U14522 (N_14522,N_7054,N_5844);
nand U14523 (N_14523,N_9788,N_9910);
nor U14524 (N_14524,N_8673,N_8605);
or U14525 (N_14525,N_9797,N_6414);
nor U14526 (N_14526,N_5434,N_9239);
or U14527 (N_14527,N_8714,N_8941);
nand U14528 (N_14528,N_7161,N_7724);
or U14529 (N_14529,N_6215,N_5335);
nor U14530 (N_14530,N_9983,N_8002);
or U14531 (N_14531,N_8346,N_8205);
or U14532 (N_14532,N_9864,N_9429);
and U14533 (N_14533,N_9651,N_9573);
nor U14534 (N_14534,N_9628,N_8874);
nor U14535 (N_14535,N_9769,N_9987);
and U14536 (N_14536,N_5756,N_8725);
or U14537 (N_14537,N_9725,N_7298);
nor U14538 (N_14538,N_8671,N_8544);
nand U14539 (N_14539,N_9913,N_5131);
xor U14540 (N_14540,N_8422,N_7318);
and U14541 (N_14541,N_6968,N_8728);
nand U14542 (N_14542,N_7870,N_6107);
and U14543 (N_14543,N_5754,N_6246);
or U14544 (N_14544,N_8535,N_8230);
nand U14545 (N_14545,N_5875,N_6139);
nand U14546 (N_14546,N_7928,N_6229);
and U14547 (N_14547,N_8702,N_7315);
nor U14548 (N_14548,N_9443,N_7416);
nor U14549 (N_14549,N_7913,N_7650);
or U14550 (N_14550,N_7011,N_8218);
xnor U14551 (N_14551,N_5645,N_8386);
and U14552 (N_14552,N_6923,N_7747);
nor U14553 (N_14553,N_9372,N_7856);
nand U14554 (N_14554,N_8930,N_8304);
and U14555 (N_14555,N_7432,N_6432);
nand U14556 (N_14556,N_9418,N_6520);
nand U14557 (N_14557,N_8291,N_7322);
and U14558 (N_14558,N_5000,N_9583);
xor U14559 (N_14559,N_8637,N_5164);
and U14560 (N_14560,N_8560,N_5633);
nand U14561 (N_14561,N_9692,N_6942);
and U14562 (N_14562,N_7830,N_9506);
or U14563 (N_14563,N_6100,N_5561);
nor U14564 (N_14564,N_5010,N_6464);
nor U14565 (N_14565,N_6815,N_7592);
xnor U14566 (N_14566,N_7471,N_5969);
nand U14567 (N_14567,N_5105,N_6253);
and U14568 (N_14568,N_6946,N_9375);
and U14569 (N_14569,N_5933,N_7642);
and U14570 (N_14570,N_7068,N_6701);
xor U14571 (N_14571,N_6961,N_6026);
and U14572 (N_14572,N_6121,N_5123);
and U14573 (N_14573,N_6762,N_9334);
nand U14574 (N_14574,N_5066,N_9138);
nand U14575 (N_14575,N_9348,N_7387);
and U14576 (N_14576,N_5049,N_6844);
nor U14577 (N_14577,N_5579,N_5293);
or U14578 (N_14578,N_7337,N_5069);
or U14579 (N_14579,N_5001,N_9658);
nor U14580 (N_14580,N_9931,N_7283);
or U14581 (N_14581,N_7892,N_6078);
nand U14582 (N_14582,N_9188,N_5722);
or U14583 (N_14583,N_5927,N_6802);
nor U14584 (N_14584,N_6128,N_8108);
nand U14585 (N_14585,N_5888,N_9156);
nand U14586 (N_14586,N_6286,N_7848);
nand U14587 (N_14587,N_8962,N_5106);
nand U14588 (N_14588,N_8883,N_7005);
xor U14589 (N_14589,N_5294,N_8375);
nor U14590 (N_14590,N_5982,N_9594);
or U14591 (N_14591,N_6600,N_5190);
nor U14592 (N_14592,N_8017,N_5772);
xnor U14593 (N_14593,N_7465,N_7505);
nand U14594 (N_14594,N_6654,N_9266);
or U14595 (N_14595,N_7757,N_9352);
xnor U14596 (N_14596,N_7690,N_8973);
or U14597 (N_14597,N_6689,N_6094);
nand U14598 (N_14598,N_7046,N_5445);
or U14599 (N_14599,N_5701,N_8230);
or U14600 (N_14600,N_8681,N_9214);
and U14601 (N_14601,N_8985,N_9579);
xor U14602 (N_14602,N_5548,N_8451);
or U14603 (N_14603,N_6128,N_9748);
nor U14604 (N_14604,N_9344,N_6499);
nor U14605 (N_14605,N_8314,N_8900);
xnor U14606 (N_14606,N_8135,N_8773);
nand U14607 (N_14607,N_9031,N_9199);
nor U14608 (N_14608,N_9527,N_6447);
nor U14609 (N_14609,N_8426,N_5529);
nand U14610 (N_14610,N_6573,N_5353);
and U14611 (N_14611,N_9981,N_9610);
nand U14612 (N_14612,N_7390,N_7658);
or U14613 (N_14613,N_9987,N_9517);
and U14614 (N_14614,N_7206,N_9041);
or U14615 (N_14615,N_7644,N_9529);
nand U14616 (N_14616,N_6762,N_5482);
and U14617 (N_14617,N_6281,N_6828);
nand U14618 (N_14618,N_6791,N_6739);
or U14619 (N_14619,N_5225,N_9653);
nor U14620 (N_14620,N_7740,N_6519);
nand U14621 (N_14621,N_7694,N_6063);
and U14622 (N_14622,N_9246,N_8722);
nor U14623 (N_14623,N_8707,N_8113);
xnor U14624 (N_14624,N_7092,N_9657);
and U14625 (N_14625,N_9085,N_7535);
nor U14626 (N_14626,N_5022,N_8467);
nand U14627 (N_14627,N_9266,N_7003);
nand U14628 (N_14628,N_5559,N_7043);
and U14629 (N_14629,N_5570,N_7013);
nor U14630 (N_14630,N_6615,N_9389);
xor U14631 (N_14631,N_8756,N_9417);
nand U14632 (N_14632,N_7433,N_5667);
or U14633 (N_14633,N_8428,N_7039);
or U14634 (N_14634,N_7125,N_9738);
and U14635 (N_14635,N_9778,N_9750);
xor U14636 (N_14636,N_5685,N_7277);
and U14637 (N_14637,N_7928,N_8496);
xnor U14638 (N_14638,N_7490,N_6667);
or U14639 (N_14639,N_5689,N_5307);
or U14640 (N_14640,N_7079,N_8129);
nor U14641 (N_14641,N_8425,N_8148);
nor U14642 (N_14642,N_9600,N_7435);
or U14643 (N_14643,N_9296,N_7292);
nor U14644 (N_14644,N_7670,N_7568);
nand U14645 (N_14645,N_7554,N_7097);
or U14646 (N_14646,N_5792,N_5438);
nand U14647 (N_14647,N_6488,N_8173);
nand U14648 (N_14648,N_9491,N_9279);
nor U14649 (N_14649,N_7981,N_5755);
or U14650 (N_14650,N_9660,N_6734);
and U14651 (N_14651,N_7477,N_5941);
and U14652 (N_14652,N_9486,N_7484);
xor U14653 (N_14653,N_5486,N_6090);
nor U14654 (N_14654,N_8128,N_9206);
xnor U14655 (N_14655,N_7795,N_9582);
and U14656 (N_14656,N_6658,N_8404);
nand U14657 (N_14657,N_5066,N_8471);
nor U14658 (N_14658,N_6125,N_9814);
nor U14659 (N_14659,N_8540,N_9996);
or U14660 (N_14660,N_8709,N_5066);
nand U14661 (N_14661,N_6364,N_9401);
nand U14662 (N_14662,N_6972,N_7391);
nand U14663 (N_14663,N_8889,N_8248);
or U14664 (N_14664,N_5596,N_5342);
or U14665 (N_14665,N_6809,N_9478);
and U14666 (N_14666,N_5916,N_5082);
nand U14667 (N_14667,N_6300,N_9116);
xnor U14668 (N_14668,N_8754,N_5917);
or U14669 (N_14669,N_9858,N_5095);
nor U14670 (N_14670,N_8745,N_8135);
and U14671 (N_14671,N_8469,N_6324);
nand U14672 (N_14672,N_8775,N_5366);
nand U14673 (N_14673,N_6173,N_9069);
nand U14674 (N_14674,N_6875,N_8820);
or U14675 (N_14675,N_5584,N_6877);
or U14676 (N_14676,N_7614,N_7686);
or U14677 (N_14677,N_6601,N_6592);
and U14678 (N_14678,N_7177,N_8924);
or U14679 (N_14679,N_6085,N_6714);
nand U14680 (N_14680,N_6257,N_6112);
nand U14681 (N_14681,N_6626,N_8812);
nor U14682 (N_14682,N_6883,N_9736);
and U14683 (N_14683,N_5283,N_5005);
and U14684 (N_14684,N_5797,N_7661);
nand U14685 (N_14685,N_8442,N_7027);
nand U14686 (N_14686,N_8301,N_8511);
and U14687 (N_14687,N_7516,N_9385);
or U14688 (N_14688,N_7726,N_8688);
nor U14689 (N_14689,N_9913,N_6710);
nor U14690 (N_14690,N_6080,N_6522);
nor U14691 (N_14691,N_6828,N_7003);
nand U14692 (N_14692,N_8064,N_6483);
or U14693 (N_14693,N_9119,N_8284);
nand U14694 (N_14694,N_7504,N_7213);
and U14695 (N_14695,N_9759,N_6505);
and U14696 (N_14696,N_8466,N_5440);
nand U14697 (N_14697,N_8776,N_7024);
or U14698 (N_14698,N_5086,N_8980);
and U14699 (N_14699,N_8663,N_7883);
or U14700 (N_14700,N_6212,N_7823);
nor U14701 (N_14701,N_6976,N_6487);
nor U14702 (N_14702,N_9859,N_6760);
nand U14703 (N_14703,N_6489,N_6754);
nor U14704 (N_14704,N_7532,N_5692);
nor U14705 (N_14705,N_7402,N_9569);
or U14706 (N_14706,N_9814,N_9492);
nor U14707 (N_14707,N_9373,N_7951);
or U14708 (N_14708,N_9395,N_5705);
xor U14709 (N_14709,N_8754,N_7604);
xor U14710 (N_14710,N_8841,N_6571);
and U14711 (N_14711,N_5342,N_7457);
and U14712 (N_14712,N_5113,N_9276);
and U14713 (N_14713,N_6376,N_9054);
nor U14714 (N_14714,N_9746,N_5951);
nor U14715 (N_14715,N_6770,N_6838);
nor U14716 (N_14716,N_5491,N_8994);
nor U14717 (N_14717,N_7856,N_9309);
and U14718 (N_14718,N_5033,N_7852);
or U14719 (N_14719,N_7678,N_9671);
nand U14720 (N_14720,N_9764,N_7123);
and U14721 (N_14721,N_9216,N_8245);
nand U14722 (N_14722,N_5442,N_6088);
or U14723 (N_14723,N_5771,N_6066);
nor U14724 (N_14724,N_7461,N_7049);
and U14725 (N_14725,N_6563,N_5640);
and U14726 (N_14726,N_5447,N_6145);
and U14727 (N_14727,N_7306,N_7356);
and U14728 (N_14728,N_6401,N_5310);
nor U14729 (N_14729,N_5482,N_6960);
or U14730 (N_14730,N_8345,N_6749);
or U14731 (N_14731,N_8125,N_7225);
nand U14732 (N_14732,N_6102,N_6365);
xor U14733 (N_14733,N_6000,N_9235);
xnor U14734 (N_14734,N_5225,N_6590);
or U14735 (N_14735,N_9625,N_8250);
nor U14736 (N_14736,N_7232,N_9894);
and U14737 (N_14737,N_8047,N_7956);
or U14738 (N_14738,N_6438,N_8383);
nor U14739 (N_14739,N_9509,N_6354);
nand U14740 (N_14740,N_5554,N_5801);
or U14741 (N_14741,N_9570,N_5348);
nor U14742 (N_14742,N_7994,N_6947);
xor U14743 (N_14743,N_7629,N_5909);
xor U14744 (N_14744,N_5931,N_7685);
or U14745 (N_14745,N_6667,N_7508);
and U14746 (N_14746,N_9493,N_8179);
or U14747 (N_14747,N_6048,N_7951);
nor U14748 (N_14748,N_8761,N_6362);
nor U14749 (N_14749,N_8256,N_8610);
and U14750 (N_14750,N_7086,N_8240);
nor U14751 (N_14751,N_9765,N_6611);
xor U14752 (N_14752,N_6344,N_9160);
and U14753 (N_14753,N_9457,N_6168);
nand U14754 (N_14754,N_7426,N_6305);
nand U14755 (N_14755,N_5624,N_9766);
xnor U14756 (N_14756,N_5222,N_6505);
and U14757 (N_14757,N_5988,N_8054);
and U14758 (N_14758,N_6462,N_9771);
and U14759 (N_14759,N_9091,N_9219);
and U14760 (N_14760,N_7521,N_9879);
nor U14761 (N_14761,N_9895,N_6521);
nand U14762 (N_14762,N_8533,N_6279);
xnor U14763 (N_14763,N_9976,N_9712);
and U14764 (N_14764,N_6534,N_6492);
or U14765 (N_14765,N_5994,N_8946);
and U14766 (N_14766,N_6650,N_8893);
nand U14767 (N_14767,N_8687,N_5813);
or U14768 (N_14768,N_7790,N_5491);
and U14769 (N_14769,N_5363,N_7012);
or U14770 (N_14770,N_6548,N_6883);
nor U14771 (N_14771,N_6443,N_8224);
and U14772 (N_14772,N_6006,N_6925);
and U14773 (N_14773,N_6743,N_6995);
nor U14774 (N_14774,N_8724,N_6176);
or U14775 (N_14775,N_8055,N_8813);
xor U14776 (N_14776,N_9639,N_5884);
nand U14777 (N_14777,N_5498,N_9513);
nand U14778 (N_14778,N_7125,N_7983);
nor U14779 (N_14779,N_5099,N_7569);
or U14780 (N_14780,N_5845,N_7444);
nor U14781 (N_14781,N_6269,N_8191);
xor U14782 (N_14782,N_5744,N_7231);
and U14783 (N_14783,N_5836,N_8935);
nor U14784 (N_14784,N_7918,N_7829);
and U14785 (N_14785,N_5716,N_5128);
or U14786 (N_14786,N_7243,N_5741);
and U14787 (N_14787,N_5331,N_8517);
nor U14788 (N_14788,N_8601,N_8606);
and U14789 (N_14789,N_5754,N_5124);
nor U14790 (N_14790,N_6324,N_5487);
nand U14791 (N_14791,N_8728,N_8322);
or U14792 (N_14792,N_8750,N_7804);
and U14793 (N_14793,N_7670,N_6155);
nor U14794 (N_14794,N_8328,N_6743);
xor U14795 (N_14795,N_7328,N_8218);
and U14796 (N_14796,N_5259,N_8442);
nor U14797 (N_14797,N_6892,N_8143);
nand U14798 (N_14798,N_7952,N_7372);
xor U14799 (N_14799,N_5117,N_6885);
nand U14800 (N_14800,N_8153,N_6654);
and U14801 (N_14801,N_8690,N_7962);
or U14802 (N_14802,N_7862,N_6572);
nand U14803 (N_14803,N_9360,N_9366);
and U14804 (N_14804,N_6621,N_8422);
and U14805 (N_14805,N_7415,N_8826);
xor U14806 (N_14806,N_6632,N_7813);
or U14807 (N_14807,N_6342,N_7652);
nand U14808 (N_14808,N_6276,N_7854);
and U14809 (N_14809,N_9988,N_9943);
and U14810 (N_14810,N_8367,N_7590);
or U14811 (N_14811,N_5516,N_8409);
and U14812 (N_14812,N_6889,N_9178);
or U14813 (N_14813,N_8790,N_9686);
and U14814 (N_14814,N_9466,N_5985);
nand U14815 (N_14815,N_9107,N_7851);
or U14816 (N_14816,N_7730,N_5202);
nor U14817 (N_14817,N_5824,N_5109);
or U14818 (N_14818,N_6275,N_7662);
nor U14819 (N_14819,N_9789,N_5956);
nor U14820 (N_14820,N_6848,N_9647);
nor U14821 (N_14821,N_5100,N_8464);
or U14822 (N_14822,N_9622,N_5135);
and U14823 (N_14823,N_7172,N_7114);
nor U14824 (N_14824,N_6382,N_9593);
or U14825 (N_14825,N_7745,N_5747);
nor U14826 (N_14826,N_9172,N_5345);
and U14827 (N_14827,N_9415,N_5297);
and U14828 (N_14828,N_7643,N_6178);
and U14829 (N_14829,N_7956,N_6663);
nor U14830 (N_14830,N_5729,N_7161);
or U14831 (N_14831,N_9102,N_5504);
nor U14832 (N_14832,N_7762,N_9142);
and U14833 (N_14833,N_8359,N_5225);
and U14834 (N_14834,N_8141,N_7187);
xnor U14835 (N_14835,N_8105,N_5023);
and U14836 (N_14836,N_7991,N_6034);
nand U14837 (N_14837,N_5322,N_5674);
or U14838 (N_14838,N_5655,N_9139);
and U14839 (N_14839,N_9230,N_5810);
or U14840 (N_14840,N_8655,N_6077);
or U14841 (N_14841,N_8896,N_7778);
or U14842 (N_14842,N_8693,N_6201);
nand U14843 (N_14843,N_7901,N_9228);
or U14844 (N_14844,N_7973,N_9071);
xor U14845 (N_14845,N_9974,N_8472);
or U14846 (N_14846,N_5002,N_5416);
or U14847 (N_14847,N_8561,N_8693);
nor U14848 (N_14848,N_9281,N_9650);
nand U14849 (N_14849,N_8886,N_9661);
or U14850 (N_14850,N_6483,N_7774);
or U14851 (N_14851,N_6796,N_9104);
nand U14852 (N_14852,N_7251,N_6723);
nor U14853 (N_14853,N_5066,N_8811);
nor U14854 (N_14854,N_6343,N_9880);
and U14855 (N_14855,N_6028,N_6869);
nor U14856 (N_14856,N_8057,N_6179);
or U14857 (N_14857,N_9956,N_5891);
nor U14858 (N_14858,N_9909,N_7419);
nand U14859 (N_14859,N_9088,N_9862);
nand U14860 (N_14860,N_5463,N_8877);
nor U14861 (N_14861,N_9790,N_7716);
and U14862 (N_14862,N_6901,N_7679);
or U14863 (N_14863,N_8083,N_5374);
nand U14864 (N_14864,N_7932,N_7389);
xnor U14865 (N_14865,N_7809,N_9780);
and U14866 (N_14866,N_5325,N_5287);
xnor U14867 (N_14867,N_8666,N_5395);
and U14868 (N_14868,N_6666,N_9744);
nor U14869 (N_14869,N_5119,N_8261);
and U14870 (N_14870,N_6294,N_8602);
nor U14871 (N_14871,N_5138,N_9216);
and U14872 (N_14872,N_8033,N_8965);
nor U14873 (N_14873,N_5008,N_7832);
nor U14874 (N_14874,N_6568,N_9356);
nor U14875 (N_14875,N_6601,N_8164);
or U14876 (N_14876,N_9917,N_5371);
nor U14877 (N_14877,N_9629,N_7809);
or U14878 (N_14878,N_5542,N_9668);
xnor U14879 (N_14879,N_6125,N_9046);
nand U14880 (N_14880,N_7764,N_7187);
nand U14881 (N_14881,N_7638,N_5722);
or U14882 (N_14882,N_6542,N_5379);
or U14883 (N_14883,N_6728,N_5156);
or U14884 (N_14884,N_8260,N_8620);
or U14885 (N_14885,N_5542,N_5954);
nor U14886 (N_14886,N_9649,N_9145);
and U14887 (N_14887,N_5049,N_5943);
and U14888 (N_14888,N_6231,N_9886);
and U14889 (N_14889,N_8037,N_7177);
nor U14890 (N_14890,N_8376,N_6572);
nand U14891 (N_14891,N_6479,N_5403);
nand U14892 (N_14892,N_8348,N_8706);
xor U14893 (N_14893,N_9099,N_9306);
or U14894 (N_14894,N_8532,N_7489);
or U14895 (N_14895,N_9730,N_9764);
or U14896 (N_14896,N_7626,N_6289);
nor U14897 (N_14897,N_7335,N_6756);
nand U14898 (N_14898,N_8912,N_7020);
nand U14899 (N_14899,N_6155,N_5383);
nand U14900 (N_14900,N_7949,N_6343);
nor U14901 (N_14901,N_5018,N_8681);
or U14902 (N_14902,N_8864,N_5895);
xor U14903 (N_14903,N_8639,N_9401);
and U14904 (N_14904,N_5496,N_8982);
and U14905 (N_14905,N_7929,N_8498);
or U14906 (N_14906,N_5219,N_9327);
nand U14907 (N_14907,N_5670,N_9157);
and U14908 (N_14908,N_7045,N_7399);
or U14909 (N_14909,N_7689,N_6491);
or U14910 (N_14910,N_9106,N_7604);
nand U14911 (N_14911,N_9787,N_8356);
xnor U14912 (N_14912,N_6170,N_5216);
or U14913 (N_14913,N_6383,N_9942);
xor U14914 (N_14914,N_8504,N_6127);
or U14915 (N_14915,N_9980,N_5307);
and U14916 (N_14916,N_8780,N_5153);
nand U14917 (N_14917,N_9870,N_7590);
nand U14918 (N_14918,N_8932,N_9207);
nand U14919 (N_14919,N_5054,N_5467);
and U14920 (N_14920,N_7751,N_8944);
or U14921 (N_14921,N_7358,N_9208);
and U14922 (N_14922,N_6238,N_5992);
and U14923 (N_14923,N_9235,N_8712);
nor U14924 (N_14924,N_5163,N_9719);
nor U14925 (N_14925,N_6138,N_9879);
nor U14926 (N_14926,N_5241,N_9794);
and U14927 (N_14927,N_8334,N_8683);
nand U14928 (N_14928,N_9193,N_7286);
nor U14929 (N_14929,N_9382,N_6851);
and U14930 (N_14930,N_5431,N_5083);
nand U14931 (N_14931,N_7643,N_8003);
nor U14932 (N_14932,N_7269,N_6804);
or U14933 (N_14933,N_8802,N_5361);
or U14934 (N_14934,N_7943,N_7537);
nand U14935 (N_14935,N_7526,N_9412);
and U14936 (N_14936,N_9152,N_9414);
nand U14937 (N_14937,N_8434,N_9932);
nand U14938 (N_14938,N_7764,N_8088);
xnor U14939 (N_14939,N_9612,N_7029);
or U14940 (N_14940,N_5618,N_9236);
or U14941 (N_14941,N_8726,N_9176);
xor U14942 (N_14942,N_5605,N_7209);
nand U14943 (N_14943,N_5011,N_7002);
nand U14944 (N_14944,N_5313,N_9669);
xnor U14945 (N_14945,N_5108,N_5206);
or U14946 (N_14946,N_6735,N_5430);
nor U14947 (N_14947,N_6960,N_5101);
nand U14948 (N_14948,N_9277,N_5076);
xnor U14949 (N_14949,N_7046,N_8080);
or U14950 (N_14950,N_5499,N_8809);
nand U14951 (N_14951,N_9379,N_9017);
or U14952 (N_14952,N_6528,N_5080);
xor U14953 (N_14953,N_7426,N_8332);
or U14954 (N_14954,N_8849,N_9263);
or U14955 (N_14955,N_8218,N_6249);
and U14956 (N_14956,N_9699,N_7461);
nand U14957 (N_14957,N_6230,N_9709);
or U14958 (N_14958,N_7837,N_6369);
nand U14959 (N_14959,N_9507,N_7853);
or U14960 (N_14960,N_8677,N_5432);
nand U14961 (N_14961,N_6650,N_5586);
nand U14962 (N_14962,N_9379,N_9162);
nor U14963 (N_14963,N_8082,N_8407);
nor U14964 (N_14964,N_5460,N_6947);
nand U14965 (N_14965,N_6154,N_6075);
or U14966 (N_14966,N_6777,N_6112);
xnor U14967 (N_14967,N_8059,N_7678);
nand U14968 (N_14968,N_5445,N_6873);
or U14969 (N_14969,N_6662,N_9697);
nor U14970 (N_14970,N_6353,N_7859);
nand U14971 (N_14971,N_6683,N_5475);
or U14972 (N_14972,N_8145,N_7057);
xor U14973 (N_14973,N_5891,N_7680);
nand U14974 (N_14974,N_5533,N_7071);
nor U14975 (N_14975,N_9453,N_5092);
or U14976 (N_14976,N_8045,N_8260);
or U14977 (N_14977,N_8050,N_6024);
nor U14978 (N_14978,N_6387,N_7421);
nor U14979 (N_14979,N_6245,N_5844);
nor U14980 (N_14980,N_9567,N_7943);
nand U14981 (N_14981,N_7444,N_5818);
xor U14982 (N_14982,N_9901,N_8069);
or U14983 (N_14983,N_9200,N_7872);
and U14984 (N_14984,N_5088,N_7135);
or U14985 (N_14985,N_7469,N_5257);
and U14986 (N_14986,N_8448,N_5187);
or U14987 (N_14987,N_9067,N_9155);
and U14988 (N_14988,N_7013,N_7489);
and U14989 (N_14989,N_9896,N_8760);
nand U14990 (N_14990,N_9089,N_5605);
and U14991 (N_14991,N_7878,N_5156);
and U14992 (N_14992,N_5026,N_8176);
nand U14993 (N_14993,N_6498,N_8613);
and U14994 (N_14994,N_9532,N_8467);
and U14995 (N_14995,N_7783,N_7613);
nor U14996 (N_14996,N_9970,N_6424);
and U14997 (N_14997,N_6164,N_9896);
nand U14998 (N_14998,N_6285,N_6281);
nand U14999 (N_14999,N_5213,N_9515);
xor U15000 (N_15000,N_14490,N_13497);
or U15001 (N_15001,N_13565,N_13586);
nor U15002 (N_15002,N_13871,N_11280);
and U15003 (N_15003,N_12582,N_14056);
nand U15004 (N_15004,N_11504,N_13368);
or U15005 (N_15005,N_13474,N_13700);
or U15006 (N_15006,N_12029,N_13215);
nor U15007 (N_15007,N_14463,N_14637);
and U15008 (N_15008,N_12228,N_10132);
and U15009 (N_15009,N_14100,N_14603);
nor U15010 (N_15010,N_13008,N_11164);
nand U15011 (N_15011,N_14210,N_10529);
xnor U15012 (N_15012,N_14966,N_11069);
and U15013 (N_15013,N_13346,N_14990);
or U15014 (N_15014,N_14604,N_13694);
and U15015 (N_15015,N_14267,N_10844);
nor U15016 (N_15016,N_14938,N_12539);
and U15017 (N_15017,N_14118,N_12400);
nor U15018 (N_15018,N_13438,N_13333);
nor U15019 (N_15019,N_11867,N_12177);
and U15020 (N_15020,N_10145,N_12363);
or U15021 (N_15021,N_10937,N_11927);
nor U15022 (N_15022,N_11200,N_13145);
nor U15023 (N_15023,N_14211,N_14883);
or U15024 (N_15024,N_14716,N_11852);
nand U15025 (N_15025,N_12050,N_12927);
nor U15026 (N_15026,N_10900,N_14583);
nor U15027 (N_15027,N_11766,N_10488);
nand U15028 (N_15028,N_14703,N_10958);
nand U15029 (N_15029,N_13712,N_12425);
nand U15030 (N_15030,N_13951,N_13257);
nor U15031 (N_15031,N_12312,N_13983);
and U15032 (N_15032,N_14536,N_14471);
and U15033 (N_15033,N_14892,N_10765);
and U15034 (N_15034,N_11144,N_12951);
or U15035 (N_15035,N_11547,N_11061);
nand U15036 (N_15036,N_11509,N_12007);
nand U15037 (N_15037,N_13006,N_10184);
or U15038 (N_15038,N_11461,N_10157);
or U15039 (N_15039,N_13188,N_11954);
and U15040 (N_15040,N_12067,N_13042);
nand U15041 (N_15041,N_11009,N_14717);
and U15042 (N_15042,N_12465,N_11578);
nand U15043 (N_15043,N_11301,N_12702);
nand U15044 (N_15044,N_13773,N_12795);
or U15045 (N_15045,N_10377,N_11843);
or U15046 (N_15046,N_14364,N_13220);
nor U15047 (N_15047,N_11646,N_10589);
nand U15048 (N_15048,N_13915,N_10244);
and U15049 (N_15049,N_10693,N_11528);
and U15050 (N_15050,N_11500,N_12506);
nor U15051 (N_15051,N_10829,N_11266);
nand U15052 (N_15052,N_13293,N_12227);
nor U15053 (N_15053,N_11659,N_10426);
nand U15054 (N_15054,N_12397,N_12743);
or U15055 (N_15055,N_14707,N_13051);
and U15056 (N_15056,N_12804,N_13989);
nand U15057 (N_15057,N_12975,N_13945);
xnor U15058 (N_15058,N_11366,N_11903);
or U15059 (N_15059,N_13988,N_14189);
nor U15060 (N_15060,N_11580,N_14355);
xnor U15061 (N_15061,N_14578,N_14154);
or U15062 (N_15062,N_12877,N_13764);
or U15063 (N_15063,N_12640,N_12149);
and U15064 (N_15064,N_11238,N_10740);
nor U15065 (N_15065,N_13500,N_11541);
and U15066 (N_15066,N_14550,N_14077);
or U15067 (N_15067,N_11221,N_11998);
xnor U15068 (N_15068,N_11950,N_14470);
nand U15069 (N_15069,N_11126,N_10977);
nor U15070 (N_15070,N_14382,N_14448);
nand U15071 (N_15071,N_12655,N_10782);
nor U15072 (N_15072,N_14008,N_14513);
or U15073 (N_15073,N_11846,N_12457);
and U15074 (N_15074,N_12623,N_11579);
nor U15075 (N_15075,N_13771,N_14696);
nor U15076 (N_15076,N_14875,N_10151);
xor U15077 (N_15077,N_12490,N_13807);
nand U15078 (N_15078,N_11475,N_10487);
nand U15079 (N_15079,N_13931,N_12738);
nand U15080 (N_15080,N_10970,N_12864);
nor U15081 (N_15081,N_13611,N_13696);
nor U15082 (N_15082,N_11218,N_13503);
nand U15083 (N_15083,N_12176,N_14303);
nor U15084 (N_15084,N_10554,N_11811);
nand U15085 (N_15085,N_13413,N_14796);
nor U15086 (N_15086,N_13964,N_12357);
nor U15087 (N_15087,N_12476,N_13318);
nand U15088 (N_15088,N_11133,N_14447);
nand U15089 (N_15089,N_11123,N_12204);
and U15090 (N_15090,N_12258,N_14278);
xnor U15091 (N_15091,N_11535,N_14418);
nand U15092 (N_15092,N_10428,N_11293);
xor U15093 (N_15093,N_12172,N_12447);
nand U15094 (N_15094,N_11864,N_10431);
nor U15095 (N_15095,N_11545,N_12139);
nor U15096 (N_15096,N_13820,N_14620);
nand U15097 (N_15097,N_10203,N_12599);
nand U15098 (N_15098,N_13162,N_10147);
and U15099 (N_15099,N_11125,N_13806);
or U15100 (N_15100,N_10657,N_14395);
and U15101 (N_15101,N_14083,N_10037);
and U15102 (N_15102,N_12800,N_10646);
or U15103 (N_15103,N_11084,N_13765);
and U15104 (N_15104,N_14544,N_14192);
nor U15105 (N_15105,N_14459,N_11631);
nor U15106 (N_15106,N_13585,N_13045);
nand U15107 (N_15107,N_14389,N_12358);
or U15108 (N_15108,N_12513,N_10619);
nor U15109 (N_15109,N_11319,N_13038);
and U15110 (N_15110,N_13824,N_12614);
nand U15111 (N_15111,N_10139,N_13419);
nand U15112 (N_15112,N_11268,N_12711);
or U15113 (N_15113,N_10754,N_14239);
nand U15114 (N_15114,N_14230,N_14237);
nand U15115 (N_15115,N_12212,N_14798);
or U15116 (N_15116,N_10158,N_13448);
nor U15117 (N_15117,N_12373,N_11727);
nor U15118 (N_15118,N_13398,N_10557);
nor U15119 (N_15119,N_14374,N_13434);
nand U15120 (N_15120,N_10853,N_10018);
or U15121 (N_15121,N_10186,N_12040);
or U15122 (N_15122,N_11434,N_10768);
and U15123 (N_15123,N_10008,N_12769);
nor U15124 (N_15124,N_10289,N_10834);
and U15125 (N_15125,N_12809,N_12379);
nor U15126 (N_15126,N_11561,N_14831);
nor U15127 (N_15127,N_11926,N_11039);
xor U15128 (N_15128,N_13062,N_11312);
and U15129 (N_15129,N_10884,N_11106);
xnor U15130 (N_15130,N_11432,N_11600);
nor U15131 (N_15131,N_12266,N_12863);
xor U15132 (N_15132,N_11670,N_13677);
nor U15133 (N_15133,N_11994,N_10163);
xor U15134 (N_15134,N_13278,N_11627);
nor U15135 (N_15135,N_13054,N_10407);
or U15136 (N_15136,N_12386,N_14288);
and U15137 (N_15137,N_14869,N_13439);
nor U15138 (N_15138,N_14203,N_10763);
and U15139 (N_15139,N_14932,N_14882);
or U15140 (N_15140,N_14337,N_11937);
and U15141 (N_15141,N_10176,N_10368);
nor U15142 (N_15142,N_11618,N_13132);
nor U15143 (N_15143,N_10796,N_12383);
and U15144 (N_15144,N_13866,N_14152);
xor U15145 (N_15145,N_10755,N_13627);
and U15146 (N_15146,N_11724,N_11699);
and U15147 (N_15147,N_14030,N_14296);
nor U15148 (N_15148,N_11054,N_14336);
nor U15149 (N_15149,N_14429,N_12362);
or U15150 (N_15150,N_13337,N_12536);
and U15151 (N_15151,N_10106,N_11323);
nor U15152 (N_15152,N_12246,N_11657);
or U15153 (N_15153,N_14481,N_11350);
nor U15154 (N_15154,N_14137,N_12325);
nor U15155 (N_15155,N_14553,N_10563);
nand U15156 (N_15156,N_14794,N_11310);
or U15157 (N_15157,N_14036,N_12264);
and U15158 (N_15158,N_14049,N_10596);
or U15159 (N_15159,N_11826,N_13378);
or U15160 (N_15160,N_13247,N_14423);
and U15161 (N_15161,N_14482,N_14075);
nor U15162 (N_15162,N_13332,N_13354);
nor U15163 (N_15163,N_13834,N_14994);
or U15164 (N_15164,N_13809,N_10086);
or U15165 (N_15165,N_11370,N_10373);
xor U15166 (N_15166,N_13213,N_13266);
or U15167 (N_15167,N_10445,N_11154);
or U15168 (N_15168,N_13542,N_11676);
nor U15169 (N_15169,N_12081,N_14308);
or U15170 (N_15170,N_14939,N_10581);
and U15171 (N_15171,N_12956,N_13007);
nor U15172 (N_15172,N_11785,N_12840);
nor U15173 (N_15173,N_13265,N_13335);
and U15174 (N_15174,N_12774,N_14750);
and U15175 (N_15175,N_10659,N_12044);
nand U15176 (N_15176,N_12468,N_14416);
and U15177 (N_15177,N_10997,N_13846);
nor U15178 (N_15178,N_11316,N_13851);
nor U15179 (N_15179,N_12662,N_13157);
or U15180 (N_15180,N_13636,N_12962);
or U15181 (N_15181,N_14785,N_14934);
nand U15182 (N_15182,N_12894,N_14726);
nor U15183 (N_15183,N_14368,N_14045);
nor U15184 (N_15184,N_10486,N_13167);
and U15185 (N_15185,N_14038,N_13424);
nor U15186 (N_15186,N_11795,N_10943);
xnor U15187 (N_15187,N_12281,N_10936);
or U15188 (N_15188,N_13343,N_11990);
nand U15189 (N_15189,N_10118,N_11562);
nor U15190 (N_15190,N_12178,N_13023);
and U15191 (N_15191,N_11853,N_11524);
or U15192 (N_15192,N_13447,N_14779);
and U15193 (N_15193,N_11099,N_12347);
or U15194 (N_15194,N_14819,N_11866);
and U15195 (N_15195,N_12461,N_14908);
nand U15196 (N_15196,N_10211,N_11018);
and U15197 (N_15197,N_13260,N_14357);
or U15198 (N_15198,N_11745,N_10980);
nand U15199 (N_15199,N_12251,N_13466);
xnor U15200 (N_15200,N_14193,N_11711);
or U15201 (N_15201,N_14034,N_10714);
nand U15202 (N_15202,N_12168,N_11495);
nor U15203 (N_15203,N_13305,N_12806);
nand U15204 (N_15204,N_12742,N_14351);
xnor U15205 (N_15205,N_12480,N_10371);
nand U15206 (N_15206,N_13856,N_13217);
nor U15207 (N_15207,N_11656,N_14834);
and U15208 (N_15208,N_13750,N_10042);
and U15209 (N_15209,N_14111,N_11428);
and U15210 (N_15210,N_12729,N_12699);
nor U15211 (N_15211,N_13746,N_11622);
nor U15212 (N_15212,N_14041,N_14621);
nor U15213 (N_15213,N_11128,N_13129);
or U15214 (N_15214,N_10511,N_12815);
xnor U15215 (N_15215,N_10722,N_14913);
nor U15216 (N_15216,N_12637,N_11245);
xor U15217 (N_15217,N_13292,N_12531);
and U15218 (N_15218,N_12186,N_13966);
nand U15219 (N_15219,N_12035,N_10221);
and U15220 (N_15220,N_11258,N_11251);
or U15221 (N_15221,N_12252,N_14283);
nor U15222 (N_15222,N_14635,N_14112);
or U15223 (N_15223,N_13853,N_10237);
and U15224 (N_15224,N_14234,N_10205);
and U15225 (N_15225,N_13529,N_10811);
nand U15226 (N_15226,N_11959,N_14841);
nand U15227 (N_15227,N_14775,N_11454);
nand U15228 (N_15228,N_13114,N_11151);
nand U15229 (N_15229,N_13982,N_10329);
xor U15230 (N_15230,N_13436,N_14977);
or U15231 (N_15231,N_10406,N_13494);
and U15232 (N_15232,N_10833,N_13168);
or U15233 (N_15233,N_10481,N_13546);
and U15234 (N_15234,N_10872,N_12590);
nand U15235 (N_15235,N_11894,N_14624);
and U15236 (N_15236,N_10700,N_10769);
nor U15237 (N_15237,N_10102,N_10799);
or U15238 (N_15238,N_11713,N_13313);
and U15239 (N_15239,N_13645,N_11592);
nor U15240 (N_15240,N_14533,N_14832);
nand U15241 (N_15241,N_13796,N_12270);
and U15242 (N_15242,N_12508,N_12153);
nor U15243 (N_15243,N_13862,N_10709);
and U15244 (N_15244,N_13884,N_10886);
xor U15245 (N_15245,N_10122,N_12914);
and U15246 (N_15246,N_14371,N_10572);
and U15247 (N_15247,N_14269,N_14091);
or U15248 (N_15248,N_14125,N_10832);
and U15249 (N_15249,N_10593,N_11334);
or U15250 (N_15250,N_12603,N_10328);
nand U15251 (N_15251,N_13226,N_10934);
or U15252 (N_15252,N_10335,N_12514);
and U15253 (N_15253,N_11022,N_13949);
and U15254 (N_15254,N_13705,N_11246);
or U15255 (N_15255,N_10501,N_12160);
xor U15256 (N_15256,N_10615,N_11920);
nand U15257 (N_15257,N_14331,N_11593);
nand U15258 (N_15258,N_13976,N_12409);
xor U15259 (N_15259,N_10874,N_12672);
nor U15260 (N_15260,N_11325,N_13601);
nand U15261 (N_15261,N_11042,N_13271);
nand U15262 (N_15262,N_11513,N_14453);
or U15263 (N_15263,N_10046,N_10418);
nor U15264 (N_15264,N_11764,N_10766);
or U15265 (N_15265,N_10978,N_12656);
or U15266 (N_15266,N_11427,N_10772);
nand U15267 (N_15267,N_13723,N_11736);
or U15268 (N_15268,N_10524,N_10167);
and U15269 (N_15269,N_10424,N_12763);
xnor U15270 (N_15270,N_11911,N_13917);
and U15271 (N_15271,N_13321,N_13633);
nand U15272 (N_15272,N_10869,N_11778);
and U15273 (N_15273,N_14174,N_13507);
or U15274 (N_15274,N_10344,N_12203);
or U15275 (N_15275,N_12229,N_11263);
nor U15276 (N_15276,N_12456,N_13566);
and U15277 (N_15277,N_11322,N_13160);
or U15278 (N_15278,N_12563,N_11922);
nand U15279 (N_15279,N_10553,N_10278);
nor U15280 (N_15280,N_11207,N_12671);
nor U15281 (N_15281,N_12568,N_10004);
or U15282 (N_15282,N_12922,N_12693);
xor U15283 (N_15283,N_10419,N_13786);
nor U15284 (N_15284,N_14712,N_14721);
nand U15285 (N_15285,N_13197,N_11633);
nor U15286 (N_15286,N_13960,N_13756);
or U15287 (N_15287,N_13681,N_14282);
nand U15288 (N_15288,N_14015,N_10116);
nand U15289 (N_15289,N_11566,N_14881);
nand U15290 (N_15290,N_12355,N_10045);
and U15291 (N_15291,N_10764,N_11146);
and U15292 (N_15292,N_13429,N_10105);
nor U15293 (N_15293,N_10504,N_14467);
xor U15294 (N_15294,N_14220,N_12963);
nor U15295 (N_15295,N_10255,N_13821);
nand U15296 (N_15296,N_10349,N_12198);
xor U15297 (N_15297,N_11835,N_11871);
and U15298 (N_15298,N_14911,N_11723);
nor U15299 (N_15299,N_12071,N_14080);
or U15300 (N_15300,N_14062,N_11443);
or U15301 (N_15301,N_14872,N_14275);
nand U15302 (N_15302,N_13901,N_12485);
or U15303 (N_15303,N_14692,N_14623);
nor U15304 (N_15304,N_14148,N_11411);
and U15305 (N_15305,N_12020,N_11138);
nand U15306 (N_15306,N_13185,N_12601);
and U15307 (N_15307,N_14260,N_11987);
nor U15308 (N_15308,N_14666,N_12961);
and U15309 (N_15309,N_14085,N_13300);
xor U15310 (N_15310,N_11342,N_12710);
or U15311 (N_15311,N_14534,N_11530);
and U15312 (N_15312,N_12643,N_14212);
nand U15313 (N_15313,N_12593,N_11445);
nand U15314 (N_15314,N_13048,N_10707);
and U15315 (N_15315,N_14529,N_11722);
xnor U15316 (N_15316,N_13516,N_13477);
nor U15317 (N_15317,N_11584,N_10254);
nand U15318 (N_15318,N_13968,N_13452);
and U15319 (N_15319,N_14329,N_14215);
or U15320 (N_15320,N_11650,N_12300);
and U15321 (N_15321,N_12886,N_12881);
nand U15322 (N_15322,N_14359,N_13534);
nand U15323 (N_15323,N_14307,N_12544);
or U15324 (N_15324,N_14110,N_10442);
nor U15325 (N_15325,N_12371,N_11611);
xor U15326 (N_15326,N_12089,N_13172);
and U15327 (N_15327,N_12045,N_13034);
and U15328 (N_15328,N_10220,N_13621);
or U15329 (N_15329,N_13433,N_13944);
nand U15330 (N_15330,N_13721,N_12124);
nand U15331 (N_15331,N_14243,N_14739);
or U15332 (N_15332,N_12992,N_13872);
and U15333 (N_15333,N_13563,N_14475);
nand U15334 (N_15334,N_12427,N_12552);
nand U15335 (N_15335,N_11698,N_11721);
nand U15336 (N_15336,N_10346,N_11825);
nand U15337 (N_15337,N_10726,N_14185);
nor U15338 (N_15338,N_14986,N_12547);
nand U15339 (N_15339,N_13275,N_13582);
xnor U15340 (N_15340,N_10571,N_11977);
or U15341 (N_15341,N_13341,N_11328);
nor U15342 (N_15342,N_11729,N_11073);
and U15343 (N_15343,N_11753,N_12833);
nor U15344 (N_15344,N_13900,N_12759);
nand U15345 (N_15345,N_12688,N_12489);
or U15346 (N_15346,N_11204,N_14172);
or U15347 (N_15347,N_12407,N_12648);
nand U15348 (N_15348,N_10223,N_13191);
nor U15349 (N_15349,N_11652,N_13060);
or U15350 (N_15350,N_11837,N_12673);
nor U15351 (N_15351,N_14647,N_12669);
nand U15352 (N_15352,N_14035,N_11969);
and U15353 (N_15353,N_12471,N_14017);
and U15354 (N_15354,N_14762,N_11161);
nand U15355 (N_15355,N_10603,N_11953);
nor U15356 (N_15356,N_11743,N_13124);
or U15357 (N_15357,N_13064,N_10236);
xor U15358 (N_15358,N_11260,N_10492);
xnor U15359 (N_15359,N_14093,N_14936);
and U15360 (N_15360,N_12694,N_13784);
nand U15361 (N_15361,N_14037,N_10066);
and U15362 (N_15362,N_14019,N_13282);
and U15363 (N_15363,N_12005,N_14432);
or U15364 (N_15364,N_10140,N_10174);
or U15365 (N_15365,N_11171,N_14235);
nand U15366 (N_15366,N_10698,N_13830);
and U15367 (N_15367,N_11700,N_13810);
nand U15368 (N_15368,N_12432,N_13925);
nand U15369 (N_15369,N_11363,N_13311);
nor U15370 (N_15370,N_10271,N_10331);
or U15371 (N_15371,N_10587,N_12746);
nor U15372 (N_15372,N_11080,N_11224);
nand U15373 (N_15373,N_11886,N_11636);
nor U15374 (N_15374,N_12319,N_11938);
and U15375 (N_15375,N_10912,N_14146);
or U15376 (N_15376,N_13152,N_11348);
and U15377 (N_15377,N_14771,N_10425);
xnor U15378 (N_15378,N_11993,N_14948);
xor U15379 (N_15379,N_11872,N_11111);
and U15380 (N_15380,N_11857,N_11282);
or U15381 (N_15381,N_14598,N_10154);
and U15382 (N_15382,N_11150,N_11256);
nor U15383 (N_15383,N_13342,N_13614);
and U15384 (N_15384,N_10882,N_13564);
nor U15385 (N_15385,N_10232,N_13244);
and U15386 (N_15386,N_10392,N_11349);
and U15387 (N_15387,N_10704,N_14128);
and U15388 (N_15388,N_11112,N_10576);
or U15389 (N_15389,N_13175,N_12380);
and U15390 (N_15390,N_14362,N_12757);
or U15391 (N_15391,N_10090,N_12521);
nor U15392 (N_15392,N_10667,N_11796);
nand U15393 (N_15393,N_12872,N_11693);
nand U15394 (N_15394,N_14570,N_13262);
and U15395 (N_15395,N_11661,N_13643);
or U15396 (N_15396,N_10910,N_10069);
or U15397 (N_15397,N_10518,N_10862);
nor U15398 (N_15398,N_11912,N_14622);
and U15399 (N_15399,N_13298,N_11897);
nand U15400 (N_15400,N_12062,N_14360);
and U15401 (N_15401,N_13122,N_14667);
nand U15402 (N_15402,N_11616,N_13431);
nor U15403 (N_15403,N_11962,N_11046);
nor U15404 (N_15404,N_11197,N_13626);
and U15405 (N_15405,N_10399,N_14201);
and U15406 (N_15406,N_14495,N_10183);
nor U15407 (N_15407,N_12243,N_12902);
nor U15408 (N_15408,N_10218,N_14033);
nor U15409 (N_15409,N_11095,N_12910);
or U15410 (N_15410,N_12762,N_14079);
nand U15411 (N_15411,N_12683,N_12685);
or U15412 (N_15412,N_10453,N_11553);
nor U15413 (N_15413,N_10573,N_10771);
nand U15414 (N_15414,N_11540,N_10676);
nor U15415 (N_15415,N_13894,N_13230);
nor U15416 (N_15416,N_10143,N_14391);
nor U15417 (N_15417,N_13923,N_11441);
nand U15418 (N_15418,N_14006,N_14643);
and U15419 (N_15419,N_14424,N_12888);
and U15420 (N_15420,N_10133,N_13314);
nand U15421 (N_15421,N_11410,N_10949);
nor U15422 (N_15422,N_11253,N_12965);
xnor U15423 (N_15423,N_11534,N_13281);
xor U15424 (N_15424,N_13423,N_13610);
and U15425 (N_15425,N_12684,N_14926);
and U15426 (N_15426,N_12487,N_14025);
nand U15427 (N_15427,N_11444,N_14340);
and U15428 (N_15428,N_13603,N_10767);
or U15429 (N_15429,N_10124,N_10716);
nand U15430 (N_15430,N_12324,N_13555);
nand U15431 (N_15431,N_12583,N_12787);
or U15432 (N_15432,N_10552,N_13100);
nor U15433 (N_15433,N_12706,N_12848);
nand U15434 (N_15434,N_12498,N_14129);
nor U15435 (N_15435,N_13324,N_10993);
nand U15436 (N_15436,N_10473,N_10495);
nand U15437 (N_15437,N_14064,N_11744);
and U15438 (N_15438,N_13941,N_14565);
nor U15439 (N_15439,N_13470,N_11810);
or U15440 (N_15440,N_13315,N_12402);
nand U15441 (N_15441,N_10224,N_14508);
or U15442 (N_15442,N_14465,N_14690);
or U15443 (N_15443,N_10068,N_11552);
nor U15444 (N_15444,N_12517,N_12618);
nand U15445 (N_15445,N_14259,N_10134);
nand U15446 (N_15446,N_11103,N_12895);
nor U15447 (N_15447,N_11004,N_13927);
nand U15448 (N_15448,N_12730,N_14594);
nor U15449 (N_15449,N_12318,N_12764);
nor U15450 (N_15450,N_10359,N_14339);
or U15451 (N_15451,N_11264,N_14270);
or U15452 (N_15452,N_10959,N_10918);
or U15453 (N_15453,N_13914,N_13693);
nor U15454 (N_15454,N_13939,N_12190);
and U15455 (N_15455,N_11588,N_10979);
or U15456 (N_15456,N_10779,N_10188);
nor U15457 (N_15457,N_10355,N_14907);
nand U15458 (N_15458,N_10826,N_14488);
or U15459 (N_15459,N_14317,N_14390);
xor U15460 (N_15460,N_11373,N_11120);
and U15461 (N_15461,N_12234,N_14719);
nand U15462 (N_15462,N_14833,N_14625);
and U15463 (N_15463,N_12296,N_14225);
nand U15464 (N_15464,N_11070,N_10966);
and U15465 (N_15465,N_10955,N_13734);
nor U15466 (N_15466,N_14676,N_10522);
nand U15467 (N_15467,N_12707,N_10762);
or U15468 (N_15468,N_11533,N_13779);
or U15469 (N_15469,N_14009,N_12056);
nor U15470 (N_15470,N_12150,N_10376);
and U15471 (N_15471,N_10230,N_12891);
nand U15472 (N_15472,N_10297,N_14258);
nor U15473 (N_15473,N_11964,N_12835);
nand U15474 (N_15474,N_10210,N_10911);
or U15475 (N_15475,N_14228,N_10701);
or U15476 (N_15476,N_14957,N_13417);
and U15477 (N_15477,N_10540,N_14186);
and U15478 (N_15478,N_10320,N_10200);
nand U15479 (N_15479,N_14250,N_13128);
or U15480 (N_15480,N_13033,N_12173);
and U15481 (N_15481,N_10257,N_12812);
and U15482 (N_15482,N_10692,N_14286);
or U15483 (N_15483,N_14683,N_11333);
and U15484 (N_15484,N_10469,N_12556);
and U15485 (N_15485,N_14793,N_11367);
nor U15486 (N_15486,N_12401,N_13004);
or U15487 (N_15487,N_11905,N_12330);
xor U15488 (N_15488,N_13743,N_10337);
nor U15489 (N_15489,N_11130,N_12540);
or U15490 (N_15490,N_14401,N_11672);
or U15491 (N_15491,N_11025,N_14864);
nor U15492 (N_15492,N_12464,N_13295);
nand U15493 (N_15493,N_13171,N_10561);
nand U15494 (N_15494,N_11467,N_14124);
and U15495 (N_15495,N_12924,N_13081);
or U15496 (N_15496,N_13016,N_13532);
xnor U15497 (N_15497,N_13604,N_14044);
and U15498 (N_15498,N_14956,N_13969);
xor U15499 (N_15499,N_11414,N_13683);
nand U15500 (N_15500,N_14849,N_12095);
xnor U15501 (N_15501,N_11907,N_14933);
or U15502 (N_15502,N_13813,N_13833);
xor U15503 (N_15503,N_10400,N_13937);
and U15504 (N_15504,N_10715,N_13403);
nand U15505 (N_15505,N_14218,N_11285);
nand U15506 (N_15506,N_11673,N_14051);
and U15507 (N_15507,N_10856,N_11274);
xor U15508 (N_15508,N_11376,N_11353);
or U15509 (N_15509,N_13783,N_11447);
nand U15510 (N_15510,N_11386,N_11807);
or U15511 (N_15511,N_10791,N_12575);
nor U15512 (N_15512,N_10354,N_11747);
or U15513 (N_15513,N_10204,N_11402);
or U15514 (N_15514,N_13459,N_10845);
nand U15515 (N_15515,N_10888,N_12183);
and U15516 (N_15516,N_12057,N_14396);
or U15517 (N_15517,N_12253,N_10577);
nor U15518 (N_15518,N_14657,N_13581);
nor U15519 (N_15519,N_12876,N_12093);
or U15520 (N_15520,N_10010,N_10616);
and U15521 (N_15521,N_11780,N_10780);
nor U15522 (N_15522,N_10879,N_14522);
nor U15523 (N_15523,N_10284,N_12128);
xor U15524 (N_15524,N_14047,N_14815);
and U15525 (N_15525,N_10758,N_10027);
xor U15526 (N_15526,N_13530,N_14605);
nand U15527 (N_15527,N_13551,N_13501);
and U15528 (N_15528,N_10530,N_10808);
or U15529 (N_15529,N_14332,N_14078);
or U15530 (N_15530,N_14310,N_12580);
and U15531 (N_15531,N_14528,N_14191);
and U15532 (N_15532,N_11862,N_12534);
or U15533 (N_15533,N_11819,N_12748);
or U15534 (N_15534,N_11684,N_13568);
nor U15535 (N_15535,N_13210,N_13950);
and U15536 (N_15536,N_13442,N_11758);
and U15537 (N_15537,N_10677,N_13410);
or U15538 (N_15538,N_12169,N_13699);
nand U15539 (N_15539,N_10155,N_11804);
nand U15540 (N_15540,N_10868,N_14411);
or U15541 (N_15541,N_10520,N_14805);
xor U15542 (N_15542,N_13112,N_14817);
nand U15543 (N_15543,N_13817,N_13299);
and U15544 (N_15544,N_11557,N_12101);
nand U15545 (N_15545,N_13445,N_12100);
and U15546 (N_15546,N_12799,N_12529);
xor U15547 (N_15547,N_12143,N_13382);
nand U15548 (N_15548,N_11664,N_13316);
nand U15549 (N_15549,N_12133,N_14344);
or U15550 (N_15550,N_12449,N_12107);
and U15551 (N_15551,N_13754,N_14407);
nor U15552 (N_15552,N_10401,N_11590);
and U15553 (N_15553,N_10272,N_13562);
nand U15554 (N_15554,N_14698,N_10731);
or U15555 (N_15555,N_10984,N_12032);
nor U15556 (N_15556,N_11321,N_13076);
nor U15557 (N_15557,N_12713,N_13874);
nand U15558 (N_15558,N_11893,N_12548);
xnor U15559 (N_15559,N_13182,N_13913);
nand U15560 (N_15560,N_10033,N_13524);
nor U15561 (N_15561,N_13912,N_12156);
nand U15562 (N_15562,N_13485,N_11273);
or U15563 (N_15563,N_13331,N_14782);
or U15564 (N_15564,N_11910,N_12930);
nor U15565 (N_15565,N_13059,N_10509);
or U15566 (N_15566,N_14468,N_10216);
nand U15567 (N_15567,N_12006,N_13646);
nor U15568 (N_15568,N_14969,N_13977);
nand U15569 (N_15569,N_13044,N_14223);
or U15570 (N_15570,N_13702,N_13548);
and U15571 (N_15571,N_11470,N_13165);
nand U15572 (N_15572,N_14410,N_10545);
nand U15573 (N_15573,N_10823,N_14338);
nand U15574 (N_15574,N_14646,N_13103);
nor U15575 (N_15575,N_14399,N_10538);
or U15576 (N_15576,N_11383,N_14850);
nor U15577 (N_15577,N_13078,N_14004);
nor U15578 (N_15578,N_13632,N_12736);
xor U15579 (N_15579,N_14539,N_12511);
and U15580 (N_15580,N_10528,N_14485);
nand U15581 (N_15581,N_10374,N_11431);
and U15582 (N_15582,N_11787,N_13737);
nand U15583 (N_15583,N_10521,N_11538);
nor U15584 (N_15584,N_10222,N_12408);
and U15585 (N_15585,N_13030,N_10642);
nor U15586 (N_15586,N_11141,N_13499);
or U15587 (N_15587,N_10123,N_10268);
nor U15588 (N_15588,N_10519,N_14415);
and U15589 (N_15589,N_13066,N_10003);
nor U15590 (N_15590,N_10468,N_12154);
nor U15591 (N_15591,N_10575,N_12374);
and U15592 (N_15592,N_10971,N_12953);
nor U15593 (N_15593,N_14134,N_11392);
nor U15594 (N_15594,N_10774,N_13506);
or U15595 (N_15595,N_13091,N_13056);
or U15596 (N_15596,N_11728,N_14991);
xor U15597 (N_15597,N_14089,N_10365);
and U15598 (N_15598,N_13446,N_11275);
or U15599 (N_15599,N_13596,N_10662);
nor U15600 (N_15600,N_12825,N_10280);
and U15601 (N_15601,N_11842,N_10381);
nor U15602 (N_15602,N_12182,N_12061);
nor U15603 (N_15603,N_13767,N_14175);
nand U15604 (N_15604,N_12528,N_11619);
or U15605 (N_15605,N_14050,N_10475);
or U15606 (N_15606,N_11032,N_12267);
nor U15607 (N_15607,N_14507,N_12798);
nand U15608 (N_15608,N_13787,N_10989);
nand U15609 (N_15609,N_11786,N_11760);
nand U15610 (N_15610,N_13306,N_14677);
and U15611 (N_15611,N_10742,N_13461);
and U15612 (N_15612,N_12375,N_12564);
or U15613 (N_15613,N_12846,N_12900);
or U15614 (N_15614,N_13854,N_12370);
and U15615 (N_15615,N_14545,N_11291);
or U15616 (N_15616,N_11045,N_14799);
or U15617 (N_15617,N_13101,N_14856);
and U15618 (N_15618,N_12999,N_12268);
and U15619 (N_15619,N_11526,N_11696);
or U15620 (N_15620,N_13684,N_12219);
and U15621 (N_15621,N_13744,N_12192);
nand U15622 (N_15622,N_10113,N_13327);
nor U15623 (N_15623,N_11477,N_11879);
and U15624 (N_15624,N_14126,N_13231);
nor U15625 (N_15625,N_11830,N_11848);
and U15626 (N_15626,N_10566,N_14807);
nor U15627 (N_15627,N_10942,N_11554);
and U15628 (N_15628,N_13531,N_12075);
nand U15629 (N_15629,N_12613,N_12467);
nand U15630 (N_15630,N_12767,N_14886);
nand U15631 (N_15631,N_11388,N_10802);
nor U15632 (N_15632,N_10635,N_10041);
or U15633 (N_15633,N_14665,N_13496);
or U15634 (N_15634,N_10382,N_11941);
and U15635 (N_15635,N_13963,N_12577);
nand U15636 (N_15636,N_12286,N_13987);
nand U15637 (N_15637,N_12441,N_12650);
xor U15638 (N_15638,N_13308,N_14524);
nand U15639 (N_15639,N_10023,N_12983);
nor U15640 (N_15640,N_11725,N_14527);
or U15641 (N_15641,N_10975,N_11719);
nor U15642 (N_15642,N_13381,N_13414);
and U15643 (N_15643,N_12157,N_13498);
nand U15644 (N_15644,N_12741,N_12678);
nor U15645 (N_15645,N_14177,N_11522);
nor U15646 (N_15646,N_13943,N_10843);
or U15647 (N_15647,N_13706,N_11613);
nand U15648 (N_15648,N_10851,N_13092);
xnor U15649 (N_15649,N_12652,N_12274);
and U15650 (N_15650,N_14742,N_10703);
or U15651 (N_15651,N_10253,N_13200);
nand U15652 (N_15652,N_12248,N_11471);
nor U15653 (N_15653,N_10474,N_12586);
nand U15654 (N_15654,N_14963,N_11916);
nand U15655 (N_15655,N_14301,N_13844);
or U15656 (N_15656,N_13204,N_11259);
and U15657 (N_15657,N_13973,N_11418);
or U15658 (N_15658,N_12078,N_14952);
nand U15659 (N_15659,N_11763,N_13367);
nand U15660 (N_15660,N_14865,N_11845);
xnor U15661 (N_15661,N_12976,N_12413);
and U15662 (N_15662,N_10015,N_14574);
and U15663 (N_15663,N_14800,N_12995);
nor U15664 (N_15664,N_12131,N_10044);
nor U15665 (N_15665,N_10672,N_12209);
nor U15666 (N_15666,N_12737,N_12340);
nor U15667 (N_15667,N_14060,N_11387);
nand U15668 (N_15668,N_14139,N_11924);
or U15669 (N_15669,N_10953,N_11029);
and U15670 (N_15670,N_13179,N_10075);
or U15671 (N_15671,N_12695,N_10505);
and U15672 (N_15672,N_13249,N_13263);
xor U15673 (N_15673,N_10836,N_14942);
and U15674 (N_15674,N_10206,N_14610);
xnor U15675 (N_15675,N_10070,N_14688);
nand U15676 (N_15676,N_13893,N_11002);
nor U15677 (N_15677,N_10290,N_12604);
or U15678 (N_15678,N_13922,N_12272);
and U15679 (N_15679,N_14503,N_12970);
and U15680 (N_15680,N_10624,N_14947);
nor U15681 (N_15681,N_11460,N_11284);
nor U15682 (N_15682,N_10161,N_10219);
nor U15683 (N_15683,N_13889,N_13954);
nor U15684 (N_15684,N_13493,N_12507);
nor U15685 (N_15685,N_13253,N_11060);
or U15686 (N_15686,N_12306,N_10778);
nor U15687 (N_15687,N_10586,N_11358);
xor U15688 (N_15688,N_13036,N_11355);
nor U15689 (N_15689,N_13233,N_13471);
or U15690 (N_15690,N_12641,N_12796);
nor U15691 (N_15691,N_14117,N_14232);
nor U15692 (N_15692,N_10270,N_12185);
and U15693 (N_15693,N_11571,N_14076);
nor U15694 (N_15694,N_11359,N_11733);
nor U15695 (N_15695,N_12037,N_12181);
nor U15696 (N_15696,N_12273,N_11306);
or U15697 (N_15697,N_10433,N_12415);
and U15698 (N_15698,N_11174,N_11170);
nand U15699 (N_15699,N_13109,N_12921);
nor U15700 (N_15700,N_12072,N_11462);
nand U15701 (N_15701,N_12745,N_12942);
xor U15702 (N_15702,N_12038,N_14001);
nor U15703 (N_15703,N_12946,N_12170);
nand U15704 (N_15704,N_11908,N_11021);
or U15705 (N_15705,N_13992,N_12708);
nand U15706 (N_15706,N_13274,N_14561);
and U15707 (N_15707,N_14949,N_12929);
xnor U15708 (N_15708,N_10588,N_12290);
or U15709 (N_15709,N_12043,N_11199);
nor U15710 (N_15710,N_11092,N_13400);
or U15711 (N_15711,N_14548,N_14923);
and U15712 (N_15712,N_14897,N_14366);
and U15713 (N_15713,N_14182,N_14104);
xor U15714 (N_15714,N_14109,N_13863);
or U15715 (N_15715,N_10721,N_13974);
and U15716 (N_15716,N_13364,N_11789);
or U15717 (N_15717,N_12931,N_11081);
nand U15718 (N_15718,N_14102,N_12444);
and U15719 (N_15719,N_14914,N_10322);
and U15720 (N_15720,N_14101,N_13219);
and U15721 (N_15721,N_11463,N_14213);
and U15722 (N_15722,N_12653,N_11071);
nor U15723 (N_15723,N_11189,N_14797);
nand U15724 (N_15724,N_10922,N_11623);
and U15725 (N_15725,N_10112,N_14378);
or U15726 (N_15726,N_12416,N_13686);
and U15727 (N_15727,N_13225,N_10562);
or U15728 (N_15728,N_11399,N_11364);
nand U15729 (N_15729,N_12682,N_14026);
and U15730 (N_15730,N_14551,N_12205);
nand U15731 (N_15731,N_10120,N_11716);
nand U15732 (N_15732,N_13541,N_13223);
nand U15733 (N_15733,N_14274,N_13328);
or U15734 (N_15734,N_10465,N_10092);
and U15735 (N_15735,N_10367,N_10181);
xor U15736 (N_15736,N_13956,N_11691);
xnor U15737 (N_15737,N_12391,N_12440);
and U15738 (N_15738,N_10100,N_14502);
or U15739 (N_15739,N_10925,N_11803);
nand U15740 (N_15740,N_12147,N_13248);
or U15741 (N_15741,N_13443,N_13803);
xnor U15742 (N_15742,N_12570,N_11237);
nand U15743 (N_15743,N_12632,N_12609);
or U15744 (N_15744,N_13680,N_11570);
and U15745 (N_15745,N_12821,N_12732);
nand U15746 (N_15746,N_11186,N_10476);
nand U15747 (N_15747,N_14010,N_10686);
nor U15748 (N_15748,N_13352,N_12889);
nor U15749 (N_15749,N_14613,N_13173);
xnor U15750 (N_15750,N_12257,N_14760);
or U15751 (N_15751,N_10546,N_10103);
and U15752 (N_15752,N_10914,N_11761);
and U15753 (N_15753,N_14320,N_14299);
nand U15754 (N_15754,N_13365,N_11741);
nand U15755 (N_15755,N_10854,N_12530);
and U15756 (N_15756,N_10281,N_12819);
nor U15757 (N_15757,N_10054,N_11109);
or U15758 (N_15758,N_14759,N_11091);
nor U15759 (N_15759,N_11946,N_14711);
or U15760 (N_15760,N_10050,N_13455);
nor U15761 (N_15761,N_11455,N_12002);
nor U15762 (N_15762,N_10598,N_12916);
xor U15763 (N_15763,N_12781,N_14729);
or U15764 (N_15764,N_10067,N_10480);
and U15765 (N_15765,N_12989,N_10450);
nor U15766 (N_15766,N_10114,N_10164);
or U15767 (N_15767,N_12994,N_13591);
and U15768 (N_15768,N_13991,N_11357);
nor U15769 (N_15769,N_11209,N_13155);
and U15770 (N_15770,N_13184,N_14653);
nor U15771 (N_15771,N_13793,N_14600);
nor U15772 (N_15772,N_14290,N_10606);
nor U15773 (N_15773,N_14494,N_11233);
and U15774 (N_15774,N_12661,N_13726);
nand U15775 (N_15775,N_10776,N_10414);
nand U15776 (N_15776,N_12724,N_12854);
nor U15777 (N_15777,N_10477,N_10683);
nand U15778 (N_15778,N_12715,N_10275);
or U15779 (N_15779,N_11678,N_14055);
xor U15780 (N_15780,N_11970,N_12103);
nor U15781 (N_15781,N_14577,N_13587);
or U15782 (N_15782,N_12602,N_11704);
and U15783 (N_15783,N_13641,N_12353);
or U15784 (N_15784,N_14571,N_12138);
and U15785 (N_15785,N_14706,N_11685);
nand U15786 (N_15786,N_12352,N_11662);
nor U15787 (N_15787,N_10962,N_14745);
or U15788 (N_15788,N_14874,N_14708);
or U15789 (N_15789,N_14648,N_13676);
or U15790 (N_15790,N_10751,N_14962);
nor U15791 (N_15791,N_13629,N_10691);
or U15792 (N_15792,N_13488,N_11324);
nor U15793 (N_15793,N_13896,N_10370);
and U15794 (N_15794,N_12197,N_13933);
nor U15795 (N_15795,N_11505,N_13383);
nor U15796 (N_15796,N_12058,N_10904);
nand U15797 (N_15797,N_11824,N_14919);
xor U15798 (N_15798,N_12086,N_12410);
or U15799 (N_15799,N_14801,N_11605);
and U15800 (N_15800,N_10544,N_12200);
nand U15801 (N_15801,N_12558,N_14951);
nand U15802 (N_15802,N_11430,N_13287);
nor U15803 (N_15803,N_10276,N_11229);
nand U15804 (N_15804,N_11595,N_13148);
nor U15805 (N_15805,N_11003,N_10411);
and U15806 (N_15806,N_13648,N_13462);
nand U15807 (N_15807,N_10787,N_12878);
xor U15808 (N_15808,N_12013,N_14954);
or U15809 (N_15809,N_12665,N_14000);
nand U15810 (N_15810,N_10121,N_14857);
xnor U15811 (N_15811,N_14005,N_14145);
or U15812 (N_15812,N_12859,N_13877);
nor U15813 (N_15813,N_10543,N_12940);
nand U15814 (N_15814,N_11979,N_13458);
and U15815 (N_15815,N_13183,N_11928);
or U15816 (N_15816,N_10141,N_13637);
nand U15817 (N_15817,N_11612,N_10287);
or U15818 (N_15818,N_13782,N_14372);
and U15819 (N_15819,N_12261,N_12225);
xor U15820 (N_15820,N_13518,N_14159);
nor U15821 (N_15821,N_14998,N_14200);
nor U15822 (N_15822,N_10215,N_14208);
nand U15823 (N_15823,N_12275,N_14756);
nor U15824 (N_15824,N_14972,N_14538);
and U15825 (N_15825,N_11774,N_11602);
nand U15826 (N_15826,N_10458,N_12398);
nor U15827 (N_15827,N_14157,N_14024);
or U15828 (N_15828,N_11874,N_13067);
or U15829 (N_15829,N_12003,N_13840);
nor U15830 (N_15830,N_13280,N_11031);
and U15831 (N_15831,N_14066,N_11531);
nand U15832 (N_15832,N_12497,N_14105);
and U15833 (N_15833,N_13740,N_13942);
nor U15834 (N_15834,N_14164,N_11630);
nor U15835 (N_15835,N_10889,N_11191);
and U15836 (N_15836,N_14725,N_10098);
nor U15837 (N_15837,N_12562,N_10748);
and U15838 (N_15838,N_13254,N_10747);
nand U15839 (N_15839,N_12850,N_11219);
xnor U15840 (N_15840,N_14498,N_11380);
or U15841 (N_15841,N_12145,N_14700);
xnor U15842 (N_15842,N_14392,N_11784);
or U15843 (N_15843,N_12220,N_13357);
or U15844 (N_15844,N_11020,N_14061);
nand U15845 (N_15845,N_11314,N_11851);
xnor U15846 (N_15846,N_13692,N_14268);
nor U15847 (N_15847,N_11738,N_13577);
nand U15848 (N_15848,N_10138,N_13940);
xnor U15849 (N_15849,N_10148,N_14630);
nand U15850 (N_15850,N_10739,N_11469);
nand U15851 (N_15851,N_12303,N_10082);
nand U15852 (N_15852,N_14753,N_10383);
nand U15853 (N_15853,N_10895,N_13144);
nand U15854 (N_15854,N_11078,N_10570);
nand U15855 (N_15855,N_14818,N_14489);
and U15856 (N_15856,N_13887,N_13098);
or U15857 (N_15857,N_10256,N_12165);
or U15858 (N_15858,N_13961,N_14901);
and U15859 (N_15859,N_11405,N_12000);
and U15860 (N_15860,N_10187,N_12551);
or U15861 (N_15861,N_11913,N_14714);
or U15862 (N_15862,N_12968,N_13593);
nor U15863 (N_15863,N_10422,N_13608);
or U15864 (N_15864,N_13412,N_13682);
nand U15865 (N_15865,N_12188,N_11261);
nor U15866 (N_15866,N_13360,N_13640);
nand U15867 (N_15867,N_11569,N_11242);
xor U15868 (N_15868,N_10641,N_12986);
or U15869 (N_15869,N_12856,N_11288);
nor U15870 (N_15870,N_14219,N_12378);
or U15871 (N_15871,N_13671,N_14787);
nor U15872 (N_15872,N_14450,N_10024);
and U15873 (N_15873,N_10578,N_14149);
nor U15874 (N_15874,N_10002,N_12755);
nand U15875 (N_15875,N_11601,N_12099);
or U15876 (N_15876,N_12144,N_11389);
or U15877 (N_15877,N_12175,N_12797);
nand U15878 (N_15878,N_12634,N_12780);
or U15879 (N_15879,N_14546,N_11558);
nand U15880 (N_15880,N_10246,N_13599);
nor U15881 (N_15881,N_11821,N_13768);
nor U15882 (N_15882,N_10296,N_14876);
nand U15883 (N_15883,N_12024,N_12102);
nor U15884 (N_15884,N_10434,N_13766);
nor U15885 (N_15885,N_13201,N_14555);
nor U15886 (N_15886,N_14645,N_14661);
and U15887 (N_15887,N_12055,N_10944);
nor U15888 (N_15888,N_10960,N_13955);
xnor U15889 (N_15889,N_13207,N_11692);
nand U15890 (N_15890,N_10435,N_11436);
and U15891 (N_15891,N_10012,N_13831);
nand U15892 (N_15892,N_11423,N_14743);
nor U15893 (N_15893,N_14007,N_12596);
and U15894 (N_15894,N_10301,N_13617);
nand U15895 (N_15895,N_11508,N_11024);
and U15896 (N_15896,N_11110,N_13178);
and U15897 (N_15897,N_14830,N_11658);
and U15898 (N_15898,N_14058,N_10678);
or U15899 (N_15899,N_13240,N_10583);
nand U15900 (N_15900,N_13380,N_14795);
or U15901 (N_15901,N_13811,N_14361);
or U15902 (N_15902,N_13967,N_14904);
nand U15903 (N_15903,N_13797,N_13957);
nand U15904 (N_15904,N_11037,N_14373);
xor U15905 (N_15905,N_10348,N_14224);
nand U15906 (N_15906,N_14788,N_14915);
nand U15907 (N_15907,N_12893,N_10077);
nor U15908 (N_15908,N_13325,N_13574);
or U15909 (N_15909,N_11902,N_14567);
nor U15910 (N_15910,N_10109,N_10760);
nor U15911 (N_15911,N_11882,N_10074);
and U15912 (N_15912,N_12892,N_12113);
nand U15913 (N_15913,N_11492,N_12046);
and U15914 (N_15914,N_13134,N_14890);
xnor U15915 (N_15915,N_10170,N_11488);
or U15916 (N_15916,N_10169,N_12884);
nand U15917 (N_15917,N_12813,N_10968);
nor U15918 (N_15918,N_10656,N_14178);
nand U15919 (N_15919,N_14297,N_12794);
and U15920 (N_15920,N_14569,N_14096);
nand U15921 (N_15921,N_13652,N_10896);
xor U15922 (N_15922,N_11643,N_13822);
nor U15923 (N_15923,N_10099,N_13427);
or U15924 (N_15924,N_13732,N_12070);
and U15925 (N_15925,N_12028,N_11849);
nand U15926 (N_15926,N_11577,N_11490);
or U15927 (N_15927,N_10119,N_14214);
nor U15928 (N_15928,N_12187,N_10841);
xnor U15929 (N_15929,N_14910,N_13505);
nor U15930 (N_15930,N_10352,N_11012);
nor U15931 (N_15931,N_10166,N_12022);
nand U15932 (N_15932,N_13972,N_12853);
nand U15933 (N_15933,N_13291,N_14414);
and U15934 (N_15934,N_14027,N_11818);
nor U15935 (N_15935,N_14241,N_13550);
or U15936 (N_15936,N_14652,N_13035);
nor U15937 (N_15937,N_11779,N_10743);
nand U15938 (N_15938,N_14040,N_10423);
nand U15939 (N_15939,N_13024,N_13769);
xnor U15940 (N_15940,N_13946,N_11708);
nor U15941 (N_15941,N_14918,N_13011);
nor U15942 (N_15942,N_13138,N_10753);
or U15943 (N_15943,N_11269,N_10330);
or U15944 (N_15944,N_13284,N_14902);
nor U15945 (N_15945,N_14161,N_12422);
nor U15946 (N_15946,N_12404,N_11093);
nand U15947 (N_15947,N_10732,N_14153);
nor U15948 (N_15948,N_10192,N_13347);
xor U15949 (N_15949,N_14086,N_12051);
nor U15950 (N_15950,N_13620,N_13290);
or U15951 (N_15951,N_14967,N_14221);
nand U15952 (N_15952,N_11991,N_14931);
and U15953 (N_15953,N_10837,N_13077);
or U15954 (N_15954,N_14930,N_11576);
and U15955 (N_15955,N_11175,N_14599);
or U15956 (N_15956,N_10650,N_14961);
and U15957 (N_15957,N_14678,N_10795);
or U15958 (N_15958,N_10420,N_13948);
nor U15959 (N_15959,N_14573,N_14597);
nand U15960 (N_15960,N_12826,N_12063);
nand U15961 (N_15961,N_11885,N_10614);
or U15962 (N_15962,N_13146,N_10775);
and U15963 (N_15963,N_12206,N_12923);
or U15964 (N_15964,N_11244,N_12073);
nor U15965 (N_15965,N_10865,N_12472);
xnor U15966 (N_15966,N_13040,N_10891);
and U15967 (N_15967,N_14393,N_12428);
or U15968 (N_15968,N_14379,N_13312);
nor U15969 (N_15969,N_14701,N_10021);
nand U15970 (N_15970,N_12376,N_12333);
xnor U15971 (N_15971,N_11210,N_14568);
or U15972 (N_15972,N_12244,N_11292);
nor U15973 (N_15973,N_12222,N_13021);
nand U15974 (N_15974,N_13984,N_13259);
xnor U15975 (N_15975,N_10020,N_13580);
nor U15976 (N_15976,N_11485,N_14852);
and U15977 (N_15977,N_11396,N_10718);
or U15978 (N_15978,N_14322,N_10441);
or U15979 (N_15979,N_14069,N_14641);
nor U15980 (N_15980,N_14738,N_12933);
nand U15981 (N_15981,N_13962,N_14755);
xor U15982 (N_15982,N_12179,N_12526);
and U15983 (N_15983,N_11982,N_10523);
xnor U15984 (N_15984,N_14084,N_14560);
xnor U15985 (N_15985,N_10403,N_13052);
or U15986 (N_15986,N_13037,N_10017);
nor U15987 (N_15987,N_11527,N_10484);
xor U15988 (N_15988,N_14216,N_12919);
nor U15989 (N_15989,N_12280,N_10638);
nand U15990 (N_15990,N_13776,N_14272);
nor U15991 (N_15991,N_13425,N_14113);
and U15992 (N_15992,N_10610,N_12442);
or U15993 (N_15993,N_10179,N_12782);
or U15994 (N_15994,N_11823,N_11139);
or U15995 (N_15995,N_12313,N_10001);
and U15996 (N_15996,N_14877,N_12322);
or U15997 (N_15997,N_14018,N_10019);
nand U15998 (N_15998,N_10720,N_13921);
or U15999 (N_15999,N_11925,N_10909);
xnor U16000 (N_16000,N_14443,N_14032);
and U16001 (N_16001,N_11214,N_11575);
or U16002 (N_16002,N_11435,N_11064);
xnor U16003 (N_16003,N_13029,N_11548);
xor U16004 (N_16004,N_10706,N_10752);
nor U16005 (N_16005,N_11313,N_11227);
nor U16006 (N_16006,N_13986,N_10674);
or U16007 (N_16007,N_11473,N_12849);
nor U16008 (N_16008,N_13691,N_12474);
and U16009 (N_16009,N_13835,N_12451);
nor U16010 (N_16010,N_10369,N_11005);
xnor U16011 (N_16011,N_10160,N_10663);
xnor U16012 (N_16012,N_12475,N_12725);
nor U16013 (N_16013,N_13363,N_10648);
xnor U16014 (N_16014,N_14905,N_13539);
or U16015 (N_16015,N_11401,N_14675);
or U16016 (N_16016,N_13514,N_10006);
xor U16017 (N_16017,N_11539,N_14380);
or U16018 (N_16018,N_11281,N_12218);
or U16019 (N_16019,N_10671,N_13801);
xnor U16020 (N_16020,N_10548,N_11914);
nand U16021 (N_16021,N_12837,N_13276);
xor U16022 (N_16022,N_10264,N_14629);
nor U16023 (N_16023,N_13490,N_11317);
or U16024 (N_16024,N_10858,N_13657);
and U16025 (N_16025,N_14757,N_12098);
nand U16026 (N_16026,N_11489,N_12576);
nand U16027 (N_16027,N_14277,N_14167);
and U16028 (N_16028,N_14885,N_11628);
nor U16029 (N_16029,N_14642,N_13886);
or U16030 (N_16030,N_10235,N_13465);
or U16031 (N_16031,N_13196,N_13252);
or U16032 (N_16032,N_10195,N_12036);
nor U16033 (N_16033,N_12566,N_12532);
xnor U16034 (N_16034,N_12896,N_12166);
or U16035 (N_16035,N_14868,N_10389);
nand U16036 (N_16036,N_12194,N_11816);
and U16037 (N_16037,N_14435,N_10675);
or U16038 (N_16038,N_14291,N_10807);
or U16039 (N_16039,N_10729,N_12161);
nor U16040 (N_16040,N_14484,N_10507);
nand U16041 (N_16041,N_12831,N_13336);
or U16042 (N_16042,N_13739,N_13839);
or U16043 (N_16043,N_11063,N_10059);
or U16044 (N_16044,N_11184,N_10866);
nor U16045 (N_16045,N_14761,N_12982);
nor U16046 (N_16046,N_11320,N_11407);
nor U16047 (N_16047,N_12704,N_12744);
nand U16048 (N_16048,N_13142,N_12344);
or U16049 (N_16049,N_10814,N_13788);
or U16050 (N_16050,N_13523,N_11720);
or U16051 (N_16051,N_13826,N_10696);
or U16052 (N_16052,N_14858,N_14444);
or U16053 (N_16053,N_13478,N_12025);
and U16054 (N_16054,N_14871,N_10240);
nand U16055 (N_16055,N_13222,N_14853);
nand U16056 (N_16056,N_11781,N_12309);
nor U16057 (N_16057,N_13307,N_12783);
nand U16058 (N_16058,N_14824,N_10880);
xnor U16059 (N_16059,N_12317,N_12950);
or U16060 (N_16060,N_13805,N_11000);
nor U16061 (N_16061,N_10629,N_13838);
and U16062 (N_16062,N_10258,N_11503);
nand U16063 (N_16063,N_14896,N_11252);
nand U16064 (N_16064,N_11583,N_12984);
nand U16065 (N_16065,N_13107,N_12106);
or U16066 (N_16066,N_13212,N_11768);
xor U16067 (N_16067,N_10948,N_13123);
nand U16068 (N_16068,N_14406,N_14511);
or U16069 (N_16069,N_13025,N_11290);
and U16070 (N_16070,N_11368,N_11878);
or U16071 (N_16071,N_13905,N_11655);
and U16072 (N_16072,N_11059,N_12610);
or U16073 (N_16073,N_10390,N_11299);
nor U16074 (N_16074,N_13393,N_13444);
and U16075 (N_16075,N_14898,N_14873);
and U16076 (N_16076,N_13559,N_13359);
xnor U16077 (N_16077,N_13689,N_14487);
xnor U16078 (N_16078,N_11884,N_13221);
xor U16079 (N_16079,N_10637,N_10983);
nand U16080 (N_16080,N_10781,N_10062);
or U16081 (N_16081,N_14592,N_10084);
xor U16082 (N_16082,N_11155,N_14845);
nand U16083 (N_16083,N_12751,N_12247);
nor U16084 (N_16084,N_14964,N_10622);
or U16085 (N_16085,N_11801,N_14764);
or U16086 (N_16086,N_12749,N_11216);
or U16087 (N_16087,N_14011,N_14273);
nor U16088 (N_16088,N_11930,N_12712);
nor U16089 (N_16089,N_11249,N_12687);
nand U16090 (N_16090,N_14514,N_13117);
nand U16091 (N_16091,N_12210,N_14632);
nor U16092 (N_16092,N_10695,N_10579);
and U16093 (N_16093,N_11466,N_11235);
or U16094 (N_16094,N_14252,N_13061);
nand U16095 (N_16095,N_12041,N_14644);
and U16096 (N_16096,N_12311,N_13068);
nand U16097 (N_16097,N_11265,N_12329);
nor U16098 (N_16098,N_12944,N_10185);
nor U16099 (N_16099,N_13089,N_12481);
nand U16100 (N_16100,N_11890,N_13920);
xnor U16101 (N_16101,N_10180,N_12486);
xnor U16102 (N_16102,N_10850,N_12777);
nand U16103 (N_16103,N_14417,N_14521);
or U16104 (N_16104,N_11944,N_11814);
or U16105 (N_16105,N_13647,N_13374);
and U16106 (N_16106,N_12512,N_14016);
and U16107 (N_16107,N_14087,N_11074);
and U16108 (N_16108,N_10459,N_11574);
and U16109 (N_16109,N_14183,N_14803);
nand U16110 (N_16110,N_13339,N_14162);
nor U16111 (N_16111,N_13735,N_14168);
xnor U16112 (N_16112,N_13170,N_14928);
nand U16113 (N_16113,N_14305,N_14970);
and U16114 (N_16114,N_14449,N_14433);
xor U16115 (N_16115,N_14585,N_11337);
nor U16116 (N_16116,N_13661,N_13356);
nand U16117 (N_16117,N_12869,N_12943);
nor U16118 (N_16118,N_13454,N_11891);
nor U16119 (N_16119,N_14263,N_11955);
and U16120 (N_16120,N_11104,N_10438);
and U16121 (N_16121,N_13003,N_10661);
or U16122 (N_16122,N_13286,N_12882);
nor U16123 (N_16123,N_13340,N_11769);
nand U16124 (N_16124,N_13131,N_14115);
nor U16125 (N_16125,N_13527,N_14618);
and U16126 (N_16126,N_10260,N_10245);
and U16127 (N_16127,N_11113,N_14098);
xor U16128 (N_16128,N_11496,N_10226);
nor U16129 (N_16129,N_10613,N_14323);
or U16130 (N_16130,N_11163,N_11817);
nand U16131 (N_16131,N_13483,N_12589);
or U16132 (N_16132,N_14184,N_10199);
nand U16133 (N_16133,N_10311,N_13362);
or U16134 (N_16134,N_11550,N_13174);
nand U16135 (N_16135,N_12717,N_12162);
or U16136 (N_16136,N_10871,N_10655);
and U16137 (N_16137,N_12852,N_12786);
nor U16138 (N_16138,N_12448,N_12174);
or U16139 (N_16139,N_13935,N_12277);
nor U16140 (N_16140,N_10567,N_14912);
xor U16141 (N_16141,N_11178,N_12328);
and U16142 (N_16142,N_12125,N_14251);
nor U16143 (N_16143,N_10490,N_11514);
or U16144 (N_16144,N_14617,N_10372);
and U16145 (N_16145,N_14043,N_11984);
nor U16146 (N_16146,N_10556,N_12011);
xnor U16147 (N_16147,N_14627,N_12450);
nor U16148 (N_16148,N_11206,N_12510);
and U16149 (N_16149,N_12594,N_11296);
nor U16150 (N_16150,N_11438,N_13557);
and U16151 (N_16151,N_11481,N_12913);
and U16152 (N_16152,N_10049,N_13869);
or U16153 (N_16153,N_10198,N_10599);
xnor U16154 (N_16154,N_12969,N_12585);
nand U16155 (N_16155,N_12802,N_10687);
or U16156 (N_16156,N_10804,N_13031);
and U16157 (N_16157,N_10972,N_10773);
nand U16158 (N_16158,N_11660,N_13521);
nand U16159 (N_16159,N_11748,N_12158);
or U16160 (N_16160,N_14068,N_12626);
nand U16161 (N_16161,N_12624,N_10309);
nor U16162 (N_16162,N_12954,N_10360);
or U16163 (N_16163,N_10825,N_10535);
nor U16164 (N_16164,N_14811,N_14123);
and U16165 (N_16165,N_13093,N_12348);
or U16166 (N_16166,N_12754,N_13001);
nand U16167 (N_16167,N_13104,N_11549);
nor U16168 (N_16168,N_13659,N_13837);
xor U16169 (N_16169,N_12136,N_12433);
xor U16170 (N_16170,N_11075,N_10690);
and U16171 (N_16171,N_11542,N_10633);
and U16172 (N_16172,N_10048,N_10994);
and U16173 (N_16173,N_13584,N_10584);
nor U16174 (N_16174,N_11996,N_10489);
or U16175 (N_16175,N_13453,N_12233);
and U16176 (N_16176,N_11520,N_10043);
nor U16177 (N_16177,N_13069,N_14891);
nor U16178 (N_16178,N_11271,N_12042);
or U16179 (N_16179,N_12533,N_10417);
or U16180 (N_16180,N_14823,N_13251);
nor U16181 (N_16181,N_10565,N_14279);
nand U16182 (N_16182,N_10515,N_10085);
nor U16183 (N_16183,N_11083,N_10876);
or U16184 (N_16184,N_12034,N_12395);
nand U16185 (N_16185,N_12299,N_13792);
or U16186 (N_16186,N_10908,N_11805);
nor U16187 (N_16187,N_14071,N_11203);
or U16188 (N_16188,N_11859,N_13985);
or U16189 (N_16189,N_10712,N_14691);
and U16190 (N_16190,N_11497,N_14960);
nand U16191 (N_16191,N_12048,N_14002);
nand U16192 (N_16192,N_12958,N_11205);
or U16193 (N_16193,N_10711,N_12980);
and U16194 (N_16194,N_12155,N_12691);
nand U16195 (N_16195,N_12284,N_12360);
nand U16196 (N_16196,N_14013,N_10078);
and U16197 (N_16197,N_12616,N_13202);
and U16198 (N_16198,N_11833,N_11608);
and U16199 (N_16199,N_12332,N_10430);
nor U16200 (N_16200,N_12615,N_13072);
and U16201 (N_16201,N_14781,N_14684);
and U16202 (N_16202,N_14767,N_13892);
nand U16203 (N_16203,N_12697,N_12535);
or U16204 (N_16204,N_11114,N_10087);
xor U16205 (N_16205,N_14469,N_10736);
nor U16206 (N_16206,N_10785,N_12207);
and U16207 (N_16207,N_11587,N_14820);
nor U16208 (N_16208,N_10626,N_11829);
and U16209 (N_16209,N_14616,N_10136);
nor U16210 (N_16210,N_12001,N_14206);
or U16211 (N_16211,N_11677,N_13186);
nor U16212 (N_16212,N_12617,N_10517);
or U16213 (N_16213,N_10455,N_12838);
and U16214 (N_16214,N_11393,N_10597);
and U16215 (N_16215,N_10104,N_13602);
nor U16216 (N_16216,N_12973,N_14638);
xnor U16217 (N_16217,N_13097,N_11201);
and U16218 (N_16218,N_14595,N_12285);
or U16219 (N_16219,N_10427,N_11202);
xnor U16220 (N_16220,N_11049,N_14846);
nor U16221 (N_16221,N_10028,N_11965);
or U16222 (N_16222,N_13317,N_10353);
nand U16223 (N_16223,N_10713,N_13389);
nand U16224 (N_16224,N_11255,N_13799);
xnor U16225 (N_16225,N_13304,N_10965);
nand U16226 (N_16226,N_10534,N_10660);
and U16227 (N_16227,N_14477,N_12808);
or U16228 (N_16228,N_13755,N_12004);
or U16229 (N_16229,N_11706,N_11762);
or U16230 (N_16230,N_12584,N_11105);
and U16231 (N_16231,N_12334,N_14584);
and U16232 (N_16232,N_11194,N_10047);
or U16233 (N_16233,N_11169,N_12775);
xor U16234 (N_16234,N_13710,N_11369);
or U16235 (N_16235,N_11157,N_11225);
or U16236 (N_16236,N_12345,N_14309);
nand U16237 (N_16237,N_12670,N_10498);
or U16238 (N_16238,N_12855,N_13147);
nor U16239 (N_16239,N_14097,N_12463);
nor U16240 (N_16240,N_12770,N_11502);
or U16241 (N_16241,N_13338,N_12722);
or U16242 (N_16242,N_14445,N_11351);
xnor U16243 (N_16243,N_10746,N_11966);
nand U16244 (N_16244,N_11160,N_14709);
and U16245 (N_16245,N_12629,N_10875);
xnor U16246 (N_16246,N_11961,N_12555);
nand U16247 (N_16247,N_14980,N_13473);
xnor U16248 (N_16248,N_10094,N_13589);
and U16249 (N_16249,N_10899,N_11147);
nor U16250 (N_16250,N_10356,N_12239);
xnor U16251 (N_16251,N_11262,N_11958);
xnor U16252 (N_16252,N_13492,N_11122);
nand U16253 (N_16253,N_13050,N_11464);
nor U16254 (N_16254,N_12901,N_12703);
or U16255 (N_16255,N_12949,N_12298);
nand U16256 (N_16256,N_10820,N_10801);
xnor U16257 (N_16257,N_10654,N_14879);
and U16258 (N_16258,N_13032,N_14776);
nand U16259 (N_16259,N_12117,N_11865);
or U16260 (N_16260,N_14518,N_13409);
xnor U16261 (N_16261,N_14840,N_10483);
nor U16262 (N_16262,N_13216,N_10303);
or U16263 (N_16263,N_11390,N_12436);
nand U16264 (N_16264,N_14562,N_10717);
and U16265 (N_16265,N_11896,N_13055);
and U16266 (N_16266,N_12446,N_13607);
or U16267 (N_16267,N_14261,N_14039);
or U16268 (N_16268,N_13772,N_10921);
nor U16269 (N_16269,N_12016,N_12226);
and U16270 (N_16270,N_13088,N_13116);
nor U16271 (N_16271,N_11921,N_10855);
and U16272 (N_16272,N_10719,N_14749);
and U16273 (N_16273,N_14633,N_10189);
and U16274 (N_16274,N_13469,N_14993);
nor U16275 (N_16275,N_13708,N_14386);
nand U16276 (N_16276,N_11563,N_10680);
nor U16277 (N_16277,N_13947,N_12494);
and U16278 (N_16278,N_11840,N_11379);
and U16279 (N_16279,N_12979,N_11211);
nand U16280 (N_16280,N_14431,N_14133);
nand U16281 (N_16281,N_10022,N_10810);
nand U16282 (N_16282,N_11521,N_13685);
nor U16283 (N_16283,N_14367,N_11935);
and U16284 (N_16284,N_13804,N_12276);
nor U16285 (N_16285,N_14227,N_12885);
or U16286 (N_16286,N_13763,N_13544);
xor U16287 (N_16287,N_12680,N_14249);
xor U16288 (N_16288,N_10702,N_14483);
nand U16289 (N_16289,N_11934,N_10541);
or U16290 (N_16290,N_13760,N_10601);
and U16291 (N_16291,N_14012,N_12265);
and U16292 (N_16292,N_10986,N_10595);
nand U16293 (N_16293,N_11371,N_12918);
and U16294 (N_16294,N_10551,N_10292);
or U16295 (N_16295,N_14654,N_11304);
or U16296 (N_16296,N_14384,N_14313);
nor U16297 (N_16297,N_11972,N_12939);
xor U16298 (N_16298,N_11585,N_14586);
nand U16299 (N_16299,N_12971,N_10594);
or U16300 (N_16300,N_12473,N_10125);
xor U16301 (N_16301,N_12294,N_12231);
nor U16302 (N_16302,N_14839,N_13176);
xnor U16303 (N_16303,N_10890,N_14181);
nor U16304 (N_16304,N_12359,N_10318);
nor U16305 (N_16305,N_10549,N_10324);
nand U16306 (N_16306,N_13569,N_10783);
nor U16307 (N_16307,N_11222,N_10282);
and U16308 (N_16308,N_10788,N_14821);
nand U16309 (N_16309,N_10857,N_13415);
or U16310 (N_16310,N_11860,N_11767);
nor U16311 (N_16311,N_12690,N_10229);
nor U16312 (N_16312,N_10673,N_12110);
nand U16313 (N_16313,N_11638,N_10816);
or U16314 (N_16314,N_10265,N_13020);
nand U16315 (N_16315,N_11732,N_13227);
xnor U16316 (N_16316,N_12496,N_11038);
and U16317 (N_16317,N_13828,N_10060);
nand U16318 (N_16318,N_10126,N_13242);
or U16319 (N_16319,N_10725,N_10034);
nor U16320 (N_16320,N_12996,N_14142);
xnor U16321 (N_16321,N_11472,N_11854);
nand U16322 (N_16322,N_12723,N_13426);
nor U16323 (N_16323,N_13511,N_12470);
xor U16324 (N_16324,N_12114,N_14413);
nor U16325 (N_16325,N_10397,N_13238);
nor U16326 (N_16326,N_10496,N_13592);
and U16327 (N_16327,N_14319,N_13656);
and U16328 (N_16328,N_12438,N_12642);
and U16329 (N_16329,N_13345,N_13858);
or U16330 (N_16330,N_10923,N_12459);
nor U16331 (N_16331,N_12674,N_12377);
or U16332 (N_16332,N_12163,N_12587);
nand U16333 (N_16333,N_11968,N_10494);
and U16334 (N_16334,N_11456,N_11459);
nand U16335 (N_16335,N_12017,N_11543);
or U16336 (N_16336,N_12753,N_10749);
nand U16337 (N_16337,N_12660,N_14813);
or U16338 (N_16338,N_13159,N_14702);
xor U16339 (N_16339,N_14778,N_10512);
nand U16340 (N_16340,N_12297,N_13576);
or U16341 (N_16341,N_14244,N_10699);
or U16342 (N_16342,N_13651,N_14063);
and U16343 (N_16343,N_11270,N_14981);
and U16344 (N_16344,N_10878,N_12747);
nand U16345 (N_16345,N_11448,N_11757);
nand U16346 (N_16346,N_11519,N_13781);
and U16347 (N_16347,N_11043,N_11062);
and U16348 (N_16348,N_14114,N_12709);
or U16349 (N_16349,N_11695,N_11420);
or U16350 (N_16350,N_12142,N_12820);
nor U16351 (N_16351,N_12911,N_12054);
or U16352 (N_16352,N_14705,N_14523);
or U16353 (N_16353,N_12304,N_11347);
nor U16354 (N_16354,N_14848,N_12651);
nand U16355 (N_16355,N_10283,N_10502);
nor U16356 (N_16356,N_14658,N_13819);
nor U16357 (N_16357,N_13890,N_14505);
or U16358 (N_16358,N_14222,N_10926);
nand U16359 (N_16359,N_14321,N_11957);
nand U16360 (N_16360,N_12771,N_10307);
nor U16361 (N_16361,N_10756,N_14072);
and U16362 (N_16362,N_10590,N_12720);
nand U16363 (N_16363,N_10930,N_11152);
nor U16364 (N_16364,N_11040,N_12335);
and U16365 (N_16365,N_10096,N_10321);
or U16366 (N_16366,N_13401,N_14304);
nor U16367 (N_16367,N_14975,N_14383);
or U16368 (N_16368,N_14280,N_13420);
and U16369 (N_16369,N_12906,N_11117);
xor U16370 (N_16370,N_10177,N_12361);
xnor U16371 (N_16371,N_12477,N_11058);
nor U16372 (N_16372,N_14144,N_13158);
xnor U16373 (N_16373,N_12033,N_11875);
or U16374 (N_16374,N_13404,N_11635);
or U16375 (N_16375,N_10471,N_14878);
and U16376 (N_16376,N_14751,N_10416);
or U16377 (N_16377,N_12466,N_12912);
or U16378 (N_16378,N_11667,N_12341);
nand U16379 (N_16379,N_13808,N_12947);
and U16380 (N_16380,N_14941,N_12242);
and U16381 (N_16381,N_10797,N_12199);
nand U16382 (N_16382,N_12096,N_10658);
or U16383 (N_16383,N_13909,N_14298);
nand U16384 (N_16384,N_11649,N_11429);
xnor U16385 (N_16385,N_11408,N_13387);
xnor U16386 (N_16386,N_14559,N_13268);
xnor U16387 (N_16387,N_11568,N_14722);
nand U16388 (N_16388,N_10460,N_13126);
nor U16389 (N_16389,N_12790,N_11315);
nand U16390 (N_16390,N_12326,N_14204);
and U16391 (N_16391,N_12692,N_12418);
or U16392 (N_16392,N_13264,N_11793);
and U16393 (N_16393,N_11506,N_10150);
and U16394 (N_16394,N_11701,N_10171);
nor U16395 (N_16395,N_13269,N_11135);
or U16396 (N_16396,N_11028,N_13881);
or U16397 (N_16397,N_10451,N_13619);
or U16398 (N_16398,N_14179,N_13934);
nand U16399 (N_16399,N_13888,N_10437);
xor U16400 (N_16400,N_14579,N_14580);
nand U16401 (N_16401,N_14660,N_10089);
nand U16402 (N_16402,N_13829,N_14537);
or U16403 (N_16403,N_12735,N_11877);
nor U16404 (N_16404,N_10285,N_10585);
nand U16405 (N_16405,N_14059,N_11050);
nand U16406 (N_16406,N_13902,N_13392);
nor U16407 (N_16407,N_10175,N_13695);
or U16408 (N_16408,N_12727,N_12728);
or U16409 (N_16409,N_12630,N_10761);
or U16410 (N_16410,N_11036,N_13753);
or U16411 (N_16411,N_14659,N_13533);
and U16412 (N_16412,N_14937,N_11510);
or U16413 (N_16413,N_14385,N_10093);
and U16414 (N_16414,N_10688,N_13919);
nor U16415 (N_16415,N_12559,N_10981);
nor U16416 (N_16416,N_13785,N_12573);
xor U16417 (N_16417,N_14333,N_10159);
or U16418 (N_16418,N_14615,N_11799);
and U16419 (N_16419,N_12612,N_10592);
nand U16420 (N_16420,N_12292,N_10649);
and U16421 (N_16421,N_11669,N_12429);
nor U16422 (N_16422,N_11703,N_14003);
or U16423 (N_16423,N_12622,N_14663);
and U16424 (N_16424,N_12606,N_10409);
or U16425 (N_16425,N_14828,N_11231);
xnor U16426 (N_16426,N_13111,N_12832);
nor U16427 (N_16427,N_10144,N_11378);
and U16428 (N_16428,N_12959,N_13351);
or U16429 (N_16429,N_13084,N_13519);
or U16430 (N_16430,N_12030,N_10961);
xor U16431 (N_16431,N_14207,N_11047);
and U16432 (N_16432,N_14394,N_10313);
or U16433 (N_16433,N_12538,N_11052);
and U16434 (N_16434,N_12793,N_12112);
and U16435 (N_16435,N_10063,N_11889);
nor U16436 (N_16436,N_11560,N_14356);
and U16437 (N_16437,N_14116,N_13898);
nor U16438 (N_16438,N_12116,N_13718);
and U16439 (N_16439,N_13394,N_10366);
and U16440 (N_16440,N_11599,N_14127);
xnor U16441 (N_16441,N_12647,N_13791);
and U16442 (N_16442,N_12844,N_14451);
and U16443 (N_16443,N_11832,N_13558);
and U16444 (N_16444,N_13115,N_14893);
or U16445 (N_16445,N_10443,N_13463);
or U16446 (N_16446,N_13738,N_11360);
nor U16447 (N_16447,N_12184,N_12491);
or U16448 (N_16448,N_12331,N_14458);
and U16449 (N_16449,N_12282,N_12077);
nand U16450 (N_16450,N_10503,N_12082);
nand U16451 (N_16451,N_12293,N_13228);
and U16452 (N_16452,N_13218,N_12115);
nand U16453 (N_16453,N_13662,N_11134);
or U16454 (N_16454,N_11834,N_10279);
and U16455 (N_16455,N_12423,N_10393);
or U16456 (N_16456,N_10784,N_12998);
nor U16457 (N_16457,N_13715,N_12988);
nand U16458 (N_16458,N_10727,N_14141);
or U16459 (N_16459,N_11847,N_10466);
nor U16460 (N_16460,N_14053,N_13320);
nor U16461 (N_16461,N_11188,N_11179);
and U16462 (N_16462,N_12053,N_11085);
or U16463 (N_16463,N_13598,N_13041);
nand U16464 (N_16464,N_10259,N_12667);
nand U16465 (N_16465,N_14325,N_13508);
nand U16466 (N_16466,N_12104,N_10470);
nor U16467 (N_16467,N_12217,N_11705);
nor U16468 (N_16468,N_12600,N_11220);
and U16469 (N_16469,N_14456,N_14067);
nand U16470 (N_16470,N_10681,N_10973);
nand U16471 (N_16471,N_11565,N_11581);
nand U16472 (N_16472,N_13717,N_10669);
and U16473 (N_16473,N_12132,N_13832);
or U16474 (N_16474,N_10117,N_11409);
or U16475 (N_16475,N_10830,N_12019);
and U16476 (N_16476,N_10903,N_12936);
nor U16477 (N_16477,N_12865,N_13849);
and U16478 (N_16478,N_12779,N_10190);
nand U16479 (N_16479,N_12654,N_11346);
xor U16480 (N_16480,N_10867,N_11257);
and U16481 (N_16481,N_14945,N_11989);
nor U16482 (N_16482,N_11149,N_12120);
xnor U16483 (N_16483,N_14530,N_10609);
or U16484 (N_16484,N_11683,N_14350);
or U16485 (N_16485,N_14163,N_13166);
or U16486 (N_16486,N_10274,N_10627);
nor U16487 (N_16487,N_12645,N_12126);
and U16488 (N_16488,N_12686,N_10057);
or U16489 (N_16489,N_11808,N_13996);
nand U16490 (N_16490,N_14486,N_11501);
and U16491 (N_16491,N_10813,N_14151);
or U16492 (N_16492,N_13396,N_10202);
nor U16493 (N_16493,N_13018,N_12778);
or U16494 (N_16494,N_13150,N_13437);
or U16495 (N_16495,N_10333,N_11338);
or U16496 (N_16496,N_14953,N_10439);
nand U16497 (N_16497,N_12830,N_11906);
xnor U16498 (N_16498,N_12920,N_12412);
and U16499 (N_16499,N_11394,N_13449);
and U16500 (N_16500,N_14165,N_14438);
or U16501 (N_16501,N_12941,N_12839);
xor U16502 (N_16502,N_14780,N_10840);
nand U16503 (N_16503,N_12012,N_14670);
and U16504 (N_16504,N_13724,N_13475);
and U16505 (N_16505,N_10061,N_13998);
and U16506 (N_16506,N_12452,N_10847);
nand U16507 (N_16507,N_14982,N_11710);
nand U16508 (N_16508,N_12052,N_14436);
and U16509 (N_16509,N_12437,N_13981);
and U16510 (N_16510,N_13842,N_13669);
and U16511 (N_16511,N_12705,N_10824);
or U16512 (N_16512,N_12365,N_11181);
and U16513 (N_16513,N_10030,N_13929);
or U16514 (N_16514,N_14735,N_12631);
or U16515 (N_16515,N_11735,N_11680);
and U16516 (N_16516,N_10817,N_11856);
or U16517 (N_16517,N_13102,N_12084);
nor U16518 (N_16518,N_14649,N_14827);
xor U16519 (N_16519,N_14662,N_10846);
xnor U16520 (N_16520,N_12860,N_10913);
nand U16521 (N_16521,N_11176,N_14838);
and U16522 (N_16522,N_12469,N_14314);
or U16523 (N_16523,N_11400,N_10724);
and U16524 (N_16524,N_14065,N_11468);
or U16525 (N_16525,N_13644,N_13047);
and U16526 (N_16526,N_13430,N_14197);
nor U16527 (N_16527,N_10738,N_14842);
nor U16528 (N_16528,N_13549,N_14388);
nor U16529 (N_16529,N_14466,N_12488);
or U16530 (N_16530,N_11715,N_14720);
nand U16531 (N_16531,N_11289,N_10315);
nor U16532 (N_16532,N_10759,N_13719);
or U16533 (N_16533,N_14188,N_11356);
or U16534 (N_16534,N_11686,N_12829);
or U16535 (N_16535,N_12064,N_10071);
and U16536 (N_16536,N_13301,N_11165);
or U16537 (N_16537,N_11494,N_11551);
and U16538 (N_16538,N_10009,N_13609);
or U16539 (N_16539,N_10651,N_13594);
xor U16540 (N_16540,N_12721,N_14903);
nor U16541 (N_16541,N_14255,N_13258);
nand U16542 (N_16542,N_11901,N_11751);
and U16543 (N_16543,N_14996,N_11644);
or U16544 (N_16544,N_14899,N_10472);
nand U16545 (N_16545,N_14596,N_10000);
or U16546 (N_16546,N_14324,N_10940);
nand U16547 (N_16547,N_13707,N_12887);
nand U16548 (N_16548,N_11066,N_11088);
nor U16549 (N_16549,N_13106,N_11248);
nor U16550 (N_16550,N_11674,N_10231);
and U16551 (N_16551,N_13323,N_10679);
or U16552 (N_16552,N_14345,N_13105);
nor U16553 (N_16553,N_12240,N_11931);
or U16554 (N_16554,N_13395,N_14347);
nor U16555 (N_16555,N_10266,N_12504);
or U16556 (N_16556,N_11688,N_12816);
or U16557 (N_16557,N_14806,N_11734);
and U16558 (N_16558,N_13504,N_14816);
and U16559 (N_16559,N_11836,N_13575);
and U16560 (N_16560,N_12392,N_12565);
and U16561 (N_16561,N_13229,N_13095);
or U16562 (N_16562,N_11499,N_12842);
xnor U16563 (N_16563,N_11007,N_10319);
nand U16564 (N_16564,N_10640,N_13198);
xnor U16565 (N_16565,N_14812,N_10812);
nand U16566 (N_16566,N_14682,N_11718);
or U16567 (N_16567,N_14349,N_10375);
and U16568 (N_16568,N_10870,N_11107);
nor U16569 (N_16569,N_12069,N_10893);
nand U16570 (N_16570,N_11681,N_14256);
nor U16571 (N_16571,N_10305,N_13897);
nor U16572 (N_16572,N_11416,N_12700);
nand U16573 (N_16573,N_14976,N_10744);
nor U16574 (N_16574,N_11486,N_11948);
and U16575 (N_16575,N_13074,N_10464);
nor U16576 (N_16576,N_14809,N_13741);
or U16577 (N_16577,N_12382,N_14131);
or U16578 (N_16578,N_13203,N_14090);
xnor U16579 (N_16579,N_11626,N_12349);
xnor U16580 (N_16580,N_10386,N_13606);
nand U16581 (N_16581,N_14971,N_14334);
and U16582 (N_16582,N_14777,N_11142);
or U16583 (N_16583,N_11512,N_10634);
or U16584 (N_16584,N_14589,N_11391);
or U16585 (N_16585,N_12788,N_14107);
nor U16586 (N_16586,N_12195,N_13205);
nand U16587 (N_16587,N_13468,N_10357);
and U16588 (N_16588,N_13774,N_14656);
nand U16589 (N_16589,N_14515,N_14474);
nor U16590 (N_16590,N_13867,N_14602);
nor U16591 (N_16591,N_10560,N_12074);
nor U16592 (N_16592,N_13553,N_10182);
and U16593 (N_16593,N_10864,N_11936);
and U16594 (N_16594,N_10327,N_12458);
and U16595 (N_16595,N_14187,N_13703);
and U16596 (N_16596,N_10065,N_10317);
nand U16597 (N_16597,N_11654,N_14387);
nand U16598 (N_16598,N_10786,N_13751);
nor U16599 (N_16599,N_14607,N_11336);
and U16600 (N_16600,N_14916,N_13373);
and U16601 (N_16601,N_14532,N_12237);
or U16602 (N_16602,N_13232,N_13255);
and U16603 (N_16603,N_11572,N_10905);
nand U16604 (N_16604,N_11952,N_11213);
nand U16605 (N_16605,N_10447,N_12411);
or U16606 (N_16606,N_12581,N_12828);
xnor U16607 (N_16607,N_11422,N_10920);
and U16608 (N_16608,N_11424,N_13545);
nor U16609 (N_16609,N_12394,N_10623);
and U16610 (N_16610,N_11812,N_13536);
nor U16611 (N_16611,N_13958,N_11498);
or U16612 (N_16612,N_12560,N_12021);
and U16613 (N_16613,N_11666,N_13775);
nand U16614 (N_16614,N_12008,N_13163);
nand U16615 (N_16615,N_12620,N_14264);
or U16616 (N_16616,N_12905,N_10415);
nor U16617 (N_16617,N_13177,N_11532);
and U16618 (N_16618,N_10351,N_13297);
nand U16619 (N_16619,N_11480,N_14925);
nand U16620 (N_16620,N_14499,N_13722);
or U16621 (N_16621,N_14588,N_12509);
nor U16622 (N_16622,N_11341,N_14108);
xor U16623 (N_16623,N_11690,N_14122);
or U16624 (N_16624,N_12338,N_13547);
and U16625 (N_16625,N_12628,N_13279);
nand U16626 (N_16626,N_11413,N_12818);
nand U16627 (N_16627,N_13876,N_10456);
xor U16628 (N_16628,N_13537,N_14922);
or U16629 (N_16629,N_13371,N_13628);
xnor U16630 (N_16630,N_12636,N_11694);
and U16631 (N_16631,N_11973,N_10011);
nor U16632 (N_16632,N_12550,N_14293);
or U16633 (N_16633,N_13285,N_11287);
xnor U16634 (N_16634,N_12571,N_11663);
or U16635 (N_16635,N_10252,N_13823);
or U16636 (N_16636,N_11559,N_12426);
nor U16637 (N_16637,N_13528,N_11440);
nor U16638 (N_16638,N_13903,N_10178);
or U16639 (N_16639,N_12123,N_14989);
or U16640 (N_16640,N_12180,N_12351);
and U16641 (N_16641,N_13572,N_14884);
nand U16642 (N_16642,N_11986,N_14446);
or U16643 (N_16643,N_12431,N_10621);
or U16644 (N_16644,N_14985,N_12343);
and U16645 (N_16645,N_13727,N_12140);
nand U16646 (N_16646,N_12625,N_10402);
nand U16647 (N_16647,N_10745,N_12023);
and U16648 (N_16648,N_13411,N_14376);
nor U16649 (N_16649,N_13309,N_10806);
or U16650 (N_16650,N_11838,N_11286);
nand U16651 (N_16651,N_12388,N_11094);
and U16652 (N_16652,N_14992,N_12675);
nand U16653 (N_16653,N_11034,N_12271);
nand U16654 (N_16654,N_10239,N_12454);
nor U16655 (N_16655,N_10340,N_12518);
xnor U16656 (N_16656,N_13733,N_13590);
or U16657 (N_16657,N_11951,N_12760);
nor U16658 (N_16658,N_10542,N_11679);
and U16659 (N_16659,N_10838,N_12937);
or U16660 (N_16660,N_11949,N_11915);
nor U16661 (N_16661,N_10625,N_10902);
nand U16662 (N_16662,N_10362,N_12733);
and U16663 (N_16663,N_13464,N_12479);
and U16664 (N_16664,N_12834,N_10286);
nand U16665 (N_16665,N_10842,N_12406);
nor U16666 (N_16666,N_10582,N_11182);
and U16667 (N_16667,N_11250,N_11148);
or U16668 (N_16668,N_12546,N_11307);
xor U16669 (N_16669,N_12091,N_10800);
and U16670 (N_16670,N_12105,N_10604);
nand U16671 (N_16671,N_14855,N_10479);
nor U16672 (N_16672,N_13798,N_14674);
nor U16673 (N_16673,N_10039,N_13481);
nand U16674 (N_16674,N_13156,N_12214);
nor U16675 (N_16675,N_14810,N_11403);
nor U16676 (N_16676,N_12758,N_11707);
nor U16677 (N_16677,N_12792,N_13510);
nand U16678 (N_16678,N_11898,N_10446);
and U16679 (N_16679,N_11839,N_13502);
nor U16680 (N_16680,N_12907,N_11041);
nor U16681 (N_16681,N_11983,N_10408);
or U16682 (N_16682,N_12542,N_12801);
xor U16683 (N_16683,N_11415,N_13745);
nor U16684 (N_16684,N_12364,N_13027);
xnor U16685 (N_16685,N_14281,N_13918);
or U16686 (N_16686,N_12097,N_12639);
or U16687 (N_16687,N_12342,N_11086);
nand U16688 (N_16688,N_11417,N_10129);
or U16689 (N_16689,N_10939,N_10915);
xor U16690 (N_16690,N_12369,N_10267);
xnor U16691 (N_16691,N_10516,N_13195);
and U16692 (N_16692,N_12283,N_11239);
and U16693 (N_16693,N_10251,N_10277);
or U16694 (N_16694,N_13860,N_12525);
nor U16695 (N_16695,N_10338,N_10938);
nor U16696 (N_16696,N_12726,N_13137);
or U16697 (N_16697,N_10835,N_14727);
nor U16698 (N_16698,N_10935,N_12484);
xor U16699 (N_16699,N_11124,N_14176);
nand U16700 (N_16700,N_11870,N_11311);
nand U16701 (N_16701,N_11023,N_11006);
nor U16702 (N_16702,N_10379,N_13391);
or U16703 (N_16703,N_13495,N_11001);
nand U16704 (N_16704,N_12847,N_11437);
and U16705 (N_16705,N_12701,N_10448);
nand U16706 (N_16706,N_13141,N_12810);
and U16707 (N_16707,N_14427,N_11515);
nor U16708 (N_16708,N_14073,N_14022);
nor U16709 (N_16709,N_13816,N_14457);
or U16710 (N_16710,N_12714,N_14262);
and U16711 (N_16711,N_11923,N_12047);
nand U16712 (N_16712,N_13836,N_13043);
nand U16713 (N_16713,N_10873,N_14023);
and U16714 (N_16714,N_14276,N_11740);
and U16715 (N_16715,N_14713,N_12756);
nor U16716 (N_16716,N_11918,N_11484);
xnor U16717 (N_16717,N_11507,N_10887);
nand U16718 (N_16718,N_12776,N_10985);
and U16719 (N_16719,N_12851,N_14836);
or U16720 (N_16720,N_10031,N_10697);
nand U16721 (N_16721,N_13467,N_11140);
nor U16722 (N_16722,N_12430,N_14020);
and U16723 (N_16723,N_14479,N_13484);
nor U16724 (N_16724,N_14870,N_14944);
and U16725 (N_16725,N_12768,N_12236);
nand U16726 (N_16726,N_11119,N_12858);
nor U16727 (N_16727,N_14369,N_12553);
xor U16728 (N_16728,N_10095,N_13605);
xor U16729 (N_16729,N_14581,N_10664);
and U16730 (N_16730,N_12635,N_14791);
and U16731 (N_16731,N_14217,N_13878);
nor U16732 (N_16732,N_13193,N_13698);
nand U16733 (N_16733,N_11712,N_11048);
nand U16734 (N_16734,N_11056,N_10945);
nor U16735 (N_16735,N_10991,N_13353);
nor U16736 (N_16736,N_11226,N_14572);
nand U16737 (N_16737,N_13432,N_12991);
nor U16738 (N_16738,N_12316,N_10974);
or U16739 (N_16739,N_13234,N_13911);
or U16740 (N_16740,N_12862,N_12805);
and U16741 (N_16741,N_10072,N_14564);
and U16742 (N_16742,N_12301,N_13579);
or U16743 (N_16743,N_14103,N_14099);
nor U16744 (N_16744,N_11880,N_11971);
nand U16745 (N_16745,N_11820,N_13907);
nand U16746 (N_16746,N_13938,N_13802);
nand U16747 (N_16747,N_12087,N_10630);
nor U16748 (N_16748,N_13658,N_13192);
nand U16749 (N_16749,N_11339,N_14512);
and U16750 (N_16750,N_14405,N_14979);
nor U16751 (N_16751,N_14520,N_14847);
xnor U16752 (N_16752,N_10454,N_10013);
nor U16753 (N_16753,N_13953,N_13749);
nor U16754 (N_16754,N_12215,N_13895);
and U16755 (N_16755,N_13418,N_10079);
nand U16756 (N_16756,N_14476,N_12460);
xor U16757 (N_16757,N_10152,N_12567);
nand U16758 (N_16758,N_12523,N_11129);
or U16759 (N_16759,N_13673,N_14634);
and U16760 (N_16760,N_13538,N_10798);
or U16761 (N_16761,N_11621,N_11665);
nor U16762 (N_16762,N_13730,N_13113);
or U16763 (N_16763,N_13143,N_12520);
and U16764 (N_16764,N_11195,N_12904);
nand U16765 (N_16765,N_11143,N_11247);
and U16766 (N_16766,N_13979,N_10861);
nor U16767 (N_16767,N_11992,N_10111);
and U16768 (N_16768,N_13668,N_11573);
xor U16769 (N_16769,N_14766,N_12827);
or U16770 (N_16770,N_13075,N_13057);
nand U16771 (N_16771,N_12679,N_11381);
nor U16772 (N_16772,N_10342,N_10493);
or U16773 (N_16773,N_14439,N_13597);
nand U16774 (N_16774,N_11755,N_11243);
and U16775 (N_16775,N_11750,N_10014);
nor U16776 (N_16776,N_14442,N_10385);
or U16777 (N_16777,N_13928,N_13361);
nor U16778 (N_16778,N_13688,N_14680);
or U16779 (N_16779,N_13046,N_12663);
nand U16780 (N_16780,N_10631,N_11236);
nand U16781 (N_16781,N_14209,N_10213);
and U16782 (N_16782,N_12861,N_12060);
and U16783 (N_16783,N_12148,N_13366);
and U16784 (N_16784,N_11158,N_14628);
nor U16785 (N_16785,N_10197,N_13472);
and U16786 (N_16786,N_13679,N_14768);
nor U16787 (N_16787,N_14978,N_12083);
nand U16788 (N_16788,N_11011,N_14195);
and U16789 (N_16789,N_12734,N_10611);
nor U16790 (N_16790,N_10108,N_12841);
or U16791 (N_16791,N_14180,N_12903);
nor U16792 (N_16792,N_11132,N_13672);
nor U16793 (N_16793,N_14478,N_14460);
nand U16794 (N_16794,N_13416,N_13778);
and U16795 (N_16795,N_10710,N_12094);
and U16796 (N_16796,N_12278,N_10173);
xnor U16797 (N_16797,N_12681,N_14461);
or U16798 (N_16798,N_10907,N_12354);
nor U16799 (N_16799,N_12250,N_14143);
or U16800 (N_16800,N_12807,N_13017);
nor U16801 (N_16801,N_11634,N_13667);
nand U16802 (N_16802,N_14626,N_12873);
nand U16803 (N_16803,N_10395,N_14887);
or U16804 (N_16804,N_13543,N_14888);
and U16805 (N_16805,N_10803,N_11975);
nand U16806 (N_16806,N_14772,N_11079);
nand U16807 (N_16807,N_13079,N_10463);
and U16808 (N_16808,N_10608,N_12619);
nor U16809 (N_16809,N_11254,N_11689);
nor U16810 (N_16810,N_12291,N_11876);
and U16811 (N_16811,N_13397,N_13615);
nor U16812 (N_16812,N_10332,N_11887);
nand U16813 (N_16813,N_10685,N_11279);
or U16814 (N_16814,N_12879,N_12932);
xnor U16815 (N_16815,N_11121,N_11297);
and U16816 (N_16816,N_11791,N_11167);
and U16817 (N_16817,N_14651,N_10076);
nor U16818 (N_16818,N_11303,N_11340);
and U16819 (N_16819,N_12987,N_11895);
nand U16820 (N_16820,N_13790,N_14999);
or U16821 (N_16821,N_13310,N_11335);
and U16822 (N_16822,N_10569,N_13709);
nand U16823 (N_16823,N_13847,N_12595);
and U16824 (N_16824,N_10885,N_10056);
nor U16825 (N_16825,N_14549,N_11776);
nand U16826 (N_16826,N_11089,N_10917);
nor U16827 (N_16827,N_12478,N_13789);
nand U16828 (N_16828,N_13322,N_14671);
or U16829 (N_16829,N_10526,N_14880);
and U16830 (N_16830,N_13690,N_12597);
nor U16831 (N_16831,N_14328,N_12644);
nand U16832 (N_16832,N_11230,N_10491);
and U16833 (N_16833,N_13026,N_13635);
or U16834 (N_16834,N_12483,N_14844);
nor U16835 (N_16835,N_14057,N_11775);
nor U16836 (N_16836,N_12718,N_12372);
and U16837 (N_16837,N_12164,N_10249);
and U16838 (N_16838,N_10302,N_12638);
and U16839 (N_16839,N_11277,N_10026);
and U16840 (N_16840,N_11101,N_10574);
and U16841 (N_16841,N_11985,N_12719);
xor U16842 (N_16842,N_13235,N_12957);
xor U16843 (N_16843,N_14959,N_12092);
nor U16844 (N_16844,N_11881,N_12898);
nand U16845 (N_16845,N_11374,N_12381);
xor U16846 (N_16846,N_10877,N_14516);
nand U16847 (N_16847,N_10294,N_13870);
nor U16848 (N_16848,N_10988,N_14464);
nand U16849 (N_16849,N_13859,N_13267);
nor U16850 (N_16850,N_13236,N_11087);
or U16851 (N_16851,N_14758,N_10793);
and U16852 (N_16852,N_11589,N_14563);
or U16853 (N_16853,N_12890,N_10750);
nand U16854 (N_16854,N_12981,N_11625);
or U16855 (N_16855,N_14655,N_14741);
nor U16856 (N_16856,N_10436,N_11127);
nor U16857 (N_16857,N_12249,N_10967);
nor U16858 (N_16858,N_11726,N_13390);
and U16859 (N_16859,N_12193,N_13302);
or U16860 (N_16860,N_14921,N_13065);
nor U16861 (N_16861,N_12588,N_12611);
or U16862 (N_16862,N_13650,N_13015);
and U16863 (N_16863,N_11717,N_13082);
nor U16864 (N_16864,N_14199,N_11425);
xor U16865 (N_16865,N_13479,N_14557);
nand U16866 (N_16866,N_14381,N_13561);
xor U16867 (N_16867,N_13108,N_14497);
and U16868 (N_16868,N_14422,N_14302);
or U16869 (N_16869,N_14789,N_11610);
nor U16870 (N_16870,N_13169,N_11956);
and U16871 (N_16871,N_12814,N_11478);
xnor U16872 (N_16872,N_13180,N_11067);
and U16873 (N_16873,N_10269,N_11653);
and U16874 (N_16874,N_14746,N_14397);
nand U16875 (N_16875,N_12320,N_13670);
or U16876 (N_16876,N_10733,N_12159);
or U16877 (N_16877,N_11746,N_11177);
nand U16878 (N_16878,N_12871,N_13554);
nand U16879 (N_16879,N_11858,N_13777);
nor U16880 (N_16880,N_14636,N_10536);
nor U16881 (N_16881,N_14121,N_14246);
nor U16882 (N_16882,N_10449,N_10035);
or U16883 (N_16883,N_13063,N_14718);
nor U16884 (N_16884,N_13526,N_11813);
and U16885 (N_16885,N_10225,N_14335);
nor U16886 (N_16886,N_14704,N_14590);
and U16887 (N_16887,N_14346,N_10982);
nor U16888 (N_16888,N_13012,N_12387);
nand U16889 (N_16889,N_10191,N_13206);
nor U16890 (N_16890,N_14906,N_12766);
and U16891 (N_16891,N_11802,N_14686);
nand U16892 (N_16892,N_13277,N_10146);
or U16893 (N_16893,N_14404,N_12899);
or U16894 (N_16894,N_12129,N_12135);
nor U16895 (N_16895,N_13818,N_14517);
nor U16896 (N_16896,N_10207,N_11809);
or U16897 (N_16897,N_12505,N_13486);
nand U16898 (N_16898,N_11044,N_12403);
nand U16899 (N_16899,N_11241,N_11668);
or U16900 (N_16900,N_13971,N_13515);
and U16901 (N_16901,N_14238,N_12118);
and U16902 (N_16902,N_12545,N_10467);
and U16903 (N_16903,N_13513,N_14547);
xor U16904 (N_16904,N_11792,N_14752);
nand U16905 (N_16905,N_14326,N_11917);
nand U16906 (N_16906,N_11797,N_11614);
and U16907 (N_16907,N_12578,N_11929);
and U16908 (N_16908,N_12262,N_11730);
or U16909 (N_16909,N_13994,N_12137);
and U16910 (N_16910,N_13460,N_14997);
nand U16911 (N_16911,N_11988,N_12453);
xnor U16912 (N_16912,N_11395,N_14496);
nor U16913 (N_16913,N_13552,N_12191);
and U16914 (N_16914,N_12649,N_10580);
nor U16915 (N_16915,N_13595,N_10091);
or U16916 (N_16916,N_13714,N_11375);
nand U16917 (N_16917,N_14531,N_10741);
and U16918 (N_16918,N_13080,N_13978);
and U16919 (N_16919,N_10947,N_14859);
and U16920 (N_16920,N_10730,N_13049);
or U16921 (N_16921,N_14611,N_10898);
xnor U16922 (N_16922,N_14318,N_13348);
nor U16923 (N_16923,N_14229,N_11739);
nor U16924 (N_16924,N_11055,N_10819);
nand U16925 (N_16925,N_11742,N_13214);
and U16926 (N_16926,N_11754,N_12065);
nand U16927 (N_16927,N_10083,N_10273);
nor U16928 (N_16928,N_11597,N_10387);
nand U16929 (N_16929,N_12646,N_10233);
nor U16930 (N_16930,N_10682,N_13711);
or U16931 (N_16931,N_11397,N_14242);
xnor U16932 (N_16932,N_11945,N_10398);
nand U16933 (N_16933,N_10956,N_13916);
nor U16934 (N_16934,N_13435,N_12260);
nor U16935 (N_16935,N_14851,N_13660);
nand U16936 (N_16936,N_10291,N_13154);
and U16937 (N_16937,N_14315,N_13457);
nor U16938 (N_16938,N_11053,N_10848);
nor U16939 (N_16939,N_13571,N_14608);
nand U16940 (N_16940,N_13762,N_13855);
or U16941 (N_16941,N_13489,N_10196);
or U16942 (N_16942,N_10723,N_10088);
and U16943 (N_16943,N_10016,N_12230);
nand U16944 (N_16944,N_14082,N_14412);
or U16945 (N_16945,N_12167,N_11841);
xor U16946 (N_16946,N_13239,N_14783);
xnor U16947 (N_16947,N_11398,N_13583);
nand U16948 (N_16948,N_13071,N_11180);
nand U16949 (N_16949,N_10217,N_10954);
or U16950 (N_16950,N_13355,N_14867);
or U16951 (N_16951,N_13164,N_13864);
nand U16952 (N_16952,N_13476,N_14029);
nand U16953 (N_16953,N_11976,N_11193);
xor U16954 (N_16954,N_14327,N_13256);
xor U16955 (N_16955,N_10995,N_11168);
or U16956 (N_16956,N_12399,N_14240);
or U16957 (N_16957,N_12845,N_14452);
nor U16958 (N_16958,N_10777,N_12739);
or U16959 (N_16959,N_12689,N_10308);
or U16960 (N_16960,N_10208,N_13250);
nand U16961 (N_16961,N_12978,N_10919);
and U16962 (N_16962,N_10999,N_10537);
xnor U16963 (N_16963,N_11035,N_12515);
or U16964 (N_16964,N_12111,N_12633);
and U16965 (N_16965,N_10510,N_14074);
or U16966 (N_16966,N_13211,N_13450);
and U16967 (N_16967,N_10792,N_13906);
nor U16968 (N_16968,N_14170,N_13570);
nand U16969 (N_16969,N_13385,N_13402);
or U16970 (N_16970,N_14710,N_11153);
or U16971 (N_16971,N_14226,N_12659);
xor U16972 (N_16972,N_13736,N_14965);
and U16973 (N_16973,N_14155,N_13729);
nor U16974 (N_16974,N_13926,N_13491);
nor U16975 (N_16975,N_10963,N_11234);
or U16976 (N_16976,N_14826,N_14506);
nand U16977 (N_16977,N_12791,N_14862);
nor U16978 (N_16978,N_13634,N_12314);
and U16979 (N_16979,N_11372,N_11332);
and U16980 (N_16980,N_14409,N_14860);
or U16981 (N_16981,N_14774,N_14554);
or U16982 (N_16982,N_12390,N_13241);
or U16983 (N_16983,N_11318,N_10478);
or U16984 (N_16984,N_13631,N_11223);
nand U16985 (N_16985,N_10852,N_11137);
nand U16986 (N_16986,N_14526,N_14542);
nand U16987 (N_16987,N_14894,N_12569);
xnor U16988 (N_16988,N_12811,N_14472);
nand U16989 (N_16989,N_12598,N_13408);
or U16990 (N_16990,N_12424,N_14070);
nor U16991 (N_16991,N_14837,N_10300);
nand U16992 (N_16992,N_11187,N_11995);
nor U16993 (N_16993,N_14614,N_13270);
nand U16994 (N_16994,N_10380,N_13930);
nor U16995 (N_16995,N_13110,N_12350);
or U16996 (N_16996,N_10378,N_14150);
and U16997 (N_16997,N_13970,N_13540);
or U16998 (N_16998,N_13814,N_12664);
xnor U16999 (N_16999,N_13388,N_11212);
nand U17000 (N_17000,N_10821,N_13421);
or U17001 (N_17001,N_13675,N_11909);
or U17002 (N_17002,N_11974,N_13995);
and U17003 (N_17003,N_10128,N_10462);
and U17004 (N_17004,N_10497,N_13406);
or U17005 (N_17005,N_14054,N_10941);
nand U17006 (N_17006,N_10306,N_14311);
xnor U17007 (N_17007,N_12141,N_10193);
nor U17008 (N_17008,N_12221,N_14375);
nor U17009 (N_17009,N_10946,N_14728);
nor U17010 (N_17010,N_11385,N_14031);
and U17011 (N_17011,N_10347,N_13087);
nor U17012 (N_17012,N_10527,N_10860);
nor U17013 (N_17013,N_12605,N_11645);
or U17014 (N_17014,N_13720,N_11482);
nand U17015 (N_17015,N_11594,N_13199);
xor U17016 (N_17016,N_10525,N_12419);
nand U17017 (N_17017,N_11033,N_11331);
and U17018 (N_17018,N_14740,N_11639);
nor U17019 (N_17019,N_11065,N_13010);
nor U17020 (N_17020,N_10929,N_12287);
and U17021 (N_17021,N_11697,N_10933);
nand U17022 (N_17022,N_14619,N_13480);
nand U17023 (N_17023,N_10558,N_10172);
nor U17024 (N_17024,N_10931,N_10928);
or U17025 (N_17025,N_13891,N_14265);
nor U17026 (N_17026,N_10336,N_14462);
nor U17027 (N_17027,N_10384,N_12366);
and U17028 (N_17028,N_14088,N_13133);
nand U17029 (N_17029,N_10097,N_10135);
or U17030 (N_17030,N_14927,N_12405);
and U17031 (N_17031,N_14430,N_11102);
nand U17032 (N_17032,N_12773,N_11546);
and U17033 (N_17033,N_14566,N_10794);
nand U17034 (N_17034,N_10555,N_14420);
nor U17035 (N_17035,N_14733,N_13344);
nand U17036 (N_17036,N_11190,N_10906);
nand U17037 (N_17037,N_12068,N_14535);
nor U17038 (N_17038,N_11603,N_13296);
or U17039 (N_17039,N_13618,N_12874);
xnor U17040 (N_17040,N_10293,N_14909);
nor U17041 (N_17041,N_12527,N_13070);
nand U17042 (N_17042,N_12666,N_13405);
nand U17043 (N_17043,N_12731,N_10396);
and U17044 (N_17044,N_14247,N_10863);
and U17045 (N_17045,N_10410,N_12336);
or U17046 (N_17046,N_13330,N_11861);
or U17047 (N_17047,N_10343,N_12238);
and U17048 (N_17048,N_11098,N_10670);
or U17049 (N_17049,N_13578,N_10358);
or U17050 (N_17050,N_10325,N_10298);
nor U17051 (N_17051,N_14501,N_14330);
nand U17052 (N_17052,N_13019,N_11173);
nand U17053 (N_17053,N_13085,N_12591);
and U17054 (N_17054,N_10334,N_10345);
or U17055 (N_17055,N_14973,N_10115);
nand U17056 (N_17056,N_10894,N_11097);
and U17057 (N_17057,N_12315,N_14306);
or U17058 (N_17058,N_12130,N_12420);
and U17059 (N_17059,N_11709,N_11516);
nor U17060 (N_17060,N_14968,N_12524);
nor U17061 (N_17061,N_12189,N_10957);
nor U17062 (N_17062,N_14773,N_14292);
and U17063 (N_17063,N_12817,N_13625);
nor U17064 (N_17064,N_13613,N_13747);
nor U17065 (N_17065,N_13573,N_14822);
nand U17066 (N_17066,N_13451,N_14575);
and U17067 (N_17067,N_10647,N_14754);
xor U17068 (N_17068,N_14940,N_11145);
nand U17069 (N_17069,N_11166,N_13399);
and U17070 (N_17070,N_12305,N_13090);
and U17071 (N_17071,N_12417,N_11382);
and U17072 (N_17072,N_10058,N_13600);
xnor U17073 (N_17073,N_14748,N_11997);
nand U17074 (N_17074,N_12935,N_10992);
and U17075 (N_17075,N_13642,N_11017);
nor U17076 (N_17076,N_13002,N_12960);
or U17077 (N_17077,N_11759,N_10243);
nand U17078 (N_17078,N_11637,N_10620);
xor U17079 (N_17079,N_14156,N_12455);
nor U17080 (N_17080,N_12621,N_11345);
and U17081 (N_17081,N_10262,N_11671);
nor U17082 (N_17082,N_13384,N_12543);
nor U17083 (N_17083,N_11354,N_13153);
or U17084 (N_17084,N_13377,N_13376);
and U17085 (N_17085,N_12439,N_12263);
xor U17086 (N_17086,N_14342,N_14769);
and U17087 (N_17087,N_13073,N_13827);
nand U17088 (N_17088,N_14693,N_13509);
nand U17089 (N_17089,N_13622,N_12608);
xor U17090 (N_17090,N_13752,N_12938);
nor U17091 (N_17091,N_12974,N_12824);
or U17092 (N_17092,N_13780,N_12822);
nor U17093 (N_17093,N_11108,N_11476);
nor U17094 (N_17094,N_14863,N_11919);
or U17095 (N_17095,N_12592,N_10666);
nor U17096 (N_17096,N_10617,N_12337);
nor U17097 (N_17097,N_13742,N_10612);
xor U17098 (N_17098,N_13407,N_13841);
nor U17099 (N_17099,N_10341,N_13713);
and U17100 (N_17100,N_14895,N_10131);
or U17101 (N_17101,N_12435,N_12288);
nand U17102 (N_17102,N_14202,N_13812);
and U17103 (N_17103,N_14408,N_12928);
nor U17104 (N_17104,N_13868,N_14639);
or U17105 (N_17105,N_10550,N_14398);
nand U17106 (N_17106,N_13440,N_10591);
and U17107 (N_17107,N_10080,N_12857);
nand U17108 (N_17108,N_12368,N_13623);
nand U17109 (N_17109,N_12109,N_11770);
xnor U17110 (N_17110,N_14341,N_12772);
nand U17111 (N_17111,N_11453,N_12495);
nor U17112 (N_17112,N_11217,N_10127);
nand U17113 (N_17113,N_14606,N_13630);
nor U17114 (N_17114,N_11183,N_11208);
and U17115 (N_17115,N_10559,N_13588);
nor U17116 (N_17116,N_10299,N_13149);
or U17117 (N_17117,N_13999,N_14300);
nor U17118 (N_17118,N_13639,N_13135);
nand U17119 (N_17119,N_10452,N_12010);
and U17120 (N_17120,N_10568,N_12211);
nand U17121 (N_17121,N_13624,N_10149);
and U17122 (N_17122,N_10737,N_12676);
nand U17123 (N_17123,N_14744,N_14492);
xnor U17124 (N_17124,N_13273,N_12516);
xor U17125 (N_17125,N_11640,N_14593);
nand U17126 (N_17126,N_14287,N_14253);
and U17127 (N_17127,N_11714,N_13704);
nand U17128 (N_17128,N_14974,N_10137);
and U17129 (N_17129,N_11978,N_13350);
nor U17130 (N_17130,N_12443,N_14480);
and U17131 (N_17131,N_12389,N_12088);
nand U17132 (N_17132,N_11115,N_12421);
nor U17133 (N_17133,N_14400,N_12945);
or U17134 (N_17134,N_10916,N_11844);
nand U17135 (N_17135,N_14935,N_12917);
xor U17136 (N_17136,N_11198,N_10809);
and U17137 (N_17137,N_10990,N_12356);
nand U17138 (N_17138,N_10665,N_14541);
nand U17139 (N_17139,N_13845,N_13209);
nand U17140 (N_17140,N_11900,N_10110);
nand U17141 (N_17141,N_10632,N_11162);
and U17142 (N_17142,N_14835,N_11555);
nand U17143 (N_17143,N_13666,N_13283);
nor U17144 (N_17144,N_12289,N_14147);
or U17145 (N_17145,N_14353,N_14271);
nand U17146 (N_17146,N_10652,N_13181);
nand U17147 (N_17147,N_11536,N_13261);
nor U17148 (N_17148,N_12119,N_13725);
and U17149 (N_17149,N_10849,N_13616);
nand U17150 (N_17150,N_14995,N_12384);
nor U17151 (N_17151,N_11831,N_10513);
and U17152 (N_17152,N_14540,N_13795);
or U17153 (N_17153,N_12985,N_12090);
nor U17154 (N_17154,N_10051,N_10326);
or U17155 (N_17155,N_11215,N_14140);
or U17156 (N_17156,N_10822,N_11863);
nand U17157 (N_17157,N_14348,N_12909);
and U17158 (N_17158,N_12501,N_11586);
nor U17159 (N_17159,N_14120,N_11419);
nor U17160 (N_17160,N_10168,N_14092);
and U17161 (N_17161,N_11771,N_11624);
or U17162 (N_17162,N_11019,N_10040);
xnor U17163 (N_17163,N_14924,N_13422);
nand U17164 (N_17164,N_14790,N_12039);
and U17165 (N_17165,N_10500,N_14695);
or U17166 (N_17166,N_14509,N_14983);
nor U17167 (N_17167,N_12561,N_12295);
or U17168 (N_17168,N_14171,N_14132);
or U17169 (N_17169,N_14664,N_11647);
nor U17170 (N_17170,N_12346,N_14441);
or U17171 (N_17171,N_11426,N_14119);
xor U17172 (N_17172,N_11090,N_12223);
and U17173 (N_17173,N_14736,N_13612);
nor U17174 (N_17174,N_13560,N_10684);
or U17175 (N_17175,N_14543,N_13319);
or U17176 (N_17176,N_10927,N_14829);
or U17177 (N_17177,N_14285,N_13245);
nor U17178 (N_17178,N_13096,N_14792);
nand U17179 (N_17179,N_12966,N_12434);
nor U17180 (N_17180,N_11783,N_10757);
or U17181 (N_17181,N_14889,N_13000);
nor U17182 (N_17182,N_10316,N_11790);
or U17183 (N_17183,N_11326,N_11136);
nor U17184 (N_17184,N_10055,N_11458);
and U17185 (N_17185,N_10005,N_14236);
nand U17186 (N_17186,N_10323,N_13517);
xor U17187 (N_17187,N_11451,N_10828);
or U17188 (N_17188,N_12339,N_10644);
and U17189 (N_17189,N_11629,N_11788);
or U17190 (N_17190,N_13748,N_14737);
nand U17191 (N_17191,N_13761,N_10339);
nor U17192 (N_17192,N_11651,N_10227);
xnor U17193 (N_17193,N_14987,N_11525);
nor U17194 (N_17194,N_12031,N_12658);
nand U17195 (N_17195,N_11300,N_14731);
nor U17196 (N_17196,N_12254,N_12948);
nor U17197 (N_17197,N_12307,N_11873);
and U17198 (N_17198,N_13879,N_13663);
nor U17199 (N_17199,N_10029,N_11933);
and U17200 (N_17200,N_10987,N_11960);
nor U17201 (N_17201,N_14747,N_11604);
nor U17202 (N_17202,N_10897,N_11131);
and U17203 (N_17203,N_12202,N_10461);
nor U17204 (N_17204,N_14095,N_14765);
or U17205 (N_17205,N_14437,N_14428);
nand U17206 (N_17206,N_12866,N_11465);
nand U17207 (N_17207,N_13924,N_12323);
nor U17208 (N_17208,N_13885,N_13975);
or U17209 (N_17209,N_11479,N_14312);
or U17210 (N_17210,N_12499,N_14042);
xor U17211 (N_17211,N_14955,N_12972);
nand U17212 (N_17212,N_13358,N_11883);
or U17213 (N_17213,N_13952,N_10295);
and U17214 (N_17214,N_11172,N_12026);
or U17215 (N_17215,N_10412,N_12952);
and U17216 (N_17216,N_10248,N_11567);
or U17217 (N_17217,N_14284,N_10314);
or U17218 (N_17218,N_13272,N_14403);
nand U17219 (N_17219,N_12213,N_13379);
or U17220 (N_17220,N_14094,N_13678);
nand U17221 (N_17221,N_14601,N_14419);
nor U17222 (N_17222,N_12607,N_13375);
or U17223 (N_17223,N_12868,N_12993);
nor U17224 (N_17224,N_11015,N_10734);
and U17225 (N_17225,N_13130,N_14681);
nand U17226 (N_17226,N_13794,N_13140);
and U17227 (N_17227,N_10007,N_14136);
or U17228 (N_17228,N_14365,N_14558);
or U17229 (N_17229,N_12579,N_11283);
or U17230 (N_17230,N_11449,N_14048);
nor U17231 (N_17231,N_10976,N_13965);
nor U17232 (N_17232,N_13151,N_13664);
nor U17233 (N_17233,N_14158,N_11943);
and U17234 (N_17234,N_12245,N_12492);
or U17235 (N_17235,N_13731,N_12883);
and U17236 (N_17236,N_11981,N_12627);
or U17237 (N_17237,N_14687,N_11159);
or U17238 (N_17238,N_12066,N_12549);
or U17239 (N_17239,N_12836,N_13456);
or U17240 (N_17240,N_11196,N_10950);
nor U17241 (N_17241,N_10770,N_12122);
nor U17242 (N_17242,N_10032,N_14363);
or U17243 (N_17243,N_12955,N_12750);
nor U17244 (N_17244,N_14734,N_11648);
and U17245 (N_17245,N_11344,N_13303);
xnor U17246 (N_17246,N_13852,N_10952);
and U17247 (N_17247,N_13099,N_12977);
or U17248 (N_17248,N_14248,N_13349);
or U17249 (N_17249,N_10130,N_13522);
xor U17250 (N_17250,N_14316,N_11487);
and U17251 (N_17251,N_14640,N_11278);
and U17252 (N_17252,N_14257,N_12085);
or U17253 (N_17253,N_13487,N_11298);
nand U17254 (N_17254,N_13208,N_13997);
nand U17255 (N_17255,N_12027,N_14377);
and U17256 (N_17256,N_11118,N_12572);
or U17257 (N_17257,N_10639,N_14587);
or U17258 (N_17258,N_10964,N_12255);
nor U17259 (N_17259,N_10201,N_14631);
nor U17260 (N_17260,N_11511,N_12843);
xor U17261 (N_17261,N_11765,N_13674);
nand U17262 (N_17262,N_13990,N_12171);
nor U17263 (N_17263,N_13882,N_14958);
or U17264 (N_17264,N_12049,N_13039);
or U17265 (N_17265,N_10547,N_14804);
nor U17266 (N_17266,N_10081,N_13005);
or U17267 (N_17267,N_11632,N_14454);
xor U17268 (N_17268,N_13697,N_12241);
nor U17269 (N_17269,N_10064,N_11433);
nor U17270 (N_17270,N_11100,N_12785);
nand U17271 (N_17271,N_11947,N_11362);
nand U17272 (N_17272,N_11850,N_13535);
xor U17273 (N_17273,N_13653,N_10694);
and U17274 (N_17274,N_12557,N_13329);
nor U17275 (N_17275,N_12080,N_10499);
and U17276 (N_17276,N_13441,N_11855);
and U17277 (N_17277,N_10194,N_13334);
nor U17278 (N_17278,N_14843,N_14724);
nor U17279 (N_17279,N_10214,N_14245);
nor U17280 (N_17280,N_13800,N_12152);
or U17281 (N_17281,N_14021,N_11932);
nor U17282 (N_17282,N_11026,N_12259);
or U17283 (N_17283,N_11330,N_13899);
nor U17284 (N_17284,N_11072,N_11737);
nand U17285 (N_17285,N_10815,N_10234);
and U17286 (N_17286,N_14917,N_10038);
nand U17287 (N_17287,N_10107,N_10394);
nor U17288 (N_17288,N_10156,N_14689);
and U17289 (N_17289,N_13294,N_12327);
nand U17290 (N_17290,N_14679,N_12009);
nor U17291 (N_17291,N_11615,N_11068);
or U17292 (N_17292,N_11361,N_11752);
nand U17293 (N_17293,N_11384,N_11687);
and U17294 (N_17294,N_10242,N_10413);
xor U17295 (N_17295,N_11675,N_12500);
nor U17296 (N_17296,N_12915,N_11116);
or U17297 (N_17297,N_14434,N_12803);
and U17298 (N_17298,N_11421,N_11272);
nor U17299 (N_17299,N_13649,N_11295);
or U17300 (N_17300,N_14135,N_12108);
xor U17301 (N_17301,N_14556,N_13288);
nand U17302 (N_17302,N_11309,N_13136);
xor U17303 (N_17303,N_12541,N_11868);
or U17304 (N_17304,N_11523,N_10932);
or U17305 (N_17305,N_10789,N_11008);
xnor U17306 (N_17306,N_13556,N_11702);
and U17307 (N_17307,N_14784,N_10969);
nand U17308 (N_17308,N_14504,N_10827);
xnor U17309 (N_17309,N_14455,N_13687);
xnor U17310 (N_17310,N_10728,N_13757);
nand U17311 (N_17311,N_14106,N_14294);
or U17312 (N_17312,N_12445,N_11888);
nor U17313 (N_17313,N_13127,N_14493);
and U17314 (N_17314,N_11777,N_11756);
xor U17315 (N_17315,N_12308,N_14130);
and U17316 (N_17316,N_11474,N_12926);
nand U17317 (N_17317,N_12789,N_10363);
and U17318 (N_17318,N_10883,N_11731);
xor U17319 (N_17319,N_10901,N_13370);
xor U17320 (N_17320,N_10432,N_13326);
and U17321 (N_17321,N_12462,N_11939);
and U17322 (N_17322,N_13815,N_14591);
nor U17323 (N_17323,N_11491,N_12554);
or U17324 (N_17324,N_10996,N_13857);
xor U17325 (N_17325,N_13825,N_13013);
nor U17326 (N_17326,N_11749,N_11450);
nand U17327 (N_17327,N_13861,N_14196);
xnor U17328 (N_17328,N_11773,N_12385);
nor U17329 (N_17329,N_12146,N_13369);
nor U17330 (N_17330,N_11327,N_12151);
xnor U17331 (N_17331,N_11899,N_12493);
nor U17332 (N_17332,N_13094,N_13873);
nand U17333 (N_17333,N_11013,N_13386);
xnor U17334 (N_17334,N_14081,N_14295);
and U17335 (N_17335,N_11302,N_11980);
xnor U17336 (N_17336,N_11606,N_10404);
nor U17337 (N_17337,N_10350,N_10831);
and U17338 (N_17338,N_10607,N_11192);
nor U17339 (N_17339,N_11027,N_12224);
nor U17340 (N_17340,N_13189,N_13638);
or U17341 (N_17341,N_13980,N_12414);
nand U17342 (N_17342,N_13843,N_13758);
xnor U17343 (N_17343,N_10859,N_12897);
or U17344 (N_17344,N_12964,N_13083);
xor U17345 (N_17345,N_12784,N_12201);
and U17346 (N_17346,N_14694,N_10531);
or U17347 (N_17347,N_13655,N_12393);
and U17348 (N_17348,N_14950,N_12321);
and U17349 (N_17349,N_13139,N_11591);
nor U17350 (N_17350,N_14582,N_10364);
nand U17351 (N_17351,N_14205,N_12716);
nand U17352 (N_17352,N_10705,N_10288);
and U17353 (N_17353,N_13865,N_13118);
xnor U17354 (N_17354,N_10312,N_14233);
nor U17355 (N_17355,N_14198,N_10053);
nand U17356 (N_17356,N_12502,N_14668);
xor U17357 (N_17357,N_10052,N_13716);
nor U17358 (N_17358,N_10533,N_14028);
and U17359 (N_17359,N_14370,N_12059);
nor U17360 (N_17360,N_11082,N_11442);
nand U17361 (N_17361,N_14473,N_14046);
and U17362 (N_17362,N_11942,N_12908);
nor U17363 (N_17363,N_10457,N_10532);
nand U17364 (N_17364,N_13187,N_12079);
or U17365 (N_17365,N_10636,N_14825);
nand U17366 (N_17366,N_10643,N_14194);
xor U17367 (N_17367,N_10735,N_12925);
nor U17368 (N_17368,N_11240,N_14491);
or U17369 (N_17369,N_11564,N_12279);
and U17370 (N_17370,N_14984,N_10165);
nor U17371 (N_17371,N_12076,N_11457);
and U17372 (N_17372,N_11794,N_12014);
and U17373 (N_17373,N_14425,N_11782);
nand U17374 (N_17374,N_11076,N_10892);
and U17375 (N_17375,N_10539,N_10388);
and U17376 (N_17376,N_10153,N_13759);
or U17377 (N_17377,N_13665,N_14802);
or U17378 (N_17378,N_10506,N_11963);
or U17379 (N_17379,N_14861,N_14231);
nand U17380 (N_17380,N_11815,N_11483);
and U17381 (N_17381,N_11556,N_11308);
or U17382 (N_17382,N_13372,N_13053);
or U17383 (N_17383,N_13009,N_13289);
and U17384 (N_17384,N_11030,N_13086);
xnor U17385 (N_17385,N_11352,N_10600);
xor U17386 (N_17386,N_14988,N_14500);
nor U17387 (N_17387,N_13161,N_10429);
xor U17388 (N_17388,N_12875,N_10805);
nor U17389 (N_17389,N_10228,N_14519);
and U17390 (N_17390,N_11305,N_12880);
and U17391 (N_17391,N_11016,N_14052);
and U17392 (N_17392,N_11406,N_10250);
nand U17393 (N_17393,N_11294,N_13120);
and U17394 (N_17394,N_12668,N_11365);
nor U17395 (N_17395,N_12870,N_14685);
xnor U17396 (N_17396,N_10162,N_12997);
and U17397 (N_17397,N_10951,N_14421);
or U17398 (N_17398,N_11598,N_11682);
nor U17399 (N_17399,N_12134,N_11537);
and U17400 (N_17400,N_14929,N_14920);
and U17401 (N_17401,N_12208,N_10668);
nor U17402 (N_17402,N_14440,N_14673);
nand U17403 (N_17403,N_11609,N_11582);
or U17404 (N_17404,N_11641,N_13848);
nand U17405 (N_17405,N_13119,N_10405);
nor U17406 (N_17406,N_11827,N_14190);
nand U17407 (N_17407,N_14266,N_12823);
nor U17408 (N_17408,N_14354,N_10241);
and U17409 (N_17409,N_11377,N_14763);
nand U17410 (N_17410,N_10605,N_12015);
and U17411 (N_17411,N_14609,N_14669);
and U17412 (N_17412,N_12934,N_12396);
nand U17413 (N_17413,N_10261,N_10421);
nor U17414 (N_17414,N_12310,N_12196);
xnor U17415 (N_17415,N_11828,N_10602);
and U17416 (N_17416,N_11806,N_11999);
and U17417 (N_17417,N_12367,N_13237);
nand U17418 (N_17418,N_13224,N_10073);
nor U17419 (N_17419,N_11772,N_13936);
or U17420 (N_17420,N_14426,N_11267);
nand U17421 (N_17421,N_12967,N_11051);
and U17422 (N_17422,N_10485,N_13850);
nor U17423 (N_17423,N_11822,N_10247);
or U17424 (N_17424,N_14169,N_12765);
nand U17425 (N_17425,N_12256,N_10818);
nand U17426 (N_17426,N_11228,N_11329);
and U17427 (N_17427,N_14612,N_11892);
or U17428 (N_17428,N_14770,N_12269);
xor U17429 (N_17429,N_10790,N_11869);
and U17430 (N_17430,N_14854,N_12752);
nor U17431 (N_17431,N_14166,N_10689);
xor U17432 (N_17432,N_14943,N_13959);
or U17433 (N_17433,N_10924,N_10482);
and U17434 (N_17434,N_14289,N_10508);
xor U17435 (N_17435,N_13243,N_14699);
and U17436 (N_17436,N_11544,N_13014);
nand U17437 (N_17437,N_13883,N_12018);
and U17438 (N_17438,N_11077,N_13932);
nor U17439 (N_17439,N_13246,N_11185);
or U17440 (N_17440,N_12121,N_13654);
and U17441 (N_17441,N_12657,N_10564);
nor U17442 (N_17442,N_10514,N_13875);
and U17443 (N_17443,N_13910,N_12677);
nor U17444 (N_17444,N_14814,N_10263);
nor U17445 (N_17445,N_13482,N_11452);
and U17446 (N_17446,N_14730,N_14650);
or U17447 (N_17447,N_12761,N_14946);
or U17448 (N_17448,N_13567,N_14697);
nor U17449 (N_17449,N_10310,N_10839);
xnor U17450 (N_17450,N_12216,N_14358);
or U17451 (N_17451,N_10361,N_10708);
nand U17452 (N_17452,N_13121,N_10645);
nor U17453 (N_17453,N_13904,N_13125);
xor U17454 (N_17454,N_14808,N_11517);
xnor U17455 (N_17455,N_11800,N_12482);
nand U17456 (N_17456,N_13908,N_14014);
or U17457 (N_17457,N_11057,N_11798);
nand U17458 (N_17458,N_11617,N_10025);
or U17459 (N_17459,N_14866,N_14900);
nand U17460 (N_17460,N_14343,N_13701);
xnor U17461 (N_17461,N_10881,N_11607);
xnor U17462 (N_17462,N_14173,N_13520);
nor U17463 (N_17463,N_11412,N_12232);
nand U17464 (N_17464,N_11343,N_14732);
and U17465 (N_17465,N_11096,N_12522);
and U17466 (N_17466,N_11493,N_12302);
nand U17467 (N_17467,N_10998,N_12696);
nor U17468 (N_17468,N_11232,N_10209);
nor U17469 (N_17469,N_11518,N_10440);
nand U17470 (N_17470,N_11276,N_12867);
nand U17471 (N_17471,N_14254,N_13058);
nand U17472 (N_17472,N_14715,N_12127);
and U17473 (N_17473,N_14402,N_11967);
or U17474 (N_17474,N_14576,N_13194);
or U17475 (N_17475,N_12574,N_10101);
nand U17476 (N_17476,N_12698,N_14160);
nand U17477 (N_17477,N_11940,N_13880);
and U17478 (N_17478,N_12503,N_13770);
nand U17479 (N_17479,N_11904,N_10036);
or U17480 (N_17480,N_10142,N_13512);
or U17481 (N_17481,N_11596,N_10628);
nand U17482 (N_17482,N_10391,N_10212);
nor U17483 (N_17483,N_11446,N_14352);
nand U17484 (N_17484,N_12235,N_13022);
nor U17485 (N_17485,N_13993,N_14138);
nand U17486 (N_17486,N_11014,N_14672);
nor U17487 (N_17487,N_10238,N_12537);
or U17488 (N_17488,N_13525,N_11642);
xor U17489 (N_17489,N_11404,N_14552);
nor U17490 (N_17490,N_10653,N_10444);
nor U17491 (N_17491,N_14525,N_10304);
or U17492 (N_17492,N_11156,N_10618);
nand U17493 (N_17493,N_12990,N_12740);
nand U17494 (N_17494,N_14723,N_14786);
nor U17495 (N_17495,N_13028,N_11620);
or U17496 (N_17496,N_11439,N_13728);
nand U17497 (N_17497,N_13428,N_12519);
nand U17498 (N_17498,N_11010,N_13190);
nand U17499 (N_17499,N_14510,N_11529);
and U17500 (N_17500,N_10446,N_12663);
nand U17501 (N_17501,N_12643,N_11359);
and U17502 (N_17502,N_14622,N_10108);
or U17503 (N_17503,N_13906,N_11655);
nor U17504 (N_17504,N_13723,N_10001);
nand U17505 (N_17505,N_10055,N_10142);
nor U17506 (N_17506,N_14094,N_12104);
xnor U17507 (N_17507,N_10232,N_10159);
or U17508 (N_17508,N_13210,N_13606);
and U17509 (N_17509,N_13525,N_13585);
xnor U17510 (N_17510,N_10185,N_10568);
xnor U17511 (N_17511,N_13562,N_12116);
and U17512 (N_17512,N_10367,N_13824);
and U17513 (N_17513,N_10123,N_10719);
nand U17514 (N_17514,N_14666,N_12135);
and U17515 (N_17515,N_14289,N_10513);
and U17516 (N_17516,N_13168,N_13680);
nand U17517 (N_17517,N_12024,N_10570);
and U17518 (N_17518,N_12933,N_11213);
xor U17519 (N_17519,N_13002,N_14759);
nor U17520 (N_17520,N_13488,N_11243);
nand U17521 (N_17521,N_13557,N_12317);
and U17522 (N_17522,N_12817,N_14040);
and U17523 (N_17523,N_11380,N_14075);
xnor U17524 (N_17524,N_13817,N_13336);
xor U17525 (N_17525,N_10869,N_12800);
nand U17526 (N_17526,N_10152,N_11128);
nor U17527 (N_17527,N_12302,N_12334);
or U17528 (N_17528,N_10904,N_14072);
or U17529 (N_17529,N_13676,N_11542);
and U17530 (N_17530,N_11994,N_12310);
and U17531 (N_17531,N_12412,N_14195);
nand U17532 (N_17532,N_10729,N_14096);
xor U17533 (N_17533,N_14734,N_12577);
nor U17534 (N_17534,N_12329,N_11150);
nand U17535 (N_17535,N_12642,N_11611);
nor U17536 (N_17536,N_11594,N_12743);
or U17537 (N_17537,N_12798,N_13569);
xnor U17538 (N_17538,N_12220,N_11789);
xor U17539 (N_17539,N_10912,N_13658);
or U17540 (N_17540,N_12146,N_11294);
nand U17541 (N_17541,N_14363,N_14627);
nand U17542 (N_17542,N_14444,N_13784);
or U17543 (N_17543,N_14187,N_11732);
and U17544 (N_17544,N_14505,N_10431);
nor U17545 (N_17545,N_13287,N_14143);
and U17546 (N_17546,N_10421,N_12475);
nor U17547 (N_17547,N_11773,N_11709);
and U17548 (N_17548,N_10378,N_11519);
and U17549 (N_17549,N_14540,N_13842);
and U17550 (N_17550,N_14434,N_13554);
and U17551 (N_17551,N_11146,N_11258);
or U17552 (N_17552,N_10219,N_13479);
nor U17553 (N_17553,N_14893,N_12270);
and U17554 (N_17554,N_11903,N_12089);
or U17555 (N_17555,N_11755,N_14741);
xor U17556 (N_17556,N_11169,N_13391);
nor U17557 (N_17557,N_12884,N_12297);
or U17558 (N_17558,N_13360,N_10808);
nand U17559 (N_17559,N_13721,N_12118);
xor U17560 (N_17560,N_10560,N_13478);
and U17561 (N_17561,N_12980,N_10913);
nand U17562 (N_17562,N_10727,N_14964);
or U17563 (N_17563,N_10699,N_11239);
and U17564 (N_17564,N_13949,N_14330);
nand U17565 (N_17565,N_13400,N_13232);
and U17566 (N_17566,N_12151,N_14574);
nor U17567 (N_17567,N_13709,N_11116);
nor U17568 (N_17568,N_13161,N_12258);
and U17569 (N_17569,N_13491,N_10749);
nor U17570 (N_17570,N_14103,N_10085);
and U17571 (N_17571,N_14032,N_11186);
or U17572 (N_17572,N_11235,N_12834);
and U17573 (N_17573,N_10521,N_13524);
and U17574 (N_17574,N_14228,N_14664);
nor U17575 (N_17575,N_10889,N_13246);
nor U17576 (N_17576,N_13419,N_10556);
and U17577 (N_17577,N_14158,N_13416);
nand U17578 (N_17578,N_12863,N_13889);
nor U17579 (N_17579,N_14472,N_12923);
nand U17580 (N_17580,N_12514,N_14321);
nor U17581 (N_17581,N_12602,N_13204);
and U17582 (N_17582,N_11754,N_12487);
or U17583 (N_17583,N_14362,N_12278);
nand U17584 (N_17584,N_14126,N_12219);
and U17585 (N_17585,N_12018,N_10018);
or U17586 (N_17586,N_14542,N_14500);
nand U17587 (N_17587,N_12906,N_14045);
nand U17588 (N_17588,N_13092,N_14419);
and U17589 (N_17589,N_10336,N_10736);
or U17590 (N_17590,N_12456,N_12202);
and U17591 (N_17591,N_13270,N_14042);
nand U17592 (N_17592,N_12963,N_10934);
nor U17593 (N_17593,N_14062,N_14257);
and U17594 (N_17594,N_14893,N_13018);
or U17595 (N_17595,N_12880,N_10115);
and U17596 (N_17596,N_12683,N_11091);
nor U17597 (N_17597,N_11589,N_13495);
or U17598 (N_17598,N_14973,N_12570);
and U17599 (N_17599,N_12105,N_13563);
xnor U17600 (N_17600,N_14629,N_10514);
nor U17601 (N_17601,N_13036,N_13263);
nor U17602 (N_17602,N_11065,N_14369);
and U17603 (N_17603,N_14349,N_13147);
nand U17604 (N_17604,N_11610,N_10702);
nand U17605 (N_17605,N_13663,N_11071);
or U17606 (N_17606,N_11893,N_13255);
nor U17607 (N_17607,N_11233,N_13063);
nor U17608 (N_17608,N_13101,N_11068);
or U17609 (N_17609,N_14168,N_10464);
and U17610 (N_17610,N_14541,N_10732);
or U17611 (N_17611,N_12762,N_11946);
and U17612 (N_17612,N_10156,N_11769);
nand U17613 (N_17613,N_10797,N_14893);
and U17614 (N_17614,N_11251,N_10826);
nor U17615 (N_17615,N_11963,N_13613);
xnor U17616 (N_17616,N_12516,N_12491);
or U17617 (N_17617,N_11060,N_12737);
or U17618 (N_17618,N_11254,N_13554);
nand U17619 (N_17619,N_14744,N_10023);
or U17620 (N_17620,N_12646,N_11778);
nand U17621 (N_17621,N_10484,N_12066);
and U17622 (N_17622,N_10973,N_11303);
nand U17623 (N_17623,N_14980,N_13349);
nor U17624 (N_17624,N_14757,N_13367);
or U17625 (N_17625,N_14106,N_11875);
or U17626 (N_17626,N_11331,N_10851);
and U17627 (N_17627,N_14350,N_14009);
nor U17628 (N_17628,N_13473,N_12955);
and U17629 (N_17629,N_11094,N_13704);
or U17630 (N_17630,N_13688,N_12467);
or U17631 (N_17631,N_12284,N_14926);
and U17632 (N_17632,N_11296,N_13574);
nand U17633 (N_17633,N_13079,N_11932);
or U17634 (N_17634,N_12368,N_14086);
nor U17635 (N_17635,N_10293,N_14878);
and U17636 (N_17636,N_10922,N_14730);
nor U17637 (N_17637,N_14138,N_11552);
nand U17638 (N_17638,N_10109,N_14693);
and U17639 (N_17639,N_14085,N_12461);
nand U17640 (N_17640,N_14531,N_14449);
and U17641 (N_17641,N_10693,N_11315);
or U17642 (N_17642,N_13834,N_14893);
or U17643 (N_17643,N_13103,N_13213);
xnor U17644 (N_17644,N_10879,N_13040);
nand U17645 (N_17645,N_10276,N_11405);
xnor U17646 (N_17646,N_13315,N_13168);
and U17647 (N_17647,N_14468,N_11047);
or U17648 (N_17648,N_10672,N_10875);
or U17649 (N_17649,N_11205,N_11670);
and U17650 (N_17650,N_13736,N_11917);
nor U17651 (N_17651,N_14572,N_10495);
or U17652 (N_17652,N_10439,N_10662);
nor U17653 (N_17653,N_14527,N_14271);
nand U17654 (N_17654,N_10899,N_14184);
and U17655 (N_17655,N_12636,N_13236);
nand U17656 (N_17656,N_11522,N_14173);
nand U17657 (N_17657,N_14863,N_11200);
nor U17658 (N_17658,N_13445,N_11746);
nand U17659 (N_17659,N_13030,N_10349);
and U17660 (N_17660,N_12282,N_11313);
nand U17661 (N_17661,N_13356,N_14067);
and U17662 (N_17662,N_12538,N_14925);
nor U17663 (N_17663,N_14584,N_10063);
xnor U17664 (N_17664,N_14609,N_12198);
nor U17665 (N_17665,N_11545,N_14152);
and U17666 (N_17666,N_14289,N_10167);
nand U17667 (N_17667,N_12762,N_10863);
nor U17668 (N_17668,N_14755,N_10672);
nor U17669 (N_17669,N_12723,N_10857);
xor U17670 (N_17670,N_12134,N_13565);
nand U17671 (N_17671,N_14765,N_14911);
or U17672 (N_17672,N_10788,N_13123);
and U17673 (N_17673,N_13291,N_11092);
nand U17674 (N_17674,N_12082,N_10315);
xnor U17675 (N_17675,N_10775,N_11945);
xor U17676 (N_17676,N_11833,N_13868);
or U17677 (N_17677,N_10855,N_14916);
xor U17678 (N_17678,N_11683,N_10010);
and U17679 (N_17679,N_11394,N_10226);
nor U17680 (N_17680,N_11916,N_10528);
nor U17681 (N_17681,N_10335,N_11727);
nor U17682 (N_17682,N_10914,N_10771);
or U17683 (N_17683,N_11038,N_11576);
nor U17684 (N_17684,N_14148,N_14874);
xor U17685 (N_17685,N_10748,N_13285);
or U17686 (N_17686,N_12873,N_14447);
or U17687 (N_17687,N_11835,N_11074);
nor U17688 (N_17688,N_13384,N_10404);
and U17689 (N_17689,N_12253,N_14300);
nand U17690 (N_17690,N_10216,N_12584);
or U17691 (N_17691,N_14436,N_12485);
nand U17692 (N_17692,N_13655,N_11111);
and U17693 (N_17693,N_12744,N_11076);
and U17694 (N_17694,N_10900,N_11462);
and U17695 (N_17695,N_10155,N_14005);
and U17696 (N_17696,N_10575,N_10765);
nand U17697 (N_17697,N_10527,N_10490);
and U17698 (N_17698,N_11134,N_10995);
nor U17699 (N_17699,N_13084,N_10108);
or U17700 (N_17700,N_13908,N_10710);
and U17701 (N_17701,N_14873,N_12735);
nand U17702 (N_17702,N_10021,N_12932);
or U17703 (N_17703,N_10610,N_13092);
nand U17704 (N_17704,N_12312,N_11935);
nor U17705 (N_17705,N_11823,N_10514);
nor U17706 (N_17706,N_11544,N_10818);
and U17707 (N_17707,N_14812,N_12289);
or U17708 (N_17708,N_14162,N_14993);
and U17709 (N_17709,N_10351,N_13803);
nor U17710 (N_17710,N_14638,N_13198);
or U17711 (N_17711,N_14793,N_14158);
nor U17712 (N_17712,N_11634,N_10580);
and U17713 (N_17713,N_11502,N_14515);
xor U17714 (N_17714,N_13186,N_12995);
or U17715 (N_17715,N_13013,N_12432);
nand U17716 (N_17716,N_11944,N_12913);
nand U17717 (N_17717,N_13962,N_10589);
and U17718 (N_17718,N_13061,N_13855);
or U17719 (N_17719,N_11588,N_13872);
or U17720 (N_17720,N_13258,N_10228);
nor U17721 (N_17721,N_14741,N_12920);
or U17722 (N_17722,N_13770,N_11956);
or U17723 (N_17723,N_10846,N_13929);
nand U17724 (N_17724,N_12685,N_10028);
xnor U17725 (N_17725,N_14098,N_14954);
or U17726 (N_17726,N_14105,N_10885);
nand U17727 (N_17727,N_10146,N_12906);
nand U17728 (N_17728,N_12429,N_12346);
xor U17729 (N_17729,N_12698,N_12384);
and U17730 (N_17730,N_13191,N_11584);
nand U17731 (N_17731,N_13851,N_10355);
xor U17732 (N_17732,N_12428,N_13690);
xor U17733 (N_17733,N_11520,N_13293);
nor U17734 (N_17734,N_13419,N_14313);
xnor U17735 (N_17735,N_10292,N_12142);
or U17736 (N_17736,N_10184,N_11143);
and U17737 (N_17737,N_12272,N_13249);
nor U17738 (N_17738,N_12806,N_10520);
xnor U17739 (N_17739,N_11990,N_13179);
or U17740 (N_17740,N_13007,N_13641);
nor U17741 (N_17741,N_14466,N_12658);
or U17742 (N_17742,N_12398,N_10058);
xnor U17743 (N_17743,N_10558,N_14775);
xnor U17744 (N_17744,N_12185,N_10919);
xor U17745 (N_17745,N_12019,N_13811);
xor U17746 (N_17746,N_14402,N_11505);
nor U17747 (N_17747,N_13224,N_14397);
nand U17748 (N_17748,N_10085,N_13315);
or U17749 (N_17749,N_11101,N_10339);
and U17750 (N_17750,N_13302,N_10004);
nand U17751 (N_17751,N_14277,N_13466);
and U17752 (N_17752,N_13928,N_13793);
nand U17753 (N_17753,N_13688,N_11542);
nor U17754 (N_17754,N_10036,N_14332);
nand U17755 (N_17755,N_11621,N_13989);
and U17756 (N_17756,N_10443,N_13351);
nand U17757 (N_17757,N_14800,N_14533);
or U17758 (N_17758,N_12608,N_12050);
or U17759 (N_17759,N_12498,N_11652);
nor U17760 (N_17760,N_14444,N_13132);
or U17761 (N_17761,N_14094,N_14794);
and U17762 (N_17762,N_13588,N_12241);
nor U17763 (N_17763,N_13913,N_12798);
nor U17764 (N_17764,N_12339,N_10920);
and U17765 (N_17765,N_10348,N_14906);
or U17766 (N_17766,N_13263,N_14373);
nand U17767 (N_17767,N_11155,N_14617);
or U17768 (N_17768,N_12031,N_11440);
and U17769 (N_17769,N_12503,N_10914);
nand U17770 (N_17770,N_10973,N_14656);
and U17771 (N_17771,N_11828,N_10338);
nor U17772 (N_17772,N_10706,N_11665);
xnor U17773 (N_17773,N_11466,N_11198);
or U17774 (N_17774,N_10793,N_13938);
or U17775 (N_17775,N_11200,N_14144);
nor U17776 (N_17776,N_13891,N_10543);
or U17777 (N_17777,N_11582,N_14025);
nand U17778 (N_17778,N_14517,N_11302);
nand U17779 (N_17779,N_13683,N_12349);
xnor U17780 (N_17780,N_14640,N_13537);
and U17781 (N_17781,N_13294,N_13382);
or U17782 (N_17782,N_11853,N_13419);
or U17783 (N_17783,N_11945,N_13457);
and U17784 (N_17784,N_10578,N_13454);
nand U17785 (N_17785,N_12268,N_11250);
and U17786 (N_17786,N_12681,N_13673);
nand U17787 (N_17787,N_12740,N_11198);
xnor U17788 (N_17788,N_14179,N_11628);
and U17789 (N_17789,N_10334,N_10772);
or U17790 (N_17790,N_13793,N_14835);
nor U17791 (N_17791,N_10752,N_13236);
or U17792 (N_17792,N_13106,N_11497);
xnor U17793 (N_17793,N_11437,N_11294);
nor U17794 (N_17794,N_12555,N_11167);
or U17795 (N_17795,N_11075,N_12315);
or U17796 (N_17796,N_13892,N_10317);
nand U17797 (N_17797,N_11665,N_12687);
and U17798 (N_17798,N_13303,N_11549);
xor U17799 (N_17799,N_13065,N_12004);
and U17800 (N_17800,N_10103,N_12193);
or U17801 (N_17801,N_10660,N_13473);
and U17802 (N_17802,N_14019,N_14037);
or U17803 (N_17803,N_11745,N_12007);
xnor U17804 (N_17804,N_11148,N_13625);
xor U17805 (N_17805,N_13641,N_10306);
nor U17806 (N_17806,N_11344,N_14884);
nor U17807 (N_17807,N_12135,N_13653);
and U17808 (N_17808,N_14133,N_12183);
and U17809 (N_17809,N_13386,N_10175);
nand U17810 (N_17810,N_10837,N_12550);
or U17811 (N_17811,N_10132,N_11709);
and U17812 (N_17812,N_11010,N_10899);
and U17813 (N_17813,N_12380,N_12425);
nand U17814 (N_17814,N_14835,N_11782);
xnor U17815 (N_17815,N_12846,N_14264);
nand U17816 (N_17816,N_13707,N_14827);
and U17817 (N_17817,N_11313,N_13873);
or U17818 (N_17818,N_11382,N_14599);
nand U17819 (N_17819,N_11735,N_11772);
or U17820 (N_17820,N_10689,N_12511);
nand U17821 (N_17821,N_10081,N_10269);
xnor U17822 (N_17822,N_10328,N_10165);
and U17823 (N_17823,N_11582,N_13952);
nand U17824 (N_17824,N_11212,N_13949);
xnor U17825 (N_17825,N_13154,N_11188);
nor U17826 (N_17826,N_11683,N_11328);
nor U17827 (N_17827,N_11573,N_12306);
and U17828 (N_17828,N_14008,N_10085);
or U17829 (N_17829,N_10033,N_10660);
nand U17830 (N_17830,N_14808,N_12313);
nand U17831 (N_17831,N_13506,N_13553);
nor U17832 (N_17832,N_10163,N_14508);
nand U17833 (N_17833,N_10374,N_14186);
nand U17834 (N_17834,N_10206,N_14422);
and U17835 (N_17835,N_10340,N_12795);
or U17836 (N_17836,N_12579,N_10020);
and U17837 (N_17837,N_11271,N_12725);
nand U17838 (N_17838,N_14468,N_12770);
or U17839 (N_17839,N_14908,N_14931);
or U17840 (N_17840,N_14184,N_12875);
nor U17841 (N_17841,N_10875,N_14822);
nor U17842 (N_17842,N_11682,N_10001);
and U17843 (N_17843,N_10516,N_14290);
or U17844 (N_17844,N_10182,N_13719);
or U17845 (N_17845,N_10081,N_13122);
xnor U17846 (N_17846,N_13401,N_13045);
nor U17847 (N_17847,N_14207,N_12297);
and U17848 (N_17848,N_10107,N_14372);
and U17849 (N_17849,N_11123,N_13507);
xor U17850 (N_17850,N_11991,N_12854);
nor U17851 (N_17851,N_14846,N_10508);
nor U17852 (N_17852,N_13614,N_13887);
or U17853 (N_17853,N_14321,N_10571);
or U17854 (N_17854,N_13663,N_10266);
nand U17855 (N_17855,N_14040,N_12918);
nand U17856 (N_17856,N_10081,N_14263);
nor U17857 (N_17857,N_14994,N_13082);
nor U17858 (N_17858,N_10212,N_12362);
nand U17859 (N_17859,N_14029,N_13491);
nand U17860 (N_17860,N_13007,N_14360);
nor U17861 (N_17861,N_13437,N_11564);
nor U17862 (N_17862,N_11347,N_11386);
nor U17863 (N_17863,N_11393,N_10970);
or U17864 (N_17864,N_10290,N_10671);
or U17865 (N_17865,N_12079,N_10747);
and U17866 (N_17866,N_13249,N_13361);
or U17867 (N_17867,N_11286,N_10004);
nor U17868 (N_17868,N_14268,N_11970);
or U17869 (N_17869,N_14830,N_13070);
nor U17870 (N_17870,N_13926,N_11816);
or U17871 (N_17871,N_14040,N_11040);
nor U17872 (N_17872,N_10023,N_13983);
nor U17873 (N_17873,N_12976,N_14676);
and U17874 (N_17874,N_11876,N_12915);
or U17875 (N_17875,N_12741,N_10335);
nor U17876 (N_17876,N_14913,N_10707);
or U17877 (N_17877,N_14739,N_12206);
or U17878 (N_17878,N_12710,N_11869);
and U17879 (N_17879,N_12065,N_10100);
nand U17880 (N_17880,N_13684,N_11356);
nor U17881 (N_17881,N_13152,N_13623);
and U17882 (N_17882,N_11009,N_12692);
nor U17883 (N_17883,N_10726,N_13142);
nand U17884 (N_17884,N_10070,N_10150);
or U17885 (N_17885,N_10718,N_13639);
nor U17886 (N_17886,N_11251,N_13614);
nand U17887 (N_17887,N_13059,N_14585);
or U17888 (N_17888,N_11288,N_14534);
or U17889 (N_17889,N_11856,N_12110);
or U17890 (N_17890,N_12975,N_12974);
nand U17891 (N_17891,N_12280,N_10977);
nor U17892 (N_17892,N_12344,N_12950);
or U17893 (N_17893,N_12812,N_10962);
and U17894 (N_17894,N_13315,N_13046);
nor U17895 (N_17895,N_11234,N_12340);
and U17896 (N_17896,N_11566,N_10211);
nor U17897 (N_17897,N_14213,N_10592);
nand U17898 (N_17898,N_13884,N_13276);
and U17899 (N_17899,N_13964,N_14330);
or U17900 (N_17900,N_12161,N_11467);
or U17901 (N_17901,N_10241,N_10417);
nand U17902 (N_17902,N_14163,N_12952);
nor U17903 (N_17903,N_13809,N_10930);
and U17904 (N_17904,N_13833,N_13279);
nand U17905 (N_17905,N_11254,N_10134);
or U17906 (N_17906,N_13208,N_14237);
and U17907 (N_17907,N_14202,N_12838);
nor U17908 (N_17908,N_10912,N_12980);
xor U17909 (N_17909,N_14217,N_14444);
xnor U17910 (N_17910,N_10245,N_12538);
nor U17911 (N_17911,N_14676,N_12178);
or U17912 (N_17912,N_14167,N_10079);
and U17913 (N_17913,N_11835,N_10808);
and U17914 (N_17914,N_14078,N_10629);
xor U17915 (N_17915,N_12876,N_10084);
nor U17916 (N_17916,N_13765,N_13700);
xor U17917 (N_17917,N_14250,N_11001);
and U17918 (N_17918,N_14596,N_10087);
or U17919 (N_17919,N_14822,N_14048);
or U17920 (N_17920,N_12449,N_12667);
or U17921 (N_17921,N_11240,N_14735);
nor U17922 (N_17922,N_13028,N_12451);
nand U17923 (N_17923,N_12402,N_14756);
xor U17924 (N_17924,N_10224,N_11138);
and U17925 (N_17925,N_14841,N_14493);
and U17926 (N_17926,N_10720,N_14046);
nand U17927 (N_17927,N_13085,N_10066);
and U17928 (N_17928,N_13636,N_12116);
nor U17929 (N_17929,N_13312,N_13622);
or U17930 (N_17930,N_12161,N_11967);
nand U17931 (N_17931,N_14853,N_11168);
or U17932 (N_17932,N_11232,N_10295);
xnor U17933 (N_17933,N_14664,N_14459);
nor U17934 (N_17934,N_12289,N_13886);
or U17935 (N_17935,N_11366,N_10783);
or U17936 (N_17936,N_14261,N_11978);
nand U17937 (N_17937,N_14521,N_11311);
nor U17938 (N_17938,N_11955,N_11039);
nor U17939 (N_17939,N_13217,N_13154);
xnor U17940 (N_17940,N_13032,N_11944);
nand U17941 (N_17941,N_14387,N_11863);
and U17942 (N_17942,N_14073,N_13474);
and U17943 (N_17943,N_11519,N_12891);
and U17944 (N_17944,N_10559,N_12859);
nand U17945 (N_17945,N_14941,N_10076);
nand U17946 (N_17946,N_12507,N_11238);
nand U17947 (N_17947,N_10541,N_13017);
nor U17948 (N_17948,N_12606,N_13725);
or U17949 (N_17949,N_10282,N_14735);
nand U17950 (N_17950,N_12859,N_14551);
nor U17951 (N_17951,N_13838,N_13539);
xnor U17952 (N_17952,N_11271,N_14304);
and U17953 (N_17953,N_12442,N_11665);
nor U17954 (N_17954,N_10787,N_11877);
or U17955 (N_17955,N_10529,N_13495);
nand U17956 (N_17956,N_10699,N_14957);
and U17957 (N_17957,N_12781,N_11952);
nand U17958 (N_17958,N_12319,N_14540);
nand U17959 (N_17959,N_11573,N_10020);
nor U17960 (N_17960,N_13224,N_10338);
nand U17961 (N_17961,N_13340,N_12727);
and U17962 (N_17962,N_12008,N_11568);
or U17963 (N_17963,N_12349,N_14161);
nor U17964 (N_17964,N_12636,N_12348);
nor U17965 (N_17965,N_14919,N_13869);
and U17966 (N_17966,N_13899,N_11593);
nor U17967 (N_17967,N_13627,N_14463);
and U17968 (N_17968,N_10564,N_11150);
nand U17969 (N_17969,N_13922,N_14256);
nand U17970 (N_17970,N_12568,N_13203);
and U17971 (N_17971,N_14632,N_11084);
and U17972 (N_17972,N_10744,N_12981);
nand U17973 (N_17973,N_11661,N_12947);
nor U17974 (N_17974,N_10665,N_11627);
or U17975 (N_17975,N_14297,N_13397);
and U17976 (N_17976,N_11504,N_14581);
nand U17977 (N_17977,N_10466,N_13992);
nand U17978 (N_17978,N_14337,N_13664);
and U17979 (N_17979,N_10306,N_10224);
and U17980 (N_17980,N_10615,N_11935);
or U17981 (N_17981,N_14572,N_12145);
and U17982 (N_17982,N_10953,N_10640);
or U17983 (N_17983,N_10181,N_13949);
nor U17984 (N_17984,N_10087,N_11711);
nor U17985 (N_17985,N_13452,N_10403);
or U17986 (N_17986,N_10735,N_11048);
nor U17987 (N_17987,N_10209,N_11136);
nor U17988 (N_17988,N_14286,N_10842);
and U17989 (N_17989,N_12689,N_10053);
nand U17990 (N_17990,N_13499,N_14725);
xor U17991 (N_17991,N_10117,N_14416);
or U17992 (N_17992,N_11442,N_14842);
nor U17993 (N_17993,N_12705,N_14272);
or U17994 (N_17994,N_14373,N_14755);
nand U17995 (N_17995,N_14110,N_14152);
nand U17996 (N_17996,N_10220,N_11524);
nor U17997 (N_17997,N_12766,N_11964);
nor U17998 (N_17998,N_11754,N_10664);
or U17999 (N_17999,N_12648,N_12792);
and U18000 (N_18000,N_11034,N_13100);
or U18001 (N_18001,N_11585,N_14196);
and U18002 (N_18002,N_13259,N_12244);
and U18003 (N_18003,N_13700,N_13060);
nand U18004 (N_18004,N_12118,N_10905);
nand U18005 (N_18005,N_10828,N_13479);
nand U18006 (N_18006,N_12721,N_13678);
xor U18007 (N_18007,N_14797,N_11455);
xor U18008 (N_18008,N_14285,N_14456);
nor U18009 (N_18009,N_11883,N_10574);
and U18010 (N_18010,N_14801,N_11743);
or U18011 (N_18011,N_12735,N_10068);
nor U18012 (N_18012,N_11091,N_12585);
and U18013 (N_18013,N_11825,N_13640);
or U18014 (N_18014,N_14501,N_12066);
or U18015 (N_18015,N_14320,N_12037);
xor U18016 (N_18016,N_13358,N_11532);
or U18017 (N_18017,N_11836,N_14492);
nand U18018 (N_18018,N_12616,N_11423);
nand U18019 (N_18019,N_11079,N_11362);
nand U18020 (N_18020,N_11770,N_10422);
nand U18021 (N_18021,N_13270,N_12673);
and U18022 (N_18022,N_12928,N_13907);
nand U18023 (N_18023,N_14945,N_12855);
nand U18024 (N_18024,N_13500,N_13601);
or U18025 (N_18025,N_11370,N_14699);
nor U18026 (N_18026,N_10920,N_10279);
and U18027 (N_18027,N_12601,N_10290);
and U18028 (N_18028,N_13149,N_12103);
nand U18029 (N_18029,N_14314,N_10161);
or U18030 (N_18030,N_10863,N_13416);
nand U18031 (N_18031,N_10454,N_10923);
or U18032 (N_18032,N_13679,N_13594);
and U18033 (N_18033,N_13754,N_13047);
xnor U18034 (N_18034,N_13537,N_14405);
xor U18035 (N_18035,N_11018,N_12026);
and U18036 (N_18036,N_12623,N_12666);
xnor U18037 (N_18037,N_13029,N_12269);
xnor U18038 (N_18038,N_13288,N_10448);
nor U18039 (N_18039,N_12722,N_12323);
and U18040 (N_18040,N_11032,N_12942);
or U18041 (N_18041,N_11497,N_14603);
and U18042 (N_18042,N_10430,N_10194);
nand U18043 (N_18043,N_12970,N_14817);
nand U18044 (N_18044,N_13976,N_12023);
or U18045 (N_18045,N_12287,N_11031);
nor U18046 (N_18046,N_13187,N_11025);
nor U18047 (N_18047,N_14542,N_11133);
nor U18048 (N_18048,N_11240,N_10936);
or U18049 (N_18049,N_10349,N_11211);
and U18050 (N_18050,N_14209,N_10093);
xor U18051 (N_18051,N_11225,N_13250);
nor U18052 (N_18052,N_11318,N_10395);
and U18053 (N_18053,N_11808,N_12754);
and U18054 (N_18054,N_10993,N_12752);
nand U18055 (N_18055,N_14773,N_10393);
and U18056 (N_18056,N_11332,N_13106);
xor U18057 (N_18057,N_14639,N_14606);
nor U18058 (N_18058,N_10118,N_11946);
or U18059 (N_18059,N_10620,N_14790);
nand U18060 (N_18060,N_11597,N_12311);
nor U18061 (N_18061,N_14893,N_11282);
nor U18062 (N_18062,N_13521,N_12093);
nor U18063 (N_18063,N_14986,N_12639);
nor U18064 (N_18064,N_12768,N_11192);
nor U18065 (N_18065,N_14391,N_10355);
nand U18066 (N_18066,N_11251,N_14710);
or U18067 (N_18067,N_11810,N_12734);
and U18068 (N_18068,N_14098,N_13075);
nor U18069 (N_18069,N_11311,N_14881);
or U18070 (N_18070,N_10693,N_13595);
nor U18071 (N_18071,N_10016,N_10329);
nand U18072 (N_18072,N_12801,N_14040);
xor U18073 (N_18073,N_14927,N_14112);
or U18074 (N_18074,N_11938,N_13593);
nor U18075 (N_18075,N_11502,N_10083);
and U18076 (N_18076,N_14406,N_10052);
and U18077 (N_18077,N_14824,N_14613);
and U18078 (N_18078,N_12883,N_10463);
nor U18079 (N_18079,N_10400,N_14206);
or U18080 (N_18080,N_12213,N_10311);
nand U18081 (N_18081,N_11315,N_14502);
or U18082 (N_18082,N_14202,N_14746);
nor U18083 (N_18083,N_13738,N_14533);
or U18084 (N_18084,N_13746,N_10488);
nand U18085 (N_18085,N_10436,N_10719);
and U18086 (N_18086,N_11717,N_13331);
nor U18087 (N_18087,N_13259,N_14875);
or U18088 (N_18088,N_13084,N_12055);
and U18089 (N_18089,N_11032,N_14700);
nor U18090 (N_18090,N_14563,N_10584);
or U18091 (N_18091,N_14173,N_14188);
nand U18092 (N_18092,N_14491,N_11616);
and U18093 (N_18093,N_13862,N_12363);
nand U18094 (N_18094,N_11417,N_11998);
or U18095 (N_18095,N_13718,N_10227);
and U18096 (N_18096,N_10776,N_10262);
or U18097 (N_18097,N_10846,N_12596);
nand U18098 (N_18098,N_10432,N_11726);
nor U18099 (N_18099,N_12216,N_13046);
and U18100 (N_18100,N_14855,N_12723);
and U18101 (N_18101,N_11454,N_10647);
or U18102 (N_18102,N_10529,N_12664);
nor U18103 (N_18103,N_13416,N_14757);
xor U18104 (N_18104,N_12268,N_12918);
nor U18105 (N_18105,N_11616,N_13581);
nand U18106 (N_18106,N_12123,N_10478);
nand U18107 (N_18107,N_13427,N_11056);
or U18108 (N_18108,N_13030,N_11101);
or U18109 (N_18109,N_10697,N_14458);
or U18110 (N_18110,N_10246,N_10261);
and U18111 (N_18111,N_14272,N_13801);
xnor U18112 (N_18112,N_14934,N_12317);
nand U18113 (N_18113,N_11969,N_14000);
or U18114 (N_18114,N_11755,N_13909);
xor U18115 (N_18115,N_12646,N_13783);
nor U18116 (N_18116,N_12493,N_10186);
or U18117 (N_18117,N_13311,N_13897);
nand U18118 (N_18118,N_14587,N_14659);
nor U18119 (N_18119,N_10606,N_11704);
nor U18120 (N_18120,N_12464,N_10522);
or U18121 (N_18121,N_10707,N_10728);
nand U18122 (N_18122,N_12598,N_14255);
and U18123 (N_18123,N_11067,N_13862);
nand U18124 (N_18124,N_13420,N_11108);
nor U18125 (N_18125,N_13578,N_11091);
xor U18126 (N_18126,N_11821,N_12154);
nor U18127 (N_18127,N_12536,N_13767);
and U18128 (N_18128,N_10240,N_10841);
and U18129 (N_18129,N_12890,N_10930);
xnor U18130 (N_18130,N_10976,N_14976);
or U18131 (N_18131,N_12556,N_11670);
or U18132 (N_18132,N_12324,N_10958);
and U18133 (N_18133,N_10429,N_14932);
or U18134 (N_18134,N_14364,N_12695);
and U18135 (N_18135,N_10188,N_10544);
nor U18136 (N_18136,N_13496,N_12296);
and U18137 (N_18137,N_10049,N_10439);
or U18138 (N_18138,N_12769,N_14252);
nor U18139 (N_18139,N_12504,N_10916);
nand U18140 (N_18140,N_12217,N_11695);
nand U18141 (N_18141,N_10723,N_13309);
xnor U18142 (N_18142,N_12272,N_14032);
nand U18143 (N_18143,N_12126,N_13629);
and U18144 (N_18144,N_14574,N_11692);
nor U18145 (N_18145,N_13224,N_13413);
nor U18146 (N_18146,N_12726,N_12666);
nand U18147 (N_18147,N_13852,N_13827);
or U18148 (N_18148,N_13852,N_12414);
nand U18149 (N_18149,N_10483,N_11869);
nor U18150 (N_18150,N_14368,N_13094);
and U18151 (N_18151,N_13288,N_10570);
and U18152 (N_18152,N_12597,N_10219);
or U18153 (N_18153,N_14717,N_10944);
xnor U18154 (N_18154,N_10260,N_11717);
or U18155 (N_18155,N_11082,N_12820);
xor U18156 (N_18156,N_12667,N_12800);
or U18157 (N_18157,N_11072,N_14807);
and U18158 (N_18158,N_11854,N_12485);
nand U18159 (N_18159,N_14394,N_10737);
and U18160 (N_18160,N_10429,N_14863);
nor U18161 (N_18161,N_10934,N_11741);
and U18162 (N_18162,N_10878,N_10587);
or U18163 (N_18163,N_13916,N_11233);
nor U18164 (N_18164,N_10649,N_10341);
and U18165 (N_18165,N_12778,N_14899);
or U18166 (N_18166,N_11663,N_14139);
nor U18167 (N_18167,N_10412,N_14935);
and U18168 (N_18168,N_13469,N_11608);
nor U18169 (N_18169,N_10142,N_11996);
or U18170 (N_18170,N_10606,N_12648);
nand U18171 (N_18171,N_14801,N_13896);
and U18172 (N_18172,N_14788,N_14438);
nand U18173 (N_18173,N_12105,N_12566);
nand U18174 (N_18174,N_14669,N_13763);
nor U18175 (N_18175,N_11010,N_11222);
and U18176 (N_18176,N_11020,N_14660);
nor U18177 (N_18177,N_13042,N_14151);
xnor U18178 (N_18178,N_11646,N_13864);
nor U18179 (N_18179,N_10478,N_14939);
xor U18180 (N_18180,N_13728,N_13268);
nand U18181 (N_18181,N_13897,N_14014);
or U18182 (N_18182,N_12985,N_11657);
nand U18183 (N_18183,N_12248,N_12616);
and U18184 (N_18184,N_12598,N_13759);
nand U18185 (N_18185,N_14385,N_10374);
nand U18186 (N_18186,N_10098,N_12730);
and U18187 (N_18187,N_14807,N_11654);
or U18188 (N_18188,N_14415,N_10637);
and U18189 (N_18189,N_10280,N_12313);
nand U18190 (N_18190,N_13391,N_11487);
nand U18191 (N_18191,N_14485,N_11506);
nand U18192 (N_18192,N_12893,N_10977);
nor U18193 (N_18193,N_10625,N_12029);
or U18194 (N_18194,N_11717,N_10531);
xnor U18195 (N_18195,N_13160,N_13799);
or U18196 (N_18196,N_13768,N_11622);
or U18197 (N_18197,N_14689,N_13223);
or U18198 (N_18198,N_10367,N_12452);
xor U18199 (N_18199,N_14867,N_13359);
nor U18200 (N_18200,N_12441,N_12027);
nor U18201 (N_18201,N_11037,N_10801);
nor U18202 (N_18202,N_11846,N_11235);
and U18203 (N_18203,N_14257,N_13060);
nand U18204 (N_18204,N_10547,N_14050);
nand U18205 (N_18205,N_13310,N_14637);
and U18206 (N_18206,N_10373,N_10521);
xor U18207 (N_18207,N_10005,N_14453);
and U18208 (N_18208,N_12704,N_14526);
nor U18209 (N_18209,N_12092,N_14269);
nor U18210 (N_18210,N_11287,N_12367);
or U18211 (N_18211,N_10920,N_11853);
or U18212 (N_18212,N_14179,N_11248);
nor U18213 (N_18213,N_12691,N_11118);
and U18214 (N_18214,N_14308,N_12264);
nand U18215 (N_18215,N_11671,N_14466);
and U18216 (N_18216,N_14798,N_10959);
nor U18217 (N_18217,N_14013,N_10479);
nand U18218 (N_18218,N_13301,N_12874);
nor U18219 (N_18219,N_14974,N_10290);
nand U18220 (N_18220,N_14391,N_14868);
or U18221 (N_18221,N_13460,N_11332);
or U18222 (N_18222,N_11266,N_12934);
nor U18223 (N_18223,N_14777,N_12155);
and U18224 (N_18224,N_13111,N_10003);
nand U18225 (N_18225,N_14597,N_11424);
nand U18226 (N_18226,N_10220,N_14157);
or U18227 (N_18227,N_14103,N_10069);
and U18228 (N_18228,N_10772,N_13065);
or U18229 (N_18229,N_12339,N_12092);
nand U18230 (N_18230,N_10508,N_13842);
nor U18231 (N_18231,N_14733,N_13996);
nand U18232 (N_18232,N_14197,N_14989);
or U18233 (N_18233,N_13301,N_14988);
or U18234 (N_18234,N_10128,N_11427);
or U18235 (N_18235,N_13485,N_13126);
nor U18236 (N_18236,N_14664,N_11755);
nand U18237 (N_18237,N_13347,N_10924);
nand U18238 (N_18238,N_11775,N_10601);
and U18239 (N_18239,N_14934,N_13498);
nand U18240 (N_18240,N_13628,N_11019);
nor U18241 (N_18241,N_12298,N_12365);
and U18242 (N_18242,N_11189,N_10046);
nor U18243 (N_18243,N_13288,N_12532);
and U18244 (N_18244,N_13728,N_12861);
xnor U18245 (N_18245,N_10020,N_14685);
xor U18246 (N_18246,N_14975,N_14337);
and U18247 (N_18247,N_14972,N_12441);
nand U18248 (N_18248,N_11025,N_11599);
and U18249 (N_18249,N_14347,N_10426);
or U18250 (N_18250,N_13050,N_14568);
nor U18251 (N_18251,N_12751,N_10251);
or U18252 (N_18252,N_10040,N_14333);
or U18253 (N_18253,N_11561,N_10054);
and U18254 (N_18254,N_14243,N_12652);
and U18255 (N_18255,N_11630,N_13574);
or U18256 (N_18256,N_12485,N_10545);
and U18257 (N_18257,N_12418,N_12795);
or U18258 (N_18258,N_11152,N_13892);
nand U18259 (N_18259,N_12720,N_11990);
or U18260 (N_18260,N_13299,N_12892);
nor U18261 (N_18261,N_13572,N_11030);
and U18262 (N_18262,N_10014,N_14554);
or U18263 (N_18263,N_13515,N_14268);
nor U18264 (N_18264,N_13063,N_12868);
nor U18265 (N_18265,N_12150,N_10388);
and U18266 (N_18266,N_10550,N_10960);
and U18267 (N_18267,N_10339,N_10242);
nand U18268 (N_18268,N_12824,N_12589);
nand U18269 (N_18269,N_11703,N_12574);
or U18270 (N_18270,N_11918,N_13496);
nor U18271 (N_18271,N_12124,N_10844);
or U18272 (N_18272,N_11284,N_14442);
xor U18273 (N_18273,N_11639,N_10050);
or U18274 (N_18274,N_10392,N_11538);
nand U18275 (N_18275,N_14164,N_10683);
and U18276 (N_18276,N_14439,N_10938);
nand U18277 (N_18277,N_12885,N_11294);
or U18278 (N_18278,N_10875,N_11294);
xnor U18279 (N_18279,N_13452,N_10752);
nor U18280 (N_18280,N_14118,N_12673);
nand U18281 (N_18281,N_11088,N_10616);
nand U18282 (N_18282,N_12135,N_12063);
nor U18283 (N_18283,N_13157,N_10315);
nor U18284 (N_18284,N_12909,N_11734);
or U18285 (N_18285,N_10024,N_14774);
nor U18286 (N_18286,N_14345,N_12834);
nand U18287 (N_18287,N_10811,N_11538);
or U18288 (N_18288,N_10650,N_11111);
nor U18289 (N_18289,N_11290,N_11145);
and U18290 (N_18290,N_13092,N_12776);
nor U18291 (N_18291,N_11631,N_11473);
and U18292 (N_18292,N_12489,N_12687);
nor U18293 (N_18293,N_13448,N_12307);
or U18294 (N_18294,N_13312,N_10144);
or U18295 (N_18295,N_11049,N_10558);
and U18296 (N_18296,N_13102,N_14650);
and U18297 (N_18297,N_10784,N_10404);
nor U18298 (N_18298,N_10893,N_13897);
and U18299 (N_18299,N_13079,N_10212);
nand U18300 (N_18300,N_13218,N_12542);
nor U18301 (N_18301,N_13852,N_12250);
and U18302 (N_18302,N_12887,N_12956);
or U18303 (N_18303,N_14392,N_11150);
nor U18304 (N_18304,N_14199,N_10501);
nor U18305 (N_18305,N_12385,N_10582);
xor U18306 (N_18306,N_12330,N_10200);
and U18307 (N_18307,N_14879,N_10466);
or U18308 (N_18308,N_14296,N_10552);
and U18309 (N_18309,N_10603,N_11960);
nor U18310 (N_18310,N_10949,N_13580);
xnor U18311 (N_18311,N_13749,N_13986);
and U18312 (N_18312,N_13146,N_12337);
and U18313 (N_18313,N_12567,N_14122);
and U18314 (N_18314,N_13338,N_12674);
nand U18315 (N_18315,N_14636,N_11985);
xor U18316 (N_18316,N_11413,N_10043);
nor U18317 (N_18317,N_13288,N_13128);
nand U18318 (N_18318,N_14841,N_14363);
nand U18319 (N_18319,N_14768,N_14441);
or U18320 (N_18320,N_11250,N_10295);
nor U18321 (N_18321,N_12998,N_13335);
xnor U18322 (N_18322,N_13030,N_13802);
xnor U18323 (N_18323,N_10132,N_13622);
nand U18324 (N_18324,N_10652,N_10334);
nor U18325 (N_18325,N_10398,N_10144);
and U18326 (N_18326,N_13874,N_14829);
nor U18327 (N_18327,N_13074,N_14484);
or U18328 (N_18328,N_12263,N_14016);
nor U18329 (N_18329,N_11317,N_10521);
nand U18330 (N_18330,N_14701,N_14714);
or U18331 (N_18331,N_14241,N_13375);
and U18332 (N_18332,N_10675,N_11736);
nor U18333 (N_18333,N_12426,N_11182);
nor U18334 (N_18334,N_12049,N_11143);
nand U18335 (N_18335,N_12659,N_11847);
or U18336 (N_18336,N_11940,N_12575);
nand U18337 (N_18337,N_13057,N_11866);
nor U18338 (N_18338,N_14011,N_12257);
nor U18339 (N_18339,N_12895,N_10944);
nor U18340 (N_18340,N_11660,N_14258);
xnor U18341 (N_18341,N_12520,N_13042);
nand U18342 (N_18342,N_13527,N_14664);
or U18343 (N_18343,N_14811,N_13347);
and U18344 (N_18344,N_13291,N_13461);
and U18345 (N_18345,N_12096,N_10377);
or U18346 (N_18346,N_13547,N_14832);
or U18347 (N_18347,N_12450,N_11190);
nand U18348 (N_18348,N_10347,N_11334);
or U18349 (N_18349,N_14083,N_11118);
nand U18350 (N_18350,N_11165,N_13468);
nand U18351 (N_18351,N_12932,N_11909);
and U18352 (N_18352,N_10881,N_12074);
nand U18353 (N_18353,N_11448,N_14076);
nand U18354 (N_18354,N_10861,N_12144);
nand U18355 (N_18355,N_14924,N_13070);
or U18356 (N_18356,N_11252,N_10888);
nand U18357 (N_18357,N_12967,N_14146);
nand U18358 (N_18358,N_11491,N_13235);
xnor U18359 (N_18359,N_12667,N_12555);
nand U18360 (N_18360,N_12788,N_14382);
xnor U18361 (N_18361,N_14632,N_10493);
or U18362 (N_18362,N_12220,N_14251);
nand U18363 (N_18363,N_13669,N_11995);
or U18364 (N_18364,N_12580,N_10470);
or U18365 (N_18365,N_12034,N_10393);
or U18366 (N_18366,N_12661,N_14719);
or U18367 (N_18367,N_12022,N_10028);
and U18368 (N_18368,N_12664,N_13086);
nand U18369 (N_18369,N_14581,N_11186);
nand U18370 (N_18370,N_10191,N_12714);
or U18371 (N_18371,N_13938,N_11935);
nand U18372 (N_18372,N_14599,N_11800);
nand U18373 (N_18373,N_10044,N_13383);
and U18374 (N_18374,N_12438,N_14506);
xor U18375 (N_18375,N_11064,N_13581);
nand U18376 (N_18376,N_13956,N_14109);
nor U18377 (N_18377,N_12127,N_10922);
xnor U18378 (N_18378,N_10032,N_13886);
and U18379 (N_18379,N_11796,N_14903);
or U18380 (N_18380,N_14679,N_11757);
or U18381 (N_18381,N_11026,N_12884);
or U18382 (N_18382,N_10393,N_11288);
or U18383 (N_18383,N_11563,N_14210);
or U18384 (N_18384,N_13809,N_13586);
and U18385 (N_18385,N_11038,N_13644);
nand U18386 (N_18386,N_14044,N_10315);
nand U18387 (N_18387,N_10865,N_14249);
and U18388 (N_18388,N_13433,N_10221);
or U18389 (N_18389,N_12555,N_11348);
or U18390 (N_18390,N_11701,N_12551);
nor U18391 (N_18391,N_12045,N_11677);
or U18392 (N_18392,N_12091,N_13661);
or U18393 (N_18393,N_11451,N_11780);
nand U18394 (N_18394,N_13949,N_11370);
and U18395 (N_18395,N_11651,N_11822);
nand U18396 (N_18396,N_14282,N_11316);
nand U18397 (N_18397,N_14302,N_10961);
xor U18398 (N_18398,N_14451,N_12400);
or U18399 (N_18399,N_11892,N_10876);
xor U18400 (N_18400,N_11977,N_14284);
nand U18401 (N_18401,N_13934,N_14531);
nor U18402 (N_18402,N_14261,N_14027);
nand U18403 (N_18403,N_13534,N_10894);
nand U18404 (N_18404,N_12316,N_12680);
nor U18405 (N_18405,N_14853,N_11523);
nor U18406 (N_18406,N_11300,N_11770);
and U18407 (N_18407,N_11279,N_12507);
xor U18408 (N_18408,N_10524,N_13607);
or U18409 (N_18409,N_13063,N_14001);
and U18410 (N_18410,N_10669,N_13968);
nand U18411 (N_18411,N_13052,N_13864);
and U18412 (N_18412,N_12403,N_11524);
nor U18413 (N_18413,N_11695,N_14632);
or U18414 (N_18414,N_11471,N_11522);
xor U18415 (N_18415,N_13272,N_14640);
nand U18416 (N_18416,N_11906,N_12978);
xnor U18417 (N_18417,N_10983,N_13788);
nand U18418 (N_18418,N_13964,N_14957);
nand U18419 (N_18419,N_11344,N_12330);
or U18420 (N_18420,N_11947,N_13197);
or U18421 (N_18421,N_12203,N_14535);
nor U18422 (N_18422,N_11450,N_10429);
or U18423 (N_18423,N_12084,N_11776);
nor U18424 (N_18424,N_10595,N_13859);
nor U18425 (N_18425,N_13500,N_14755);
and U18426 (N_18426,N_12005,N_12080);
nand U18427 (N_18427,N_13726,N_14947);
or U18428 (N_18428,N_14445,N_11621);
and U18429 (N_18429,N_14759,N_14832);
nand U18430 (N_18430,N_13012,N_11531);
nor U18431 (N_18431,N_10586,N_10416);
and U18432 (N_18432,N_14594,N_14456);
and U18433 (N_18433,N_13648,N_13429);
and U18434 (N_18434,N_12488,N_10121);
or U18435 (N_18435,N_14516,N_10558);
or U18436 (N_18436,N_11917,N_11856);
or U18437 (N_18437,N_14639,N_13353);
and U18438 (N_18438,N_10407,N_13489);
nor U18439 (N_18439,N_11658,N_11220);
xor U18440 (N_18440,N_10661,N_13364);
nand U18441 (N_18441,N_12010,N_14384);
xor U18442 (N_18442,N_11442,N_10579);
or U18443 (N_18443,N_12097,N_13545);
xnor U18444 (N_18444,N_10545,N_11024);
nand U18445 (N_18445,N_14819,N_14850);
nand U18446 (N_18446,N_11191,N_11248);
nor U18447 (N_18447,N_13347,N_12711);
and U18448 (N_18448,N_14574,N_10569);
xnor U18449 (N_18449,N_11624,N_11507);
or U18450 (N_18450,N_10424,N_11783);
or U18451 (N_18451,N_11981,N_13699);
and U18452 (N_18452,N_14873,N_11319);
or U18453 (N_18453,N_12831,N_10610);
nand U18454 (N_18454,N_12936,N_11490);
nand U18455 (N_18455,N_13603,N_14709);
nor U18456 (N_18456,N_13481,N_12932);
and U18457 (N_18457,N_14689,N_12263);
nand U18458 (N_18458,N_10752,N_11031);
or U18459 (N_18459,N_10985,N_10229);
and U18460 (N_18460,N_12535,N_11307);
and U18461 (N_18461,N_13785,N_13039);
nand U18462 (N_18462,N_10268,N_13925);
nor U18463 (N_18463,N_12267,N_12321);
and U18464 (N_18464,N_11241,N_14778);
nand U18465 (N_18465,N_10613,N_11209);
and U18466 (N_18466,N_12568,N_13880);
and U18467 (N_18467,N_11492,N_12979);
xnor U18468 (N_18468,N_10329,N_12572);
and U18469 (N_18469,N_11520,N_13781);
nor U18470 (N_18470,N_11723,N_11690);
nor U18471 (N_18471,N_11254,N_14308);
and U18472 (N_18472,N_11332,N_13197);
or U18473 (N_18473,N_13359,N_11800);
nor U18474 (N_18474,N_11922,N_10838);
nand U18475 (N_18475,N_10222,N_14083);
nand U18476 (N_18476,N_13626,N_11697);
nand U18477 (N_18477,N_12223,N_14048);
nor U18478 (N_18478,N_10390,N_11253);
nor U18479 (N_18479,N_10041,N_14232);
and U18480 (N_18480,N_14649,N_12736);
or U18481 (N_18481,N_12384,N_12626);
nor U18482 (N_18482,N_10360,N_14840);
nand U18483 (N_18483,N_12874,N_11858);
nand U18484 (N_18484,N_13903,N_14633);
or U18485 (N_18485,N_12737,N_14415);
or U18486 (N_18486,N_11079,N_14413);
or U18487 (N_18487,N_14194,N_11314);
and U18488 (N_18488,N_13949,N_11559);
nand U18489 (N_18489,N_10145,N_10455);
and U18490 (N_18490,N_14010,N_10933);
or U18491 (N_18491,N_11819,N_14322);
nand U18492 (N_18492,N_11855,N_12441);
or U18493 (N_18493,N_13471,N_12769);
nand U18494 (N_18494,N_10728,N_14353);
nor U18495 (N_18495,N_14068,N_12458);
nand U18496 (N_18496,N_12473,N_14723);
xnor U18497 (N_18497,N_13601,N_11862);
nand U18498 (N_18498,N_10047,N_12038);
or U18499 (N_18499,N_12849,N_13333);
xor U18500 (N_18500,N_10038,N_11140);
nor U18501 (N_18501,N_14828,N_13213);
nor U18502 (N_18502,N_14453,N_11953);
and U18503 (N_18503,N_12095,N_11092);
nor U18504 (N_18504,N_14593,N_12679);
and U18505 (N_18505,N_13657,N_10778);
and U18506 (N_18506,N_11008,N_11595);
or U18507 (N_18507,N_10596,N_13656);
or U18508 (N_18508,N_13813,N_14167);
or U18509 (N_18509,N_10524,N_11324);
or U18510 (N_18510,N_10123,N_14324);
and U18511 (N_18511,N_10802,N_11858);
xnor U18512 (N_18512,N_10351,N_13563);
and U18513 (N_18513,N_12479,N_13251);
or U18514 (N_18514,N_10781,N_11975);
and U18515 (N_18515,N_14701,N_11386);
nand U18516 (N_18516,N_14084,N_14604);
nand U18517 (N_18517,N_13426,N_10107);
nand U18518 (N_18518,N_10602,N_14231);
or U18519 (N_18519,N_10084,N_14556);
nor U18520 (N_18520,N_14044,N_14031);
or U18521 (N_18521,N_11059,N_13247);
or U18522 (N_18522,N_10087,N_10942);
and U18523 (N_18523,N_11867,N_14240);
or U18524 (N_18524,N_10227,N_12415);
or U18525 (N_18525,N_12352,N_10393);
or U18526 (N_18526,N_10648,N_13183);
nand U18527 (N_18527,N_12448,N_14715);
nand U18528 (N_18528,N_12252,N_13641);
nor U18529 (N_18529,N_12572,N_14997);
and U18530 (N_18530,N_13121,N_12309);
and U18531 (N_18531,N_11904,N_11671);
nand U18532 (N_18532,N_14946,N_13729);
and U18533 (N_18533,N_11773,N_13288);
or U18534 (N_18534,N_11906,N_11330);
and U18535 (N_18535,N_10269,N_12307);
or U18536 (N_18536,N_13670,N_13637);
or U18537 (N_18537,N_10142,N_14222);
nor U18538 (N_18538,N_14273,N_14609);
nand U18539 (N_18539,N_14384,N_12189);
or U18540 (N_18540,N_11189,N_13610);
nand U18541 (N_18541,N_13503,N_13473);
nor U18542 (N_18542,N_13022,N_13636);
or U18543 (N_18543,N_12692,N_10419);
nand U18544 (N_18544,N_10487,N_11507);
or U18545 (N_18545,N_11418,N_10993);
or U18546 (N_18546,N_14528,N_13627);
nor U18547 (N_18547,N_10429,N_14940);
and U18548 (N_18548,N_12158,N_13739);
nor U18549 (N_18549,N_11850,N_14797);
or U18550 (N_18550,N_10288,N_14171);
xnor U18551 (N_18551,N_12603,N_11949);
xnor U18552 (N_18552,N_11783,N_14863);
nor U18553 (N_18553,N_14858,N_13477);
nor U18554 (N_18554,N_12209,N_10278);
or U18555 (N_18555,N_13955,N_14278);
nor U18556 (N_18556,N_13590,N_14362);
and U18557 (N_18557,N_13165,N_11544);
nand U18558 (N_18558,N_10526,N_10801);
and U18559 (N_18559,N_12197,N_14047);
xnor U18560 (N_18560,N_11575,N_13052);
xor U18561 (N_18561,N_14941,N_12106);
and U18562 (N_18562,N_11587,N_14034);
nand U18563 (N_18563,N_13276,N_11344);
nand U18564 (N_18564,N_12542,N_13837);
nor U18565 (N_18565,N_14733,N_12385);
nor U18566 (N_18566,N_12770,N_14666);
xor U18567 (N_18567,N_13829,N_13333);
and U18568 (N_18568,N_10239,N_11599);
nor U18569 (N_18569,N_13717,N_14568);
or U18570 (N_18570,N_13283,N_13106);
or U18571 (N_18571,N_13127,N_12155);
and U18572 (N_18572,N_14078,N_14264);
or U18573 (N_18573,N_14717,N_12655);
nor U18574 (N_18574,N_13525,N_13264);
and U18575 (N_18575,N_11089,N_13902);
nand U18576 (N_18576,N_14006,N_13954);
nor U18577 (N_18577,N_11264,N_14755);
and U18578 (N_18578,N_12344,N_14504);
and U18579 (N_18579,N_13517,N_12963);
or U18580 (N_18580,N_11408,N_14028);
nand U18581 (N_18581,N_12886,N_10825);
nor U18582 (N_18582,N_14107,N_12701);
nor U18583 (N_18583,N_11835,N_10292);
nor U18584 (N_18584,N_14980,N_12710);
nor U18585 (N_18585,N_13088,N_13015);
and U18586 (N_18586,N_13141,N_10665);
and U18587 (N_18587,N_11463,N_11591);
xnor U18588 (N_18588,N_11346,N_13376);
nor U18589 (N_18589,N_10627,N_11229);
nand U18590 (N_18590,N_13223,N_12559);
xor U18591 (N_18591,N_14783,N_11365);
or U18592 (N_18592,N_10169,N_12209);
and U18593 (N_18593,N_14947,N_10307);
nand U18594 (N_18594,N_14890,N_13313);
nor U18595 (N_18595,N_14178,N_14203);
nand U18596 (N_18596,N_13881,N_14434);
and U18597 (N_18597,N_12327,N_11775);
and U18598 (N_18598,N_10627,N_10163);
xnor U18599 (N_18599,N_12931,N_14900);
and U18600 (N_18600,N_14121,N_10727);
nand U18601 (N_18601,N_12197,N_11105);
and U18602 (N_18602,N_13917,N_14421);
nand U18603 (N_18603,N_12475,N_11841);
nor U18604 (N_18604,N_10489,N_13477);
nand U18605 (N_18605,N_11563,N_13099);
nand U18606 (N_18606,N_10262,N_11663);
and U18607 (N_18607,N_13506,N_14313);
and U18608 (N_18608,N_14727,N_14374);
and U18609 (N_18609,N_12598,N_13624);
and U18610 (N_18610,N_14365,N_12968);
nand U18611 (N_18611,N_14724,N_11932);
or U18612 (N_18612,N_10115,N_11941);
or U18613 (N_18613,N_12755,N_14053);
nand U18614 (N_18614,N_13718,N_10088);
nand U18615 (N_18615,N_11092,N_14788);
nor U18616 (N_18616,N_13314,N_13005);
nor U18617 (N_18617,N_13152,N_12215);
nand U18618 (N_18618,N_14900,N_13673);
nand U18619 (N_18619,N_11796,N_10455);
and U18620 (N_18620,N_10760,N_14273);
nor U18621 (N_18621,N_14273,N_10089);
nor U18622 (N_18622,N_11591,N_14966);
or U18623 (N_18623,N_10743,N_10521);
nor U18624 (N_18624,N_12594,N_12197);
or U18625 (N_18625,N_14370,N_13955);
nand U18626 (N_18626,N_10242,N_10438);
nand U18627 (N_18627,N_13402,N_11278);
or U18628 (N_18628,N_12308,N_10207);
nor U18629 (N_18629,N_11033,N_14541);
nand U18630 (N_18630,N_12440,N_14060);
or U18631 (N_18631,N_14875,N_11365);
or U18632 (N_18632,N_11615,N_11492);
nor U18633 (N_18633,N_13159,N_12130);
nand U18634 (N_18634,N_11184,N_13580);
nor U18635 (N_18635,N_11359,N_11754);
or U18636 (N_18636,N_13088,N_14936);
and U18637 (N_18637,N_10356,N_11654);
nand U18638 (N_18638,N_11740,N_14662);
and U18639 (N_18639,N_12116,N_13720);
and U18640 (N_18640,N_13381,N_12090);
nor U18641 (N_18641,N_11526,N_11978);
and U18642 (N_18642,N_10787,N_11896);
nand U18643 (N_18643,N_12808,N_14074);
and U18644 (N_18644,N_10402,N_12552);
or U18645 (N_18645,N_12462,N_14526);
and U18646 (N_18646,N_13972,N_14455);
nor U18647 (N_18647,N_13537,N_10396);
xor U18648 (N_18648,N_13508,N_10346);
nor U18649 (N_18649,N_11942,N_13411);
nand U18650 (N_18650,N_14220,N_10645);
xor U18651 (N_18651,N_14610,N_11408);
nand U18652 (N_18652,N_13852,N_14725);
or U18653 (N_18653,N_13144,N_10032);
and U18654 (N_18654,N_13492,N_11120);
nor U18655 (N_18655,N_11472,N_12805);
or U18656 (N_18656,N_14354,N_13977);
nor U18657 (N_18657,N_10324,N_12333);
nor U18658 (N_18658,N_12488,N_11620);
nand U18659 (N_18659,N_10418,N_13027);
or U18660 (N_18660,N_14694,N_12274);
xor U18661 (N_18661,N_12889,N_11955);
nor U18662 (N_18662,N_14102,N_11025);
nor U18663 (N_18663,N_10754,N_13250);
and U18664 (N_18664,N_13608,N_10561);
nand U18665 (N_18665,N_13996,N_11845);
nor U18666 (N_18666,N_12094,N_11818);
and U18667 (N_18667,N_13055,N_11734);
or U18668 (N_18668,N_12487,N_12548);
nand U18669 (N_18669,N_13908,N_10818);
nor U18670 (N_18670,N_11207,N_12633);
nor U18671 (N_18671,N_12234,N_10909);
and U18672 (N_18672,N_11168,N_12285);
xnor U18673 (N_18673,N_13889,N_14575);
nand U18674 (N_18674,N_14290,N_10711);
and U18675 (N_18675,N_10426,N_14424);
nand U18676 (N_18676,N_12320,N_11688);
nand U18677 (N_18677,N_11846,N_12444);
and U18678 (N_18678,N_10982,N_11867);
nor U18679 (N_18679,N_11477,N_11616);
and U18680 (N_18680,N_11024,N_12533);
or U18681 (N_18681,N_13653,N_12703);
xor U18682 (N_18682,N_10579,N_13037);
nand U18683 (N_18683,N_10577,N_13614);
or U18684 (N_18684,N_14476,N_14545);
and U18685 (N_18685,N_12189,N_12858);
and U18686 (N_18686,N_13309,N_12742);
nor U18687 (N_18687,N_14015,N_10935);
nand U18688 (N_18688,N_13527,N_11765);
or U18689 (N_18689,N_14310,N_12517);
nand U18690 (N_18690,N_14308,N_10729);
nor U18691 (N_18691,N_10243,N_10814);
or U18692 (N_18692,N_10338,N_13758);
or U18693 (N_18693,N_14409,N_12391);
nor U18694 (N_18694,N_14954,N_14415);
nand U18695 (N_18695,N_10216,N_11347);
nand U18696 (N_18696,N_13949,N_10451);
nor U18697 (N_18697,N_11228,N_12618);
and U18698 (N_18698,N_11812,N_12565);
nand U18699 (N_18699,N_12095,N_12590);
and U18700 (N_18700,N_14084,N_13950);
and U18701 (N_18701,N_13306,N_14787);
nand U18702 (N_18702,N_11517,N_12502);
and U18703 (N_18703,N_12864,N_10446);
nand U18704 (N_18704,N_14903,N_10659);
nand U18705 (N_18705,N_12474,N_10095);
or U18706 (N_18706,N_10052,N_13496);
and U18707 (N_18707,N_11756,N_12228);
nor U18708 (N_18708,N_14379,N_12346);
nor U18709 (N_18709,N_10962,N_10005);
and U18710 (N_18710,N_14141,N_10135);
and U18711 (N_18711,N_14446,N_10161);
or U18712 (N_18712,N_12317,N_12592);
and U18713 (N_18713,N_10105,N_13457);
nor U18714 (N_18714,N_14692,N_12626);
nand U18715 (N_18715,N_10380,N_10644);
or U18716 (N_18716,N_14200,N_11747);
or U18717 (N_18717,N_11197,N_14626);
and U18718 (N_18718,N_10912,N_10145);
nand U18719 (N_18719,N_13279,N_10670);
nor U18720 (N_18720,N_12968,N_10423);
and U18721 (N_18721,N_13604,N_14157);
or U18722 (N_18722,N_11402,N_10755);
xor U18723 (N_18723,N_14780,N_12409);
xor U18724 (N_18724,N_12785,N_12074);
and U18725 (N_18725,N_10937,N_14722);
nor U18726 (N_18726,N_13329,N_12218);
nand U18727 (N_18727,N_14950,N_10597);
or U18728 (N_18728,N_12441,N_10629);
and U18729 (N_18729,N_11860,N_10184);
nor U18730 (N_18730,N_10741,N_12721);
or U18731 (N_18731,N_11619,N_11755);
nand U18732 (N_18732,N_13473,N_14881);
xor U18733 (N_18733,N_11376,N_12987);
nor U18734 (N_18734,N_10259,N_11325);
nor U18735 (N_18735,N_12252,N_12449);
nor U18736 (N_18736,N_11817,N_11107);
or U18737 (N_18737,N_11126,N_10471);
or U18738 (N_18738,N_12452,N_12109);
and U18739 (N_18739,N_11675,N_11881);
nor U18740 (N_18740,N_10433,N_12272);
nor U18741 (N_18741,N_14834,N_13605);
and U18742 (N_18742,N_12357,N_11712);
and U18743 (N_18743,N_14646,N_11543);
nand U18744 (N_18744,N_13622,N_13568);
or U18745 (N_18745,N_10629,N_13109);
and U18746 (N_18746,N_12545,N_10663);
xnor U18747 (N_18747,N_12331,N_10548);
and U18748 (N_18748,N_12277,N_10270);
nor U18749 (N_18749,N_11416,N_10803);
and U18750 (N_18750,N_11228,N_14350);
or U18751 (N_18751,N_11149,N_12856);
or U18752 (N_18752,N_12085,N_14414);
or U18753 (N_18753,N_10809,N_13108);
or U18754 (N_18754,N_13665,N_12208);
nand U18755 (N_18755,N_12030,N_13699);
nor U18756 (N_18756,N_12390,N_13663);
or U18757 (N_18757,N_14148,N_10432);
or U18758 (N_18758,N_12673,N_12607);
nand U18759 (N_18759,N_14139,N_12332);
xnor U18760 (N_18760,N_14474,N_10267);
or U18761 (N_18761,N_10257,N_11868);
nand U18762 (N_18762,N_10350,N_11250);
and U18763 (N_18763,N_14765,N_14455);
and U18764 (N_18764,N_10282,N_10854);
nand U18765 (N_18765,N_10627,N_14137);
xnor U18766 (N_18766,N_14754,N_13663);
and U18767 (N_18767,N_12516,N_12660);
xnor U18768 (N_18768,N_11870,N_10714);
or U18769 (N_18769,N_11212,N_12604);
nor U18770 (N_18770,N_10174,N_11568);
nand U18771 (N_18771,N_11170,N_12284);
nor U18772 (N_18772,N_11261,N_12545);
nand U18773 (N_18773,N_13900,N_12903);
or U18774 (N_18774,N_13224,N_13159);
xnor U18775 (N_18775,N_13411,N_14075);
nor U18776 (N_18776,N_14392,N_12680);
and U18777 (N_18777,N_11373,N_12564);
nand U18778 (N_18778,N_12259,N_13733);
nand U18779 (N_18779,N_13937,N_11320);
xnor U18780 (N_18780,N_14308,N_13075);
or U18781 (N_18781,N_12461,N_11323);
nor U18782 (N_18782,N_12995,N_12688);
and U18783 (N_18783,N_10324,N_11683);
nand U18784 (N_18784,N_10398,N_14346);
and U18785 (N_18785,N_10305,N_10291);
and U18786 (N_18786,N_10576,N_12619);
xnor U18787 (N_18787,N_12397,N_11909);
nand U18788 (N_18788,N_10693,N_12096);
or U18789 (N_18789,N_10172,N_12900);
and U18790 (N_18790,N_10437,N_11090);
nand U18791 (N_18791,N_12144,N_12005);
nand U18792 (N_18792,N_12652,N_12141);
nor U18793 (N_18793,N_12583,N_13228);
and U18794 (N_18794,N_14984,N_10148);
or U18795 (N_18795,N_11071,N_13684);
or U18796 (N_18796,N_12798,N_13777);
nand U18797 (N_18797,N_12586,N_10344);
nor U18798 (N_18798,N_13465,N_11672);
xnor U18799 (N_18799,N_12688,N_10269);
or U18800 (N_18800,N_13315,N_12535);
and U18801 (N_18801,N_11494,N_12357);
or U18802 (N_18802,N_12806,N_13220);
xnor U18803 (N_18803,N_13218,N_14063);
and U18804 (N_18804,N_10214,N_13389);
nor U18805 (N_18805,N_13727,N_14643);
nor U18806 (N_18806,N_10880,N_14468);
nor U18807 (N_18807,N_10939,N_10611);
or U18808 (N_18808,N_13064,N_12991);
and U18809 (N_18809,N_14970,N_11589);
nand U18810 (N_18810,N_12964,N_11428);
nand U18811 (N_18811,N_13012,N_13647);
or U18812 (N_18812,N_12428,N_13629);
or U18813 (N_18813,N_10780,N_11865);
nor U18814 (N_18814,N_12530,N_11041);
and U18815 (N_18815,N_11966,N_13649);
and U18816 (N_18816,N_10502,N_11169);
nand U18817 (N_18817,N_11072,N_11732);
nand U18818 (N_18818,N_12135,N_10812);
or U18819 (N_18819,N_13651,N_11363);
nor U18820 (N_18820,N_13053,N_12709);
and U18821 (N_18821,N_14767,N_11637);
and U18822 (N_18822,N_13783,N_12826);
nor U18823 (N_18823,N_14123,N_10860);
nand U18824 (N_18824,N_14220,N_13420);
nor U18825 (N_18825,N_11023,N_14738);
or U18826 (N_18826,N_10275,N_12333);
or U18827 (N_18827,N_13540,N_13956);
or U18828 (N_18828,N_11697,N_14247);
and U18829 (N_18829,N_13376,N_13552);
xor U18830 (N_18830,N_11534,N_14915);
nor U18831 (N_18831,N_13272,N_14487);
or U18832 (N_18832,N_14488,N_13481);
and U18833 (N_18833,N_11358,N_12531);
or U18834 (N_18834,N_12623,N_10253);
xnor U18835 (N_18835,N_14646,N_11036);
and U18836 (N_18836,N_14762,N_12381);
nor U18837 (N_18837,N_14375,N_10693);
and U18838 (N_18838,N_11472,N_13544);
nand U18839 (N_18839,N_10916,N_14130);
nor U18840 (N_18840,N_14032,N_12610);
or U18841 (N_18841,N_10102,N_12770);
nand U18842 (N_18842,N_11261,N_12784);
nor U18843 (N_18843,N_13448,N_13868);
and U18844 (N_18844,N_12619,N_10645);
or U18845 (N_18845,N_11986,N_10053);
or U18846 (N_18846,N_12051,N_10746);
or U18847 (N_18847,N_10848,N_13378);
and U18848 (N_18848,N_14108,N_12344);
nand U18849 (N_18849,N_12683,N_10207);
and U18850 (N_18850,N_11693,N_11240);
nor U18851 (N_18851,N_14297,N_14928);
and U18852 (N_18852,N_13362,N_14976);
or U18853 (N_18853,N_14609,N_14480);
nor U18854 (N_18854,N_10919,N_14335);
and U18855 (N_18855,N_10255,N_12753);
nor U18856 (N_18856,N_12421,N_13873);
and U18857 (N_18857,N_14985,N_13146);
or U18858 (N_18858,N_11624,N_14406);
or U18859 (N_18859,N_11386,N_11965);
xor U18860 (N_18860,N_11928,N_13946);
or U18861 (N_18861,N_12200,N_10855);
nand U18862 (N_18862,N_13087,N_10029);
nor U18863 (N_18863,N_10633,N_10109);
and U18864 (N_18864,N_11738,N_12965);
and U18865 (N_18865,N_11081,N_11919);
xor U18866 (N_18866,N_12226,N_14274);
nand U18867 (N_18867,N_13141,N_12300);
nor U18868 (N_18868,N_11915,N_11746);
nand U18869 (N_18869,N_14408,N_12606);
nor U18870 (N_18870,N_10901,N_10191);
or U18871 (N_18871,N_13302,N_13101);
nor U18872 (N_18872,N_14130,N_11925);
xor U18873 (N_18873,N_12466,N_13793);
nand U18874 (N_18874,N_11400,N_11738);
or U18875 (N_18875,N_13954,N_14622);
nor U18876 (N_18876,N_10184,N_13939);
or U18877 (N_18877,N_13140,N_14994);
or U18878 (N_18878,N_14109,N_12010);
nor U18879 (N_18879,N_12362,N_12788);
and U18880 (N_18880,N_11143,N_13555);
xnor U18881 (N_18881,N_12272,N_14752);
or U18882 (N_18882,N_14539,N_14725);
nand U18883 (N_18883,N_14672,N_12554);
and U18884 (N_18884,N_13828,N_14458);
nand U18885 (N_18885,N_11411,N_10909);
and U18886 (N_18886,N_13086,N_14535);
or U18887 (N_18887,N_12491,N_10547);
and U18888 (N_18888,N_13307,N_14639);
nor U18889 (N_18889,N_10763,N_14929);
nor U18890 (N_18890,N_13388,N_12551);
and U18891 (N_18891,N_11182,N_11504);
or U18892 (N_18892,N_11588,N_13785);
xnor U18893 (N_18893,N_13938,N_11004);
nand U18894 (N_18894,N_13853,N_12555);
nor U18895 (N_18895,N_14852,N_11171);
and U18896 (N_18896,N_14358,N_11273);
nand U18897 (N_18897,N_14479,N_14846);
and U18898 (N_18898,N_14557,N_13745);
or U18899 (N_18899,N_14111,N_12897);
nand U18900 (N_18900,N_14031,N_14437);
nand U18901 (N_18901,N_12014,N_12759);
nor U18902 (N_18902,N_10627,N_11539);
nand U18903 (N_18903,N_11707,N_11943);
nand U18904 (N_18904,N_10974,N_10802);
and U18905 (N_18905,N_10372,N_13553);
nand U18906 (N_18906,N_11452,N_11665);
or U18907 (N_18907,N_11518,N_10195);
or U18908 (N_18908,N_10347,N_14044);
or U18909 (N_18909,N_13379,N_10257);
nand U18910 (N_18910,N_12706,N_13511);
nand U18911 (N_18911,N_13116,N_10234);
xnor U18912 (N_18912,N_12594,N_13747);
and U18913 (N_18913,N_11650,N_10949);
or U18914 (N_18914,N_11470,N_12446);
and U18915 (N_18915,N_10621,N_13625);
or U18916 (N_18916,N_12080,N_14845);
nand U18917 (N_18917,N_13227,N_14734);
and U18918 (N_18918,N_11408,N_12196);
nor U18919 (N_18919,N_11038,N_11531);
and U18920 (N_18920,N_10020,N_11701);
and U18921 (N_18921,N_10830,N_14696);
nor U18922 (N_18922,N_11780,N_11231);
nor U18923 (N_18923,N_12574,N_13457);
or U18924 (N_18924,N_13511,N_11289);
or U18925 (N_18925,N_13900,N_10310);
nand U18926 (N_18926,N_12579,N_13550);
or U18927 (N_18927,N_14787,N_12526);
xnor U18928 (N_18928,N_10628,N_13631);
nand U18929 (N_18929,N_12419,N_11243);
nor U18930 (N_18930,N_10802,N_11190);
nand U18931 (N_18931,N_13927,N_13456);
and U18932 (N_18932,N_10341,N_11714);
nor U18933 (N_18933,N_13712,N_10999);
xnor U18934 (N_18934,N_12989,N_14714);
and U18935 (N_18935,N_14311,N_14885);
nand U18936 (N_18936,N_11037,N_11916);
nor U18937 (N_18937,N_10744,N_10265);
nand U18938 (N_18938,N_11566,N_11801);
and U18939 (N_18939,N_11056,N_10357);
nand U18940 (N_18940,N_13156,N_13374);
nand U18941 (N_18941,N_12093,N_14642);
nand U18942 (N_18942,N_13668,N_14211);
nor U18943 (N_18943,N_14912,N_10749);
nor U18944 (N_18944,N_13173,N_11991);
nand U18945 (N_18945,N_11168,N_13146);
or U18946 (N_18946,N_13692,N_11271);
nor U18947 (N_18947,N_10181,N_12292);
xor U18948 (N_18948,N_10629,N_13451);
nor U18949 (N_18949,N_12431,N_10321);
and U18950 (N_18950,N_12862,N_11005);
and U18951 (N_18951,N_13775,N_11639);
and U18952 (N_18952,N_10052,N_12112);
nand U18953 (N_18953,N_10609,N_11810);
and U18954 (N_18954,N_12506,N_13027);
nand U18955 (N_18955,N_12357,N_10278);
or U18956 (N_18956,N_10311,N_10746);
nand U18957 (N_18957,N_13199,N_12138);
nor U18958 (N_18958,N_13936,N_12416);
nand U18959 (N_18959,N_14392,N_11799);
nand U18960 (N_18960,N_12497,N_10860);
and U18961 (N_18961,N_14270,N_13792);
nor U18962 (N_18962,N_11064,N_13634);
nor U18963 (N_18963,N_12827,N_13430);
or U18964 (N_18964,N_13435,N_14288);
and U18965 (N_18965,N_12663,N_12939);
nand U18966 (N_18966,N_11277,N_14523);
and U18967 (N_18967,N_11604,N_11801);
and U18968 (N_18968,N_11456,N_13225);
or U18969 (N_18969,N_10003,N_10486);
or U18970 (N_18970,N_11762,N_10899);
nor U18971 (N_18971,N_12862,N_11693);
and U18972 (N_18972,N_11732,N_11556);
nand U18973 (N_18973,N_13992,N_10325);
xnor U18974 (N_18974,N_12655,N_14323);
xor U18975 (N_18975,N_10081,N_13926);
and U18976 (N_18976,N_12749,N_13439);
and U18977 (N_18977,N_13825,N_12961);
and U18978 (N_18978,N_12971,N_11365);
nor U18979 (N_18979,N_10344,N_10456);
and U18980 (N_18980,N_10652,N_11734);
nand U18981 (N_18981,N_14974,N_13043);
nand U18982 (N_18982,N_10275,N_11057);
nor U18983 (N_18983,N_14274,N_13654);
nor U18984 (N_18984,N_14724,N_11975);
nand U18985 (N_18985,N_14234,N_14408);
and U18986 (N_18986,N_14070,N_10024);
and U18987 (N_18987,N_11941,N_13250);
and U18988 (N_18988,N_11334,N_14094);
nand U18989 (N_18989,N_13494,N_10977);
xnor U18990 (N_18990,N_10737,N_10030);
nor U18991 (N_18991,N_11902,N_14811);
or U18992 (N_18992,N_12479,N_10811);
and U18993 (N_18993,N_12417,N_14192);
nor U18994 (N_18994,N_10086,N_11568);
nor U18995 (N_18995,N_14178,N_12667);
and U18996 (N_18996,N_14753,N_11308);
nand U18997 (N_18997,N_14223,N_12400);
xor U18998 (N_18998,N_13452,N_11903);
or U18999 (N_18999,N_11683,N_13191);
nor U19000 (N_19000,N_14839,N_14027);
xor U19001 (N_19001,N_13030,N_11466);
xnor U19002 (N_19002,N_12832,N_12410);
and U19003 (N_19003,N_12000,N_13070);
or U19004 (N_19004,N_12878,N_13031);
nand U19005 (N_19005,N_11473,N_13126);
or U19006 (N_19006,N_13175,N_12693);
nor U19007 (N_19007,N_12714,N_11392);
nor U19008 (N_19008,N_14631,N_10909);
and U19009 (N_19009,N_11173,N_11347);
xnor U19010 (N_19010,N_14621,N_11911);
nor U19011 (N_19011,N_11767,N_11823);
nor U19012 (N_19012,N_11400,N_13462);
nor U19013 (N_19013,N_11687,N_10121);
and U19014 (N_19014,N_11603,N_13706);
nand U19015 (N_19015,N_12653,N_11261);
nand U19016 (N_19016,N_14672,N_10402);
xor U19017 (N_19017,N_10772,N_14800);
nor U19018 (N_19018,N_14113,N_11674);
and U19019 (N_19019,N_11645,N_12227);
or U19020 (N_19020,N_12658,N_14800);
nand U19021 (N_19021,N_10817,N_14109);
or U19022 (N_19022,N_11103,N_12089);
and U19023 (N_19023,N_10745,N_11563);
and U19024 (N_19024,N_13646,N_13936);
and U19025 (N_19025,N_13104,N_12450);
nor U19026 (N_19026,N_14874,N_12379);
or U19027 (N_19027,N_10865,N_14716);
nand U19028 (N_19028,N_10322,N_11838);
and U19029 (N_19029,N_13428,N_12893);
and U19030 (N_19030,N_11297,N_12826);
nand U19031 (N_19031,N_12618,N_12693);
or U19032 (N_19032,N_11014,N_13917);
or U19033 (N_19033,N_13870,N_13135);
xnor U19034 (N_19034,N_12011,N_11493);
or U19035 (N_19035,N_13366,N_11312);
nor U19036 (N_19036,N_14371,N_10745);
or U19037 (N_19037,N_13234,N_11555);
or U19038 (N_19038,N_10915,N_11595);
nand U19039 (N_19039,N_12432,N_11508);
nand U19040 (N_19040,N_12636,N_14670);
nor U19041 (N_19041,N_10966,N_13156);
and U19042 (N_19042,N_14050,N_14624);
or U19043 (N_19043,N_12538,N_12344);
and U19044 (N_19044,N_10063,N_12639);
nand U19045 (N_19045,N_12124,N_11065);
nand U19046 (N_19046,N_11614,N_13242);
nor U19047 (N_19047,N_12131,N_12909);
or U19048 (N_19048,N_11128,N_12702);
or U19049 (N_19049,N_11194,N_13141);
nand U19050 (N_19050,N_10534,N_11772);
nor U19051 (N_19051,N_12341,N_12509);
or U19052 (N_19052,N_10558,N_12881);
nor U19053 (N_19053,N_11301,N_11031);
nor U19054 (N_19054,N_12491,N_11394);
nor U19055 (N_19055,N_11275,N_12705);
or U19056 (N_19056,N_14345,N_11951);
nand U19057 (N_19057,N_10042,N_14307);
or U19058 (N_19058,N_12147,N_11011);
or U19059 (N_19059,N_12757,N_11186);
and U19060 (N_19060,N_14206,N_10618);
nor U19061 (N_19061,N_12165,N_12590);
or U19062 (N_19062,N_11639,N_13015);
and U19063 (N_19063,N_14061,N_11081);
or U19064 (N_19064,N_11894,N_12719);
and U19065 (N_19065,N_11429,N_12097);
or U19066 (N_19066,N_14118,N_10043);
and U19067 (N_19067,N_14134,N_10851);
or U19068 (N_19068,N_14473,N_10012);
xnor U19069 (N_19069,N_11369,N_12986);
nor U19070 (N_19070,N_14140,N_11811);
nand U19071 (N_19071,N_12768,N_12675);
nand U19072 (N_19072,N_12617,N_14086);
nor U19073 (N_19073,N_12411,N_13185);
or U19074 (N_19074,N_12593,N_10366);
xor U19075 (N_19075,N_12101,N_11527);
xnor U19076 (N_19076,N_10140,N_14209);
xor U19077 (N_19077,N_12193,N_14345);
nand U19078 (N_19078,N_12388,N_13576);
xor U19079 (N_19079,N_14414,N_12186);
or U19080 (N_19080,N_10630,N_10323);
nand U19081 (N_19081,N_10762,N_14882);
or U19082 (N_19082,N_12995,N_11542);
nor U19083 (N_19083,N_13966,N_12664);
xnor U19084 (N_19084,N_11099,N_13306);
nand U19085 (N_19085,N_14663,N_12139);
nor U19086 (N_19086,N_13332,N_12153);
nand U19087 (N_19087,N_14670,N_11045);
or U19088 (N_19088,N_12004,N_14715);
and U19089 (N_19089,N_12011,N_12995);
nand U19090 (N_19090,N_13585,N_11240);
nor U19091 (N_19091,N_13479,N_14890);
xnor U19092 (N_19092,N_10396,N_11560);
nand U19093 (N_19093,N_10956,N_14152);
and U19094 (N_19094,N_10453,N_13289);
nor U19095 (N_19095,N_14706,N_11895);
and U19096 (N_19096,N_14466,N_13075);
nand U19097 (N_19097,N_14220,N_12222);
or U19098 (N_19098,N_11786,N_13010);
nand U19099 (N_19099,N_13991,N_10857);
nand U19100 (N_19100,N_13760,N_11821);
nand U19101 (N_19101,N_13090,N_10245);
or U19102 (N_19102,N_14905,N_10473);
nand U19103 (N_19103,N_10748,N_13008);
nand U19104 (N_19104,N_11440,N_13082);
nor U19105 (N_19105,N_13666,N_11771);
nor U19106 (N_19106,N_12923,N_14100);
xnor U19107 (N_19107,N_14005,N_12208);
and U19108 (N_19108,N_12901,N_13354);
and U19109 (N_19109,N_12192,N_11965);
and U19110 (N_19110,N_10869,N_12514);
and U19111 (N_19111,N_12805,N_12011);
and U19112 (N_19112,N_12383,N_10883);
xnor U19113 (N_19113,N_14026,N_14488);
nand U19114 (N_19114,N_11921,N_12817);
and U19115 (N_19115,N_10814,N_10764);
or U19116 (N_19116,N_10832,N_12927);
nor U19117 (N_19117,N_14554,N_11286);
nor U19118 (N_19118,N_13653,N_10206);
and U19119 (N_19119,N_10868,N_13857);
nor U19120 (N_19120,N_10639,N_13017);
nand U19121 (N_19121,N_13475,N_14200);
nand U19122 (N_19122,N_13033,N_14942);
and U19123 (N_19123,N_13574,N_14774);
or U19124 (N_19124,N_14265,N_10296);
and U19125 (N_19125,N_12421,N_12020);
or U19126 (N_19126,N_12577,N_13529);
or U19127 (N_19127,N_10279,N_14350);
and U19128 (N_19128,N_10883,N_14679);
xnor U19129 (N_19129,N_13515,N_10968);
or U19130 (N_19130,N_11512,N_10775);
xor U19131 (N_19131,N_11566,N_11843);
xor U19132 (N_19132,N_12294,N_11211);
nor U19133 (N_19133,N_13434,N_13025);
or U19134 (N_19134,N_12812,N_11343);
nand U19135 (N_19135,N_12764,N_11929);
xor U19136 (N_19136,N_13493,N_13963);
or U19137 (N_19137,N_14385,N_14650);
nand U19138 (N_19138,N_12054,N_10960);
nor U19139 (N_19139,N_12647,N_14984);
and U19140 (N_19140,N_11141,N_13251);
and U19141 (N_19141,N_10457,N_11743);
and U19142 (N_19142,N_11797,N_10860);
xor U19143 (N_19143,N_12762,N_13305);
or U19144 (N_19144,N_11875,N_10087);
nor U19145 (N_19145,N_14475,N_11846);
xnor U19146 (N_19146,N_14243,N_10243);
and U19147 (N_19147,N_13947,N_11726);
and U19148 (N_19148,N_14493,N_12703);
or U19149 (N_19149,N_13540,N_14909);
or U19150 (N_19150,N_14031,N_14630);
nand U19151 (N_19151,N_13829,N_12821);
nand U19152 (N_19152,N_11021,N_14406);
and U19153 (N_19153,N_10761,N_13588);
and U19154 (N_19154,N_13074,N_11319);
or U19155 (N_19155,N_10148,N_12469);
nand U19156 (N_19156,N_14768,N_14478);
nor U19157 (N_19157,N_13718,N_12607);
xor U19158 (N_19158,N_11986,N_13149);
nor U19159 (N_19159,N_10321,N_12811);
or U19160 (N_19160,N_13963,N_10670);
and U19161 (N_19161,N_12286,N_12570);
or U19162 (N_19162,N_11623,N_11414);
xor U19163 (N_19163,N_12750,N_13336);
or U19164 (N_19164,N_12428,N_12780);
nand U19165 (N_19165,N_13058,N_13764);
or U19166 (N_19166,N_12502,N_13777);
or U19167 (N_19167,N_12128,N_11146);
xor U19168 (N_19168,N_12305,N_13437);
and U19169 (N_19169,N_12494,N_12257);
nand U19170 (N_19170,N_14844,N_14569);
or U19171 (N_19171,N_14713,N_12134);
nand U19172 (N_19172,N_11944,N_13932);
nand U19173 (N_19173,N_12162,N_10385);
xnor U19174 (N_19174,N_12800,N_13689);
nor U19175 (N_19175,N_13764,N_11850);
nor U19176 (N_19176,N_10535,N_11667);
nand U19177 (N_19177,N_10182,N_13943);
nand U19178 (N_19178,N_10440,N_14134);
nand U19179 (N_19179,N_11156,N_12562);
nor U19180 (N_19180,N_13657,N_10783);
xor U19181 (N_19181,N_10494,N_11836);
nand U19182 (N_19182,N_14957,N_10151);
or U19183 (N_19183,N_13871,N_10598);
nand U19184 (N_19184,N_13373,N_10200);
or U19185 (N_19185,N_12723,N_12987);
nor U19186 (N_19186,N_11239,N_11169);
and U19187 (N_19187,N_14334,N_10221);
or U19188 (N_19188,N_14632,N_13626);
nand U19189 (N_19189,N_13945,N_11959);
or U19190 (N_19190,N_10806,N_13642);
and U19191 (N_19191,N_11301,N_11624);
and U19192 (N_19192,N_13878,N_10675);
and U19193 (N_19193,N_12437,N_10683);
nor U19194 (N_19194,N_11619,N_11502);
and U19195 (N_19195,N_12213,N_10229);
or U19196 (N_19196,N_12612,N_11902);
and U19197 (N_19197,N_13904,N_14938);
and U19198 (N_19198,N_11687,N_13729);
nor U19199 (N_19199,N_13570,N_10721);
or U19200 (N_19200,N_12218,N_12570);
xor U19201 (N_19201,N_12230,N_12476);
nor U19202 (N_19202,N_12279,N_12408);
nor U19203 (N_19203,N_10157,N_13243);
and U19204 (N_19204,N_14277,N_14615);
and U19205 (N_19205,N_13589,N_14519);
nor U19206 (N_19206,N_14399,N_14759);
nor U19207 (N_19207,N_14370,N_10370);
xor U19208 (N_19208,N_13593,N_11118);
nor U19209 (N_19209,N_14246,N_13520);
nor U19210 (N_19210,N_11659,N_10844);
nor U19211 (N_19211,N_12198,N_11219);
or U19212 (N_19212,N_13670,N_14910);
and U19213 (N_19213,N_13463,N_12791);
xnor U19214 (N_19214,N_10001,N_10897);
and U19215 (N_19215,N_12123,N_10216);
or U19216 (N_19216,N_12765,N_10274);
or U19217 (N_19217,N_10927,N_13653);
nand U19218 (N_19218,N_10878,N_14315);
xnor U19219 (N_19219,N_13515,N_11701);
nor U19220 (N_19220,N_11808,N_14187);
nor U19221 (N_19221,N_13962,N_11676);
or U19222 (N_19222,N_14764,N_12462);
nand U19223 (N_19223,N_13568,N_12063);
and U19224 (N_19224,N_12516,N_10591);
nor U19225 (N_19225,N_10672,N_11155);
and U19226 (N_19226,N_12959,N_14541);
nor U19227 (N_19227,N_13012,N_12652);
xor U19228 (N_19228,N_13480,N_11220);
nand U19229 (N_19229,N_14706,N_10669);
nor U19230 (N_19230,N_12982,N_12482);
or U19231 (N_19231,N_12907,N_12333);
and U19232 (N_19232,N_10789,N_13898);
xnor U19233 (N_19233,N_11762,N_10591);
xor U19234 (N_19234,N_14722,N_13292);
xnor U19235 (N_19235,N_10517,N_12423);
nor U19236 (N_19236,N_12237,N_11357);
and U19237 (N_19237,N_12622,N_10983);
nor U19238 (N_19238,N_13570,N_12846);
and U19239 (N_19239,N_13289,N_12620);
or U19240 (N_19240,N_13193,N_13389);
and U19241 (N_19241,N_11624,N_14335);
nand U19242 (N_19242,N_12805,N_11981);
xor U19243 (N_19243,N_11774,N_12520);
nand U19244 (N_19244,N_13706,N_12364);
and U19245 (N_19245,N_13351,N_12626);
nand U19246 (N_19246,N_10221,N_11822);
nor U19247 (N_19247,N_10799,N_14432);
nand U19248 (N_19248,N_14859,N_13221);
nor U19249 (N_19249,N_14017,N_13374);
or U19250 (N_19250,N_10048,N_11317);
xor U19251 (N_19251,N_11459,N_11110);
nand U19252 (N_19252,N_14490,N_10235);
and U19253 (N_19253,N_13137,N_12030);
or U19254 (N_19254,N_13146,N_12173);
nor U19255 (N_19255,N_13934,N_11946);
nand U19256 (N_19256,N_14659,N_10318);
nor U19257 (N_19257,N_13574,N_10411);
nand U19258 (N_19258,N_13918,N_14610);
and U19259 (N_19259,N_11089,N_11092);
and U19260 (N_19260,N_12159,N_14975);
or U19261 (N_19261,N_11804,N_10837);
nand U19262 (N_19262,N_14383,N_10964);
nand U19263 (N_19263,N_13654,N_13481);
or U19264 (N_19264,N_13628,N_10340);
nand U19265 (N_19265,N_14949,N_13592);
nor U19266 (N_19266,N_12575,N_14918);
or U19267 (N_19267,N_10118,N_11524);
nor U19268 (N_19268,N_12761,N_12644);
nand U19269 (N_19269,N_11341,N_12632);
and U19270 (N_19270,N_11951,N_12635);
nor U19271 (N_19271,N_13307,N_13237);
nand U19272 (N_19272,N_12623,N_14577);
xnor U19273 (N_19273,N_10192,N_10424);
xor U19274 (N_19274,N_11249,N_11093);
and U19275 (N_19275,N_14311,N_12357);
or U19276 (N_19276,N_11390,N_13477);
nor U19277 (N_19277,N_10344,N_12246);
nand U19278 (N_19278,N_11593,N_11471);
nor U19279 (N_19279,N_13203,N_12908);
or U19280 (N_19280,N_13430,N_10081);
and U19281 (N_19281,N_14359,N_13792);
and U19282 (N_19282,N_11216,N_11869);
nand U19283 (N_19283,N_10357,N_12773);
and U19284 (N_19284,N_14569,N_11052);
nor U19285 (N_19285,N_14006,N_11021);
or U19286 (N_19286,N_14349,N_14984);
and U19287 (N_19287,N_10194,N_12043);
nand U19288 (N_19288,N_10952,N_14385);
or U19289 (N_19289,N_14133,N_11911);
or U19290 (N_19290,N_13097,N_11026);
xor U19291 (N_19291,N_11453,N_11245);
nand U19292 (N_19292,N_11480,N_14558);
nor U19293 (N_19293,N_10830,N_13951);
nand U19294 (N_19294,N_13055,N_13634);
nand U19295 (N_19295,N_14450,N_14026);
nand U19296 (N_19296,N_11634,N_12907);
xor U19297 (N_19297,N_12004,N_11412);
and U19298 (N_19298,N_10864,N_11378);
nand U19299 (N_19299,N_11499,N_10704);
or U19300 (N_19300,N_10909,N_11908);
nand U19301 (N_19301,N_10448,N_13377);
nand U19302 (N_19302,N_14149,N_13203);
or U19303 (N_19303,N_13653,N_11919);
and U19304 (N_19304,N_14876,N_10087);
and U19305 (N_19305,N_11673,N_14276);
xnor U19306 (N_19306,N_10622,N_11435);
or U19307 (N_19307,N_12333,N_12751);
xor U19308 (N_19308,N_12001,N_12952);
nand U19309 (N_19309,N_11954,N_11267);
nand U19310 (N_19310,N_12351,N_12043);
or U19311 (N_19311,N_11593,N_14868);
xor U19312 (N_19312,N_11806,N_10749);
nand U19313 (N_19313,N_12340,N_13110);
and U19314 (N_19314,N_12004,N_14510);
nor U19315 (N_19315,N_12511,N_14621);
nand U19316 (N_19316,N_14640,N_10878);
nor U19317 (N_19317,N_12202,N_14402);
and U19318 (N_19318,N_11827,N_10604);
xnor U19319 (N_19319,N_13929,N_11092);
nor U19320 (N_19320,N_14459,N_12802);
nor U19321 (N_19321,N_11996,N_10664);
nor U19322 (N_19322,N_12399,N_10128);
nand U19323 (N_19323,N_10174,N_14980);
nor U19324 (N_19324,N_11873,N_11350);
nor U19325 (N_19325,N_12241,N_14158);
and U19326 (N_19326,N_12996,N_10339);
or U19327 (N_19327,N_14361,N_14154);
or U19328 (N_19328,N_10965,N_12914);
xor U19329 (N_19329,N_10775,N_10905);
nand U19330 (N_19330,N_13339,N_13592);
nand U19331 (N_19331,N_12091,N_13436);
nand U19332 (N_19332,N_11741,N_13955);
nand U19333 (N_19333,N_13548,N_12429);
xnor U19334 (N_19334,N_11876,N_12156);
nand U19335 (N_19335,N_12439,N_13533);
and U19336 (N_19336,N_11193,N_14080);
xor U19337 (N_19337,N_13176,N_12026);
nor U19338 (N_19338,N_13598,N_10416);
nand U19339 (N_19339,N_10155,N_14329);
and U19340 (N_19340,N_10518,N_14800);
nand U19341 (N_19341,N_11599,N_13340);
xnor U19342 (N_19342,N_12646,N_12491);
nor U19343 (N_19343,N_11884,N_12033);
or U19344 (N_19344,N_13596,N_13708);
and U19345 (N_19345,N_14918,N_11887);
or U19346 (N_19346,N_11254,N_14865);
or U19347 (N_19347,N_14659,N_11065);
or U19348 (N_19348,N_11528,N_10930);
nor U19349 (N_19349,N_13762,N_14181);
and U19350 (N_19350,N_14202,N_11443);
nor U19351 (N_19351,N_11850,N_14838);
and U19352 (N_19352,N_12544,N_12097);
nor U19353 (N_19353,N_10089,N_13142);
or U19354 (N_19354,N_14441,N_12997);
or U19355 (N_19355,N_13501,N_10889);
nand U19356 (N_19356,N_10862,N_11376);
xor U19357 (N_19357,N_11170,N_11480);
and U19358 (N_19358,N_14914,N_11693);
and U19359 (N_19359,N_14678,N_10901);
nand U19360 (N_19360,N_10536,N_12493);
or U19361 (N_19361,N_10910,N_13144);
nand U19362 (N_19362,N_10659,N_10069);
xor U19363 (N_19363,N_13972,N_11686);
nand U19364 (N_19364,N_11487,N_12891);
nand U19365 (N_19365,N_10821,N_13084);
or U19366 (N_19366,N_14518,N_12124);
nor U19367 (N_19367,N_14837,N_13318);
nor U19368 (N_19368,N_13157,N_14001);
nand U19369 (N_19369,N_11606,N_10957);
nor U19370 (N_19370,N_10598,N_11306);
nand U19371 (N_19371,N_14994,N_14337);
and U19372 (N_19372,N_11388,N_10874);
nor U19373 (N_19373,N_13329,N_11349);
nand U19374 (N_19374,N_13506,N_10493);
and U19375 (N_19375,N_14356,N_11620);
or U19376 (N_19376,N_13670,N_14529);
nor U19377 (N_19377,N_12354,N_12555);
nor U19378 (N_19378,N_11435,N_11114);
nor U19379 (N_19379,N_13776,N_12817);
and U19380 (N_19380,N_10007,N_11467);
or U19381 (N_19381,N_12693,N_11698);
nand U19382 (N_19382,N_11716,N_10882);
nor U19383 (N_19383,N_11276,N_14735);
nand U19384 (N_19384,N_12465,N_12887);
and U19385 (N_19385,N_13935,N_11519);
nand U19386 (N_19386,N_10355,N_10375);
or U19387 (N_19387,N_11947,N_14015);
or U19388 (N_19388,N_14174,N_11116);
nand U19389 (N_19389,N_10405,N_11694);
xnor U19390 (N_19390,N_12676,N_10023);
nor U19391 (N_19391,N_14457,N_11269);
nand U19392 (N_19392,N_10178,N_13617);
nor U19393 (N_19393,N_14007,N_12737);
or U19394 (N_19394,N_10825,N_13944);
xor U19395 (N_19395,N_12964,N_14906);
nand U19396 (N_19396,N_10765,N_14914);
nor U19397 (N_19397,N_12329,N_13861);
or U19398 (N_19398,N_14381,N_12709);
or U19399 (N_19399,N_11094,N_14307);
nor U19400 (N_19400,N_10878,N_12573);
nand U19401 (N_19401,N_11099,N_14765);
nand U19402 (N_19402,N_13182,N_10756);
or U19403 (N_19403,N_12942,N_14414);
nor U19404 (N_19404,N_10127,N_10964);
nand U19405 (N_19405,N_13869,N_14573);
nand U19406 (N_19406,N_12300,N_12263);
nand U19407 (N_19407,N_14082,N_10676);
xor U19408 (N_19408,N_11237,N_14756);
nor U19409 (N_19409,N_12364,N_11061);
nand U19410 (N_19410,N_10121,N_12081);
and U19411 (N_19411,N_12144,N_12296);
nand U19412 (N_19412,N_12368,N_13704);
or U19413 (N_19413,N_11966,N_12778);
and U19414 (N_19414,N_11096,N_10499);
xnor U19415 (N_19415,N_12811,N_13862);
and U19416 (N_19416,N_12792,N_10159);
xnor U19417 (N_19417,N_10762,N_14430);
xnor U19418 (N_19418,N_10697,N_11592);
xor U19419 (N_19419,N_10066,N_11595);
and U19420 (N_19420,N_10332,N_13049);
xor U19421 (N_19421,N_13750,N_14055);
nor U19422 (N_19422,N_14085,N_13469);
or U19423 (N_19423,N_12137,N_11057);
nor U19424 (N_19424,N_11237,N_12209);
nand U19425 (N_19425,N_14237,N_10918);
or U19426 (N_19426,N_13480,N_11914);
or U19427 (N_19427,N_14211,N_11955);
or U19428 (N_19428,N_11742,N_12734);
nor U19429 (N_19429,N_13058,N_10476);
and U19430 (N_19430,N_10974,N_11841);
and U19431 (N_19431,N_12510,N_13686);
xnor U19432 (N_19432,N_11451,N_13360);
nor U19433 (N_19433,N_11602,N_11841);
or U19434 (N_19434,N_10852,N_10536);
and U19435 (N_19435,N_11409,N_11947);
and U19436 (N_19436,N_11238,N_13058);
nand U19437 (N_19437,N_11350,N_12088);
xor U19438 (N_19438,N_11496,N_13363);
and U19439 (N_19439,N_13477,N_13990);
xor U19440 (N_19440,N_11587,N_12465);
nor U19441 (N_19441,N_11772,N_10514);
nor U19442 (N_19442,N_11489,N_10719);
nand U19443 (N_19443,N_14976,N_11305);
nand U19444 (N_19444,N_14787,N_13237);
nor U19445 (N_19445,N_11995,N_12958);
or U19446 (N_19446,N_12316,N_13800);
and U19447 (N_19447,N_13159,N_12713);
and U19448 (N_19448,N_14776,N_10502);
nand U19449 (N_19449,N_11390,N_10678);
and U19450 (N_19450,N_13649,N_12484);
nand U19451 (N_19451,N_13677,N_12228);
or U19452 (N_19452,N_12190,N_13589);
xor U19453 (N_19453,N_12605,N_13866);
or U19454 (N_19454,N_13834,N_13334);
or U19455 (N_19455,N_12515,N_14225);
nor U19456 (N_19456,N_13933,N_14809);
or U19457 (N_19457,N_10488,N_14857);
and U19458 (N_19458,N_12166,N_11638);
nor U19459 (N_19459,N_14128,N_11958);
and U19460 (N_19460,N_13471,N_13577);
or U19461 (N_19461,N_11632,N_13320);
nand U19462 (N_19462,N_11208,N_12465);
xor U19463 (N_19463,N_13652,N_11366);
or U19464 (N_19464,N_13676,N_10589);
nor U19465 (N_19465,N_12406,N_13051);
xor U19466 (N_19466,N_11311,N_10894);
and U19467 (N_19467,N_12626,N_13938);
and U19468 (N_19468,N_14585,N_10673);
nor U19469 (N_19469,N_10075,N_12935);
nor U19470 (N_19470,N_10400,N_13873);
or U19471 (N_19471,N_13299,N_12010);
or U19472 (N_19472,N_14969,N_10101);
nand U19473 (N_19473,N_12400,N_11776);
nor U19474 (N_19474,N_12919,N_11333);
nand U19475 (N_19475,N_10179,N_12572);
nor U19476 (N_19476,N_13769,N_12831);
nand U19477 (N_19477,N_10877,N_11650);
xnor U19478 (N_19478,N_11963,N_10249);
and U19479 (N_19479,N_10042,N_13983);
and U19480 (N_19480,N_12088,N_13188);
or U19481 (N_19481,N_11963,N_12791);
or U19482 (N_19482,N_10270,N_12216);
or U19483 (N_19483,N_14708,N_12200);
or U19484 (N_19484,N_14158,N_13809);
or U19485 (N_19485,N_12054,N_10818);
nor U19486 (N_19486,N_13353,N_10185);
or U19487 (N_19487,N_13992,N_11282);
nor U19488 (N_19488,N_12159,N_12355);
or U19489 (N_19489,N_13505,N_13039);
or U19490 (N_19490,N_13937,N_14163);
nand U19491 (N_19491,N_10815,N_11505);
xor U19492 (N_19492,N_11374,N_14852);
or U19493 (N_19493,N_13974,N_11302);
nand U19494 (N_19494,N_10146,N_12442);
and U19495 (N_19495,N_14636,N_11400);
and U19496 (N_19496,N_14861,N_14824);
or U19497 (N_19497,N_13704,N_12194);
and U19498 (N_19498,N_10950,N_12670);
and U19499 (N_19499,N_12183,N_11258);
or U19500 (N_19500,N_11067,N_11812);
nand U19501 (N_19501,N_14176,N_11607);
or U19502 (N_19502,N_13518,N_12204);
or U19503 (N_19503,N_14906,N_12336);
or U19504 (N_19504,N_10514,N_10202);
nor U19505 (N_19505,N_14224,N_12457);
nor U19506 (N_19506,N_14024,N_14072);
xnor U19507 (N_19507,N_14425,N_14158);
nor U19508 (N_19508,N_14433,N_13033);
or U19509 (N_19509,N_13657,N_10370);
or U19510 (N_19510,N_11598,N_10958);
xor U19511 (N_19511,N_11714,N_14328);
nor U19512 (N_19512,N_11651,N_13293);
xor U19513 (N_19513,N_14702,N_13775);
or U19514 (N_19514,N_13987,N_13936);
and U19515 (N_19515,N_13674,N_11502);
or U19516 (N_19516,N_14134,N_13810);
or U19517 (N_19517,N_14818,N_11081);
nand U19518 (N_19518,N_10489,N_13190);
or U19519 (N_19519,N_13374,N_14575);
and U19520 (N_19520,N_13411,N_11963);
nand U19521 (N_19521,N_13026,N_10536);
and U19522 (N_19522,N_10166,N_10886);
nand U19523 (N_19523,N_13361,N_10330);
or U19524 (N_19524,N_10254,N_13368);
xor U19525 (N_19525,N_14801,N_14759);
and U19526 (N_19526,N_13364,N_10828);
nor U19527 (N_19527,N_11841,N_11911);
nand U19528 (N_19528,N_10320,N_13164);
xor U19529 (N_19529,N_12359,N_14219);
and U19530 (N_19530,N_14122,N_11647);
and U19531 (N_19531,N_13643,N_12380);
nor U19532 (N_19532,N_14759,N_14222);
and U19533 (N_19533,N_10623,N_11965);
nor U19534 (N_19534,N_11034,N_14118);
nand U19535 (N_19535,N_13359,N_14977);
or U19536 (N_19536,N_12018,N_10217);
and U19537 (N_19537,N_11955,N_14910);
and U19538 (N_19538,N_12777,N_14894);
xnor U19539 (N_19539,N_10862,N_14882);
nor U19540 (N_19540,N_13916,N_10341);
or U19541 (N_19541,N_13525,N_10853);
and U19542 (N_19542,N_14181,N_11755);
or U19543 (N_19543,N_13760,N_13881);
nand U19544 (N_19544,N_11204,N_11480);
or U19545 (N_19545,N_12664,N_13030);
nor U19546 (N_19546,N_10262,N_12497);
nand U19547 (N_19547,N_13119,N_11452);
xor U19548 (N_19548,N_10272,N_12281);
and U19549 (N_19549,N_13269,N_12751);
or U19550 (N_19550,N_10970,N_14951);
and U19551 (N_19551,N_12292,N_14095);
and U19552 (N_19552,N_13441,N_14010);
nand U19553 (N_19553,N_12894,N_12825);
xor U19554 (N_19554,N_14759,N_13969);
nand U19555 (N_19555,N_13151,N_14048);
nor U19556 (N_19556,N_10315,N_10003);
and U19557 (N_19557,N_12025,N_10813);
and U19558 (N_19558,N_13021,N_14161);
nor U19559 (N_19559,N_10473,N_11314);
nand U19560 (N_19560,N_13642,N_12694);
and U19561 (N_19561,N_14661,N_12427);
and U19562 (N_19562,N_11966,N_14430);
nor U19563 (N_19563,N_11522,N_12989);
nand U19564 (N_19564,N_13002,N_13614);
or U19565 (N_19565,N_10079,N_11785);
nor U19566 (N_19566,N_11555,N_14279);
xor U19567 (N_19567,N_11461,N_12959);
nor U19568 (N_19568,N_10502,N_12638);
and U19569 (N_19569,N_11875,N_11071);
nor U19570 (N_19570,N_13853,N_13192);
and U19571 (N_19571,N_12471,N_10907);
and U19572 (N_19572,N_13862,N_13341);
and U19573 (N_19573,N_12717,N_13501);
or U19574 (N_19574,N_11780,N_12944);
xnor U19575 (N_19575,N_14550,N_13448);
xnor U19576 (N_19576,N_14662,N_11849);
nand U19577 (N_19577,N_13297,N_10511);
or U19578 (N_19578,N_11836,N_11498);
and U19579 (N_19579,N_11811,N_13194);
or U19580 (N_19580,N_13570,N_12415);
nand U19581 (N_19581,N_14915,N_11924);
nor U19582 (N_19582,N_13725,N_10904);
nand U19583 (N_19583,N_11099,N_14785);
nand U19584 (N_19584,N_13247,N_11756);
or U19585 (N_19585,N_13489,N_14215);
or U19586 (N_19586,N_11371,N_11999);
or U19587 (N_19587,N_11395,N_11358);
or U19588 (N_19588,N_11218,N_11874);
nor U19589 (N_19589,N_11412,N_14504);
and U19590 (N_19590,N_13365,N_14259);
nand U19591 (N_19591,N_13623,N_10290);
and U19592 (N_19592,N_13444,N_12549);
and U19593 (N_19593,N_11537,N_14871);
xor U19594 (N_19594,N_13358,N_10054);
xnor U19595 (N_19595,N_13975,N_10724);
nor U19596 (N_19596,N_10505,N_10852);
or U19597 (N_19597,N_13921,N_13414);
or U19598 (N_19598,N_12912,N_11017);
nand U19599 (N_19599,N_11286,N_11003);
and U19600 (N_19600,N_11569,N_14116);
and U19601 (N_19601,N_10397,N_12393);
or U19602 (N_19602,N_11339,N_11155);
or U19603 (N_19603,N_11731,N_11574);
and U19604 (N_19604,N_13317,N_12566);
nand U19605 (N_19605,N_12639,N_14596);
or U19606 (N_19606,N_11325,N_13837);
nor U19607 (N_19607,N_10047,N_13337);
nor U19608 (N_19608,N_11452,N_13709);
or U19609 (N_19609,N_13633,N_11412);
or U19610 (N_19610,N_10774,N_10876);
nand U19611 (N_19611,N_13883,N_13389);
and U19612 (N_19612,N_10989,N_10956);
or U19613 (N_19613,N_12511,N_10546);
xor U19614 (N_19614,N_11122,N_10376);
and U19615 (N_19615,N_11259,N_14748);
and U19616 (N_19616,N_11468,N_11572);
and U19617 (N_19617,N_12338,N_12782);
nor U19618 (N_19618,N_10689,N_14517);
or U19619 (N_19619,N_10800,N_11320);
nand U19620 (N_19620,N_13627,N_12566);
or U19621 (N_19621,N_12505,N_13732);
nor U19622 (N_19622,N_11931,N_12934);
nand U19623 (N_19623,N_13247,N_13045);
or U19624 (N_19624,N_11415,N_10295);
or U19625 (N_19625,N_10575,N_11208);
xor U19626 (N_19626,N_11931,N_13649);
or U19627 (N_19627,N_14881,N_14175);
or U19628 (N_19628,N_13514,N_10439);
or U19629 (N_19629,N_14097,N_12723);
and U19630 (N_19630,N_12609,N_13318);
or U19631 (N_19631,N_12157,N_14625);
and U19632 (N_19632,N_13997,N_10334);
and U19633 (N_19633,N_14638,N_12913);
or U19634 (N_19634,N_12627,N_14999);
nand U19635 (N_19635,N_14428,N_12136);
nor U19636 (N_19636,N_11411,N_13626);
and U19637 (N_19637,N_12539,N_13241);
or U19638 (N_19638,N_13552,N_12198);
and U19639 (N_19639,N_12233,N_12388);
and U19640 (N_19640,N_11577,N_13751);
nand U19641 (N_19641,N_14495,N_12092);
nand U19642 (N_19642,N_11939,N_10118);
nand U19643 (N_19643,N_10690,N_10896);
nor U19644 (N_19644,N_14634,N_10255);
nand U19645 (N_19645,N_11709,N_10158);
or U19646 (N_19646,N_14539,N_12670);
or U19647 (N_19647,N_14049,N_13100);
and U19648 (N_19648,N_13714,N_11628);
nor U19649 (N_19649,N_13003,N_13476);
nand U19650 (N_19650,N_12527,N_11810);
nor U19651 (N_19651,N_11108,N_12320);
nand U19652 (N_19652,N_11391,N_10157);
or U19653 (N_19653,N_13475,N_11302);
nor U19654 (N_19654,N_10764,N_12929);
xor U19655 (N_19655,N_11807,N_13753);
and U19656 (N_19656,N_12085,N_14447);
or U19657 (N_19657,N_13150,N_12752);
nand U19658 (N_19658,N_14770,N_14712);
and U19659 (N_19659,N_12115,N_11774);
nand U19660 (N_19660,N_11797,N_14680);
xor U19661 (N_19661,N_13305,N_10081);
or U19662 (N_19662,N_10314,N_10381);
nor U19663 (N_19663,N_14076,N_14889);
or U19664 (N_19664,N_10211,N_11271);
nor U19665 (N_19665,N_10446,N_14565);
nor U19666 (N_19666,N_10674,N_11296);
nor U19667 (N_19667,N_10434,N_12510);
nand U19668 (N_19668,N_12098,N_11622);
xor U19669 (N_19669,N_13653,N_11826);
and U19670 (N_19670,N_12540,N_10389);
and U19671 (N_19671,N_13034,N_14694);
or U19672 (N_19672,N_10696,N_12304);
nor U19673 (N_19673,N_12589,N_14064);
nor U19674 (N_19674,N_11793,N_13517);
nand U19675 (N_19675,N_14351,N_11246);
nand U19676 (N_19676,N_12387,N_12480);
nand U19677 (N_19677,N_14118,N_14491);
and U19678 (N_19678,N_14454,N_10670);
xnor U19679 (N_19679,N_11946,N_11842);
nand U19680 (N_19680,N_11385,N_14763);
or U19681 (N_19681,N_11366,N_13464);
nand U19682 (N_19682,N_14083,N_11492);
xnor U19683 (N_19683,N_11620,N_10788);
xor U19684 (N_19684,N_10970,N_12779);
nand U19685 (N_19685,N_12770,N_13381);
nor U19686 (N_19686,N_13457,N_14588);
nand U19687 (N_19687,N_14480,N_12403);
or U19688 (N_19688,N_10634,N_14388);
or U19689 (N_19689,N_11184,N_10381);
nand U19690 (N_19690,N_14851,N_14458);
xnor U19691 (N_19691,N_10452,N_10611);
xnor U19692 (N_19692,N_14931,N_14194);
nor U19693 (N_19693,N_14776,N_13138);
and U19694 (N_19694,N_10568,N_13800);
and U19695 (N_19695,N_14735,N_10440);
or U19696 (N_19696,N_14768,N_13741);
and U19697 (N_19697,N_14574,N_11592);
nor U19698 (N_19698,N_14314,N_11548);
or U19699 (N_19699,N_13096,N_11406);
nor U19700 (N_19700,N_13204,N_11075);
nor U19701 (N_19701,N_12330,N_13120);
nand U19702 (N_19702,N_14976,N_11903);
or U19703 (N_19703,N_12170,N_11782);
and U19704 (N_19704,N_14844,N_14484);
nor U19705 (N_19705,N_14083,N_13956);
and U19706 (N_19706,N_12876,N_13470);
nor U19707 (N_19707,N_11236,N_11603);
nor U19708 (N_19708,N_12786,N_12726);
or U19709 (N_19709,N_10995,N_13564);
nor U19710 (N_19710,N_13771,N_10168);
or U19711 (N_19711,N_14683,N_13233);
or U19712 (N_19712,N_10322,N_10663);
or U19713 (N_19713,N_12738,N_14265);
or U19714 (N_19714,N_10686,N_10636);
and U19715 (N_19715,N_10716,N_11770);
xor U19716 (N_19716,N_14350,N_13197);
and U19717 (N_19717,N_14563,N_12115);
or U19718 (N_19718,N_11987,N_13610);
nand U19719 (N_19719,N_10547,N_11843);
and U19720 (N_19720,N_11988,N_13254);
nor U19721 (N_19721,N_11535,N_13844);
nand U19722 (N_19722,N_10911,N_12362);
and U19723 (N_19723,N_12318,N_12399);
nand U19724 (N_19724,N_10706,N_10961);
or U19725 (N_19725,N_13172,N_11865);
and U19726 (N_19726,N_11091,N_14191);
nand U19727 (N_19727,N_14259,N_12081);
nand U19728 (N_19728,N_14104,N_14359);
and U19729 (N_19729,N_14865,N_14034);
and U19730 (N_19730,N_10671,N_10961);
nor U19731 (N_19731,N_14385,N_11730);
or U19732 (N_19732,N_14030,N_14288);
or U19733 (N_19733,N_11005,N_11050);
nand U19734 (N_19734,N_13050,N_13325);
xnor U19735 (N_19735,N_14917,N_12042);
or U19736 (N_19736,N_14537,N_13395);
and U19737 (N_19737,N_14232,N_13585);
xnor U19738 (N_19738,N_11476,N_14865);
nand U19739 (N_19739,N_13156,N_11306);
or U19740 (N_19740,N_12182,N_13140);
nor U19741 (N_19741,N_13317,N_13754);
and U19742 (N_19742,N_13028,N_12403);
nand U19743 (N_19743,N_12741,N_12368);
nor U19744 (N_19744,N_13967,N_13208);
and U19745 (N_19745,N_13467,N_11069);
or U19746 (N_19746,N_14894,N_14645);
xor U19747 (N_19747,N_12839,N_13689);
nor U19748 (N_19748,N_14991,N_11610);
nand U19749 (N_19749,N_13920,N_14009);
and U19750 (N_19750,N_10617,N_10350);
nor U19751 (N_19751,N_14544,N_10342);
nand U19752 (N_19752,N_12145,N_11206);
nor U19753 (N_19753,N_11462,N_10988);
xnor U19754 (N_19754,N_12516,N_11128);
nor U19755 (N_19755,N_10535,N_13155);
nand U19756 (N_19756,N_12738,N_13037);
nor U19757 (N_19757,N_12807,N_12750);
and U19758 (N_19758,N_14047,N_10862);
nand U19759 (N_19759,N_13338,N_13001);
nor U19760 (N_19760,N_13913,N_11146);
and U19761 (N_19761,N_14001,N_11129);
and U19762 (N_19762,N_13686,N_13471);
and U19763 (N_19763,N_12567,N_13565);
and U19764 (N_19764,N_13095,N_12827);
nor U19765 (N_19765,N_12496,N_11724);
xnor U19766 (N_19766,N_12639,N_11684);
or U19767 (N_19767,N_10767,N_11807);
and U19768 (N_19768,N_12640,N_14769);
or U19769 (N_19769,N_14292,N_10342);
and U19770 (N_19770,N_12250,N_13867);
nor U19771 (N_19771,N_10808,N_10132);
nand U19772 (N_19772,N_13812,N_11842);
nand U19773 (N_19773,N_10951,N_11166);
nor U19774 (N_19774,N_10699,N_11033);
or U19775 (N_19775,N_13589,N_12962);
nor U19776 (N_19776,N_13917,N_12947);
and U19777 (N_19777,N_14535,N_11609);
or U19778 (N_19778,N_12114,N_12102);
or U19779 (N_19779,N_10538,N_11121);
nand U19780 (N_19780,N_14893,N_14487);
nand U19781 (N_19781,N_11815,N_14392);
xnor U19782 (N_19782,N_14203,N_13445);
xnor U19783 (N_19783,N_12352,N_12467);
or U19784 (N_19784,N_14484,N_10613);
nor U19785 (N_19785,N_11868,N_13838);
nor U19786 (N_19786,N_11560,N_13490);
nand U19787 (N_19787,N_14726,N_14606);
or U19788 (N_19788,N_14936,N_11872);
nand U19789 (N_19789,N_14018,N_11917);
nand U19790 (N_19790,N_14726,N_10670);
and U19791 (N_19791,N_12424,N_10926);
nor U19792 (N_19792,N_14516,N_14358);
nand U19793 (N_19793,N_12442,N_11064);
and U19794 (N_19794,N_11870,N_10393);
or U19795 (N_19795,N_10685,N_12553);
or U19796 (N_19796,N_10350,N_11796);
nand U19797 (N_19797,N_12982,N_11372);
or U19798 (N_19798,N_10078,N_10337);
nand U19799 (N_19799,N_11203,N_13214);
or U19800 (N_19800,N_10598,N_12385);
nor U19801 (N_19801,N_12932,N_12188);
and U19802 (N_19802,N_12885,N_11759);
or U19803 (N_19803,N_10587,N_10535);
nand U19804 (N_19804,N_12636,N_14920);
nand U19805 (N_19805,N_13451,N_10347);
xor U19806 (N_19806,N_14217,N_14265);
nand U19807 (N_19807,N_13292,N_10228);
and U19808 (N_19808,N_11417,N_10031);
nand U19809 (N_19809,N_11838,N_11981);
xor U19810 (N_19810,N_12606,N_13935);
or U19811 (N_19811,N_14420,N_14516);
and U19812 (N_19812,N_11976,N_10806);
nand U19813 (N_19813,N_14119,N_14096);
nor U19814 (N_19814,N_10576,N_13762);
nor U19815 (N_19815,N_12317,N_12863);
nand U19816 (N_19816,N_12648,N_11364);
nor U19817 (N_19817,N_10740,N_13432);
nand U19818 (N_19818,N_11003,N_14834);
or U19819 (N_19819,N_12684,N_13735);
nand U19820 (N_19820,N_12226,N_11933);
or U19821 (N_19821,N_11436,N_11664);
or U19822 (N_19822,N_13963,N_14523);
nand U19823 (N_19823,N_12015,N_11031);
nand U19824 (N_19824,N_12194,N_14954);
nor U19825 (N_19825,N_10223,N_12581);
nor U19826 (N_19826,N_14951,N_13862);
nand U19827 (N_19827,N_14277,N_12350);
or U19828 (N_19828,N_13187,N_14117);
or U19829 (N_19829,N_12907,N_13254);
or U19830 (N_19830,N_12888,N_12701);
nand U19831 (N_19831,N_14247,N_11768);
and U19832 (N_19832,N_14941,N_12941);
xor U19833 (N_19833,N_13064,N_14950);
nor U19834 (N_19834,N_12078,N_13156);
or U19835 (N_19835,N_11298,N_14384);
or U19836 (N_19836,N_10569,N_10363);
xor U19837 (N_19837,N_14199,N_13170);
or U19838 (N_19838,N_14015,N_10456);
and U19839 (N_19839,N_11003,N_14843);
nor U19840 (N_19840,N_14562,N_10842);
or U19841 (N_19841,N_12636,N_13242);
nand U19842 (N_19842,N_11476,N_13386);
or U19843 (N_19843,N_10745,N_14333);
and U19844 (N_19844,N_14058,N_12893);
or U19845 (N_19845,N_11641,N_11019);
and U19846 (N_19846,N_14140,N_13692);
xor U19847 (N_19847,N_14804,N_10184);
and U19848 (N_19848,N_11854,N_12195);
and U19849 (N_19849,N_14074,N_14829);
and U19850 (N_19850,N_10311,N_14392);
nand U19851 (N_19851,N_13271,N_12910);
nand U19852 (N_19852,N_14739,N_13557);
or U19853 (N_19853,N_11532,N_13187);
nand U19854 (N_19854,N_10448,N_14500);
or U19855 (N_19855,N_13042,N_11634);
and U19856 (N_19856,N_12588,N_13656);
nand U19857 (N_19857,N_14314,N_11704);
and U19858 (N_19858,N_10286,N_13293);
and U19859 (N_19859,N_12459,N_12175);
nor U19860 (N_19860,N_13146,N_14002);
nor U19861 (N_19861,N_10200,N_12645);
nor U19862 (N_19862,N_14335,N_10616);
nor U19863 (N_19863,N_10024,N_11555);
nand U19864 (N_19864,N_12476,N_12712);
nor U19865 (N_19865,N_12961,N_12722);
xnor U19866 (N_19866,N_14907,N_12690);
and U19867 (N_19867,N_10416,N_14398);
and U19868 (N_19868,N_12185,N_10975);
nor U19869 (N_19869,N_10899,N_13774);
nor U19870 (N_19870,N_14315,N_13348);
nor U19871 (N_19871,N_14470,N_12514);
nand U19872 (N_19872,N_11238,N_11030);
nand U19873 (N_19873,N_14656,N_14861);
nor U19874 (N_19874,N_12146,N_12826);
nand U19875 (N_19875,N_13920,N_11093);
nand U19876 (N_19876,N_12877,N_11681);
nor U19877 (N_19877,N_11201,N_13407);
or U19878 (N_19878,N_13394,N_13041);
and U19879 (N_19879,N_10491,N_11338);
nor U19880 (N_19880,N_10295,N_14349);
nor U19881 (N_19881,N_12308,N_13929);
nor U19882 (N_19882,N_11304,N_12930);
and U19883 (N_19883,N_10598,N_10894);
or U19884 (N_19884,N_10077,N_13073);
and U19885 (N_19885,N_10231,N_14183);
and U19886 (N_19886,N_10029,N_13475);
and U19887 (N_19887,N_11367,N_14760);
and U19888 (N_19888,N_13096,N_10057);
xnor U19889 (N_19889,N_10152,N_11924);
or U19890 (N_19890,N_14328,N_10628);
nor U19891 (N_19891,N_11806,N_10472);
and U19892 (N_19892,N_12719,N_13707);
or U19893 (N_19893,N_13680,N_12673);
nand U19894 (N_19894,N_10580,N_14609);
nor U19895 (N_19895,N_14477,N_13533);
nor U19896 (N_19896,N_10514,N_13601);
nor U19897 (N_19897,N_13196,N_14697);
or U19898 (N_19898,N_11434,N_12798);
and U19899 (N_19899,N_12510,N_13901);
nand U19900 (N_19900,N_13275,N_12928);
nor U19901 (N_19901,N_13481,N_10752);
nand U19902 (N_19902,N_13782,N_13369);
nand U19903 (N_19903,N_10413,N_12252);
or U19904 (N_19904,N_14924,N_14048);
xnor U19905 (N_19905,N_11903,N_14205);
nor U19906 (N_19906,N_13239,N_14753);
or U19907 (N_19907,N_11228,N_11030);
nand U19908 (N_19908,N_13701,N_11228);
nor U19909 (N_19909,N_10807,N_13391);
and U19910 (N_19910,N_11809,N_13357);
nand U19911 (N_19911,N_10770,N_11183);
or U19912 (N_19912,N_12355,N_11251);
or U19913 (N_19913,N_11742,N_14674);
or U19914 (N_19914,N_10267,N_10105);
nand U19915 (N_19915,N_12287,N_11643);
nor U19916 (N_19916,N_10388,N_14748);
or U19917 (N_19917,N_10610,N_14420);
nor U19918 (N_19918,N_13341,N_11585);
nor U19919 (N_19919,N_11088,N_12386);
or U19920 (N_19920,N_10411,N_13147);
and U19921 (N_19921,N_13000,N_13444);
or U19922 (N_19922,N_13478,N_10029);
nand U19923 (N_19923,N_11316,N_10245);
or U19924 (N_19924,N_12736,N_14674);
or U19925 (N_19925,N_10996,N_12822);
nor U19926 (N_19926,N_14794,N_13286);
and U19927 (N_19927,N_14468,N_12726);
nand U19928 (N_19928,N_14645,N_11691);
and U19929 (N_19929,N_11958,N_13341);
and U19930 (N_19930,N_13753,N_12137);
nand U19931 (N_19931,N_14885,N_10085);
or U19932 (N_19932,N_14731,N_11702);
or U19933 (N_19933,N_11485,N_13231);
or U19934 (N_19934,N_10756,N_12615);
or U19935 (N_19935,N_12710,N_10671);
nand U19936 (N_19936,N_10308,N_13832);
and U19937 (N_19937,N_10863,N_12133);
nand U19938 (N_19938,N_14300,N_12995);
xnor U19939 (N_19939,N_12447,N_13489);
nor U19940 (N_19940,N_12693,N_10120);
nor U19941 (N_19941,N_10439,N_10227);
xnor U19942 (N_19942,N_14015,N_10653);
or U19943 (N_19943,N_11424,N_10769);
and U19944 (N_19944,N_14552,N_10828);
nor U19945 (N_19945,N_13300,N_11030);
nand U19946 (N_19946,N_11069,N_10855);
and U19947 (N_19947,N_13487,N_13984);
nand U19948 (N_19948,N_11215,N_11356);
nand U19949 (N_19949,N_10054,N_13925);
nand U19950 (N_19950,N_14496,N_12880);
or U19951 (N_19951,N_12089,N_10047);
or U19952 (N_19952,N_10910,N_13273);
nand U19953 (N_19953,N_13038,N_10859);
nand U19954 (N_19954,N_12953,N_11913);
and U19955 (N_19955,N_14678,N_13803);
nor U19956 (N_19956,N_12368,N_13283);
nand U19957 (N_19957,N_10716,N_12982);
or U19958 (N_19958,N_11530,N_13435);
nor U19959 (N_19959,N_10759,N_11406);
and U19960 (N_19960,N_10418,N_10078);
or U19961 (N_19961,N_10631,N_10948);
nand U19962 (N_19962,N_10084,N_14007);
and U19963 (N_19963,N_14536,N_14445);
nor U19964 (N_19964,N_12408,N_12291);
or U19965 (N_19965,N_12027,N_10448);
nand U19966 (N_19966,N_13088,N_13002);
nor U19967 (N_19967,N_12813,N_10558);
nand U19968 (N_19968,N_11888,N_14402);
and U19969 (N_19969,N_12347,N_10072);
nand U19970 (N_19970,N_14462,N_14165);
nand U19971 (N_19971,N_10750,N_11719);
and U19972 (N_19972,N_14570,N_10345);
xnor U19973 (N_19973,N_10492,N_11843);
or U19974 (N_19974,N_11247,N_10380);
nor U19975 (N_19975,N_10368,N_12307);
or U19976 (N_19976,N_12164,N_10129);
or U19977 (N_19977,N_11788,N_13033);
nor U19978 (N_19978,N_14194,N_11563);
nor U19979 (N_19979,N_11061,N_14887);
nand U19980 (N_19980,N_10580,N_13174);
or U19981 (N_19981,N_12296,N_13246);
or U19982 (N_19982,N_10762,N_13269);
and U19983 (N_19983,N_14462,N_14528);
and U19984 (N_19984,N_10903,N_12032);
xor U19985 (N_19985,N_14718,N_12343);
nand U19986 (N_19986,N_10990,N_11172);
and U19987 (N_19987,N_12860,N_12630);
and U19988 (N_19988,N_14476,N_12629);
nand U19989 (N_19989,N_10785,N_12061);
and U19990 (N_19990,N_11237,N_10150);
nand U19991 (N_19991,N_13424,N_11256);
nor U19992 (N_19992,N_10872,N_14708);
or U19993 (N_19993,N_13985,N_12383);
nor U19994 (N_19994,N_12915,N_14900);
nor U19995 (N_19995,N_12512,N_10966);
and U19996 (N_19996,N_12393,N_12754);
nand U19997 (N_19997,N_11528,N_12624);
and U19998 (N_19998,N_10014,N_12162);
and U19999 (N_19999,N_13744,N_12390);
or U20000 (N_20000,N_18562,N_15927);
or U20001 (N_20001,N_16901,N_16746);
or U20002 (N_20002,N_18569,N_19682);
nand U20003 (N_20003,N_17487,N_15644);
nor U20004 (N_20004,N_19087,N_17667);
and U20005 (N_20005,N_16864,N_18210);
and U20006 (N_20006,N_18791,N_17654);
and U20007 (N_20007,N_18732,N_17794);
nor U20008 (N_20008,N_17536,N_19191);
nand U20009 (N_20009,N_18522,N_18276);
nand U20010 (N_20010,N_19127,N_16650);
or U20011 (N_20011,N_16114,N_19203);
nor U20012 (N_20012,N_18837,N_18311);
or U20013 (N_20013,N_17953,N_18401);
nand U20014 (N_20014,N_18334,N_19985);
nand U20015 (N_20015,N_17223,N_15460);
or U20016 (N_20016,N_16818,N_19181);
nand U20017 (N_20017,N_16172,N_19495);
xnor U20018 (N_20018,N_15033,N_16899);
nor U20019 (N_20019,N_19205,N_16151);
or U20020 (N_20020,N_17323,N_15404);
nand U20021 (N_20021,N_18788,N_15590);
or U20022 (N_20022,N_18068,N_15826);
nand U20023 (N_20023,N_15022,N_19404);
or U20024 (N_20024,N_18138,N_19328);
or U20025 (N_20025,N_15709,N_15768);
xor U20026 (N_20026,N_15700,N_15915);
xnor U20027 (N_20027,N_17244,N_18187);
nand U20028 (N_20028,N_16401,N_16195);
or U20029 (N_20029,N_18353,N_18190);
xnor U20030 (N_20030,N_15438,N_17203);
nor U20031 (N_20031,N_15668,N_17152);
and U20032 (N_20032,N_16801,N_15426);
xor U20033 (N_20033,N_17760,N_16597);
or U20034 (N_20034,N_18978,N_16963);
nor U20035 (N_20035,N_15048,N_19422);
and U20036 (N_20036,N_16196,N_17922);
or U20037 (N_20037,N_15511,N_17142);
nand U20038 (N_20038,N_19009,N_16904);
nand U20039 (N_20039,N_18680,N_16451);
nand U20040 (N_20040,N_19669,N_19490);
and U20041 (N_20041,N_18727,N_19355);
nor U20042 (N_20042,N_18629,N_18163);
or U20043 (N_20043,N_16360,N_15820);
nor U20044 (N_20044,N_18537,N_17039);
and U20045 (N_20045,N_19762,N_16435);
xnor U20046 (N_20046,N_19760,N_19510);
nor U20047 (N_20047,N_15228,N_17421);
nand U20048 (N_20048,N_16197,N_17617);
nand U20049 (N_20049,N_15948,N_15113);
or U20050 (N_20050,N_18570,N_17878);
and U20051 (N_20051,N_15951,N_17567);
and U20052 (N_20052,N_19357,N_16079);
and U20053 (N_20053,N_17026,N_15373);
nand U20054 (N_20054,N_19242,N_19256);
xor U20055 (N_20055,N_19236,N_15970);
and U20056 (N_20056,N_18478,N_19953);
or U20057 (N_20057,N_18760,N_19292);
or U20058 (N_20058,N_18656,N_16124);
nand U20059 (N_20059,N_17797,N_19403);
or U20060 (N_20060,N_15338,N_17798);
or U20061 (N_20061,N_19830,N_18740);
and U20062 (N_20062,N_15221,N_17159);
nand U20063 (N_20063,N_18500,N_17360);
nand U20064 (N_20064,N_18599,N_15642);
nor U20065 (N_20065,N_18563,N_16638);
or U20066 (N_20066,N_15576,N_17095);
nor U20067 (N_20067,N_18855,N_15300);
nor U20068 (N_20068,N_16331,N_15715);
nor U20069 (N_20069,N_16406,N_17538);
nand U20070 (N_20070,N_16300,N_19590);
nor U20071 (N_20071,N_16689,N_15660);
nand U20072 (N_20072,N_17201,N_16341);
or U20073 (N_20073,N_18256,N_19136);
nor U20074 (N_20074,N_19179,N_19920);
nor U20075 (N_20075,N_18428,N_18008);
nor U20076 (N_20076,N_18691,N_17022);
or U20077 (N_20077,N_15043,N_17348);
nand U20078 (N_20078,N_16103,N_16775);
nor U20079 (N_20079,N_18636,N_16890);
and U20080 (N_20080,N_18745,N_19877);
or U20081 (N_20081,N_19408,N_16003);
or U20082 (N_20082,N_16660,N_17818);
and U20083 (N_20083,N_19588,N_16387);
and U20084 (N_20084,N_18280,N_19980);
nand U20085 (N_20085,N_17997,N_16822);
and U20086 (N_20086,N_16722,N_17415);
or U20087 (N_20087,N_16239,N_16572);
or U20088 (N_20088,N_19098,N_15215);
or U20089 (N_20089,N_15764,N_15792);
or U20090 (N_20090,N_15110,N_18083);
nor U20091 (N_20091,N_15123,N_19166);
nand U20092 (N_20092,N_18771,N_18447);
nor U20093 (N_20093,N_18886,N_16519);
nand U20094 (N_20094,N_15530,N_16998);
nor U20095 (N_20095,N_15706,N_17719);
nor U20096 (N_20096,N_17626,N_18889);
nand U20097 (N_20097,N_18031,N_18956);
nor U20098 (N_20098,N_17989,N_17119);
nor U20099 (N_20099,N_18526,N_17551);
or U20100 (N_20100,N_17046,N_16781);
nand U20101 (N_20101,N_17769,N_15767);
nand U20102 (N_20102,N_18647,N_18934);
xnor U20103 (N_20103,N_15988,N_16821);
or U20104 (N_20104,N_19230,N_18191);
xnor U20105 (N_20105,N_17849,N_15995);
or U20106 (N_20106,N_17508,N_16525);
nor U20107 (N_20107,N_19022,N_17168);
or U20108 (N_20108,N_17546,N_16643);
nor U20109 (N_20109,N_18899,N_18726);
nand U20110 (N_20110,N_17107,N_18523);
and U20111 (N_20111,N_16679,N_17104);
or U20112 (N_20112,N_17629,N_16208);
nand U20113 (N_20113,N_18486,N_19167);
or U20114 (N_20114,N_19708,N_17262);
or U20115 (N_20115,N_16811,N_19197);
nor U20116 (N_20116,N_18768,N_19827);
nand U20117 (N_20117,N_15039,N_15934);
or U20118 (N_20118,N_19971,N_15065);
or U20119 (N_20119,N_19067,N_16556);
nand U20120 (N_20120,N_19778,N_19632);
and U20121 (N_20121,N_16375,N_17275);
nand U20122 (N_20122,N_16099,N_19802);
nand U20123 (N_20123,N_15651,N_17854);
nand U20124 (N_20124,N_19846,N_16492);
and U20125 (N_20125,N_18451,N_17186);
or U20126 (N_20126,N_19469,N_15190);
nand U20127 (N_20127,N_17164,N_19329);
and U20128 (N_20128,N_19973,N_19515);
nand U20129 (N_20129,N_16886,N_15814);
and U20130 (N_20130,N_18274,N_16215);
and U20131 (N_20131,N_18742,N_19186);
nand U20132 (N_20132,N_16130,N_18764);
nor U20133 (N_20133,N_18998,N_18655);
nand U20134 (N_20134,N_19202,N_17547);
nor U20135 (N_20135,N_16039,N_16471);
or U20136 (N_20136,N_15072,N_15509);
nand U20137 (N_20137,N_15913,N_15773);
nor U20138 (N_20138,N_17606,N_19033);
nor U20139 (N_20139,N_17529,N_19351);
and U20140 (N_20140,N_16437,N_15038);
xor U20141 (N_20141,N_18149,N_15243);
or U20142 (N_20142,N_16956,N_16873);
and U20143 (N_20143,N_15318,N_16533);
or U20144 (N_20144,N_18125,N_15894);
nor U20145 (N_20145,N_15099,N_18627);
nand U20146 (N_20146,N_15153,N_19925);
nor U20147 (N_20147,N_18813,N_18057);
xor U20148 (N_20148,N_17933,N_15275);
nand U20149 (N_20149,N_18923,N_18392);
nor U20150 (N_20150,N_16286,N_18250);
or U20151 (N_20151,N_18953,N_19438);
nor U20152 (N_20152,N_17634,N_17057);
xor U20153 (N_20153,N_16859,N_18734);
nor U20154 (N_20154,N_15950,N_18044);
xor U20155 (N_20155,N_18491,N_18403);
nand U20156 (N_20156,N_15866,N_15455);
or U20157 (N_20157,N_17489,N_19058);
and U20158 (N_20158,N_18612,N_18183);
nand U20159 (N_20159,N_17803,N_15782);
nand U20160 (N_20160,N_16808,N_15128);
nand U20161 (N_20161,N_17841,N_19024);
xor U20162 (N_20162,N_18283,N_16405);
or U20163 (N_20163,N_18912,N_18897);
and U20164 (N_20164,N_17288,N_16007);
and U20165 (N_20165,N_15398,N_16919);
nand U20166 (N_20166,N_16252,N_17900);
and U20167 (N_20167,N_19286,N_16692);
and U20168 (N_20168,N_19577,N_16125);
xor U20169 (N_20169,N_16303,N_15091);
nand U20170 (N_20170,N_19341,N_17903);
nor U20171 (N_20171,N_18129,N_17093);
and U20172 (N_20172,N_17731,N_19534);
nand U20173 (N_20173,N_19752,N_16381);
or U20174 (N_20174,N_18939,N_17315);
nand U20175 (N_20175,N_15062,N_15966);
and U20176 (N_20176,N_18985,N_16984);
xnor U20177 (N_20177,N_19235,N_15074);
and U20178 (N_20178,N_17603,N_18871);
nor U20179 (N_20179,N_17272,N_15562);
or U20180 (N_20180,N_15536,N_17694);
and U20181 (N_20181,N_15628,N_17054);
xnor U20182 (N_20182,N_15365,N_18851);
and U20183 (N_20183,N_17209,N_17276);
xor U20184 (N_20184,N_19531,N_19527);
xnor U20185 (N_20185,N_15832,N_18517);
nor U20186 (N_20186,N_17174,N_16687);
nand U20187 (N_20187,N_17886,N_17190);
nand U20188 (N_20188,N_18059,N_15159);
xor U20189 (N_20189,N_19903,N_18494);
and U20190 (N_20190,N_19620,N_15273);
nand U20191 (N_20191,N_16973,N_19715);
and U20192 (N_20192,N_15103,N_17306);
and U20193 (N_20193,N_15648,N_17779);
or U20194 (N_20194,N_16646,N_17340);
nor U20195 (N_20195,N_19733,N_17586);
nand U20196 (N_20196,N_15681,N_15361);
nand U20197 (N_20197,N_19754,N_16227);
nand U20198 (N_20198,N_17085,N_16674);
or U20199 (N_20199,N_15104,N_18549);
nand U20200 (N_20200,N_17053,N_19445);
and U20201 (N_20201,N_19786,N_17532);
nand U20202 (N_20202,N_19453,N_15075);
or U20203 (N_20203,N_19625,N_15801);
or U20204 (N_20204,N_19301,N_16657);
nand U20205 (N_20205,N_18385,N_18436);
nand U20206 (N_20206,N_15376,N_16779);
nand U20207 (N_20207,N_16320,N_17239);
and U20208 (N_20208,N_17250,N_19141);
nand U20209 (N_20209,N_15886,N_15984);
or U20210 (N_20210,N_15750,N_15108);
nand U20211 (N_20211,N_19201,N_16926);
xnor U20212 (N_20212,N_16898,N_16837);
or U20213 (N_20213,N_16199,N_17359);
nand U20214 (N_20214,N_15212,N_17060);
and U20215 (N_20215,N_15557,N_18863);
nand U20216 (N_20216,N_17335,N_19129);
nor U20217 (N_20217,N_15483,N_19711);
nand U20218 (N_20218,N_15541,N_17047);
nand U20219 (N_20219,N_15486,N_16520);
or U20220 (N_20220,N_18587,N_18744);
nand U20221 (N_20221,N_17902,N_18807);
xnor U20222 (N_20222,N_15823,N_19251);
or U20223 (N_20223,N_19838,N_16272);
nor U20224 (N_20224,N_17863,N_17191);
nor U20225 (N_20225,N_16183,N_15819);
or U20226 (N_20226,N_17304,N_15513);
or U20227 (N_20227,N_16983,N_15555);
nand U20228 (N_20228,N_15446,N_16587);
nor U20229 (N_20229,N_19709,N_19358);
or U20230 (N_20230,N_15539,N_16670);
nor U20231 (N_20231,N_18381,N_15315);
nand U20232 (N_20232,N_19163,N_16596);
nor U20233 (N_20233,N_16051,N_15058);
nor U20234 (N_20234,N_16672,N_19419);
or U20235 (N_20235,N_17237,N_18121);
nor U20236 (N_20236,N_17836,N_15860);
and U20237 (N_20237,N_18172,N_16876);
xnor U20238 (N_20238,N_15342,N_18586);
nor U20239 (N_20239,N_16551,N_17358);
and U20240 (N_20240,N_15107,N_18783);
and U20241 (N_20241,N_16884,N_17459);
nor U20242 (N_20242,N_17789,N_17349);
nor U20243 (N_20243,N_17762,N_19983);
nand U20244 (N_20244,N_18509,N_15919);
nor U20245 (N_20245,N_16394,N_18193);
or U20246 (N_20246,N_16961,N_17638);
nor U20247 (N_20247,N_16091,N_18520);
xor U20248 (N_20248,N_15267,N_15185);
xor U20249 (N_20249,N_15864,N_15410);
and U20250 (N_20250,N_16085,N_19513);
nor U20251 (N_20251,N_15291,N_17757);
or U20252 (N_20252,N_15904,N_17919);
nor U20253 (N_20253,N_15122,N_16554);
or U20254 (N_20254,N_19421,N_19505);
nor U20255 (N_20255,N_19415,N_15090);
nand U20256 (N_20256,N_19208,N_19641);
or U20257 (N_20257,N_18424,N_19935);
nand U20258 (N_20258,N_19011,N_19958);
nand U20259 (N_20259,N_16621,N_15770);
nor U20260 (N_20260,N_19907,N_18574);
and U20261 (N_20261,N_19747,N_17745);
nor U20262 (N_20262,N_19145,N_17950);
and U20263 (N_20263,N_15269,N_17535);
nand U20264 (N_20264,N_19743,N_17160);
nor U20265 (N_20265,N_19342,N_16511);
nor U20266 (N_20266,N_16680,N_17228);
or U20267 (N_20267,N_17523,N_18235);
and U20268 (N_20268,N_18521,N_18104);
or U20269 (N_20269,N_18463,N_17741);
nand U20270 (N_20270,N_18262,N_18833);
nand U20271 (N_20271,N_17647,N_18358);
nand U20272 (N_20272,N_15493,N_15355);
xnor U20273 (N_20273,N_17596,N_19676);
xnor U20274 (N_20274,N_19370,N_19439);
and U20275 (N_20275,N_15925,N_16359);
and U20276 (N_20276,N_16046,N_15000);
and U20277 (N_20277,N_15730,N_16757);
and U20278 (N_20278,N_19858,N_17435);
or U20279 (N_20279,N_17067,N_17777);
nand U20280 (N_20280,N_15045,N_17485);
and U20281 (N_20281,N_18961,N_18759);
nand U20282 (N_20282,N_18747,N_19442);
nor U20283 (N_20283,N_18921,N_16855);
or U20284 (N_20284,N_15635,N_19290);
or U20285 (N_20285,N_18838,N_19356);
and U20286 (N_20286,N_17370,N_15161);
and U20287 (N_20287,N_15353,N_18093);
nand U20288 (N_20288,N_18665,N_16794);
and U20289 (N_20289,N_18800,N_19714);
or U20290 (N_20290,N_18927,N_17312);
nor U20291 (N_20291,N_16964,N_17087);
or U20292 (N_20292,N_18885,N_19956);
or U20293 (N_20293,N_19690,N_15392);
or U20294 (N_20294,N_19928,N_16610);
nor U20295 (N_20295,N_16463,N_18308);
nor U20296 (N_20296,N_17328,N_16349);
or U20297 (N_20297,N_16311,N_19680);
or U20298 (N_20298,N_16531,N_16369);
nor U20299 (N_20299,N_15765,N_16231);
nand U20300 (N_20300,N_16688,N_15031);
or U20301 (N_20301,N_16421,N_16496);
and U20302 (N_20302,N_17280,N_18307);
and U20303 (N_20303,N_15462,N_16897);
nand U20304 (N_20304,N_16999,N_16947);
nand U20305 (N_20305,N_16974,N_19600);
nor U20306 (N_20306,N_15689,N_17940);
and U20307 (N_20307,N_17357,N_19930);
nand U20308 (N_20308,N_16719,N_17491);
and U20309 (N_20309,N_16426,N_15333);
nor U20310 (N_20310,N_15716,N_18730);
nand U20311 (N_20311,N_16266,N_18495);
nand U20312 (N_20312,N_15224,N_18369);
xor U20313 (N_20313,N_19918,N_19536);
nand U20314 (N_20314,N_16662,N_18198);
or U20315 (N_20315,N_15727,N_17249);
or U20316 (N_20316,N_17981,N_17808);
xnor U20317 (N_20317,N_18527,N_18414);
and U20318 (N_20318,N_18713,N_19405);
and U20319 (N_20319,N_19798,N_18065);
nand U20320 (N_20320,N_17901,N_16154);
and U20321 (N_20321,N_18364,N_19966);
and U20322 (N_20322,N_19835,N_16251);
and U20323 (N_20323,N_19997,N_17828);
nor U20324 (N_20324,N_16173,N_18061);
xor U20325 (N_20325,N_18383,N_16347);
nor U20326 (N_20326,N_19327,N_16432);
or U20327 (N_20327,N_18556,N_19793);
or U20328 (N_20328,N_18404,N_19042);
xnor U20329 (N_20329,N_16411,N_16615);
and U20330 (N_20330,N_19943,N_19895);
or U20331 (N_20331,N_18666,N_19099);
and U20332 (N_20332,N_15946,N_15210);
nor U20333 (N_20333,N_16379,N_18014);
nor U20334 (N_20334,N_17507,N_19002);
nor U20335 (N_20335,N_15573,N_17610);
nor U20336 (N_20336,N_19307,N_15027);
nor U20337 (N_20337,N_16691,N_19570);
or U20338 (N_20338,N_16913,N_18565);
or U20339 (N_20339,N_16412,N_19744);
nand U20340 (N_20340,N_15593,N_17395);
nand U20341 (N_20341,N_18166,N_16774);
and U20342 (N_20342,N_17213,N_15235);
nor U20343 (N_20343,N_17948,N_16976);
and U20344 (N_20344,N_17602,N_19257);
nor U20345 (N_20345,N_16419,N_17082);
and U20346 (N_20346,N_18762,N_15640);
nor U20347 (N_20347,N_15817,N_16015);
nand U20348 (N_20348,N_16285,N_15985);
nor U20349 (N_20349,N_15976,N_15258);
nand U20350 (N_20350,N_17454,N_16966);
nand U20351 (N_20351,N_17627,N_16380);
or U20352 (N_20352,N_15816,N_18937);
nand U20353 (N_20353,N_16056,N_17545);
or U20354 (N_20354,N_18547,N_15092);
nand U20355 (N_20355,N_15605,N_15588);
nand U20356 (N_20356,N_16539,N_19876);
nor U20357 (N_20357,N_16844,N_19056);
and U20358 (N_20358,N_18711,N_18094);
nand U20359 (N_20359,N_19432,N_18442);
or U20360 (N_20360,N_18047,N_19111);
or U20361 (N_20361,N_16850,N_18880);
or U20362 (N_20362,N_17908,N_17063);
nand U20363 (N_20363,N_17230,N_17582);
nand U20364 (N_20364,N_18092,N_19345);
and U20365 (N_20365,N_18366,N_16290);
nand U20366 (N_20366,N_16348,N_15245);
and U20367 (N_20367,N_15967,N_18461);
nand U20368 (N_20368,N_16198,N_19554);
nor U20369 (N_20369,N_17319,N_16701);
or U20370 (N_20370,N_17193,N_16737);
nand U20371 (N_20371,N_19659,N_18237);
nand U20372 (N_20372,N_19678,N_18236);
nand U20373 (N_20373,N_17826,N_18096);
xor U20374 (N_20374,N_15013,N_17562);
or U20375 (N_20375,N_17804,N_17221);
nand U20376 (N_20376,N_15587,N_18470);
or U20377 (N_20377,N_16392,N_15563);
and U20378 (N_20378,N_17955,N_18702);
nor U20379 (N_20379,N_19774,N_16676);
and U20380 (N_20380,N_15930,N_16281);
and U20381 (N_20381,N_17450,N_15880);
and U20382 (N_20382,N_19146,N_19520);
or U20383 (N_20383,N_17317,N_17163);
or U20384 (N_20384,N_19599,N_19539);
nor U20385 (N_20385,N_17853,N_15179);
and U20386 (N_20386,N_19948,N_18258);
or U20387 (N_20387,N_18192,N_19053);
and U20388 (N_20388,N_16212,N_19396);
and U20389 (N_20389,N_15599,N_19607);
nor U20390 (N_20390,N_19325,N_19249);
or U20391 (N_20391,N_18652,N_19551);
and U20392 (N_20392,N_17464,N_16371);
nor U20393 (N_20393,N_19522,N_17162);
xnor U20394 (N_20394,N_17265,N_17271);
and U20395 (N_20395,N_18071,N_16237);
nand U20396 (N_20396,N_16295,N_15592);
and U20397 (N_20397,N_17023,N_15134);
nor U20398 (N_20398,N_18834,N_16766);
xnor U20399 (N_20399,N_15786,N_15066);
nor U20400 (N_20400,N_15920,N_17720);
nor U20401 (N_20401,N_18602,N_17279);
nand U20402 (N_20402,N_15182,N_16761);
and U20403 (N_20403,N_15690,N_18216);
or U20404 (N_20404,N_19223,N_19265);
or U20405 (N_20405,N_16078,N_15533);
nand U20406 (N_20406,N_18878,N_16684);
and U20407 (N_20407,N_19565,N_16324);
nor U20408 (N_20408,N_16936,N_16072);
or U20409 (N_20409,N_15676,N_19999);
and U20410 (N_20410,N_16865,N_17921);
nand U20411 (N_20411,N_17716,N_19095);
nand U20412 (N_20412,N_15901,N_15808);
and U20413 (N_20413,N_16819,N_15725);
nor U20414 (N_20414,N_17575,N_19957);
nand U20415 (N_20415,N_19078,N_19110);
xnor U20416 (N_20416,N_19464,N_18393);
xnor U20417 (N_20417,N_17263,N_19961);
or U20418 (N_20418,N_16980,N_16110);
or U20419 (N_20419,N_15325,N_19789);
nor U20420 (N_20420,N_17870,N_15559);
nor U20421 (N_20421,N_15314,N_18203);
nor U20422 (N_20422,N_17469,N_15169);
or U20423 (N_20423,N_19449,N_19380);
or U20424 (N_20424,N_15375,N_15330);
or U20425 (N_20425,N_19691,N_17994);
and U20426 (N_20426,N_16927,N_16929);
and U20427 (N_20427,N_15841,N_19746);
nor U20428 (N_20428,N_17412,N_19123);
or U20429 (N_20429,N_17588,N_19335);
and U20430 (N_20430,N_17300,N_17036);
and U20431 (N_20431,N_19508,N_17897);
nand U20432 (N_20432,N_17765,N_17081);
and U20433 (N_20433,N_17631,N_18089);
xnor U20434 (N_20434,N_19742,N_15465);
nor U20435 (N_20435,N_15222,N_15630);
or U20436 (N_20436,N_19093,N_16230);
or U20437 (N_20437,N_19502,N_17728);
xor U20438 (N_20438,N_15641,N_16438);
nor U20439 (N_20439,N_19074,N_19549);
and U20440 (N_20440,N_17600,N_17909);
nand U20441 (N_20441,N_18330,N_15759);
and U20442 (N_20442,N_17446,N_16699);
nor U20443 (N_20443,N_17194,N_18184);
xor U20444 (N_20444,N_16054,N_16301);
and U20445 (N_20445,N_17356,N_16755);
and U20446 (N_20446,N_18958,N_16875);
or U20447 (N_20447,N_15658,N_17079);
or U20448 (N_20448,N_15263,N_18471);
or U20449 (N_20449,N_19900,N_17855);
or U20450 (N_20450,N_18892,N_18038);
or U20451 (N_20451,N_18991,N_16445);
or U20452 (N_20452,N_18981,N_19564);
nand U20453 (N_20453,N_15220,N_17956);
or U20454 (N_20454,N_16218,N_15526);
nor U20455 (N_20455,N_16476,N_17211);
nor U20456 (N_20456,N_18162,N_15067);
xnor U20457 (N_20457,N_17264,N_17861);
and U20458 (N_20458,N_16970,N_19289);
or U20459 (N_20459,N_19981,N_18368);
xor U20460 (N_20460,N_15132,N_18024);
xor U20461 (N_20461,N_17383,N_19211);
or U20462 (N_20462,N_18968,N_19317);
nand U20463 (N_20463,N_19113,N_15352);
nor U20464 (N_20464,N_16249,N_16705);
nor U20465 (N_20465,N_16446,N_17261);
nand U20466 (N_20466,N_19117,N_19269);
nor U20467 (N_20467,N_18165,N_16627);
nor U20468 (N_20468,N_17455,N_17011);
or U20469 (N_20469,N_16810,N_15824);
nand U20470 (N_20470,N_16002,N_16613);
and U20471 (N_20471,N_18538,N_15116);
nor U20472 (N_20472,N_18941,N_19275);
nand U20473 (N_20473,N_19761,N_18072);
and U20474 (N_20474,N_15802,N_17216);
nand U20475 (N_20475,N_16134,N_15232);
or U20476 (N_20476,N_19114,N_19169);
nor U20477 (N_20477,N_17408,N_19456);
nor U20478 (N_20478,N_16881,N_16618);
nand U20479 (N_20479,N_15532,N_17324);
or U20480 (N_20480,N_19112,N_15769);
nor U20481 (N_20481,N_15804,N_15961);
or U20482 (N_20482,N_18205,N_19812);
or U20483 (N_20483,N_17645,N_16452);
nor U20484 (N_20484,N_16122,N_15124);
or U20485 (N_20485,N_19331,N_17552);
nor U20486 (N_20486,N_18412,N_19982);
nor U20487 (N_20487,N_19283,N_17714);
and U20488 (N_20488,N_16259,N_16343);
and U20489 (N_20489,N_17659,N_17810);
nor U20490 (N_20490,N_16758,N_19817);
and U20491 (N_20491,N_17373,N_19891);
or U20492 (N_20492,N_18737,N_18106);
or U20493 (N_20493,N_19601,N_15496);
nor U20494 (N_20494,N_16542,N_18722);
or U20495 (N_20495,N_16846,N_19751);
or U20496 (N_20496,N_16637,N_16254);
and U20497 (N_20497,N_18137,N_16514);
nor U20498 (N_20498,N_18676,N_16447);
or U20499 (N_20499,N_18896,N_17530);
or U20500 (N_20500,N_19597,N_17198);
nor U20501 (N_20501,N_15618,N_19972);
xor U20502 (N_20502,N_19330,N_17511);
nor U20503 (N_20503,N_19689,N_18700);
or U20504 (N_20504,N_16767,N_15514);
and U20505 (N_20505,N_15088,N_15005);
xor U20506 (N_20506,N_15647,N_16565);
or U20507 (N_20507,N_19149,N_18815);
or U20508 (N_20508,N_19963,N_15677);
and U20509 (N_20509,N_16776,N_15854);
xnor U20510 (N_20510,N_19836,N_19947);
nor U20511 (N_20511,N_16709,N_15233);
nand U20512 (N_20512,N_19702,N_17493);
xor U20513 (N_20513,N_18945,N_17170);
or U20514 (N_20514,N_18035,N_16283);
and U20515 (N_20515,N_15891,N_17549);
nor U20516 (N_20516,N_19189,N_19813);
or U20517 (N_20517,N_15746,N_17608);
nor U20518 (N_20518,N_19021,N_15519);
nand U20519 (N_20519,N_17771,N_18926);
xor U20520 (N_20520,N_18197,N_16345);
and U20521 (N_20521,N_17709,N_19046);
or U20522 (N_20522,N_18097,N_16829);
xor U20523 (N_20523,N_16835,N_15733);
nor U20524 (N_20524,N_18354,N_17813);
or U20525 (N_20525,N_15780,N_16457);
nand U20526 (N_20526,N_16243,N_15244);
xor U20527 (N_20527,N_16989,N_19069);
or U20528 (N_20528,N_18975,N_19267);
nand U20529 (N_20529,N_18820,N_15458);
or U20530 (N_20530,N_19974,N_18150);
nor U20531 (N_20531,N_17831,N_17243);
or U20532 (N_20532,N_16111,N_18518);
and U20533 (N_20533,N_18131,N_18803);
nand U20534 (N_20534,N_16860,N_15678);
and U20535 (N_20535,N_19165,N_15348);
nor U20536 (N_20536,N_15408,N_19444);
or U20537 (N_20537,N_18427,N_19511);
nand U20538 (N_20538,N_17180,N_16096);
nor U20539 (N_20539,N_16226,N_19652);
or U20540 (N_20540,N_16490,N_18614);
nand U20541 (N_20541,N_17411,N_19667);
nand U20542 (N_20542,N_16651,N_19417);
or U20543 (N_20543,N_18534,N_18753);
nand U20544 (N_20544,N_15308,N_17422);
nor U20545 (N_20545,N_18906,N_17114);
nor U20546 (N_20546,N_17460,N_16410);
or U20547 (N_20547,N_18861,N_19596);
and U20548 (N_20548,N_16557,N_15580);
and U20549 (N_20549,N_19583,N_15707);
nor U20550 (N_20550,N_15763,N_15518);
nand U20551 (N_20551,N_18255,N_16076);
nor U20552 (N_20552,N_17403,N_16495);
nand U20553 (N_20553,N_18633,N_15391);
nand U20554 (N_20554,N_16512,N_15540);
nor U20555 (N_20555,N_17787,N_15164);
and U20556 (N_20556,N_18430,N_18501);
xnor U20557 (N_20557,N_15246,N_19132);
or U20558 (N_20558,N_16499,N_15735);
nor U20559 (N_20559,N_15059,N_15848);
or U20560 (N_20560,N_19929,N_17005);
nand U20561 (N_20561,N_16214,N_15550);
nand U20562 (N_20562,N_15168,N_15306);
nand U20563 (N_20563,N_19277,N_18959);
nor U20564 (N_20564,N_19212,N_19825);
or U20565 (N_20565,N_19578,N_19631);
nor U20566 (N_20566,N_19883,N_15418);
and U20567 (N_20567,N_18819,N_17740);
nor U20568 (N_20568,N_19579,N_18770);
and U20569 (N_20569,N_15299,N_16477);
nand U20570 (N_20570,N_18238,N_18752);
or U20571 (N_20571,N_18624,N_15449);
and U20572 (N_20572,N_15111,N_17123);
or U20573 (N_20573,N_16711,N_17345);
and U20574 (N_20574,N_18876,N_17429);
xnor U20575 (N_20575,N_15929,N_19102);
xnor U20576 (N_20576,N_18832,N_19363);
nor U20577 (N_20577,N_15638,N_16792);
and U20578 (N_20578,N_16304,N_15397);
and U20579 (N_20579,N_19416,N_19575);
nor U20580 (N_20580,N_18589,N_16784);
xnor U20581 (N_20581,N_18847,N_19284);
nor U20582 (N_20582,N_18936,N_16487);
nand U20583 (N_20583,N_17303,N_18003);
or U20584 (N_20584,N_15345,N_19729);
xnor U20585 (N_20585,N_18472,N_17374);
or U20586 (N_20586,N_19035,N_19898);
xnor U20587 (N_20587,N_19657,N_19576);
nor U20588 (N_20588,N_16965,N_17027);
and U20589 (N_20589,N_19845,N_19855);
or U20590 (N_20590,N_16544,N_19862);
and U20591 (N_20591,N_19787,N_16202);
or U20592 (N_20592,N_15283,N_15902);
xnor U20593 (N_20593,N_17154,N_17031);
and U20594 (N_20594,N_15024,N_19306);
or U20595 (N_20595,N_15922,N_19081);
nor U20596 (N_20596,N_17817,N_18467);
and U20597 (N_20597,N_16738,N_18693);
or U20598 (N_20598,N_19460,N_19716);
and U20599 (N_20599,N_16753,N_18305);
or U20600 (N_20600,N_19362,N_18454);
or U20601 (N_20601,N_15251,N_17792);
xor U20602 (N_20602,N_15015,N_17254);
nand U20603 (N_20603,N_19500,N_17166);
or U20604 (N_20604,N_15130,N_16723);
or U20605 (N_20605,N_15225,N_15173);
xor U20606 (N_20606,N_17431,N_15019);
xnor U20607 (N_20607,N_18306,N_19366);
xor U20608 (N_20608,N_15044,N_15692);
and U20609 (N_20609,N_18111,N_19645);
and U20610 (N_20610,N_17376,N_17483);
and U20611 (N_20611,N_19246,N_18365);
nor U20612 (N_20612,N_16184,N_18609);
and U20613 (N_20613,N_17492,N_19964);
xnor U20614 (N_20614,N_19668,N_19232);
and U20615 (N_20615,N_18729,N_17895);
nand U20616 (N_20616,N_18450,N_15619);
and U20617 (N_20617,N_19382,N_19470);
nand U20618 (N_20618,N_18304,N_18037);
nor U20619 (N_20619,N_19848,N_18887);
nor U20620 (N_20620,N_19717,N_17975);
nand U20621 (N_20621,N_17543,N_15419);
nand U20622 (N_20622,N_18716,N_18018);
and U20623 (N_20623,N_15368,N_18708);
and U20624 (N_20624,N_15278,N_16635);
and U20625 (N_20625,N_19017,N_19504);
or U20626 (N_20626,N_15600,N_18139);
xor U20627 (N_20627,N_15311,N_15734);
nand U20628 (N_20628,N_17963,N_19905);
xor U20629 (N_20629,N_18043,N_17208);
nor U20630 (N_20630,N_18888,N_15217);
or U20631 (N_20631,N_16942,N_15320);
and U20632 (N_20632,N_17815,N_19350);
nor U20633 (N_20633,N_18914,N_16194);
nor U20634 (N_20634,N_15608,N_17430);
nor U20635 (N_20635,N_19650,N_15319);
nand U20636 (N_20636,N_15457,N_19940);
or U20637 (N_20637,N_15811,N_19244);
nand U20638 (N_20638,N_17313,N_19750);
and U20639 (N_20639,N_16567,N_17465);
nor U20640 (N_20640,N_16242,N_19661);
xnor U20641 (N_20641,N_16697,N_15788);
and U20642 (N_20642,N_19378,N_15433);
or U20643 (N_20643,N_16485,N_16741);
or U20644 (N_20644,N_17480,N_18473);
nor U20645 (N_20645,N_19840,N_17476);
xor U20646 (N_20646,N_16024,N_17028);
xnor U20647 (N_20647,N_19766,N_16036);
or U20648 (N_20648,N_15080,N_17297);
or U20649 (N_20649,N_15505,N_15036);
and U20650 (N_20650,N_17516,N_18970);
nand U20651 (N_20651,N_16474,N_15203);
nor U20652 (N_20652,N_18388,N_18146);
nand U20653 (N_20653,N_16402,N_15545);
xnor U20654 (N_20654,N_15156,N_19180);
nand U20655 (N_20655,N_15176,N_18377);
nor U20656 (N_20656,N_19685,N_17743);
nand U20657 (N_20657,N_17871,N_17220);
nand U20658 (N_20658,N_16772,N_19734);
xnor U20659 (N_20659,N_16883,N_18775);
or U20660 (N_20660,N_15622,N_16949);
nor U20661 (N_20661,N_18134,N_16486);
and U20662 (N_20662,N_16997,N_15959);
xor U20663 (N_20663,N_19218,N_17661);
or U20664 (N_20664,N_18830,N_18706);
xnor U20665 (N_20665,N_15719,N_16287);
or U20666 (N_20666,N_17010,N_18592);
nand U20667 (N_20667,N_15525,N_17913);
nor U20668 (N_20668,N_15907,N_19901);
and U20669 (N_20669,N_16484,N_15583);
or U20670 (N_20670,N_15478,N_15501);
or U20671 (N_20671,N_15052,N_17917);
and U20672 (N_20672,N_18384,N_15442);
and U20673 (N_20673,N_15893,N_16097);
nor U20674 (N_20674,N_17601,N_19466);
nor U20675 (N_20675,N_15004,N_15118);
nor U20676 (N_20676,N_15010,N_19931);
nor U20677 (N_20677,N_16466,N_16291);
nor U20678 (N_20678,N_19850,N_16169);
xnor U20679 (N_20679,N_17730,N_18079);
nand U20680 (N_20680,N_16357,N_17103);
nand U20681 (N_20681,N_18772,N_15631);
nand U20682 (N_20682,N_18133,N_18661);
and U20683 (N_20683,N_16820,N_15827);
nand U20684 (N_20684,N_18854,N_16423);
and U20685 (N_20685,N_19538,N_17781);
nand U20686 (N_20686,N_15369,N_15850);
nand U20687 (N_20687,N_18606,N_19209);
or U20688 (N_20688,N_15793,N_16494);
and U20689 (N_20689,N_16752,N_18850);
nand U20690 (N_20690,N_15791,N_15684);
nor U20691 (N_20691,N_19624,N_17088);
and U20692 (N_20692,N_17353,N_17287);
nand U20693 (N_20693,N_17066,N_17615);
nand U20694 (N_20694,N_17859,N_19192);
or U20695 (N_20695,N_18504,N_16972);
and U20696 (N_20696,N_17077,N_19261);
nor U20697 (N_20697,N_16649,N_17628);
and U20698 (N_20698,N_18884,N_18425);
nor U20699 (N_20699,N_17996,N_15851);
or U20700 (N_20700,N_16622,N_18199);
and U20701 (N_20701,N_17334,N_16659);
nor U20702 (N_20702,N_19343,N_19150);
nor U20703 (N_20703,N_15479,N_17482);
and U20704 (N_20704,N_18584,N_19871);
or U20705 (N_20705,N_19448,N_16827);
nand U20706 (N_20706,N_15194,N_15842);
and U20707 (N_20707,N_15771,N_19373);
nor U20708 (N_20708,N_19133,N_15249);
and U20709 (N_20709,N_18848,N_17832);
or U20710 (N_20710,N_18405,N_15524);
or U20711 (N_20711,N_18546,N_17248);
nor U20712 (N_20712,N_17528,N_19731);
and U20713 (N_20713,N_18053,N_17674);
nor U20714 (N_20714,N_17542,N_19227);
nor U20715 (N_20715,N_19605,N_17522);
and U20716 (N_20716,N_19833,N_17121);
and U20717 (N_20717,N_16853,N_17326);
and U20718 (N_20718,N_17096,N_18797);
or U20719 (N_20719,N_16880,N_17069);
nand U20720 (N_20720,N_18416,N_17205);
and U20721 (N_20721,N_18535,N_19319);
xor U20722 (N_20722,N_16205,N_17509);
or U20723 (N_20723,N_16147,N_17434);
and U20724 (N_20724,N_18761,N_19034);
nor U20725 (N_20725,N_16167,N_19302);
xnor U20726 (N_20726,N_16455,N_18479);
xnor U20727 (N_20727,N_18039,N_18705);
nor U20728 (N_20728,N_19516,N_16937);
nor U20729 (N_20729,N_16316,N_18558);
nand U20730 (N_20730,N_17158,N_19673);
and U20731 (N_20731,N_15853,N_17165);
nand U20732 (N_20732,N_15412,N_16872);
nand U20733 (N_20733,N_16607,N_16830);
nor U20734 (N_20734,N_15666,N_15077);
or U20735 (N_20735,N_16459,N_16161);
or U20736 (N_20736,N_17710,N_17461);
xor U20737 (N_20737,N_19326,N_16895);
nand U20738 (N_20738,N_18751,N_16793);
nand U20739 (N_20739,N_17844,N_18312);
nor U20740 (N_20740,N_15507,N_17864);
or U20741 (N_20741,N_15882,N_19899);
xor U20742 (N_20742,N_18605,N_19792);
xnor U20743 (N_20743,N_15991,N_18386);
xnor U20744 (N_20744,N_19921,N_18278);
nor U20745 (N_20745,N_16770,N_19160);
and U20746 (N_20746,N_15710,N_15553);
xor U20747 (N_20747,N_17712,N_18194);
nand U20748 (N_20748,N_15779,N_15441);
and U20749 (N_20749,N_18625,N_18901);
nand U20750 (N_20750,N_15713,N_19591);
or U20751 (N_20751,N_16922,N_15965);
nand U20752 (N_20752,N_16906,N_17969);
and U20753 (N_20753,N_17515,N_17576);
or U20754 (N_20754,N_15937,N_17080);
xor U20755 (N_20755,N_15564,N_18767);
nand U20756 (N_20756,N_15888,N_15172);
or U20757 (N_20757,N_19364,N_17640);
nand U20758 (N_20758,N_17468,N_18810);
nand U20759 (N_20759,N_15476,N_15900);
xnor U20760 (N_20760,N_19248,N_16902);
or U20761 (N_20761,N_16247,N_17229);
xor U20762 (N_20762,N_16307,N_18785);
and U20763 (N_20763,N_17887,N_19153);
and U20764 (N_20764,N_19476,N_17100);
nor U20765 (N_20765,N_17409,N_15910);
and U20766 (N_20766,N_18391,N_19478);
and U20767 (N_20767,N_17993,N_19990);
nor U20768 (N_20768,N_15790,N_18110);
and U20769 (N_20769,N_15060,N_19634);
or U20770 (N_20770,N_15796,N_19126);
and U20771 (N_20771,N_15679,N_17819);
and U20772 (N_20772,N_19927,N_15056);
and U20773 (N_20773,N_15974,N_19352);
xnor U20774 (N_20774,N_19161,N_19424);
and U20775 (N_20775,N_15189,N_19736);
nand U20776 (N_20776,N_18511,N_19867);
xor U20777 (N_20777,N_16433,N_17266);
xnor U20778 (N_20778,N_17591,N_19799);
or U20779 (N_20779,N_19945,N_16867);
nor U20780 (N_20780,N_15183,N_19305);
xnor U20781 (N_20781,N_16632,N_18786);
nor U20782 (N_20782,N_15905,N_15223);
or U20783 (N_20783,N_15783,N_15467);
and U20784 (N_20784,N_19910,N_19572);
nor U20785 (N_20785,N_18006,N_17389);
xor U20786 (N_20786,N_17330,N_15034);
nand U20787 (N_20787,N_16717,N_16127);
or U20788 (N_20788,N_18294,N_19671);
nand U20789 (N_20789,N_17307,N_16150);
and U20790 (N_20790,N_16745,N_15862);
nand U20791 (N_20791,N_19237,N_15821);
or U20792 (N_20792,N_17845,N_16269);
or U20793 (N_20793,N_15197,N_19440);
nand U20794 (N_20794,N_15589,N_16958);
nor U20795 (N_20795,N_17478,N_15731);
nor U20796 (N_20796,N_16203,N_15326);
xnor U20797 (N_20797,N_16488,N_16050);
xnor U20798 (N_20798,N_19627,N_16264);
nand U20799 (N_20799,N_17466,N_15008);
nand U20800 (N_20800,N_16465,N_18550);
nor U20801 (N_20801,N_19839,N_19801);
nand U20802 (N_20802,N_19418,N_17043);
or U20803 (N_20803,N_16177,N_15825);
nand U20804 (N_20804,N_16732,N_18052);
or U20805 (N_20805,N_19065,N_16744);
nor U20806 (N_20806,N_18220,N_16944);
or U20807 (N_20807,N_16534,N_18575);
and U20808 (N_20808,N_16467,N_17574);
and U20809 (N_20809,N_17884,N_18357);
or U20810 (N_20810,N_15415,N_17061);
and U20811 (N_20811,N_17892,N_16441);
and U20812 (N_20812,N_15781,N_17497);
nor U20813 (N_20813,N_18362,N_16460);
nor U20814 (N_20814,N_16378,N_18682);
or U20815 (N_20815,N_16892,N_18545);
nor U20816 (N_20816,N_16142,N_16991);
nand U20817 (N_20817,N_17814,N_16258);
nor U20818 (N_20818,N_19003,N_15815);
xor U20819 (N_20819,N_16735,N_18977);
nor U20820 (N_20820,N_19392,N_17526);
nand U20821 (N_20821,N_18685,N_17512);
or U20822 (N_20822,N_16284,N_17417);
nor U20823 (N_20823,N_15294,N_17184);
nand U20824 (N_20824,N_16322,N_19279);
and U20825 (N_20825,N_18516,N_16720);
nand U20826 (N_20826,N_18173,N_17687);
and U20827 (N_20827,N_19699,N_15818);
or U20828 (N_20828,N_17504,N_19558);
or U20829 (N_20829,N_17559,N_16959);
nand U20830 (N_20830,N_15953,N_16510);
and U20831 (N_20831,N_18023,N_16953);
nand U20832 (N_20832,N_15949,N_16592);
or U20833 (N_20833,N_19749,N_18108);
nand U20834 (N_20834,N_16787,N_19915);
and U20835 (N_20835,N_16417,N_19610);
xor U20836 (N_20836,N_16361,N_16005);
nor U20837 (N_20837,N_18204,N_15548);
and U20838 (N_20838,N_15696,N_18314);
nand U20839 (N_20839,N_15312,N_18440);
or U20840 (N_20840,N_16868,N_15136);
nor U20841 (N_20841,N_19321,N_19805);
and U20842 (N_20842,N_19049,N_18174);
or U20843 (N_20843,N_15270,N_19347);
nor U20844 (N_20844,N_17748,N_15906);
or U20845 (N_20845,N_16568,N_15865);
xor U20846 (N_20846,N_19276,N_17109);
nor U20847 (N_20847,N_18328,N_16031);
xor U20848 (N_20848,N_17355,N_19333);
nor U20849 (N_20849,N_18313,N_17879);
nor U20850 (N_20850,N_15617,N_18646);
or U20851 (N_20851,N_18206,N_19051);
and U20852 (N_20852,N_15627,N_19340);
nor U20853 (N_20853,N_18144,N_18648);
nor U20854 (N_20854,N_18673,N_19630);
or U20855 (N_20855,N_18468,N_16483);
nor U20856 (N_20856,N_18567,N_16546);
nand U20857 (N_20857,N_19474,N_15899);
xor U20858 (N_20858,N_16882,N_18297);
nor U20859 (N_20859,N_19759,N_17827);
nor U20860 (N_20860,N_16413,N_19696);
nor U20861 (N_20861,N_19188,N_16093);
and U20862 (N_20862,N_18159,N_17846);
nor U20863 (N_20863,N_15646,N_15171);
and U20864 (N_20864,N_15924,N_19296);
or U20865 (N_20865,N_16278,N_15911);
or U20866 (N_20866,N_16903,N_18859);
or U20867 (N_20867,N_16756,N_19528);
nor U20868 (N_20868,N_18724,N_19991);
nor U20869 (N_20869,N_17225,N_16235);
and U20870 (N_20870,N_18882,N_17392);
nand U20871 (N_20871,N_16552,N_17669);
nor U20872 (N_20872,N_18374,N_17044);
xor U20873 (N_20873,N_19540,N_17569);
or U20874 (N_20874,N_17891,N_15542);
nand U20875 (N_20875,N_17783,N_18485);
nand U20876 (N_20876,N_18662,N_17382);
nand U20877 (N_20877,N_17928,N_18823);
or U20878 (N_20878,N_16299,N_17030);
nand U20879 (N_20879,N_16677,N_16448);
nand U20880 (N_20880,N_19563,N_18678);
or U20881 (N_20881,N_19441,N_17311);
nor U20882 (N_20882,N_15135,N_15761);
nor U20883 (N_20883,N_18063,N_17727);
and U20884 (N_20884,N_19323,N_19410);
nand U20885 (N_20885,N_18041,N_17073);
nor U20886 (N_20886,N_18582,N_15076);
xnor U20887 (N_20887,N_15289,N_18654);
or U20888 (N_20888,N_18382,N_15322);
nor U20889 (N_20889,N_18227,N_19219);
and U20890 (N_20890,N_17413,N_17679);
nor U20891 (N_20891,N_18733,N_16336);
and U20892 (N_20892,N_15175,N_17014);
and U20893 (N_20893,N_17553,N_16731);
or U20894 (N_20894,N_15337,N_17557);
nor U20895 (N_20895,N_17078,N_17344);
and U20896 (N_20896,N_15502,N_19735);
nor U20897 (N_20897,N_15166,N_19338);
nand U20898 (N_20898,N_15279,N_17354);
and U20899 (N_20899,N_18074,N_19636);
and U20900 (N_20900,N_17943,N_15872);
nand U20901 (N_20901,N_17579,N_15238);
nand U20902 (N_20902,N_15983,N_19185);
xnor U20903 (N_20903,N_16832,N_16453);
nand U20904 (N_20904,N_15234,N_17032);
nand U20905 (N_20905,N_19052,N_19581);
nor U20906 (N_20906,N_15624,N_15282);
or U20907 (N_20907,N_18608,N_18686);
and U20908 (N_20908,N_18017,N_16323);
and U20909 (N_20909,N_19841,N_15797);
and U20910 (N_20910,N_19303,N_17724);
nand U20911 (N_20911,N_16149,N_15803);
nor U20912 (N_20912,N_16306,N_19626);
and U20913 (N_20913,N_17232,N_16121);
nor U20914 (N_20914,N_19767,N_19791);
nor U20915 (N_20915,N_19250,N_19446);
nor U20916 (N_20916,N_19459,N_16095);
nor U20917 (N_20917,N_17977,N_18573);
nand U20918 (N_20918,N_15682,N_17663);
and U20919 (N_20919,N_15359,N_15354);
nor U20920 (N_20920,N_17099,N_18356);
xnor U20921 (N_20921,N_16302,N_15921);
nand U20922 (N_20922,N_15158,N_15316);
or U20923 (N_20923,N_18157,N_18230);
nand U20924 (N_20924,N_17233,N_18963);
or U20925 (N_20925,N_19006,N_19014);
and U20926 (N_20926,N_18275,N_16367);
xnor U20927 (N_20927,N_19196,N_17944);
and U20928 (N_20928,N_16312,N_17915);
or U20929 (N_20929,N_19609,N_15659);
nand U20930 (N_20930,N_15523,N_18852);
and U20931 (N_20931,N_18400,N_16089);
or U20932 (N_20932,N_19015,N_18212);
nand U20933 (N_20933,N_16905,N_15277);
xor U20934 (N_20934,N_17785,N_19486);
nor U20935 (N_20935,N_19007,N_19116);
and U20936 (N_20936,N_17682,N_16934);
or U20937 (N_20937,N_17390,N_19737);
nand U20938 (N_20938,N_17420,N_16373);
or U20939 (N_20939,N_15049,N_18793);
xor U20940 (N_20940,N_16620,N_16425);
nand U20941 (N_20941,N_15471,N_16363);
nor U20942 (N_20942,N_18746,N_19496);
and U20943 (N_20943,N_19954,N_16275);
and U20944 (N_20944,N_15372,N_17842);
nand U20945 (N_20945,N_17337,N_19295);
xor U20946 (N_20946,N_18343,N_16225);
xor U20947 (N_20947,N_17428,N_15652);
nand U20948 (N_20948,N_16444,N_19887);
xnor U20949 (N_20949,N_17185,N_15002);
xor U20950 (N_20950,N_19675,N_15503);
or U20951 (N_20951,N_18642,N_18156);
and U20952 (N_20952,N_17075,N_18459);
xor U20953 (N_20953,N_18080,N_18272);
or U20954 (N_20954,N_15789,N_15405);
and U20955 (N_20955,N_19142,N_15364);
nor U20956 (N_20956,N_15150,N_18635);
nand U20957 (N_20957,N_15680,N_19262);
nand U20958 (N_20958,N_16190,N_16308);
nand U20959 (N_20959,N_18273,N_17999);
nor U20960 (N_20960,N_16981,N_18415);
nor U20961 (N_20961,N_17677,N_15157);
nor U20962 (N_20962,N_19885,N_15611);
nand U20963 (N_20963,N_19875,N_16858);
and U20964 (N_20964,N_15068,N_18736);
nor U20965 (N_20965,N_17277,N_16368);
nand U20966 (N_20966,N_16967,N_17135);
or U20967 (N_20967,N_17404,N_19986);
xnor U20968 (N_20968,N_17204,N_15812);
nand U20969 (N_20969,N_16912,N_15009);
and U20970 (N_20970,N_16751,N_18084);
nand U20971 (N_20971,N_17865,N_19880);
and U20972 (N_20972,N_17234,N_19660);
nor U20973 (N_20973,N_16049,N_16780);
or U20974 (N_20974,N_18141,N_17505);
nor U20975 (N_20975,N_15098,N_17816);
xor U20976 (N_20976,N_15952,N_17336);
nor U20977 (N_20977,N_18943,N_16132);
nand U20978 (N_20978,N_18801,N_18152);
nor U20979 (N_20979,N_18644,N_17990);
xnor U20980 (N_20980,N_15561,N_15990);
and U20981 (N_20981,N_18809,N_19001);
nor U20982 (N_20982,N_16480,N_18630);
or U20983 (N_20983,N_17690,N_15163);
nor U20984 (N_20984,N_19243,N_18143);
and U20985 (N_20985,N_16270,N_18571);
nor U20986 (N_20986,N_17361,N_17501);
nand U20987 (N_20987,N_19407,N_19374);
xor U20988 (N_20988,N_16995,N_19371);
nor U20989 (N_20989,N_16569,N_16029);
and U20990 (N_20990,N_15014,N_15199);
nand U20991 (N_20991,N_18542,N_16473);
nor U20992 (N_20992,N_16653,N_15055);
and U20993 (N_20993,N_15491,N_17825);
or U20994 (N_20994,N_19454,N_17695);
and U20995 (N_20995,N_18554,N_15046);
and U20996 (N_20996,N_15849,N_16931);
or U20997 (N_20997,N_15003,N_18905);
and U20998 (N_20998,N_16690,N_18101);
and U20999 (N_20999,N_15954,N_19904);
nor U21000 (N_21000,N_18723,N_15942);
or U21001 (N_21001,N_16219,N_16536);
or U21002 (N_21002,N_18596,N_17754);
or U21003 (N_21003,N_15538,N_19806);
or U21004 (N_21004,N_16059,N_17747);
or U21005 (N_21005,N_19450,N_19765);
or U21006 (N_21006,N_17936,N_15728);
and U21007 (N_21007,N_16543,N_19688);
or U21008 (N_21008,N_17172,N_15450);
or U21009 (N_21009,N_18808,N_18514);
or U21010 (N_21010,N_18107,N_16518);
nand U21011 (N_21011,N_17766,N_15029);
or U21012 (N_21012,N_17982,N_17688);
and U21013 (N_21013,N_18413,N_19134);
and U21014 (N_21014,N_17343,N_18831);
or U21015 (N_21015,N_18098,N_16532);
xor U21016 (N_21016,N_16245,N_17017);
nand U21017 (N_21017,N_16600,N_18720);
nand U21018 (N_21018,N_18302,N_17834);
nor U21019 (N_21019,N_16156,N_15451);
nor U21020 (N_21020,N_16938,N_15256);
and U21021 (N_21021,N_19861,N_15537);
or U21022 (N_21022,N_18869,N_19233);
or U21023 (N_21023,N_19048,N_18949);
nor U21024 (N_21024,N_19782,N_16939);
or U21025 (N_21025,N_18251,N_16502);
or U21026 (N_21026,N_16458,N_17656);
or U21027 (N_21027,N_19823,N_17732);
and U21028 (N_21028,N_15070,N_19187);
and U21029 (N_21029,N_17432,N_16769);
or U21030 (N_21030,N_15633,N_17672);
or U21031 (N_21031,N_15293,N_18016);
or U21032 (N_21032,N_16739,N_15469);
and U21033 (N_21033,N_16911,N_16207);
nor U21034 (N_21034,N_19176,N_18619);
nor U21035 (N_21035,N_15625,N_19937);
xor U21036 (N_21036,N_17644,N_18533);
xnor U21037 (N_21037,N_16839,N_17914);
nand U21038 (N_21038,N_18865,N_18651);
or U21039 (N_21039,N_18883,N_17954);
nor U21040 (N_21040,N_17623,N_17224);
or U21041 (N_21041,N_17033,N_18339);
nor U21042 (N_21042,N_15464,N_18360);
or U21043 (N_21043,N_18983,N_18390);
and U21044 (N_21044,N_18408,N_15394);
or U21045 (N_21045,N_18699,N_17882);
and U21046 (N_21046,N_15993,N_16748);
nor U21047 (N_21047,N_15807,N_15423);
nand U21048 (N_21048,N_17188,N_16294);
or U21049 (N_21049,N_18060,N_15453);
nand U21050 (N_21050,N_19512,N_17338);
nor U21051 (N_21051,N_16468,N_15434);
or U21052 (N_21052,N_17885,N_19533);
and U21053 (N_21053,N_15498,N_18689);
nor U21054 (N_21054,N_15711,N_17298);
nor U21055 (N_21055,N_15378,N_16351);
nand U21056 (N_21056,N_16740,N_18288);
xnor U21057 (N_21057,N_19044,N_19060);
and U21058 (N_21058,N_15152,N_19253);
or U21059 (N_21059,N_17833,N_15626);
nand U21060 (N_21060,N_16038,N_16559);
or U21061 (N_21061,N_19063,N_17377);
and U21062 (N_21062,N_19411,N_17531);
nand U21063 (N_21063,N_17089,N_15620);
or U21064 (N_21064,N_15632,N_16698);
and U21065 (N_21065,N_18158,N_17086);
nor U21066 (N_21066,N_17735,N_16317);
and U21067 (N_21067,N_19758,N_18410);
nor U21068 (N_21068,N_15896,N_17076);
nor U21069 (N_21069,N_16788,N_17560);
nand U21070 (N_21070,N_16145,N_16352);
nand U21071 (N_21071,N_18663,N_18637);
or U21072 (N_21072,N_17147,N_16608);
and U21073 (N_21073,N_15490,N_16601);
nor U21074 (N_21074,N_15597,N_17883);
and U21075 (N_21075,N_16968,N_17675);
or U21076 (N_21076,N_16727,N_15810);
or U21077 (N_21077,N_18639,N_16575);
xor U21078 (N_21078,N_16012,N_16508);
and U21079 (N_21079,N_19756,N_15466);
or U21080 (N_21080,N_17065,N_16986);
nand U21081 (N_21081,N_18930,N_17533);
nor U21082 (N_21082,N_15858,N_17452);
xor U21083 (N_21083,N_15100,N_18576);
nand U21084 (N_21084,N_19546,N_17342);
nor U21085 (N_21085,N_18007,N_18536);
and U21086 (N_21086,N_17419,N_19526);
nor U21087 (N_21087,N_17958,N_19831);
nor U21088 (N_21088,N_15084,N_18421);
and U21089 (N_21089,N_18645,N_16069);
and U21090 (N_21090,N_16545,N_18242);
xnor U21091 (N_21091,N_16146,N_19911);
nand U21092 (N_21092,N_16128,N_15339);
or U21093 (N_21093,N_17097,N_17259);
nor U21094 (N_21094,N_18164,N_16656);
nand U21095 (N_21095,N_16614,N_18260);
or U21096 (N_21096,N_19088,N_19156);
and U21097 (N_21097,N_17169,N_18480);
nor U21098 (N_21098,N_16652,N_17302);
and U21099 (N_21099,N_17256,N_18493);
xor U21100 (N_21100,N_18361,N_15139);
xor U21101 (N_21101,N_15776,N_17925);
nand U21102 (N_21102,N_15477,N_18245);
or U21103 (N_21103,N_15760,N_17425);
and U21104 (N_21104,N_18231,N_18277);
nor U21105 (N_21105,N_16914,N_17241);
nand U21106 (N_21106,N_17018,N_15962);
nor U21107 (N_21107,N_19479,N_15884);
nand U21108 (N_21108,N_18626,N_17835);
and U21109 (N_21109,N_19518,N_19569);
or U21110 (N_21110,N_19780,N_16987);
nor U21111 (N_21111,N_17976,N_15382);
xnor U21112 (N_21112,N_16975,N_17481);
nand U21113 (N_21113,N_16851,N_19119);
or U21114 (N_21114,N_19507,N_17962);
and U21115 (N_21115,N_16527,N_18224);
nor U21116 (N_21116,N_17471,N_15078);
xor U21117 (N_21117,N_17285,N_17502);
and U21118 (N_21118,N_19288,N_16889);
nor U21119 (N_21119,N_18758,N_19842);
nand U21120 (N_21120,N_17680,N_18160);
nor U21121 (N_21121,N_17857,N_17091);
nor U21122 (N_21122,N_15305,N_17381);
nand U21123 (N_21123,N_18553,N_18240);
and U21124 (N_21124,N_17758,N_17607);
xor U21125 (N_21125,N_15259,N_17375);
nor U21126 (N_21126,N_15813,N_17772);
nor U21127 (N_21127,N_18119,N_19103);
or U21128 (N_21128,N_19638,N_16338);
nand U21129 (N_21129,N_18351,N_17102);
or U21130 (N_21130,N_16500,N_19790);
and U21131 (N_21131,N_19621,N_19728);
nand U21132 (N_21132,N_18902,N_15909);
and U21133 (N_21133,N_18077,N_18512);
or U21134 (N_21134,N_18115,N_18794);
or U21135 (N_21135,N_15650,N_16108);
nor U21136 (N_21136,N_18317,N_18117);
or U21137 (N_21137,N_17346,N_17380);
nand U21138 (N_21138,N_18239,N_15145);
xnor U21139 (N_21139,N_16957,N_19025);
or U21140 (N_21140,N_16189,N_17685);
or U21141 (N_21141,N_16060,N_16240);
and U21142 (N_21142,N_17665,N_19154);
nand U21143 (N_21143,N_15744,N_19828);
or U21144 (N_21144,N_15454,N_19748);
xnor U21145 (N_21145,N_16389,N_17177);
and U21146 (N_21146,N_18694,N_19482);
xor U21147 (N_21147,N_16782,N_18142);
nand U21148 (N_21148,N_15839,N_16442);
and U21149 (N_21149,N_19152,N_17705);
xor U21150 (N_21150,N_17167,N_17822);
and U21151 (N_21151,N_17770,N_15131);
nand U21152 (N_21152,N_15527,N_18022);
and U21153 (N_21153,N_17368,N_19037);
nor U21154 (N_21154,N_17133,N_15895);
and U21155 (N_21155,N_18515,N_15025);
nand U21156 (N_21156,N_19072,N_19228);
or U21157 (N_21157,N_15276,N_19977);
and U21158 (N_21158,N_16700,N_19658);
nor U21159 (N_21159,N_15272,N_15688);
and U21160 (N_21160,N_17796,N_17024);
and U21161 (N_21161,N_16064,N_19753);
nor U21162 (N_21162,N_18757,N_18067);
nor U21163 (N_21163,N_19216,N_18130);
and U21164 (N_21164,N_15262,N_15999);
xor U21165 (N_21165,N_18818,N_18920);
nand U21166 (N_21166,N_15574,N_16703);
nor U21167 (N_21167,N_18387,N_17247);
nand U21168 (N_21168,N_18046,N_19062);
nand U21169 (N_21169,N_18458,N_17824);
and U21170 (N_21170,N_19130,N_16070);
nor U21171 (N_21171,N_18703,N_18618);
xnor U21172 (N_21172,N_16549,N_18460);
and U21173 (N_21173,N_16100,N_15500);
nor U21174 (N_21174,N_17283,N_16362);
and U21175 (N_21175,N_17594,N_16253);
or U21176 (N_21176,N_19229,N_15694);
or U21177 (N_21177,N_19281,N_18432);
nor U21178 (N_21178,N_15439,N_16566);
nor U21179 (N_21179,N_15127,N_15488);
and U21180 (N_21180,N_17333,N_15357);
nand U21181 (N_21181,N_15829,N_17410);
nor U21182 (N_21182,N_16400,N_18717);
and U21183 (N_21183,N_16422,N_19308);
and U21184 (N_21184,N_17155,N_16469);
nand U21185 (N_21185,N_16427,N_15073);
or U21186 (N_21186,N_16418,N_16353);
nor U21187 (N_21187,N_18507,N_15017);
or U21188 (N_21188,N_18714,N_19816);
nor U21189 (N_21189,N_18105,N_15785);
or U21190 (N_21190,N_19368,N_17207);
xnor U21191 (N_21191,N_15529,N_19679);
nor U21192 (N_21192,N_17517,N_15346);
nor U21193 (N_21193,N_16734,N_16619);
or U21194 (N_21194,N_16119,N_17880);
and U21195 (N_21195,N_15799,N_19698);
nand U21196 (N_21196,N_16988,N_15285);
nand U21197 (N_21197,N_19989,N_19183);
and U21198 (N_21198,N_19498,N_19666);
and U21199 (N_21199,N_18331,N_18568);
nor U21200 (N_21200,N_19492,N_18034);
or U21201 (N_21201,N_15470,N_18456);
or U21202 (N_21202,N_16856,N_17837);
nor U21203 (N_21203,N_15609,N_19354);
nand U21204 (N_21204,N_17524,N_17858);
or U21205 (N_21205,N_17440,N_18580);
and U21206 (N_21206,N_16796,N_16315);
or U21207 (N_21207,N_18449,N_19138);
nand U21208 (N_21208,N_16581,N_17414);
nor U21209 (N_21209,N_19171,N_19968);
and U21210 (N_21210,N_16712,N_15675);
nand U21211 (N_21211,N_17255,N_16863);
xor U21212 (N_21212,N_19594,N_16979);
xor U21213 (N_21213,N_18103,N_15480);
nand U21214 (N_21214,N_18679,N_18303);
and U21215 (N_21215,N_17286,N_16682);
or U21216 (N_21216,N_19959,N_16725);
and U21217 (N_21217,N_15358,N_16573);
xor U21218 (N_21218,N_15674,N_17565);
xor U21219 (N_21219,N_19560,N_17369);
and U21220 (N_21220,N_15655,N_15591);
and U21221 (N_21221,N_19582,N_16742);
and U21222 (N_21222,N_17749,N_18965);
or U21223 (N_21223,N_18529,N_18178);
or U21224 (N_21224,N_16870,N_19934);
or U21225 (N_21225,N_15041,N_18603);
or U21226 (N_21226,N_16661,N_18915);
and U21227 (N_21227,N_15964,N_17918);
nor U21228 (N_21228,N_16826,N_16023);
xnor U21229 (N_21229,N_16475,N_18419);
and U21230 (N_21230,N_15331,N_15054);
nand U21231 (N_21231,N_18151,N_18195);
nor U21232 (N_21232,N_19173,N_19745);
and U21233 (N_21233,N_18113,N_17998);
or U21234 (N_21234,N_17912,N_16082);
nand U21235 (N_21235,N_15687,N_15380);
nand U21236 (N_21236,N_16354,N_18244);
or U21237 (N_21237,N_15543,N_16599);
nor U21238 (N_21238,N_19040,N_16704);
and U21239 (N_21239,N_15363,N_18170);
nand U21240 (N_21240,N_18907,N_16928);
nor U21241 (N_21241,N_18054,N_19951);
or U21242 (N_21242,N_15083,N_18243);
or U21243 (N_21243,N_19854,N_17074);
or U21244 (N_21244,N_15649,N_15495);
or U21245 (N_21245,N_18066,N_18042);
or U21246 (N_21246,N_18476,N_19955);
or U21247 (N_21247,N_19917,N_16261);
nor U21248 (N_21248,N_17125,N_15211);
and U21249 (N_21249,N_16052,N_16168);
nor U21250 (N_21250,N_18944,N_16164);
and U21251 (N_21251,N_16383,N_16577);
nor U21252 (N_21252,N_19384,N_15916);
nand U21253 (N_21253,N_17439,N_16153);
or U21254 (N_21254,N_18657,N_19190);
and U21255 (N_21255,N_15643,N_15936);
nor U21256 (N_21256,N_17707,N_17519);
nor U21257 (N_21257,N_18225,N_16666);
nand U21258 (N_21258,N_15437,N_15389);
or U21259 (N_21259,N_19298,N_17876);
nor U21260 (N_21260,N_17467,N_17025);
nand U21261 (N_21261,N_18201,N_17128);
xor U21262 (N_21262,N_19712,N_17739);
nand U21263 (N_21263,N_17700,N_19402);
and U21264 (N_21264,N_16479,N_19874);
nor U21265 (N_21265,N_15436,N_16160);
and U21266 (N_21266,N_18816,N_18281);
nand U21267 (N_21267,N_19623,N_19975);
nor U21268 (N_21268,N_16985,N_18099);
and U21269 (N_21269,N_19085,N_17946);
or U21270 (N_21270,N_18903,N_18168);
nand U21271 (N_21271,N_18799,N_17935);
or U21272 (N_21272,N_19413,N_18379);
nand U21273 (N_21273,N_18116,N_15387);
and U21274 (N_21274,N_19556,N_16120);
or U21275 (N_21275,N_19725,N_16058);
nor U21276 (N_21276,N_17438,N_17111);
and U21277 (N_21277,N_19278,N_16416);
nand U21278 (N_21278,N_15472,N_19214);
or U21279 (N_21279,N_16391,N_18091);
nor U21280 (N_21280,N_16166,N_19435);
or U21281 (N_21281,N_17151,N_15487);
xnor U21282 (N_21282,N_16155,N_15683);
or U21283 (N_21283,N_18435,N_16538);
nand U21284 (N_21284,N_15309,N_17006);
xor U21285 (N_21285,N_16206,N_17558);
nand U21286 (N_21286,N_17860,N_15497);
xnor U21287 (N_21287,N_15360,N_15063);
or U21288 (N_21288,N_17181,N_16129);
xor U21289 (N_21289,N_15366,N_17974);
and U21290 (N_21290,N_17945,N_18916);
nor U21291 (N_21291,N_17924,N_17776);
nor U21292 (N_21292,N_18318,N_16365);
or U21293 (N_21293,N_17295,N_16063);
nor U21294 (N_21294,N_16246,N_17363);
nor U21295 (N_21295,N_17738,N_19047);
or U21296 (N_21296,N_19434,N_18585);
nand U21297 (N_21297,N_16326,N_19800);
and U21298 (N_21298,N_15756,N_18765);
and U21299 (N_21299,N_19182,N_19285);
nand U21300 (N_21300,N_19506,N_19274);
or U21301 (N_21301,N_17117,N_18879);
and U21302 (N_21302,N_19803,N_18933);
xnor U21303 (N_21303,N_15155,N_17761);
nand U21304 (N_21304,N_18778,N_18488);
nand U21305 (N_21305,N_17246,N_18445);
nand U21306 (N_21306,N_19960,N_19155);
nor U21307 (N_21307,N_16642,N_18844);
nand U21308 (N_21308,N_16126,N_17775);
xor U21309 (N_21309,N_15032,N_17585);
and U21310 (N_21310,N_17584,N_15621);
nor U21311 (N_21311,N_18806,N_18784);
nor U21312 (N_21312,N_15603,N_16255);
and U21313 (N_21313,N_18594,N_17045);
nand U21314 (N_21314,N_15021,N_16356);
nor U21315 (N_21315,N_19603,N_19829);
or U21316 (N_21316,N_19485,N_17821);
or U21317 (N_21317,N_17038,N_19239);
nand U21318 (N_21318,N_18519,N_15835);
or U21319 (N_21319,N_19207,N_15914);
nand U21320 (N_21320,N_19451,N_15255);
xnor U21321 (N_21321,N_15112,N_18234);
nor U21322 (N_21322,N_17293,N_15343);
nor U21323 (N_21323,N_17652,N_15546);
nand U21324 (N_21324,N_16482,N_15520);
or U21325 (N_21325,N_19465,N_15468);
xnor U21326 (N_21326,N_17083,N_18670);
nor U21327 (N_21327,N_17391,N_18466);
xor U21328 (N_21328,N_19730,N_18925);
and U21329 (N_21329,N_16229,N_18423);
nand U21330 (N_21330,N_17251,N_17514);
and U21331 (N_21331,N_15740,N_18781);
and U21332 (N_21332,N_17463,N_19952);
and U21333 (N_21333,N_18598,N_15889);
xor U21334 (N_21334,N_15671,N_19139);
or U21335 (N_21335,N_19517,N_17889);
xnor U21336 (N_21336,N_18177,N_17378);
nor U21337 (N_21337,N_16026,N_17683);
or U21338 (N_21338,N_15772,N_16795);
nand U21339 (N_21339,N_15616,N_15474);
and U21340 (N_21340,N_16923,N_15572);
nor U21341 (N_21341,N_17721,N_19304);
and U21342 (N_21342,N_19054,N_16954);
nand U21343 (N_21343,N_16384,N_18299);
or U21344 (N_21344,N_15395,N_19713);
nor U21345 (N_21345,N_15637,N_18264);
and U21346 (N_21346,N_17218,N_17988);
nor U21347 (N_21347,N_19706,N_15064);
nand U21348 (N_21348,N_19394,N_19879);
xor U21349 (N_21349,N_19083,N_16721);
or U21350 (N_21350,N_18263,N_16008);
and U21351 (N_21351,N_18986,N_15504);
or U21352 (N_21352,N_16289,N_15302);
nand U21353 (N_21353,N_18829,N_19949);
nor U21354 (N_21354,N_16436,N_15702);
and U21355 (N_21355,N_18126,N_19886);
and U21356 (N_21356,N_15101,N_16917);
nand U21357 (N_21357,N_15006,N_17612);
or U21358 (N_21358,N_16629,N_19079);
nor U21359 (N_21359,N_18579,N_19431);
nor U21360 (N_21360,N_19938,N_18497);
and U21361 (N_21361,N_18996,N_18551);
and U21362 (N_21362,N_18180,N_18482);
and U21363 (N_21363,N_19013,N_16223);
and U21364 (N_21364,N_19471,N_15011);
or U21365 (N_21365,N_17347,N_18290);
nor U21366 (N_21366,N_16665,N_15329);
or U21367 (N_21367,N_17670,N_15867);
or U21368 (N_21368,N_19896,N_15379);
and U21369 (N_21369,N_18908,N_17566);
nor U21370 (N_21370,N_18223,N_17979);
nor U21371 (N_21371,N_17639,N_18161);
nor U21372 (N_21372,N_15508,N_16935);
and U21373 (N_21373,N_16809,N_15047);
or U21374 (N_21374,N_19562,N_16814);
and U21375 (N_21375,N_16982,N_16724);
xnor U21376 (N_21376,N_19779,N_17790);
nand U21377 (N_21377,N_18960,N_16553);
nand U21378 (N_21378,N_16990,N_18487);
xnor U21379 (N_21379,N_19168,N_17573);
xor U21380 (N_21380,N_16481,N_16852);
nor U21381 (N_21381,N_15833,N_19653);
and U21382 (N_21382,N_19164,N_19537);
nand U21383 (N_21383,N_17447,N_18481);
nand U21384 (N_21384,N_19622,N_15510);
or U21385 (N_21385,N_15307,N_15698);
nor U21386 (N_21386,N_16854,N_19718);
nand U21387 (N_21387,N_15120,N_17698);
and U21388 (N_21388,N_19092,N_17418);
nand U21389 (N_21389,N_17957,N_15374);
nor U21390 (N_21390,N_19395,N_19425);
nor U21391 (N_21391,N_17759,N_16605);
nor U21392 (N_21392,N_18649,N_19220);
nand U21393 (N_21393,N_18616,N_17474);
or U21394 (N_21394,N_19016,N_19617);
xnor U21395 (N_21395,N_16754,N_19457);
xnor U21396 (N_21396,N_18929,N_19039);
or U21397 (N_21397,N_19654,N_15400);
nor U21398 (N_21398,N_18552,N_16358);
or U21399 (N_21399,N_17405,N_19264);
xor U21400 (N_21400,N_18588,N_16018);
and U21401 (N_21401,N_18864,N_16513);
and U21402 (N_21402,N_17144,N_15241);
nand U21403 (N_21403,N_15137,N_19226);
nor U21404 (N_21404,N_17106,N_15661);
and U21405 (N_21405,N_17678,N_19856);
nand U21406 (N_21406,N_19477,N_18029);
nand U21407 (N_21407,N_16595,N_17807);
nand U21408 (N_21408,N_16537,N_18189);
or U21409 (N_21409,N_19473,N_17189);
xnor U21410 (N_21410,N_16420,N_16313);
xor U21411 (N_21411,N_15714,N_16350);
nand U21412 (N_21412,N_15837,N_17364);
or U21413 (N_21413,N_18857,N_18675);
xnor U21414 (N_21414,N_18332,N_18229);
and U21415 (N_21415,N_17856,N_15310);
nand U21416 (N_21416,N_15115,N_18846);
and U21417 (N_21417,N_18561,N_18340);
and U21418 (N_21418,N_18992,N_15822);
or U21419 (N_21419,N_18632,N_16641);
nor U21420 (N_21420,N_19665,N_18989);
and U21421 (N_21421,N_15492,N_19287);
nor U21422 (N_21422,N_17379,N_19241);
or U21423 (N_21423,N_16503,N_16702);
nand U21424 (N_21424,N_19962,N_18269);
or U21425 (N_21425,N_19864,N_17153);
or U21426 (N_21426,N_18502,N_18398);
nor U21427 (N_21427,N_16388,N_18457);
or U21428 (N_21428,N_16113,N_17518);
and U21429 (N_21429,N_18082,N_15762);
nand U21430 (N_21430,N_16799,N_18805);
nor U21431 (N_21431,N_16644,N_19436);
or U21432 (N_21432,N_15432,N_19946);
nand U21433 (N_21433,N_18073,N_15288);
and U21434 (N_21434,N_15425,N_19619);
nand U21435 (N_21435,N_15944,N_18267);
or U21436 (N_21436,N_17555,N_18595);
xor U21437 (N_21437,N_16636,N_16836);
or U21438 (N_21438,N_17795,N_17984);
and U21439 (N_21439,N_18541,N_15705);
nor U21440 (N_21440,N_17630,N_16920);
or U21441 (N_21441,N_18344,N_15552);
xnor U21442 (N_21442,N_15778,N_16669);
and U21443 (N_21443,N_15016,N_16736);
or U21444 (N_21444,N_15857,N_17236);
or U21445 (N_21445,N_19853,N_15494);
or U21446 (N_21446,N_18352,N_15230);
or U21447 (N_21447,N_18548,N_16088);
and U21448 (N_21448,N_19847,N_16522);
and U21449 (N_21449,N_17947,N_19020);
and U21450 (N_21450,N_18601,N_18058);
or U21451 (N_21451,N_17215,N_19462);
and U21452 (N_21452,N_16849,N_16028);
and U21453 (N_21453,N_16778,N_15140);
nand U21454 (N_21454,N_19768,N_18355);
and U21455 (N_21455,N_16658,N_19120);
and U21456 (N_21456,N_17021,N_16234);
or U21457 (N_21457,N_15265,N_15093);
or U21458 (N_21458,N_16159,N_15370);
or U21459 (N_21459,N_18167,N_15247);
and U21460 (N_21460,N_16866,N_16148);
or U21461 (N_21461,N_17896,N_18342);
and U21462 (N_21462,N_19041,N_18593);
nand U21463 (N_21463,N_18531,N_19585);
nand U21464 (N_21464,N_15475,N_17108);
nand U21465 (N_21465,N_15577,N_19481);
and U21466 (N_21466,N_17388,N_19535);
or U21467 (N_21467,N_19038,N_19979);
nor U21468 (N_21468,N_16429,N_17084);
xor U21469 (N_21469,N_17938,N_19687);
or U21470 (N_21470,N_19503,N_18659);
nor U21471 (N_21471,N_17424,N_17127);
and U21472 (N_21472,N_19525,N_16144);
and U21473 (N_21473,N_19776,N_19969);
nor U21474 (N_21474,N_16449,N_15385);
and U21475 (N_21475,N_17510,N_18658);
xnor U21476 (N_21476,N_15420,N_19172);
nor U21477 (N_21477,N_15209,N_18684);
or U21478 (N_21478,N_17406,N_15938);
or U21479 (N_21479,N_18773,N_15053);
or U21480 (N_21480,N_17637,N_18499);
nor U21481 (N_21481,N_19475,N_18026);
or U21482 (N_21482,N_19703,N_15388);
nor U21483 (N_21483,N_16053,N_19467);
and U21484 (N_21484,N_19994,N_18295);
nand U21485 (N_21485,N_15371,N_19559);
nand U21486 (N_21486,N_19259,N_17278);
and U21487 (N_21487,N_19162,N_19375);
nor U21488 (N_21488,N_17862,N_19221);
and U21489 (N_21489,N_16562,N_17290);
or U21490 (N_21490,N_17673,N_19339);
nand U21491 (N_21491,N_19561,N_19032);
and U21492 (N_21492,N_15586,N_17116);
nand U21493 (N_21493,N_15424,N_16817);
nand U21494 (N_21494,N_18241,N_16370);
nand U21495 (N_21495,N_18320,N_17197);
or U21496 (N_21496,N_19834,N_17967);
and U21497 (N_21497,N_18249,N_16894);
nor U21498 (N_21498,N_17407,N_18721);
and U21499 (N_21499,N_19260,N_15237);
nand U21500 (N_21500,N_18690,N_17470);
and U21501 (N_21501,N_16090,N_15846);
or U21502 (N_21502,N_15026,N_16530);
or U21503 (N_21503,N_19073,N_19217);
nand U21504 (N_21504,N_17282,N_17520);
nand U21505 (N_21505,N_19649,N_17595);
nand U21506 (N_21506,N_15843,N_19942);
or U21507 (N_21507,N_15585,N_18446);
or U21508 (N_21508,N_19293,N_18090);
nand U21509 (N_21509,N_16221,N_15383);
nand U21510 (N_21510,N_15673,N_19064);
nand U21511 (N_21511,N_16816,N_17592);
nand U21512 (N_21512,N_19643,N_16296);
nand U21513 (N_21513,N_17916,N_17513);
nand U21514 (N_21514,N_15704,N_15654);
or U21515 (N_21515,N_18505,N_15407);
nand U21516 (N_21516,N_18755,N_15236);
nor U21517 (N_21517,N_16910,N_19501);
nand U21518 (N_21518,N_16094,N_19090);
and U21519 (N_21519,N_15390,N_18455);
and U21520 (N_21520,N_19695,N_17200);
or U21521 (N_21521,N_15177,N_19771);
and U21522 (N_21522,N_15517,N_19012);
xnor U21523 (N_21523,N_18268,N_18710);
and U21524 (N_21524,N_18976,N_19589);
or U21525 (N_21525,N_15736,N_18298);
and U21526 (N_21526,N_16021,N_19391);
nor U21527 (N_21527,N_15522,N_16933);
and U21528 (N_21528,N_17643,N_15160);
and U21529 (N_21529,N_15151,N_18019);
or U21530 (N_21530,N_17867,N_17541);
nor U21531 (N_21531,N_16878,N_15881);
nor U21532 (N_21532,N_15174,N_16501);
nor U21533 (N_21533,N_17146,N_16335);
nand U21534 (N_21534,N_15757,N_16162);
nor U21535 (N_21535,N_19291,N_15859);
nor U21536 (N_21536,N_15805,N_16424);
nor U21537 (N_21537,N_19987,N_16798);
or U21538 (N_21538,N_17873,N_16708);
or U21539 (N_21539,N_17869,N_16555);
and U21540 (N_21540,N_15351,N_16857);
or U21541 (N_21541,N_17851,N_17132);
and U21542 (N_21542,N_15295,N_15602);
and U21543 (N_21543,N_16464,N_16797);
or U21544 (N_21544,N_19245,N_17192);
nor U21545 (N_21545,N_17008,N_18539);
or U21546 (N_21546,N_18681,N_17001);
or U21547 (N_21547,N_18564,N_15037);
xor U21548 (N_21548,N_17809,N_18954);
or U21549 (N_21549,N_19772,N_17112);
nand U21550 (N_21550,N_19455,N_15409);
and U21551 (N_21551,N_18769,N_18692);
nand U21552 (N_21552,N_18739,N_16216);
nand U21553 (N_21553,N_15699,N_17456);
or U21554 (N_21554,N_19819,N_17477);
or U21555 (N_21555,N_17042,N_17260);
and U21556 (N_21556,N_17176,N_17619);
xor U21557 (N_21557,N_19433,N_19348);
and U21558 (N_21558,N_18012,N_15087);
nor U21559 (N_21559,N_18667,N_18433);
and U21560 (N_21560,N_17137,N_18974);
and U21561 (N_21561,N_17521,N_17636);
and U21562 (N_21562,N_16624,N_18490);
or U21563 (N_21563,N_16186,N_19868);
nand U21564 (N_21564,N_19458,N_18020);
or U21565 (N_21565,N_15181,N_19420);
nor U21566 (N_21566,N_17401,N_17571);
or U21567 (N_21567,N_15506,N_15726);
nand U21568 (N_21568,N_16783,N_19312);
xor U21569 (N_21569,N_15645,N_19272);
or U21570 (N_21570,N_18056,N_16397);
nor U21571 (N_21571,N_17506,N_17540);
nand U21572 (N_21572,N_19224,N_19252);
or U21573 (N_21573,N_15554,N_18957);
nor U21574 (N_21574,N_17496,N_17331);
nand U21575 (N_21575,N_17071,N_19135);
nor U21576 (N_21576,N_19633,N_17318);
nand U21577 (N_21577,N_15670,N_15154);
nor U21578 (N_21578,N_17416,N_17581);
xor U21579 (N_21579,N_18741,N_18600);
and U21580 (N_21580,N_16561,N_19019);
nor U21581 (N_21581,N_18050,N_15435);
xnor U21582 (N_21582,N_17175,N_18856);
nand U21583 (N_21583,N_18417,N_19642);
nand U21584 (N_21584,N_19686,N_18169);
nand U21585 (N_21585,N_16871,N_16804);
nand U21586 (N_21586,N_19028,N_15831);
and U21587 (N_21587,N_16541,N_18842);
nand U21588 (N_21588,N_16640,N_17839);
nand U21589 (N_21589,N_17847,N_15443);
xnor U21590 (N_21590,N_16065,N_15421);
nor U21591 (N_21591,N_17723,N_18946);
nand U21592 (N_21592,N_15558,N_15051);
nand U21593 (N_21593,N_19324,N_15126);
nor U21594 (N_21594,N_17402,N_16521);
nand U21595 (N_21595,N_15105,N_15440);
nor U21596 (N_21596,N_19499,N_16182);
and U21597 (N_21597,N_17755,N_16176);
xor U21598 (N_21598,N_17624,N_18707);
xnor U21599 (N_21599,N_18774,N_18687);
or U21600 (N_21600,N_17658,N_19390);
and U21601 (N_21601,N_16743,N_19826);
nor U21602 (N_21602,N_16941,N_19913);
nor U21603 (N_21603,N_16263,N_19337);
or U21604 (N_21604,N_19944,N_15208);
and U21605 (N_21605,N_16408,N_19646);
or U21606 (N_21606,N_17713,N_15784);
xor U21607 (N_21607,N_17767,N_18893);
or U21608 (N_21608,N_19300,N_16655);
nor U21609 (N_21609,N_18555,N_16713);
or U21610 (N_21610,N_18011,N_15662);
nor U21611 (N_21611,N_18429,N_15028);
and U21612 (N_21612,N_16152,N_18973);
or U21613 (N_21613,N_17004,N_18439);
nor U21614 (N_21614,N_18664,N_16840);
and U21615 (N_21615,N_16623,N_15324);
nor U21616 (N_21616,N_16768,N_17561);
xnor U21617 (N_21617,N_19721,N_19379);
and U21618 (N_21618,N_18610,N_16439);
and U21619 (N_21619,N_18345,N_18048);
or U21620 (N_21620,N_17877,N_17722);
xor U21621 (N_21621,N_18611,N_15653);
xnor U21622 (N_21622,N_15723,N_19200);
or U21623 (N_21623,N_16333,N_15202);
nor U21624 (N_21624,N_18728,N_18406);
and U21625 (N_21625,N_16580,N_17734);
or U21626 (N_21626,N_16506,N_18064);
nor U21627 (N_21627,N_18033,N_19194);
nor U21628 (N_21628,N_18252,N_15184);
or U21629 (N_21629,N_17939,N_16800);
nand U21630 (N_21630,N_15377,N_19970);
and U21631 (N_21631,N_15551,N_16232);
and U21632 (N_21632,N_19108,N_16626);
xnor U21633 (N_21633,N_16916,N_18701);
and U21634 (N_21634,N_17942,N_17676);
nand U21635 (N_21635,N_19884,N_16407);
xnor U21636 (N_21636,N_16055,N_19726);
or U21637 (N_21637,N_17866,N_18140);
nand U21638 (N_21638,N_15356,N_16115);
nor U21639 (N_21639,N_16187,N_16434);
nand U21640 (N_21640,N_19683,N_17875);
and U21641 (N_21641,N_18100,N_17253);
nand U21642 (N_21642,N_19359,N_15214);
xor U21643 (N_21643,N_18120,N_18214);
or U21644 (N_21644,N_16560,N_15106);
nor U21645 (N_21645,N_18154,N_16978);
or U21646 (N_21646,N_15323,N_16044);
or U21647 (N_21647,N_16086,N_15399);
nor U21648 (N_21648,N_15334,N_16683);
xnor U21649 (N_21649,N_15971,N_16710);
and U21650 (N_21650,N_18270,N_19004);
and U21651 (N_21651,N_15741,N_16321);
or U21652 (N_21652,N_16133,N_17015);
or U21653 (N_21653,N_15567,N_15777);
or U21654 (N_21654,N_17550,N_17398);
nor U21655 (N_21655,N_18881,N_17310);
nand U21656 (N_21656,N_17648,N_17563);
or U21657 (N_21657,N_15737,N_17704);
nor U21658 (N_21658,N_16273,N_18782);
and U21659 (N_21659,N_19719,N_19509);
or U21660 (N_21660,N_19639,N_18102);
or U21661 (N_21661,N_19075,N_19870);
or U21662 (N_21662,N_17650,N_15213);
nor U21663 (N_21663,N_16066,N_16563);
xnor U21664 (N_21664,N_15912,N_16462);
nor U21665 (N_21665,N_15749,N_17427);
and U21666 (N_21666,N_15191,N_19692);
nor U21667 (N_21667,N_17934,N_15753);
nand U21668 (N_21668,N_17983,N_18300);
xor U21669 (N_21669,N_19811,N_19268);
and U21670 (N_21670,N_15109,N_17141);
nor U21671 (N_21671,N_15610,N_16276);
nor U21672 (N_21672,N_17503,N_15743);
and U21673 (N_21673,N_16080,N_16578);
and U21674 (N_21674,N_17699,N_18338);
or U21675 (N_21675,N_16828,N_15629);
or U21676 (N_21676,N_18289,N_16293);
xor U21677 (N_21677,N_17689,N_16908);
xnor U21678 (N_21678,N_16022,N_17143);
or U21679 (N_21679,N_17725,N_18836);
nor U21680 (N_21680,N_18615,N_19255);
nor U21681 (N_21681,N_18789,N_17784);
nand U21682 (N_21682,N_15975,N_18279);
nand U21683 (N_21683,N_15301,N_15198);
and U21684 (N_21684,N_15852,N_17556);
nand U21685 (N_21685,N_17609,N_15582);
nand U21686 (N_21686,N_19299,N_16256);
nor U21687 (N_21687,N_18669,N_18872);
and U21688 (N_21688,N_17003,N_17906);
and U21689 (N_21689,N_17219,N_16591);
nand U21690 (N_21690,N_15960,N_19552);
and U21691 (N_21691,N_16067,N_15096);
or U21692 (N_21692,N_19131,N_17611);
nor U21693 (N_21693,N_17034,N_18891);
and U21694 (N_21694,N_17426,N_15739);
and U21695 (N_21695,N_15665,N_17668);
nor U21696 (N_21696,N_17199,N_16714);
or U21697 (N_21697,N_17240,N_15240);
or U21698 (N_21698,N_18904,N_19389);
or U21699 (N_21699,N_18219,N_18465);
nand U21700 (N_21700,N_17703,N_19122);
or U21701 (N_21701,N_16179,N_17070);
or U21702 (N_21702,N_17296,N_18969);
and U21703 (N_21703,N_16888,N_18176);
or U21704 (N_21704,N_19483,N_18873);
or U21705 (N_21705,N_15729,N_18021);
or U21706 (N_21706,N_19280,N_19157);
and U21707 (N_21707,N_15142,N_15560);
nor U21708 (N_21708,N_15512,N_17621);
nor U21709 (N_21709,N_17397,N_19796);
nand U21710 (N_21710,N_16918,N_18590);
or U21711 (N_21711,N_17708,N_18070);
nand U21712 (N_21712,N_17041,N_17978);
and U21713 (N_21713,N_16877,N_16386);
or U21714 (N_21714,N_17905,N_15745);
and U21715 (N_21715,N_19494,N_16729);
and U21716 (N_21716,N_17441,N_16771);
nand U21717 (N_21717,N_19369,N_19732);
xnor U21718 (N_21718,N_18293,N_16654);
and U21719 (N_21719,N_18286,N_16504);
or U21720 (N_21720,N_15672,N_17157);
nand U21721 (N_21721,N_18181,N_16962);
nand U21722 (N_21722,N_19555,N_16075);
nand U21723 (N_21723,N_16328,N_16013);
nand U21724 (N_21724,N_17453,N_17499);
or U21725 (N_21725,N_17037,N_17838);
or U21726 (N_21726,N_15167,N_15403);
and U21727 (N_21727,N_19000,N_19066);
xor U21728 (N_21728,N_16803,N_15417);
and U21729 (N_21729,N_15528,N_17161);
nor U21730 (N_21730,N_19857,N_17202);
nand U21731 (N_21731,N_18319,N_16617);
and U21732 (N_21732,N_17040,N_19724);
nor U21733 (N_21733,N_18825,N_16140);
and U21734 (N_21734,N_19206,N_18931);
nand U21735 (N_21735,N_17210,N_15747);
nand U21736 (N_21736,N_18078,N_16310);
nor U21737 (N_21737,N_15094,N_17284);
and U21738 (N_21738,N_16630,N_19757);
nor U21739 (N_21739,N_19029,N_15775);
xor U21740 (N_21740,N_16946,N_18898);
xor U21741 (N_21741,N_15239,N_17926);
or U21742 (N_21742,N_17484,N_17372);
nand U21743 (N_21743,N_16257,N_18508);
nand U21744 (N_21744,N_17995,N_19273);
nand U21745 (N_21745,N_15125,N_17599);
and U21746 (N_21746,N_18337,N_15485);
or U21747 (N_21747,N_16616,N_17094);
and U21748 (N_21748,N_18323,N_19198);
nand U21749 (N_21749,N_19906,N_17105);
nor U21750 (N_21750,N_18370,N_18866);
or U21751 (N_21751,N_18217,N_19144);
or U21752 (N_21752,N_18779,N_17965);
and U21753 (N_21753,N_15887,N_15097);
nor U21754 (N_21754,N_16395,N_17498);
nor U21755 (N_21755,N_17445,N_18402);
or U21756 (N_21756,N_19635,N_15030);
nor U21757 (N_21757,N_17016,N_18474);
nor U21758 (N_21758,N_15598,N_19543);
nand U21759 (N_21759,N_18604,N_15188);
or U21760 (N_21760,N_16952,N_19204);
and U21761 (N_21761,N_16279,N_17007);
nor U21762 (N_21762,N_17437,N_16777);
or U21763 (N_21763,N_17715,N_16590);
nand U21764 (N_21764,N_15809,N_15917);
nand U21765 (N_21765,N_19213,N_19878);
nand U21766 (N_21766,N_16271,N_15143);
nand U21767 (N_21767,N_19080,N_17692);
and U21768 (N_21768,N_18327,N_17742);
nor U21769 (N_21769,N_18613,N_15928);
nor U21770 (N_21770,N_16523,N_19818);
and U21771 (N_21771,N_17572,N_18207);
or U21772 (N_21772,N_18776,N_19595);
xor U21773 (N_21773,N_18221,N_15717);
nor U21774 (N_21774,N_18828,N_17649);
and U21775 (N_21775,N_18964,N_17268);
or U21776 (N_21776,N_18988,N_16664);
nand U21777 (N_21777,N_16035,N_18798);
or U21778 (N_21778,N_15973,N_18477);
nor U21779 (N_21779,N_19105,N_18971);
or U21780 (N_21780,N_18434,N_18951);
or U21781 (N_21781,N_16633,N_18009);
nand U21782 (N_21782,N_18321,N_16319);
and U21783 (N_21783,N_16921,N_17072);
nand U21784 (N_21784,N_18310,N_17458);
xnor U21785 (N_21785,N_15579,N_16209);
or U21786 (N_21786,N_15431,N_15069);
nor U21787 (N_21787,N_15800,N_15268);
or U21788 (N_21788,N_19344,N_17589);
and U21789 (N_21789,N_18085,N_15963);
nand U21790 (N_21790,N_16057,N_16790);
nor U21791 (N_21791,N_17587,N_16993);
xnor U21792 (N_21792,N_17848,N_15830);
and U21793 (N_21793,N_18208,N_15347);
nand U21794 (N_21794,N_16891,N_19648);
nand U21795 (N_21795,N_16841,N_19376);
nor U21796 (N_21796,N_18247,N_19922);
nand U21797 (N_21797,N_17778,N_19710);
nand U21798 (N_21798,N_16403,N_18950);
and U21799 (N_21799,N_19872,N_18540);
nand U21800 (N_21800,N_19892,N_17635);
or U21801 (N_21801,N_16332,N_19544);
or U21802 (N_21802,N_16265,N_17178);
or U21803 (N_21803,N_17583,N_15362);
nand U21804 (N_21804,N_17068,N_16454);
xnor U21805 (N_21805,N_19215,N_18000);
or U21806 (N_21806,N_17222,N_17399);
and U21807 (N_21807,N_18841,N_19919);
nand U21808 (N_21808,N_15206,N_18222);
and U21809 (N_21809,N_16298,N_15664);
and U21810 (N_21810,N_19810,N_19571);
nor U21811 (N_21811,N_18259,N_15061);
and U21812 (N_21812,N_15321,N_17931);
nand U21813 (N_21813,N_18171,N_16428);
or U21814 (N_21814,N_18114,N_17020);
nand U21815 (N_21815,N_18266,N_18913);
and U21816 (N_21816,N_15327,N_18287);
nor U21817 (N_21817,N_18796,N_16224);
xnor U21818 (N_21818,N_17212,N_18695);
or U21819 (N_21819,N_15798,N_15515);
nand U21820 (N_21820,N_17136,N_15636);
and U21821 (N_21821,N_18135,N_16034);
or U21822 (N_21822,N_17371,N_18431);
or U21823 (N_21823,N_15748,N_18704);
nor U21824 (N_21824,N_19656,N_15724);
or U21825 (N_21825,N_16812,N_17299);
nand U21826 (N_21826,N_19143,N_19158);
nor U21827 (N_21827,N_16009,N_19914);
nor U21828 (N_21828,N_19967,N_17693);
nor U21829 (N_21829,N_18030,N_17800);
and U21830 (N_21830,N_15977,N_17604);
and U21831 (N_21831,N_18560,N_18411);
xor U21832 (N_21832,N_18325,N_16334);
nand U21833 (N_21833,N_16576,N_16813);
or U21834 (N_21834,N_15384,N_19452);
or U21835 (N_21835,N_18376,N_15615);
nand U21836 (N_21836,N_18640,N_16930);
nor U21837 (N_21837,N_19773,N_19026);
or U21838 (N_21838,N_19177,N_18641);
xnor U21839 (N_21839,N_15286,N_19101);
and U21840 (N_21840,N_19353,N_16807);
or U21841 (N_21841,N_19426,N_15086);
nor U21842 (N_21842,N_18814,N_19071);
nand U21843 (N_21843,N_16083,N_16845);
and U21844 (N_21844,N_16558,N_16838);
or U21845 (N_21845,N_16625,N_18226);
nand U21846 (N_21846,N_16602,N_17941);
nand U21847 (N_21847,N_19644,N_15192);
nor U21848 (N_21848,N_19852,N_16529);
or U21849 (N_21849,N_17537,N_19409);
xnor U21850 (N_21850,N_19193,N_15144);
xor U21851 (N_21851,N_18683,N_19010);
nor U21852 (N_21852,N_15732,N_16374);
and U21853 (N_21853,N_17544,N_16893);
nor U21854 (N_21854,N_16547,N_15196);
xor U21855 (N_21855,N_16498,N_15499);
nor U21856 (N_21856,N_16762,N_19788);
and U21857 (N_21857,N_17118,N_15604);
or U21858 (N_21858,N_15634,N_15187);
and U21859 (N_21859,N_16340,N_15274);
nand U21860 (N_21860,N_18634,N_16047);
and U21861 (N_21861,N_19586,N_17696);
nand U21862 (N_21862,N_15349,N_16526);
nor U21863 (N_21863,N_16461,N_15947);
and U21864 (N_21864,N_19542,N_19124);
or U21865 (N_21865,N_17090,N_16175);
nor U21866 (N_21866,N_15856,N_16706);
nor U21867 (N_21867,N_16107,N_18677);
or U21868 (N_21868,N_18475,N_16157);
and U21869 (N_21869,N_15242,N_16493);
or U21870 (N_21870,N_15082,N_19614);
nor U21871 (N_21871,N_17578,N_15861);
nor U21872 (N_21872,N_18845,N_15595);
or U21873 (N_21873,N_19807,N_19738);
or U21874 (N_21874,N_16171,N_19109);
nand U21875 (N_21875,N_17273,N_19677);
xor U21876 (N_21876,N_18211,N_15863);
nor U21877 (N_21877,N_19939,N_19727);
nand U21878 (N_21878,N_18506,N_17332);
nand U21879 (N_21879,N_15253,N_15195);
nand U21880 (N_21880,N_16440,N_15639);
xnor U21881 (N_21881,N_17457,N_16327);
and U21882 (N_21882,N_16045,N_18972);
or U21883 (N_21883,N_17140,N_19140);
xor U21884 (N_21884,N_17726,N_15102);
nor U21885 (N_21885,N_18578,N_15303);
and U21886 (N_21886,N_18316,N_17733);
or U21887 (N_21887,N_16027,N_15340);
and U21888 (N_21888,N_16515,N_16996);
nor U21889 (N_21889,N_19541,N_15712);
nor U21890 (N_21890,N_16062,N_17490);
nor U21891 (N_21891,N_16584,N_18572);
or U21892 (N_21892,N_19128,N_18373);
nor U21893 (N_21893,N_19923,N_15226);
nand U21894 (N_21894,N_17750,N_17325);
or U21895 (N_21895,N_15252,N_18935);
or U21896 (N_21896,N_19372,N_17666);
and U21897 (N_21897,N_16847,N_15050);
nor U21898 (N_21898,N_15931,N_19077);
and U21899 (N_21899,N_19545,N_15584);
nand U21900 (N_21900,N_16017,N_15945);
and U21901 (N_21901,N_17367,N_16915);
nand U21902 (N_21902,N_18843,N_19694);
and U21903 (N_21903,N_15367,N_16037);
nor U21904 (N_21904,N_15081,N_18375);
or U21905 (N_21905,N_19036,N_17196);
and U21906 (N_21906,N_19824,N_19598);
and U21907 (N_21907,N_16141,N_17899);
and U21908 (N_21908,N_19849,N_15578);
and U21909 (N_21909,N_17973,N_16785);
nor U21910 (N_21910,N_17971,N_19270);
nor U21911 (N_21911,N_16763,N_16399);
nor U21912 (N_21912,N_15178,N_15933);
nand U21913 (N_21913,N_16540,N_16131);
nor U21914 (N_21914,N_15926,N_17570);
nand U21915 (N_21915,N_15071,N_19672);
or U21916 (N_21916,N_18122,N_17500);
nand U21917 (N_21917,N_19222,N_19777);
xor U21918 (N_21918,N_19068,N_18322);
and U21919 (N_21919,N_19367,N_17717);
and U21920 (N_21920,N_16165,N_17171);
or U21921 (N_21921,N_18979,N_18780);
and U21922 (N_21922,N_18952,N_17183);
and U21923 (N_21923,N_19195,N_19315);
nand U21924 (N_21924,N_18291,N_19988);
nand U21925 (N_21925,N_16862,N_19612);
or U21926 (N_21926,N_19637,N_16109);
nor U21927 (N_21927,N_19640,N_15018);
and U21928 (N_21928,N_16718,N_19832);
or U21929 (N_21929,N_16668,N_17444);
nor U21930 (N_21930,N_16645,N_17227);
nand U21931 (N_21931,N_15336,N_16193);
nand U21932 (N_21932,N_16588,N_19414);
or U21933 (N_21933,N_16789,N_15774);
nor U21934 (N_21934,N_18827,N_17257);
and U21935 (N_21935,N_15138,N_18725);
nor U21936 (N_21936,N_18597,N_19493);
nor U21937 (N_21937,N_16773,N_17554);
or U21938 (N_21938,N_19996,N_17843);
nor U21939 (N_21939,N_15085,N_15845);
xor U21940 (N_21940,N_19430,N_16377);
or U21941 (N_21941,N_18622,N_15998);
or U21942 (N_21942,N_16443,N_19995);
nand U21943 (N_21943,N_19863,N_16951);
nand U21944 (N_21944,N_18285,N_18282);
and U21945 (N_21945,N_18188,N_16524);
nor U21946 (N_21946,N_17092,N_19574);
nand U21947 (N_21947,N_15254,N_18218);
nand U21948 (N_21948,N_19381,N_18394);
and U21949 (N_21949,N_15935,N_16305);
and U21950 (N_21950,N_18409,N_17633);
nand U21951 (N_21951,N_18069,N_19106);
or U21952 (N_21952,N_15141,N_17686);
xor U21953 (N_21953,N_19148,N_18049);
nor U21954 (N_21954,N_17820,N_18712);
and U21955 (N_21955,N_15669,N_19427);
and U21956 (N_21956,N_16805,N_15752);
nor U21957 (N_21957,N_18001,N_19400);
or U21958 (N_21958,N_16314,N_17002);
nor U21959 (N_21959,N_15874,N_18719);
or U21960 (N_21960,N_18987,N_16574);
and U21961 (N_21961,N_18643,N_17488);
nor U21962 (N_21962,N_15271,N_18257);
nand U21963 (N_21963,N_16579,N_19741);
nand U21964 (N_21964,N_15547,N_17214);
and U21965 (N_21965,N_17657,N_15607);
and U21966 (N_21966,N_15855,N_17616);
and U21967 (N_21967,N_16238,N_19468);
or U21968 (N_21968,N_18051,N_16548);
or U21969 (N_21969,N_17029,N_16277);
and U21970 (N_21970,N_16178,N_19785);
nor U21971 (N_21971,N_19593,N_17968);
nor U21972 (N_21972,N_18955,N_17327);
nor U21973 (N_21973,N_15969,N_18821);
and U21974 (N_21974,N_17064,N_15892);
and U21975 (N_21975,N_17605,N_18822);
nor U21976 (N_21976,N_19018,N_19775);
or U21977 (N_21977,N_17052,N_19580);
and U21978 (N_21978,N_18718,N_18697);
or U21979 (N_21979,N_18924,N_15227);
and U21980 (N_21980,N_19491,N_17972);
nor U21981 (N_21981,N_18389,N_15957);
nand U21982 (N_21982,N_17751,N_19089);
or U21983 (N_21983,N_17231,N_16583);
and U21984 (N_21984,N_16025,N_19472);
and U21985 (N_21985,N_19707,N_19933);
and U21986 (N_21986,N_17991,N_18448);
or U21987 (N_21987,N_18525,N_15996);
nand U21988 (N_21988,N_15871,N_15001);
xor U21989 (N_21989,N_19159,N_19234);
or U21990 (N_21990,N_17655,N_18628);
nand U21991 (N_21991,N_15284,N_17949);
and U21992 (N_21992,N_19488,N_19231);
and U21993 (N_21993,N_16118,N_16815);
and U21994 (N_21994,N_17486,N_16825);
or U21995 (N_21995,N_18696,N_19137);
or U21996 (N_21996,N_17653,N_18124);
nor U21997 (N_21997,N_18015,N_17245);
nor U21998 (N_21998,N_19664,N_18967);
nand U21999 (N_21999,N_16450,N_16010);
and U22000 (N_22000,N_16330,N_16309);
or U22001 (N_22001,N_18395,N_18623);
or U22002 (N_22002,N_19783,N_17773);
and U22003 (N_22003,N_15332,N_17035);
nand U22004 (N_22004,N_17763,N_19100);
nand U22005 (N_22005,N_17322,N_19310);
and U22006 (N_22006,N_17013,N_15482);
and U22007 (N_22007,N_16707,N_18324);
nor U22008 (N_22008,N_15411,N_15879);
or U22009 (N_22009,N_15994,N_16192);
or U22010 (N_22010,N_16137,N_18577);
nand U22011 (N_22011,N_16104,N_19399);
nand U22012 (N_22012,N_16117,N_15568);
and U22013 (N_22013,N_17662,N_15298);
and U22014 (N_22014,N_16267,N_18738);
nand U22015 (N_22015,N_17881,N_16663);
xnor U22016 (N_22016,N_17805,N_16040);
nor U22017 (N_22017,N_18326,N_18607);
or U22018 (N_22018,N_15386,N_18027);
and U22019 (N_22019,N_18862,N_15989);
nand U22020 (N_22020,N_18443,N_17874);
or U22021 (N_22021,N_15721,N_19170);
or U22022 (N_22022,N_16678,N_18438);
or U22023 (N_22023,N_17632,N_19822);
and U22024 (N_22024,N_16585,N_15986);
nor U22025 (N_22025,N_15997,N_15932);
nand U22026 (N_22026,N_17664,N_18858);
nand U22027 (N_22027,N_15834,N_18621);
nand U22028 (N_22028,N_18498,N_16900);
xor U22029 (N_22029,N_16344,N_16749);
nand U22030 (N_22030,N_16081,N_18462);
nor U22031 (N_22031,N_18232,N_15452);
nand U22032 (N_22032,N_18292,N_19238);
and U22033 (N_22033,N_15613,N_15766);
nand U22034 (N_22034,N_19629,N_19313);
nor U22035 (N_22035,N_15445,N_17660);
nand U22036 (N_22036,N_17182,N_19647);
or U22037 (N_22037,N_18200,N_16228);
or U22038 (N_22038,N_19125,N_16200);
xnor U22039 (N_22039,N_18982,N_16932);
or U22040 (N_22040,N_16517,N_15473);
nor U22041 (N_22041,N_19282,N_17959);
nor U22042 (N_22042,N_17443,N_18918);
nor U22043 (N_22043,N_16509,N_18248);
nor U22044 (N_22044,N_17872,N_16834);
or U22045 (N_22045,N_15165,N_16715);
nor U22046 (N_22046,N_18464,N_18254);
and U22047 (N_22047,N_18581,N_18380);
or U22048 (N_22048,N_15755,N_15121);
and U22049 (N_22049,N_16404,N_15264);
and U22050 (N_22050,N_19821,N_19781);
nor U22051 (N_22051,N_16586,N_18874);
and U22052 (N_22052,N_15257,N_19722);
and U22053 (N_22053,N_17970,N_15581);
xnor U22054 (N_22054,N_18870,N_17961);
or U22055 (N_22055,N_15876,N_17301);
nor U22056 (N_22056,N_18123,N_19008);
or U22057 (N_22057,N_18437,N_18329);
nor U22058 (N_22058,N_15885,N_19057);
xnor U22059 (N_22059,N_19311,N_18617);
or U22060 (N_22060,N_17129,N_18088);
and U22061 (N_22061,N_19843,N_17473);
nand U22062 (N_22062,N_18543,N_15057);
nand U22063 (N_22063,N_17597,N_15350);
and U22064 (N_22064,N_19615,N_15758);
and U22065 (N_22065,N_18013,N_18132);
xnor U22066 (N_22066,N_17539,N_17436);
nor U22067 (N_22067,N_19769,N_19889);
or U22068 (N_22068,N_19086,N_17472);
and U22069 (N_22069,N_16030,N_19723);
nor U22070 (N_22070,N_18559,N_17920);
or U22071 (N_22071,N_19115,N_18349);
and U22072 (N_22072,N_17101,N_17702);
nor U22073 (N_22073,N_18910,N_19059);
xnor U22074 (N_22074,N_17448,N_16372);
and U22075 (N_22075,N_18754,N_16019);
and U22076 (N_22076,N_15193,N_15691);
and U22077 (N_22077,N_17788,N_16940);
xnor U22078 (N_22078,N_17352,N_18583);
and U22079 (N_22079,N_18371,N_15535);
nand U22080 (N_22080,N_15708,N_19763);
and U22081 (N_22081,N_18890,N_18179);
nand U22082 (N_22082,N_15556,N_19548);
and U22083 (N_22083,N_18948,N_15940);
nand U22084 (N_22084,N_17019,N_17274);
nor U22085 (N_22085,N_19844,N_19334);
nor U22086 (N_22086,N_18909,N_19514);
and U22087 (N_22087,N_15287,N_18271);
nand U22088 (N_22088,N_18004,N_19524);
or U22089 (N_22089,N_16297,N_18025);
or U22090 (N_22090,N_19147,N_17139);
nand U22091 (N_22091,N_17525,N_16382);
and U22092 (N_22092,N_19873,N_18940);
or U22093 (N_22093,N_16823,N_17622);
nor U22094 (N_22094,N_18372,N_16733);
nand U22095 (N_22095,N_16611,N_18399);
and U22096 (N_22096,N_18186,N_18175);
or U22097 (N_22097,N_19530,N_17124);
xor U22098 (N_22098,N_16598,N_17593);
xnor U22099 (N_22099,N_15020,N_18984);
or U22100 (N_22100,N_17423,N_16181);
nor U22101 (N_22101,N_16750,N_16456);
nand U22102 (N_22102,N_17433,N_17156);
xnor U22103 (N_22103,N_16639,N_15292);
nor U22104 (N_22104,N_18136,N_19487);
and U22105 (N_22105,N_17316,N_17187);
and U22106 (N_22106,N_18777,N_17898);
nand U22107 (N_22107,N_17009,N_16101);
or U22108 (N_22108,N_16589,N_17329);
nor U22109 (N_22109,N_17281,N_16032);
or U22110 (N_22110,N_18544,N_17062);
and U22111 (N_22111,N_15042,N_17150);
nand U22112 (N_22112,N_16606,N_16696);
or U22113 (N_22113,N_16833,N_15923);
nor U22114 (N_22114,N_15570,N_18895);
and U22115 (N_22115,N_17289,N_17799);
nor U22116 (N_22116,N_18418,N_16528);
and U22117 (N_22117,N_19837,N_19461);
xor U22118 (N_22118,N_19897,N_16842);
nor U22119 (N_22119,N_16824,N_16366);
nand U22120 (N_22120,N_16631,N_19592);
nand U22121 (N_22121,N_16390,N_18378);
or U22122 (N_22122,N_16594,N_16236);
nand U22123 (N_22123,N_17829,N_16105);
xnor U22124 (N_22124,N_15612,N_17449);
nand U22125 (N_22125,N_18309,N_15204);
nand U22126 (N_22126,N_17149,N_16138);
nand U22127 (N_22127,N_16233,N_17987);
nand U22128 (N_22128,N_16318,N_19662);
nand U22129 (N_22129,N_19670,N_17706);
and U22130 (N_22130,N_16992,N_16288);
nor U22131 (N_22131,N_15119,N_15079);
or U22132 (N_22132,N_19894,N_18182);
nand U22133 (N_22133,N_16217,N_19523);
or U22134 (N_22134,N_17932,N_17442);
or U22135 (N_22135,N_19397,N_19584);
nand U22136 (N_22136,N_18109,N_18922);
nand U22137 (N_22137,N_16006,N_17840);
and U22138 (N_22138,N_17226,N_16325);
nor U22139 (N_22139,N_16673,N_17314);
and U22140 (N_22140,N_16728,N_19423);
nand U22141 (N_22141,N_15427,N_19869);
or U22142 (N_22142,N_18246,N_18668);
or U22143 (N_22143,N_16628,N_19094);
nor U22144 (N_22144,N_17494,N_16675);
nand U22145 (N_22145,N_19401,N_16204);
nor U22146 (N_22146,N_17780,N_19784);
nor U22147 (N_22147,N_18202,N_15313);
nor U22148 (N_22148,N_15549,N_15787);
nand U22149 (N_22149,N_16346,N_17980);
and U22150 (N_22150,N_19393,N_18396);
or U22151 (N_22151,N_19484,N_15667);
nand U22152 (N_22152,N_19851,N_17625);
nor U22153 (N_22153,N_17131,N_19309);
nor U22154 (N_22154,N_16603,N_19091);
and U22155 (N_22155,N_19820,N_19497);
xor U22156 (N_22156,N_17235,N_16061);
or U22157 (N_22157,N_18086,N_19104);
nand U22158 (N_22158,N_17120,N_18928);
nor U22159 (N_22159,N_17098,N_19608);
nand U22160 (N_22160,N_18367,N_16364);
nor U22161 (N_22161,N_16869,N_17339);
and U22162 (N_22162,N_17786,N_18735);
nand U22163 (N_22163,N_18860,N_17564);
and U22164 (N_22164,N_15416,N_17642);
and U22165 (N_22165,N_16430,N_15982);
nand U22166 (N_22166,N_16907,N_17126);
nor U22167 (N_22167,N_16571,N_17951);
or U22168 (N_22168,N_15941,N_19385);
or U22169 (N_22169,N_19361,N_17752);
or U22170 (N_22170,N_16004,N_19199);
or U22171 (N_22171,N_17394,N_19704);
and U22172 (N_22172,N_19519,N_18802);
nor U22173 (N_22173,N_19070,N_17173);
and U22174 (N_22174,N_17217,N_19387);
nand U22175 (N_22175,N_18875,N_17267);
or U22176 (N_22176,N_19557,N_19674);
nand U22177 (N_22177,N_16342,N_16896);
xnor U22178 (N_22178,N_16885,N_18524);
xor U22179 (N_22179,N_19428,N_16248);
nand U22180 (N_22180,N_17350,N_15751);
nor U22181 (N_22181,N_17756,N_15461);
and U22182 (N_22182,N_16414,N_18036);
and U22183 (N_22183,N_18253,N_17753);
or U22184 (N_22184,N_15981,N_15304);
nand U22185 (N_22185,N_18995,N_19651);
nor U22186 (N_22186,N_18919,N_19463);
or U22187 (N_22187,N_16385,N_19258);
or U22188 (N_22188,N_17614,N_19118);
nand U22189 (N_22189,N_19316,N_17580);
xor U22190 (N_22190,N_17134,N_18483);
xor U22191 (N_22191,N_17701,N_16960);
xnor U22192 (N_22192,N_19978,N_19881);
or U22193 (N_22193,N_17671,N_16507);
nand U22194 (N_22194,N_18145,N_19739);
xor U22195 (N_22195,N_18672,N_19437);
or U22196 (N_22196,N_18849,N_15422);
xnor U22197 (N_22197,N_16201,N_17930);
and U22198 (N_22198,N_16136,N_19628);
and U22199 (N_22199,N_16950,N_19429);
nor U22200 (N_22200,N_17590,N_15873);
or U22201 (N_22201,N_19532,N_15958);
or U22202 (N_22202,N_15531,N_16831);
nor U22203 (N_22203,N_15806,N_16582);
nor U22204 (N_22204,N_17386,N_19443);
or U22205 (N_22205,N_16848,N_19386);
nor U22206 (N_22206,N_17890,N_16667);
and U22207 (N_22207,N_18196,N_16077);
and U22208 (N_22208,N_19184,N_17929);
or U22209 (N_22209,N_16139,N_17801);
or U22210 (N_22210,N_19926,N_19076);
nor U22211 (N_22211,N_18336,N_17048);
nand U22212 (N_22212,N_17122,N_16685);
and U22213 (N_22213,N_19882,N_16001);
and U22214 (N_22214,N_17145,N_15229);
nor U22215 (N_22215,N_17242,N_17568);
nand U22216 (N_22216,N_17462,N_18062);
nor U22217 (N_22217,N_15956,N_15890);
and U22218 (N_22218,N_17495,N_15657);
and U22219 (N_22219,N_15117,N_16174);
or U22220 (N_22220,N_19573,N_15381);
or U22221 (N_22221,N_15201,N_17684);
and U22222 (N_22222,N_19859,N_16470);
and U22223 (N_22223,N_16943,N_18566);
or U22224 (N_22224,N_18185,N_15429);
and U22225 (N_22225,N_17252,N_15663);
nand U22226 (N_22226,N_19701,N_16033);
nand U22227 (N_22227,N_18911,N_18005);
or U22228 (N_22228,N_19336,N_17737);
nand U22229 (N_22229,N_19005,N_17793);
and U22230 (N_22230,N_18350,N_17768);
or U22231 (N_22231,N_19332,N_15898);
xnor U22232 (N_22232,N_16158,N_15089);
or U22233 (N_22233,N_18128,N_16222);
nand U22234 (N_22234,N_17055,N_16210);
nand U22235 (N_22235,N_17927,N_16244);
or U22236 (N_22236,N_15686,N_17056);
nor U22237 (N_22237,N_16909,N_15007);
nand U22238 (N_22238,N_16730,N_16431);
xor U22239 (N_22239,N_15484,N_17548);
nand U22240 (N_22240,N_19263,N_15250);
nor U22241 (N_22241,N_18938,N_15992);
nor U22242 (N_22242,N_15012,N_19447);
or U22243 (N_22243,N_15463,N_19383);
nand U22244 (N_22244,N_19965,N_15844);
nand U22245 (N_22245,N_19210,N_18817);
and U22246 (N_22246,N_16041,N_15516);
or U22247 (N_22247,N_15393,N_18743);
nor U22248 (N_22248,N_15180,N_16415);
xnor U22249 (N_22249,N_19398,N_19890);
or U22250 (N_22250,N_15413,N_19697);
nand U22251 (N_22251,N_18055,N_18839);
or U22252 (N_22252,N_17049,N_15718);
and U22253 (N_22253,N_18962,N_18010);
and U22254 (N_22254,N_18660,N_18028);
nor U22255 (N_22255,N_15335,N_16686);
and U22256 (N_22256,N_15869,N_17960);
and U22257 (N_22257,N_19349,N_19663);
and U22258 (N_22258,N_17366,N_19681);
and U22259 (N_22259,N_18333,N_18966);
nand U22260 (N_22260,N_15147,N_19521);
or U22261 (N_22261,N_15396,N_15170);
or U22262 (N_22262,N_19814,N_17986);
or U22263 (N_22263,N_15738,N_15344);
or U22264 (N_22264,N_17113,N_17729);
nor U22265 (N_22265,N_17294,N_15939);
nand U22266 (N_22266,N_15133,N_15968);
or U22267 (N_22267,N_18341,N_17258);
nand U22268 (N_22268,N_16074,N_18265);
nand U22269 (N_22269,N_15987,N_17059);
and U22270 (N_22270,N_17269,N_17904);
nor U22271 (N_22271,N_19902,N_18469);
or U22272 (N_22272,N_19705,N_19266);
nor U22273 (N_22273,N_17852,N_16948);
and U22274 (N_22274,N_16292,N_18811);
and U22275 (N_22275,N_17305,N_19030);
nand U22276 (N_22276,N_16042,N_15877);
nor U22277 (N_22277,N_18492,N_18296);
and U22278 (N_22278,N_17195,N_15401);
and U22279 (N_22279,N_18087,N_16969);
and U22280 (N_22280,N_16716,N_18993);
or U22281 (N_22281,N_16143,N_16084);
nand U22282 (N_22282,N_19480,N_17341);
and U22283 (N_22283,N_16634,N_19529);
xor U22284 (N_22284,N_18489,N_16879);
nor U22285 (N_22285,N_19684,N_15742);
or U22286 (N_22286,N_17681,N_16887);
and U22287 (N_22287,N_16260,N_18826);
nor U22288 (N_22288,N_15290,N_17321);
nand U22289 (N_22289,N_19377,N_15297);
xnor U22290 (N_22290,N_15596,N_19655);
nand U22291 (N_22291,N_18444,N_18766);
and U22292 (N_22292,N_17964,N_16011);
and U22293 (N_22293,N_18748,N_16250);
xor U22294 (N_22294,N_18650,N_18496);
nor U22295 (N_22295,N_17888,N_16339);
nor U22296 (N_22296,N_16048,N_15448);
nor U22297 (N_22297,N_16791,N_19693);
nand U22298 (N_22298,N_16393,N_18118);
nand U22299 (N_22299,N_15571,N_18075);
or U22300 (N_22300,N_16180,N_19992);
xnor U22301 (N_22301,N_18868,N_16695);
nand U22302 (N_22302,N_18709,N_19998);
nand U22303 (N_22303,N_17115,N_16671);
nor U22304 (N_22304,N_19755,N_18947);
and U22305 (N_22305,N_15566,N_17620);
or U22306 (N_22306,N_16604,N_17320);
or U22307 (N_22307,N_19804,N_15903);
and U22308 (N_22308,N_18942,N_16491);
nor U22309 (N_22309,N_17830,N_15955);
or U22310 (N_22310,N_15534,N_19097);
and U22311 (N_22311,N_18441,N_18631);
xnor U22312 (N_22312,N_16802,N_18040);
or U22313 (N_22313,N_15838,N_19107);
xnor U22314 (N_22314,N_17292,N_18804);
or U22315 (N_22315,N_18335,N_18877);
and U22316 (N_22316,N_18530,N_19993);
nand U22317 (N_22317,N_18756,N_18426);
nand U22318 (N_22318,N_15296,N_16786);
nand U22319 (N_22319,N_19893,N_18284);
nor U22320 (N_22320,N_17736,N_18715);
and U22321 (N_22321,N_17764,N_17894);
nor U22322 (N_22322,N_16000,N_19346);
nand U22323 (N_22323,N_17985,N_18795);
and U22324 (N_22324,N_19740,N_18112);
or U22325 (N_22325,N_19924,N_15248);
nor U22326 (N_22326,N_18407,N_16211);
nor U22327 (N_22327,N_19616,N_18148);
or U22328 (N_22328,N_16016,N_17051);
nand U22329 (N_22329,N_17613,N_19412);
or U22330 (N_22330,N_19225,N_15521);
and U22331 (N_22331,N_15875,N_16806);
nor U22332 (N_22332,N_17393,N_15897);
xnor U22333 (N_22333,N_18233,N_16241);
nor U22334 (N_22334,N_15481,N_18997);
or U22335 (N_22335,N_17577,N_17050);
xnor U22336 (N_22336,N_17479,N_18397);
nor U22337 (N_22337,N_17138,N_16163);
and U22338 (N_22338,N_16955,N_18513);
or U22339 (N_22339,N_17911,N_18980);
and U22340 (N_22340,N_15218,N_15701);
nor U22341 (N_22341,N_15868,N_17791);
or U22342 (N_22342,N_17534,N_15979);
nor U22343 (N_22343,N_19096,N_16102);
and U22344 (N_22344,N_18315,N_17385);
nor U22345 (N_22345,N_19084,N_15280);
or U22346 (N_22346,N_17362,N_17384);
nor U22347 (N_22347,N_16747,N_15972);
and U22348 (N_22348,N_19314,N_18853);
and U22349 (N_22349,N_16396,N_16489);
nor U22350 (N_22350,N_15870,N_18045);
and U22351 (N_22351,N_16329,N_15095);
or U22352 (N_22352,N_16268,N_19865);
xor U22353 (N_22353,N_19795,N_16020);
and U22354 (N_22354,N_15114,N_18917);
or U22355 (N_22355,N_16185,N_16282);
nor U22356 (N_22356,N_18638,N_18671);
nand U22357 (N_22357,N_18510,N_19254);
nor U22358 (N_22358,N_19023,N_17351);
nand U22359 (N_22359,N_16398,N_16874);
nand U22360 (N_22360,N_19909,N_16765);
nor U22361 (N_22361,N_18484,N_17012);
nand U22362 (N_22362,N_19322,N_15703);
or U22363 (N_22363,N_18787,N_19604);
nor U22364 (N_22364,N_15978,N_19055);
or U22365 (N_22365,N_19606,N_16274);
or U22366 (N_22366,N_15205,N_19043);
nor U22367 (N_22367,N_16112,N_17774);
xnor U22368 (N_22368,N_18359,N_17744);
or U22369 (N_22369,N_15459,N_15146);
nor U22370 (N_22370,N_19553,N_17806);
or U22371 (N_22371,N_18215,N_15836);
or U22372 (N_22372,N_18127,N_16924);
nor U22373 (N_22373,N_19045,N_18002);
or U22374 (N_22374,N_18763,N_19547);
nor U22375 (N_22375,N_16043,N_16681);
nand U22376 (N_22376,N_17646,N_18209);
nor U22377 (N_22377,N_16280,N_15569);
nor U22378 (N_22378,N_17691,N_19031);
and U22379 (N_22379,N_15720,N_19808);
or U22380 (N_22380,N_15216,N_16535);
and U22381 (N_22381,N_18674,N_18812);
nand U22382 (N_22382,N_16073,N_19294);
xnor U22383 (N_22383,N_15828,N_16925);
and U22384 (N_22384,N_15722,N_18528);
or U22385 (N_22385,N_19121,N_15129);
nor U22386 (N_22386,N_18153,N_18990);
or U22387 (N_22387,N_15656,N_15430);
or U22388 (N_22388,N_19613,N_15794);
nor U22389 (N_22389,N_15456,N_17812);
or U22390 (N_22390,N_15260,N_17697);
or U22391 (N_22391,N_15231,N_17992);
nor U22392 (N_22392,N_19365,N_16861);
nand U22393 (N_22393,N_18032,N_15040);
xnor U22394 (N_22394,N_19602,N_15261);
or U22395 (N_22395,N_18557,N_15428);
and U22396 (N_22396,N_16098,N_16843);
and U22397 (N_22397,N_19550,N_19297);
nor U22398 (N_22398,N_19082,N_17451);
and U22399 (N_22399,N_19815,N_15402);
xor U22400 (N_22400,N_18348,N_16213);
nor U22401 (N_22401,N_16612,N_17711);
and U22402 (N_22402,N_16472,N_17206);
nand U22403 (N_22403,N_16760,N_17823);
or U22404 (N_22404,N_18731,N_15023);
or U22405 (N_22405,N_17387,N_18363);
nor U22406 (N_22406,N_15281,N_18824);
and U22407 (N_22407,N_19912,N_19720);
or U22408 (N_22408,N_15207,N_15447);
nand U22409 (N_22409,N_17110,N_15918);
and U22410 (N_22410,N_19489,N_15840);
or U22411 (N_22411,N_19027,N_18301);
nand U22412 (N_22412,N_19611,N_15219);
nand U22413 (N_22413,N_17400,N_17811);
nor U22414 (N_22414,N_19240,N_16648);
and U22415 (N_22415,N_18213,N_15685);
nand U22416 (N_22416,N_19587,N_17309);
and U22417 (N_22417,N_16516,N_18750);
xor U22418 (N_22418,N_19797,N_17148);
or U22419 (N_22419,N_18346,N_19950);
nor U22420 (N_22420,N_18790,N_15943);
or U22421 (N_22421,N_18261,N_17802);
xor U22422 (N_22422,N_19866,N_17718);
or U22423 (N_22423,N_15878,N_18792);
and U22424 (N_22424,N_16106,N_18095);
or U22425 (N_22425,N_17291,N_19174);
nand U22426 (N_22426,N_17130,N_19151);
nand U22427 (N_22427,N_15695,N_18894);
and U22428 (N_22428,N_16123,N_18932);
or U22429 (N_22429,N_15575,N_19860);
and U22430 (N_22430,N_17966,N_16994);
or U22431 (N_22431,N_16337,N_15149);
nor U22432 (N_22432,N_17475,N_16759);
nor U22433 (N_22433,N_18653,N_18620);
nor U22434 (N_22434,N_16220,N_18999);
nand U22435 (N_22435,N_15693,N_17365);
nand U22436 (N_22436,N_17952,N_15406);
xor U22437 (N_22437,N_16135,N_16170);
and U22438 (N_22438,N_16478,N_17000);
xor U22439 (N_22439,N_19568,N_15847);
and U22440 (N_22440,N_16693,N_19320);
or U22441 (N_22441,N_19809,N_19984);
and U22442 (N_22442,N_17923,N_19700);
xnor U22443 (N_22443,N_19908,N_19175);
and U22444 (N_22444,N_18867,N_16764);
or U22445 (N_22445,N_19566,N_19888);
or U22446 (N_22446,N_19271,N_19976);
nand U22447 (N_22447,N_15414,N_18422);
nand U22448 (N_22448,N_17937,N_15162);
or U22449 (N_22449,N_18081,N_15489);
and U22450 (N_22450,N_19941,N_19916);
nand U22451 (N_22451,N_16087,N_19764);
and U22452 (N_22452,N_18688,N_19178);
nor U22453 (N_22453,N_19794,N_15883);
and U22454 (N_22454,N_17396,N_19318);
or U22455 (N_22455,N_16570,N_16609);
nor U22456 (N_22456,N_18147,N_19050);
nor U22457 (N_22457,N_15908,N_17308);
nor U22458 (N_22458,N_17641,N_17868);
nor U22459 (N_22459,N_17058,N_17782);
nor U22460 (N_22460,N_17746,N_18155);
xor U22461 (N_22461,N_19247,N_16977);
xnor U22462 (N_22462,N_16505,N_16593);
or U22463 (N_22463,N_15317,N_15980);
nor U22464 (N_22464,N_16945,N_18347);
xnor U22465 (N_22465,N_17850,N_19567);
or U22466 (N_22466,N_19406,N_17893);
nor U22467 (N_22467,N_18900,N_15035);
or U22468 (N_22468,N_15623,N_19936);
and U22469 (N_22469,N_18840,N_15594);
nor U22470 (N_22470,N_18835,N_16409);
nand U22471 (N_22471,N_16355,N_17910);
or U22472 (N_22472,N_15341,N_16262);
xor U22473 (N_22473,N_16694,N_15544);
and U22474 (N_22474,N_18420,N_19388);
and U22475 (N_22475,N_16014,N_15565);
or U22476 (N_22476,N_15186,N_18591);
nor U22477 (N_22477,N_19770,N_16726);
and U22478 (N_22478,N_17527,N_17618);
and U22479 (N_22479,N_15328,N_19061);
or U22480 (N_22480,N_17270,N_15606);
nand U22481 (N_22481,N_18452,N_15614);
nand U22482 (N_22482,N_15148,N_15697);
and U22483 (N_22483,N_18503,N_18532);
or U22484 (N_22484,N_18994,N_16191);
or U22485 (N_22485,N_19618,N_16092);
or U22486 (N_22486,N_17907,N_15266);
and U22487 (N_22487,N_16971,N_18749);
or U22488 (N_22488,N_16376,N_17651);
nor U22489 (N_22489,N_15795,N_16071);
or U22490 (N_22490,N_15444,N_16116);
nand U22491 (N_22491,N_16188,N_18076);
and U22492 (N_22492,N_16497,N_16564);
or U22493 (N_22493,N_16068,N_16647);
and U22494 (N_22494,N_16550,N_18698);
or U22495 (N_22495,N_17598,N_17238);
nand U22496 (N_22496,N_19932,N_15601);
xor U22497 (N_22497,N_15200,N_15754);
or U22498 (N_22498,N_17179,N_19360);
nor U22499 (N_22499,N_18228,N_18453);
and U22500 (N_22500,N_15727,N_18977);
or U22501 (N_22501,N_15668,N_18893);
and U22502 (N_22502,N_16010,N_15640);
and U22503 (N_22503,N_16472,N_19435);
nor U22504 (N_22504,N_15843,N_19416);
nand U22505 (N_22505,N_17928,N_17522);
nor U22506 (N_22506,N_16196,N_17930);
nand U22507 (N_22507,N_15690,N_18267);
nor U22508 (N_22508,N_17730,N_19300);
and U22509 (N_22509,N_18145,N_18825);
nor U22510 (N_22510,N_15235,N_17226);
nand U22511 (N_22511,N_17266,N_19591);
nand U22512 (N_22512,N_19808,N_18509);
nand U22513 (N_22513,N_19877,N_15347);
and U22514 (N_22514,N_17127,N_15194);
nand U22515 (N_22515,N_16760,N_16026);
nand U22516 (N_22516,N_15518,N_19646);
xor U22517 (N_22517,N_17152,N_15219);
nor U22518 (N_22518,N_18995,N_16454);
nand U22519 (N_22519,N_15658,N_19199);
nand U22520 (N_22520,N_17611,N_19679);
xor U22521 (N_22521,N_17219,N_15126);
or U22522 (N_22522,N_16419,N_19563);
or U22523 (N_22523,N_16038,N_17982);
xor U22524 (N_22524,N_19797,N_19197);
and U22525 (N_22525,N_19407,N_15686);
and U22526 (N_22526,N_19902,N_19937);
nor U22527 (N_22527,N_15909,N_15151);
nand U22528 (N_22528,N_15103,N_17399);
or U22529 (N_22529,N_17548,N_19439);
nand U22530 (N_22530,N_16690,N_16763);
nor U22531 (N_22531,N_18728,N_18533);
nor U22532 (N_22532,N_19241,N_15182);
and U22533 (N_22533,N_15932,N_18148);
nor U22534 (N_22534,N_15256,N_19075);
xor U22535 (N_22535,N_16444,N_19262);
and U22536 (N_22536,N_18821,N_16748);
nor U22537 (N_22537,N_18636,N_15139);
nand U22538 (N_22538,N_19995,N_17733);
nand U22539 (N_22539,N_18608,N_17816);
and U22540 (N_22540,N_19045,N_15061);
or U22541 (N_22541,N_19945,N_15452);
nand U22542 (N_22542,N_16635,N_19871);
and U22543 (N_22543,N_17381,N_16547);
xnor U22544 (N_22544,N_16228,N_17611);
nor U22545 (N_22545,N_16602,N_15615);
and U22546 (N_22546,N_15024,N_15297);
or U22547 (N_22547,N_17954,N_18790);
nor U22548 (N_22548,N_16379,N_15387);
or U22549 (N_22549,N_19729,N_18735);
nor U22550 (N_22550,N_15203,N_15065);
and U22551 (N_22551,N_18624,N_15296);
nand U22552 (N_22552,N_15501,N_15127);
nor U22553 (N_22553,N_15406,N_15096);
or U22554 (N_22554,N_15693,N_17401);
or U22555 (N_22555,N_19613,N_15026);
or U22556 (N_22556,N_16943,N_16609);
or U22557 (N_22557,N_17983,N_16745);
nor U22558 (N_22558,N_17494,N_15133);
nor U22559 (N_22559,N_18004,N_15713);
nor U22560 (N_22560,N_18700,N_18078);
nand U22561 (N_22561,N_16489,N_15729);
nor U22562 (N_22562,N_15080,N_18182);
nor U22563 (N_22563,N_18801,N_16787);
nand U22564 (N_22564,N_17818,N_16209);
nand U22565 (N_22565,N_17976,N_16598);
nand U22566 (N_22566,N_16986,N_15139);
or U22567 (N_22567,N_18749,N_19104);
nand U22568 (N_22568,N_18947,N_18422);
and U22569 (N_22569,N_15715,N_15223);
or U22570 (N_22570,N_17110,N_18514);
or U22571 (N_22571,N_15500,N_19873);
nand U22572 (N_22572,N_19171,N_17658);
or U22573 (N_22573,N_16760,N_18815);
and U22574 (N_22574,N_18824,N_18338);
nor U22575 (N_22575,N_16833,N_19765);
nor U22576 (N_22576,N_15720,N_15697);
nor U22577 (N_22577,N_19723,N_15656);
and U22578 (N_22578,N_18355,N_17614);
and U22579 (N_22579,N_18028,N_17985);
nor U22580 (N_22580,N_17264,N_15846);
and U22581 (N_22581,N_18444,N_18716);
or U22582 (N_22582,N_19025,N_15779);
nand U22583 (N_22583,N_18958,N_19464);
xor U22584 (N_22584,N_19218,N_16161);
nor U22585 (N_22585,N_19798,N_18920);
xor U22586 (N_22586,N_15115,N_16009);
nand U22587 (N_22587,N_18372,N_19330);
or U22588 (N_22588,N_17386,N_16011);
nor U22589 (N_22589,N_18194,N_15882);
nand U22590 (N_22590,N_15473,N_17023);
xnor U22591 (N_22591,N_15429,N_18478);
xnor U22592 (N_22592,N_15579,N_15760);
nand U22593 (N_22593,N_15042,N_18418);
xnor U22594 (N_22594,N_15792,N_15342);
xnor U22595 (N_22595,N_18629,N_15476);
and U22596 (N_22596,N_15745,N_16335);
and U22597 (N_22597,N_18696,N_15086);
nor U22598 (N_22598,N_19282,N_19565);
xor U22599 (N_22599,N_18519,N_15716);
nand U22600 (N_22600,N_18724,N_19030);
and U22601 (N_22601,N_19143,N_17057);
xor U22602 (N_22602,N_18928,N_19307);
and U22603 (N_22603,N_15349,N_15714);
and U22604 (N_22604,N_17691,N_18631);
and U22605 (N_22605,N_17457,N_18434);
and U22606 (N_22606,N_16019,N_16951);
or U22607 (N_22607,N_17472,N_18247);
and U22608 (N_22608,N_18179,N_17574);
nand U22609 (N_22609,N_16053,N_15052);
and U22610 (N_22610,N_19433,N_19696);
or U22611 (N_22611,N_16488,N_15683);
nand U22612 (N_22612,N_18368,N_19003);
xor U22613 (N_22613,N_15649,N_15295);
or U22614 (N_22614,N_17178,N_17193);
and U22615 (N_22615,N_15298,N_19186);
and U22616 (N_22616,N_16740,N_16528);
or U22617 (N_22617,N_18013,N_17374);
xor U22618 (N_22618,N_19554,N_16071);
nor U22619 (N_22619,N_19278,N_17990);
xnor U22620 (N_22620,N_19538,N_18986);
and U22621 (N_22621,N_16522,N_15517);
or U22622 (N_22622,N_18783,N_17485);
nand U22623 (N_22623,N_17058,N_16521);
or U22624 (N_22624,N_17101,N_15158);
or U22625 (N_22625,N_15209,N_17417);
xor U22626 (N_22626,N_19492,N_18544);
and U22627 (N_22627,N_15644,N_18439);
nor U22628 (N_22628,N_19351,N_16990);
and U22629 (N_22629,N_15947,N_17135);
nand U22630 (N_22630,N_17056,N_15160);
nor U22631 (N_22631,N_15722,N_19972);
or U22632 (N_22632,N_16054,N_18900);
nor U22633 (N_22633,N_19715,N_18410);
nand U22634 (N_22634,N_19288,N_18986);
nand U22635 (N_22635,N_18996,N_19319);
or U22636 (N_22636,N_16834,N_15940);
nand U22637 (N_22637,N_18344,N_19018);
nand U22638 (N_22638,N_17273,N_19330);
nand U22639 (N_22639,N_16958,N_15628);
and U22640 (N_22640,N_15021,N_17374);
nand U22641 (N_22641,N_19479,N_18879);
nand U22642 (N_22642,N_16089,N_18772);
xnor U22643 (N_22643,N_15765,N_17616);
and U22644 (N_22644,N_17583,N_17481);
and U22645 (N_22645,N_16402,N_16269);
and U22646 (N_22646,N_18839,N_19603);
or U22647 (N_22647,N_16182,N_19465);
nand U22648 (N_22648,N_17935,N_19112);
or U22649 (N_22649,N_17445,N_18503);
or U22650 (N_22650,N_16839,N_15476);
xor U22651 (N_22651,N_15231,N_15158);
and U22652 (N_22652,N_15163,N_17287);
xnor U22653 (N_22653,N_15992,N_18547);
and U22654 (N_22654,N_15953,N_17758);
or U22655 (N_22655,N_16497,N_16678);
nand U22656 (N_22656,N_17726,N_17500);
or U22657 (N_22657,N_18371,N_15589);
nand U22658 (N_22658,N_17540,N_15174);
and U22659 (N_22659,N_19786,N_17536);
or U22660 (N_22660,N_19321,N_16369);
or U22661 (N_22661,N_18501,N_15674);
and U22662 (N_22662,N_17856,N_17194);
and U22663 (N_22663,N_15640,N_18906);
xor U22664 (N_22664,N_18704,N_19773);
or U22665 (N_22665,N_15578,N_19495);
or U22666 (N_22666,N_16600,N_16601);
nor U22667 (N_22667,N_17446,N_17154);
and U22668 (N_22668,N_16339,N_19685);
and U22669 (N_22669,N_17406,N_17059);
nand U22670 (N_22670,N_15838,N_16012);
xnor U22671 (N_22671,N_17453,N_17969);
nor U22672 (N_22672,N_17039,N_16696);
or U22673 (N_22673,N_18970,N_17488);
nor U22674 (N_22674,N_19873,N_19098);
or U22675 (N_22675,N_16065,N_15951);
nand U22676 (N_22676,N_19179,N_17373);
nor U22677 (N_22677,N_18047,N_18897);
or U22678 (N_22678,N_18160,N_18785);
or U22679 (N_22679,N_19077,N_15992);
or U22680 (N_22680,N_15836,N_16587);
nand U22681 (N_22681,N_16309,N_16841);
and U22682 (N_22682,N_15793,N_19204);
nor U22683 (N_22683,N_15725,N_15416);
and U22684 (N_22684,N_17296,N_17823);
nor U22685 (N_22685,N_19781,N_18776);
or U22686 (N_22686,N_18781,N_17092);
and U22687 (N_22687,N_19210,N_15076);
and U22688 (N_22688,N_17791,N_19749);
or U22689 (N_22689,N_17485,N_18935);
nand U22690 (N_22690,N_16323,N_17253);
nor U22691 (N_22691,N_17645,N_19584);
nor U22692 (N_22692,N_18363,N_17197);
and U22693 (N_22693,N_16519,N_19873);
nor U22694 (N_22694,N_15202,N_18275);
nand U22695 (N_22695,N_18098,N_19652);
or U22696 (N_22696,N_19503,N_18259);
nand U22697 (N_22697,N_19151,N_15477);
nor U22698 (N_22698,N_19754,N_17586);
xor U22699 (N_22699,N_17336,N_18079);
xnor U22700 (N_22700,N_19256,N_16007);
and U22701 (N_22701,N_17634,N_17771);
nor U22702 (N_22702,N_19930,N_15872);
xnor U22703 (N_22703,N_17258,N_17022);
nor U22704 (N_22704,N_16829,N_17457);
and U22705 (N_22705,N_18690,N_18524);
and U22706 (N_22706,N_17475,N_17137);
or U22707 (N_22707,N_17295,N_16658);
and U22708 (N_22708,N_16086,N_15981);
and U22709 (N_22709,N_17742,N_15457);
or U22710 (N_22710,N_17779,N_15553);
nor U22711 (N_22711,N_15665,N_18300);
and U22712 (N_22712,N_15390,N_18867);
and U22713 (N_22713,N_16625,N_15675);
and U22714 (N_22714,N_16967,N_19239);
and U22715 (N_22715,N_18370,N_17270);
xnor U22716 (N_22716,N_19780,N_15552);
and U22717 (N_22717,N_15582,N_18470);
and U22718 (N_22718,N_16033,N_19299);
xor U22719 (N_22719,N_15125,N_16697);
and U22720 (N_22720,N_19493,N_18891);
nand U22721 (N_22721,N_18694,N_16833);
or U22722 (N_22722,N_16503,N_17685);
or U22723 (N_22723,N_16781,N_18939);
or U22724 (N_22724,N_17689,N_16528);
nor U22725 (N_22725,N_15911,N_15539);
nor U22726 (N_22726,N_15654,N_15133);
and U22727 (N_22727,N_19875,N_16771);
xor U22728 (N_22728,N_16812,N_15219);
and U22729 (N_22729,N_17162,N_18623);
xnor U22730 (N_22730,N_18364,N_19155);
nand U22731 (N_22731,N_15581,N_17627);
and U22732 (N_22732,N_16762,N_17607);
or U22733 (N_22733,N_17361,N_15966);
nor U22734 (N_22734,N_17925,N_16143);
and U22735 (N_22735,N_16653,N_16649);
nor U22736 (N_22736,N_15906,N_18971);
or U22737 (N_22737,N_16340,N_16195);
and U22738 (N_22738,N_19399,N_15375);
xor U22739 (N_22739,N_19086,N_15613);
and U22740 (N_22740,N_18989,N_16430);
and U22741 (N_22741,N_17395,N_18972);
nor U22742 (N_22742,N_16566,N_18482);
or U22743 (N_22743,N_17973,N_19520);
nor U22744 (N_22744,N_17859,N_15685);
xnor U22745 (N_22745,N_17196,N_19805);
and U22746 (N_22746,N_18668,N_19809);
and U22747 (N_22747,N_18158,N_17343);
or U22748 (N_22748,N_15679,N_19123);
nor U22749 (N_22749,N_16547,N_18641);
nand U22750 (N_22750,N_16358,N_19954);
nand U22751 (N_22751,N_16340,N_15504);
and U22752 (N_22752,N_16690,N_15966);
and U22753 (N_22753,N_17379,N_17487);
nor U22754 (N_22754,N_19155,N_19117);
nand U22755 (N_22755,N_16261,N_16834);
nand U22756 (N_22756,N_15668,N_15402);
or U22757 (N_22757,N_19701,N_15344);
nor U22758 (N_22758,N_19980,N_15716);
or U22759 (N_22759,N_16337,N_16074);
xnor U22760 (N_22760,N_15988,N_16110);
or U22761 (N_22761,N_15645,N_17599);
nand U22762 (N_22762,N_17119,N_18478);
xnor U22763 (N_22763,N_16383,N_15501);
nor U22764 (N_22764,N_17979,N_15699);
or U22765 (N_22765,N_17561,N_18436);
xnor U22766 (N_22766,N_17526,N_15544);
or U22767 (N_22767,N_15834,N_17465);
nor U22768 (N_22768,N_16472,N_18912);
nor U22769 (N_22769,N_16837,N_19870);
and U22770 (N_22770,N_19800,N_17948);
and U22771 (N_22771,N_17811,N_16109);
nand U22772 (N_22772,N_18423,N_16049);
or U22773 (N_22773,N_16694,N_18561);
or U22774 (N_22774,N_15332,N_16609);
and U22775 (N_22775,N_16782,N_19651);
nor U22776 (N_22776,N_18840,N_19475);
xnor U22777 (N_22777,N_15195,N_15317);
nand U22778 (N_22778,N_19260,N_16010);
and U22779 (N_22779,N_17761,N_19048);
nor U22780 (N_22780,N_16721,N_16649);
nor U22781 (N_22781,N_19390,N_19544);
nor U22782 (N_22782,N_19435,N_15459);
nor U22783 (N_22783,N_16175,N_17187);
and U22784 (N_22784,N_16416,N_15708);
and U22785 (N_22785,N_19836,N_15606);
xnor U22786 (N_22786,N_19302,N_19777);
or U22787 (N_22787,N_16101,N_16608);
xor U22788 (N_22788,N_18951,N_17769);
and U22789 (N_22789,N_15530,N_17547);
nor U22790 (N_22790,N_18562,N_18782);
and U22791 (N_22791,N_17250,N_19345);
nand U22792 (N_22792,N_16008,N_19974);
or U22793 (N_22793,N_19889,N_17438);
nor U22794 (N_22794,N_15392,N_18128);
nand U22795 (N_22795,N_19570,N_15968);
or U22796 (N_22796,N_15254,N_15110);
or U22797 (N_22797,N_16979,N_19055);
and U22798 (N_22798,N_19900,N_16389);
nor U22799 (N_22799,N_16790,N_16429);
nor U22800 (N_22800,N_17001,N_17610);
xnor U22801 (N_22801,N_18925,N_19787);
nand U22802 (N_22802,N_17787,N_19160);
and U22803 (N_22803,N_18754,N_15640);
or U22804 (N_22804,N_17506,N_16168);
xnor U22805 (N_22805,N_19170,N_19213);
nand U22806 (N_22806,N_18227,N_19158);
nor U22807 (N_22807,N_17845,N_15502);
or U22808 (N_22808,N_15694,N_19421);
and U22809 (N_22809,N_15203,N_18425);
nor U22810 (N_22810,N_18157,N_18518);
xor U22811 (N_22811,N_18352,N_17475);
nand U22812 (N_22812,N_17534,N_18612);
nor U22813 (N_22813,N_19636,N_16620);
nand U22814 (N_22814,N_18904,N_17019);
or U22815 (N_22815,N_15371,N_18541);
nor U22816 (N_22816,N_19217,N_19730);
nor U22817 (N_22817,N_18766,N_15184);
nand U22818 (N_22818,N_19897,N_17333);
and U22819 (N_22819,N_17027,N_19367);
and U22820 (N_22820,N_19256,N_18074);
or U22821 (N_22821,N_19148,N_15145);
xnor U22822 (N_22822,N_15140,N_19821);
nand U22823 (N_22823,N_18083,N_17891);
xor U22824 (N_22824,N_15382,N_15859);
and U22825 (N_22825,N_18845,N_16117);
nor U22826 (N_22826,N_16942,N_15498);
and U22827 (N_22827,N_15947,N_16486);
nor U22828 (N_22828,N_15391,N_18933);
nand U22829 (N_22829,N_16899,N_19923);
nor U22830 (N_22830,N_16228,N_15331);
nand U22831 (N_22831,N_15732,N_17157);
and U22832 (N_22832,N_16801,N_15350);
and U22833 (N_22833,N_19397,N_17380);
nor U22834 (N_22834,N_17697,N_18540);
or U22835 (N_22835,N_17978,N_16148);
xnor U22836 (N_22836,N_17877,N_19740);
xnor U22837 (N_22837,N_16412,N_18706);
or U22838 (N_22838,N_19061,N_19202);
nor U22839 (N_22839,N_19945,N_18890);
and U22840 (N_22840,N_19856,N_17951);
nand U22841 (N_22841,N_15084,N_19520);
xor U22842 (N_22842,N_15563,N_19688);
nor U22843 (N_22843,N_16587,N_19717);
nor U22844 (N_22844,N_19547,N_16372);
xnor U22845 (N_22845,N_19263,N_15665);
nand U22846 (N_22846,N_15417,N_18086);
nand U22847 (N_22847,N_15191,N_17559);
or U22848 (N_22848,N_18536,N_17509);
and U22849 (N_22849,N_18113,N_17987);
nand U22850 (N_22850,N_16412,N_16278);
nor U22851 (N_22851,N_16432,N_16273);
xor U22852 (N_22852,N_15854,N_17314);
nand U22853 (N_22853,N_15673,N_19522);
or U22854 (N_22854,N_17262,N_16210);
and U22855 (N_22855,N_15569,N_19383);
and U22856 (N_22856,N_18632,N_17766);
xor U22857 (N_22857,N_18943,N_18927);
xnor U22858 (N_22858,N_19232,N_16550);
nor U22859 (N_22859,N_16663,N_17205);
and U22860 (N_22860,N_16432,N_17829);
nand U22861 (N_22861,N_19708,N_18878);
or U22862 (N_22862,N_18960,N_16580);
nand U22863 (N_22863,N_18747,N_17794);
nand U22864 (N_22864,N_19995,N_19720);
and U22865 (N_22865,N_15653,N_19329);
xor U22866 (N_22866,N_18374,N_19130);
nand U22867 (N_22867,N_19550,N_18434);
nor U22868 (N_22868,N_17544,N_15479);
and U22869 (N_22869,N_17360,N_17544);
nor U22870 (N_22870,N_16306,N_19125);
nand U22871 (N_22871,N_17729,N_18410);
and U22872 (N_22872,N_17307,N_16996);
or U22873 (N_22873,N_18796,N_19042);
or U22874 (N_22874,N_19762,N_19691);
xor U22875 (N_22875,N_19101,N_19088);
nand U22876 (N_22876,N_18404,N_15859);
xor U22877 (N_22877,N_18043,N_18670);
nor U22878 (N_22878,N_19419,N_16328);
or U22879 (N_22879,N_17726,N_19144);
nand U22880 (N_22880,N_18755,N_16974);
nand U22881 (N_22881,N_19248,N_15024);
nor U22882 (N_22882,N_17898,N_18549);
or U22883 (N_22883,N_15738,N_16975);
or U22884 (N_22884,N_18330,N_18194);
nand U22885 (N_22885,N_15387,N_17385);
or U22886 (N_22886,N_18631,N_16500);
or U22887 (N_22887,N_16641,N_19925);
and U22888 (N_22888,N_17979,N_18189);
and U22889 (N_22889,N_18944,N_19470);
or U22890 (N_22890,N_19276,N_15554);
nand U22891 (N_22891,N_15123,N_19079);
or U22892 (N_22892,N_19429,N_18577);
and U22893 (N_22893,N_18443,N_19229);
nor U22894 (N_22894,N_15069,N_19729);
nand U22895 (N_22895,N_16766,N_15719);
and U22896 (N_22896,N_19249,N_16788);
nor U22897 (N_22897,N_16239,N_16664);
nand U22898 (N_22898,N_18507,N_18622);
or U22899 (N_22899,N_17423,N_19633);
and U22900 (N_22900,N_15764,N_16893);
nor U22901 (N_22901,N_19687,N_18630);
nor U22902 (N_22902,N_18550,N_19418);
and U22903 (N_22903,N_17170,N_16692);
nand U22904 (N_22904,N_18001,N_16454);
xor U22905 (N_22905,N_18023,N_17763);
nor U22906 (N_22906,N_17758,N_19176);
xor U22907 (N_22907,N_17542,N_17200);
nor U22908 (N_22908,N_19729,N_16196);
nand U22909 (N_22909,N_18469,N_18972);
and U22910 (N_22910,N_19246,N_16244);
nand U22911 (N_22911,N_16888,N_17268);
and U22912 (N_22912,N_17207,N_17859);
and U22913 (N_22913,N_17659,N_15864);
and U22914 (N_22914,N_15761,N_19055);
or U22915 (N_22915,N_18546,N_19749);
and U22916 (N_22916,N_18168,N_17731);
xor U22917 (N_22917,N_19575,N_18799);
or U22918 (N_22918,N_19506,N_16856);
nand U22919 (N_22919,N_18105,N_19118);
and U22920 (N_22920,N_16026,N_17744);
nor U22921 (N_22921,N_17324,N_16059);
or U22922 (N_22922,N_18803,N_19129);
and U22923 (N_22923,N_17646,N_18354);
or U22924 (N_22924,N_17662,N_16563);
and U22925 (N_22925,N_15668,N_15215);
nor U22926 (N_22926,N_19811,N_17180);
nand U22927 (N_22927,N_15168,N_17775);
or U22928 (N_22928,N_19104,N_19008);
nand U22929 (N_22929,N_17226,N_16539);
nand U22930 (N_22930,N_16088,N_18791);
and U22931 (N_22931,N_15341,N_17745);
nand U22932 (N_22932,N_15784,N_15400);
and U22933 (N_22933,N_17167,N_17998);
and U22934 (N_22934,N_18545,N_16841);
and U22935 (N_22935,N_16637,N_17143);
and U22936 (N_22936,N_16033,N_16844);
xor U22937 (N_22937,N_18017,N_18808);
nor U22938 (N_22938,N_16997,N_19814);
or U22939 (N_22939,N_19233,N_18911);
or U22940 (N_22940,N_16488,N_16373);
nor U22941 (N_22941,N_16475,N_16198);
nand U22942 (N_22942,N_17885,N_15706);
nor U22943 (N_22943,N_16069,N_17869);
and U22944 (N_22944,N_19597,N_19902);
xnor U22945 (N_22945,N_17149,N_15315);
and U22946 (N_22946,N_17946,N_15573);
nor U22947 (N_22947,N_18335,N_16656);
nor U22948 (N_22948,N_16463,N_17587);
or U22949 (N_22949,N_16061,N_16102);
and U22950 (N_22950,N_16819,N_16616);
and U22951 (N_22951,N_19722,N_18281);
or U22952 (N_22952,N_19341,N_18193);
or U22953 (N_22953,N_19886,N_16611);
nor U22954 (N_22954,N_16585,N_18811);
nand U22955 (N_22955,N_18405,N_15600);
nor U22956 (N_22956,N_16545,N_18922);
nand U22957 (N_22957,N_16532,N_17384);
or U22958 (N_22958,N_19796,N_16397);
nor U22959 (N_22959,N_16030,N_18907);
nand U22960 (N_22960,N_15825,N_19867);
nor U22961 (N_22961,N_17180,N_16101);
and U22962 (N_22962,N_17301,N_19813);
xnor U22963 (N_22963,N_19377,N_16294);
nor U22964 (N_22964,N_19906,N_16293);
nor U22965 (N_22965,N_18917,N_16361);
xor U22966 (N_22966,N_15916,N_19437);
nand U22967 (N_22967,N_15342,N_15016);
and U22968 (N_22968,N_17964,N_15691);
nor U22969 (N_22969,N_17720,N_17986);
and U22970 (N_22970,N_16930,N_15726);
and U22971 (N_22971,N_16674,N_19212);
or U22972 (N_22972,N_19564,N_19221);
nand U22973 (N_22973,N_17031,N_16785);
xnor U22974 (N_22974,N_15944,N_18771);
and U22975 (N_22975,N_19087,N_17510);
nand U22976 (N_22976,N_18577,N_17632);
or U22977 (N_22977,N_19481,N_16991);
nand U22978 (N_22978,N_15756,N_15844);
nor U22979 (N_22979,N_17612,N_17607);
or U22980 (N_22980,N_18215,N_18488);
or U22981 (N_22981,N_15847,N_15493);
and U22982 (N_22982,N_19529,N_15853);
nand U22983 (N_22983,N_19731,N_15380);
nand U22984 (N_22984,N_17402,N_19689);
nand U22985 (N_22985,N_19685,N_17423);
nor U22986 (N_22986,N_17899,N_15026);
or U22987 (N_22987,N_17291,N_18098);
or U22988 (N_22988,N_19584,N_15091);
xor U22989 (N_22989,N_15009,N_15721);
xnor U22990 (N_22990,N_16683,N_18150);
or U22991 (N_22991,N_16659,N_15068);
xor U22992 (N_22992,N_16331,N_16134);
xnor U22993 (N_22993,N_16325,N_18222);
nand U22994 (N_22994,N_17829,N_17835);
and U22995 (N_22995,N_18075,N_19701);
nand U22996 (N_22996,N_16871,N_18793);
and U22997 (N_22997,N_15377,N_17958);
or U22998 (N_22998,N_18015,N_18108);
nor U22999 (N_22999,N_18071,N_19264);
or U23000 (N_23000,N_17919,N_16029);
nor U23001 (N_23001,N_18072,N_15021);
nand U23002 (N_23002,N_17134,N_18850);
or U23003 (N_23003,N_16772,N_15823);
nor U23004 (N_23004,N_17605,N_19650);
and U23005 (N_23005,N_18874,N_15584);
and U23006 (N_23006,N_17468,N_15185);
nand U23007 (N_23007,N_16595,N_16143);
xnor U23008 (N_23008,N_19472,N_17369);
xnor U23009 (N_23009,N_16361,N_19334);
xor U23010 (N_23010,N_18543,N_17456);
or U23011 (N_23011,N_15068,N_16433);
and U23012 (N_23012,N_18068,N_15703);
nand U23013 (N_23013,N_18697,N_15308);
and U23014 (N_23014,N_17616,N_18578);
nor U23015 (N_23015,N_18589,N_16355);
and U23016 (N_23016,N_17019,N_16153);
nand U23017 (N_23017,N_18941,N_15898);
nor U23018 (N_23018,N_15835,N_19240);
or U23019 (N_23019,N_15354,N_16313);
nand U23020 (N_23020,N_15000,N_15600);
and U23021 (N_23021,N_15637,N_19448);
nor U23022 (N_23022,N_19927,N_15733);
nand U23023 (N_23023,N_16926,N_15678);
nor U23024 (N_23024,N_18300,N_17583);
nor U23025 (N_23025,N_18450,N_19583);
and U23026 (N_23026,N_18922,N_16796);
and U23027 (N_23027,N_18518,N_18571);
and U23028 (N_23028,N_18418,N_16406);
or U23029 (N_23029,N_17033,N_17970);
and U23030 (N_23030,N_16980,N_17480);
nor U23031 (N_23031,N_18220,N_15256);
or U23032 (N_23032,N_17889,N_15970);
and U23033 (N_23033,N_19700,N_15362);
or U23034 (N_23034,N_19459,N_18895);
xnor U23035 (N_23035,N_16288,N_16667);
nand U23036 (N_23036,N_18423,N_15088);
or U23037 (N_23037,N_15987,N_17783);
or U23038 (N_23038,N_17317,N_15582);
nor U23039 (N_23039,N_17822,N_17129);
nor U23040 (N_23040,N_19301,N_15427);
and U23041 (N_23041,N_15184,N_15530);
nand U23042 (N_23042,N_15654,N_19288);
xor U23043 (N_23043,N_15435,N_18192);
and U23044 (N_23044,N_15722,N_18898);
nor U23045 (N_23045,N_18856,N_15700);
or U23046 (N_23046,N_18893,N_18789);
nor U23047 (N_23047,N_17451,N_19479);
nor U23048 (N_23048,N_17749,N_15724);
xor U23049 (N_23049,N_17897,N_15569);
or U23050 (N_23050,N_17877,N_18229);
nand U23051 (N_23051,N_19000,N_17462);
xnor U23052 (N_23052,N_18636,N_16577);
or U23053 (N_23053,N_16978,N_18117);
and U23054 (N_23054,N_15848,N_15773);
nor U23055 (N_23055,N_19828,N_16911);
xor U23056 (N_23056,N_16402,N_19092);
nor U23057 (N_23057,N_17144,N_19378);
nand U23058 (N_23058,N_15350,N_17896);
nand U23059 (N_23059,N_19726,N_19908);
and U23060 (N_23060,N_18828,N_15368);
nor U23061 (N_23061,N_19103,N_18406);
nand U23062 (N_23062,N_19001,N_16429);
nand U23063 (N_23063,N_16871,N_16026);
nor U23064 (N_23064,N_17228,N_15889);
nor U23065 (N_23065,N_15958,N_18645);
or U23066 (N_23066,N_15670,N_15773);
nor U23067 (N_23067,N_15238,N_15674);
and U23068 (N_23068,N_15986,N_15738);
or U23069 (N_23069,N_18304,N_16331);
and U23070 (N_23070,N_18198,N_17854);
nand U23071 (N_23071,N_15176,N_19091);
nand U23072 (N_23072,N_16610,N_16058);
and U23073 (N_23073,N_16084,N_19987);
nor U23074 (N_23074,N_19221,N_19678);
and U23075 (N_23075,N_17183,N_19984);
and U23076 (N_23076,N_18100,N_18782);
and U23077 (N_23077,N_15505,N_17741);
and U23078 (N_23078,N_16802,N_19358);
nand U23079 (N_23079,N_17370,N_19282);
nor U23080 (N_23080,N_17884,N_18442);
and U23081 (N_23081,N_15578,N_16558);
nor U23082 (N_23082,N_18130,N_15363);
xnor U23083 (N_23083,N_18969,N_17037);
nand U23084 (N_23084,N_18435,N_19497);
xnor U23085 (N_23085,N_18203,N_15771);
xor U23086 (N_23086,N_16971,N_15428);
nor U23087 (N_23087,N_18165,N_18153);
or U23088 (N_23088,N_16131,N_18267);
nor U23089 (N_23089,N_15709,N_18804);
or U23090 (N_23090,N_16564,N_18030);
nand U23091 (N_23091,N_18871,N_17929);
xor U23092 (N_23092,N_17542,N_19910);
or U23093 (N_23093,N_19887,N_15651);
or U23094 (N_23094,N_17664,N_19303);
nand U23095 (N_23095,N_17475,N_16673);
or U23096 (N_23096,N_15766,N_18326);
nor U23097 (N_23097,N_18810,N_15927);
or U23098 (N_23098,N_15683,N_16243);
or U23099 (N_23099,N_18858,N_18168);
nand U23100 (N_23100,N_17512,N_19541);
nor U23101 (N_23101,N_17939,N_17168);
and U23102 (N_23102,N_18819,N_15979);
nand U23103 (N_23103,N_15787,N_18029);
nor U23104 (N_23104,N_19004,N_19097);
xnor U23105 (N_23105,N_19317,N_16635);
xnor U23106 (N_23106,N_17957,N_16441);
and U23107 (N_23107,N_15868,N_18748);
xor U23108 (N_23108,N_15986,N_15755);
nor U23109 (N_23109,N_18902,N_17553);
nor U23110 (N_23110,N_16917,N_18489);
and U23111 (N_23111,N_18313,N_15902);
and U23112 (N_23112,N_19595,N_19391);
nand U23113 (N_23113,N_16322,N_18616);
nand U23114 (N_23114,N_15719,N_16078);
or U23115 (N_23115,N_19321,N_16395);
or U23116 (N_23116,N_15655,N_18972);
or U23117 (N_23117,N_18783,N_17919);
or U23118 (N_23118,N_15340,N_17815);
and U23119 (N_23119,N_17672,N_17554);
nor U23120 (N_23120,N_15530,N_16343);
xor U23121 (N_23121,N_17420,N_19638);
nor U23122 (N_23122,N_19677,N_17835);
nor U23123 (N_23123,N_15006,N_17360);
nand U23124 (N_23124,N_19954,N_19994);
or U23125 (N_23125,N_15456,N_19018);
and U23126 (N_23126,N_16463,N_15015);
or U23127 (N_23127,N_18491,N_17597);
nand U23128 (N_23128,N_17019,N_17101);
or U23129 (N_23129,N_16134,N_19532);
and U23130 (N_23130,N_17760,N_15987);
nand U23131 (N_23131,N_16011,N_15407);
and U23132 (N_23132,N_16414,N_19820);
nor U23133 (N_23133,N_19844,N_19655);
or U23134 (N_23134,N_19516,N_15263);
or U23135 (N_23135,N_15637,N_15780);
and U23136 (N_23136,N_15702,N_16420);
and U23137 (N_23137,N_19494,N_15249);
and U23138 (N_23138,N_19082,N_18366);
or U23139 (N_23139,N_17241,N_18498);
or U23140 (N_23140,N_19657,N_15343);
nor U23141 (N_23141,N_15191,N_17043);
nand U23142 (N_23142,N_16393,N_15910);
nand U23143 (N_23143,N_15618,N_16651);
and U23144 (N_23144,N_16903,N_15801);
nand U23145 (N_23145,N_15303,N_16191);
and U23146 (N_23146,N_19802,N_17126);
xor U23147 (N_23147,N_15486,N_19447);
and U23148 (N_23148,N_16898,N_15038);
nor U23149 (N_23149,N_18750,N_19549);
and U23150 (N_23150,N_16328,N_16577);
nor U23151 (N_23151,N_15798,N_16903);
or U23152 (N_23152,N_18900,N_19733);
nor U23153 (N_23153,N_15382,N_15544);
xor U23154 (N_23154,N_15106,N_17989);
or U23155 (N_23155,N_16922,N_15390);
nand U23156 (N_23156,N_16516,N_15525);
or U23157 (N_23157,N_16198,N_18293);
and U23158 (N_23158,N_18275,N_19656);
and U23159 (N_23159,N_15193,N_15335);
or U23160 (N_23160,N_15320,N_19089);
nand U23161 (N_23161,N_18675,N_17958);
or U23162 (N_23162,N_17068,N_18308);
nand U23163 (N_23163,N_15006,N_16195);
nor U23164 (N_23164,N_15203,N_15515);
nand U23165 (N_23165,N_17633,N_19936);
nand U23166 (N_23166,N_17201,N_15221);
nand U23167 (N_23167,N_16153,N_16434);
or U23168 (N_23168,N_17063,N_16974);
nand U23169 (N_23169,N_17107,N_16151);
or U23170 (N_23170,N_18073,N_17540);
and U23171 (N_23171,N_19617,N_16461);
xnor U23172 (N_23172,N_17082,N_15012);
xor U23173 (N_23173,N_15093,N_17167);
nor U23174 (N_23174,N_17109,N_17680);
and U23175 (N_23175,N_19929,N_18286);
nand U23176 (N_23176,N_15744,N_18840);
or U23177 (N_23177,N_16393,N_17873);
nor U23178 (N_23178,N_18856,N_16726);
xnor U23179 (N_23179,N_17878,N_18733);
or U23180 (N_23180,N_18298,N_18248);
nand U23181 (N_23181,N_18722,N_19417);
nor U23182 (N_23182,N_18625,N_19345);
nor U23183 (N_23183,N_17913,N_16776);
nor U23184 (N_23184,N_16666,N_18527);
and U23185 (N_23185,N_18990,N_19150);
or U23186 (N_23186,N_15357,N_16079);
nor U23187 (N_23187,N_17152,N_15637);
or U23188 (N_23188,N_15981,N_17063);
and U23189 (N_23189,N_15459,N_15901);
nor U23190 (N_23190,N_15100,N_17434);
nand U23191 (N_23191,N_19247,N_18155);
and U23192 (N_23192,N_15410,N_16378);
or U23193 (N_23193,N_18443,N_16167);
or U23194 (N_23194,N_17796,N_17737);
and U23195 (N_23195,N_17862,N_15966);
and U23196 (N_23196,N_17917,N_16419);
xor U23197 (N_23197,N_15685,N_18150);
or U23198 (N_23198,N_18493,N_18762);
nand U23199 (N_23199,N_16525,N_19339);
nor U23200 (N_23200,N_15221,N_18137);
and U23201 (N_23201,N_18332,N_18407);
or U23202 (N_23202,N_19371,N_17787);
and U23203 (N_23203,N_17765,N_18557);
nor U23204 (N_23204,N_15070,N_18559);
nand U23205 (N_23205,N_19391,N_16840);
or U23206 (N_23206,N_16978,N_18283);
and U23207 (N_23207,N_15312,N_19454);
nand U23208 (N_23208,N_17458,N_16379);
nand U23209 (N_23209,N_16100,N_15402);
xor U23210 (N_23210,N_16186,N_15687);
or U23211 (N_23211,N_17038,N_17504);
nor U23212 (N_23212,N_16521,N_18551);
and U23213 (N_23213,N_18949,N_17121);
or U23214 (N_23214,N_18257,N_16733);
nand U23215 (N_23215,N_16002,N_17636);
nor U23216 (N_23216,N_15213,N_17388);
nand U23217 (N_23217,N_19848,N_17569);
nand U23218 (N_23218,N_17861,N_18506);
and U23219 (N_23219,N_19853,N_15774);
nor U23220 (N_23220,N_17316,N_17454);
xnor U23221 (N_23221,N_15006,N_19173);
or U23222 (N_23222,N_19679,N_19422);
nand U23223 (N_23223,N_16437,N_16093);
or U23224 (N_23224,N_19902,N_19442);
xnor U23225 (N_23225,N_18546,N_18939);
or U23226 (N_23226,N_17434,N_19084);
nand U23227 (N_23227,N_16340,N_15177);
or U23228 (N_23228,N_18549,N_16327);
xor U23229 (N_23229,N_17904,N_16626);
nor U23230 (N_23230,N_16541,N_17205);
nand U23231 (N_23231,N_19440,N_19745);
nand U23232 (N_23232,N_15065,N_16447);
and U23233 (N_23233,N_16465,N_16623);
nand U23234 (N_23234,N_17278,N_17143);
or U23235 (N_23235,N_15573,N_15304);
nor U23236 (N_23236,N_19715,N_18145);
or U23237 (N_23237,N_15938,N_15658);
xnor U23238 (N_23238,N_18433,N_19309);
nand U23239 (N_23239,N_17267,N_17717);
or U23240 (N_23240,N_19814,N_18347);
nor U23241 (N_23241,N_17977,N_18172);
or U23242 (N_23242,N_16887,N_15880);
nand U23243 (N_23243,N_16000,N_19439);
nand U23244 (N_23244,N_15406,N_19263);
or U23245 (N_23245,N_18640,N_16137);
nor U23246 (N_23246,N_17009,N_16022);
xor U23247 (N_23247,N_15141,N_19817);
and U23248 (N_23248,N_18206,N_15594);
nor U23249 (N_23249,N_15739,N_19187);
or U23250 (N_23250,N_16581,N_19938);
nor U23251 (N_23251,N_17599,N_17472);
and U23252 (N_23252,N_15225,N_17243);
nand U23253 (N_23253,N_15830,N_19685);
xor U23254 (N_23254,N_15287,N_15404);
and U23255 (N_23255,N_19380,N_16181);
nand U23256 (N_23256,N_19061,N_16122);
xor U23257 (N_23257,N_18536,N_16495);
and U23258 (N_23258,N_19827,N_15007);
and U23259 (N_23259,N_17965,N_17435);
or U23260 (N_23260,N_17420,N_17615);
or U23261 (N_23261,N_15349,N_16799);
nand U23262 (N_23262,N_19113,N_15006);
nor U23263 (N_23263,N_16922,N_19911);
nand U23264 (N_23264,N_16577,N_18679);
or U23265 (N_23265,N_18519,N_15640);
nor U23266 (N_23266,N_16081,N_16463);
xor U23267 (N_23267,N_18668,N_17396);
nand U23268 (N_23268,N_16071,N_19493);
and U23269 (N_23269,N_19320,N_17273);
and U23270 (N_23270,N_17826,N_17036);
nand U23271 (N_23271,N_17080,N_18875);
nand U23272 (N_23272,N_19974,N_15634);
nor U23273 (N_23273,N_19959,N_18509);
nor U23274 (N_23274,N_19945,N_19707);
or U23275 (N_23275,N_19678,N_19350);
and U23276 (N_23276,N_17613,N_18076);
and U23277 (N_23277,N_17745,N_19924);
nor U23278 (N_23278,N_18811,N_16248);
or U23279 (N_23279,N_17177,N_16376);
nand U23280 (N_23280,N_17681,N_15835);
nor U23281 (N_23281,N_16421,N_17605);
xor U23282 (N_23282,N_16702,N_17063);
and U23283 (N_23283,N_19548,N_18435);
and U23284 (N_23284,N_15709,N_19671);
or U23285 (N_23285,N_15125,N_15916);
nor U23286 (N_23286,N_19321,N_15134);
or U23287 (N_23287,N_15657,N_18969);
nand U23288 (N_23288,N_15447,N_17234);
nand U23289 (N_23289,N_16537,N_19050);
nand U23290 (N_23290,N_18126,N_18859);
or U23291 (N_23291,N_16510,N_19441);
or U23292 (N_23292,N_17532,N_18623);
nor U23293 (N_23293,N_19587,N_16406);
or U23294 (N_23294,N_18260,N_18539);
or U23295 (N_23295,N_19763,N_18513);
xnor U23296 (N_23296,N_15508,N_17719);
or U23297 (N_23297,N_19107,N_15254);
and U23298 (N_23298,N_15734,N_18178);
and U23299 (N_23299,N_15352,N_15968);
nand U23300 (N_23300,N_17081,N_16857);
xor U23301 (N_23301,N_15839,N_15302);
and U23302 (N_23302,N_15128,N_16207);
or U23303 (N_23303,N_18943,N_19089);
and U23304 (N_23304,N_18725,N_17348);
nor U23305 (N_23305,N_19727,N_15339);
nand U23306 (N_23306,N_17845,N_17147);
and U23307 (N_23307,N_18681,N_15840);
or U23308 (N_23308,N_15358,N_16413);
and U23309 (N_23309,N_18253,N_17500);
nor U23310 (N_23310,N_15049,N_19413);
and U23311 (N_23311,N_16102,N_17202);
and U23312 (N_23312,N_19384,N_17179);
or U23313 (N_23313,N_15557,N_19528);
and U23314 (N_23314,N_18281,N_15117);
xnor U23315 (N_23315,N_18819,N_15541);
nor U23316 (N_23316,N_19210,N_15123);
or U23317 (N_23317,N_17544,N_16843);
nor U23318 (N_23318,N_19553,N_17724);
and U23319 (N_23319,N_18059,N_19384);
nand U23320 (N_23320,N_18350,N_19826);
nand U23321 (N_23321,N_19019,N_16930);
nor U23322 (N_23322,N_19242,N_17482);
and U23323 (N_23323,N_19372,N_17999);
and U23324 (N_23324,N_19565,N_16026);
and U23325 (N_23325,N_17077,N_19808);
nor U23326 (N_23326,N_17748,N_16256);
xor U23327 (N_23327,N_16847,N_16027);
and U23328 (N_23328,N_16312,N_16339);
or U23329 (N_23329,N_15429,N_15857);
and U23330 (N_23330,N_19798,N_17259);
nor U23331 (N_23331,N_19415,N_17234);
nor U23332 (N_23332,N_16650,N_17122);
xor U23333 (N_23333,N_15642,N_16931);
xor U23334 (N_23334,N_16124,N_18403);
and U23335 (N_23335,N_18529,N_18054);
nand U23336 (N_23336,N_17285,N_17774);
nor U23337 (N_23337,N_16420,N_17885);
or U23338 (N_23338,N_19466,N_18979);
nor U23339 (N_23339,N_17553,N_17176);
nor U23340 (N_23340,N_19994,N_15520);
and U23341 (N_23341,N_15919,N_15555);
or U23342 (N_23342,N_18454,N_15783);
and U23343 (N_23343,N_16769,N_17122);
nor U23344 (N_23344,N_18299,N_15844);
xnor U23345 (N_23345,N_18819,N_19594);
nand U23346 (N_23346,N_17105,N_17979);
nor U23347 (N_23347,N_17447,N_19566);
nand U23348 (N_23348,N_17191,N_15910);
nor U23349 (N_23349,N_18353,N_16068);
nand U23350 (N_23350,N_15412,N_17627);
or U23351 (N_23351,N_19085,N_17054);
or U23352 (N_23352,N_15571,N_15302);
and U23353 (N_23353,N_19174,N_19302);
xnor U23354 (N_23354,N_19334,N_18534);
and U23355 (N_23355,N_19323,N_19382);
or U23356 (N_23356,N_15464,N_18505);
and U23357 (N_23357,N_17203,N_15723);
nand U23358 (N_23358,N_15417,N_19073);
nor U23359 (N_23359,N_16583,N_16506);
xnor U23360 (N_23360,N_17232,N_18909);
nand U23361 (N_23361,N_15405,N_16004);
and U23362 (N_23362,N_16315,N_16419);
and U23363 (N_23363,N_16681,N_16311);
xnor U23364 (N_23364,N_16864,N_19887);
nand U23365 (N_23365,N_18295,N_18933);
nor U23366 (N_23366,N_19552,N_19426);
nor U23367 (N_23367,N_18355,N_18373);
nand U23368 (N_23368,N_19660,N_19002);
nor U23369 (N_23369,N_17097,N_16952);
nor U23370 (N_23370,N_19444,N_15250);
or U23371 (N_23371,N_15750,N_19459);
and U23372 (N_23372,N_17266,N_16470);
or U23373 (N_23373,N_16843,N_17391);
nand U23374 (N_23374,N_17536,N_19695);
or U23375 (N_23375,N_16680,N_16990);
nor U23376 (N_23376,N_16985,N_19179);
nand U23377 (N_23377,N_17691,N_15517);
nand U23378 (N_23378,N_17495,N_17948);
nor U23379 (N_23379,N_15557,N_19898);
xnor U23380 (N_23380,N_15783,N_19660);
nor U23381 (N_23381,N_16392,N_18746);
nand U23382 (N_23382,N_19119,N_18688);
nor U23383 (N_23383,N_18370,N_17301);
and U23384 (N_23384,N_15880,N_17308);
nand U23385 (N_23385,N_17197,N_19012);
or U23386 (N_23386,N_16741,N_15199);
or U23387 (N_23387,N_19075,N_16488);
nand U23388 (N_23388,N_16602,N_16327);
nand U23389 (N_23389,N_15484,N_15001);
or U23390 (N_23390,N_19295,N_17117);
nand U23391 (N_23391,N_15424,N_19876);
nor U23392 (N_23392,N_16156,N_17723);
nand U23393 (N_23393,N_17989,N_16882);
and U23394 (N_23394,N_18315,N_18769);
xor U23395 (N_23395,N_19487,N_16448);
and U23396 (N_23396,N_18615,N_16970);
and U23397 (N_23397,N_19636,N_18250);
and U23398 (N_23398,N_18201,N_17691);
nor U23399 (N_23399,N_16531,N_18788);
or U23400 (N_23400,N_15943,N_15348);
nor U23401 (N_23401,N_16832,N_18971);
nand U23402 (N_23402,N_18755,N_17033);
nand U23403 (N_23403,N_15840,N_18896);
and U23404 (N_23404,N_16806,N_16332);
or U23405 (N_23405,N_17966,N_16100);
and U23406 (N_23406,N_19139,N_17474);
nor U23407 (N_23407,N_19847,N_15033);
xnor U23408 (N_23408,N_16597,N_17345);
xor U23409 (N_23409,N_18825,N_18053);
and U23410 (N_23410,N_16709,N_17003);
nand U23411 (N_23411,N_19421,N_16397);
nand U23412 (N_23412,N_15696,N_19182);
and U23413 (N_23413,N_16764,N_19697);
or U23414 (N_23414,N_19260,N_17489);
or U23415 (N_23415,N_17401,N_15408);
or U23416 (N_23416,N_19504,N_19033);
nand U23417 (N_23417,N_18034,N_17273);
nor U23418 (N_23418,N_19493,N_17838);
nand U23419 (N_23419,N_18759,N_15147);
xor U23420 (N_23420,N_19156,N_16071);
nand U23421 (N_23421,N_18861,N_16006);
xnor U23422 (N_23422,N_17034,N_19453);
nand U23423 (N_23423,N_19548,N_16979);
nand U23424 (N_23424,N_17804,N_19187);
nand U23425 (N_23425,N_16898,N_17832);
and U23426 (N_23426,N_16106,N_19594);
xor U23427 (N_23427,N_15971,N_19480);
nor U23428 (N_23428,N_15466,N_19738);
nor U23429 (N_23429,N_15650,N_18273);
nor U23430 (N_23430,N_17406,N_15777);
or U23431 (N_23431,N_19895,N_18365);
or U23432 (N_23432,N_15788,N_19940);
nand U23433 (N_23433,N_18192,N_16680);
or U23434 (N_23434,N_15005,N_16342);
xor U23435 (N_23435,N_15661,N_16762);
or U23436 (N_23436,N_19990,N_19637);
nor U23437 (N_23437,N_17500,N_17417);
and U23438 (N_23438,N_18492,N_19008);
nand U23439 (N_23439,N_16446,N_18239);
and U23440 (N_23440,N_17734,N_15072);
nor U23441 (N_23441,N_18584,N_16938);
nor U23442 (N_23442,N_19619,N_18268);
or U23443 (N_23443,N_19715,N_16391);
nor U23444 (N_23444,N_17862,N_15683);
or U23445 (N_23445,N_16130,N_19420);
nand U23446 (N_23446,N_19406,N_18942);
nor U23447 (N_23447,N_15970,N_17691);
or U23448 (N_23448,N_17394,N_17728);
nor U23449 (N_23449,N_18360,N_16988);
nand U23450 (N_23450,N_18231,N_17883);
nor U23451 (N_23451,N_17807,N_15255);
nand U23452 (N_23452,N_18269,N_17427);
nor U23453 (N_23453,N_15557,N_16500);
nor U23454 (N_23454,N_18201,N_18990);
nand U23455 (N_23455,N_18642,N_18697);
or U23456 (N_23456,N_19404,N_19648);
nand U23457 (N_23457,N_19032,N_18163);
or U23458 (N_23458,N_18345,N_16923);
and U23459 (N_23459,N_18348,N_19367);
nand U23460 (N_23460,N_16235,N_17403);
or U23461 (N_23461,N_19532,N_19446);
and U23462 (N_23462,N_15086,N_17826);
and U23463 (N_23463,N_19938,N_17270);
nand U23464 (N_23464,N_18778,N_19574);
nor U23465 (N_23465,N_17828,N_18764);
or U23466 (N_23466,N_18079,N_15962);
nand U23467 (N_23467,N_17048,N_17211);
nand U23468 (N_23468,N_19748,N_19699);
or U23469 (N_23469,N_15098,N_16530);
xnor U23470 (N_23470,N_17005,N_18974);
nand U23471 (N_23471,N_16835,N_16494);
nor U23472 (N_23472,N_17641,N_19793);
nand U23473 (N_23473,N_17672,N_19728);
xnor U23474 (N_23474,N_16037,N_17943);
and U23475 (N_23475,N_19258,N_15983);
xor U23476 (N_23476,N_18693,N_15276);
nor U23477 (N_23477,N_17434,N_17855);
and U23478 (N_23478,N_18996,N_18246);
nor U23479 (N_23479,N_18756,N_18604);
xor U23480 (N_23480,N_15483,N_17566);
nand U23481 (N_23481,N_15223,N_15452);
or U23482 (N_23482,N_18223,N_15359);
and U23483 (N_23483,N_19616,N_18778);
nor U23484 (N_23484,N_15232,N_18720);
xnor U23485 (N_23485,N_17583,N_18529);
nor U23486 (N_23486,N_18515,N_17905);
nor U23487 (N_23487,N_19333,N_16893);
nand U23488 (N_23488,N_18591,N_18882);
and U23489 (N_23489,N_15772,N_19598);
and U23490 (N_23490,N_16502,N_19455);
and U23491 (N_23491,N_17364,N_17624);
nand U23492 (N_23492,N_18683,N_17525);
or U23493 (N_23493,N_18544,N_17126);
xnor U23494 (N_23494,N_16069,N_17742);
and U23495 (N_23495,N_17578,N_15278);
or U23496 (N_23496,N_17538,N_17757);
and U23497 (N_23497,N_17219,N_18414);
or U23498 (N_23498,N_17335,N_19414);
nor U23499 (N_23499,N_17413,N_18067);
xnor U23500 (N_23500,N_17754,N_17530);
nor U23501 (N_23501,N_19348,N_17603);
or U23502 (N_23502,N_19504,N_18739);
nor U23503 (N_23503,N_18050,N_17412);
nand U23504 (N_23504,N_19261,N_15260);
and U23505 (N_23505,N_18613,N_17515);
and U23506 (N_23506,N_16515,N_19678);
nand U23507 (N_23507,N_15728,N_17071);
or U23508 (N_23508,N_16380,N_19461);
nand U23509 (N_23509,N_16895,N_18573);
nand U23510 (N_23510,N_18870,N_15283);
nand U23511 (N_23511,N_18572,N_15526);
nor U23512 (N_23512,N_15214,N_17656);
nor U23513 (N_23513,N_18405,N_16896);
xor U23514 (N_23514,N_17398,N_18073);
nor U23515 (N_23515,N_17163,N_19640);
xnor U23516 (N_23516,N_15729,N_16089);
xor U23517 (N_23517,N_18222,N_15286);
nand U23518 (N_23518,N_16614,N_15084);
or U23519 (N_23519,N_15198,N_18765);
nand U23520 (N_23520,N_19072,N_15814);
and U23521 (N_23521,N_16821,N_16116);
nand U23522 (N_23522,N_18420,N_18918);
nor U23523 (N_23523,N_16956,N_15871);
nor U23524 (N_23524,N_19359,N_19859);
and U23525 (N_23525,N_17583,N_19290);
nand U23526 (N_23526,N_17021,N_15094);
nand U23527 (N_23527,N_17150,N_19472);
xnor U23528 (N_23528,N_15963,N_18099);
or U23529 (N_23529,N_16556,N_15735);
nor U23530 (N_23530,N_15034,N_19803);
nand U23531 (N_23531,N_15072,N_19976);
and U23532 (N_23532,N_17583,N_17440);
or U23533 (N_23533,N_17779,N_19281);
nand U23534 (N_23534,N_16736,N_17435);
or U23535 (N_23535,N_19682,N_15754);
nor U23536 (N_23536,N_15867,N_19411);
and U23537 (N_23537,N_18405,N_18488);
nand U23538 (N_23538,N_15100,N_15317);
nor U23539 (N_23539,N_15960,N_19604);
xnor U23540 (N_23540,N_18740,N_18003);
nand U23541 (N_23541,N_17269,N_15863);
or U23542 (N_23542,N_18448,N_15300);
and U23543 (N_23543,N_18135,N_19684);
nor U23544 (N_23544,N_16880,N_16860);
and U23545 (N_23545,N_17905,N_15888);
xnor U23546 (N_23546,N_15322,N_19466);
or U23547 (N_23547,N_18154,N_15763);
and U23548 (N_23548,N_18712,N_18918);
nand U23549 (N_23549,N_17918,N_19729);
xor U23550 (N_23550,N_15540,N_17316);
nand U23551 (N_23551,N_18581,N_17949);
nor U23552 (N_23552,N_18253,N_16170);
or U23553 (N_23553,N_15068,N_17819);
and U23554 (N_23554,N_19653,N_17683);
or U23555 (N_23555,N_19867,N_16978);
and U23556 (N_23556,N_19976,N_17111);
and U23557 (N_23557,N_19953,N_15406);
and U23558 (N_23558,N_15606,N_17698);
and U23559 (N_23559,N_15015,N_19320);
nor U23560 (N_23560,N_17617,N_19659);
xor U23561 (N_23561,N_15598,N_18220);
nor U23562 (N_23562,N_17749,N_19526);
and U23563 (N_23563,N_16606,N_16265);
or U23564 (N_23564,N_16547,N_18942);
nor U23565 (N_23565,N_18129,N_15782);
nor U23566 (N_23566,N_16405,N_17174);
nor U23567 (N_23567,N_18123,N_19567);
nand U23568 (N_23568,N_16758,N_19513);
and U23569 (N_23569,N_19887,N_15566);
and U23570 (N_23570,N_18085,N_15187);
nor U23571 (N_23571,N_19834,N_16522);
xnor U23572 (N_23572,N_18888,N_18565);
or U23573 (N_23573,N_17554,N_19142);
and U23574 (N_23574,N_17398,N_18103);
nor U23575 (N_23575,N_15063,N_15211);
and U23576 (N_23576,N_18939,N_17613);
or U23577 (N_23577,N_18293,N_17782);
and U23578 (N_23578,N_16083,N_17061);
and U23579 (N_23579,N_19197,N_16270);
or U23580 (N_23580,N_19826,N_19324);
nor U23581 (N_23581,N_17325,N_18851);
and U23582 (N_23582,N_15565,N_16376);
and U23583 (N_23583,N_18714,N_15191);
nand U23584 (N_23584,N_18458,N_17558);
and U23585 (N_23585,N_16185,N_17478);
nand U23586 (N_23586,N_17245,N_15465);
and U23587 (N_23587,N_16351,N_19308);
or U23588 (N_23588,N_15489,N_15469);
and U23589 (N_23589,N_17489,N_16448);
xnor U23590 (N_23590,N_17283,N_17367);
nor U23591 (N_23591,N_16555,N_16559);
and U23592 (N_23592,N_17672,N_18030);
or U23593 (N_23593,N_17541,N_18069);
nor U23594 (N_23594,N_15479,N_19635);
and U23595 (N_23595,N_17755,N_17568);
or U23596 (N_23596,N_18003,N_16872);
or U23597 (N_23597,N_17142,N_18948);
nor U23598 (N_23598,N_19606,N_19496);
or U23599 (N_23599,N_18624,N_19477);
nor U23600 (N_23600,N_18825,N_19262);
nor U23601 (N_23601,N_15288,N_16049);
nor U23602 (N_23602,N_19163,N_16738);
and U23603 (N_23603,N_18234,N_18962);
xor U23604 (N_23604,N_16774,N_16459);
or U23605 (N_23605,N_19291,N_17323);
or U23606 (N_23606,N_18590,N_15611);
nor U23607 (N_23607,N_15175,N_16706);
nor U23608 (N_23608,N_16865,N_15187);
nor U23609 (N_23609,N_16213,N_16693);
nor U23610 (N_23610,N_18819,N_15394);
or U23611 (N_23611,N_16128,N_16549);
nand U23612 (N_23612,N_17911,N_17076);
or U23613 (N_23613,N_18639,N_19713);
or U23614 (N_23614,N_16445,N_19659);
and U23615 (N_23615,N_15279,N_16317);
nor U23616 (N_23616,N_19251,N_15400);
and U23617 (N_23617,N_16329,N_15968);
or U23618 (N_23618,N_17824,N_15904);
or U23619 (N_23619,N_18759,N_16178);
nor U23620 (N_23620,N_19161,N_16267);
nand U23621 (N_23621,N_16199,N_19255);
nand U23622 (N_23622,N_18823,N_19171);
nand U23623 (N_23623,N_15046,N_18529);
xnor U23624 (N_23624,N_15532,N_17893);
nor U23625 (N_23625,N_17263,N_17318);
xor U23626 (N_23626,N_19258,N_17970);
or U23627 (N_23627,N_17829,N_17988);
and U23628 (N_23628,N_18934,N_17568);
and U23629 (N_23629,N_17296,N_15457);
nand U23630 (N_23630,N_16890,N_17309);
and U23631 (N_23631,N_15492,N_19307);
or U23632 (N_23632,N_16857,N_17597);
nor U23633 (N_23633,N_18820,N_17227);
nor U23634 (N_23634,N_18869,N_18630);
and U23635 (N_23635,N_16785,N_18038);
nand U23636 (N_23636,N_17428,N_19304);
nand U23637 (N_23637,N_19953,N_16401);
nand U23638 (N_23638,N_19005,N_19659);
nand U23639 (N_23639,N_16222,N_16249);
nor U23640 (N_23640,N_17717,N_18648);
xor U23641 (N_23641,N_18395,N_19593);
nand U23642 (N_23642,N_17794,N_19560);
or U23643 (N_23643,N_18694,N_16427);
or U23644 (N_23644,N_18959,N_19170);
or U23645 (N_23645,N_17167,N_18706);
nor U23646 (N_23646,N_18410,N_17035);
nor U23647 (N_23647,N_18986,N_19151);
and U23648 (N_23648,N_15463,N_18556);
and U23649 (N_23649,N_16705,N_17680);
and U23650 (N_23650,N_19802,N_15431);
and U23651 (N_23651,N_16159,N_16337);
or U23652 (N_23652,N_15133,N_17971);
xor U23653 (N_23653,N_17224,N_17120);
or U23654 (N_23654,N_17765,N_18651);
nand U23655 (N_23655,N_15407,N_17100);
nor U23656 (N_23656,N_18843,N_16373);
nor U23657 (N_23657,N_16726,N_17359);
nor U23658 (N_23658,N_18822,N_17791);
or U23659 (N_23659,N_15097,N_17448);
and U23660 (N_23660,N_15695,N_16322);
and U23661 (N_23661,N_15105,N_19862);
or U23662 (N_23662,N_17589,N_17593);
and U23663 (N_23663,N_18704,N_16688);
nand U23664 (N_23664,N_15448,N_15013);
or U23665 (N_23665,N_16227,N_19680);
nor U23666 (N_23666,N_15449,N_15096);
or U23667 (N_23667,N_18333,N_15230);
or U23668 (N_23668,N_18841,N_15153);
or U23669 (N_23669,N_18945,N_19031);
and U23670 (N_23670,N_15292,N_15737);
nor U23671 (N_23671,N_19819,N_19473);
or U23672 (N_23672,N_17426,N_18112);
and U23673 (N_23673,N_19551,N_15440);
nand U23674 (N_23674,N_16299,N_19521);
or U23675 (N_23675,N_17217,N_15489);
and U23676 (N_23676,N_16878,N_17147);
nor U23677 (N_23677,N_15972,N_15281);
xor U23678 (N_23678,N_15193,N_16535);
nand U23679 (N_23679,N_18131,N_18361);
nor U23680 (N_23680,N_19078,N_19587);
and U23681 (N_23681,N_19909,N_17111);
xnor U23682 (N_23682,N_16475,N_19814);
and U23683 (N_23683,N_18001,N_15413);
xnor U23684 (N_23684,N_18944,N_18964);
or U23685 (N_23685,N_15986,N_19980);
nor U23686 (N_23686,N_15946,N_17273);
nor U23687 (N_23687,N_18250,N_19477);
and U23688 (N_23688,N_18632,N_16647);
and U23689 (N_23689,N_18596,N_17075);
nor U23690 (N_23690,N_15971,N_18129);
or U23691 (N_23691,N_18834,N_17931);
and U23692 (N_23692,N_15717,N_19977);
or U23693 (N_23693,N_16598,N_16278);
nor U23694 (N_23694,N_15449,N_16101);
or U23695 (N_23695,N_17662,N_19666);
and U23696 (N_23696,N_19492,N_19332);
nand U23697 (N_23697,N_15770,N_16487);
and U23698 (N_23698,N_15786,N_19150);
nand U23699 (N_23699,N_19961,N_17061);
or U23700 (N_23700,N_15417,N_19208);
nor U23701 (N_23701,N_15137,N_19360);
and U23702 (N_23702,N_15777,N_17950);
xor U23703 (N_23703,N_15265,N_19634);
nand U23704 (N_23704,N_15957,N_19784);
or U23705 (N_23705,N_15150,N_15689);
xor U23706 (N_23706,N_15675,N_15290);
and U23707 (N_23707,N_16734,N_19247);
or U23708 (N_23708,N_15739,N_17572);
nand U23709 (N_23709,N_15689,N_17268);
or U23710 (N_23710,N_15038,N_19741);
or U23711 (N_23711,N_17877,N_19541);
and U23712 (N_23712,N_19585,N_17560);
or U23713 (N_23713,N_16718,N_16618);
or U23714 (N_23714,N_15110,N_19306);
nor U23715 (N_23715,N_17090,N_19860);
nand U23716 (N_23716,N_19141,N_15163);
and U23717 (N_23717,N_15110,N_19625);
nor U23718 (N_23718,N_19607,N_16553);
nor U23719 (N_23719,N_19273,N_16574);
xnor U23720 (N_23720,N_18236,N_19246);
or U23721 (N_23721,N_17639,N_16046);
and U23722 (N_23722,N_19823,N_19856);
xor U23723 (N_23723,N_18755,N_16771);
or U23724 (N_23724,N_19978,N_17810);
nand U23725 (N_23725,N_19767,N_17625);
nor U23726 (N_23726,N_15414,N_19698);
nand U23727 (N_23727,N_19585,N_18283);
and U23728 (N_23728,N_19017,N_16178);
and U23729 (N_23729,N_17045,N_18073);
or U23730 (N_23730,N_17400,N_15308);
nand U23731 (N_23731,N_17924,N_16649);
and U23732 (N_23732,N_19922,N_15331);
and U23733 (N_23733,N_18391,N_17138);
nor U23734 (N_23734,N_18733,N_19550);
nor U23735 (N_23735,N_19030,N_17225);
or U23736 (N_23736,N_15970,N_16819);
nor U23737 (N_23737,N_19110,N_17040);
and U23738 (N_23738,N_17102,N_18966);
xor U23739 (N_23739,N_15740,N_19673);
nor U23740 (N_23740,N_15158,N_16525);
and U23741 (N_23741,N_16754,N_18714);
nor U23742 (N_23742,N_17292,N_15764);
xnor U23743 (N_23743,N_17286,N_19003);
xor U23744 (N_23744,N_15994,N_18446);
and U23745 (N_23745,N_18549,N_17939);
nand U23746 (N_23746,N_16371,N_15268);
and U23747 (N_23747,N_18440,N_19867);
nand U23748 (N_23748,N_18082,N_15578);
nor U23749 (N_23749,N_16351,N_15465);
nor U23750 (N_23750,N_15857,N_15256);
nand U23751 (N_23751,N_17475,N_18330);
nand U23752 (N_23752,N_17152,N_15077);
or U23753 (N_23753,N_15813,N_15080);
nor U23754 (N_23754,N_18144,N_18820);
and U23755 (N_23755,N_15154,N_16760);
nand U23756 (N_23756,N_18521,N_18420);
and U23757 (N_23757,N_16278,N_18718);
and U23758 (N_23758,N_17794,N_16693);
and U23759 (N_23759,N_16593,N_17206);
nand U23760 (N_23760,N_16848,N_17318);
nor U23761 (N_23761,N_15554,N_19393);
or U23762 (N_23762,N_18640,N_18019);
nor U23763 (N_23763,N_15750,N_15831);
or U23764 (N_23764,N_18024,N_19633);
xnor U23765 (N_23765,N_17400,N_16136);
or U23766 (N_23766,N_15050,N_19186);
nand U23767 (N_23767,N_17981,N_15288);
nor U23768 (N_23768,N_16827,N_16402);
nand U23769 (N_23769,N_19419,N_18371);
and U23770 (N_23770,N_18995,N_17544);
nor U23771 (N_23771,N_18640,N_17368);
and U23772 (N_23772,N_15630,N_17576);
nor U23773 (N_23773,N_15124,N_18165);
nor U23774 (N_23774,N_17685,N_19990);
xor U23775 (N_23775,N_17647,N_15079);
xnor U23776 (N_23776,N_18997,N_16739);
nand U23777 (N_23777,N_16031,N_15506);
xor U23778 (N_23778,N_16961,N_17185);
and U23779 (N_23779,N_19133,N_17018);
nor U23780 (N_23780,N_18263,N_16232);
nor U23781 (N_23781,N_18130,N_19085);
nand U23782 (N_23782,N_19558,N_17778);
nand U23783 (N_23783,N_15623,N_15108);
xor U23784 (N_23784,N_15688,N_17172);
nor U23785 (N_23785,N_19272,N_18314);
nor U23786 (N_23786,N_17314,N_18248);
nand U23787 (N_23787,N_18389,N_19440);
and U23788 (N_23788,N_17845,N_15855);
nor U23789 (N_23789,N_19401,N_17763);
xnor U23790 (N_23790,N_17080,N_17530);
xnor U23791 (N_23791,N_18464,N_15431);
xnor U23792 (N_23792,N_15367,N_18473);
nor U23793 (N_23793,N_17239,N_15458);
nand U23794 (N_23794,N_16008,N_18700);
or U23795 (N_23795,N_19095,N_18701);
nor U23796 (N_23796,N_17676,N_17191);
nor U23797 (N_23797,N_15802,N_19314);
xor U23798 (N_23798,N_18013,N_18399);
and U23799 (N_23799,N_17779,N_15149);
nor U23800 (N_23800,N_15212,N_18731);
or U23801 (N_23801,N_19736,N_19213);
nand U23802 (N_23802,N_18075,N_17172);
nor U23803 (N_23803,N_15064,N_19989);
or U23804 (N_23804,N_17048,N_15336);
nor U23805 (N_23805,N_16108,N_19611);
nand U23806 (N_23806,N_17399,N_17272);
nand U23807 (N_23807,N_15062,N_18884);
nand U23808 (N_23808,N_18938,N_15847);
nor U23809 (N_23809,N_19502,N_19133);
xnor U23810 (N_23810,N_16858,N_18436);
xnor U23811 (N_23811,N_19632,N_15174);
nor U23812 (N_23812,N_19999,N_17862);
and U23813 (N_23813,N_18992,N_15747);
xor U23814 (N_23814,N_19153,N_16565);
nand U23815 (N_23815,N_15697,N_19183);
xor U23816 (N_23816,N_19485,N_18047);
or U23817 (N_23817,N_17196,N_19032);
nor U23818 (N_23818,N_16040,N_15098);
and U23819 (N_23819,N_18552,N_17518);
nand U23820 (N_23820,N_17417,N_18501);
xnor U23821 (N_23821,N_18660,N_15215);
or U23822 (N_23822,N_19719,N_16008);
nor U23823 (N_23823,N_16951,N_19389);
nor U23824 (N_23824,N_18312,N_19909);
and U23825 (N_23825,N_17186,N_18954);
nor U23826 (N_23826,N_19376,N_18717);
or U23827 (N_23827,N_15649,N_15988);
nor U23828 (N_23828,N_17356,N_17868);
nand U23829 (N_23829,N_15839,N_16601);
nor U23830 (N_23830,N_16574,N_19660);
xor U23831 (N_23831,N_16488,N_17369);
or U23832 (N_23832,N_18983,N_17551);
or U23833 (N_23833,N_18254,N_16498);
nor U23834 (N_23834,N_15972,N_17793);
and U23835 (N_23835,N_17421,N_19959);
nand U23836 (N_23836,N_17748,N_15764);
nor U23837 (N_23837,N_19421,N_18479);
or U23838 (N_23838,N_15406,N_15216);
nand U23839 (N_23839,N_16320,N_15105);
or U23840 (N_23840,N_19718,N_19807);
nor U23841 (N_23841,N_16307,N_17313);
nand U23842 (N_23842,N_16977,N_18183);
nand U23843 (N_23843,N_19425,N_17691);
and U23844 (N_23844,N_17649,N_18724);
nand U23845 (N_23845,N_15387,N_18139);
xnor U23846 (N_23846,N_16103,N_16343);
nand U23847 (N_23847,N_17788,N_16059);
nand U23848 (N_23848,N_19368,N_18195);
nor U23849 (N_23849,N_16241,N_18301);
and U23850 (N_23850,N_18158,N_19397);
nor U23851 (N_23851,N_18588,N_18794);
and U23852 (N_23852,N_15057,N_18342);
nand U23853 (N_23853,N_17884,N_18422);
and U23854 (N_23854,N_17472,N_15161);
or U23855 (N_23855,N_17601,N_16054);
and U23856 (N_23856,N_17759,N_15361);
nor U23857 (N_23857,N_15790,N_15745);
and U23858 (N_23858,N_18210,N_18390);
nand U23859 (N_23859,N_19730,N_17770);
nand U23860 (N_23860,N_15136,N_16084);
or U23861 (N_23861,N_17031,N_16362);
or U23862 (N_23862,N_18223,N_18703);
or U23863 (N_23863,N_16591,N_15686);
and U23864 (N_23864,N_15779,N_18650);
or U23865 (N_23865,N_17192,N_16844);
nand U23866 (N_23866,N_18871,N_17777);
and U23867 (N_23867,N_16034,N_17350);
or U23868 (N_23868,N_18488,N_19280);
and U23869 (N_23869,N_16112,N_15989);
and U23870 (N_23870,N_18247,N_15542);
nand U23871 (N_23871,N_17955,N_17372);
nand U23872 (N_23872,N_15454,N_17725);
nand U23873 (N_23873,N_19985,N_15507);
nand U23874 (N_23874,N_19899,N_15518);
xnor U23875 (N_23875,N_17654,N_15616);
or U23876 (N_23876,N_19383,N_19537);
nand U23877 (N_23877,N_19354,N_17755);
nor U23878 (N_23878,N_17988,N_16521);
xor U23879 (N_23879,N_18611,N_15380);
xor U23880 (N_23880,N_18899,N_17377);
or U23881 (N_23881,N_17828,N_17729);
nand U23882 (N_23882,N_18578,N_18684);
nand U23883 (N_23883,N_16443,N_17530);
and U23884 (N_23884,N_15787,N_16092);
and U23885 (N_23885,N_17026,N_16044);
and U23886 (N_23886,N_18798,N_15434);
nand U23887 (N_23887,N_18751,N_19882);
nor U23888 (N_23888,N_15310,N_19106);
or U23889 (N_23889,N_15014,N_16486);
and U23890 (N_23890,N_15919,N_18947);
and U23891 (N_23891,N_18783,N_19789);
or U23892 (N_23892,N_15038,N_17821);
xnor U23893 (N_23893,N_18064,N_17315);
nor U23894 (N_23894,N_18169,N_17114);
or U23895 (N_23895,N_16708,N_17857);
and U23896 (N_23896,N_15599,N_17646);
and U23897 (N_23897,N_19386,N_19940);
xnor U23898 (N_23898,N_19187,N_18438);
nand U23899 (N_23899,N_16614,N_19986);
or U23900 (N_23900,N_17378,N_19850);
nand U23901 (N_23901,N_19585,N_19374);
nor U23902 (N_23902,N_18830,N_16073);
nor U23903 (N_23903,N_15258,N_19982);
nor U23904 (N_23904,N_18894,N_16274);
nor U23905 (N_23905,N_16143,N_15492);
nor U23906 (N_23906,N_15769,N_17997);
nand U23907 (N_23907,N_19469,N_15657);
nor U23908 (N_23908,N_15959,N_15875);
nor U23909 (N_23909,N_18532,N_15856);
or U23910 (N_23910,N_16333,N_19358);
nor U23911 (N_23911,N_16823,N_18797);
and U23912 (N_23912,N_16375,N_17045);
or U23913 (N_23913,N_18192,N_17291);
or U23914 (N_23914,N_15663,N_15844);
nor U23915 (N_23915,N_19826,N_17312);
nand U23916 (N_23916,N_16051,N_17076);
nand U23917 (N_23917,N_19741,N_18858);
and U23918 (N_23918,N_17707,N_19366);
nor U23919 (N_23919,N_19943,N_18744);
or U23920 (N_23920,N_15191,N_15628);
and U23921 (N_23921,N_19848,N_16606);
and U23922 (N_23922,N_15683,N_15938);
and U23923 (N_23923,N_19090,N_19079);
nor U23924 (N_23924,N_17370,N_15654);
xor U23925 (N_23925,N_17367,N_15342);
or U23926 (N_23926,N_19470,N_18493);
nor U23927 (N_23927,N_19158,N_16011);
xor U23928 (N_23928,N_18067,N_17088);
or U23929 (N_23929,N_16106,N_17954);
nand U23930 (N_23930,N_15698,N_17156);
and U23931 (N_23931,N_19101,N_16735);
xor U23932 (N_23932,N_18372,N_18108);
nor U23933 (N_23933,N_17025,N_15106);
nand U23934 (N_23934,N_16757,N_16724);
nand U23935 (N_23935,N_17243,N_19747);
or U23936 (N_23936,N_19736,N_17490);
nor U23937 (N_23937,N_15604,N_15841);
and U23938 (N_23938,N_18521,N_17192);
or U23939 (N_23939,N_15621,N_18706);
nor U23940 (N_23940,N_16447,N_18602);
or U23941 (N_23941,N_18442,N_15428);
or U23942 (N_23942,N_17082,N_16417);
and U23943 (N_23943,N_17977,N_16753);
or U23944 (N_23944,N_15686,N_18681);
nand U23945 (N_23945,N_17809,N_16147);
nor U23946 (N_23946,N_19448,N_16951);
nand U23947 (N_23947,N_18247,N_19210);
xor U23948 (N_23948,N_19147,N_18355);
and U23949 (N_23949,N_19307,N_16355);
and U23950 (N_23950,N_19139,N_19840);
nand U23951 (N_23951,N_18055,N_18526);
or U23952 (N_23952,N_15009,N_16139);
or U23953 (N_23953,N_16135,N_19558);
nand U23954 (N_23954,N_15878,N_15002);
or U23955 (N_23955,N_17806,N_19472);
nor U23956 (N_23956,N_15015,N_17436);
nor U23957 (N_23957,N_18666,N_19863);
nor U23958 (N_23958,N_16451,N_18372);
nand U23959 (N_23959,N_16188,N_19011);
and U23960 (N_23960,N_19282,N_16213);
nor U23961 (N_23961,N_18685,N_15723);
nor U23962 (N_23962,N_18694,N_15773);
and U23963 (N_23963,N_19112,N_19588);
or U23964 (N_23964,N_19577,N_18732);
and U23965 (N_23965,N_18900,N_19204);
nand U23966 (N_23966,N_15179,N_16159);
and U23967 (N_23967,N_18273,N_16171);
or U23968 (N_23968,N_16811,N_15180);
nor U23969 (N_23969,N_18596,N_18376);
nor U23970 (N_23970,N_15763,N_16473);
nor U23971 (N_23971,N_19842,N_18449);
nand U23972 (N_23972,N_17045,N_16790);
nor U23973 (N_23973,N_17956,N_16006);
xor U23974 (N_23974,N_15550,N_18908);
xnor U23975 (N_23975,N_17815,N_19190);
nand U23976 (N_23976,N_15447,N_15022);
nand U23977 (N_23977,N_19551,N_16756);
and U23978 (N_23978,N_15476,N_15336);
nor U23979 (N_23979,N_16492,N_19820);
or U23980 (N_23980,N_15824,N_15471);
nor U23981 (N_23981,N_16609,N_17377);
or U23982 (N_23982,N_16675,N_19297);
nor U23983 (N_23983,N_15780,N_19772);
or U23984 (N_23984,N_15583,N_16707);
nor U23985 (N_23985,N_18668,N_19189);
nand U23986 (N_23986,N_18887,N_19491);
nor U23987 (N_23987,N_18322,N_19052);
nand U23988 (N_23988,N_19067,N_15513);
nor U23989 (N_23989,N_16048,N_17672);
or U23990 (N_23990,N_18256,N_19306);
nor U23991 (N_23991,N_15156,N_18711);
or U23992 (N_23992,N_15194,N_16212);
nand U23993 (N_23993,N_17777,N_17305);
nand U23994 (N_23994,N_15872,N_17516);
nand U23995 (N_23995,N_17125,N_19130);
nand U23996 (N_23996,N_15208,N_15216);
or U23997 (N_23997,N_18119,N_15029);
nor U23998 (N_23998,N_19360,N_15269);
or U23999 (N_23999,N_17598,N_19447);
nand U24000 (N_24000,N_17349,N_16503);
nand U24001 (N_24001,N_19857,N_17849);
nand U24002 (N_24002,N_18902,N_18601);
nand U24003 (N_24003,N_19367,N_16369);
nor U24004 (N_24004,N_16035,N_16238);
xor U24005 (N_24005,N_15474,N_15390);
and U24006 (N_24006,N_15078,N_15382);
nor U24007 (N_24007,N_15634,N_17013);
and U24008 (N_24008,N_16719,N_17726);
nor U24009 (N_24009,N_16380,N_18388);
xor U24010 (N_24010,N_15635,N_15103);
and U24011 (N_24011,N_16933,N_15430);
or U24012 (N_24012,N_16805,N_15320);
or U24013 (N_24013,N_16105,N_19555);
and U24014 (N_24014,N_17288,N_16393);
nand U24015 (N_24015,N_19575,N_15158);
nand U24016 (N_24016,N_18666,N_19627);
nand U24017 (N_24017,N_18430,N_19875);
nor U24018 (N_24018,N_18875,N_16094);
and U24019 (N_24019,N_15241,N_15539);
or U24020 (N_24020,N_19510,N_17730);
and U24021 (N_24021,N_15891,N_17414);
or U24022 (N_24022,N_18792,N_15148);
or U24023 (N_24023,N_17586,N_17608);
and U24024 (N_24024,N_15661,N_19507);
nand U24025 (N_24025,N_16600,N_18081);
nand U24026 (N_24026,N_15912,N_18497);
or U24027 (N_24027,N_16310,N_16300);
or U24028 (N_24028,N_17436,N_17000);
nor U24029 (N_24029,N_15126,N_16823);
nor U24030 (N_24030,N_18234,N_17650);
or U24031 (N_24031,N_17642,N_19731);
or U24032 (N_24032,N_19957,N_18065);
xnor U24033 (N_24033,N_18478,N_18363);
nand U24034 (N_24034,N_16162,N_18814);
or U24035 (N_24035,N_17816,N_16875);
nor U24036 (N_24036,N_16327,N_19335);
nand U24037 (N_24037,N_19459,N_19769);
nand U24038 (N_24038,N_18177,N_16762);
and U24039 (N_24039,N_15560,N_19853);
nand U24040 (N_24040,N_15438,N_19176);
nor U24041 (N_24041,N_17770,N_17458);
nand U24042 (N_24042,N_16477,N_15158);
nor U24043 (N_24043,N_18784,N_18599);
xnor U24044 (N_24044,N_19772,N_17874);
and U24045 (N_24045,N_16074,N_15102);
nor U24046 (N_24046,N_15451,N_19551);
nand U24047 (N_24047,N_18234,N_15973);
or U24048 (N_24048,N_19031,N_16074);
and U24049 (N_24049,N_17247,N_17413);
nor U24050 (N_24050,N_16369,N_18461);
nor U24051 (N_24051,N_15574,N_17074);
or U24052 (N_24052,N_16960,N_15821);
or U24053 (N_24053,N_19931,N_18386);
and U24054 (N_24054,N_15617,N_19406);
nor U24055 (N_24055,N_17065,N_19753);
or U24056 (N_24056,N_19580,N_16225);
or U24057 (N_24057,N_19141,N_19194);
nand U24058 (N_24058,N_17588,N_19196);
nand U24059 (N_24059,N_16855,N_15775);
and U24060 (N_24060,N_15967,N_17564);
and U24061 (N_24061,N_15064,N_18434);
nor U24062 (N_24062,N_16664,N_15191);
and U24063 (N_24063,N_19171,N_17157);
or U24064 (N_24064,N_18214,N_19741);
nor U24065 (N_24065,N_17171,N_15285);
or U24066 (N_24066,N_17346,N_19120);
or U24067 (N_24067,N_17543,N_17640);
nand U24068 (N_24068,N_15138,N_19127);
or U24069 (N_24069,N_18349,N_17861);
or U24070 (N_24070,N_17339,N_15869);
nor U24071 (N_24071,N_15381,N_15805);
and U24072 (N_24072,N_15170,N_16826);
and U24073 (N_24073,N_19181,N_19672);
nand U24074 (N_24074,N_15353,N_15426);
or U24075 (N_24075,N_19396,N_19309);
nand U24076 (N_24076,N_15324,N_16611);
or U24077 (N_24077,N_17094,N_17384);
nor U24078 (N_24078,N_16077,N_18785);
or U24079 (N_24079,N_15895,N_16003);
nand U24080 (N_24080,N_19121,N_17670);
nand U24081 (N_24081,N_17516,N_18221);
and U24082 (N_24082,N_19204,N_16938);
and U24083 (N_24083,N_15761,N_17746);
and U24084 (N_24084,N_15580,N_17722);
or U24085 (N_24085,N_16563,N_19020);
or U24086 (N_24086,N_16187,N_16064);
or U24087 (N_24087,N_17649,N_17605);
or U24088 (N_24088,N_16374,N_17468);
and U24089 (N_24089,N_17381,N_17358);
and U24090 (N_24090,N_19508,N_16174);
and U24091 (N_24091,N_15644,N_16252);
or U24092 (N_24092,N_19237,N_15925);
and U24093 (N_24093,N_15825,N_16109);
nor U24094 (N_24094,N_16893,N_18882);
xnor U24095 (N_24095,N_18661,N_19709);
or U24096 (N_24096,N_18201,N_15665);
xnor U24097 (N_24097,N_18642,N_19874);
or U24098 (N_24098,N_18546,N_15237);
nor U24099 (N_24099,N_18103,N_18225);
nor U24100 (N_24100,N_16175,N_18840);
nor U24101 (N_24101,N_15097,N_17570);
and U24102 (N_24102,N_16858,N_18449);
nor U24103 (N_24103,N_15964,N_16904);
and U24104 (N_24104,N_15417,N_19594);
or U24105 (N_24105,N_15133,N_17796);
or U24106 (N_24106,N_15040,N_18536);
nand U24107 (N_24107,N_17950,N_16827);
nor U24108 (N_24108,N_19609,N_16734);
nor U24109 (N_24109,N_18495,N_18553);
or U24110 (N_24110,N_17606,N_19025);
and U24111 (N_24111,N_18732,N_16483);
and U24112 (N_24112,N_15592,N_15143);
nand U24113 (N_24113,N_19058,N_18891);
and U24114 (N_24114,N_15700,N_17325);
xor U24115 (N_24115,N_15693,N_17939);
nand U24116 (N_24116,N_19846,N_15983);
nand U24117 (N_24117,N_16764,N_16845);
nor U24118 (N_24118,N_19453,N_15939);
and U24119 (N_24119,N_16288,N_16496);
and U24120 (N_24120,N_17783,N_18593);
nor U24121 (N_24121,N_15392,N_15540);
and U24122 (N_24122,N_19546,N_18212);
nor U24123 (N_24123,N_16919,N_18812);
nand U24124 (N_24124,N_15718,N_15367);
nor U24125 (N_24125,N_19595,N_19387);
nand U24126 (N_24126,N_18342,N_15382);
or U24127 (N_24127,N_17639,N_17429);
and U24128 (N_24128,N_17836,N_19131);
nor U24129 (N_24129,N_17862,N_17552);
nor U24130 (N_24130,N_18063,N_19428);
nor U24131 (N_24131,N_19224,N_18263);
xor U24132 (N_24132,N_15128,N_17669);
nand U24133 (N_24133,N_19665,N_17240);
nand U24134 (N_24134,N_16440,N_17912);
nand U24135 (N_24135,N_18967,N_16920);
and U24136 (N_24136,N_15800,N_17507);
nor U24137 (N_24137,N_17288,N_19548);
nor U24138 (N_24138,N_18893,N_19541);
or U24139 (N_24139,N_19822,N_15606);
nor U24140 (N_24140,N_16247,N_19692);
nor U24141 (N_24141,N_18898,N_16461);
nor U24142 (N_24142,N_18250,N_18377);
nor U24143 (N_24143,N_19631,N_19166);
nand U24144 (N_24144,N_17474,N_16066);
nand U24145 (N_24145,N_19410,N_19794);
and U24146 (N_24146,N_17187,N_19163);
or U24147 (N_24147,N_15751,N_16054);
and U24148 (N_24148,N_15666,N_15487);
or U24149 (N_24149,N_19132,N_17511);
or U24150 (N_24150,N_19110,N_15225);
and U24151 (N_24151,N_15857,N_19693);
nand U24152 (N_24152,N_17820,N_18608);
and U24153 (N_24153,N_15857,N_15968);
nand U24154 (N_24154,N_17566,N_17577);
nand U24155 (N_24155,N_19847,N_16184);
nor U24156 (N_24156,N_18107,N_17327);
nor U24157 (N_24157,N_17815,N_19078);
xor U24158 (N_24158,N_17982,N_15148);
and U24159 (N_24159,N_17849,N_19211);
nand U24160 (N_24160,N_18117,N_19863);
xor U24161 (N_24161,N_17153,N_18587);
or U24162 (N_24162,N_17326,N_19713);
nand U24163 (N_24163,N_19413,N_18396);
and U24164 (N_24164,N_17581,N_18953);
or U24165 (N_24165,N_19260,N_15293);
nand U24166 (N_24166,N_19834,N_15480);
nand U24167 (N_24167,N_19671,N_17403);
nor U24168 (N_24168,N_15885,N_18084);
nand U24169 (N_24169,N_16187,N_17477);
xnor U24170 (N_24170,N_15824,N_17032);
nor U24171 (N_24171,N_17874,N_17596);
nand U24172 (N_24172,N_17357,N_17873);
nand U24173 (N_24173,N_16716,N_16143);
nand U24174 (N_24174,N_17303,N_17432);
nand U24175 (N_24175,N_17745,N_17108);
or U24176 (N_24176,N_15588,N_15691);
and U24177 (N_24177,N_18700,N_19386);
nor U24178 (N_24178,N_16202,N_19072);
or U24179 (N_24179,N_16853,N_16538);
xor U24180 (N_24180,N_16315,N_19746);
and U24181 (N_24181,N_18369,N_16045);
xor U24182 (N_24182,N_16081,N_15335);
nor U24183 (N_24183,N_18527,N_16447);
nand U24184 (N_24184,N_15260,N_17693);
or U24185 (N_24185,N_19272,N_17853);
and U24186 (N_24186,N_15457,N_17978);
and U24187 (N_24187,N_17147,N_17188);
or U24188 (N_24188,N_15204,N_16698);
or U24189 (N_24189,N_16605,N_17603);
nand U24190 (N_24190,N_19017,N_17693);
or U24191 (N_24191,N_15341,N_19925);
and U24192 (N_24192,N_18121,N_16902);
nand U24193 (N_24193,N_15275,N_18876);
and U24194 (N_24194,N_19273,N_16148);
or U24195 (N_24195,N_15618,N_15067);
nor U24196 (N_24196,N_17928,N_15638);
or U24197 (N_24197,N_19774,N_17492);
and U24198 (N_24198,N_18569,N_17802);
nor U24199 (N_24199,N_18253,N_16958);
nor U24200 (N_24200,N_18650,N_18130);
nor U24201 (N_24201,N_17837,N_15787);
nand U24202 (N_24202,N_15224,N_17243);
or U24203 (N_24203,N_19771,N_16218);
or U24204 (N_24204,N_15891,N_19565);
or U24205 (N_24205,N_17368,N_15164);
and U24206 (N_24206,N_17550,N_19566);
nor U24207 (N_24207,N_16819,N_15611);
or U24208 (N_24208,N_15473,N_19084);
nand U24209 (N_24209,N_17414,N_18392);
and U24210 (N_24210,N_17448,N_16682);
nor U24211 (N_24211,N_16086,N_16829);
and U24212 (N_24212,N_18853,N_15936);
nand U24213 (N_24213,N_19901,N_15066);
nor U24214 (N_24214,N_15524,N_19811);
nor U24215 (N_24215,N_15093,N_15930);
and U24216 (N_24216,N_18724,N_18997);
or U24217 (N_24217,N_19388,N_17453);
or U24218 (N_24218,N_15214,N_17964);
and U24219 (N_24219,N_15776,N_15347);
nand U24220 (N_24220,N_16676,N_16475);
or U24221 (N_24221,N_18680,N_17357);
nand U24222 (N_24222,N_15036,N_18105);
xor U24223 (N_24223,N_16103,N_15481);
nand U24224 (N_24224,N_16414,N_15817);
and U24225 (N_24225,N_19939,N_17137);
or U24226 (N_24226,N_15351,N_18746);
nand U24227 (N_24227,N_16520,N_18438);
and U24228 (N_24228,N_19425,N_18087);
or U24229 (N_24229,N_18427,N_17316);
xor U24230 (N_24230,N_18507,N_18439);
nand U24231 (N_24231,N_17487,N_19385);
nor U24232 (N_24232,N_19599,N_16592);
nor U24233 (N_24233,N_16134,N_15997);
nor U24234 (N_24234,N_17113,N_15286);
or U24235 (N_24235,N_17080,N_18061);
and U24236 (N_24236,N_18129,N_17946);
nand U24237 (N_24237,N_18671,N_15958);
nor U24238 (N_24238,N_19753,N_16817);
or U24239 (N_24239,N_15729,N_19298);
nor U24240 (N_24240,N_15660,N_15961);
or U24241 (N_24241,N_16576,N_15858);
or U24242 (N_24242,N_18885,N_15582);
and U24243 (N_24243,N_19060,N_19493);
nor U24244 (N_24244,N_15567,N_15678);
nand U24245 (N_24245,N_17973,N_15738);
nand U24246 (N_24246,N_17648,N_17468);
xnor U24247 (N_24247,N_17174,N_18445);
nor U24248 (N_24248,N_19866,N_18599);
and U24249 (N_24249,N_16892,N_18227);
or U24250 (N_24250,N_16468,N_16836);
and U24251 (N_24251,N_17956,N_16344);
nor U24252 (N_24252,N_15219,N_19981);
and U24253 (N_24253,N_16129,N_18005);
or U24254 (N_24254,N_18676,N_16551);
and U24255 (N_24255,N_15797,N_17577);
nor U24256 (N_24256,N_16897,N_19321);
nand U24257 (N_24257,N_18283,N_16091);
xor U24258 (N_24258,N_17316,N_16399);
or U24259 (N_24259,N_16238,N_17738);
nor U24260 (N_24260,N_17154,N_17974);
or U24261 (N_24261,N_19346,N_17803);
nor U24262 (N_24262,N_18393,N_16630);
xnor U24263 (N_24263,N_19831,N_17248);
nand U24264 (N_24264,N_19943,N_17825);
and U24265 (N_24265,N_15818,N_15060);
nor U24266 (N_24266,N_15278,N_19643);
and U24267 (N_24267,N_18623,N_18308);
nor U24268 (N_24268,N_17573,N_18610);
nor U24269 (N_24269,N_18527,N_16869);
nor U24270 (N_24270,N_19811,N_18969);
nand U24271 (N_24271,N_18912,N_15804);
or U24272 (N_24272,N_16001,N_17643);
nand U24273 (N_24273,N_19201,N_19924);
or U24274 (N_24274,N_18696,N_15776);
and U24275 (N_24275,N_17102,N_19148);
and U24276 (N_24276,N_15748,N_19969);
and U24277 (N_24277,N_17899,N_15713);
and U24278 (N_24278,N_19010,N_15747);
xnor U24279 (N_24279,N_16617,N_16109);
nand U24280 (N_24280,N_15083,N_16621);
or U24281 (N_24281,N_18920,N_19231);
nor U24282 (N_24282,N_16253,N_19850);
or U24283 (N_24283,N_16071,N_17601);
nand U24284 (N_24284,N_16015,N_15428);
or U24285 (N_24285,N_17918,N_17942);
nand U24286 (N_24286,N_19361,N_18954);
or U24287 (N_24287,N_15628,N_17966);
nand U24288 (N_24288,N_19079,N_19097);
or U24289 (N_24289,N_17963,N_18067);
nor U24290 (N_24290,N_18535,N_19259);
nor U24291 (N_24291,N_16022,N_17068);
nor U24292 (N_24292,N_17861,N_17141);
xnor U24293 (N_24293,N_16423,N_16266);
nor U24294 (N_24294,N_18873,N_17918);
or U24295 (N_24295,N_17839,N_18682);
nand U24296 (N_24296,N_19682,N_18939);
nand U24297 (N_24297,N_17017,N_16658);
and U24298 (N_24298,N_19321,N_19585);
xor U24299 (N_24299,N_16349,N_19142);
nor U24300 (N_24300,N_19384,N_19898);
or U24301 (N_24301,N_17546,N_17951);
or U24302 (N_24302,N_18999,N_16765);
and U24303 (N_24303,N_19675,N_19576);
or U24304 (N_24304,N_16439,N_19845);
nor U24305 (N_24305,N_15390,N_15355);
xor U24306 (N_24306,N_15386,N_17838);
xnor U24307 (N_24307,N_17723,N_15809);
xor U24308 (N_24308,N_17146,N_18420);
or U24309 (N_24309,N_15911,N_16192);
nand U24310 (N_24310,N_16666,N_18768);
nor U24311 (N_24311,N_16652,N_18295);
nand U24312 (N_24312,N_16958,N_17186);
nor U24313 (N_24313,N_18867,N_15665);
and U24314 (N_24314,N_17899,N_19753);
nand U24315 (N_24315,N_18335,N_19798);
nand U24316 (N_24316,N_17513,N_16847);
nor U24317 (N_24317,N_17319,N_15202);
xor U24318 (N_24318,N_19343,N_17165);
or U24319 (N_24319,N_15139,N_16595);
nand U24320 (N_24320,N_16873,N_17305);
nand U24321 (N_24321,N_17965,N_18675);
nor U24322 (N_24322,N_15259,N_18120);
nand U24323 (N_24323,N_16621,N_16816);
or U24324 (N_24324,N_17740,N_15307);
nand U24325 (N_24325,N_19319,N_19738);
and U24326 (N_24326,N_15228,N_16268);
xor U24327 (N_24327,N_15771,N_16765);
nor U24328 (N_24328,N_18118,N_15803);
or U24329 (N_24329,N_16236,N_16260);
nor U24330 (N_24330,N_15528,N_19634);
or U24331 (N_24331,N_16642,N_17545);
nor U24332 (N_24332,N_18885,N_19231);
xnor U24333 (N_24333,N_15547,N_15808);
xnor U24334 (N_24334,N_18279,N_18714);
xor U24335 (N_24335,N_18319,N_17197);
or U24336 (N_24336,N_18542,N_15244);
or U24337 (N_24337,N_17095,N_19872);
and U24338 (N_24338,N_17494,N_18357);
and U24339 (N_24339,N_17870,N_19495);
nor U24340 (N_24340,N_17215,N_15914);
and U24341 (N_24341,N_16146,N_17988);
nand U24342 (N_24342,N_15499,N_17592);
nand U24343 (N_24343,N_19638,N_17755);
or U24344 (N_24344,N_18092,N_17013);
or U24345 (N_24345,N_16583,N_18254);
or U24346 (N_24346,N_19010,N_15841);
or U24347 (N_24347,N_19803,N_16219);
or U24348 (N_24348,N_17965,N_16141);
xor U24349 (N_24349,N_17569,N_17319);
or U24350 (N_24350,N_19118,N_15970);
or U24351 (N_24351,N_19882,N_15627);
or U24352 (N_24352,N_15296,N_15810);
and U24353 (N_24353,N_15707,N_15841);
and U24354 (N_24354,N_16812,N_18158);
and U24355 (N_24355,N_18696,N_17143);
nand U24356 (N_24356,N_18396,N_17234);
nand U24357 (N_24357,N_16085,N_18258);
and U24358 (N_24358,N_16755,N_18809);
and U24359 (N_24359,N_17579,N_18863);
nand U24360 (N_24360,N_16472,N_18864);
nand U24361 (N_24361,N_19616,N_19842);
nand U24362 (N_24362,N_19935,N_19225);
nor U24363 (N_24363,N_19067,N_16178);
nor U24364 (N_24364,N_18376,N_19072);
or U24365 (N_24365,N_15861,N_17990);
nor U24366 (N_24366,N_15185,N_16759);
xnor U24367 (N_24367,N_18409,N_19420);
xor U24368 (N_24368,N_18768,N_17375);
or U24369 (N_24369,N_16114,N_17682);
nor U24370 (N_24370,N_16812,N_17696);
nor U24371 (N_24371,N_15215,N_15743);
nor U24372 (N_24372,N_19490,N_15996);
or U24373 (N_24373,N_18645,N_18831);
or U24374 (N_24374,N_16128,N_19656);
nand U24375 (N_24375,N_15654,N_17554);
nand U24376 (N_24376,N_15457,N_16588);
nand U24377 (N_24377,N_19768,N_17126);
xor U24378 (N_24378,N_15300,N_17078);
nor U24379 (N_24379,N_16686,N_16362);
or U24380 (N_24380,N_16758,N_18735);
nand U24381 (N_24381,N_15882,N_15756);
xnor U24382 (N_24382,N_16686,N_18615);
nand U24383 (N_24383,N_15606,N_19305);
or U24384 (N_24384,N_15547,N_19347);
nand U24385 (N_24385,N_18136,N_17762);
nand U24386 (N_24386,N_17361,N_19000);
nor U24387 (N_24387,N_15261,N_16563);
xor U24388 (N_24388,N_16367,N_18100);
or U24389 (N_24389,N_17618,N_18994);
nor U24390 (N_24390,N_18752,N_15703);
nor U24391 (N_24391,N_17884,N_19805);
or U24392 (N_24392,N_16422,N_19138);
or U24393 (N_24393,N_16533,N_16682);
nor U24394 (N_24394,N_16384,N_16302);
or U24395 (N_24395,N_18471,N_17754);
nand U24396 (N_24396,N_17477,N_18253);
and U24397 (N_24397,N_19949,N_15316);
nand U24398 (N_24398,N_18006,N_15090);
nor U24399 (N_24399,N_19688,N_19099);
nand U24400 (N_24400,N_18470,N_15243);
nor U24401 (N_24401,N_15393,N_15311);
and U24402 (N_24402,N_17943,N_17420);
nand U24403 (N_24403,N_17996,N_16823);
or U24404 (N_24404,N_17004,N_17655);
nand U24405 (N_24405,N_19369,N_19306);
nor U24406 (N_24406,N_16684,N_18027);
xor U24407 (N_24407,N_15339,N_18559);
or U24408 (N_24408,N_16823,N_19180);
nand U24409 (N_24409,N_15970,N_19184);
and U24410 (N_24410,N_16636,N_19616);
xor U24411 (N_24411,N_16053,N_18153);
and U24412 (N_24412,N_17894,N_16451);
nand U24413 (N_24413,N_18578,N_17754);
nor U24414 (N_24414,N_18973,N_17343);
nor U24415 (N_24415,N_19490,N_18103);
and U24416 (N_24416,N_16837,N_17255);
nand U24417 (N_24417,N_16124,N_18134);
and U24418 (N_24418,N_18101,N_18817);
nor U24419 (N_24419,N_15349,N_15180);
and U24420 (N_24420,N_16431,N_16425);
and U24421 (N_24421,N_16597,N_17056);
xnor U24422 (N_24422,N_15608,N_18879);
or U24423 (N_24423,N_19173,N_18425);
nor U24424 (N_24424,N_16540,N_16961);
and U24425 (N_24425,N_18620,N_19333);
nor U24426 (N_24426,N_19735,N_17703);
nand U24427 (N_24427,N_17565,N_19686);
nor U24428 (N_24428,N_18745,N_17395);
xor U24429 (N_24429,N_15809,N_19591);
or U24430 (N_24430,N_18339,N_16061);
and U24431 (N_24431,N_17388,N_17400);
and U24432 (N_24432,N_15028,N_17128);
and U24433 (N_24433,N_16128,N_17602);
or U24434 (N_24434,N_15861,N_16313);
nand U24435 (N_24435,N_15392,N_16565);
nand U24436 (N_24436,N_17178,N_16662);
nand U24437 (N_24437,N_16288,N_17875);
nand U24438 (N_24438,N_19830,N_18594);
nand U24439 (N_24439,N_15057,N_15937);
nor U24440 (N_24440,N_15715,N_18453);
nand U24441 (N_24441,N_19922,N_18140);
nor U24442 (N_24442,N_19422,N_18166);
nor U24443 (N_24443,N_15751,N_19308);
and U24444 (N_24444,N_19621,N_16592);
or U24445 (N_24445,N_15422,N_19812);
or U24446 (N_24446,N_17508,N_18922);
nand U24447 (N_24447,N_15241,N_15161);
nand U24448 (N_24448,N_17808,N_17497);
xnor U24449 (N_24449,N_17588,N_18183);
or U24450 (N_24450,N_15246,N_19613);
and U24451 (N_24451,N_15934,N_15330);
nor U24452 (N_24452,N_15452,N_17183);
nor U24453 (N_24453,N_15654,N_17385);
nand U24454 (N_24454,N_16149,N_17211);
nor U24455 (N_24455,N_18196,N_17259);
nand U24456 (N_24456,N_17243,N_17628);
or U24457 (N_24457,N_18057,N_17091);
nand U24458 (N_24458,N_17868,N_19793);
nor U24459 (N_24459,N_19967,N_19050);
and U24460 (N_24460,N_15761,N_17889);
nor U24461 (N_24461,N_19325,N_16865);
xnor U24462 (N_24462,N_18063,N_16478);
xnor U24463 (N_24463,N_16326,N_17568);
nor U24464 (N_24464,N_16919,N_15906);
and U24465 (N_24465,N_15641,N_18350);
nand U24466 (N_24466,N_15592,N_19334);
and U24467 (N_24467,N_17371,N_16233);
nor U24468 (N_24468,N_16799,N_19235);
nand U24469 (N_24469,N_16181,N_18332);
xnor U24470 (N_24470,N_15917,N_15643);
nand U24471 (N_24471,N_15765,N_19859);
nand U24472 (N_24472,N_17840,N_16565);
or U24473 (N_24473,N_17014,N_19163);
nand U24474 (N_24474,N_16992,N_17428);
or U24475 (N_24475,N_19637,N_17226);
nor U24476 (N_24476,N_17532,N_16723);
and U24477 (N_24477,N_16515,N_17409);
xnor U24478 (N_24478,N_18145,N_16349);
nand U24479 (N_24479,N_19433,N_18950);
or U24480 (N_24480,N_16244,N_18180);
nor U24481 (N_24481,N_17399,N_19287);
nand U24482 (N_24482,N_19858,N_16484);
nor U24483 (N_24483,N_19022,N_15730);
and U24484 (N_24484,N_18315,N_18502);
nor U24485 (N_24485,N_15340,N_17249);
nand U24486 (N_24486,N_17627,N_16625);
or U24487 (N_24487,N_16176,N_19682);
and U24488 (N_24488,N_19906,N_18687);
or U24489 (N_24489,N_18133,N_16401);
nor U24490 (N_24490,N_15138,N_19746);
or U24491 (N_24491,N_16571,N_15964);
nand U24492 (N_24492,N_18154,N_16618);
and U24493 (N_24493,N_15534,N_19507);
nor U24494 (N_24494,N_18148,N_17817);
nor U24495 (N_24495,N_19314,N_15479);
nor U24496 (N_24496,N_15487,N_16553);
and U24497 (N_24497,N_18330,N_19132);
xor U24498 (N_24498,N_19305,N_16318);
xnor U24499 (N_24499,N_15586,N_18449);
nor U24500 (N_24500,N_17086,N_19941);
nor U24501 (N_24501,N_17832,N_16743);
or U24502 (N_24502,N_19229,N_15308);
and U24503 (N_24503,N_18285,N_18593);
or U24504 (N_24504,N_18936,N_16684);
and U24505 (N_24505,N_15705,N_17811);
nand U24506 (N_24506,N_15676,N_16845);
nor U24507 (N_24507,N_18742,N_15209);
and U24508 (N_24508,N_16322,N_17231);
or U24509 (N_24509,N_15752,N_18327);
and U24510 (N_24510,N_18621,N_17305);
nand U24511 (N_24511,N_19562,N_15888);
and U24512 (N_24512,N_17499,N_19242);
or U24513 (N_24513,N_16335,N_17631);
and U24514 (N_24514,N_18676,N_16140);
and U24515 (N_24515,N_15338,N_16815);
or U24516 (N_24516,N_15093,N_19569);
nor U24517 (N_24517,N_18882,N_16505);
nor U24518 (N_24518,N_16408,N_19300);
and U24519 (N_24519,N_17636,N_18313);
or U24520 (N_24520,N_15033,N_16216);
or U24521 (N_24521,N_19301,N_16701);
nor U24522 (N_24522,N_16103,N_18793);
nor U24523 (N_24523,N_19294,N_19461);
nor U24524 (N_24524,N_15241,N_16697);
or U24525 (N_24525,N_19915,N_15382);
or U24526 (N_24526,N_16425,N_17563);
nand U24527 (N_24527,N_16875,N_17070);
and U24528 (N_24528,N_19531,N_17224);
or U24529 (N_24529,N_19542,N_19037);
nor U24530 (N_24530,N_16891,N_15557);
nand U24531 (N_24531,N_16535,N_15857);
nor U24532 (N_24532,N_19646,N_17598);
nor U24533 (N_24533,N_17534,N_15820);
or U24534 (N_24534,N_15833,N_16900);
or U24535 (N_24535,N_18129,N_18396);
nor U24536 (N_24536,N_18909,N_15178);
nor U24537 (N_24537,N_19887,N_18555);
nor U24538 (N_24538,N_18402,N_18454);
and U24539 (N_24539,N_15720,N_16850);
nand U24540 (N_24540,N_15460,N_18206);
nand U24541 (N_24541,N_19929,N_19946);
nand U24542 (N_24542,N_17893,N_17158);
and U24543 (N_24543,N_15886,N_18000);
nor U24544 (N_24544,N_16773,N_19599);
nand U24545 (N_24545,N_17622,N_17713);
nor U24546 (N_24546,N_16382,N_17503);
or U24547 (N_24547,N_19935,N_15089);
or U24548 (N_24548,N_16472,N_15105);
xnor U24549 (N_24549,N_16516,N_18375);
and U24550 (N_24550,N_16891,N_19308);
nor U24551 (N_24551,N_15928,N_17241);
or U24552 (N_24552,N_18314,N_16311);
or U24553 (N_24553,N_18387,N_19937);
nor U24554 (N_24554,N_15519,N_19983);
nand U24555 (N_24555,N_19038,N_19278);
and U24556 (N_24556,N_16593,N_18972);
or U24557 (N_24557,N_17547,N_16693);
and U24558 (N_24558,N_18554,N_19028);
or U24559 (N_24559,N_19638,N_18249);
nand U24560 (N_24560,N_16009,N_19476);
and U24561 (N_24561,N_15211,N_15740);
and U24562 (N_24562,N_15392,N_16779);
nand U24563 (N_24563,N_15313,N_16387);
or U24564 (N_24564,N_18815,N_19570);
nand U24565 (N_24565,N_15060,N_19117);
xor U24566 (N_24566,N_16778,N_18375);
nor U24567 (N_24567,N_15764,N_16505);
nand U24568 (N_24568,N_16711,N_17589);
nor U24569 (N_24569,N_15427,N_17157);
or U24570 (N_24570,N_18692,N_19807);
or U24571 (N_24571,N_17437,N_18190);
or U24572 (N_24572,N_17779,N_17775);
and U24573 (N_24573,N_17676,N_19040);
nor U24574 (N_24574,N_19259,N_16908);
or U24575 (N_24575,N_18904,N_15867);
or U24576 (N_24576,N_18097,N_15158);
nand U24577 (N_24577,N_17218,N_15654);
nand U24578 (N_24578,N_16570,N_15900);
xor U24579 (N_24579,N_19727,N_18496);
nand U24580 (N_24580,N_15210,N_19807);
xnor U24581 (N_24581,N_17934,N_15717);
nor U24582 (N_24582,N_17025,N_17874);
nand U24583 (N_24583,N_19344,N_18500);
nand U24584 (N_24584,N_19179,N_18583);
and U24585 (N_24585,N_18309,N_18705);
xor U24586 (N_24586,N_17072,N_19013);
xor U24587 (N_24587,N_19177,N_17680);
nor U24588 (N_24588,N_16240,N_17600);
xnor U24589 (N_24589,N_18576,N_16674);
or U24590 (N_24590,N_18613,N_17322);
and U24591 (N_24591,N_17994,N_16788);
nand U24592 (N_24592,N_18386,N_17397);
nand U24593 (N_24593,N_16698,N_19493);
and U24594 (N_24594,N_18426,N_15789);
nor U24595 (N_24595,N_17004,N_15044);
nor U24596 (N_24596,N_18520,N_16606);
nor U24597 (N_24597,N_18734,N_19859);
or U24598 (N_24598,N_15062,N_16672);
and U24599 (N_24599,N_19097,N_15294);
and U24600 (N_24600,N_17808,N_16911);
nand U24601 (N_24601,N_19302,N_16416);
and U24602 (N_24602,N_19891,N_19965);
nor U24603 (N_24603,N_15434,N_18951);
or U24604 (N_24604,N_15460,N_15577);
or U24605 (N_24605,N_19322,N_18889);
or U24606 (N_24606,N_19441,N_17076);
nand U24607 (N_24607,N_15759,N_18373);
nor U24608 (N_24608,N_19583,N_16561);
or U24609 (N_24609,N_16202,N_18927);
or U24610 (N_24610,N_19067,N_15518);
or U24611 (N_24611,N_17112,N_18948);
nor U24612 (N_24612,N_19866,N_15099);
nand U24613 (N_24613,N_15258,N_16013);
nor U24614 (N_24614,N_19256,N_16635);
and U24615 (N_24615,N_16330,N_18078);
and U24616 (N_24616,N_18818,N_18040);
nand U24617 (N_24617,N_18817,N_19895);
nor U24618 (N_24618,N_15719,N_15164);
nand U24619 (N_24619,N_17936,N_18944);
or U24620 (N_24620,N_18504,N_17198);
nor U24621 (N_24621,N_19718,N_16083);
nand U24622 (N_24622,N_16195,N_17777);
and U24623 (N_24623,N_16380,N_15218);
nor U24624 (N_24624,N_17095,N_19994);
or U24625 (N_24625,N_16576,N_18550);
nand U24626 (N_24626,N_17075,N_17258);
nor U24627 (N_24627,N_16045,N_17161);
xor U24628 (N_24628,N_17944,N_15069);
or U24629 (N_24629,N_17943,N_18462);
or U24630 (N_24630,N_16733,N_17551);
nand U24631 (N_24631,N_17926,N_17792);
and U24632 (N_24632,N_19410,N_16334);
and U24633 (N_24633,N_19173,N_17043);
or U24634 (N_24634,N_16024,N_15572);
nand U24635 (N_24635,N_19377,N_19267);
nand U24636 (N_24636,N_15740,N_19696);
and U24637 (N_24637,N_19386,N_19041);
or U24638 (N_24638,N_17804,N_15037);
xor U24639 (N_24639,N_16116,N_18454);
nor U24640 (N_24640,N_17564,N_15766);
and U24641 (N_24641,N_19096,N_17592);
nand U24642 (N_24642,N_15565,N_15937);
nand U24643 (N_24643,N_15003,N_16578);
nor U24644 (N_24644,N_18150,N_17019);
nand U24645 (N_24645,N_16520,N_15856);
or U24646 (N_24646,N_15909,N_17314);
nand U24647 (N_24647,N_15849,N_16425);
or U24648 (N_24648,N_17208,N_17682);
xnor U24649 (N_24649,N_16065,N_19737);
nand U24650 (N_24650,N_15044,N_15408);
and U24651 (N_24651,N_18099,N_18514);
nand U24652 (N_24652,N_16632,N_19476);
nand U24653 (N_24653,N_17615,N_19954);
or U24654 (N_24654,N_17277,N_17825);
and U24655 (N_24655,N_16028,N_16250);
nor U24656 (N_24656,N_15318,N_18042);
nor U24657 (N_24657,N_16696,N_18330);
and U24658 (N_24658,N_16425,N_19953);
nor U24659 (N_24659,N_16012,N_19958);
nand U24660 (N_24660,N_17469,N_16895);
nand U24661 (N_24661,N_17544,N_18391);
nor U24662 (N_24662,N_15047,N_19196);
or U24663 (N_24663,N_19038,N_17950);
xnor U24664 (N_24664,N_19755,N_17667);
nor U24665 (N_24665,N_16151,N_18954);
and U24666 (N_24666,N_16501,N_15354);
nand U24667 (N_24667,N_16988,N_17206);
nor U24668 (N_24668,N_17313,N_19318);
or U24669 (N_24669,N_18163,N_18025);
or U24670 (N_24670,N_15658,N_18866);
or U24671 (N_24671,N_17912,N_18477);
and U24672 (N_24672,N_15615,N_15839);
nand U24673 (N_24673,N_18143,N_18900);
nand U24674 (N_24674,N_16846,N_16799);
or U24675 (N_24675,N_16482,N_18882);
nor U24676 (N_24676,N_17825,N_16460);
nor U24677 (N_24677,N_18436,N_15269);
nand U24678 (N_24678,N_16004,N_15795);
or U24679 (N_24679,N_18770,N_15082);
nand U24680 (N_24680,N_15072,N_18222);
nand U24681 (N_24681,N_16892,N_16354);
and U24682 (N_24682,N_19387,N_19033);
or U24683 (N_24683,N_17296,N_16129);
nor U24684 (N_24684,N_18500,N_18611);
nand U24685 (N_24685,N_19366,N_15518);
nor U24686 (N_24686,N_15853,N_15743);
and U24687 (N_24687,N_17895,N_18784);
or U24688 (N_24688,N_16860,N_16269);
and U24689 (N_24689,N_15424,N_15997);
or U24690 (N_24690,N_15430,N_19295);
and U24691 (N_24691,N_16432,N_19783);
or U24692 (N_24692,N_15465,N_15220);
or U24693 (N_24693,N_18047,N_15350);
and U24694 (N_24694,N_15223,N_17849);
nor U24695 (N_24695,N_19132,N_17464);
or U24696 (N_24696,N_17716,N_19266);
and U24697 (N_24697,N_19033,N_19931);
and U24698 (N_24698,N_17715,N_15446);
xnor U24699 (N_24699,N_15565,N_18330);
nand U24700 (N_24700,N_19689,N_17450);
nand U24701 (N_24701,N_17028,N_18180);
nor U24702 (N_24702,N_15613,N_18786);
or U24703 (N_24703,N_16594,N_16539);
nand U24704 (N_24704,N_18644,N_19161);
nor U24705 (N_24705,N_18351,N_15215);
and U24706 (N_24706,N_19386,N_15454);
or U24707 (N_24707,N_17883,N_16558);
nor U24708 (N_24708,N_16523,N_18285);
or U24709 (N_24709,N_19397,N_19592);
nand U24710 (N_24710,N_15495,N_19762);
xor U24711 (N_24711,N_15428,N_19008);
and U24712 (N_24712,N_18472,N_17056);
nor U24713 (N_24713,N_18671,N_16335);
and U24714 (N_24714,N_17686,N_15857);
and U24715 (N_24715,N_18394,N_19197);
nand U24716 (N_24716,N_16835,N_19369);
or U24717 (N_24717,N_18430,N_16424);
nand U24718 (N_24718,N_17100,N_19299);
or U24719 (N_24719,N_15159,N_18215);
nand U24720 (N_24720,N_17825,N_17684);
nor U24721 (N_24721,N_18528,N_19216);
and U24722 (N_24722,N_15710,N_17266);
or U24723 (N_24723,N_16170,N_16023);
nand U24724 (N_24724,N_18546,N_16960);
xor U24725 (N_24725,N_15324,N_19416);
and U24726 (N_24726,N_17492,N_19175);
and U24727 (N_24727,N_16478,N_16738);
xor U24728 (N_24728,N_17809,N_15974);
or U24729 (N_24729,N_18162,N_17052);
or U24730 (N_24730,N_15032,N_18115);
xor U24731 (N_24731,N_17365,N_16756);
nand U24732 (N_24732,N_16898,N_19093);
xor U24733 (N_24733,N_18658,N_16791);
nand U24734 (N_24734,N_19602,N_15680);
nor U24735 (N_24735,N_19339,N_17576);
nor U24736 (N_24736,N_15126,N_16753);
nand U24737 (N_24737,N_17352,N_16385);
xnor U24738 (N_24738,N_18035,N_18113);
nand U24739 (N_24739,N_19865,N_18865);
or U24740 (N_24740,N_16413,N_17582);
and U24741 (N_24741,N_17588,N_16809);
xnor U24742 (N_24742,N_17109,N_17475);
nand U24743 (N_24743,N_19888,N_19835);
and U24744 (N_24744,N_18015,N_18371);
or U24745 (N_24745,N_15122,N_19284);
and U24746 (N_24746,N_18736,N_18837);
nand U24747 (N_24747,N_15377,N_18894);
nand U24748 (N_24748,N_17961,N_16846);
and U24749 (N_24749,N_15657,N_17741);
nand U24750 (N_24750,N_18572,N_16185);
nand U24751 (N_24751,N_17608,N_18905);
or U24752 (N_24752,N_16507,N_17612);
and U24753 (N_24753,N_16101,N_17913);
nand U24754 (N_24754,N_16127,N_15334);
nor U24755 (N_24755,N_17267,N_16494);
nor U24756 (N_24756,N_16599,N_15339);
nand U24757 (N_24757,N_19134,N_17461);
nand U24758 (N_24758,N_16599,N_17980);
or U24759 (N_24759,N_18135,N_19622);
and U24760 (N_24760,N_15502,N_19397);
xor U24761 (N_24761,N_19359,N_17523);
or U24762 (N_24762,N_15712,N_15001);
nand U24763 (N_24763,N_19906,N_15398);
or U24764 (N_24764,N_16261,N_16278);
or U24765 (N_24765,N_15612,N_17098);
nor U24766 (N_24766,N_18753,N_16322);
and U24767 (N_24767,N_18838,N_15672);
and U24768 (N_24768,N_18535,N_19323);
and U24769 (N_24769,N_17560,N_18576);
nor U24770 (N_24770,N_18654,N_16707);
or U24771 (N_24771,N_15424,N_19921);
and U24772 (N_24772,N_17690,N_18914);
nor U24773 (N_24773,N_19084,N_15193);
nor U24774 (N_24774,N_18739,N_19984);
and U24775 (N_24775,N_15239,N_18412);
nand U24776 (N_24776,N_16644,N_17537);
xor U24777 (N_24777,N_15228,N_18435);
nand U24778 (N_24778,N_15478,N_17853);
and U24779 (N_24779,N_19368,N_18693);
nand U24780 (N_24780,N_15866,N_17170);
nand U24781 (N_24781,N_16660,N_15279);
nor U24782 (N_24782,N_15076,N_17869);
xor U24783 (N_24783,N_18122,N_15382);
nor U24784 (N_24784,N_18478,N_17780);
nor U24785 (N_24785,N_19510,N_17658);
or U24786 (N_24786,N_17267,N_18769);
nor U24787 (N_24787,N_17212,N_18003);
nor U24788 (N_24788,N_15856,N_19799);
nand U24789 (N_24789,N_15412,N_15254);
and U24790 (N_24790,N_19864,N_15877);
nor U24791 (N_24791,N_16661,N_17765);
or U24792 (N_24792,N_17094,N_15806);
xnor U24793 (N_24793,N_17780,N_15810);
or U24794 (N_24794,N_18902,N_16410);
nand U24795 (N_24795,N_18073,N_18302);
and U24796 (N_24796,N_18778,N_17967);
or U24797 (N_24797,N_17131,N_19176);
nor U24798 (N_24798,N_19852,N_18664);
or U24799 (N_24799,N_17934,N_17499);
nor U24800 (N_24800,N_17349,N_17364);
or U24801 (N_24801,N_19325,N_18251);
and U24802 (N_24802,N_15342,N_17329);
nor U24803 (N_24803,N_19186,N_17860);
xnor U24804 (N_24804,N_19173,N_15524);
nand U24805 (N_24805,N_19309,N_19989);
and U24806 (N_24806,N_18597,N_16417);
or U24807 (N_24807,N_18495,N_18592);
and U24808 (N_24808,N_15821,N_15977);
nand U24809 (N_24809,N_16727,N_16404);
nor U24810 (N_24810,N_15525,N_19922);
nor U24811 (N_24811,N_18559,N_19771);
nand U24812 (N_24812,N_16206,N_15764);
nor U24813 (N_24813,N_17148,N_18561);
nor U24814 (N_24814,N_19864,N_19400);
nand U24815 (N_24815,N_18592,N_19168);
nand U24816 (N_24816,N_18943,N_15674);
nor U24817 (N_24817,N_19808,N_15193);
and U24818 (N_24818,N_15204,N_19265);
nand U24819 (N_24819,N_16676,N_19819);
nand U24820 (N_24820,N_17335,N_16807);
or U24821 (N_24821,N_16714,N_16890);
or U24822 (N_24822,N_16463,N_18127);
nand U24823 (N_24823,N_15810,N_18886);
nor U24824 (N_24824,N_19568,N_18250);
nor U24825 (N_24825,N_15981,N_16899);
or U24826 (N_24826,N_16136,N_16229);
nor U24827 (N_24827,N_17533,N_19595);
or U24828 (N_24828,N_15032,N_19880);
and U24829 (N_24829,N_19542,N_19715);
or U24830 (N_24830,N_19800,N_15077);
nor U24831 (N_24831,N_18455,N_18995);
nand U24832 (N_24832,N_17884,N_15616);
xnor U24833 (N_24833,N_15887,N_18289);
or U24834 (N_24834,N_16356,N_18629);
and U24835 (N_24835,N_17435,N_17451);
or U24836 (N_24836,N_18848,N_15551);
and U24837 (N_24837,N_16967,N_18592);
or U24838 (N_24838,N_19431,N_18005);
or U24839 (N_24839,N_17401,N_16096);
nand U24840 (N_24840,N_16768,N_19203);
nor U24841 (N_24841,N_17562,N_19813);
or U24842 (N_24842,N_17900,N_16230);
nor U24843 (N_24843,N_16552,N_19346);
nand U24844 (N_24844,N_18357,N_17299);
nor U24845 (N_24845,N_16431,N_17998);
and U24846 (N_24846,N_17433,N_16755);
nor U24847 (N_24847,N_16093,N_16354);
nor U24848 (N_24848,N_15128,N_19665);
nand U24849 (N_24849,N_15995,N_18205);
and U24850 (N_24850,N_17485,N_19560);
and U24851 (N_24851,N_17091,N_17416);
or U24852 (N_24852,N_16421,N_17066);
nand U24853 (N_24853,N_19481,N_19307);
nor U24854 (N_24854,N_16467,N_19588);
nand U24855 (N_24855,N_17193,N_19779);
nor U24856 (N_24856,N_17092,N_18832);
nor U24857 (N_24857,N_18407,N_18475);
and U24858 (N_24858,N_16663,N_15404);
or U24859 (N_24859,N_18806,N_15350);
nand U24860 (N_24860,N_18522,N_19270);
nor U24861 (N_24861,N_19438,N_16792);
and U24862 (N_24862,N_17938,N_16065);
nand U24863 (N_24863,N_16982,N_17366);
and U24864 (N_24864,N_15416,N_17269);
nand U24865 (N_24865,N_17129,N_18448);
nand U24866 (N_24866,N_15583,N_15716);
nand U24867 (N_24867,N_15659,N_16564);
and U24868 (N_24868,N_19194,N_17233);
or U24869 (N_24869,N_15384,N_15694);
nand U24870 (N_24870,N_19533,N_16617);
and U24871 (N_24871,N_16533,N_18186);
or U24872 (N_24872,N_15727,N_15197);
nor U24873 (N_24873,N_16264,N_17692);
nand U24874 (N_24874,N_15564,N_16366);
nand U24875 (N_24875,N_16616,N_15938);
nand U24876 (N_24876,N_16163,N_16104);
xnor U24877 (N_24877,N_17618,N_16681);
nand U24878 (N_24878,N_17261,N_18698);
nand U24879 (N_24879,N_16138,N_15559);
xnor U24880 (N_24880,N_18892,N_18906);
nor U24881 (N_24881,N_19207,N_19291);
xor U24882 (N_24882,N_16317,N_17573);
and U24883 (N_24883,N_19655,N_15683);
xnor U24884 (N_24884,N_16983,N_18982);
nor U24885 (N_24885,N_19352,N_15614);
or U24886 (N_24886,N_17802,N_17519);
or U24887 (N_24887,N_19906,N_17760);
and U24888 (N_24888,N_16051,N_19699);
and U24889 (N_24889,N_19619,N_19297);
nor U24890 (N_24890,N_15377,N_18925);
or U24891 (N_24891,N_18499,N_17562);
nor U24892 (N_24892,N_18986,N_17216);
and U24893 (N_24893,N_18229,N_15718);
xnor U24894 (N_24894,N_19368,N_19179);
or U24895 (N_24895,N_19816,N_15208);
xor U24896 (N_24896,N_17331,N_16287);
nor U24897 (N_24897,N_17391,N_19413);
and U24898 (N_24898,N_18690,N_19015);
nor U24899 (N_24899,N_18986,N_15116);
nand U24900 (N_24900,N_18933,N_16610);
or U24901 (N_24901,N_16357,N_15031);
xnor U24902 (N_24902,N_18695,N_17879);
and U24903 (N_24903,N_17728,N_17582);
nand U24904 (N_24904,N_17957,N_17032);
nor U24905 (N_24905,N_17685,N_16427);
nor U24906 (N_24906,N_19756,N_17166);
nor U24907 (N_24907,N_17529,N_18328);
xnor U24908 (N_24908,N_15521,N_18150);
nand U24909 (N_24909,N_15584,N_19295);
nand U24910 (N_24910,N_16313,N_17198);
nand U24911 (N_24911,N_17157,N_18130);
and U24912 (N_24912,N_18747,N_18489);
nand U24913 (N_24913,N_18212,N_15407);
nor U24914 (N_24914,N_18301,N_19454);
nand U24915 (N_24915,N_15296,N_17506);
and U24916 (N_24916,N_19376,N_17721);
nand U24917 (N_24917,N_18868,N_17315);
or U24918 (N_24918,N_15397,N_18375);
nor U24919 (N_24919,N_15877,N_15817);
xor U24920 (N_24920,N_19573,N_15471);
nand U24921 (N_24921,N_16656,N_19841);
nand U24922 (N_24922,N_17425,N_19158);
and U24923 (N_24923,N_16881,N_18409);
and U24924 (N_24924,N_15908,N_15904);
nand U24925 (N_24925,N_17092,N_16113);
or U24926 (N_24926,N_19627,N_19643);
and U24927 (N_24927,N_16700,N_19584);
nor U24928 (N_24928,N_16832,N_16147);
nand U24929 (N_24929,N_19591,N_17531);
or U24930 (N_24930,N_19241,N_16906);
nor U24931 (N_24931,N_18920,N_19121);
nor U24932 (N_24932,N_18786,N_19318);
nand U24933 (N_24933,N_15719,N_17404);
nor U24934 (N_24934,N_17318,N_16454);
xor U24935 (N_24935,N_18665,N_16242);
nand U24936 (N_24936,N_19528,N_18664);
nand U24937 (N_24937,N_17741,N_18608);
nor U24938 (N_24938,N_19333,N_15202);
or U24939 (N_24939,N_17177,N_16283);
or U24940 (N_24940,N_19997,N_15622);
and U24941 (N_24941,N_18764,N_15135);
or U24942 (N_24942,N_19633,N_16120);
and U24943 (N_24943,N_19660,N_18673);
or U24944 (N_24944,N_17709,N_16810);
nor U24945 (N_24945,N_15788,N_18387);
xnor U24946 (N_24946,N_15045,N_17439);
or U24947 (N_24947,N_19442,N_16344);
nand U24948 (N_24948,N_15366,N_17825);
nand U24949 (N_24949,N_15817,N_16068);
nor U24950 (N_24950,N_16038,N_18187);
nor U24951 (N_24951,N_17175,N_15875);
nor U24952 (N_24952,N_16854,N_17734);
nor U24953 (N_24953,N_16547,N_16571);
xnor U24954 (N_24954,N_18497,N_17924);
nand U24955 (N_24955,N_17014,N_18281);
and U24956 (N_24956,N_19414,N_16011);
xor U24957 (N_24957,N_17055,N_19871);
and U24958 (N_24958,N_18999,N_18828);
nor U24959 (N_24959,N_15617,N_18695);
or U24960 (N_24960,N_16572,N_15157);
or U24961 (N_24961,N_15254,N_17779);
or U24962 (N_24962,N_16246,N_15595);
or U24963 (N_24963,N_15187,N_17486);
nor U24964 (N_24964,N_17149,N_15326);
nand U24965 (N_24965,N_17115,N_16702);
and U24966 (N_24966,N_15626,N_18129);
or U24967 (N_24967,N_17056,N_15201);
or U24968 (N_24968,N_18846,N_18629);
and U24969 (N_24969,N_19383,N_15686);
or U24970 (N_24970,N_18833,N_16042);
and U24971 (N_24971,N_15838,N_16572);
nand U24972 (N_24972,N_18306,N_15905);
and U24973 (N_24973,N_19243,N_16164);
or U24974 (N_24974,N_16770,N_19982);
and U24975 (N_24975,N_18367,N_15256);
nor U24976 (N_24976,N_15884,N_17715);
or U24977 (N_24977,N_19865,N_19944);
and U24978 (N_24978,N_17314,N_16631);
xnor U24979 (N_24979,N_17266,N_15750);
and U24980 (N_24980,N_18458,N_19138);
xor U24981 (N_24981,N_15808,N_18305);
nand U24982 (N_24982,N_17070,N_19167);
nor U24983 (N_24983,N_19429,N_15404);
nor U24984 (N_24984,N_19168,N_19282);
or U24985 (N_24985,N_19904,N_18088);
or U24986 (N_24986,N_17490,N_17537);
and U24987 (N_24987,N_18217,N_19392);
and U24988 (N_24988,N_19713,N_16499);
nor U24989 (N_24989,N_18138,N_19029);
xnor U24990 (N_24990,N_16782,N_17022);
and U24991 (N_24991,N_16869,N_19396);
nor U24992 (N_24992,N_19364,N_17462);
and U24993 (N_24993,N_15810,N_18149);
nand U24994 (N_24994,N_15297,N_17502);
and U24995 (N_24995,N_17725,N_16521);
nor U24996 (N_24996,N_19753,N_17653);
and U24997 (N_24997,N_16712,N_17508);
and U24998 (N_24998,N_15041,N_18198);
or U24999 (N_24999,N_17857,N_16136);
nor U25000 (N_25000,N_24236,N_23776);
nand U25001 (N_25001,N_22603,N_21643);
nor U25002 (N_25002,N_22755,N_21163);
or U25003 (N_25003,N_20666,N_22747);
nor U25004 (N_25004,N_23125,N_22231);
or U25005 (N_25005,N_21709,N_20795);
or U25006 (N_25006,N_20099,N_24521);
and U25007 (N_25007,N_23740,N_20202);
and U25008 (N_25008,N_20293,N_22452);
xor U25009 (N_25009,N_24422,N_23062);
or U25010 (N_25010,N_22919,N_20005);
and U25011 (N_25011,N_20451,N_20053);
xnor U25012 (N_25012,N_22869,N_21903);
or U25013 (N_25013,N_22376,N_23605);
nor U25014 (N_25014,N_24279,N_22709);
xnor U25015 (N_25015,N_24974,N_22162);
or U25016 (N_25016,N_24057,N_20253);
and U25017 (N_25017,N_21500,N_24770);
nor U25018 (N_25018,N_22959,N_21898);
xor U25019 (N_25019,N_23826,N_23811);
and U25020 (N_25020,N_23500,N_22088);
nand U25021 (N_25021,N_22722,N_20204);
xnor U25022 (N_25022,N_21043,N_20529);
nor U25023 (N_25023,N_21371,N_22170);
or U25024 (N_25024,N_24217,N_21368);
and U25025 (N_25025,N_22768,N_23029);
nor U25026 (N_25026,N_20872,N_23867);
or U25027 (N_25027,N_20558,N_20238);
nand U25028 (N_25028,N_22730,N_20320);
and U25029 (N_25029,N_22699,N_24448);
xnor U25030 (N_25030,N_22202,N_24443);
nor U25031 (N_25031,N_21394,N_21991);
nand U25032 (N_25032,N_23434,N_23839);
and U25033 (N_25033,N_23172,N_24640);
nand U25034 (N_25034,N_24728,N_21621);
or U25035 (N_25035,N_24717,N_20598);
nand U25036 (N_25036,N_22431,N_20746);
and U25037 (N_25037,N_24153,N_23326);
and U25038 (N_25038,N_23938,N_21876);
or U25039 (N_25039,N_20607,N_22296);
nor U25040 (N_25040,N_22106,N_23520);
or U25041 (N_25041,N_20941,N_23182);
or U25042 (N_25042,N_22800,N_21782);
nand U25043 (N_25043,N_20863,N_22311);
and U25044 (N_25044,N_23561,N_24827);
or U25045 (N_25045,N_23374,N_22200);
nand U25046 (N_25046,N_23307,N_20290);
nor U25047 (N_25047,N_21370,N_21383);
and U25048 (N_25048,N_21421,N_23926);
and U25049 (N_25049,N_24987,N_24199);
nor U25050 (N_25050,N_22134,N_24470);
or U25051 (N_25051,N_22551,N_24067);
nor U25052 (N_25052,N_20868,N_22865);
nor U25053 (N_25053,N_24274,N_20312);
and U25054 (N_25054,N_20562,N_24201);
xnor U25055 (N_25055,N_22460,N_20057);
nand U25056 (N_25056,N_21946,N_24505);
nor U25057 (N_25057,N_20786,N_23211);
nand U25058 (N_25058,N_21183,N_21753);
nor U25059 (N_25059,N_22986,N_20142);
and U25060 (N_25060,N_20192,N_21649);
nand U25061 (N_25061,N_24726,N_24400);
nor U25062 (N_25062,N_21377,N_21061);
nor U25063 (N_25063,N_23831,N_24925);
nor U25064 (N_25064,N_20663,N_23693);
and U25065 (N_25065,N_24897,N_22928);
nor U25066 (N_25066,N_23198,N_20223);
or U25067 (N_25067,N_22856,N_22258);
and U25068 (N_25068,N_20844,N_21119);
or U25069 (N_25069,N_24347,N_21286);
or U25070 (N_25070,N_24024,N_22118);
nor U25071 (N_25071,N_24808,N_20662);
and U25072 (N_25072,N_21622,N_24494);
nor U25073 (N_25073,N_21954,N_21740);
nand U25074 (N_25074,N_21335,N_22314);
xnor U25075 (N_25075,N_22562,N_22904);
nor U25076 (N_25076,N_22353,N_20186);
or U25077 (N_25077,N_22802,N_20788);
nor U25078 (N_25078,N_20163,N_22899);
or U25079 (N_25079,N_22714,N_24797);
nand U25080 (N_25080,N_20027,N_22135);
or U25081 (N_25081,N_23636,N_20028);
nor U25082 (N_25082,N_20035,N_24791);
nand U25083 (N_25083,N_20898,N_20498);
nand U25084 (N_25084,N_23408,N_23643);
and U25085 (N_25085,N_23228,N_24957);
or U25086 (N_25086,N_20535,N_20675);
nor U25087 (N_25087,N_20507,N_20782);
or U25088 (N_25088,N_22557,N_24600);
and U25089 (N_25089,N_24331,N_24625);
or U25090 (N_25090,N_20383,N_24014);
and U25091 (N_25091,N_24094,N_20148);
and U25092 (N_25092,N_22401,N_23541);
nand U25093 (N_25093,N_23925,N_21730);
nand U25094 (N_25094,N_21262,N_22574);
and U25095 (N_25095,N_23240,N_22512);
or U25096 (N_25096,N_21748,N_21463);
nand U25097 (N_25097,N_23470,N_20232);
nor U25098 (N_25098,N_20984,N_23503);
nand U25099 (N_25099,N_24363,N_23004);
or U25100 (N_25100,N_20358,N_21322);
or U25101 (N_25101,N_20780,N_20632);
or U25102 (N_25102,N_24139,N_21582);
xnor U25103 (N_25103,N_24665,N_22659);
nand U25104 (N_25104,N_20551,N_22068);
or U25105 (N_25105,N_24003,N_20974);
nor U25106 (N_25106,N_23622,N_21082);
and U25107 (N_25107,N_24305,N_24580);
nor U25108 (N_25108,N_23401,N_22408);
and U25109 (N_25109,N_22176,N_23331);
nand U25110 (N_25110,N_24106,N_22742);
xnor U25111 (N_25111,N_22708,N_23412);
nand U25112 (N_25112,N_24446,N_20855);
nor U25113 (N_25113,N_24175,N_24992);
nand U25114 (N_25114,N_24899,N_21080);
and U25115 (N_25115,N_21710,N_21382);
nor U25116 (N_25116,N_22195,N_22846);
nor U25117 (N_25117,N_21442,N_24032);
and U25118 (N_25118,N_21102,N_22977);
or U25119 (N_25119,N_24645,N_20416);
nand U25120 (N_25120,N_22395,N_21074);
nor U25121 (N_25121,N_23480,N_22837);
or U25122 (N_25122,N_20015,N_21677);
and U25123 (N_25123,N_23661,N_21881);
nand U25124 (N_25124,N_24076,N_24068);
nor U25125 (N_25125,N_23965,N_22669);
or U25126 (N_25126,N_24491,N_23651);
xor U25127 (N_25127,N_24434,N_24906);
or U25128 (N_25128,N_24504,N_22500);
nand U25129 (N_25129,N_22864,N_24046);
or U25130 (N_25130,N_21676,N_21819);
or U25131 (N_25131,N_24315,N_24870);
nand U25132 (N_25132,N_20145,N_21591);
nor U25133 (N_25133,N_21755,N_24276);
nand U25134 (N_25134,N_22850,N_22234);
nor U25135 (N_25135,N_23532,N_22434);
nand U25136 (N_25136,N_24069,N_20164);
or U25137 (N_25137,N_21540,N_22984);
nand U25138 (N_25138,N_23519,N_24981);
or U25139 (N_25139,N_22109,N_24136);
nand U25140 (N_25140,N_22302,N_24253);
or U25141 (N_25141,N_22858,N_22441);
nor U25142 (N_25142,N_22995,N_23473);
and U25143 (N_25143,N_24700,N_21957);
and U25144 (N_25144,N_22792,N_22037);
nor U25145 (N_25145,N_22006,N_20930);
nand U25146 (N_25146,N_22498,N_24519);
or U25147 (N_25147,N_22748,N_21804);
xor U25148 (N_25148,N_22767,N_21026);
and U25149 (N_25149,N_21662,N_20591);
nand U25150 (N_25150,N_24296,N_22256);
nand U25151 (N_25151,N_24609,N_21426);
or U25152 (N_25152,N_20268,N_24666);
nor U25153 (N_25153,N_24402,N_20157);
nor U25154 (N_25154,N_20621,N_23289);
and U25155 (N_25155,N_24747,N_24690);
nand U25156 (N_25156,N_21469,N_20450);
and U25157 (N_25157,N_21556,N_21428);
or U25158 (N_25158,N_21384,N_21337);
xor U25159 (N_25159,N_20087,N_20995);
or U25160 (N_25160,N_22644,N_22320);
nor U25161 (N_25161,N_20261,N_23175);
nor U25162 (N_25162,N_23159,N_23834);
nor U25163 (N_25163,N_24919,N_21277);
nor U25164 (N_25164,N_21240,N_24156);
xnor U25165 (N_25165,N_23620,N_21635);
xor U25166 (N_25166,N_23549,N_21310);
or U25167 (N_25167,N_24261,N_21243);
and U25168 (N_25168,N_22657,N_22681);
xnor U25169 (N_25169,N_24123,N_20395);
nand U25170 (N_25170,N_20805,N_20103);
nor U25171 (N_25171,N_20224,N_23189);
or U25172 (N_25172,N_24869,N_20902);
and U25173 (N_25173,N_21933,N_22443);
nand U25174 (N_25174,N_20994,N_22797);
and U25175 (N_25175,N_24181,N_21419);
and U25176 (N_25176,N_24859,N_21809);
or U25177 (N_25177,N_20615,N_21153);
nand U25178 (N_25178,N_23214,N_20532);
nor U25179 (N_25179,N_23564,N_22961);
or U25180 (N_25180,N_22964,N_21772);
and U25181 (N_25181,N_20199,N_24221);
and U25182 (N_25182,N_23625,N_21056);
xnor U25183 (N_25183,N_23663,N_20243);
nor U25184 (N_25184,N_21927,N_23601);
nor U25185 (N_25185,N_20673,N_20424);
and U25186 (N_25186,N_22972,N_24984);
and U25187 (N_25187,N_23317,N_20874);
or U25188 (N_25188,N_23298,N_20712);
and U25189 (N_25189,N_24497,N_22830);
or U25190 (N_25190,N_20381,N_21914);
and U25191 (N_25191,N_24496,N_24349);
or U25192 (N_25192,N_21767,N_20038);
nor U25193 (N_25193,N_23124,N_24738);
nand U25194 (N_25194,N_23980,N_20740);
nand U25195 (N_25195,N_23059,N_21568);
nor U25196 (N_25196,N_24733,N_20309);
nor U25197 (N_25197,N_22705,N_21269);
nor U25198 (N_25198,N_23443,N_20116);
nand U25199 (N_25199,N_21615,N_23810);
nor U25200 (N_25200,N_22516,N_24380);
or U25201 (N_25201,N_22870,N_20329);
and U25202 (N_25202,N_22586,N_21923);
or U25203 (N_25203,N_20139,N_24427);
nor U25204 (N_25204,N_21038,N_21467);
and U25205 (N_25205,N_24202,N_24663);
nand U25206 (N_25206,N_24595,N_24748);
and U25207 (N_25207,N_22221,N_23696);
xor U25208 (N_25208,N_23243,N_21438);
nand U25209 (N_25209,N_20561,N_21155);
xor U25210 (N_25210,N_21793,N_20614);
nor U25211 (N_25211,N_24614,N_22808);
and U25212 (N_25212,N_23452,N_20431);
nor U25213 (N_25213,N_21339,N_22423);
nor U25214 (N_25214,N_23596,N_21612);
nand U25215 (N_25215,N_21184,N_20603);
nor U25216 (N_25216,N_24072,N_20684);
and U25217 (N_25217,N_21319,N_22341);
nand U25218 (N_25218,N_22154,N_21255);
or U25219 (N_25219,N_22673,N_20314);
or U25220 (N_25220,N_21349,N_24518);
and U25221 (N_25221,N_24036,N_23691);
nand U25222 (N_25222,N_23567,N_21641);
or U25223 (N_25223,N_24035,N_20828);
and U25224 (N_25224,N_21374,N_20373);
or U25225 (N_25225,N_21219,N_20034);
or U25226 (N_25226,N_23019,N_22587);
xor U25227 (N_25227,N_21227,N_24982);
and U25228 (N_25228,N_22346,N_22655);
and U25229 (N_25229,N_20773,N_23474);
or U25230 (N_25230,N_22746,N_23460);
nand U25231 (N_25231,N_22736,N_23285);
or U25232 (N_25232,N_21258,N_20337);
nor U25233 (N_25233,N_20839,N_21817);
nor U25234 (N_25234,N_24359,N_21395);
or U25235 (N_25235,N_22652,N_20600);
nand U25236 (N_25236,N_23013,N_20079);
nand U25237 (N_25237,N_20935,N_23162);
and U25238 (N_25238,N_21504,N_23351);
and U25239 (N_25239,N_24148,N_21529);
and U25240 (N_25240,N_22955,N_24693);
nor U25241 (N_25241,N_20411,N_22740);
and U25242 (N_25242,N_21758,N_24922);
xnor U25243 (N_25243,N_20412,N_21328);
nor U25244 (N_25244,N_22847,N_20407);
and U25245 (N_25245,N_21937,N_20924);
or U25246 (N_25246,N_21168,N_21416);
nor U25247 (N_25247,N_24712,N_23263);
nor U25248 (N_25248,N_23377,N_20587);
or U25249 (N_25249,N_22712,N_23830);
nand U25250 (N_25250,N_20187,N_22476);
nor U25251 (N_25251,N_21808,N_20915);
and U25252 (N_25252,N_20408,N_24033);
and U25253 (N_25253,N_22578,N_23328);
nor U25254 (N_25254,N_22464,N_20612);
or U25255 (N_25255,N_23442,N_22217);
or U25256 (N_25256,N_21317,N_22071);
nand U25257 (N_25257,N_22172,N_21502);
xor U25258 (N_25258,N_23606,N_23276);
nor U25259 (N_25259,N_20521,N_21062);
or U25260 (N_25260,N_20182,N_20723);
or U25261 (N_25261,N_24127,N_21108);
or U25262 (N_25262,N_24097,N_20732);
nand U25263 (N_25263,N_24746,N_23015);
and U25264 (N_25264,N_21208,N_23146);
and U25265 (N_25265,N_24223,N_24684);
nor U25266 (N_25266,N_20791,N_21813);
nand U25267 (N_25267,N_22776,N_22735);
and U25268 (N_25268,N_22110,N_21324);
and U25269 (N_25269,N_22305,N_21949);
nor U25270 (N_25270,N_20398,N_20808);
and U25271 (N_25271,N_22835,N_23914);
nor U25272 (N_25272,N_22707,N_23267);
and U25273 (N_25273,N_22160,N_20331);
nand U25274 (N_25274,N_20807,N_23427);
nand U25275 (N_25275,N_20447,N_24927);
xnor U25276 (N_25276,N_21883,N_23381);
or U25277 (N_25277,N_22621,N_23270);
or U25278 (N_25278,N_23388,N_23048);
nor U25279 (N_25279,N_24342,N_22422);
nor U25280 (N_25280,N_20810,N_22488);
xor U25281 (N_25281,N_23988,N_23154);
or U25282 (N_25282,N_21856,N_24087);
or U25283 (N_25283,N_24037,N_24424);
and U25284 (N_25284,N_23086,N_21194);
nand U25285 (N_25285,N_20517,N_24725);
nand U25286 (N_25286,N_21474,N_20346);
or U25287 (N_25287,N_21186,N_23805);
or U25288 (N_25288,N_24163,N_22946);
nor U25289 (N_25289,N_24379,N_20066);
and U25290 (N_25290,N_21241,N_22169);
nand U25291 (N_25291,N_21990,N_22080);
or U25292 (N_25292,N_20129,N_22140);
nor U25293 (N_25293,N_20633,N_24109);
or U25294 (N_25294,N_21228,N_24893);
nand U25295 (N_25295,N_22349,N_24479);
nor U25296 (N_25296,N_24405,N_23734);
and U25297 (N_25297,N_23424,N_23612);
nor U25298 (N_25298,N_21961,N_23624);
and U25299 (N_25299,N_24555,N_20772);
and U25300 (N_25300,N_20235,N_22090);
or U25301 (N_25301,N_21664,N_24288);
nand U25302 (N_25302,N_20648,N_21563);
nor U25303 (N_25303,N_24207,N_21489);
nor U25304 (N_25304,N_23425,N_23778);
nand U25305 (N_25305,N_22882,N_24147);
or U25306 (N_25306,N_20288,N_20365);
nor U25307 (N_25307,N_24762,N_21123);
nand U25308 (N_25308,N_24432,N_23562);
or U25309 (N_25309,N_20503,N_24940);
or U25310 (N_25310,N_20165,N_22375);
xor U25311 (N_25311,N_20231,N_24088);
nor U25312 (N_25312,N_23065,N_21652);
and U25313 (N_25313,N_21202,N_21908);
and U25314 (N_25314,N_22251,N_23171);
nor U25315 (N_25315,N_20246,N_24007);
and U25316 (N_25316,N_24309,N_24648);
or U25317 (N_25317,N_21072,N_23730);
nand U25318 (N_25318,N_21539,N_22437);
and U25319 (N_25319,N_20506,N_24611);
nor U25320 (N_25320,N_22785,N_24115);
nor U25321 (N_25321,N_23126,N_24294);
and U25322 (N_25322,N_24326,N_20977);
and U25323 (N_25323,N_20778,N_20100);
or U25324 (N_25324,N_21475,N_22891);
or U25325 (N_25325,N_23650,N_21737);
nor U25326 (N_25326,N_23828,N_21389);
xor U25327 (N_25327,N_20885,N_22590);
and U25328 (N_25328,N_24247,N_23832);
nor U25329 (N_25329,N_22252,N_24935);
xnor U25330 (N_25330,N_20043,N_23613);
xor U25331 (N_25331,N_21207,N_24742);
nor U25332 (N_25332,N_22824,N_22149);
or U25333 (N_25333,N_22128,N_21769);
nor U25334 (N_25334,N_20735,N_24038);
nand U25335 (N_25335,N_22348,N_23658);
nor U25336 (N_25336,N_23618,N_21846);
and U25337 (N_25337,N_23708,N_23397);
xor U25338 (N_25338,N_24104,N_22241);
nand U25339 (N_25339,N_23698,N_24418);
and U25340 (N_25340,N_24540,N_24344);
nand U25341 (N_25341,N_24477,N_21100);
and U25342 (N_25342,N_22025,N_20641);
or U25343 (N_25343,N_22095,N_23026);
or U25344 (N_25344,N_24287,N_21367);
and U25345 (N_25345,N_21146,N_22878);
and U25346 (N_25346,N_21181,N_23716);
nor U25347 (N_25347,N_21133,N_20652);
and U25348 (N_25348,N_21402,N_24487);
nand U25349 (N_25349,N_22087,N_21642);
nor U25350 (N_25350,N_20923,N_20213);
nor U25351 (N_25351,N_21122,N_20104);
nand U25352 (N_25352,N_23761,N_22021);
or U25353 (N_25353,N_20463,N_20527);
or U25354 (N_25354,N_22816,N_24063);
and U25355 (N_25355,N_23306,N_23616);
or U25356 (N_25356,N_22299,N_23637);
nand U25357 (N_25357,N_21648,N_22286);
and U25358 (N_25358,N_21580,N_20343);
and U25359 (N_25359,N_20916,N_22888);
or U25360 (N_25360,N_20031,N_24401);
nor U25361 (N_25361,N_21350,N_20004);
nor U25362 (N_25362,N_23705,N_21040);
and U25363 (N_25363,N_21482,N_21401);
nor U25364 (N_25364,N_20635,N_23565);
and U25365 (N_25365,N_23391,N_22611);
nor U25366 (N_25366,N_24913,N_23378);
or U25367 (N_25367,N_22990,N_22383);
or U25368 (N_25368,N_24234,N_21506);
and U25369 (N_25369,N_21454,N_22849);
and U25370 (N_25370,N_20596,N_24577);
xor U25371 (N_25371,N_20921,N_21882);
and U25372 (N_25372,N_22868,N_20550);
nand U25373 (N_25373,N_24924,N_23749);
or U25374 (N_25374,N_22718,N_22190);
or U25375 (N_25375,N_23887,N_21880);
nor U25376 (N_25376,N_24850,N_21916);
and U25377 (N_25377,N_24681,N_21084);
nor U25378 (N_25378,N_22728,N_22739);
or U25379 (N_25379,N_21494,N_23063);
nand U25380 (N_25380,N_24495,N_20519);
nor U25381 (N_25381,N_23385,N_23233);
and U25382 (N_25382,N_22704,N_22379);
xnor U25383 (N_25383,N_20294,N_20300);
nor U25384 (N_25384,N_23027,N_22362);
nand U25385 (N_25385,N_24056,N_21444);
and U25386 (N_25386,N_20114,N_23354);
xnor U25387 (N_25387,N_22525,N_22207);
xor U25388 (N_25388,N_22084,N_21985);
xor U25389 (N_25389,N_22073,N_20420);
or U25390 (N_25390,N_20686,N_24709);
or U25391 (N_25391,N_21720,N_20049);
nor U25392 (N_25392,N_23795,N_24967);
nor U25393 (N_25393,N_20889,N_21185);
nor U25394 (N_25394,N_24120,N_23433);
nand U25395 (N_25395,N_22001,N_20806);
and U25396 (N_25396,N_20784,N_22651);
xor U25397 (N_25397,N_24411,N_21673);
or U25398 (N_25398,N_23219,N_20324);
nor U25399 (N_25399,N_20873,N_21744);
nor U25400 (N_25400,N_22329,N_21471);
or U25401 (N_25401,N_20443,N_21553);
and U25402 (N_25402,N_21033,N_21592);
or U25403 (N_25403,N_21131,N_23221);
or U25404 (N_25404,N_24680,N_20610);
nor U25405 (N_25405,N_20241,N_24568);
nand U25406 (N_25406,N_20616,N_20055);
or U25407 (N_25407,N_24366,N_21815);
and U25408 (N_25408,N_22642,N_24830);
nand U25409 (N_25409,N_20690,N_20291);
xnor U25410 (N_25410,N_22641,N_21997);
nand U25411 (N_25411,N_22243,N_22226);
nor U25412 (N_25412,N_22769,N_23961);
nor U25413 (N_25413,N_20319,N_24993);
and U25414 (N_25414,N_21248,N_22238);
nand U25415 (N_25415,N_23509,N_21795);
and U25416 (N_25416,N_21632,N_22445);
xnor U25417 (N_25417,N_21544,N_23569);
nand U25418 (N_25418,N_24831,N_22577);
and U25419 (N_25419,N_21654,N_20265);
nor U25420 (N_25420,N_21360,N_21728);
nand U25421 (N_25421,N_21658,N_23321);
nand U25422 (N_25422,N_20866,N_24741);
and U25423 (N_25423,N_21457,N_23692);
or U25424 (N_25424,N_22871,N_24516);
xor U25425 (N_25425,N_20894,N_22715);
and U25426 (N_25426,N_24900,N_21311);
nor U25427 (N_25427,N_21427,N_21015);
nand U25428 (N_25428,N_24244,N_21296);
and U25429 (N_25429,N_20042,N_20811);
or U25430 (N_25430,N_23318,N_24917);
nor U25431 (N_25431,N_24091,N_24541);
nor U25432 (N_25432,N_23040,N_23829);
or U25433 (N_25433,N_21724,N_20177);
nand U25434 (N_25434,N_23602,N_20283);
or U25435 (N_25435,N_20298,N_20818);
nor U25436 (N_25436,N_20709,N_24605);
or U25437 (N_25437,N_23598,N_22957);
nand U25438 (N_25438,N_23685,N_20642);
nor U25439 (N_25439,N_24006,N_23762);
nand U25440 (N_25440,N_24812,N_22047);
or U25441 (N_25441,N_23858,N_23312);
and U25442 (N_25442,N_21118,N_21137);
and U25443 (N_25443,N_23607,N_20626);
nand U25444 (N_25444,N_23502,N_22706);
and U25445 (N_25445,N_23884,N_21729);
xor U25446 (N_25446,N_23599,N_21892);
and U25447 (N_25447,N_23195,N_21942);
nor U25448 (N_25448,N_24795,N_20128);
nor U25449 (N_25449,N_24082,N_21578);
nor U25450 (N_25450,N_20619,N_23181);
nor U25451 (N_25451,N_23468,N_21530);
or U25452 (N_25452,N_21775,N_20530);
or U25453 (N_25453,N_24528,N_23809);
or U25454 (N_25454,N_20295,N_22598);
nor U25455 (N_25455,N_21045,N_23967);
nand U25456 (N_25456,N_22877,N_24551);
nand U25457 (N_25457,N_24407,N_23989);
nand U25458 (N_25458,N_23430,N_23784);
xor U25459 (N_25459,N_22316,N_20487);
or U25460 (N_25460,N_22330,N_21749);
xor U25461 (N_25461,N_20077,N_21235);
nor U25462 (N_25462,N_23669,N_23710);
nor U25463 (N_25463,N_23205,N_22895);
or U25464 (N_25464,N_23493,N_21125);
nand U25465 (N_25465,N_21060,N_21661);
and U25466 (N_25466,N_21517,N_23986);
nand U25467 (N_25467,N_24469,N_24399);
and U25468 (N_25468,N_23087,N_23255);
or U25469 (N_25469,N_22513,N_22393);
and U25470 (N_25470,N_23489,N_20414);
nand U25471 (N_25471,N_20097,N_24852);
or U25472 (N_25472,N_24289,N_23053);
and U25473 (N_25473,N_23467,N_20991);
nand U25474 (N_25474,N_21564,N_23186);
nand U25475 (N_25475,N_24675,N_20001);
nand U25476 (N_25476,N_21831,N_23837);
nor U25477 (N_25477,N_21779,N_23970);
nor U25478 (N_25478,N_22993,N_21762);
nand U25479 (N_25479,N_20460,N_24530);
nand U25480 (N_25480,N_24703,N_24849);
nand U25481 (N_25481,N_24620,N_22550);
and U25482 (N_25482,N_21915,N_21332);
nand U25483 (N_25483,N_20687,N_20470);
nor U25484 (N_25484,N_24635,N_23548);
and U25485 (N_25485,N_21009,N_23158);
nand U25486 (N_25486,N_23996,N_21187);
nand U25487 (N_25487,N_24837,N_21596);
nand U25488 (N_25488,N_21799,N_22510);
and U25489 (N_25489,N_24396,N_22494);
nor U25490 (N_25490,N_23077,N_21932);
nand U25491 (N_25491,N_21910,N_24714);
and U25492 (N_25492,N_24552,N_23251);
nand U25493 (N_25493,N_22319,N_24706);
nor U25494 (N_25494,N_22357,N_22898);
xnor U25495 (N_25495,N_22480,N_21096);
nand U25496 (N_25496,N_22732,N_21850);
xor U25497 (N_25497,N_24385,N_20590);
nand U25498 (N_25498,N_22079,N_21404);
nand U25499 (N_25499,N_23016,N_20860);
nor U25500 (N_25500,N_21928,N_20084);
nor U25501 (N_25501,N_21399,N_24892);
nand U25502 (N_25502,N_20744,N_24138);
and U25503 (N_25503,N_24929,N_22798);
and U25504 (N_25504,N_21342,N_23885);
nand U25505 (N_25505,N_24307,N_22976);
nor U25506 (N_25506,N_20392,N_20434);
nor U25507 (N_25507,N_24556,N_23177);
and U25508 (N_25508,N_22973,N_20110);
or U25509 (N_25509,N_23242,N_23123);
nand U25510 (N_25510,N_20937,N_22322);
nand U25511 (N_25511,N_20912,N_22093);
or U25512 (N_25512,N_22248,N_23098);
nand U25513 (N_25513,N_21086,N_20827);
nor U25514 (N_25514,N_24636,N_23119);
nor U25515 (N_25515,N_24691,N_20504);
and U25516 (N_25516,N_22920,N_22827);
and U25517 (N_25517,N_24618,N_22103);
or U25518 (N_25518,N_20770,N_21599);
and U25519 (N_25519,N_20852,N_23568);
and U25520 (N_25520,N_22406,N_24034);
and U25521 (N_25521,N_24464,N_24806);
nand U25522 (N_25522,N_20763,N_20625);
nand U25523 (N_25523,N_23928,N_24529);
and U25524 (N_25524,N_23253,N_24079);
xnor U25525 (N_25525,N_20260,N_24626);
nor U25526 (N_25526,N_23232,N_23372);
and U25527 (N_25527,N_21770,N_21852);
or U25528 (N_25528,N_20969,N_24510);
nor U25529 (N_25529,N_24783,N_20698);
xor U25530 (N_25530,N_23680,N_22546);
nand U25531 (N_25531,N_22165,N_22937);
nand U25532 (N_25532,N_21693,N_21351);
or U25533 (N_25533,N_22690,N_24745);
nor U25534 (N_25534,N_22325,N_21493);
and U25535 (N_25535,N_20180,N_20068);
or U25536 (N_25536,N_22520,N_20002);
and U25537 (N_25537,N_24018,N_20883);
or U25538 (N_25538,N_24149,N_22363);
and U25539 (N_25539,N_22649,N_22684);
xnor U25540 (N_25540,N_20754,N_22168);
and U25541 (N_25541,N_23426,N_21858);
and U25542 (N_25542,N_20750,N_24237);
or U25543 (N_25543,N_24085,N_24936);
nand U25544 (N_25544,N_20438,N_24751);
xor U25545 (N_25545,N_23479,N_24209);
or U25546 (N_25546,N_22428,N_22107);
and U25547 (N_25547,N_23717,N_20578);
and U25548 (N_25548,N_24398,N_21409);
nand U25549 (N_25549,N_24754,N_23133);
nor U25550 (N_25550,N_24959,N_20624);
and U25551 (N_25551,N_22822,N_23169);
and U25552 (N_25552,N_23935,N_23649);
nor U25553 (N_25553,N_22211,N_24302);
nor U25554 (N_25554,N_24823,N_24224);
and U25555 (N_25555,N_20210,N_22009);
nor U25556 (N_25556,N_21655,N_20474);
or U25557 (N_25557,N_21156,N_20716);
and U25558 (N_25558,N_24301,N_21668);
nand U25559 (N_25559,N_24769,N_21798);
or U25560 (N_25560,N_23752,N_23997);
and U25561 (N_25561,N_20918,N_23861);
nor U25562 (N_25562,N_23777,N_22790);
nand U25563 (N_25563,N_20078,N_21854);
and U25564 (N_25564,N_23787,N_20219);
and U25565 (N_25565,N_23373,N_24065);
nand U25566 (N_25566,N_20321,N_22250);
or U25567 (N_25567,N_24628,N_22522);
nand U25568 (N_25568,N_22795,N_21690);
and U25569 (N_25569,N_23954,N_21176);
xor U25570 (N_25570,N_23327,N_24585);
and U25571 (N_25571,N_24208,N_20217);
nand U25572 (N_25572,N_20236,N_22949);
xor U25573 (N_25573,N_24752,N_24832);
or U25574 (N_25574,N_24559,N_20914);
nor U25575 (N_25575,N_22469,N_21049);
nand U25576 (N_25576,N_21315,N_22386);
and U25577 (N_25577,N_20820,N_24954);
and U25578 (N_25578,N_23552,N_22179);
or U25579 (N_25579,N_20130,N_23014);
xnor U25580 (N_25580,N_21242,N_23871);
or U25581 (N_25581,N_23101,N_23486);
xor U25582 (N_25582,N_20513,N_23316);
and U25583 (N_25583,N_22019,N_21862);
and U25584 (N_25584,N_23732,N_23409);
or U25585 (N_25585,N_24019,N_20029);
nor U25586 (N_25586,N_20326,N_20394);
nand U25587 (N_25587,N_23750,N_20881);
or U25588 (N_25588,N_23690,N_22982);
nand U25589 (N_25589,N_22300,N_20205);
and U25590 (N_25590,N_21111,N_24368);
or U25591 (N_25591,N_24829,N_20476);
or U25592 (N_25592,N_22733,N_24484);
xnor U25593 (N_25593,N_24130,N_22876);
or U25594 (N_25594,N_23309,N_24269);
nor U25595 (N_25595,N_23768,N_23672);
and U25596 (N_25596,N_20785,N_21414);
nor U25597 (N_25597,N_21180,N_21260);
and U25598 (N_25598,N_23942,N_20727);
and U25599 (N_25599,N_23540,N_24860);
nor U25600 (N_25600,N_23458,N_24321);
and U25601 (N_25601,N_23659,N_22097);
nor U25602 (N_25602,N_23864,N_23157);
nor U25603 (N_25603,N_22963,N_21757);
nor U25604 (N_25604,N_20378,N_23404);
or U25605 (N_25605,N_23006,N_20948);
or U25606 (N_25606,N_22403,N_22455);
or U25607 (N_25607,N_23539,N_22032);
and U25608 (N_25608,N_23591,N_22482);
nor U25609 (N_25609,N_20299,N_24792);
nor U25610 (N_25610,N_23993,N_22442);
or U25611 (N_25611,N_23278,N_22511);
nor U25612 (N_25612,N_23588,N_24946);
nand U25613 (N_25613,N_21640,N_24844);
or U25614 (N_25614,N_22101,N_20620);
and U25615 (N_25615,N_24841,N_21273);
nor U25616 (N_25616,N_22677,N_21263);
or U25617 (N_25617,N_21116,N_21816);
nand U25618 (N_25618,N_23633,N_24020);
xnor U25619 (N_25619,N_20908,N_24674);
nand U25620 (N_25620,N_21095,N_20234);
nor U25621 (N_25621,N_21948,N_20544);
or U25622 (N_25622,N_21630,N_21088);
or U25623 (N_25623,N_20759,N_22624);
or U25624 (N_25624,N_23689,N_20528);
or U25625 (N_25625,N_24513,N_23394);
nand U25626 (N_25626,N_24679,N_21800);
nor U25627 (N_25627,N_24928,N_22879);
xor U25628 (N_25628,N_23084,N_20695);
or U25629 (N_25629,N_22317,N_20109);
or U25630 (N_25630,N_21282,N_24579);
nor U25631 (N_25631,N_24212,N_21174);
and U25632 (N_25632,N_21712,N_21909);
or U25633 (N_25633,N_21473,N_24951);
or U25634 (N_25634,N_22533,N_23824);
and U25635 (N_25635,N_24451,N_21863);
and U25636 (N_25636,N_20947,N_24651);
xor U25637 (N_25637,N_20765,N_22236);
xnor U25638 (N_25638,N_24724,N_20218);
and U25639 (N_25639,N_21004,N_20756);
nand U25640 (N_25640,N_23083,N_20580);
nand U25641 (N_25641,N_20153,N_20940);
or U25642 (N_25642,N_22030,N_21656);
xor U25643 (N_25643,N_22031,N_21000);
nand U25644 (N_25644,N_23594,N_24952);
and U25645 (N_25645,N_24966,N_24406);
nand U25646 (N_25646,N_20382,N_24732);
nand U25647 (N_25647,N_20311,N_23148);
nor U25648 (N_25648,N_22421,N_20493);
or U25649 (N_25649,N_22070,N_21205);
nor U25650 (N_25650,N_22671,N_24116);
nor U25651 (N_25651,N_22910,N_23456);
or U25652 (N_25652,N_24105,N_20357);
nor U25653 (N_25653,N_24511,N_23376);
nand U25654 (N_25654,N_21193,N_23783);
or U25655 (N_25655,N_22999,N_22223);
nand U25656 (N_25656,N_23816,N_21002);
and U25657 (N_25657,N_21306,N_20448);
nor U25658 (N_25658,N_20010,N_20602);
nand U25659 (N_25659,N_21974,N_24835);
and U25660 (N_25660,N_22082,N_20983);
or U25661 (N_25661,N_20980,N_22481);
or U25662 (N_25662,N_24676,N_22612);
nor U25663 (N_25663,N_23505,N_23034);
and U25664 (N_25664,N_22777,N_22678);
or U25665 (N_25665,N_22661,N_21265);
and U25666 (N_25666,N_23144,N_22399);
and U25667 (N_25667,N_20046,N_24332);
nor U25668 (N_25668,N_21281,N_23758);
and U25669 (N_25669,N_21216,N_24560);
nor U25670 (N_25670,N_20409,N_23976);
or U25671 (N_25671,N_24589,N_23640);
or U25672 (N_25672,N_20330,N_22108);
nand U25673 (N_25673,N_23706,N_24855);
and U25674 (N_25674,N_22013,N_22143);
nand U25675 (N_25675,N_22860,N_23981);
nand U25676 (N_25676,N_24121,N_23851);
or U25677 (N_25677,N_23512,N_22334);
xor U25678 (N_25678,N_20606,N_20896);
or U25679 (N_25679,N_20747,N_20095);
or U25680 (N_25680,N_22237,N_23417);
and U25681 (N_25681,N_22397,N_23590);
nor U25682 (N_25682,N_24668,N_22089);
or U25683 (N_25683,N_22622,N_23449);
or U25684 (N_25684,N_22425,N_22212);
or U25685 (N_25685,N_21099,N_20385);
nor U25686 (N_25686,N_20541,N_20531);
and U25687 (N_25687,N_22602,N_20170);
and U25688 (N_25688,N_22862,N_20720);
nor U25689 (N_25689,N_22763,N_20836);
nor U25690 (N_25690,N_22091,N_20882);
and U25691 (N_25691,N_21867,N_23261);
nand U25692 (N_25692,N_22630,N_22438);
or U25693 (N_25693,N_24334,N_23919);
or U25694 (N_25694,N_22038,N_24764);
xnor U25695 (N_25695,N_24319,N_20134);
nor U25696 (N_25696,N_21344,N_21812);
or U25697 (N_25697,N_22479,N_21996);
nor U25698 (N_25698,N_24171,N_23122);
xnor U25699 (N_25699,N_22873,N_21629);
nand U25700 (N_25700,N_20691,N_22628);
and U25701 (N_25701,N_22446,N_24488);
nand U25702 (N_25702,N_24089,N_22818);
nand U25703 (N_25703,N_22509,N_21534);
nor U25704 (N_25704,N_23770,N_23078);
xnor U25705 (N_25705,N_21408,N_22829);
and U25706 (N_25706,N_21618,N_24439);
xnor U25707 (N_25707,N_23866,N_24017);
or U25708 (N_25708,N_22921,N_24838);
nand U25709 (N_25709,N_20847,N_22680);
xor U25710 (N_25710,N_21784,N_22112);
nand U25711 (N_25711,N_24544,N_21291);
and U25712 (N_25712,N_22666,N_22720);
xnor U25713 (N_25713,N_22115,N_24200);
nand U25714 (N_25714,N_24872,N_22174);
xor U25715 (N_25715,N_21598,N_21508);
nand U25716 (N_25716,N_22384,N_23024);
nor U25717 (N_25717,N_24866,N_23904);
nor U25718 (N_25718,N_21220,N_21610);
nor U25719 (N_25719,N_21390,N_23438);
or U25720 (N_25720,N_24027,N_22373);
nand U25721 (N_25721,N_22692,N_22536);
or U25722 (N_25722,N_24341,N_24267);
or U25723 (N_25723,N_20814,N_20467);
nand U25724 (N_25724,N_22929,N_24028);
nor U25725 (N_25725,N_20796,N_20963);
nand U25726 (N_25726,N_21604,N_22703);
and U25727 (N_25727,N_22756,N_21076);
nand U25728 (N_25728,N_22535,N_22597);
nand U25729 (N_25729,N_23491,N_24455);
nor U25730 (N_25730,N_24145,N_21925);
nor U25731 (N_25731,N_20211,N_23344);
and U25732 (N_25732,N_22303,N_21577);
or U25733 (N_25733,N_22119,N_24820);
nor U25734 (N_25734,N_23850,N_22534);
or U25735 (N_25735,N_21393,N_22004);
or U25736 (N_25736,N_20047,N_23281);
nand U25737 (N_25737,N_21366,N_23497);
and U25738 (N_25738,N_22005,N_20008);
and U25739 (N_25739,N_24374,N_23297);
or U25740 (N_25740,N_24607,N_24062);
and U25741 (N_25741,N_22407,N_23746);
nand U25742 (N_25742,N_24239,N_23506);
or U25743 (N_25743,N_24785,N_21678);
nor U25744 (N_25744,N_24876,N_22826);
and U25745 (N_25745,N_22335,N_24367);
nand U25746 (N_25746,N_22246,N_22321);
and U25747 (N_25747,N_24167,N_20018);
and U25748 (N_25748,N_24233,N_22750);
and U25749 (N_25749,N_23005,N_23675);
or U25750 (N_25750,N_21098,N_20322);
nand U25751 (N_25751,N_20107,N_20745);
and U25752 (N_25752,N_22981,N_20567);
and U25753 (N_25753,N_20439,N_23760);
nor U25754 (N_25754,N_24969,N_20341);
or U25755 (N_25755,N_21602,N_24802);
and U25756 (N_25756,N_22259,N_21230);
and U25757 (N_25757,N_22347,N_23729);
nand U25758 (N_25758,N_23155,N_24539);
or U25759 (N_25759,N_20477,N_20340);
nor U25760 (N_25760,N_23170,N_21157);
or U25761 (N_25761,N_24462,N_23959);
nand U25762 (N_25762,N_22184,N_24029);
nand U25763 (N_25763,N_24482,N_24658);
or U25764 (N_25764,N_20987,N_23559);
or U25765 (N_25765,N_20768,N_23054);
or U25766 (N_25766,N_20427,N_20509);
xnor U25767 (N_25767,N_20359,N_23141);
and U25768 (N_25768,N_20545,N_22486);
nand U25769 (N_25769,N_23962,N_24220);
nor U25770 (N_25770,N_23990,N_24111);
nor U25771 (N_25771,N_21509,N_21703);
or U25772 (N_25772,N_24996,N_23819);
nor U25773 (N_25773,N_23523,N_22272);
and U25774 (N_25774,N_22257,N_22807);
and U25775 (N_25775,N_22245,N_21851);
nor U25776 (N_25776,N_24734,N_20195);
nand U25777 (N_25777,N_22210,N_22872);
or U25778 (N_25778,N_23128,N_21431);
or U25779 (N_25779,N_23994,N_22600);
and U25780 (N_25780,N_24814,N_24565);
nor U25781 (N_25781,N_24066,N_20864);
and U25782 (N_25782,N_20953,N_24483);
or U25783 (N_25783,N_20336,N_22517);
or U25784 (N_25784,N_20658,N_24723);
and U25785 (N_25785,N_20629,N_24578);
nor U25786 (N_25786,N_21576,N_22960);
nor U25787 (N_25787,N_20417,N_23765);
nand U25788 (N_25788,N_22206,N_24493);
nand U25789 (N_25789,N_20413,N_20830);
nor U25790 (N_25790,N_20333,N_22701);
and U25791 (N_25791,N_22966,N_23030);
or U25792 (N_25792,N_23515,N_24246);
and U25793 (N_25793,N_21837,N_20316);
and U25794 (N_25794,N_20533,N_21689);
or U25795 (N_25795,N_23849,N_21866);
and U25796 (N_25796,N_23687,N_20910);
and U25797 (N_25797,N_23507,N_20287);
nor U25798 (N_25798,N_20304,N_23872);
nor U25799 (N_25799,N_24131,N_21680);
nand U25800 (N_25800,N_21405,N_21290);
or U25801 (N_25801,N_22631,N_21058);
and U25802 (N_25802,N_22114,N_20325);
and U25803 (N_25803,N_21583,N_22368);
nor U25804 (N_25804,N_22845,N_21746);
nand U25805 (N_25805,N_24420,N_23204);
nor U25806 (N_25806,N_21543,N_24584);
or U25807 (N_25807,N_22351,N_21940);
or U25808 (N_25808,N_24177,N_20108);
or U25809 (N_25809,N_23049,N_20936);
and U25810 (N_25810,N_22572,N_22914);
xnor U25811 (N_25811,N_22825,N_23190);
nand U25812 (N_25812,N_22358,N_23067);
nand U25813 (N_25813,N_20905,N_23755);
or U25814 (N_25814,N_20518,N_20981);
nor U25815 (N_25815,N_21309,N_20693);
and U25816 (N_25816,N_23524,N_20466);
or U25817 (N_25817,N_23723,N_20683);
or U25818 (N_25818,N_21483,N_21585);
nand U25819 (N_25819,N_21570,N_21537);
or U25820 (N_25820,N_24517,N_22146);
nand U25821 (N_25821,N_22267,N_22216);
and U25822 (N_25822,N_21130,N_21177);
or U25823 (N_25823,N_23332,N_24444);
nand U25824 (N_25824,N_23905,N_20022);
or U25825 (N_25825,N_23982,N_23844);
nor U25826 (N_25826,N_21254,N_22002);
nand U25827 (N_25827,N_21379,N_23238);
and U25828 (N_25828,N_22892,N_22225);
nor U25829 (N_25829,N_20722,N_23737);
and U25830 (N_25830,N_23282,N_24938);
nand U25831 (N_25831,N_24090,N_20971);
and U25832 (N_25832,N_24948,N_24522);
or U25833 (N_25833,N_22275,N_23945);
and U25834 (N_25834,N_20557,N_23292);
nor U25835 (N_25835,N_24077,N_24475);
nand U25836 (N_25836,N_20033,N_20227);
nand U25837 (N_25837,N_22398,N_24662);
and U25838 (N_25838,N_20208,N_20592);
or U25839 (N_25839,N_20375,N_21796);
xor U25840 (N_25840,N_21605,N_22337);
nand U25841 (N_25841,N_24150,N_23407);
xor U25842 (N_25842,N_20571,N_20755);
nor U25843 (N_25843,N_20582,N_24458);
xnor U25844 (N_25844,N_22167,N_24998);
nor U25845 (N_25845,N_24886,N_21497);
xor U25846 (N_25846,N_20682,N_20258);
nor U25847 (N_25847,N_24457,N_22197);
and U25848 (N_25848,N_24526,N_20402);
and U25849 (N_25849,N_24902,N_23047);
xor U25850 (N_25850,N_22215,N_22907);
nand U25851 (N_25851,N_23504,N_23697);
nor U25852 (N_25852,N_23411,N_21455);
xor U25853 (N_25853,N_22085,N_21077);
nand U25854 (N_25854,N_24240,N_24481);
nand U25855 (N_25855,N_20577,N_22000);
and U25856 (N_25856,N_22185,N_22060);
xor U25857 (N_25857,N_20158,N_24887);
or U25858 (N_25858,N_23446,N_24161);
and U25859 (N_25859,N_22113,N_23638);
and U25860 (N_25860,N_20351,N_21357);
and U25861 (N_25861,N_22566,N_21714);
xor U25862 (N_25862,N_20415,N_20511);
or U25863 (N_25863,N_23808,N_24813);
nor U25864 (N_25864,N_22601,N_21519);
and U25865 (N_25865,N_22931,N_22637);
nand U25866 (N_25866,N_24203,N_24112);
nand U25867 (N_25867,N_24610,N_20636);
and U25868 (N_25868,N_20052,N_23574);
and U25869 (N_25869,N_23266,N_24179);
nand U25870 (N_25870,N_22388,N_23646);
or U25871 (N_25871,N_22199,N_20160);
nand U25872 (N_25872,N_20144,N_23051);
or U25873 (N_25873,N_20696,N_23930);
nor U25874 (N_25874,N_22283,N_23139);
nand U25875 (N_25875,N_23066,N_21413);
or U25876 (N_25876,N_20360,N_23224);
nand U25877 (N_25877,N_23720,N_23132);
nor U25878 (N_25878,N_24615,N_24629);
nand U25879 (N_25879,N_21251,N_21447);
nand U25880 (N_25880,N_21745,N_22024);
or U25881 (N_25881,N_20581,N_24809);
and U25882 (N_25882,N_21774,N_23764);
or U25883 (N_25883,N_23499,N_21616);
nand U25884 (N_25884,N_24816,N_23642);
or U25885 (N_25885,N_23779,N_21981);
nor U25886 (N_25886,N_20076,N_21159);
nor U25887 (N_25887,N_20920,N_23657);
or U25888 (N_25888,N_22853,N_23682);
nand U25889 (N_25889,N_21562,N_20660);
nor U25890 (N_25890,N_23718,N_23902);
and U25891 (N_25891,N_23852,N_24657);
nand U25892 (N_25892,N_21304,N_22151);
and U25893 (N_25893,N_22711,N_24453);
nor U25894 (N_25894,N_21134,N_20137);
nor U25895 (N_25895,N_23152,N_20239);
and U25896 (N_25896,N_24968,N_21603);
nand U25897 (N_25897,N_21560,N_24340);
and U25898 (N_25898,N_22308,N_23644);
nand U25899 (N_25899,N_22814,N_20242);
and U25900 (N_25900,N_22779,N_20082);
nand U25901 (N_25901,N_23002,N_24934);
nor U25902 (N_25902,N_24713,N_23296);
and U25903 (N_25903,N_21288,N_22639);
nor U25904 (N_25904,N_21926,N_22571);
and U25905 (N_25905,N_21035,N_22506);
and U25906 (N_25906,N_22626,N_20540);
and U25907 (N_25907,N_20903,N_24474);
nand U25908 (N_25908,N_20627,N_23356);
xnor U25909 (N_25909,N_22953,N_21572);
and U25910 (N_25910,N_22173,N_21320);
xnor U25911 (N_25911,N_20490,N_24489);
nand U25912 (N_25912,N_22552,N_22290);
and U25913 (N_25913,N_23653,N_23215);
or U25914 (N_25914,N_21586,N_22371);
and U25915 (N_25915,N_21822,N_22277);
nor U25916 (N_25916,N_23751,N_21947);
nand U25917 (N_25917,N_22023,N_21329);
or U25918 (N_25918,N_23241,N_22133);
and U25919 (N_25919,N_21535,N_23947);
nor U25920 (N_25920,N_20962,N_22331);
nand U25921 (N_25921,N_20749,N_24382);
nand U25922 (N_25922,N_23915,N_23121);
nand U25923 (N_25923,N_20289,N_23896);
nor U25924 (N_25924,N_21900,N_22820);
nor U25925 (N_25925,N_20539,N_21365);
or U25926 (N_25926,N_22817,N_24603);
or U25927 (N_25927,N_24317,N_24804);
nor U25928 (N_25928,N_24891,N_23978);
nand U25929 (N_25929,N_24503,N_22688);
nand U25930 (N_25930,N_23035,N_20552);
nand U25931 (N_25931,N_20703,N_21433);
nand U25932 (N_25932,N_24749,N_22063);
nand U25933 (N_25933,N_21872,N_21068);
or U25934 (N_25934,N_20120,N_20943);
or U25935 (N_25935,N_20676,N_22553);
nor U25936 (N_25936,N_24506,N_20760);
or U25937 (N_25937,N_23268,N_24588);
nor U25938 (N_25938,N_22155,N_22583);
nand U25939 (N_25939,N_21781,N_24520);
nand U25940 (N_25940,N_20892,N_24005);
and U25941 (N_25941,N_20560,N_20798);
or U25942 (N_25942,N_22978,N_21129);
and U25943 (N_25943,N_23383,N_23073);
or U25944 (N_25944,N_23563,N_22344);
and U25945 (N_25945,N_21934,N_23665);
or U25946 (N_25946,N_24963,N_20194);
nor U25947 (N_25947,N_20151,N_21647);
and U25948 (N_25948,N_20284,N_22035);
nand U25949 (N_25949,N_23741,N_22361);
and U25950 (N_25950,N_20907,N_22927);
nand U25951 (N_25951,N_22055,N_23439);
nand U25952 (N_25952,N_21106,N_23008);
or U25953 (N_25953,N_24890,N_23022);
nor U25954 (N_25954,N_22717,N_21179);
nand U25955 (N_25955,N_21300,N_20534);
nor U25956 (N_25956,N_21165,N_20584);
nor U25957 (N_25957,N_24939,N_21091);
or U25958 (N_25958,N_20059,N_21743);
nor U25959 (N_25959,N_20220,N_23011);
and U25960 (N_25960,N_23300,N_23445);
nor U25961 (N_25961,N_21792,N_23820);
nand U25962 (N_25962,N_22923,N_20964);
or U25963 (N_25963,N_20307,N_23387);
nor U25964 (N_25964,N_21161,N_22254);
or U25965 (N_25965,N_20512,N_20575);
or U25966 (N_25966,N_22209,N_23249);
and U25967 (N_25967,N_24999,N_22495);
nor U25968 (N_25968,N_23088,N_23939);
and U25969 (N_25969,N_23772,N_21982);
nor U25970 (N_25970,N_24904,N_20526);
nor U25971 (N_25971,N_24730,N_23274);
nor U25972 (N_25972,N_23586,N_24189);
nand U25973 (N_25973,N_22729,N_24377);
and U25974 (N_25974,N_23220,N_22098);
nand U25975 (N_25975,N_23330,N_20496);
or U25976 (N_25976,N_20012,N_21217);
nand U25977 (N_25977,N_21215,N_21005);
xor U25978 (N_25978,N_20070,N_20207);
and U25979 (N_25979,N_22204,N_24979);
nor U25980 (N_25980,N_23272,N_24863);
nand U25981 (N_25981,N_24361,N_22633);
xnor U25982 (N_25982,N_21238,N_21214);
nand U25983 (N_25983,N_20025,N_23286);
and U25984 (N_25984,N_21840,N_22147);
and U25985 (N_25985,N_23836,N_24569);
or U25986 (N_25986,N_20789,N_21233);
or U25987 (N_25987,N_24113,N_21257);
nand U25988 (N_25988,N_24550,N_24964);
nor U25989 (N_25989,N_22640,N_21031);
or U25990 (N_25990,N_22273,N_24972);
and U25991 (N_25991,N_20999,N_23153);
nand U25992 (N_25992,N_22230,N_20523);
nor U25993 (N_25993,N_21010,N_22340);
and U25994 (N_25994,N_20480,N_24304);
nand U25995 (N_25995,N_23614,N_24354);
nor U25996 (N_25996,N_23715,N_22507);
or U25997 (N_25997,N_23032,N_23968);
nand U25998 (N_25998,N_20481,N_20094);
nand U25999 (N_25999,N_22459,N_22288);
xor U26000 (N_26000,N_23325,N_20651);
nand U26001 (N_26001,N_21027,N_24486);
nand U26002 (N_26002,N_21638,N_23703);
and U26003 (N_26003,N_21278,N_23389);
or U26004 (N_26004,N_21929,N_23104);
and U26005 (N_26005,N_24195,N_23323);
and U26006 (N_26006,N_24756,N_21760);
and U26007 (N_26007,N_22780,N_22766);
nand U26008 (N_26008,N_21468,N_20566);
and U26009 (N_26009,N_24436,N_22696);
nor U26010 (N_26010,N_24047,N_24231);
and U26011 (N_26011,N_22069,N_23966);
and U26012 (N_26012,N_22414,N_24851);
or U26013 (N_26013,N_23420,N_24545);
xor U26014 (N_26014,N_24914,N_22328);
and U26015 (N_26015,N_23700,N_22793);
or U26016 (N_26016,N_24644,N_21039);
nor U26017 (N_26017,N_24188,N_21006);
nand U26018 (N_26018,N_23529,N_24533);
and U26019 (N_26019,N_24678,N_23531);
and U26020 (N_26020,N_23492,N_20126);
xor U26021 (N_26021,N_22909,N_23943);
nor U26022 (N_26022,N_20303,N_23382);
and U26023 (N_26023,N_21270,N_24012);
or U26024 (N_26024,N_21765,N_21145);
or U26025 (N_26025,N_22497,N_23724);
xnor U26026 (N_26026,N_20715,N_20471);
or U26027 (N_26027,N_20919,N_22989);
nor U26028 (N_26028,N_24699,N_23462);
or U26029 (N_26029,N_23950,N_20998);
nand U26030 (N_26030,N_22433,N_23604);
xnor U26031 (N_26031,N_24440,N_20949);
nand U26032 (N_26032,N_21967,N_21030);
and U26033 (N_26033,N_20403,N_21434);
and U26034 (N_26034,N_20643,N_23738);
nor U26035 (N_26035,N_24025,N_20149);
xnor U26036 (N_26036,N_23018,N_23684);
nand U26037 (N_26037,N_20733,N_23437);
nand U26038 (N_26038,N_23069,N_24977);
and U26039 (N_26039,N_24108,N_20143);
and U26040 (N_26040,N_20878,N_23535);
nand U26041 (N_26041,N_20115,N_22027);
nand U26042 (N_26042,N_21221,N_20376);
or U26043 (N_26043,N_23611,N_20266);
and U26044 (N_26044,N_21150,N_24485);
nand U26045 (N_26045,N_20380,N_21094);
nand U26046 (N_26046,N_20875,N_24023);
or U26047 (N_26047,N_21657,N_23454);
and U26048 (N_26048,N_23895,N_22549);
nor U26049 (N_26049,N_24995,N_23686);
nand U26050 (N_26050,N_21144,N_22874);
nand U26051 (N_26051,N_20668,N_24051);
nor U26052 (N_26052,N_20702,N_23271);
nor U26053 (N_26053,N_22461,N_23466);
nor U26054 (N_26054,N_24441,N_21778);
or U26055 (N_26055,N_21301,N_20654);
or U26056 (N_26056,N_24480,N_20019);
and U26057 (N_26057,N_20990,N_20520);
nor U26058 (N_26058,N_24449,N_22852);
or U26059 (N_26059,N_24688,N_23537);
nor U26060 (N_26060,N_23279,N_23333);
or U26061 (N_26061,N_23921,N_24632);
nor U26062 (N_26062,N_24308,N_24750);
and U26063 (N_26063,N_24229,N_20797);
xnor U26064 (N_26064,N_20206,N_21516);
and U26065 (N_26065,N_24898,N_21047);
or U26066 (N_26066,N_24376,N_22499);
nor U26067 (N_26067,N_22229,N_21514);
or U26068 (N_26068,N_23577,N_23440);
and U26069 (N_26069,N_22159,N_23237);
and U26070 (N_26070,N_23463,N_23358);
and U26071 (N_26071,N_20464,N_24336);
and U26072 (N_26072,N_24157,N_21975);
nor U26073 (N_26073,N_23571,N_21175);
or U26074 (N_26074,N_23825,N_21023);
xnor U26075 (N_26075,N_23522,N_20345);
and U26076 (N_26076,N_20942,N_22593);
or U26077 (N_26077,N_23583,N_22081);
nand U26078 (N_26078,N_24413,N_22634);
or U26079 (N_26079,N_24228,N_20313);
and U26080 (N_26080,N_23854,N_24270);
xnor U26081 (N_26081,N_24423,N_24442);
and U26082 (N_26082,N_21569,N_23570);
nor U26083 (N_26083,N_23149,N_23444);
nand U26084 (N_26084,N_20721,N_20292);
nor U26085 (N_26085,N_21347,N_23482);
or U26086 (N_26086,N_23192,N_23822);
xnor U26087 (N_26087,N_23436,N_21810);
or U26088 (N_26088,N_24779,N_21466);
nor U26089 (N_26089,N_23801,N_24346);
nand U26090 (N_26090,N_22323,N_23940);
or U26091 (N_26091,N_23346,N_23020);
nand U26092 (N_26092,N_22462,N_24081);
xor U26093 (N_26093,N_23818,N_22450);
or U26094 (N_26094,N_20674,N_23001);
and U26095 (N_26095,N_21597,N_22018);
and U26096 (N_26096,N_20429,N_24222);
nor U26097 (N_26097,N_23359,N_20172);
nor U26098 (N_26098,N_22514,N_21369);
or U26099 (N_26099,N_24670,N_22104);
nand U26100 (N_26100,N_22564,N_23236);
or U26101 (N_26101,N_21398,N_22489);
nor U26102 (N_26102,N_23025,N_23948);
and U26103 (N_26103,N_21950,N_22415);
nor U26104 (N_26104,N_24888,N_23260);
nand U26105 (N_26105,N_22968,N_21120);
nor U26106 (N_26106,N_20522,N_24044);
or U26107 (N_26107,N_23892,N_21397);
nor U26108 (N_26108,N_24574,N_22938);
nor U26109 (N_26109,N_22926,N_24210);
or U26110 (N_26110,N_23033,N_20812);
nor U26111 (N_26111,N_22607,N_24591);
nor U26112 (N_26112,N_22124,N_23343);
nand U26113 (N_26113,N_21430,N_20804);
nand U26114 (N_26114,N_22332,N_24466);
and U26115 (N_26115,N_23797,N_21336);
xor U26116 (N_26116,N_22806,N_20334);
nor U26117 (N_26117,N_24134,N_24291);
and U26118 (N_26118,N_21962,N_21355);
nor U26119 (N_26119,N_21001,N_21821);
and U26120 (N_26120,N_21617,N_20011);
nor U26121 (N_26121,N_20131,N_20762);
or U26122 (N_26122,N_22493,N_23566);
nand U26123 (N_26123,N_21969,N_24125);
nor U26124 (N_26124,N_20492,N_23455);
xnor U26125 (N_26125,N_21443,N_21555);
nor U26126 (N_26126,N_23342,N_20705);
or U26127 (N_26127,N_23322,N_23483);
and U26128 (N_26128,N_23911,N_21083);
xnor U26129 (N_26129,N_22467,N_22613);
or U26130 (N_26130,N_22503,N_21054);
and U26131 (N_26131,N_24937,N_23365);
nand U26132 (N_26132,N_22588,N_24083);
and U26133 (N_26133,N_24716,N_22232);
nor U26134 (N_26134,N_23095,N_21245);
nor U26135 (N_26135,N_23969,N_22447);
nor U26136 (N_26136,N_21325,N_22573);
nand U26137 (N_26137,N_21988,N_24875);
nand U26138 (N_26138,N_21521,N_21452);
and U26139 (N_26139,N_20462,N_24570);
or U26140 (N_26140,N_23244,N_21067);
nand U26141 (N_26141,N_22505,N_20397);
nand U26142 (N_26142,N_20677,N_24846);
and U26143 (N_26143,N_22689,N_22022);
and U26144 (N_26144,N_24213,N_24266);
and U26145 (N_26145,N_21613,N_24395);
and U26146 (N_26146,N_24720,N_20225);
nor U26147 (N_26147,N_22911,N_20111);
nand U26148 (N_26148,N_22697,N_20445);
nand U26149 (N_26149,N_21224,N_20605);
and U26150 (N_26150,N_24429,N_23320);
xor U26151 (N_26151,N_23127,N_22292);
or U26152 (N_26152,N_20280,N_24655);
nor U26153 (N_26153,N_21303,N_22219);
and U26154 (N_26154,N_22094,N_22676);
nor U26155 (N_26155,N_24355,N_23550);
and U26156 (N_26156,N_22887,N_20734);
or U26157 (N_26157,N_24492,N_20867);
nand U26158 (N_26158,N_24358,N_20985);
nand U26159 (N_26159,N_20886,N_22102);
nand U26160 (N_26160,N_22980,N_21832);
and U26161 (N_26161,N_23576,N_21587);
nor U26162 (N_26162,N_24215,N_24781);
or U26163 (N_26163,N_21417,N_24701);
and U26164 (N_26164,N_23475,N_23878);
nor U26165 (N_26165,N_21021,N_20593);
or U26166 (N_26166,N_22727,N_24384);
nand U26167 (N_26167,N_24983,N_24845);
nand U26168 (N_26168,N_20254,N_22743);
or U26169 (N_26169,N_22158,N_23835);
nand U26170 (N_26170,N_21448,N_24920);
or U26171 (N_26171,N_22458,N_23212);
nor U26172 (N_26172,N_23796,N_20840);
or U26173 (N_26173,N_22653,N_23245);
or U26174 (N_26174,N_22576,N_20829);
and U26175 (N_26175,N_21904,N_24042);
and U26176 (N_26176,N_20267,N_21913);
and U26177 (N_26177,N_23528,N_21188);
xor U26178 (N_26178,N_20249,N_22429);
xor U26179 (N_26179,N_21406,N_23662);
or U26180 (N_26180,N_23695,N_21773);
nand U26181 (N_26181,N_20837,N_22605);
and U26182 (N_26182,N_21044,N_22773);
and U26183 (N_26183,N_24498,N_24254);
nor U26184 (N_26184,N_21542,N_21687);
or U26185 (N_26185,N_21665,N_20761);
nor U26186 (N_26186,N_20572,N_20809);
nor U26187 (N_26187,N_24168,N_20834);
and U26188 (N_26188,N_20425,N_24022);
or U26189 (N_26189,N_20997,N_20781);
nor U26190 (N_26190,N_22985,N_23924);
or U26191 (N_26191,N_23786,N_24601);
nor U26192 (N_26192,N_22903,N_23953);
nor U26193 (N_26193,N_23265,N_22350);
nor U26194 (N_26194,N_23573,N_21066);
nand U26195 (N_26195,N_23681,N_24103);
nor U26196 (N_26196,N_22475,N_23767);
and U26197 (N_26197,N_23140,N_23656);
nor U26198 (N_26198,N_20846,N_20697);
or U26199 (N_26199,N_22775,N_21791);
nand U26200 (N_26200,N_21412,N_21353);
or U26201 (N_26201,N_22264,N_21073);
nor U26202 (N_26202,N_21019,N_22935);
or U26203 (N_26203,N_24962,N_21993);
and U26204 (N_26204,N_24777,N_24692);
and U26205 (N_26205,N_23102,N_24524);
nand U26206 (N_26206,N_21499,N_23116);
or U26207 (N_26207,N_24110,N_20040);
or U26208 (N_26208,N_21259,N_21545);
nand U26209 (N_26209,N_22313,N_22471);
nand U26210 (N_26210,N_20484,N_23889);
nand U26211 (N_26211,N_22127,N_20486);
or U26212 (N_26212,N_21028,N_22327);
and U26213 (N_26213,N_21853,N_22364);
nand U26214 (N_26214,N_24572,N_21016);
nand U26215 (N_26215,N_23575,N_24931);
or U26216 (N_26216,N_22941,N_20255);
nand U26217 (N_26217,N_22819,N_24053);
or U26218 (N_26218,N_22721,N_23788);
nand U26219 (N_26219,N_24102,N_20790);
nor U26220 (N_26220,N_22255,N_22132);
xor U26221 (N_26221,N_21024,N_23229);
or U26222 (N_26222,N_23883,N_23089);
and U26223 (N_26223,N_21750,N_22171);
nand U26224 (N_26224,N_24576,N_21136);
nor U26225 (N_26225,N_22369,N_23527);
nor U26226 (N_26226,N_21844,N_22003);
and U26227 (N_26227,N_24773,N_21912);
xnor U26228 (N_26228,N_21307,N_23641);
and U26229 (N_26229,N_23046,N_20904);
nand U26230 (N_26230,N_22295,N_22293);
nor U26231 (N_26231,N_24009,N_21305);
nor U26232 (N_26232,N_24553,N_23617);
and U26233 (N_26233,N_22531,N_20514);
nand U26234 (N_26234,N_20956,N_21788);
nand U26235 (N_26235,N_20611,N_23880);
nand U26236 (N_26236,N_23064,N_21491);
nor U26237 (N_26237,N_23235,N_22532);
or U26238 (N_26238,N_24778,N_20124);
and U26239 (N_26239,N_22519,N_20146);
nor U26240 (N_26240,N_20056,N_20657);
nor U26241 (N_26241,N_22668,N_21869);
nand U26242 (N_26242,N_22799,N_23495);
nand U26243 (N_26243,N_21204,N_21843);
or U26244 (N_26244,N_23362,N_23683);
nand U26245 (N_26245,N_20335,N_22208);
or U26246 (N_26246,N_21549,N_20906);
nor U26247 (N_26247,N_24719,N_21836);
xnor U26248 (N_26248,N_23804,N_21857);
nor U26249 (N_26249,N_23634,N_21873);
nor U26250 (N_26250,N_21685,N_23109);
or U26251 (N_26251,N_20767,N_21531);
nand U26252 (N_26252,N_24815,N_20214);
nand U26253 (N_26253,N_22744,N_20479);
or U26254 (N_26254,N_23941,N_23739);
nor U26255 (N_26255,N_24650,N_20286);
and U26256 (N_26256,N_23626,N_21284);
nand U26257 (N_26257,N_24155,N_24373);
nand U26258 (N_26258,N_21283,N_24721);
nand U26259 (N_26259,N_23511,N_21256);
nor U26260 (N_26260,N_20374,N_21887);
or U26261 (N_26261,N_21107,N_21634);
xor U26262 (N_26262,N_21200,N_24961);
or U26263 (N_26263,N_22665,N_24542);
nor U26264 (N_26264,N_24949,N_22400);
and U26265 (N_26265,N_21624,N_24502);
nor U26266 (N_26266,N_22540,N_20897);
nor U26267 (N_26267,N_22660,N_23654);
and U26268 (N_26268,N_23435,N_22504);
and U26269 (N_26269,N_24531,N_21313);
xnor U26270 (N_26270,N_21326,N_24671);
and U26271 (N_26271,N_20536,N_21436);
nor U26272 (N_26272,N_21526,N_24896);
nor U26273 (N_26273,N_21190,N_20363);
or U26274 (N_26274,N_22713,N_23366);
and U26275 (N_26275,N_23870,N_24571);
or U26276 (N_26276,N_23593,N_22950);
and U26277 (N_26277,N_24923,N_22048);
nor U26278 (N_26278,N_21487,N_23610);
nor U26279 (N_26279,N_22157,N_22011);
or U26280 (N_26280,N_24839,N_20992);
xor U26281 (N_26281,N_20458,N_20240);
xor U26282 (N_26282,N_20353,N_22944);
nor U26283 (N_26283,N_23200,N_21878);
and U26284 (N_26284,N_23193,N_24026);
or U26285 (N_26285,N_24654,N_22298);
nand U26286 (N_26286,N_20802,N_20188);
nand U26287 (N_26287,N_21814,N_20089);
and U26288 (N_26288,N_20639,N_20775);
nor U26289 (N_26289,N_23481,N_20257);
nand U26290 (N_26290,N_24310,N_20233);
and U26291 (N_26291,N_22117,N_21672);
nand U26292 (N_26292,N_23023,N_20842);
and U26293 (N_26293,N_20212,N_22409);
nor U26294 (N_26294,N_22454,N_20221);
or U26295 (N_26295,N_24169,N_22544);
nand U26296 (N_26296,N_20193,N_24438);
and U26297 (N_26297,N_23748,N_24864);
nand U26298 (N_26298,N_23056,N_20777);
nand U26299 (N_26299,N_20274,N_23208);
nor U26300 (N_26300,N_21906,N_20252);
and U26301 (N_26301,N_21048,N_23418);
nor U26302 (N_26302,N_22774,N_20787);
and U26303 (N_26303,N_23050,N_20317);
and U26304 (N_26304,N_21182,N_24322);
and U26305 (N_26305,N_23380,N_24818);
and U26306 (N_26306,N_22719,N_24512);
and U26307 (N_26307,N_20147,N_21786);
nor U26308 (N_26308,N_22194,N_23526);
and U26309 (N_26309,N_20141,N_23415);
nor U26310 (N_26310,N_21148,N_22129);
or U26311 (N_26311,N_22046,N_20459);
or U26312 (N_26312,N_21025,N_24780);
or U26313 (N_26313,N_23704,N_24561);
and U26314 (N_26314,N_20489,N_21575);
or U26315 (N_26315,N_24258,N_22595);
nor U26316 (N_26316,N_20769,N_23173);
or U26317 (N_26317,N_24878,N_24174);
nor U26318 (N_26318,N_22867,N_23094);
and U26319 (N_26319,N_21486,N_21653);
and U26320 (N_26320,N_20083,N_23250);
or U26321 (N_26321,N_22933,N_23403);
xnor U26322 (N_26322,N_22582,N_22017);
and U26323 (N_26323,N_23295,N_23667);
or U26324 (N_26324,N_22548,N_24933);
xnor U26325 (N_26325,N_23045,N_24164);
or U26326 (N_26326,N_22096,N_21966);
nor U26327 (N_26327,N_24011,N_24473);
nand U26328 (N_26328,N_20452,N_24214);
xnor U26329 (N_26329,N_20050,N_24431);
nor U26330 (N_26330,N_24416,N_20538);
nand U26331 (N_26331,N_20645,N_23668);
or U26332 (N_26332,N_21212,N_22893);
and U26333 (N_26333,N_21536,N_22274);
xnor U26334 (N_26334,N_21462,N_21600);
nor U26335 (N_26335,N_23405,N_24463);
nand U26336 (N_26336,N_21955,N_24554);
or U26337 (N_26337,N_20081,N_20168);
nand U26338 (N_26338,N_21410,N_21945);
and U26339 (N_26339,N_23226,N_21761);
and U26340 (N_26340,N_23721,N_20841);
xnor U26341 (N_26341,N_23903,N_22342);
and U26342 (N_26342,N_22758,N_23254);
xnor U26343 (N_26343,N_23726,N_24252);
and U26344 (N_26344,N_22782,N_22152);
and U26345 (N_26345,N_24205,N_24290);
nor U26346 (N_26346,N_20350,N_23197);
or U26347 (N_26347,N_22354,N_24926);
nand U26348 (N_26348,N_23079,N_23120);
nor U26349 (N_26349,N_22810,N_22136);
or U26350 (N_26350,N_22646,N_20555);
xor U26351 (N_26351,N_22141,N_24788);
and U26352 (N_26352,N_24853,N_23766);
and U26353 (N_26353,N_24807,N_21897);
nand U26354 (N_26354,N_22764,N_20508);
nor U26355 (N_26355,N_23111,N_20062);
and U26356 (N_26356,N_23399,N_24822);
or U26357 (N_26357,N_20771,N_20399);
or U26358 (N_26358,N_24538,N_23949);
nand U26359 (N_26359,N_23589,N_24868);
or U26360 (N_26360,N_24639,N_22508);
or U26361 (N_26361,N_20483,N_20054);
or U26362 (N_26362,N_23977,N_24970);
or U26363 (N_26363,N_24284,N_20730);
or U26364 (N_26364,N_20315,N_22672);
nor U26365 (N_26365,N_24408,N_21178);
nor U26366 (N_26366,N_21348,N_22635);
or U26367 (N_26367,N_23615,N_22974);
nor U26368 (N_26368,N_20023,N_21244);
nor U26369 (N_26369,N_21293,N_24004);
and U26370 (N_26370,N_21113,N_22778);
nand U26371 (N_26371,N_23936,N_24638);
nand U26372 (N_26372,N_21069,N_22083);
xor U26373 (N_26373,N_21759,N_21783);
nor U26374 (N_26374,N_22922,N_24667);
nor U26375 (N_26375,N_23194,N_24978);
nor U26376 (N_26376,N_22555,N_24980);
nor U26377 (N_26377,N_23191,N_22594);
nand U26378 (N_26378,N_23017,N_20865);
xnor U26379 (N_26379,N_21884,N_22881);
or U26380 (N_26380,N_21735,N_24905);
or U26381 (N_26381,N_24000,N_23085);
and U26382 (N_26382,N_20848,N_23081);
and U26383 (N_26383,N_21541,N_23666);
nor U26384 (N_26384,N_23857,N_21532);
and U26385 (N_26385,N_21441,N_23092);
nor U26386 (N_26386,N_20354,N_20932);
nor U26387 (N_26387,N_24272,N_21070);
nor U26388 (N_26388,N_21686,N_23906);
or U26389 (N_26389,N_23572,N_21415);
nor U26390 (N_26390,N_21169,N_24685);
and U26391 (N_26391,N_23451,N_20975);
or U26392 (N_26392,N_24881,N_20649);
and U26393 (N_26393,N_24259,N_23165);
nor U26394 (N_26394,N_24915,N_24616);
nor U26395 (N_26395,N_23218,N_21143);
nand U26396 (N_26396,N_20037,N_20965);
or U26397 (N_26397,N_22591,N_21849);
and U26398 (N_26398,N_22983,N_22527);
nand U26399 (N_26399,N_22724,N_22247);
or U26400 (N_26400,N_24735,N_22890);
nor U26401 (N_26401,N_23277,N_23501);
nand U26402 (N_26402,N_23973,N_24643);
nor U26403 (N_26403,N_20499,N_20573);
or U26404 (N_26404,N_24122,N_23457);
and U26405 (N_26405,N_20069,N_23164);
nand U26406 (N_26406,N_24099,N_22908);
nand U26407 (N_26407,N_24454,N_21496);
nor U26408 (N_26408,N_23660,N_22121);
nand U26409 (N_26409,N_24468,N_20196);
or U26410 (N_26410,N_20646,N_21935);
or U26411 (N_26411,N_20966,N_22390);
or U26412 (N_26412,N_23422,N_24790);
or U26413 (N_26413,N_20051,N_22269);
and U26414 (N_26414,N_22917,N_22367);
and U26415 (N_26415,N_23161,N_24861);
and U26416 (N_26416,N_23579,N_21524);
nor U26417 (N_26417,N_20988,N_21756);
nand U26418 (N_26418,N_23694,N_23093);
and U26419 (N_26419,N_21375,N_20473);
and U26420 (N_26420,N_24596,N_23974);
or U26421 (N_26421,N_24117,N_24218);
and U26422 (N_26422,N_23247,N_24282);
xnor U26423 (N_26423,N_24160,N_21682);
or U26424 (N_26424,N_20880,N_20516);
nand U26425 (N_26425,N_22753,N_20074);
and U26426 (N_26426,N_21092,N_20136);
nand U26427 (N_26427,N_23156,N_22861);
and U26428 (N_26428,N_23461,N_21488);
or U26429 (N_26429,N_24884,N_24093);
and U26430 (N_26430,N_20510,N_24417);
and U26431 (N_26431,N_20845,N_21896);
nor U26432 (N_26432,N_23448,N_22886);
xor U26433 (N_26433,N_23386,N_21034);
nor U26434 (N_26434,N_21877,N_24353);
nor U26435 (N_26435,N_24641,N_22656);
nor U26436 (N_26436,N_20369,N_23180);
or U26437 (N_26437,N_20200,N_24567);
nand U26438 (N_26438,N_21261,N_21331);
nor U26439 (N_26439,N_20179,N_21449);
and U26440 (N_26440,N_23744,N_24461);
nand U26441 (N_26441,N_24370,N_20039);
xnor U26442 (N_26442,N_23756,N_23413);
nor U26443 (N_26443,N_22875,N_23678);
and U26444 (N_26444,N_21584,N_22033);
nand U26445 (N_26445,N_24075,N_20090);
nor U26446 (N_26446,N_20063,N_23900);
or U26447 (N_26447,N_23113,N_24352);
xor U26448 (N_26448,N_23131,N_21593);
nor U26449 (N_26449,N_23166,N_23627);
nor U26450 (N_26450,N_22754,N_20586);
nor U26451 (N_26451,N_22894,N_24393);
and U26452 (N_26452,N_21160,N_20191);
or U26453 (N_26453,N_24722,N_20073);
and U26454 (N_26454,N_22833,N_21889);
nand U26455 (N_26455,N_21987,N_23118);
xnor U26456 (N_26456,N_22939,N_22821);
and U26457 (N_26457,N_24219,N_20440);
and U26458 (N_26458,N_21362,N_24343);
or U26459 (N_26459,N_21700,N_24536);
or U26460 (N_26460,N_23196,N_20667);
or U26461 (N_26461,N_21081,N_24129);
nor U26462 (N_26462,N_21087,N_23556);
nand U26463 (N_26463,N_21518,N_21461);
and U26464 (N_26464,N_22638,N_24404);
nand U26465 (N_26465,N_20670,N_20166);
nor U26466 (N_26466,N_20546,N_24824);
nor U26467 (N_26467,N_22969,N_22473);
xnor U26468 (N_26468,N_24456,N_24073);
nor U26469 (N_26469,N_21352,N_20739);
or U26470 (N_26470,N_21971,N_20405);
and U26471 (N_26471,N_20475,N_20656);
nand U26472 (N_26472,N_21158,N_23701);
and U26473 (N_26473,N_23803,N_22182);
nor U26474 (N_26474,N_24460,N_21726);
nor U26475 (N_26475,N_22164,N_22664);
nand U26476 (N_26476,N_22291,N_20665);
nand U26477 (N_26477,N_21361,N_24445);
or U26478 (N_26478,N_21495,N_24357);
or U26479 (N_26479,N_20014,N_23888);
or U26480 (N_26480,N_21380,N_21465);
and U26481 (N_26481,N_23469,N_23097);
nor U26482 (N_26482,N_20548,N_20589);
nand U26483 (N_26483,N_22765,N_23130);
nand U26484 (N_26484,N_20044,N_21911);
nand U26485 (N_26485,N_21147,N_24086);
nor U26486 (N_26486,N_22051,N_22253);
and U26487 (N_26487,N_24604,N_23223);
xnor U26488 (N_26488,N_24030,N_21218);
or U26489 (N_26489,N_21445,N_22997);
nand U26490 (N_26490,N_23679,N_22539);
xnor U26491 (N_26491,N_22523,N_20067);
nor U26492 (N_26492,N_23814,N_21268);
and U26493 (N_26493,N_21280,N_20377);
or U26494 (N_26494,N_22554,N_21299);
or U26495 (N_26495,N_23110,N_24766);
and U26496 (N_26496,N_22144,N_24997);
nor U26497 (N_26497,N_24689,N_23163);
nand U26498 (N_26498,N_24608,N_20794);
or U26499 (N_26499,N_24137,N_23367);
or U26500 (N_26500,N_22260,N_23868);
nand U26501 (N_26501,N_23044,N_24235);
or U26502 (N_26502,N_20075,N_23922);
xnor U26503 (N_26503,N_20390,N_22338);
nand U26504 (N_26504,N_21063,N_21895);
nand U26505 (N_26505,N_21807,N_21124);
and U26506 (N_26506,N_20710,N_21739);
nor U26507 (N_26507,N_23874,N_20003);
and U26508 (N_26508,N_23106,N_23203);
xor U26509 (N_26509,N_21823,N_23429);
or U26510 (N_26510,N_21151,N_24889);
and U26511 (N_26511,N_20608,N_24704);
nand U26512 (N_26512,N_22304,N_20911);
and U26513 (N_26513,N_22965,N_22396);
nor U26514 (N_26514,N_24784,N_24190);
nor U26515 (N_26515,N_23987,N_24049);
nand U26516 (N_26516,N_20731,N_23853);
nor U26517 (N_26517,N_21346,N_23985);
nand U26518 (N_26518,N_23671,N_22213);
nor U26519 (N_26519,N_20843,N_22844);
or U26520 (N_26520,N_24763,N_21959);
and U26521 (N_26521,N_20349,N_20700);
and U26522 (N_26522,N_24767,N_20669);
nor U26523 (N_26523,N_22148,N_23840);
nor U26524 (N_26524,N_21456,N_24096);
and U26525 (N_26525,N_21659,N_24196);
and U26526 (N_26526,N_24158,N_20132);
nor U26527 (N_26527,N_24183,N_21453);
nand U26528 (N_26528,N_21802,N_21162);
nor U26529 (N_26529,N_23533,N_23558);
nor U26530 (N_26530,N_20006,N_20013);
and U26531 (N_26531,N_21667,N_20020);
and U26532 (N_26532,N_24757,N_23960);
nor U26533 (N_26533,N_22686,N_21860);
and U26534 (N_26534,N_23991,N_22979);
and U26535 (N_26535,N_20364,N_24351);
and U26536 (N_26536,N_20853,N_21501);
nor U26537 (N_26537,N_22623,N_21848);
xor U26538 (N_26538,N_22178,N_20742);
or U26539 (N_26539,N_22240,N_20248);
nor U26540 (N_26540,N_23584,N_21298);
nand U26541 (N_26541,N_22854,N_22725);
or U26542 (N_26542,N_23178,N_22788);
and U26543 (N_26543,N_20851,N_21308);
nand U26544 (N_26544,N_20245,N_24727);
or U26545 (N_26545,N_23071,N_22426);
or U26546 (N_26546,N_21484,N_23410);
and U26547 (N_26547,N_22848,N_22650);
nor U26548 (N_26548,N_21154,N_21695);
nand U26549 (N_26549,N_23058,N_20893);
nor U26550 (N_26550,N_22420,N_24230);
and U26551 (N_26551,N_22280,N_22366);
and U26552 (N_26552,N_20928,N_22561);
nand U26553 (N_26553,N_23630,N_23688);
nand U26554 (N_26554,N_23188,N_21020);
and U26555 (N_26555,N_24467,N_21392);
or U26556 (N_26556,N_20967,N_21121);
or U26557 (N_26557,N_22530,N_24172);
nand U26558 (N_26558,N_23187,N_22061);
nor U26559 (N_26559,N_23592,N_23780);
or U26560 (N_26560,N_23560,N_20833);
nor U26561 (N_26561,N_23587,N_24295);
and U26562 (N_26562,N_20738,N_20850);
nor U26563 (N_26563,N_20386,N_20989);
nand U26564 (N_26564,N_20824,N_23517);
or U26565 (N_26565,N_21373,N_21838);
nand U26566 (N_26566,N_20634,N_24010);
nor U26567 (N_26567,N_21785,N_20813);
nor U26568 (N_26568,N_24953,N_21135);
and U26569 (N_26569,N_21764,N_24299);
xnor U26570 (N_26570,N_23485,N_22947);
or U26571 (N_26571,N_24789,N_23207);
and U26572 (N_26572,N_21302,N_22884);
nand U26573 (N_26573,N_23057,N_21356);
nand U26574 (N_26574,N_22284,N_20030);
nor U26575 (N_26575,N_22436,N_20455);
nand U26576 (N_26576,N_23488,N_22122);
nor U26577 (N_26577,N_24796,N_23931);
or U26578 (N_26578,N_22670,N_20302);
nor U26579 (N_26579,N_21719,N_23952);
nand U26580 (N_26580,N_22263,N_21490);
or U26581 (N_26581,N_24856,N_20421);
nand U26582 (N_26582,N_20680,N_23202);
xor U26583 (N_26583,N_21768,N_22326);
nand U26584 (N_26584,N_20876,N_23496);
nor U26585 (N_26585,N_24508,N_21736);
or U26586 (N_26586,N_20167,N_21477);
and U26587 (N_26587,N_23725,N_22563);
xor U26588 (N_26588,N_23041,N_20576);
nor U26589 (N_26589,N_20348,N_20228);
nand U26590 (N_26590,N_21014,N_21117);
nand U26591 (N_26591,N_20613,N_22153);
nor U26592 (N_26592,N_23759,N_21936);
xor U26593 (N_26593,N_23699,N_24659);
nand U26594 (N_26594,N_23893,N_23134);
or U26595 (N_26595,N_20946,N_22662);
nor U26596 (N_26596,N_22045,N_21110);
nand U26597 (N_26597,N_23414,N_23623);
xnor U26598 (N_26598,N_21931,N_20355);
or U26599 (N_26599,N_23375,N_21890);
and U26600 (N_26600,N_23806,N_21018);
or U26601 (N_26601,N_23799,N_21696);
nand U26602 (N_26602,N_24249,N_20938);
nand U26603 (N_26603,N_23257,N_20181);
or U26604 (N_26604,N_22074,N_21199);
and U26605 (N_26605,N_20461,N_20198);
nor U26606 (N_26606,N_21742,N_22885);
xor U26607 (N_26607,N_22658,N_22043);
and U26608 (N_26608,N_22515,N_22125);
and U26609 (N_26609,N_23812,N_24306);
nand U26610 (N_26610,N_23052,N_23239);
and U26611 (N_26611,N_20900,N_23757);
nand U26612 (N_26612,N_23719,N_22382);
or U26613 (N_26613,N_21022,N_21588);
or U26614 (N_26614,N_21636,N_20862);
xor U26615 (N_26615,N_24694,N_22731);
or U26616 (N_26616,N_21097,N_22198);
xnor U26617 (N_26617,N_21608,N_23423);
nor U26618 (N_26618,N_24135,N_22988);
and U26619 (N_26619,N_22365,N_20884);
and U26620 (N_26620,N_21893,N_24039);
nand U26621 (N_26621,N_22007,N_23000);
xor U26622 (N_26622,N_23396,N_21385);
or U26623 (N_26623,N_24637,N_21835);
nor U26624 (N_26624,N_21464,N_21528);
and U26625 (N_26625,N_24262,N_22608);
nor U26626 (N_26626,N_22092,N_22745);
nand U26627 (N_26627,N_24256,N_22823);
nor U26628 (N_26628,N_24243,N_20774);
nor U26629 (N_26629,N_24821,N_21287);
or U26630 (N_26630,N_22726,N_23677);
and U26631 (N_26631,N_24976,N_24107);
nand U26632 (N_26632,N_21924,N_24885);
and U26633 (N_26633,N_22175,N_20060);
nor U26634 (N_26634,N_23039,N_23138);
nand U26635 (N_26635,N_22075,N_24098);
nor U26636 (N_26636,N_20190,N_24391);
nor U26637 (N_26637,N_22599,N_20815);
nor U26638 (N_26638,N_20901,N_22698);
or U26639 (N_26639,N_23655,N_21192);
and U26640 (N_26640,N_21805,N_21727);
and U26641 (N_26641,N_21340,N_21871);
and U26642 (N_26642,N_24008,N_22526);
and U26643 (N_26643,N_20505,N_23908);
nor U26644 (N_26644,N_20859,N_21561);
nor U26645 (N_26645,N_20960,N_21763);
or U26646 (N_26646,N_23794,N_21079);
nor U26647 (N_26647,N_20871,N_20391);
or U26648 (N_26648,N_22483,N_21423);
nor U26649 (N_26649,N_23258,N_23301);
nor U26650 (N_26650,N_20361,N_22050);
xor U26651 (N_26651,N_21105,N_23364);
nor U26652 (N_26652,N_23753,N_21285);
nand U26653 (N_26653,N_21211,N_23676);
nor U26654 (N_26654,N_21675,N_20482);
nand U26655 (N_26655,N_21294,N_24627);
or U26656 (N_26656,N_21861,N_23823);
or U26657 (N_26657,N_20406,N_22139);
and U26658 (N_26658,N_21480,N_22565);
or U26659 (N_26659,N_24768,N_24275);
xnor U26660 (N_26660,N_23536,N_22261);
and U26661 (N_26661,N_22187,N_23105);
and U26662 (N_26662,N_22193,N_23927);
nand U26663 (N_26663,N_22741,N_23934);
or U26664 (N_26664,N_21387,N_22617);
xor U26665 (N_26665,N_21980,N_24817);
nor U26666 (N_26666,N_23918,N_20979);
or U26667 (N_26667,N_20708,N_24080);
nand U26668 (N_26668,N_21126,N_21978);
and U26669 (N_26669,N_24590,N_23416);
or U26670 (N_26670,N_21684,N_21297);
nand U26671 (N_26671,N_23234,N_21801);
nand U26672 (N_26672,N_22772,N_23100);
nand U26673 (N_26673,N_22166,N_22716);
nand U26674 (N_26674,N_24311,N_20718);
or U26675 (N_26675,N_21691,N_24283);
nor U26676 (N_26676,N_23115,N_20628);
nor U26677 (N_26677,N_22839,N_24619);
nand U26678 (N_26678,N_20801,N_24594);
or U26679 (N_26679,N_21149,N_23521);
nor U26680 (N_26680,N_24421,N_24622);
nor U26681 (N_26681,N_22606,N_22723);
and U26682 (N_26682,N_23542,N_24918);
xor U26683 (N_26683,N_21976,N_23147);
and U26684 (N_26684,N_21963,N_20588);
nor U26685 (N_26685,N_21222,N_20640);
xor U26686 (N_26686,N_24715,N_23042);
and U26687 (N_26687,N_21651,N_22391);
nor U26688 (N_26688,N_21547,N_22130);
xor U26689 (N_26689,N_22470,N_20707);
nand U26690 (N_26690,N_20996,N_20379);
nor U26691 (N_26691,N_23484,N_21378);
or U26692 (N_26692,N_23898,N_23769);
and U26693 (N_26693,N_24414,N_24617);
and U26694 (N_26694,N_22900,N_21152);
nand U26695 (N_26695,N_23848,N_21196);
or U26696 (N_26696,N_22228,N_20117);
nor U26697 (N_26697,N_21885,N_21274);
and U26698 (N_26698,N_23995,N_21995);
nand U26699 (N_26699,N_23807,N_24197);
nand U26700 (N_26700,N_21826,N_21977);
or U26701 (N_26701,N_21952,N_24335);
nand U26702 (N_26702,N_23946,N_21037);
nor U26703 (N_26703,N_23459,N_22786);
and U26704 (N_26704,N_24191,N_23964);
nor U26705 (N_26705,N_21359,N_22734);
nor U26706 (N_26706,N_23956,N_22616);
or U26707 (N_26707,N_21619,N_21707);
or U26708 (N_26708,N_24333,N_23361);
nor U26709 (N_26709,N_21886,N_20138);
or U26710 (N_26710,N_22843,N_23103);
nor U26711 (N_26711,N_22049,N_20189);
and U26712 (N_26712,N_24793,N_22975);
xnor U26713 (N_26713,N_24630,N_24774);
and U26714 (N_26714,N_21478,N_20410);
and U26715 (N_26715,N_24286,N_24642);
nand U26716 (N_26716,N_24170,N_23168);
or U26717 (N_26717,N_23545,N_21628);
or U26718 (N_26718,N_22996,N_24325);
nand U26719 (N_26719,N_24293,N_23494);
nand U26720 (N_26720,N_22405,N_24606);
or U26721 (N_26721,N_20891,N_20688);
and U26722 (N_26722,N_24329,N_24061);
or U26723 (N_26723,N_20564,N_22906);
nor U26724 (N_26724,N_20071,N_22285);
and U26725 (N_26725,N_22710,N_22831);
or U26726 (N_26726,N_21011,N_23217);
xor U26727 (N_26727,N_22076,N_23951);
and U26728 (N_26728,N_24324,N_20570);
xnor U26729 (N_26729,N_23339,N_22787);
nor U26730 (N_26730,N_21777,N_24397);
nand U26731 (N_26731,N_24599,N_24041);
xnor U26732 (N_26732,N_24437,N_20933);
or U26733 (N_26733,N_21400,N_21206);
and U26734 (N_26734,N_24582,N_20821);
nand U26735 (N_26735,N_24388,N_22310);
and U26736 (N_26736,N_24369,N_24660);
and U26737 (N_26737,N_22568,N_21460);
nor U26738 (N_26738,N_22836,N_21505);
nor U26739 (N_26739,N_20713,N_24901);
nand U26740 (N_26740,N_21797,N_24271);
nand U26741 (N_26741,N_23293,N_24348);
or U26742 (N_26742,N_24801,N_23813);
nor U26743 (N_26743,N_22487,N_20822);
nand U26744 (N_26744,N_22100,N_22163);
or U26745 (N_26745,N_21888,N_24378);
nor U26746 (N_26746,N_21627,N_22282);
nor U26747 (N_26747,N_20488,N_23763);
and U26748 (N_26748,N_20203,N_21459);
and U26749 (N_26749,N_24362,N_22099);
xor U26750 (N_26750,N_24074,N_20323);
nor U26751 (N_26751,N_23160,N_21391);
and U26752 (N_26752,N_23222,N_24206);
or U26753 (N_26753,N_20783,N_23747);
or U26754 (N_26754,N_21829,N_22970);
and U26755 (N_26755,N_23827,N_23390);
or U26756 (N_26756,N_23742,N_22934);
or U26757 (N_26757,N_21865,N_23632);
and U26758 (N_26758,N_24880,N_23635);
and U26759 (N_26759,N_20766,N_24623);
nand U26760 (N_26760,N_22570,N_20835);
nand U26761 (N_26761,N_23419,N_21013);
nand U26762 (N_26762,N_22444,N_22932);
nand U26763 (N_26763,N_23137,N_20869);
nand U26764 (N_26764,N_24776,N_21973);
nand U26765 (N_26765,N_24031,N_21752);
or U26766 (N_26766,N_21625,N_20388);
and U26767 (N_26767,N_23712,N_20800);
nor U26768 (N_26768,N_23792,N_24338);
nand U26769 (N_26769,N_24547,N_24292);
or U26770 (N_26770,N_23167,N_20453);
or U26771 (N_26771,N_21943,N_20152);
nor U26772 (N_26772,N_23313,N_20929);
nor U26773 (N_26773,N_21830,N_20704);
nand U26774 (N_26774,N_20362,N_22918);
xnor U26775 (N_26775,N_20537,N_20671);
xor U26776 (N_26776,N_23516,N_22738);
nor U26777 (N_26777,N_22702,N_21052);
nand U26778 (N_26778,N_21595,N_20617);
nor U26779 (N_26779,N_21606,N_20048);
nand U26780 (N_26780,N_21422,N_21104);
or U26781 (N_26781,N_22615,N_23290);
nor U26782 (N_26782,N_20838,N_22463);
nand U26783 (N_26783,N_22558,N_23789);
or U26784 (N_26784,N_22465,N_22991);
and U26785 (N_26785,N_21771,N_23199);
nor U26786 (N_26786,N_21292,N_23055);
nor U26787 (N_26787,N_23530,N_20970);
and U26788 (N_26788,N_22828,N_23771);
or U26789 (N_26789,N_21732,N_24848);
nor U26790 (N_26790,N_23600,N_21046);
and U26791 (N_26791,N_22372,N_24260);
or U26792 (N_26792,N_24162,N_22840);
nand U26793 (N_26793,N_20278,N_23299);
and U26794 (N_26794,N_23894,N_24871);
nand U26795 (N_26795,N_24471,N_20441);
nand U26796 (N_26796,N_21633,N_23862);
nand U26797 (N_26797,N_20685,N_21173);
and U26798 (N_26798,N_21614,N_24575);
or U26799 (N_26799,N_21650,N_20972);
xnor U26800 (N_26800,N_23999,N_24597);
and U26801 (N_26801,N_24211,N_22695);
or U26802 (N_26802,N_22289,N_22987);
or U26803 (N_26803,N_24459,N_24646);
nand U26804 (N_26804,N_23231,N_21751);
nand U26805 (N_26805,N_21103,N_20085);
and U26806 (N_26806,N_20793,N_22851);
and U26807 (N_26807,N_21075,N_23842);
nor U26808 (N_26808,N_21645,N_23582);
nand U26809 (N_26809,N_24895,N_21476);
or U26810 (N_26810,N_24132,N_24523);
nor U26811 (N_26811,N_21702,N_22196);
or U26812 (N_26812,N_22560,N_24403);
nor U26813 (N_26813,N_22584,N_24114);
nand U26814 (N_26814,N_23875,N_22942);
nor U26815 (N_26815,N_20968,N_20404);
or U26816 (N_26816,N_22377,N_23145);
and U26817 (N_26817,N_23334,N_20728);
nor U26818 (N_26818,N_24327,N_20140);
xnor U26819 (N_26819,N_22812,N_23347);
and U26820 (N_26820,N_20446,N_23363);
xor U26821 (N_26821,N_21731,N_22008);
or U26822 (N_26822,N_24708,N_20176);
nor U26823 (N_26823,N_20276,N_24490);
or U26824 (N_26824,N_23031,N_22472);
or U26825 (N_26825,N_24612,N_24710);
nand U26826 (N_26826,N_21594,N_21590);
and U26827 (N_26827,N_22339,N_21811);
nand U26828 (N_26828,N_21989,N_21567);
nor U26829 (N_26829,N_20174,N_21041);
nand U26830 (N_26830,N_21345,N_24985);
nand U26831 (N_26831,N_23379,N_21333);
or U26832 (N_26832,N_20599,N_22057);
or U26833 (N_26833,N_22180,N_22645);
nand U26834 (N_26834,N_23619,N_21716);
nor U26835 (N_26835,N_21085,N_20594);
nor U26836 (N_26836,N_23264,N_24930);
or U26837 (N_26837,N_24186,N_20086);
xor U26838 (N_26838,N_20338,N_22912);
xnor U26839 (N_26839,N_21234,N_24624);
or U26840 (N_26840,N_23932,N_24598);
nor U26841 (N_26841,N_22235,N_22556);
and U26842 (N_26842,N_20959,N_22691);
nor U26843 (N_26843,N_20711,N_20957);
or U26844 (N_26844,N_23392,N_23142);
or U26845 (N_26845,N_23259,N_22387);
or U26846 (N_26846,N_24381,N_24527);
and U26847 (N_26847,N_23735,N_20277);
and U26848 (N_26848,N_22880,N_22010);
and U26849 (N_26849,N_22757,N_22815);
nand U26850 (N_26850,N_21354,N_21051);
nor U26851 (N_26851,N_24702,N_21855);
nor U26852 (N_26852,N_21523,N_24857);
and U26853 (N_26853,N_21223,N_22191);
xor U26854 (N_26854,N_23450,N_20779);
or U26855 (N_26855,N_24216,N_20719);
nor U26856 (N_26856,N_24911,N_21388);
xnor U26857 (N_26857,N_24078,N_22053);
nor U26858 (N_26858,N_23340,N_24312);
and U26859 (N_26859,N_24602,N_22636);
nand U26860 (N_26860,N_23957,N_22029);
or U26861 (N_26861,N_24185,N_21232);
nor U26862 (N_26862,N_20272,N_22770);
nand U26863 (N_26863,N_20161,N_23886);
and U26864 (N_26864,N_22222,N_23841);
nor U26865 (N_26865,N_23248,N_20515);
nor U26866 (N_26866,N_24847,N_24772);
or U26867 (N_26867,N_21983,N_23998);
nor U26868 (N_26868,N_23009,N_21705);
or U26869 (N_26869,N_21195,N_21674);
or U26870 (N_26870,N_24435,N_24043);
xnor U26871 (N_26871,N_24877,N_21418);
or U26872 (N_26872,N_20565,N_22268);
nand U26873 (N_26873,N_20547,N_24392);
nor U26874 (N_26874,N_24786,N_20016);
or U26875 (N_26875,N_22343,N_24862);
or U26876 (N_26876,N_23963,N_22457);
and U26877 (N_26877,N_24947,N_24250);
nand U26878 (N_26878,N_20101,N_22629);
and U26879 (N_26879,N_22456,N_20432);
nor U26880 (N_26880,N_23525,N_24840);
nor U26881 (N_26881,N_20934,N_20955);
and U26882 (N_26882,N_20449,N_22052);
nand U26883 (N_26883,N_21715,N_21012);
and U26884 (N_26884,N_21271,N_23745);
and U26885 (N_26885,N_24365,N_24744);
or U26886 (N_26886,N_22693,N_22020);
nor U26887 (N_26887,N_20135,N_22312);
nand U26888 (N_26888,N_21295,N_20457);
and U26889 (N_26889,N_23227,N_21267);
or U26890 (N_26890,N_24372,N_22265);
nand U26891 (N_26891,N_22620,N_22181);
nor U26892 (N_26892,N_21902,N_23910);
nor U26893 (N_26893,N_20826,N_20112);
and U26894 (N_26894,N_23781,N_21481);
or U26895 (N_26895,N_23402,N_21708);
nand U26896 (N_26896,N_24241,N_22410);
xnor U26897 (N_26897,N_22567,N_24743);
and U26898 (N_26898,N_22962,N_20726);
xnor U26899 (N_26899,N_21999,N_22262);
or U26900 (N_26900,N_20036,N_21439);
or U26901 (N_26901,N_24587,N_21581);
nor U26902 (N_26902,N_22306,N_23096);
nor U26903 (N_26903,N_24740,N_21440);
nor U26904 (N_26904,N_22307,N_23324);
nor U26905 (N_26905,N_23736,N_22244);
nor U26906 (N_26906,N_23465,N_20725);
or U26907 (N_26907,N_23037,N_20096);
and U26908 (N_26908,N_20776,N_20297);
nand U26909 (N_26909,N_20171,N_24811);
or U26910 (N_26910,N_23754,N_20895);
and U26911 (N_26911,N_22242,N_24883);
xor U26912 (N_26912,N_21922,N_22394);
or U26913 (N_26913,N_22477,N_20400);
nand U26914 (N_26914,N_20909,N_20630);
and U26915 (N_26915,N_24320,N_20856);
or U26916 (N_26916,N_24337,N_22131);
and U26917 (N_26917,N_21198,N_21472);
nand U26918 (N_26918,N_23273,N_24945);
and U26919 (N_26919,N_21520,N_21794);
xnor U26920 (N_26920,N_20468,N_22618);
nor U26921 (N_26921,N_23043,N_21646);
nor U26922 (N_26922,N_20647,N_20308);
and U26923 (N_26923,N_21554,N_22547);
or U26924 (N_26924,N_24452,N_21507);
and U26925 (N_26925,N_23585,N_20371);
nor U26926 (N_26926,N_21429,N_20758);
nor U26927 (N_26927,N_21057,N_24557);
and U26928 (N_26928,N_20553,N_24543);
nor U26929 (N_26929,N_23702,N_22418);
nand U26930 (N_26930,N_22866,N_24350);
xor U26931 (N_26931,N_20426,N_21253);
nor U26932 (N_26932,N_20678,N_20568);
or U26933 (N_26933,N_24874,N_22440);
nor U26934 (N_26934,N_23782,N_22863);
nor U26935 (N_26935,N_22783,N_24753);
xnor U26936 (N_26936,N_20310,N_23179);
nand U26937 (N_26937,N_20156,N_22297);
nand U26938 (N_26938,N_23151,N_23847);
and U26939 (N_26939,N_24514,N_22065);
or U26940 (N_26940,N_24653,N_21571);
and U26941 (N_26941,N_23534,N_21458);
and U26942 (N_26942,N_20743,N_22072);
nand U26943 (N_26943,N_22901,N_23305);
nand U26944 (N_26944,N_22524,N_22419);
or U26945 (N_26945,N_21003,N_23003);
and U26946 (N_26946,N_21741,N_20574);
and U26947 (N_26947,N_23791,N_22545);
nand U26948 (N_26948,N_20270,N_24956);
and U26949 (N_26949,N_23674,N_24737);
nand U26950 (N_26950,N_20857,N_20816);
nor U26951 (N_26951,N_20367,N_22801);
nor U26952 (N_26952,N_23350,N_23371);
nand U26953 (N_26953,N_24045,N_20825);
nor U26954 (N_26954,N_21930,N_24805);
nor U26955 (N_26955,N_20748,N_23595);
and U26956 (N_26956,N_21552,N_20501);
nand U26957 (N_26957,N_23400,N_24613);
nor U26958 (N_26958,N_20879,N_20419);
and U26959 (N_26959,N_21747,N_24634);
nor U26960 (N_26960,N_22609,N_20263);
nor U26961 (N_26961,N_24661,N_24318);
nand U26962 (N_26962,N_20026,N_21364);
nand U26963 (N_26963,N_23090,N_20653);
and U26964 (N_26964,N_21847,N_22796);
or U26965 (N_26965,N_24013,N_23275);
and U26966 (N_26966,N_24819,N_24054);
nand U26967 (N_26967,N_24558,N_23664);
nor U26968 (N_26968,N_20736,N_22627);
and U26969 (N_26969,N_21894,N_21717);
and U26970 (N_26970,N_24826,N_23352);
and U26971 (N_26971,N_24825,N_21875);
nor U26972 (N_26972,N_22485,N_21565);
or U26973 (N_26973,N_24410,N_22490);
nor U26974 (N_26974,N_21330,N_21683);
nor U26975 (N_26975,N_21115,N_20701);
nor U26976 (N_26976,N_23348,N_24647);
nand U26977 (N_26977,N_21432,N_24119);
nor U26978 (N_26978,N_24323,N_20917);
or U26979 (N_26979,N_24278,N_24313);
nand U26980 (N_26980,N_23817,N_22318);
or U26981 (N_26981,N_20659,N_21071);
or U26982 (N_26982,N_24194,N_23815);
nand U26983 (N_26983,N_21918,N_24843);
or U26984 (N_26984,N_21032,N_23855);
xor U26985 (N_26985,N_21343,N_24500);
nand U26986 (N_26986,N_20454,N_22857);
and U26987 (N_26987,N_23185,N_23393);
nor U26988 (N_26988,N_21666,N_22012);
and U26989 (N_26989,N_24375,N_20926);
and U26990 (N_26990,N_24955,N_20469);
and U26991 (N_26991,N_20327,N_22432);
and U26992 (N_26992,N_20007,N_21766);
nor U26993 (N_26993,N_21789,N_20098);
or U26994 (N_26994,N_24390,N_24052);
and U26995 (N_26995,N_21093,N_20064);
nor U26996 (N_26996,N_21191,N_24672);
or U26997 (N_26997,N_23487,N_23800);
nor U26998 (N_26998,N_20178,N_23578);
and U26999 (N_26999,N_20175,N_24297);
or U27000 (N_27000,N_20609,N_24509);
and U27001 (N_27001,N_20549,N_20041);
nand U27002 (N_27002,N_24303,N_22385);
nand U27003 (N_27003,N_23060,N_23652);
and U27004 (N_27004,N_24941,N_23075);
or U27005 (N_27005,N_20849,N_21189);
nor U27006 (N_27006,N_24986,N_21953);
nor U27007 (N_27007,N_24687,N_20597);
or U27008 (N_27008,N_20159,N_21806);
or U27009 (N_27009,N_20169,N_23933);
nor U27010 (N_27010,N_24882,N_20422);
nand U27011 (N_27011,N_21138,N_20442);
xor U27012 (N_27012,N_24204,N_23395);
or U27013 (N_27013,N_20032,N_24562);
and U27014 (N_27014,N_23983,N_22809);
and U27015 (N_27015,N_21064,N_22760);
nor U27016 (N_27016,N_23213,N_24525);
and U27017 (N_27017,N_23288,N_21089);
or U27018 (N_27018,N_21498,N_24515);
or U27019 (N_27019,N_21776,N_20396);
nor U27020 (N_27020,N_21546,N_20344);
and U27021 (N_27021,N_22016,N_24182);
nor U27022 (N_27022,N_23711,N_23920);
nand U27023 (N_27023,N_22036,N_24060);
or U27024 (N_27024,N_22381,N_20072);
or U27025 (N_27025,N_22161,N_22042);
or U27026 (N_27026,N_20585,N_23283);
nor U27027 (N_27027,N_20764,N_23076);
or U27028 (N_27028,N_20389,N_23337);
or U27029 (N_27029,N_24971,N_20285);
nor U27030 (N_27030,N_21226,N_24910);
nor U27031 (N_27031,N_24803,N_23879);
nand U27032 (N_27032,N_23510,N_22145);
nor U27033 (N_27033,N_20250,N_22883);
nor U27034 (N_27034,N_24356,N_24765);
nor U27035 (N_27035,N_23629,N_20559);
and U27036 (N_27036,N_23899,N_24973);
and U27037 (N_27037,N_20729,N_22896);
or U27038 (N_27038,N_20986,N_23731);
or U27039 (N_27039,N_24140,N_23713);
or U27040 (N_27040,N_22925,N_22424);
or U27041 (N_27041,N_21631,N_22811);
xnor U27042 (N_27042,N_21236,N_20689);
nor U27043 (N_27043,N_20418,N_21701);
and U27044 (N_27044,N_21435,N_21053);
or U27045 (N_27045,N_20237,N_20631);
nor U27046 (N_27046,N_24711,N_20951);
nor U27047 (N_27047,N_21697,N_20244);
or U27048 (N_27048,N_20525,N_24300);
or U27049 (N_27049,N_21533,N_23099);
or U27050 (N_27050,N_21503,N_23246);
nand U27051 (N_27051,N_23937,N_22105);
nor U27052 (N_27052,N_21921,N_21859);
and U27053 (N_27053,N_22749,N_24070);
nand U27054 (N_27054,N_24387,N_23821);
nand U27055 (N_27055,N_24909,N_21166);
nand U27056 (N_27056,N_20401,N_21334);
and U27057 (N_27057,N_23341,N_20741);
nor U27058 (N_27058,N_21029,N_20247);
and U27059 (N_27059,N_20106,N_21036);
nand U27060 (N_27060,N_21626,N_24192);
nand U27061 (N_27061,N_24128,N_22413);
nand U27062 (N_27062,N_24991,N_22943);
nor U27063 (N_27063,N_22589,N_20387);
nor U27064 (N_27064,N_22249,N_24798);
nand U27065 (N_27065,N_23869,N_21172);
nand U27066 (N_27066,N_24908,N_20273);
nand U27067 (N_27067,N_20209,N_23645);
or U27068 (N_27068,N_22838,N_21557);
or U27069 (N_27069,N_22492,N_22784);
nor U27070 (N_27070,N_24761,N_22279);
nand U27071 (N_27071,N_20215,N_22186);
nand U27072 (N_27072,N_23518,N_21669);
or U27073 (N_27073,N_22189,N_22402);
nor U27074 (N_27074,N_23722,N_22992);
nor U27075 (N_27075,N_21139,N_22685);
xnor U27076 (N_27076,N_22039,N_23310);
xnor U27077 (N_27077,N_23269,N_24810);
xnor U27078 (N_27078,N_22971,N_22805);
nand U27079 (N_27079,N_23431,N_22056);
or U27080 (N_27080,N_23184,N_24916);
or U27081 (N_27081,N_20430,N_20563);
and U27082 (N_27082,N_22126,N_20102);
xnor U27083 (N_27083,N_20368,N_22123);
or U27084 (N_27084,N_22916,N_22309);
nor U27085 (N_27085,N_20306,N_23955);
nor U27086 (N_27086,N_23972,N_22333);
or U27087 (N_27087,N_21994,N_24673);
or U27088 (N_27088,N_22679,N_22336);
xor U27089 (N_27089,N_24330,N_21327);
nor U27090 (N_27090,N_21679,N_24782);
nand U27091 (N_27091,N_20230,N_20638);
or U27092 (N_27092,N_23673,N_20694);
nor U27093 (N_27093,N_20275,N_22315);
nor U27094 (N_27094,N_22192,N_20491);
or U27095 (N_27095,N_24059,N_20939);
and U27096 (N_27096,N_20125,N_20332);
and U27097 (N_27097,N_23733,N_22569);
nor U27098 (N_27098,N_23785,N_23477);
nand U27099 (N_27099,N_20370,N_23080);
nor U27100 (N_27100,N_24649,N_23873);
and U27101 (N_27101,N_24298,N_22059);
or U27102 (N_27102,N_23490,N_20222);
or U27103 (N_27103,N_23107,N_23727);
xnor U27104 (N_27104,N_24152,N_22604);
nor U27105 (N_27105,N_22518,N_22201);
and U27106 (N_27106,N_24245,N_20296);
nor U27107 (N_27107,N_20123,N_24669);
or U27108 (N_27108,N_21132,N_24265);
or U27109 (N_27109,N_21734,N_23728);
and U27110 (N_27110,N_22356,N_20952);
xnor U27111 (N_27111,N_22430,N_24394);
and U27112 (N_27112,N_22026,N_20485);
nor U27113 (N_27113,N_22271,N_22936);
nor U27114 (N_27114,N_20435,N_22041);
or U27115 (N_27115,N_21515,N_23225);
xor U27116 (N_27116,N_24124,N_20259);
nand U27117 (N_27117,N_22266,N_20226);
nand U27118 (N_27118,N_20542,N_20502);
or U27119 (N_27119,N_23979,N_23010);
xnor U27120 (N_27120,N_24412,N_21420);
nand U27121 (N_27121,N_24944,N_21574);
and U27122 (N_27122,N_24621,N_22378);
or U27123 (N_27123,N_21723,N_20093);
or U27124 (N_27124,N_24532,N_24002);
and U27125 (N_27125,N_24314,N_23551);
and U27126 (N_27126,N_20604,N_22064);
or U27127 (N_27127,N_21733,N_22648);
nor U27128 (N_27128,N_23901,N_23975);
or U27129 (N_27129,N_23360,N_20301);
or U27130 (N_27130,N_24328,N_22528);
nor U27131 (N_27131,N_23072,N_20155);
or U27132 (N_27132,N_20817,N_20554);
nor U27133 (N_27133,N_24739,N_22484);
nand U27134 (N_27134,N_20118,N_24631);
nand U27135 (N_27135,N_21210,N_23793);
and U27136 (N_27136,N_21670,N_22804);
or U27137 (N_27137,N_24360,N_22188);
and U27138 (N_27138,N_20973,N_21919);
nor U27139 (N_27139,N_22156,N_21446);
nand U27140 (N_27140,N_21059,N_24758);
nor U27141 (N_27141,N_23252,N_24465);
or U27142 (N_27142,N_21164,N_20133);
nor U27143 (N_27143,N_24994,N_23216);
nor U27144 (N_27144,N_20714,N_24371);
and U27145 (N_27145,N_22762,N_22897);
or U27146 (N_27146,N_21321,N_20982);
xnor U27147 (N_27147,N_22352,N_22521);
nor U27148 (N_27148,N_23068,N_23091);
nand U27149 (N_27149,N_24697,N_21803);
and U27150 (N_27150,N_22142,N_24425);
or U27151 (N_27151,N_22417,N_22667);
and U27152 (N_27152,N_23108,N_24165);
or U27153 (N_27153,N_21972,N_24833);
nand U27154 (N_27154,N_23923,N_24415);
nor U27155 (N_27155,N_21323,N_21425);
nand U27156 (N_27156,N_21644,N_24433);
or U27157 (N_27157,N_24430,N_20799);
xnor U27158 (N_27158,N_22067,N_21213);
and U27159 (N_27159,N_24232,N_21692);
and U27160 (N_27160,N_22355,N_23012);
xnor U27161 (N_27161,N_21589,N_24800);
and U27162 (N_27162,N_20436,N_20342);
and U27163 (N_27163,N_24865,N_21725);
nand U27164 (N_27164,N_22270,N_23773);
nor U27165 (N_27165,N_23913,N_21754);
and U27166 (N_27166,N_22889,N_20162);
nor U27167 (N_27167,N_22803,N_23628);
nand U27168 (N_27168,N_23112,N_21611);
xnor U27169 (N_27169,N_23860,N_20494);
xor U27170 (N_27170,N_20887,N_23308);
nand U27171 (N_27171,N_20751,N_21510);
nor U27172 (N_27172,N_20000,N_24990);
and U27173 (N_27173,N_23555,N_20819);
nor U27174 (N_27174,N_22451,N_20595);
nand U27175 (N_27175,N_21979,N_24858);
and U27176 (N_27176,N_24907,N_20792);
xor U27177 (N_27177,N_24187,N_22675);
or U27178 (N_27178,N_23143,N_21386);
and U27179 (N_27179,N_24682,N_21513);
nand U27180 (N_27180,N_22374,N_24573);
nor U27181 (N_27181,N_23917,N_23021);
nand U27182 (N_27182,N_21688,N_23061);
and U27183 (N_27183,N_22585,N_24942);
and U27184 (N_27184,N_21790,N_22044);
and U27185 (N_27185,N_23538,N_24799);
or U27186 (N_27186,N_21637,N_22116);
nor U27187 (N_27187,N_22496,N_22466);
and U27188 (N_27188,N_22062,N_20009);
nand U27189 (N_27189,N_24016,N_24903);
or U27190 (N_27190,N_21671,N_21699);
and U27191 (N_27191,N_24586,N_22205);
or U27192 (N_27192,N_24836,N_21042);
or U27193 (N_27193,N_24535,N_21538);
or U27194 (N_27194,N_22940,N_21007);
or U27195 (N_27195,N_22913,N_21944);
nor U27196 (N_27196,N_23546,N_21721);
xor U27197 (N_27197,N_23369,N_20650);
nor U27198 (N_27198,N_21839,N_21479);
and U27199 (N_27199,N_21941,N_22301);
xor U27200 (N_27200,N_24166,N_23303);
nor U27201 (N_27201,N_24339,N_23428);
or U27202 (N_27202,N_21396,N_21718);
nor U27203 (N_27203,N_21372,N_20823);
nand U27204 (N_27204,N_22619,N_23544);
or U27205 (N_27205,N_23743,N_23476);
and U27206 (N_27206,N_24426,N_20724);
nor U27207 (N_27207,N_21899,N_22392);
and U27208 (N_27208,N_22233,N_24705);
or U27209 (N_27209,N_23603,N_21992);
or U27210 (N_27210,N_24280,N_24867);
nand U27211 (N_27211,N_23714,N_23319);
nor U27212 (N_27212,N_20122,N_21623);
or U27213 (N_27213,N_23508,N_21492);
or U27214 (N_27214,N_24146,N_24988);
nor U27215 (N_27215,N_20543,N_21128);
nor U27216 (N_27216,N_21114,N_24143);
xnor U27217 (N_27217,N_24242,N_24226);
and U27218 (N_27218,N_22842,N_20699);
nand U27219 (N_27219,N_20384,N_24854);
and U27220 (N_27220,N_21738,N_21827);
and U27221 (N_27221,N_21833,N_23907);
nor U27222 (N_27222,N_24248,N_22537);
nor U27223 (N_27223,N_22956,N_22575);
nand U27224 (N_27224,N_22737,N_22752);
nor U27225 (N_27225,N_21246,N_22345);
nand U27226 (N_27226,N_24273,N_23621);
nor U27227 (N_27227,N_24507,N_24386);
or U27228 (N_27228,N_20366,N_24198);
or U27229 (N_27229,N_21276,N_20618);
xor U27230 (N_27230,N_21951,N_20328);
or U27231 (N_27231,N_23838,N_21907);
nor U27232 (N_27232,N_20958,N_21970);
nand U27233 (N_27233,N_24428,N_24696);
nand U27234 (N_27234,N_23036,N_24707);
nand U27235 (N_27235,N_23553,N_21938);
and U27236 (N_27236,N_23891,N_20256);
and U27237 (N_27237,N_21127,N_22077);
nand U27238 (N_27238,N_23890,N_20271);
nand U27239 (N_27239,N_22625,N_21834);
nor U27240 (N_27240,N_24389,N_23597);
nand U27241 (N_27241,N_24257,N_23709);
nand U27242 (N_27242,N_24383,N_22439);
or U27243 (N_27243,N_22359,N_22138);
xnor U27244 (N_27244,N_22491,N_24698);
or U27245 (N_27245,N_23038,N_20423);
xnor U27246 (N_27246,N_24834,N_24050);
xnor U27247 (N_27247,N_21842,N_23074);
xor U27248 (N_27248,N_22945,N_24450);
or U27249 (N_27249,N_23580,N_24193);
and U27250 (N_27250,N_23958,N_21663);
xnor U27251 (N_27251,N_23370,N_23353);
nand U27252 (N_27252,N_22066,N_22183);
nor U27253 (N_27253,N_24794,N_23992);
nor U27254 (N_27254,N_23117,N_20045);
nor U27255 (N_27255,N_22412,N_23774);
xor U27256 (N_27256,N_24118,N_23876);
and U27257 (N_27257,N_24583,N_20185);
nand U27258 (N_27258,N_21965,N_22610);
nor U27259 (N_27259,N_22654,N_20861);
or U27260 (N_27260,N_22855,N_24238);
and U27261 (N_27261,N_23557,N_24932);
nor U27262 (N_27262,N_24755,N_24960);
nand U27263 (N_27263,N_21112,N_24989);
nor U27264 (N_27264,N_21376,N_21437);
or U27265 (N_27265,N_23070,N_24021);
and U27266 (N_27266,N_24154,N_21559);
xor U27267 (N_27267,N_20976,N_22224);
and U27268 (N_27268,N_21824,N_23174);
nor U27269 (N_27269,N_23833,N_22177);
nand U27270 (N_27270,N_24064,N_20251);
nand U27271 (N_27271,N_20832,N_20113);
nor U27272 (N_27272,N_22111,N_20622);
xnor U27273 (N_27273,N_21170,N_23136);
xor U27274 (N_27274,N_22416,N_24277);
nor U27275 (N_27275,N_23441,N_22324);
nor U27276 (N_27276,N_22761,N_23856);
and U27277 (N_27277,N_20347,N_20262);
or U27278 (N_27278,N_24652,N_21197);
and U27279 (N_27279,N_22789,N_20890);
or U27280 (N_27280,N_21998,N_24084);
xor U27281 (N_27281,N_23345,N_20305);
or U27282 (N_27282,N_23513,N_20706);
or U27283 (N_27283,N_22239,N_20091);
nand U27284 (N_27284,N_22841,N_23648);
and U27285 (N_27285,N_24101,N_20569);
or U27286 (N_27286,N_21879,N_22015);
nand U27287 (N_27287,N_24144,N_22227);
nand U27288 (N_27288,N_22448,N_22287);
nor U27289 (N_27289,N_22474,N_20803);
nor U27290 (N_27290,N_22580,N_21266);
and U27291 (N_27291,N_21870,N_20088);
and U27292 (N_27292,N_21787,N_24775);
or U27293 (N_27293,N_21247,N_23135);
or U27294 (N_27294,N_21142,N_23472);
nor U27295 (N_27295,N_24950,N_21601);
or U27296 (N_27296,N_23287,N_23514);
and U27297 (N_27297,N_20854,N_21275);
nand U27298 (N_27298,N_24251,N_23007);
and U27299 (N_27299,N_23478,N_21905);
or U27300 (N_27300,N_20119,N_22502);
and U27301 (N_27301,N_22994,N_22683);
xnor U27302 (N_27302,N_22078,N_23916);
nand U27303 (N_27303,N_22905,N_20352);
nor U27304 (N_27304,N_22952,N_22751);
nand U27305 (N_27305,N_21694,N_21272);
nor U27306 (N_27306,N_24564,N_24178);
or U27307 (N_27307,N_20922,N_21171);
xor U27308 (N_27308,N_23329,N_20017);
xor U27309 (N_27309,N_22924,N_20264);
and U27310 (N_27310,N_21065,N_22220);
nand U27311 (N_27311,N_23183,N_21209);
and U27312 (N_27312,N_24015,N_21901);
nor U27313 (N_27313,N_20524,N_21958);
and U27314 (N_27314,N_20428,N_21660);
and U27315 (N_27315,N_22694,N_21289);
and U27316 (N_27316,N_24656,N_22632);
xor U27317 (N_27317,N_21239,N_23790);
nand U27318 (N_27318,N_24225,N_21403);
and U27319 (N_27319,N_23256,N_21363);
and U27320 (N_27320,N_24563,N_22278);
and U27321 (N_27321,N_23368,N_20831);
or U27322 (N_27322,N_23150,N_24759);
or U27323 (N_27323,N_21956,N_23863);
nand U27324 (N_27324,N_24264,N_21558);
nand U27325 (N_27325,N_21050,N_24364);
and U27326 (N_27326,N_21579,N_23581);
and U27327 (N_27327,N_22663,N_22453);
and U27328 (N_27328,N_23028,N_22781);
and U27329 (N_27329,N_22449,N_20184);
nor U27330 (N_27330,N_24268,N_20372);
or U27331 (N_27331,N_23338,N_24472);
nor U27332 (N_27332,N_24842,N_20393);
nor U27333 (N_27333,N_20282,N_22137);
nand U27334 (N_27334,N_20183,N_20092);
nand U27335 (N_27335,N_21681,N_20925);
nor U27336 (N_27336,N_22759,N_22771);
or U27337 (N_27337,N_23357,N_24549);
and U27338 (N_27338,N_23608,N_23881);
and U27339 (N_27339,N_24683,N_20281);
and U27340 (N_27340,N_22478,N_21868);
nand U27341 (N_27341,N_24677,N_23294);
and U27342 (N_27342,N_22859,N_22700);
nand U27343 (N_27343,N_20058,N_23280);
nor U27344 (N_27344,N_24159,N_22411);
or U27345 (N_27345,N_20279,N_21424);
nor U27346 (N_27346,N_23547,N_23639);
nand U27347 (N_27347,N_22794,N_21711);
and U27348 (N_27348,N_24095,N_24285);
nand U27349 (N_27349,N_21109,N_24501);
or U27350 (N_27350,N_21706,N_20229);
nand U27351 (N_27351,N_20637,N_22592);
xnor U27352 (N_27352,N_20655,N_20752);
and U27353 (N_27353,N_20127,N_24828);
and U27354 (N_27354,N_22427,N_21101);
xnor U27355 (N_27355,N_20456,N_22058);
nand U27356 (N_27356,N_20556,N_21078);
nand U27357 (N_27357,N_24409,N_20024);
and U27358 (N_27358,N_21229,N_24476);
and U27359 (N_27359,N_22832,N_23464);
or U27360 (N_27360,N_24548,N_22687);
xnor U27361 (N_27361,N_21986,N_21008);
nand U27362 (N_27362,N_24419,N_23262);
and U27363 (N_27363,N_21249,N_22404);
nor U27364 (N_27364,N_22541,N_20753);
nor U27365 (N_27365,N_21017,N_21511);
nor U27366 (N_27366,N_24566,N_20717);
nand U27367 (N_27367,N_23929,N_24092);
nand U27368 (N_27368,N_20495,N_23447);
and U27369 (N_27369,N_23877,N_24447);
and U27370 (N_27370,N_24879,N_24255);
or U27371 (N_27371,N_22294,N_20664);
xnor U27372 (N_27372,N_21055,N_20021);
nand U27373 (N_27373,N_20216,N_23859);
nand U27374 (N_27374,N_23114,N_23846);
xor U27375 (N_27375,N_21573,N_21450);
or U27376 (N_27376,N_23291,N_21939);
and U27377 (N_27377,N_24760,N_20105);
nand U27378 (N_27378,N_20497,N_21722);
or U27379 (N_27379,N_20318,N_22813);
nand U27380 (N_27380,N_21407,N_24633);
or U27381 (N_27381,N_23349,N_23775);
and U27382 (N_27382,N_23912,N_20931);
nor U27383 (N_27383,N_23355,N_24499);
or U27384 (N_27384,N_22468,N_21231);
nand U27385 (N_27385,N_21620,N_21140);
nor U27386 (N_27386,N_24537,N_23406);
nand U27387 (N_27387,N_22958,N_21485);
and U27388 (N_27388,N_23206,N_20197);
nor U27389 (N_27389,N_24873,N_23421);
nor U27390 (N_27390,N_21820,N_24180);
or U27391 (N_27391,N_23971,N_24894);
nand U27392 (N_27392,N_21314,N_23230);
nand U27393 (N_27393,N_24534,N_22954);
nor U27394 (N_27394,N_21818,N_21525);
and U27395 (N_27395,N_21250,N_23647);
nor U27396 (N_27396,N_24921,N_20870);
nand U27397 (N_27397,N_20433,N_20927);
nor U27398 (N_27398,N_22014,N_20679);
or U27399 (N_27399,N_20888,N_20623);
or U27400 (N_27400,N_21512,N_24943);
nand U27401 (N_27401,N_23909,N_21264);
nand U27402 (N_27402,N_21845,N_20154);
or U27403 (N_27403,N_21566,N_24975);
nor U27404 (N_27404,N_21841,N_24058);
nand U27405 (N_27405,N_20583,N_20737);
and U27406 (N_27406,N_21920,N_22542);
or U27407 (N_27407,N_24071,N_23845);
nand U27408 (N_27408,N_22218,N_20757);
nand U27409 (N_27409,N_24581,N_23798);
nor U27410 (N_27410,N_23129,N_21639);
and U27411 (N_27411,N_24592,N_21470);
nand U27412 (N_27412,N_21964,N_21864);
nor U27413 (N_27413,N_20978,N_21341);
nand U27414 (N_27414,N_21607,N_21960);
or U27415 (N_27415,N_20944,N_23176);
xnor U27416 (N_27416,N_23284,N_20269);
xnor U27417 (N_27417,N_22614,N_20444);
nor U27418 (N_27418,N_20356,N_22214);
nor U27419 (N_27419,N_23543,N_24345);
nor U27420 (N_27420,N_22559,N_20121);
xnor U27421 (N_27421,N_22647,N_22682);
nor U27422 (N_27422,N_21358,N_21201);
or U27423 (N_27423,N_21338,N_21237);
nor U27424 (N_27424,N_23336,N_22930);
and U27425 (N_27425,N_23453,N_22086);
xnor U27426 (N_27426,N_21225,N_21984);
nor U27427 (N_27427,N_24316,N_23471);
nand U27428 (N_27428,N_20080,N_21411);
nand U27429 (N_27429,N_22281,N_20437);
nor U27430 (N_27430,N_24133,N_21891);
nand U27431 (N_27431,N_22370,N_22791);
xnor U27432 (N_27432,N_24912,N_23802);
nand U27433 (N_27433,N_22643,N_20954);
nand U27434 (N_27434,N_22380,N_24695);
and U27435 (N_27435,N_21316,N_21312);
or U27436 (N_27436,N_23631,N_21713);
or U27437 (N_27437,N_23311,N_20899);
and U27438 (N_27438,N_20601,N_23882);
nand U27439 (N_27439,N_23398,N_20465);
nand U27440 (N_27440,N_20961,N_24263);
and U27441 (N_27441,N_24173,N_23209);
nor U27442 (N_27442,N_22951,N_24184);
and U27443 (N_27443,N_24664,N_24055);
nor U27444 (N_27444,N_21451,N_23335);
nor U27445 (N_27445,N_21828,N_23304);
or U27446 (N_27446,N_21522,N_24151);
nor U27447 (N_27447,N_22998,N_20681);
and U27448 (N_27448,N_21551,N_22834);
nand U27449 (N_27449,N_24176,N_23384);
nor U27450 (N_27450,N_22028,N_23843);
xor U27451 (N_27451,N_22902,N_21550);
or U27452 (N_27452,N_24100,N_22501);
or U27453 (N_27453,N_23201,N_21917);
nand U27454 (N_27454,N_20579,N_22948);
or U27455 (N_27455,N_23554,N_22276);
nand U27456 (N_27456,N_22203,N_22579);
and U27457 (N_27457,N_21381,N_22538);
or U27458 (N_27458,N_24736,N_24965);
xnor U27459 (N_27459,N_20150,N_22120);
nor U27460 (N_27460,N_22915,N_22054);
nor U27461 (N_27461,N_24771,N_24048);
nand U27462 (N_27462,N_23707,N_22581);
nor U27463 (N_27463,N_20472,N_21609);
nand U27464 (N_27464,N_24958,N_21704);
nand U27465 (N_27465,N_20339,N_24227);
nor U27466 (N_27466,N_24593,N_24546);
or U27467 (N_27467,N_21825,N_23498);
nand U27468 (N_27468,N_23670,N_22529);
and U27469 (N_27469,N_24686,N_23897);
nand U27470 (N_27470,N_23944,N_20950);
and U27471 (N_27471,N_20065,N_21698);
nand U27472 (N_27472,N_21090,N_24731);
xor U27473 (N_27473,N_23865,N_20500);
and U27474 (N_27474,N_23302,N_20201);
xnor U27475 (N_27475,N_21780,N_24126);
nand U27476 (N_27476,N_22389,N_22596);
and U27477 (N_27477,N_24729,N_23314);
nor U27478 (N_27478,N_21167,N_24040);
xnor U27479 (N_27479,N_21252,N_24787);
or U27480 (N_27480,N_23432,N_20913);
and U27481 (N_27481,N_20478,N_20661);
nor U27482 (N_27482,N_24281,N_21527);
nand U27483 (N_27483,N_21874,N_24141);
nand U27484 (N_27484,N_21548,N_20644);
and U27485 (N_27485,N_22674,N_22040);
and U27486 (N_27486,N_22543,N_23082);
xnor U27487 (N_27487,N_21968,N_23210);
or U27488 (N_27488,N_23609,N_21279);
and U27489 (N_27489,N_20993,N_24001);
or U27490 (N_27490,N_20877,N_21318);
xnor U27491 (N_27491,N_23315,N_20173);
nand U27492 (N_27492,N_22150,N_22360);
xnor U27493 (N_27493,N_24478,N_20945);
nand U27494 (N_27494,N_24718,N_23984);
nand U27495 (N_27495,N_22435,N_21203);
or U27496 (N_27496,N_21141,N_22034);
nor U27497 (N_27497,N_20672,N_24142);
nand U27498 (N_27498,N_20061,N_20692);
or U27499 (N_27499,N_22967,N_20858);
or U27500 (N_27500,N_23022,N_20049);
xor U27501 (N_27501,N_23024,N_20279);
xnor U27502 (N_27502,N_22723,N_23641);
nand U27503 (N_27503,N_21471,N_24866);
nor U27504 (N_27504,N_20601,N_24725);
and U27505 (N_27505,N_22192,N_20445);
and U27506 (N_27506,N_21933,N_24410);
xnor U27507 (N_27507,N_21228,N_24950);
nand U27508 (N_27508,N_21816,N_20289);
or U27509 (N_27509,N_20510,N_20887);
nor U27510 (N_27510,N_23683,N_20554);
nor U27511 (N_27511,N_23068,N_23789);
and U27512 (N_27512,N_21367,N_22268);
xor U27513 (N_27513,N_23027,N_21904);
nor U27514 (N_27514,N_24941,N_23649);
or U27515 (N_27515,N_20359,N_20512);
or U27516 (N_27516,N_24108,N_24627);
and U27517 (N_27517,N_22278,N_22650);
nor U27518 (N_27518,N_24918,N_21645);
and U27519 (N_27519,N_23453,N_23992);
and U27520 (N_27520,N_24327,N_23889);
and U27521 (N_27521,N_20487,N_22624);
xnor U27522 (N_27522,N_22414,N_21662);
or U27523 (N_27523,N_20291,N_23592);
and U27524 (N_27524,N_22275,N_21366);
and U27525 (N_27525,N_22316,N_23904);
or U27526 (N_27526,N_24840,N_23871);
nand U27527 (N_27527,N_21281,N_20165);
and U27528 (N_27528,N_23251,N_22797);
nor U27529 (N_27529,N_22823,N_23246);
nor U27530 (N_27530,N_20893,N_20612);
or U27531 (N_27531,N_23825,N_20292);
and U27532 (N_27532,N_21906,N_24269);
nor U27533 (N_27533,N_21434,N_24497);
and U27534 (N_27534,N_20516,N_24352);
nand U27535 (N_27535,N_23548,N_24480);
nor U27536 (N_27536,N_22546,N_22116);
or U27537 (N_27537,N_20596,N_20661);
or U27538 (N_27538,N_21918,N_22719);
or U27539 (N_27539,N_20960,N_23716);
xnor U27540 (N_27540,N_24748,N_22064);
and U27541 (N_27541,N_24478,N_23468);
or U27542 (N_27542,N_20874,N_24031);
and U27543 (N_27543,N_22402,N_23545);
nor U27544 (N_27544,N_23798,N_23566);
nand U27545 (N_27545,N_24249,N_22091);
xnor U27546 (N_27546,N_21487,N_20013);
nor U27547 (N_27547,N_23927,N_24844);
and U27548 (N_27548,N_23048,N_21785);
nand U27549 (N_27549,N_24506,N_20377);
xnor U27550 (N_27550,N_21608,N_22763);
xnor U27551 (N_27551,N_20587,N_20328);
or U27552 (N_27552,N_21403,N_21353);
nand U27553 (N_27553,N_22251,N_21696);
nor U27554 (N_27554,N_21088,N_21557);
nor U27555 (N_27555,N_21942,N_20940);
or U27556 (N_27556,N_22758,N_24396);
and U27557 (N_27557,N_24893,N_20939);
nand U27558 (N_27558,N_23660,N_22962);
and U27559 (N_27559,N_24450,N_20505);
and U27560 (N_27560,N_24002,N_23950);
xnor U27561 (N_27561,N_23268,N_21548);
or U27562 (N_27562,N_23041,N_24711);
nand U27563 (N_27563,N_24133,N_20270);
and U27564 (N_27564,N_24977,N_24957);
nor U27565 (N_27565,N_21968,N_20002);
xnor U27566 (N_27566,N_22671,N_24156);
and U27567 (N_27567,N_20940,N_24895);
or U27568 (N_27568,N_24158,N_24296);
xnor U27569 (N_27569,N_23065,N_22225);
nor U27570 (N_27570,N_21171,N_21056);
or U27571 (N_27571,N_22542,N_22042);
or U27572 (N_27572,N_24372,N_23040);
nand U27573 (N_27573,N_20371,N_21276);
xnor U27574 (N_27574,N_24475,N_21625);
and U27575 (N_27575,N_20122,N_22514);
nand U27576 (N_27576,N_21888,N_21480);
and U27577 (N_27577,N_24390,N_21999);
or U27578 (N_27578,N_23427,N_23209);
or U27579 (N_27579,N_23135,N_22320);
nand U27580 (N_27580,N_22067,N_22582);
or U27581 (N_27581,N_21784,N_22916);
or U27582 (N_27582,N_24215,N_22528);
and U27583 (N_27583,N_22832,N_20448);
and U27584 (N_27584,N_23493,N_23947);
nor U27585 (N_27585,N_20877,N_23142);
nand U27586 (N_27586,N_22577,N_23468);
xnor U27587 (N_27587,N_22639,N_24276);
or U27588 (N_27588,N_21100,N_20454);
nor U27589 (N_27589,N_20257,N_23241);
nand U27590 (N_27590,N_20966,N_23108);
nand U27591 (N_27591,N_20965,N_21740);
nor U27592 (N_27592,N_21060,N_23460);
nand U27593 (N_27593,N_20177,N_23021);
nand U27594 (N_27594,N_22892,N_24390);
nand U27595 (N_27595,N_23491,N_23401);
and U27596 (N_27596,N_21596,N_20003);
or U27597 (N_27597,N_24944,N_20981);
nand U27598 (N_27598,N_22575,N_21884);
nand U27599 (N_27599,N_23533,N_23055);
or U27600 (N_27600,N_22565,N_20673);
and U27601 (N_27601,N_21194,N_20459);
xnor U27602 (N_27602,N_23670,N_23506);
nor U27603 (N_27603,N_23323,N_24579);
nor U27604 (N_27604,N_23423,N_23111);
xnor U27605 (N_27605,N_21038,N_22296);
and U27606 (N_27606,N_22400,N_24407);
nor U27607 (N_27607,N_23899,N_22910);
nor U27608 (N_27608,N_20080,N_20524);
and U27609 (N_27609,N_24883,N_21530);
nor U27610 (N_27610,N_24460,N_24121);
or U27611 (N_27611,N_20764,N_21530);
xor U27612 (N_27612,N_24917,N_24623);
nand U27613 (N_27613,N_23643,N_21443);
nor U27614 (N_27614,N_22430,N_22655);
or U27615 (N_27615,N_21069,N_21323);
nor U27616 (N_27616,N_22364,N_23750);
nand U27617 (N_27617,N_20907,N_23139);
and U27618 (N_27618,N_21850,N_24371);
nor U27619 (N_27619,N_20975,N_20752);
xor U27620 (N_27620,N_22688,N_20868);
nand U27621 (N_27621,N_22460,N_23298);
nor U27622 (N_27622,N_20988,N_23725);
xnor U27623 (N_27623,N_20188,N_22480);
nand U27624 (N_27624,N_20152,N_21739);
and U27625 (N_27625,N_22896,N_22072);
nor U27626 (N_27626,N_23979,N_23868);
and U27627 (N_27627,N_24659,N_20173);
and U27628 (N_27628,N_21641,N_21409);
or U27629 (N_27629,N_22367,N_21610);
and U27630 (N_27630,N_22268,N_22284);
and U27631 (N_27631,N_20035,N_20847);
xor U27632 (N_27632,N_24462,N_23698);
or U27633 (N_27633,N_20571,N_20147);
xnor U27634 (N_27634,N_24982,N_21050);
nor U27635 (N_27635,N_23604,N_23237);
and U27636 (N_27636,N_22051,N_22915);
nand U27637 (N_27637,N_24788,N_24577);
and U27638 (N_27638,N_21007,N_20664);
nand U27639 (N_27639,N_22120,N_22075);
nand U27640 (N_27640,N_20572,N_22042);
nor U27641 (N_27641,N_20218,N_24211);
or U27642 (N_27642,N_21816,N_23137);
nor U27643 (N_27643,N_23480,N_23604);
and U27644 (N_27644,N_23405,N_24693);
nor U27645 (N_27645,N_23786,N_22080);
nand U27646 (N_27646,N_21229,N_23582);
and U27647 (N_27647,N_24342,N_20343);
or U27648 (N_27648,N_21636,N_24917);
nand U27649 (N_27649,N_21819,N_22598);
nand U27650 (N_27650,N_22591,N_24376);
or U27651 (N_27651,N_20961,N_23153);
or U27652 (N_27652,N_21614,N_24935);
and U27653 (N_27653,N_21875,N_20521);
or U27654 (N_27654,N_23882,N_23767);
xnor U27655 (N_27655,N_21023,N_22040);
and U27656 (N_27656,N_21281,N_22876);
xor U27657 (N_27657,N_23535,N_20898);
and U27658 (N_27658,N_23194,N_22260);
xnor U27659 (N_27659,N_20314,N_23287);
and U27660 (N_27660,N_23937,N_24395);
nand U27661 (N_27661,N_24856,N_23451);
nor U27662 (N_27662,N_21368,N_20554);
or U27663 (N_27663,N_24797,N_20777);
xor U27664 (N_27664,N_23406,N_22277);
nand U27665 (N_27665,N_22773,N_22653);
and U27666 (N_27666,N_23721,N_22804);
or U27667 (N_27667,N_22342,N_20363);
or U27668 (N_27668,N_20685,N_21117);
nand U27669 (N_27669,N_21811,N_23118);
or U27670 (N_27670,N_21151,N_20662);
and U27671 (N_27671,N_24590,N_20862);
nor U27672 (N_27672,N_24659,N_24768);
nand U27673 (N_27673,N_22192,N_22690);
or U27674 (N_27674,N_20780,N_22598);
and U27675 (N_27675,N_22453,N_23776);
and U27676 (N_27676,N_21785,N_24920);
nor U27677 (N_27677,N_24427,N_24443);
and U27678 (N_27678,N_20076,N_22782);
or U27679 (N_27679,N_20440,N_23780);
nor U27680 (N_27680,N_21834,N_23171);
nor U27681 (N_27681,N_21346,N_24592);
nand U27682 (N_27682,N_24078,N_22003);
or U27683 (N_27683,N_21531,N_21890);
nand U27684 (N_27684,N_22175,N_23968);
nand U27685 (N_27685,N_24897,N_22004);
nor U27686 (N_27686,N_22964,N_21189);
and U27687 (N_27687,N_20574,N_21363);
nand U27688 (N_27688,N_22465,N_21608);
or U27689 (N_27689,N_23982,N_21323);
nor U27690 (N_27690,N_22398,N_21138);
or U27691 (N_27691,N_20002,N_24358);
nor U27692 (N_27692,N_24840,N_20258);
nor U27693 (N_27693,N_23460,N_21448);
nand U27694 (N_27694,N_21201,N_22063);
and U27695 (N_27695,N_20890,N_24620);
nand U27696 (N_27696,N_23274,N_21462);
xnor U27697 (N_27697,N_21870,N_24377);
nor U27698 (N_27698,N_21832,N_24448);
and U27699 (N_27699,N_21068,N_20403);
xnor U27700 (N_27700,N_20461,N_24719);
nand U27701 (N_27701,N_20579,N_23185);
xnor U27702 (N_27702,N_23710,N_21283);
or U27703 (N_27703,N_24796,N_21682);
and U27704 (N_27704,N_22810,N_24756);
nor U27705 (N_27705,N_21865,N_22563);
nor U27706 (N_27706,N_21262,N_20316);
xnor U27707 (N_27707,N_24503,N_20824);
nor U27708 (N_27708,N_21761,N_21134);
and U27709 (N_27709,N_21346,N_24102);
nand U27710 (N_27710,N_22112,N_24088);
and U27711 (N_27711,N_22468,N_22845);
xnor U27712 (N_27712,N_22471,N_21670);
xnor U27713 (N_27713,N_22629,N_23600);
nand U27714 (N_27714,N_21715,N_24155);
nor U27715 (N_27715,N_24542,N_23452);
or U27716 (N_27716,N_24529,N_20407);
and U27717 (N_27717,N_22940,N_20896);
xnor U27718 (N_27718,N_24785,N_20287);
nor U27719 (N_27719,N_23580,N_23792);
nor U27720 (N_27720,N_24591,N_24153);
nand U27721 (N_27721,N_21760,N_22489);
nand U27722 (N_27722,N_20583,N_24285);
and U27723 (N_27723,N_24018,N_24743);
nor U27724 (N_27724,N_22819,N_24386);
and U27725 (N_27725,N_22629,N_22231);
nor U27726 (N_27726,N_21148,N_22464);
nor U27727 (N_27727,N_21723,N_20262);
nand U27728 (N_27728,N_20260,N_23281);
nand U27729 (N_27729,N_22419,N_20437);
nand U27730 (N_27730,N_22300,N_20562);
or U27731 (N_27731,N_24804,N_23507);
or U27732 (N_27732,N_20549,N_23920);
nor U27733 (N_27733,N_20778,N_24615);
nand U27734 (N_27734,N_20584,N_21050);
or U27735 (N_27735,N_23437,N_22617);
and U27736 (N_27736,N_24873,N_22197);
or U27737 (N_27737,N_21556,N_24112);
xnor U27738 (N_27738,N_23902,N_20585);
nor U27739 (N_27739,N_21369,N_22406);
or U27740 (N_27740,N_23114,N_23042);
or U27741 (N_27741,N_24208,N_20989);
or U27742 (N_27742,N_23217,N_23533);
or U27743 (N_27743,N_22905,N_21235);
or U27744 (N_27744,N_22701,N_21284);
nand U27745 (N_27745,N_24935,N_20825);
nor U27746 (N_27746,N_21111,N_22457);
nand U27747 (N_27747,N_22621,N_22063);
xor U27748 (N_27748,N_22883,N_22237);
xor U27749 (N_27749,N_22331,N_21150);
nand U27750 (N_27750,N_23331,N_23526);
nor U27751 (N_27751,N_22330,N_20216);
and U27752 (N_27752,N_21924,N_21724);
and U27753 (N_27753,N_23260,N_24956);
nand U27754 (N_27754,N_20864,N_20716);
nand U27755 (N_27755,N_20926,N_23941);
or U27756 (N_27756,N_21046,N_22774);
and U27757 (N_27757,N_23930,N_22006);
nand U27758 (N_27758,N_24072,N_21271);
nand U27759 (N_27759,N_23034,N_21249);
nor U27760 (N_27760,N_23140,N_21821);
nor U27761 (N_27761,N_22987,N_24462);
or U27762 (N_27762,N_20220,N_21694);
or U27763 (N_27763,N_21364,N_24425);
nand U27764 (N_27764,N_21982,N_21168);
or U27765 (N_27765,N_23588,N_24119);
nand U27766 (N_27766,N_22028,N_22383);
and U27767 (N_27767,N_22043,N_21344);
nor U27768 (N_27768,N_23153,N_23463);
and U27769 (N_27769,N_23638,N_23247);
nand U27770 (N_27770,N_21829,N_24770);
nor U27771 (N_27771,N_20229,N_20672);
and U27772 (N_27772,N_24383,N_21433);
nand U27773 (N_27773,N_21333,N_24125);
nor U27774 (N_27774,N_20625,N_23740);
nor U27775 (N_27775,N_23020,N_21532);
and U27776 (N_27776,N_20288,N_24934);
nand U27777 (N_27777,N_23672,N_24350);
nand U27778 (N_27778,N_23171,N_20910);
nor U27779 (N_27779,N_24780,N_23982);
or U27780 (N_27780,N_21924,N_23268);
or U27781 (N_27781,N_20955,N_21167);
and U27782 (N_27782,N_22530,N_24300);
nor U27783 (N_27783,N_24845,N_21436);
or U27784 (N_27784,N_22167,N_22522);
nand U27785 (N_27785,N_23390,N_22236);
nand U27786 (N_27786,N_24983,N_24073);
or U27787 (N_27787,N_20517,N_22944);
nand U27788 (N_27788,N_24603,N_23770);
or U27789 (N_27789,N_24808,N_21230);
xnor U27790 (N_27790,N_21400,N_20693);
nand U27791 (N_27791,N_24434,N_20241);
xor U27792 (N_27792,N_24080,N_21141);
or U27793 (N_27793,N_24911,N_21543);
xnor U27794 (N_27794,N_24127,N_20811);
and U27795 (N_27795,N_23365,N_23514);
xor U27796 (N_27796,N_20586,N_24568);
nand U27797 (N_27797,N_23774,N_23796);
nor U27798 (N_27798,N_24155,N_21623);
nor U27799 (N_27799,N_21163,N_22930);
nand U27800 (N_27800,N_21226,N_20706);
nor U27801 (N_27801,N_22235,N_21611);
nand U27802 (N_27802,N_22566,N_23222);
nand U27803 (N_27803,N_22274,N_23791);
nor U27804 (N_27804,N_20381,N_23090);
nor U27805 (N_27805,N_20723,N_24275);
nand U27806 (N_27806,N_22419,N_21878);
nor U27807 (N_27807,N_21693,N_22843);
nand U27808 (N_27808,N_24849,N_21131);
nor U27809 (N_27809,N_23469,N_21497);
or U27810 (N_27810,N_21238,N_24524);
nand U27811 (N_27811,N_23388,N_22544);
and U27812 (N_27812,N_24455,N_20702);
nor U27813 (N_27813,N_21067,N_23693);
nand U27814 (N_27814,N_21392,N_24081);
xor U27815 (N_27815,N_24628,N_20306);
or U27816 (N_27816,N_23543,N_20452);
or U27817 (N_27817,N_20703,N_21561);
or U27818 (N_27818,N_20453,N_22350);
nand U27819 (N_27819,N_23701,N_22226);
xnor U27820 (N_27820,N_21342,N_24646);
nand U27821 (N_27821,N_23224,N_21008);
nand U27822 (N_27822,N_21597,N_20585);
nand U27823 (N_27823,N_20132,N_21738);
xor U27824 (N_27824,N_20420,N_24106);
or U27825 (N_27825,N_23822,N_22077);
or U27826 (N_27826,N_22109,N_24405);
or U27827 (N_27827,N_21419,N_22454);
nand U27828 (N_27828,N_20656,N_20341);
or U27829 (N_27829,N_20515,N_20542);
nor U27830 (N_27830,N_21749,N_20827);
nor U27831 (N_27831,N_20345,N_21382);
nor U27832 (N_27832,N_24494,N_21777);
and U27833 (N_27833,N_22045,N_22085);
xnor U27834 (N_27834,N_23075,N_23153);
xor U27835 (N_27835,N_23000,N_20974);
and U27836 (N_27836,N_24639,N_20257);
or U27837 (N_27837,N_23728,N_21090);
xor U27838 (N_27838,N_21603,N_20900);
and U27839 (N_27839,N_22714,N_24283);
nand U27840 (N_27840,N_20109,N_23518);
or U27841 (N_27841,N_24789,N_22342);
nor U27842 (N_27842,N_23537,N_22356);
xor U27843 (N_27843,N_24771,N_22400);
or U27844 (N_27844,N_20785,N_24415);
and U27845 (N_27845,N_21522,N_20203);
xnor U27846 (N_27846,N_22817,N_21900);
nand U27847 (N_27847,N_24146,N_20862);
or U27848 (N_27848,N_24930,N_24099);
nor U27849 (N_27849,N_21046,N_22396);
nor U27850 (N_27850,N_20188,N_20466);
or U27851 (N_27851,N_22420,N_22787);
nor U27852 (N_27852,N_22110,N_24717);
nor U27853 (N_27853,N_21278,N_24902);
nor U27854 (N_27854,N_23522,N_21471);
or U27855 (N_27855,N_24388,N_22613);
nor U27856 (N_27856,N_20477,N_20408);
nor U27857 (N_27857,N_23356,N_23057);
nand U27858 (N_27858,N_22108,N_21338);
nand U27859 (N_27859,N_23884,N_24711);
nand U27860 (N_27860,N_22016,N_20224);
nand U27861 (N_27861,N_21031,N_24964);
nor U27862 (N_27862,N_20182,N_21971);
nor U27863 (N_27863,N_21115,N_23239);
xnor U27864 (N_27864,N_24981,N_22087);
nor U27865 (N_27865,N_21119,N_20587);
and U27866 (N_27866,N_21106,N_22762);
nand U27867 (N_27867,N_20774,N_20571);
nand U27868 (N_27868,N_20535,N_24962);
nand U27869 (N_27869,N_21464,N_21781);
and U27870 (N_27870,N_22397,N_21924);
or U27871 (N_27871,N_21748,N_23040);
and U27872 (N_27872,N_23759,N_22118);
or U27873 (N_27873,N_21325,N_21688);
or U27874 (N_27874,N_20806,N_24046);
and U27875 (N_27875,N_22398,N_21296);
nor U27876 (N_27876,N_22001,N_21466);
and U27877 (N_27877,N_22313,N_22896);
nand U27878 (N_27878,N_24844,N_23346);
or U27879 (N_27879,N_20990,N_23721);
and U27880 (N_27880,N_21101,N_22551);
and U27881 (N_27881,N_24383,N_24613);
xnor U27882 (N_27882,N_23279,N_21856);
nand U27883 (N_27883,N_23094,N_22420);
or U27884 (N_27884,N_23466,N_24527);
nand U27885 (N_27885,N_22821,N_24356);
nor U27886 (N_27886,N_24231,N_20284);
nand U27887 (N_27887,N_20289,N_20011);
nand U27888 (N_27888,N_24708,N_20197);
or U27889 (N_27889,N_23182,N_23080);
or U27890 (N_27890,N_20566,N_23000);
nand U27891 (N_27891,N_21179,N_23861);
xor U27892 (N_27892,N_22733,N_21080);
or U27893 (N_27893,N_20564,N_22799);
nand U27894 (N_27894,N_23281,N_23952);
xor U27895 (N_27895,N_22025,N_23727);
nor U27896 (N_27896,N_22256,N_22497);
nor U27897 (N_27897,N_22969,N_24115);
and U27898 (N_27898,N_22710,N_20482);
or U27899 (N_27899,N_22297,N_20792);
xnor U27900 (N_27900,N_20204,N_20098);
nand U27901 (N_27901,N_22412,N_24627);
and U27902 (N_27902,N_21628,N_23297);
and U27903 (N_27903,N_21936,N_21466);
nor U27904 (N_27904,N_23340,N_23775);
and U27905 (N_27905,N_21637,N_24896);
nor U27906 (N_27906,N_22970,N_20833);
nor U27907 (N_27907,N_23769,N_20978);
and U27908 (N_27908,N_20314,N_22303);
and U27909 (N_27909,N_20330,N_24314);
nor U27910 (N_27910,N_21587,N_24636);
or U27911 (N_27911,N_21439,N_22045);
or U27912 (N_27912,N_24469,N_22684);
or U27913 (N_27913,N_21333,N_22581);
xnor U27914 (N_27914,N_24193,N_22358);
and U27915 (N_27915,N_22587,N_23062);
nor U27916 (N_27916,N_20888,N_23481);
xor U27917 (N_27917,N_24102,N_24824);
nor U27918 (N_27918,N_21676,N_20730);
and U27919 (N_27919,N_22661,N_20232);
nor U27920 (N_27920,N_24332,N_21868);
nand U27921 (N_27921,N_22476,N_23400);
xnor U27922 (N_27922,N_23369,N_24602);
nor U27923 (N_27923,N_21308,N_22331);
and U27924 (N_27924,N_24440,N_24512);
nand U27925 (N_27925,N_22757,N_23730);
or U27926 (N_27926,N_23234,N_22055);
and U27927 (N_27927,N_24343,N_21244);
xor U27928 (N_27928,N_21656,N_23713);
nand U27929 (N_27929,N_24462,N_21796);
or U27930 (N_27930,N_21532,N_24253);
nor U27931 (N_27931,N_24957,N_20099);
nand U27932 (N_27932,N_21917,N_23205);
nand U27933 (N_27933,N_21763,N_21493);
nand U27934 (N_27934,N_23560,N_23593);
xnor U27935 (N_27935,N_23234,N_21456);
nand U27936 (N_27936,N_22305,N_24684);
and U27937 (N_27937,N_22038,N_21084);
or U27938 (N_27938,N_21309,N_24751);
nand U27939 (N_27939,N_20100,N_23815);
nor U27940 (N_27940,N_22223,N_22343);
and U27941 (N_27941,N_21405,N_20139);
nor U27942 (N_27942,N_21784,N_24743);
nand U27943 (N_27943,N_24579,N_24955);
or U27944 (N_27944,N_20901,N_20968);
nand U27945 (N_27945,N_23380,N_22531);
xor U27946 (N_27946,N_22562,N_22926);
nand U27947 (N_27947,N_22174,N_20126);
nand U27948 (N_27948,N_24785,N_24882);
nor U27949 (N_27949,N_20872,N_23984);
and U27950 (N_27950,N_24238,N_20634);
or U27951 (N_27951,N_24726,N_22020);
xor U27952 (N_27952,N_20118,N_24931);
or U27953 (N_27953,N_21382,N_23300);
nor U27954 (N_27954,N_20382,N_22879);
or U27955 (N_27955,N_20312,N_24800);
nand U27956 (N_27956,N_21009,N_21624);
and U27957 (N_27957,N_23174,N_24011);
xnor U27958 (N_27958,N_24698,N_22970);
nor U27959 (N_27959,N_22194,N_20462);
or U27960 (N_27960,N_22276,N_22594);
or U27961 (N_27961,N_22892,N_21800);
or U27962 (N_27962,N_21448,N_22613);
nand U27963 (N_27963,N_23559,N_21817);
nand U27964 (N_27964,N_21088,N_23867);
and U27965 (N_27965,N_23298,N_23817);
nand U27966 (N_27966,N_20984,N_21547);
or U27967 (N_27967,N_20947,N_22463);
nor U27968 (N_27968,N_22312,N_21225);
nor U27969 (N_27969,N_24996,N_23897);
or U27970 (N_27970,N_20473,N_23545);
nor U27971 (N_27971,N_21077,N_22641);
nor U27972 (N_27972,N_21775,N_21947);
nand U27973 (N_27973,N_22767,N_23620);
nand U27974 (N_27974,N_22496,N_20299);
xnor U27975 (N_27975,N_21980,N_20588);
xor U27976 (N_27976,N_22668,N_24284);
nand U27977 (N_27977,N_20869,N_22428);
nand U27978 (N_27978,N_20607,N_20933);
or U27979 (N_27979,N_24663,N_21260);
nor U27980 (N_27980,N_23253,N_22459);
nand U27981 (N_27981,N_21726,N_22115);
nand U27982 (N_27982,N_21305,N_24718);
nand U27983 (N_27983,N_23064,N_21547);
nor U27984 (N_27984,N_21111,N_22385);
or U27985 (N_27985,N_24948,N_22473);
or U27986 (N_27986,N_21665,N_21167);
nor U27987 (N_27987,N_20182,N_23214);
nand U27988 (N_27988,N_20268,N_24269);
and U27989 (N_27989,N_22683,N_21736);
xor U27990 (N_27990,N_24545,N_20953);
nor U27991 (N_27991,N_22251,N_23613);
and U27992 (N_27992,N_20020,N_21983);
and U27993 (N_27993,N_23951,N_21093);
nor U27994 (N_27994,N_20265,N_21303);
nand U27995 (N_27995,N_24341,N_22963);
nor U27996 (N_27996,N_20532,N_24593);
or U27997 (N_27997,N_23092,N_22646);
and U27998 (N_27998,N_22728,N_22525);
or U27999 (N_27999,N_21938,N_20144);
or U28000 (N_28000,N_22753,N_24122);
nor U28001 (N_28001,N_23153,N_22880);
nor U28002 (N_28002,N_22083,N_20734);
or U28003 (N_28003,N_22544,N_20626);
nor U28004 (N_28004,N_23061,N_23745);
nand U28005 (N_28005,N_22328,N_22977);
and U28006 (N_28006,N_24636,N_22837);
nand U28007 (N_28007,N_22297,N_22573);
and U28008 (N_28008,N_20393,N_23401);
or U28009 (N_28009,N_20692,N_22419);
nand U28010 (N_28010,N_23370,N_23203);
nand U28011 (N_28011,N_23680,N_24903);
or U28012 (N_28012,N_23771,N_22232);
or U28013 (N_28013,N_20417,N_24420);
nor U28014 (N_28014,N_22696,N_23580);
xor U28015 (N_28015,N_20435,N_24418);
nand U28016 (N_28016,N_20490,N_22131);
or U28017 (N_28017,N_20744,N_24789);
nor U28018 (N_28018,N_21946,N_23283);
nand U28019 (N_28019,N_24012,N_21079);
and U28020 (N_28020,N_24906,N_21682);
nand U28021 (N_28021,N_20242,N_21796);
or U28022 (N_28022,N_22939,N_23089);
and U28023 (N_28023,N_23093,N_22744);
or U28024 (N_28024,N_20446,N_22709);
xor U28025 (N_28025,N_24508,N_20094);
nor U28026 (N_28026,N_24735,N_21409);
and U28027 (N_28027,N_20471,N_23915);
nor U28028 (N_28028,N_23555,N_23987);
or U28029 (N_28029,N_23261,N_20438);
nor U28030 (N_28030,N_23969,N_24894);
nor U28031 (N_28031,N_21428,N_22859);
nor U28032 (N_28032,N_20625,N_20636);
nand U28033 (N_28033,N_20083,N_20006);
nor U28034 (N_28034,N_20132,N_21899);
xnor U28035 (N_28035,N_21724,N_23274);
nand U28036 (N_28036,N_20834,N_22041);
nand U28037 (N_28037,N_21456,N_21789);
or U28038 (N_28038,N_21080,N_20692);
nand U28039 (N_28039,N_24439,N_20335);
nand U28040 (N_28040,N_24097,N_20574);
nand U28041 (N_28041,N_21043,N_22784);
xnor U28042 (N_28042,N_20004,N_20932);
nor U28043 (N_28043,N_21818,N_20447);
and U28044 (N_28044,N_23793,N_22603);
or U28045 (N_28045,N_20798,N_24934);
nand U28046 (N_28046,N_22260,N_20100);
nor U28047 (N_28047,N_24775,N_21824);
or U28048 (N_28048,N_24214,N_22518);
or U28049 (N_28049,N_20996,N_23747);
nand U28050 (N_28050,N_22288,N_23984);
and U28051 (N_28051,N_23928,N_24741);
nor U28052 (N_28052,N_24456,N_21852);
and U28053 (N_28053,N_23457,N_23993);
or U28054 (N_28054,N_22990,N_20016);
nor U28055 (N_28055,N_21740,N_23014);
and U28056 (N_28056,N_22014,N_22267);
nor U28057 (N_28057,N_21141,N_24591);
nand U28058 (N_28058,N_21389,N_20571);
xnor U28059 (N_28059,N_20037,N_24828);
and U28060 (N_28060,N_24097,N_21930);
nor U28061 (N_28061,N_23750,N_24792);
or U28062 (N_28062,N_24956,N_23017);
or U28063 (N_28063,N_23722,N_23002);
nand U28064 (N_28064,N_24734,N_23192);
and U28065 (N_28065,N_23327,N_24556);
and U28066 (N_28066,N_21145,N_23411);
or U28067 (N_28067,N_20832,N_24354);
nand U28068 (N_28068,N_23521,N_22539);
nor U28069 (N_28069,N_21324,N_24126);
nor U28070 (N_28070,N_22510,N_23698);
and U28071 (N_28071,N_23588,N_20537);
xnor U28072 (N_28072,N_21781,N_20648);
xnor U28073 (N_28073,N_24799,N_21497);
xnor U28074 (N_28074,N_24983,N_20001);
or U28075 (N_28075,N_22026,N_21484);
nor U28076 (N_28076,N_20443,N_23760);
or U28077 (N_28077,N_20838,N_22995);
and U28078 (N_28078,N_22410,N_22058);
xnor U28079 (N_28079,N_24566,N_23451);
nor U28080 (N_28080,N_23740,N_20530);
or U28081 (N_28081,N_22500,N_20467);
nor U28082 (N_28082,N_23604,N_23627);
or U28083 (N_28083,N_22963,N_24903);
nor U28084 (N_28084,N_21591,N_21392);
or U28085 (N_28085,N_23089,N_21549);
or U28086 (N_28086,N_24109,N_21740);
or U28087 (N_28087,N_20666,N_23489);
or U28088 (N_28088,N_20409,N_24120);
nand U28089 (N_28089,N_24983,N_24646);
nand U28090 (N_28090,N_24289,N_24276);
or U28091 (N_28091,N_24618,N_24575);
nor U28092 (N_28092,N_20003,N_20410);
nand U28093 (N_28093,N_22565,N_21073);
or U28094 (N_28094,N_23434,N_21661);
or U28095 (N_28095,N_21514,N_21890);
nand U28096 (N_28096,N_22563,N_24942);
or U28097 (N_28097,N_21514,N_21939);
nand U28098 (N_28098,N_20117,N_24337);
nand U28099 (N_28099,N_22852,N_24924);
nor U28100 (N_28100,N_23913,N_24444);
nor U28101 (N_28101,N_22800,N_23013);
nor U28102 (N_28102,N_23814,N_21917);
and U28103 (N_28103,N_21473,N_20346);
nor U28104 (N_28104,N_23496,N_22560);
nand U28105 (N_28105,N_24860,N_23291);
and U28106 (N_28106,N_22209,N_21668);
xnor U28107 (N_28107,N_23432,N_21188);
nor U28108 (N_28108,N_23905,N_24206);
nand U28109 (N_28109,N_22599,N_22163);
and U28110 (N_28110,N_24010,N_22291);
nor U28111 (N_28111,N_23216,N_22284);
and U28112 (N_28112,N_20926,N_21114);
or U28113 (N_28113,N_21139,N_20056);
nand U28114 (N_28114,N_23205,N_21542);
nand U28115 (N_28115,N_22071,N_23025);
xor U28116 (N_28116,N_24636,N_20850);
or U28117 (N_28117,N_24925,N_22383);
xnor U28118 (N_28118,N_22492,N_20771);
nand U28119 (N_28119,N_21239,N_20435);
xor U28120 (N_28120,N_21145,N_22613);
nand U28121 (N_28121,N_20327,N_23294);
or U28122 (N_28122,N_24249,N_20093);
and U28123 (N_28123,N_24163,N_23436);
nor U28124 (N_28124,N_20569,N_22460);
and U28125 (N_28125,N_23424,N_21855);
nand U28126 (N_28126,N_21396,N_21232);
or U28127 (N_28127,N_22444,N_24510);
and U28128 (N_28128,N_23624,N_21291);
nand U28129 (N_28129,N_24384,N_21617);
xnor U28130 (N_28130,N_23015,N_22151);
nand U28131 (N_28131,N_22642,N_20345);
and U28132 (N_28132,N_22176,N_21014);
and U28133 (N_28133,N_21969,N_24855);
nand U28134 (N_28134,N_21304,N_21523);
nor U28135 (N_28135,N_24177,N_21820);
nor U28136 (N_28136,N_24522,N_22885);
and U28137 (N_28137,N_24015,N_20166);
nor U28138 (N_28138,N_24100,N_21138);
nand U28139 (N_28139,N_21883,N_20241);
nor U28140 (N_28140,N_22175,N_24040);
or U28141 (N_28141,N_24859,N_21509);
nor U28142 (N_28142,N_22043,N_23245);
or U28143 (N_28143,N_23929,N_22425);
xor U28144 (N_28144,N_24220,N_24497);
or U28145 (N_28145,N_20766,N_20732);
xnor U28146 (N_28146,N_23870,N_23567);
nand U28147 (N_28147,N_20627,N_20176);
nor U28148 (N_28148,N_21949,N_20464);
or U28149 (N_28149,N_23869,N_21623);
and U28150 (N_28150,N_20112,N_23941);
or U28151 (N_28151,N_21788,N_23049);
xor U28152 (N_28152,N_20744,N_24756);
xnor U28153 (N_28153,N_20369,N_22050);
nor U28154 (N_28154,N_21568,N_22422);
or U28155 (N_28155,N_23253,N_21320);
and U28156 (N_28156,N_23098,N_24900);
or U28157 (N_28157,N_21197,N_21231);
nand U28158 (N_28158,N_23965,N_24153);
nor U28159 (N_28159,N_23915,N_22547);
nand U28160 (N_28160,N_20993,N_24539);
or U28161 (N_28161,N_22322,N_23860);
or U28162 (N_28162,N_23987,N_20727);
nand U28163 (N_28163,N_23934,N_21024);
xor U28164 (N_28164,N_23200,N_24355);
and U28165 (N_28165,N_20307,N_23207);
or U28166 (N_28166,N_24821,N_20225);
and U28167 (N_28167,N_21587,N_20612);
and U28168 (N_28168,N_24163,N_23292);
nor U28169 (N_28169,N_23732,N_22503);
and U28170 (N_28170,N_23660,N_24326);
nor U28171 (N_28171,N_20021,N_24670);
or U28172 (N_28172,N_21503,N_20412);
and U28173 (N_28173,N_23804,N_22502);
or U28174 (N_28174,N_21525,N_24900);
or U28175 (N_28175,N_23431,N_20307);
nor U28176 (N_28176,N_23313,N_22196);
and U28177 (N_28177,N_20988,N_21952);
or U28178 (N_28178,N_21312,N_24358);
nand U28179 (N_28179,N_24807,N_21676);
nand U28180 (N_28180,N_24928,N_21779);
nand U28181 (N_28181,N_23765,N_24173);
xor U28182 (N_28182,N_23697,N_22023);
nand U28183 (N_28183,N_20863,N_22360);
and U28184 (N_28184,N_20564,N_22214);
and U28185 (N_28185,N_23113,N_23563);
nand U28186 (N_28186,N_20394,N_22684);
or U28187 (N_28187,N_24648,N_23299);
nand U28188 (N_28188,N_21175,N_20493);
or U28189 (N_28189,N_22502,N_20561);
nand U28190 (N_28190,N_24267,N_22278);
or U28191 (N_28191,N_23468,N_24495);
nand U28192 (N_28192,N_24349,N_22481);
or U28193 (N_28193,N_20073,N_23919);
nand U28194 (N_28194,N_22073,N_22401);
nor U28195 (N_28195,N_22486,N_24172);
nor U28196 (N_28196,N_22053,N_24470);
nor U28197 (N_28197,N_21926,N_21584);
xor U28198 (N_28198,N_24687,N_22416);
xnor U28199 (N_28199,N_22896,N_23243);
or U28200 (N_28200,N_22888,N_22255);
xor U28201 (N_28201,N_22944,N_21342);
nor U28202 (N_28202,N_24787,N_22222);
nand U28203 (N_28203,N_23635,N_24012);
or U28204 (N_28204,N_23104,N_20258);
or U28205 (N_28205,N_21419,N_23457);
nor U28206 (N_28206,N_20617,N_20334);
and U28207 (N_28207,N_22182,N_24159);
and U28208 (N_28208,N_20663,N_23948);
nand U28209 (N_28209,N_22964,N_24811);
or U28210 (N_28210,N_20489,N_20927);
nand U28211 (N_28211,N_22511,N_24735);
nor U28212 (N_28212,N_23486,N_20481);
nand U28213 (N_28213,N_24640,N_21421);
nor U28214 (N_28214,N_23924,N_22533);
nor U28215 (N_28215,N_24366,N_22990);
nor U28216 (N_28216,N_24950,N_23202);
nor U28217 (N_28217,N_20351,N_21547);
nor U28218 (N_28218,N_24535,N_22973);
nor U28219 (N_28219,N_22816,N_24625);
and U28220 (N_28220,N_21845,N_20391);
nand U28221 (N_28221,N_20100,N_22814);
nand U28222 (N_28222,N_20922,N_20126);
and U28223 (N_28223,N_21776,N_23185);
nand U28224 (N_28224,N_23076,N_20137);
and U28225 (N_28225,N_22068,N_23065);
or U28226 (N_28226,N_20328,N_22453);
or U28227 (N_28227,N_22997,N_24007);
nand U28228 (N_28228,N_22788,N_21171);
and U28229 (N_28229,N_22355,N_20001);
or U28230 (N_28230,N_22957,N_21688);
nand U28231 (N_28231,N_24332,N_23603);
nor U28232 (N_28232,N_24113,N_23161);
and U28233 (N_28233,N_23480,N_21302);
or U28234 (N_28234,N_21569,N_24999);
and U28235 (N_28235,N_21656,N_23871);
nor U28236 (N_28236,N_23291,N_21072);
nor U28237 (N_28237,N_21602,N_22806);
and U28238 (N_28238,N_24394,N_23864);
nor U28239 (N_28239,N_24269,N_22619);
nor U28240 (N_28240,N_21625,N_22811);
xor U28241 (N_28241,N_23908,N_23354);
nand U28242 (N_28242,N_24928,N_20313);
nand U28243 (N_28243,N_23251,N_22447);
xor U28244 (N_28244,N_24352,N_22155);
and U28245 (N_28245,N_23147,N_24119);
xor U28246 (N_28246,N_24949,N_23961);
and U28247 (N_28247,N_22160,N_24014);
nor U28248 (N_28248,N_22327,N_23923);
nand U28249 (N_28249,N_23280,N_22437);
and U28250 (N_28250,N_22148,N_20182);
and U28251 (N_28251,N_21603,N_21353);
or U28252 (N_28252,N_21747,N_22500);
nand U28253 (N_28253,N_24101,N_23468);
and U28254 (N_28254,N_22359,N_23521);
nand U28255 (N_28255,N_22007,N_21855);
nand U28256 (N_28256,N_20699,N_22513);
nor U28257 (N_28257,N_21218,N_22768);
and U28258 (N_28258,N_23269,N_22608);
nor U28259 (N_28259,N_23915,N_23163);
nand U28260 (N_28260,N_20161,N_24696);
nor U28261 (N_28261,N_20936,N_23325);
nand U28262 (N_28262,N_20603,N_23262);
nor U28263 (N_28263,N_20474,N_23426);
xor U28264 (N_28264,N_21631,N_22906);
nor U28265 (N_28265,N_21278,N_24140);
xor U28266 (N_28266,N_20678,N_24932);
nand U28267 (N_28267,N_21434,N_22138);
nand U28268 (N_28268,N_22650,N_22416);
nor U28269 (N_28269,N_24431,N_22278);
and U28270 (N_28270,N_23221,N_23599);
nor U28271 (N_28271,N_21615,N_24797);
nor U28272 (N_28272,N_23085,N_20688);
or U28273 (N_28273,N_24829,N_22184);
or U28274 (N_28274,N_21625,N_20932);
nand U28275 (N_28275,N_23080,N_23867);
or U28276 (N_28276,N_23978,N_21819);
xnor U28277 (N_28277,N_21770,N_21127);
nand U28278 (N_28278,N_21934,N_21727);
and U28279 (N_28279,N_21904,N_22151);
nor U28280 (N_28280,N_21900,N_20590);
and U28281 (N_28281,N_24638,N_21998);
nor U28282 (N_28282,N_23628,N_23076);
nor U28283 (N_28283,N_24603,N_23880);
nand U28284 (N_28284,N_21972,N_21736);
nor U28285 (N_28285,N_23117,N_23561);
and U28286 (N_28286,N_22901,N_20737);
or U28287 (N_28287,N_20096,N_24955);
or U28288 (N_28288,N_20773,N_23021);
and U28289 (N_28289,N_22361,N_21535);
nand U28290 (N_28290,N_22970,N_24273);
xor U28291 (N_28291,N_24113,N_20902);
and U28292 (N_28292,N_23364,N_23481);
and U28293 (N_28293,N_21958,N_23904);
and U28294 (N_28294,N_21194,N_22726);
or U28295 (N_28295,N_23522,N_24746);
or U28296 (N_28296,N_22219,N_23761);
and U28297 (N_28297,N_21708,N_20748);
and U28298 (N_28298,N_21485,N_22885);
nand U28299 (N_28299,N_24809,N_23281);
nor U28300 (N_28300,N_22150,N_23675);
nor U28301 (N_28301,N_23872,N_23249);
or U28302 (N_28302,N_20257,N_20252);
nor U28303 (N_28303,N_22948,N_20879);
or U28304 (N_28304,N_24590,N_20864);
nand U28305 (N_28305,N_21342,N_21516);
nor U28306 (N_28306,N_23661,N_23326);
or U28307 (N_28307,N_22177,N_20596);
nor U28308 (N_28308,N_23192,N_20921);
and U28309 (N_28309,N_20617,N_20249);
nand U28310 (N_28310,N_24163,N_22540);
nand U28311 (N_28311,N_20538,N_21080);
or U28312 (N_28312,N_20701,N_20303);
and U28313 (N_28313,N_24567,N_21439);
or U28314 (N_28314,N_22851,N_22910);
nand U28315 (N_28315,N_22984,N_20889);
nand U28316 (N_28316,N_24302,N_21452);
nor U28317 (N_28317,N_24160,N_21114);
or U28318 (N_28318,N_22468,N_21932);
or U28319 (N_28319,N_22051,N_21742);
nand U28320 (N_28320,N_20831,N_23906);
xnor U28321 (N_28321,N_23993,N_20693);
nor U28322 (N_28322,N_21561,N_20247);
or U28323 (N_28323,N_21871,N_24633);
or U28324 (N_28324,N_24656,N_22853);
nor U28325 (N_28325,N_24964,N_21439);
or U28326 (N_28326,N_24332,N_20032);
nand U28327 (N_28327,N_21645,N_20934);
and U28328 (N_28328,N_21321,N_20728);
or U28329 (N_28329,N_21807,N_22684);
or U28330 (N_28330,N_20969,N_24137);
or U28331 (N_28331,N_22900,N_23618);
nor U28332 (N_28332,N_21319,N_20894);
nor U28333 (N_28333,N_24332,N_20273);
nand U28334 (N_28334,N_24857,N_21223);
nand U28335 (N_28335,N_20808,N_20621);
nand U28336 (N_28336,N_24203,N_22168);
or U28337 (N_28337,N_21736,N_22351);
nor U28338 (N_28338,N_22622,N_24428);
nand U28339 (N_28339,N_23533,N_20019);
or U28340 (N_28340,N_23344,N_23805);
and U28341 (N_28341,N_20267,N_20228);
nand U28342 (N_28342,N_24356,N_21086);
nand U28343 (N_28343,N_21351,N_24371);
nor U28344 (N_28344,N_21926,N_20775);
or U28345 (N_28345,N_20135,N_21863);
nor U28346 (N_28346,N_21224,N_23764);
xnor U28347 (N_28347,N_23301,N_20499);
and U28348 (N_28348,N_20576,N_22544);
xnor U28349 (N_28349,N_24157,N_24153);
xnor U28350 (N_28350,N_22461,N_23045);
nor U28351 (N_28351,N_24392,N_21499);
nand U28352 (N_28352,N_22585,N_21463);
and U28353 (N_28353,N_20354,N_20489);
and U28354 (N_28354,N_22584,N_24289);
nor U28355 (N_28355,N_24249,N_20841);
or U28356 (N_28356,N_22657,N_22883);
or U28357 (N_28357,N_22439,N_20663);
nor U28358 (N_28358,N_23818,N_20578);
nand U28359 (N_28359,N_22487,N_21989);
and U28360 (N_28360,N_20306,N_22587);
nor U28361 (N_28361,N_20300,N_22198);
and U28362 (N_28362,N_22894,N_24198);
and U28363 (N_28363,N_23271,N_23341);
nor U28364 (N_28364,N_20162,N_22002);
or U28365 (N_28365,N_24693,N_22539);
nand U28366 (N_28366,N_23216,N_24664);
nand U28367 (N_28367,N_21002,N_21159);
nor U28368 (N_28368,N_20570,N_21460);
nand U28369 (N_28369,N_21363,N_24199);
nor U28370 (N_28370,N_20966,N_21536);
nor U28371 (N_28371,N_20089,N_24650);
and U28372 (N_28372,N_21548,N_20115);
and U28373 (N_28373,N_24160,N_20411);
and U28374 (N_28374,N_21814,N_20068);
nor U28375 (N_28375,N_21025,N_23066);
nor U28376 (N_28376,N_24973,N_24515);
or U28377 (N_28377,N_22880,N_21041);
and U28378 (N_28378,N_23650,N_24251);
nor U28379 (N_28379,N_23698,N_22924);
nand U28380 (N_28380,N_20335,N_21796);
and U28381 (N_28381,N_20928,N_24326);
nand U28382 (N_28382,N_23684,N_24193);
nor U28383 (N_28383,N_21485,N_21669);
nor U28384 (N_28384,N_23038,N_23031);
or U28385 (N_28385,N_20303,N_20741);
and U28386 (N_28386,N_24693,N_23276);
and U28387 (N_28387,N_21878,N_21056);
xor U28388 (N_28388,N_20648,N_24521);
nand U28389 (N_28389,N_21001,N_21660);
nand U28390 (N_28390,N_24065,N_20253);
nand U28391 (N_28391,N_23596,N_21922);
and U28392 (N_28392,N_24838,N_22157);
nor U28393 (N_28393,N_20586,N_21243);
nand U28394 (N_28394,N_22733,N_23949);
and U28395 (N_28395,N_23548,N_23613);
or U28396 (N_28396,N_21381,N_24975);
nor U28397 (N_28397,N_24578,N_22125);
nor U28398 (N_28398,N_20166,N_21678);
or U28399 (N_28399,N_21002,N_23323);
or U28400 (N_28400,N_22393,N_24556);
or U28401 (N_28401,N_23134,N_22095);
or U28402 (N_28402,N_21232,N_22429);
and U28403 (N_28403,N_24323,N_23688);
nor U28404 (N_28404,N_21976,N_24438);
nand U28405 (N_28405,N_21369,N_20877);
or U28406 (N_28406,N_20581,N_21077);
or U28407 (N_28407,N_21758,N_22230);
or U28408 (N_28408,N_20556,N_23795);
or U28409 (N_28409,N_22565,N_24887);
or U28410 (N_28410,N_23783,N_24983);
xnor U28411 (N_28411,N_24127,N_21945);
nor U28412 (N_28412,N_20197,N_20955);
or U28413 (N_28413,N_20390,N_23217);
or U28414 (N_28414,N_21774,N_22966);
or U28415 (N_28415,N_22435,N_20852);
nor U28416 (N_28416,N_22710,N_20937);
nor U28417 (N_28417,N_22431,N_21231);
and U28418 (N_28418,N_23044,N_23041);
nand U28419 (N_28419,N_20568,N_23792);
nand U28420 (N_28420,N_23882,N_21582);
nand U28421 (N_28421,N_23011,N_21373);
or U28422 (N_28422,N_20497,N_22107);
xnor U28423 (N_28423,N_24359,N_20238);
xnor U28424 (N_28424,N_20025,N_24057);
nor U28425 (N_28425,N_20703,N_22924);
nor U28426 (N_28426,N_21083,N_24015);
or U28427 (N_28427,N_24437,N_20486);
or U28428 (N_28428,N_23188,N_24975);
or U28429 (N_28429,N_24002,N_21092);
or U28430 (N_28430,N_20828,N_24280);
or U28431 (N_28431,N_23053,N_24355);
nor U28432 (N_28432,N_23189,N_23788);
nand U28433 (N_28433,N_21389,N_24288);
and U28434 (N_28434,N_23190,N_20228);
and U28435 (N_28435,N_24413,N_24225);
and U28436 (N_28436,N_22947,N_21283);
or U28437 (N_28437,N_20782,N_22470);
nand U28438 (N_28438,N_23897,N_22464);
nor U28439 (N_28439,N_23575,N_21425);
or U28440 (N_28440,N_20250,N_22289);
and U28441 (N_28441,N_20192,N_22131);
or U28442 (N_28442,N_23938,N_22185);
xor U28443 (N_28443,N_20520,N_22739);
and U28444 (N_28444,N_23683,N_24269);
and U28445 (N_28445,N_24035,N_20837);
and U28446 (N_28446,N_20325,N_22232);
or U28447 (N_28447,N_24584,N_22892);
nor U28448 (N_28448,N_23015,N_22634);
or U28449 (N_28449,N_20076,N_24624);
nand U28450 (N_28450,N_21844,N_23115);
nor U28451 (N_28451,N_21823,N_20011);
and U28452 (N_28452,N_21765,N_20237);
nor U28453 (N_28453,N_23806,N_24610);
or U28454 (N_28454,N_21176,N_20595);
and U28455 (N_28455,N_24195,N_21071);
nand U28456 (N_28456,N_23685,N_22546);
or U28457 (N_28457,N_20986,N_23199);
nor U28458 (N_28458,N_22874,N_24942);
and U28459 (N_28459,N_20550,N_23475);
and U28460 (N_28460,N_22603,N_21497);
and U28461 (N_28461,N_23410,N_24503);
nand U28462 (N_28462,N_20550,N_20448);
nand U28463 (N_28463,N_23542,N_24874);
or U28464 (N_28464,N_20344,N_23608);
nor U28465 (N_28465,N_24195,N_24112);
and U28466 (N_28466,N_24001,N_20504);
nor U28467 (N_28467,N_21455,N_24571);
or U28468 (N_28468,N_23654,N_24425);
and U28469 (N_28469,N_21393,N_23459);
xnor U28470 (N_28470,N_24720,N_23948);
nand U28471 (N_28471,N_21489,N_22204);
or U28472 (N_28472,N_20769,N_22402);
nand U28473 (N_28473,N_22657,N_22354);
or U28474 (N_28474,N_23737,N_21108);
and U28475 (N_28475,N_23821,N_21582);
nor U28476 (N_28476,N_21777,N_21578);
nor U28477 (N_28477,N_24507,N_21472);
nor U28478 (N_28478,N_22499,N_24040);
nor U28479 (N_28479,N_23569,N_20858);
or U28480 (N_28480,N_24523,N_24948);
or U28481 (N_28481,N_22119,N_22862);
and U28482 (N_28482,N_21863,N_23434);
nand U28483 (N_28483,N_20699,N_23546);
xnor U28484 (N_28484,N_22046,N_24302);
nor U28485 (N_28485,N_23420,N_20714);
xnor U28486 (N_28486,N_23229,N_23025);
and U28487 (N_28487,N_23998,N_24158);
or U28488 (N_28488,N_22577,N_23373);
nor U28489 (N_28489,N_23706,N_24704);
nor U28490 (N_28490,N_24783,N_23053);
and U28491 (N_28491,N_22885,N_24997);
nand U28492 (N_28492,N_23776,N_21913);
nor U28493 (N_28493,N_22397,N_20301);
nor U28494 (N_28494,N_24206,N_21375);
nor U28495 (N_28495,N_20777,N_21448);
and U28496 (N_28496,N_24836,N_24681);
or U28497 (N_28497,N_22047,N_22894);
or U28498 (N_28498,N_23254,N_20797);
or U28499 (N_28499,N_24800,N_20211);
nand U28500 (N_28500,N_22092,N_24737);
or U28501 (N_28501,N_21790,N_22646);
or U28502 (N_28502,N_23693,N_21369);
nand U28503 (N_28503,N_21005,N_24232);
xor U28504 (N_28504,N_24091,N_21677);
nor U28505 (N_28505,N_24212,N_22968);
nand U28506 (N_28506,N_22068,N_24764);
nand U28507 (N_28507,N_21581,N_23668);
nor U28508 (N_28508,N_20254,N_22597);
xor U28509 (N_28509,N_20622,N_22164);
nor U28510 (N_28510,N_21593,N_24842);
or U28511 (N_28511,N_20796,N_24912);
nor U28512 (N_28512,N_20083,N_20843);
nor U28513 (N_28513,N_22364,N_20735);
nor U28514 (N_28514,N_20258,N_24480);
nor U28515 (N_28515,N_24797,N_24529);
and U28516 (N_28516,N_24490,N_23166);
or U28517 (N_28517,N_20298,N_21941);
nand U28518 (N_28518,N_20021,N_20701);
nor U28519 (N_28519,N_24427,N_23856);
or U28520 (N_28520,N_21204,N_22124);
nor U28521 (N_28521,N_23870,N_20082);
xor U28522 (N_28522,N_22329,N_24283);
nor U28523 (N_28523,N_20963,N_20218);
or U28524 (N_28524,N_23499,N_24965);
and U28525 (N_28525,N_23682,N_24051);
or U28526 (N_28526,N_24768,N_22538);
and U28527 (N_28527,N_23354,N_23691);
nor U28528 (N_28528,N_21273,N_20177);
nor U28529 (N_28529,N_24668,N_20386);
and U28530 (N_28530,N_23579,N_22246);
or U28531 (N_28531,N_24794,N_22606);
or U28532 (N_28532,N_20955,N_23178);
or U28533 (N_28533,N_24008,N_21092);
nor U28534 (N_28534,N_20647,N_20292);
or U28535 (N_28535,N_23004,N_22999);
nor U28536 (N_28536,N_23828,N_20717);
nand U28537 (N_28537,N_20957,N_21284);
or U28538 (N_28538,N_23097,N_20046);
nor U28539 (N_28539,N_22951,N_21444);
nand U28540 (N_28540,N_24115,N_22881);
nor U28541 (N_28541,N_22538,N_21300);
and U28542 (N_28542,N_24978,N_22375);
nand U28543 (N_28543,N_22303,N_23733);
nor U28544 (N_28544,N_22500,N_21594);
xnor U28545 (N_28545,N_24479,N_23693);
or U28546 (N_28546,N_21074,N_23249);
nand U28547 (N_28547,N_20591,N_20597);
and U28548 (N_28548,N_24029,N_20070);
nor U28549 (N_28549,N_21595,N_23677);
nand U28550 (N_28550,N_23236,N_24099);
and U28551 (N_28551,N_22369,N_20684);
or U28552 (N_28552,N_21878,N_23813);
nor U28553 (N_28553,N_21479,N_22798);
and U28554 (N_28554,N_20348,N_24443);
and U28555 (N_28555,N_20658,N_23056);
and U28556 (N_28556,N_23361,N_20756);
or U28557 (N_28557,N_23236,N_20174);
nor U28558 (N_28558,N_21938,N_22730);
and U28559 (N_28559,N_22203,N_23086);
and U28560 (N_28560,N_22229,N_22381);
nand U28561 (N_28561,N_22610,N_20279);
and U28562 (N_28562,N_20928,N_22596);
nand U28563 (N_28563,N_23480,N_24492);
and U28564 (N_28564,N_20846,N_22994);
nor U28565 (N_28565,N_22000,N_20221);
and U28566 (N_28566,N_23509,N_24600);
or U28567 (N_28567,N_21455,N_20429);
or U28568 (N_28568,N_23393,N_20833);
nand U28569 (N_28569,N_21623,N_24895);
nand U28570 (N_28570,N_24463,N_20757);
nor U28571 (N_28571,N_24289,N_24999);
nand U28572 (N_28572,N_22576,N_24971);
nand U28573 (N_28573,N_23930,N_20995);
nand U28574 (N_28574,N_24206,N_23442);
nand U28575 (N_28575,N_21025,N_24557);
and U28576 (N_28576,N_23638,N_23028);
nand U28577 (N_28577,N_20109,N_23756);
nor U28578 (N_28578,N_22713,N_21386);
nand U28579 (N_28579,N_23224,N_23661);
or U28580 (N_28580,N_22632,N_21720);
and U28581 (N_28581,N_24700,N_21861);
or U28582 (N_28582,N_24626,N_23697);
nand U28583 (N_28583,N_20552,N_24446);
and U28584 (N_28584,N_22140,N_23138);
or U28585 (N_28585,N_23255,N_23130);
or U28586 (N_28586,N_20221,N_22969);
nor U28587 (N_28587,N_20296,N_23424);
or U28588 (N_28588,N_23664,N_21205);
nand U28589 (N_28589,N_23141,N_21081);
nand U28590 (N_28590,N_22637,N_20276);
xor U28591 (N_28591,N_20502,N_22313);
xor U28592 (N_28592,N_22768,N_24310);
nor U28593 (N_28593,N_20953,N_21046);
or U28594 (N_28594,N_23502,N_21359);
nor U28595 (N_28595,N_22580,N_23279);
and U28596 (N_28596,N_22844,N_23334);
nor U28597 (N_28597,N_20415,N_24537);
or U28598 (N_28598,N_20401,N_20989);
and U28599 (N_28599,N_24324,N_22012);
nand U28600 (N_28600,N_23074,N_23817);
and U28601 (N_28601,N_24938,N_23905);
and U28602 (N_28602,N_24503,N_20208);
and U28603 (N_28603,N_20037,N_24634);
and U28604 (N_28604,N_22986,N_22300);
nor U28605 (N_28605,N_21183,N_20551);
or U28606 (N_28606,N_21877,N_24603);
xnor U28607 (N_28607,N_24087,N_24385);
and U28608 (N_28608,N_22641,N_24101);
or U28609 (N_28609,N_20868,N_23365);
xor U28610 (N_28610,N_20960,N_20579);
or U28611 (N_28611,N_21310,N_22171);
nor U28612 (N_28612,N_20650,N_23991);
nand U28613 (N_28613,N_24708,N_21228);
nor U28614 (N_28614,N_24797,N_21097);
nand U28615 (N_28615,N_21755,N_21273);
nor U28616 (N_28616,N_24296,N_22872);
nand U28617 (N_28617,N_24721,N_22452);
xnor U28618 (N_28618,N_20177,N_24539);
or U28619 (N_28619,N_24094,N_21547);
and U28620 (N_28620,N_21945,N_23696);
and U28621 (N_28621,N_22088,N_21088);
nor U28622 (N_28622,N_23340,N_21918);
and U28623 (N_28623,N_24108,N_23762);
or U28624 (N_28624,N_22905,N_22856);
nand U28625 (N_28625,N_20370,N_24039);
or U28626 (N_28626,N_20749,N_20944);
xnor U28627 (N_28627,N_23982,N_20502);
and U28628 (N_28628,N_21362,N_20471);
nor U28629 (N_28629,N_22111,N_23982);
nand U28630 (N_28630,N_21390,N_21702);
or U28631 (N_28631,N_21439,N_21440);
or U28632 (N_28632,N_22217,N_23411);
nor U28633 (N_28633,N_22347,N_22411);
or U28634 (N_28634,N_23078,N_22546);
and U28635 (N_28635,N_23470,N_20933);
and U28636 (N_28636,N_20038,N_20223);
and U28637 (N_28637,N_22188,N_24530);
and U28638 (N_28638,N_22596,N_23441);
nand U28639 (N_28639,N_20016,N_21873);
or U28640 (N_28640,N_24603,N_22694);
or U28641 (N_28641,N_20893,N_21818);
nand U28642 (N_28642,N_20167,N_24656);
nor U28643 (N_28643,N_21614,N_20560);
nor U28644 (N_28644,N_21694,N_20153);
nand U28645 (N_28645,N_24851,N_21492);
nor U28646 (N_28646,N_23176,N_20375);
nor U28647 (N_28647,N_24411,N_23428);
and U28648 (N_28648,N_20803,N_20964);
or U28649 (N_28649,N_20843,N_22046);
xor U28650 (N_28650,N_23930,N_21922);
nand U28651 (N_28651,N_22517,N_23040);
xor U28652 (N_28652,N_24598,N_21393);
and U28653 (N_28653,N_21046,N_22407);
and U28654 (N_28654,N_23289,N_22971);
or U28655 (N_28655,N_21642,N_23679);
nor U28656 (N_28656,N_24261,N_21922);
xor U28657 (N_28657,N_21441,N_20089);
nand U28658 (N_28658,N_20200,N_20039);
nor U28659 (N_28659,N_20948,N_21171);
or U28660 (N_28660,N_21369,N_24484);
or U28661 (N_28661,N_21905,N_23782);
nor U28662 (N_28662,N_21650,N_21148);
nor U28663 (N_28663,N_23113,N_22144);
and U28664 (N_28664,N_22593,N_22095);
or U28665 (N_28665,N_22174,N_24874);
nor U28666 (N_28666,N_22648,N_20115);
and U28667 (N_28667,N_23358,N_20655);
xnor U28668 (N_28668,N_21147,N_22350);
or U28669 (N_28669,N_22237,N_21321);
or U28670 (N_28670,N_22140,N_23752);
or U28671 (N_28671,N_20482,N_24003);
or U28672 (N_28672,N_20171,N_20813);
nand U28673 (N_28673,N_22796,N_20551);
or U28674 (N_28674,N_20346,N_23190);
and U28675 (N_28675,N_20327,N_20644);
nor U28676 (N_28676,N_20726,N_24845);
and U28677 (N_28677,N_23717,N_23425);
and U28678 (N_28678,N_24602,N_24727);
or U28679 (N_28679,N_20610,N_21554);
nand U28680 (N_28680,N_22915,N_23537);
and U28681 (N_28681,N_22298,N_22906);
nor U28682 (N_28682,N_24417,N_24835);
xor U28683 (N_28683,N_24498,N_21420);
and U28684 (N_28684,N_22872,N_21179);
or U28685 (N_28685,N_22111,N_22481);
and U28686 (N_28686,N_20030,N_20045);
nand U28687 (N_28687,N_21690,N_24043);
nor U28688 (N_28688,N_20213,N_22172);
nand U28689 (N_28689,N_20426,N_23717);
nand U28690 (N_28690,N_23613,N_23730);
and U28691 (N_28691,N_21802,N_24002);
nor U28692 (N_28692,N_20432,N_24616);
and U28693 (N_28693,N_23486,N_23178);
or U28694 (N_28694,N_23332,N_20029);
and U28695 (N_28695,N_20643,N_22753);
nand U28696 (N_28696,N_24048,N_21681);
or U28697 (N_28697,N_20491,N_23559);
nor U28698 (N_28698,N_20419,N_23205);
or U28699 (N_28699,N_22099,N_24191);
nand U28700 (N_28700,N_23855,N_23345);
nor U28701 (N_28701,N_21614,N_22385);
xnor U28702 (N_28702,N_20677,N_24434);
and U28703 (N_28703,N_20694,N_20631);
or U28704 (N_28704,N_22546,N_23920);
and U28705 (N_28705,N_20197,N_22889);
nand U28706 (N_28706,N_21458,N_21013);
and U28707 (N_28707,N_20116,N_20022);
nor U28708 (N_28708,N_20616,N_24982);
or U28709 (N_28709,N_21180,N_20819);
xor U28710 (N_28710,N_23359,N_20416);
nor U28711 (N_28711,N_22612,N_20612);
nand U28712 (N_28712,N_24634,N_20600);
nor U28713 (N_28713,N_24525,N_20841);
nor U28714 (N_28714,N_21510,N_23337);
nor U28715 (N_28715,N_21052,N_22575);
xor U28716 (N_28716,N_24630,N_21222);
or U28717 (N_28717,N_20119,N_20970);
or U28718 (N_28718,N_24408,N_23055);
nand U28719 (N_28719,N_21750,N_24964);
nand U28720 (N_28720,N_23683,N_23477);
or U28721 (N_28721,N_21856,N_24102);
nand U28722 (N_28722,N_23662,N_20015);
nand U28723 (N_28723,N_23231,N_22187);
or U28724 (N_28724,N_21134,N_23294);
and U28725 (N_28725,N_21599,N_22322);
and U28726 (N_28726,N_22852,N_20358);
xor U28727 (N_28727,N_21880,N_20435);
or U28728 (N_28728,N_22847,N_20875);
nand U28729 (N_28729,N_24473,N_23978);
or U28730 (N_28730,N_22502,N_20558);
or U28731 (N_28731,N_21474,N_23021);
and U28732 (N_28732,N_22456,N_22208);
or U28733 (N_28733,N_20579,N_24346);
and U28734 (N_28734,N_20248,N_22262);
nand U28735 (N_28735,N_21064,N_24831);
xnor U28736 (N_28736,N_21332,N_20466);
nand U28737 (N_28737,N_22276,N_20462);
nand U28738 (N_28738,N_24589,N_20285);
nor U28739 (N_28739,N_21360,N_22870);
xor U28740 (N_28740,N_20673,N_20220);
nor U28741 (N_28741,N_20703,N_21487);
nand U28742 (N_28742,N_23829,N_20540);
nor U28743 (N_28743,N_24366,N_20625);
and U28744 (N_28744,N_22159,N_20831);
and U28745 (N_28745,N_24494,N_21271);
and U28746 (N_28746,N_22707,N_20111);
and U28747 (N_28747,N_20570,N_21952);
xor U28748 (N_28748,N_22287,N_20283);
nor U28749 (N_28749,N_21730,N_20837);
xnor U28750 (N_28750,N_20479,N_24278);
xnor U28751 (N_28751,N_20968,N_23372);
xnor U28752 (N_28752,N_21375,N_21055);
and U28753 (N_28753,N_24878,N_20457);
or U28754 (N_28754,N_23166,N_22659);
nor U28755 (N_28755,N_21200,N_21209);
and U28756 (N_28756,N_24408,N_24222);
xor U28757 (N_28757,N_24440,N_22269);
nand U28758 (N_28758,N_21107,N_21744);
nor U28759 (N_28759,N_20188,N_23893);
xor U28760 (N_28760,N_24539,N_22667);
nand U28761 (N_28761,N_20867,N_22068);
nand U28762 (N_28762,N_23915,N_20406);
nor U28763 (N_28763,N_21511,N_21132);
nand U28764 (N_28764,N_23878,N_22746);
nand U28765 (N_28765,N_22022,N_23099);
xor U28766 (N_28766,N_23740,N_23190);
or U28767 (N_28767,N_24572,N_20926);
and U28768 (N_28768,N_22119,N_22207);
or U28769 (N_28769,N_23694,N_22555);
nand U28770 (N_28770,N_24037,N_22390);
nor U28771 (N_28771,N_24131,N_24293);
xor U28772 (N_28772,N_21112,N_20916);
and U28773 (N_28773,N_23206,N_20648);
and U28774 (N_28774,N_24866,N_20970);
nor U28775 (N_28775,N_23980,N_23408);
or U28776 (N_28776,N_22872,N_22149);
nor U28777 (N_28777,N_22131,N_24473);
or U28778 (N_28778,N_20661,N_24360);
xor U28779 (N_28779,N_23997,N_21390);
xnor U28780 (N_28780,N_23456,N_21865);
nor U28781 (N_28781,N_21263,N_24037);
nand U28782 (N_28782,N_20189,N_22773);
and U28783 (N_28783,N_21802,N_24682);
nor U28784 (N_28784,N_22168,N_24448);
nand U28785 (N_28785,N_20082,N_20993);
or U28786 (N_28786,N_24192,N_24417);
and U28787 (N_28787,N_24800,N_22628);
xnor U28788 (N_28788,N_24531,N_20583);
and U28789 (N_28789,N_21230,N_23432);
and U28790 (N_28790,N_23409,N_20535);
and U28791 (N_28791,N_22404,N_24170);
nor U28792 (N_28792,N_22558,N_24653);
and U28793 (N_28793,N_22694,N_20498);
nand U28794 (N_28794,N_22549,N_20888);
nor U28795 (N_28795,N_22754,N_20524);
nor U28796 (N_28796,N_22125,N_23715);
and U28797 (N_28797,N_21501,N_21861);
and U28798 (N_28798,N_21892,N_24020);
and U28799 (N_28799,N_22576,N_20898);
or U28800 (N_28800,N_22971,N_23298);
or U28801 (N_28801,N_22322,N_20827);
and U28802 (N_28802,N_22649,N_22408);
nand U28803 (N_28803,N_22596,N_22007);
nand U28804 (N_28804,N_20878,N_20301);
and U28805 (N_28805,N_24825,N_23238);
nand U28806 (N_28806,N_23290,N_21984);
nor U28807 (N_28807,N_24580,N_20316);
and U28808 (N_28808,N_24122,N_24424);
or U28809 (N_28809,N_20256,N_23299);
nor U28810 (N_28810,N_23422,N_23845);
and U28811 (N_28811,N_20968,N_21963);
xor U28812 (N_28812,N_20447,N_23241);
nor U28813 (N_28813,N_22265,N_21219);
xor U28814 (N_28814,N_23883,N_24071);
nor U28815 (N_28815,N_22365,N_24112);
xor U28816 (N_28816,N_23782,N_24203);
and U28817 (N_28817,N_23802,N_24309);
xor U28818 (N_28818,N_20254,N_23382);
or U28819 (N_28819,N_20623,N_22417);
xnor U28820 (N_28820,N_23811,N_22882);
nor U28821 (N_28821,N_20728,N_21012);
xnor U28822 (N_28822,N_22466,N_22859);
or U28823 (N_28823,N_22688,N_24087);
or U28824 (N_28824,N_21045,N_22006);
and U28825 (N_28825,N_20443,N_21509);
or U28826 (N_28826,N_22922,N_24959);
and U28827 (N_28827,N_22419,N_23411);
and U28828 (N_28828,N_22551,N_24567);
nand U28829 (N_28829,N_20912,N_24320);
and U28830 (N_28830,N_22441,N_20595);
nand U28831 (N_28831,N_21487,N_20383);
or U28832 (N_28832,N_20486,N_21268);
nand U28833 (N_28833,N_20893,N_21278);
nor U28834 (N_28834,N_22181,N_23189);
xor U28835 (N_28835,N_23486,N_24652);
nor U28836 (N_28836,N_23442,N_23272);
xnor U28837 (N_28837,N_20345,N_23386);
and U28838 (N_28838,N_21214,N_24878);
and U28839 (N_28839,N_24444,N_21176);
and U28840 (N_28840,N_21514,N_23057);
nor U28841 (N_28841,N_20369,N_20072);
nor U28842 (N_28842,N_20396,N_24398);
nor U28843 (N_28843,N_22296,N_23620);
nor U28844 (N_28844,N_20102,N_23749);
or U28845 (N_28845,N_22848,N_23654);
nand U28846 (N_28846,N_20244,N_20699);
nand U28847 (N_28847,N_23672,N_20847);
nor U28848 (N_28848,N_24710,N_21554);
and U28849 (N_28849,N_21799,N_20495);
xor U28850 (N_28850,N_21343,N_22428);
xor U28851 (N_28851,N_20921,N_24172);
nand U28852 (N_28852,N_22681,N_21217);
and U28853 (N_28853,N_20616,N_22861);
nand U28854 (N_28854,N_23919,N_24674);
nand U28855 (N_28855,N_22110,N_21218);
and U28856 (N_28856,N_23278,N_22460);
nor U28857 (N_28857,N_23606,N_22033);
xor U28858 (N_28858,N_22526,N_22271);
and U28859 (N_28859,N_21390,N_24718);
and U28860 (N_28860,N_23435,N_23719);
nand U28861 (N_28861,N_22878,N_24580);
and U28862 (N_28862,N_20814,N_23774);
or U28863 (N_28863,N_21363,N_20824);
and U28864 (N_28864,N_20421,N_21767);
and U28865 (N_28865,N_23827,N_22595);
nor U28866 (N_28866,N_20400,N_22176);
and U28867 (N_28867,N_24896,N_21193);
or U28868 (N_28868,N_21178,N_22483);
or U28869 (N_28869,N_23939,N_22017);
or U28870 (N_28870,N_21121,N_20893);
or U28871 (N_28871,N_21932,N_23914);
and U28872 (N_28872,N_24006,N_24289);
xor U28873 (N_28873,N_24432,N_22686);
nand U28874 (N_28874,N_22156,N_24786);
or U28875 (N_28875,N_21867,N_22458);
or U28876 (N_28876,N_21652,N_23489);
xor U28877 (N_28877,N_21747,N_23254);
or U28878 (N_28878,N_23551,N_21820);
or U28879 (N_28879,N_22650,N_23295);
or U28880 (N_28880,N_21655,N_24825);
or U28881 (N_28881,N_22410,N_21928);
and U28882 (N_28882,N_21145,N_21906);
or U28883 (N_28883,N_21958,N_23880);
or U28884 (N_28884,N_22639,N_20833);
or U28885 (N_28885,N_23422,N_20277);
nand U28886 (N_28886,N_23857,N_20381);
and U28887 (N_28887,N_20679,N_21365);
nand U28888 (N_28888,N_20778,N_24701);
and U28889 (N_28889,N_24493,N_21454);
and U28890 (N_28890,N_22221,N_21262);
nand U28891 (N_28891,N_20468,N_23323);
and U28892 (N_28892,N_20689,N_22770);
or U28893 (N_28893,N_21100,N_20609);
nand U28894 (N_28894,N_22833,N_22784);
and U28895 (N_28895,N_22727,N_22160);
or U28896 (N_28896,N_21543,N_22807);
and U28897 (N_28897,N_24192,N_24243);
nand U28898 (N_28898,N_24810,N_23978);
xnor U28899 (N_28899,N_20267,N_24393);
or U28900 (N_28900,N_21546,N_23498);
nand U28901 (N_28901,N_22064,N_23413);
nand U28902 (N_28902,N_23076,N_23776);
nand U28903 (N_28903,N_21475,N_20996);
and U28904 (N_28904,N_23832,N_20709);
nand U28905 (N_28905,N_21785,N_24588);
or U28906 (N_28906,N_24515,N_21862);
or U28907 (N_28907,N_23892,N_21771);
nor U28908 (N_28908,N_20591,N_24978);
nand U28909 (N_28909,N_23216,N_24358);
and U28910 (N_28910,N_24142,N_20610);
nor U28911 (N_28911,N_20216,N_23028);
nand U28912 (N_28912,N_22480,N_22514);
and U28913 (N_28913,N_20005,N_21027);
or U28914 (N_28914,N_24744,N_22588);
nor U28915 (N_28915,N_21541,N_20386);
nand U28916 (N_28916,N_21001,N_22227);
xor U28917 (N_28917,N_20010,N_22092);
xnor U28918 (N_28918,N_20382,N_21979);
or U28919 (N_28919,N_21125,N_21023);
nor U28920 (N_28920,N_24482,N_20767);
nor U28921 (N_28921,N_24443,N_20866);
nand U28922 (N_28922,N_24807,N_24061);
nand U28923 (N_28923,N_24132,N_23073);
nor U28924 (N_28924,N_20930,N_21929);
nor U28925 (N_28925,N_22286,N_21589);
nand U28926 (N_28926,N_22278,N_24625);
and U28927 (N_28927,N_24111,N_22604);
nor U28928 (N_28928,N_20865,N_22905);
and U28929 (N_28929,N_22609,N_22162);
or U28930 (N_28930,N_21965,N_23957);
nor U28931 (N_28931,N_20507,N_22804);
or U28932 (N_28932,N_20511,N_21614);
or U28933 (N_28933,N_21190,N_22559);
nand U28934 (N_28934,N_24812,N_21571);
xor U28935 (N_28935,N_23017,N_24323);
nand U28936 (N_28936,N_22564,N_22923);
and U28937 (N_28937,N_22687,N_22496);
and U28938 (N_28938,N_21604,N_20638);
nor U28939 (N_28939,N_24975,N_23012);
or U28940 (N_28940,N_23896,N_24070);
or U28941 (N_28941,N_24418,N_22612);
xnor U28942 (N_28942,N_23395,N_21605);
xnor U28943 (N_28943,N_20311,N_21065);
nand U28944 (N_28944,N_22883,N_23194);
or U28945 (N_28945,N_24231,N_24401);
nor U28946 (N_28946,N_21970,N_24237);
and U28947 (N_28947,N_21110,N_24424);
nand U28948 (N_28948,N_22012,N_20999);
nor U28949 (N_28949,N_22006,N_22371);
nand U28950 (N_28950,N_23921,N_20083);
or U28951 (N_28951,N_20658,N_22190);
and U28952 (N_28952,N_20872,N_20824);
nor U28953 (N_28953,N_24006,N_21683);
nand U28954 (N_28954,N_23339,N_20032);
nand U28955 (N_28955,N_24530,N_24672);
or U28956 (N_28956,N_24661,N_21233);
nand U28957 (N_28957,N_22202,N_22426);
and U28958 (N_28958,N_20805,N_23959);
nor U28959 (N_28959,N_23003,N_23236);
or U28960 (N_28960,N_21280,N_23445);
xnor U28961 (N_28961,N_23822,N_23685);
nand U28962 (N_28962,N_20754,N_24607);
nor U28963 (N_28963,N_21877,N_20249);
or U28964 (N_28964,N_21028,N_21770);
xnor U28965 (N_28965,N_23658,N_23420);
and U28966 (N_28966,N_23600,N_21327);
nand U28967 (N_28967,N_22139,N_20248);
and U28968 (N_28968,N_21829,N_21311);
or U28969 (N_28969,N_24449,N_23318);
and U28970 (N_28970,N_21760,N_21769);
nand U28971 (N_28971,N_21410,N_23565);
nand U28972 (N_28972,N_21654,N_21265);
or U28973 (N_28973,N_21793,N_20702);
nor U28974 (N_28974,N_24772,N_21643);
xor U28975 (N_28975,N_23508,N_23328);
and U28976 (N_28976,N_23767,N_20859);
nand U28977 (N_28977,N_20939,N_20599);
nor U28978 (N_28978,N_20389,N_24664);
and U28979 (N_28979,N_24038,N_23849);
nand U28980 (N_28980,N_20102,N_23388);
or U28981 (N_28981,N_20844,N_24055);
nor U28982 (N_28982,N_23593,N_24432);
nand U28983 (N_28983,N_21963,N_22972);
nor U28984 (N_28984,N_22095,N_21470);
nor U28985 (N_28985,N_20316,N_23868);
nand U28986 (N_28986,N_21041,N_22575);
nand U28987 (N_28987,N_24716,N_22716);
nand U28988 (N_28988,N_23500,N_24290);
or U28989 (N_28989,N_20638,N_24775);
nand U28990 (N_28990,N_22400,N_23961);
nand U28991 (N_28991,N_24751,N_23359);
nor U28992 (N_28992,N_21150,N_21515);
nor U28993 (N_28993,N_20677,N_20722);
and U28994 (N_28994,N_24282,N_23458);
nand U28995 (N_28995,N_23119,N_24326);
xnor U28996 (N_28996,N_20728,N_20842);
or U28997 (N_28997,N_21247,N_21839);
nor U28998 (N_28998,N_22188,N_22672);
xnor U28999 (N_28999,N_21862,N_21124);
nor U29000 (N_29000,N_22068,N_23957);
and U29001 (N_29001,N_24806,N_22600);
and U29002 (N_29002,N_20848,N_23893);
nor U29003 (N_29003,N_22970,N_23851);
and U29004 (N_29004,N_23160,N_20344);
nor U29005 (N_29005,N_24527,N_23652);
nand U29006 (N_29006,N_21671,N_21499);
nand U29007 (N_29007,N_24921,N_22420);
nand U29008 (N_29008,N_24726,N_20745);
and U29009 (N_29009,N_22694,N_20503);
and U29010 (N_29010,N_21805,N_22717);
nand U29011 (N_29011,N_20291,N_24655);
or U29012 (N_29012,N_21074,N_20547);
nor U29013 (N_29013,N_24975,N_23336);
and U29014 (N_29014,N_23021,N_24294);
or U29015 (N_29015,N_21483,N_24696);
and U29016 (N_29016,N_22130,N_20123);
nor U29017 (N_29017,N_20974,N_21818);
and U29018 (N_29018,N_20494,N_24947);
and U29019 (N_29019,N_23583,N_21700);
or U29020 (N_29020,N_22240,N_23522);
or U29021 (N_29021,N_20353,N_24318);
or U29022 (N_29022,N_20362,N_23027);
or U29023 (N_29023,N_24907,N_21277);
and U29024 (N_29024,N_24285,N_20744);
and U29025 (N_29025,N_21296,N_24461);
nand U29026 (N_29026,N_24948,N_21862);
nand U29027 (N_29027,N_21967,N_20288);
or U29028 (N_29028,N_22458,N_21642);
nand U29029 (N_29029,N_21177,N_23028);
nand U29030 (N_29030,N_20236,N_21358);
and U29031 (N_29031,N_20168,N_20052);
or U29032 (N_29032,N_20727,N_23350);
or U29033 (N_29033,N_22664,N_21183);
nand U29034 (N_29034,N_24605,N_22982);
xnor U29035 (N_29035,N_21722,N_23233);
or U29036 (N_29036,N_22521,N_24737);
xnor U29037 (N_29037,N_21899,N_20981);
or U29038 (N_29038,N_24039,N_24105);
nand U29039 (N_29039,N_24716,N_20151);
nand U29040 (N_29040,N_22106,N_21614);
or U29041 (N_29041,N_20365,N_22175);
and U29042 (N_29042,N_21337,N_24477);
or U29043 (N_29043,N_22637,N_22361);
nand U29044 (N_29044,N_23121,N_21770);
and U29045 (N_29045,N_21297,N_24949);
nor U29046 (N_29046,N_21512,N_20252);
and U29047 (N_29047,N_22636,N_22519);
nor U29048 (N_29048,N_22158,N_20014);
nor U29049 (N_29049,N_20726,N_22402);
and U29050 (N_29050,N_23997,N_21296);
or U29051 (N_29051,N_23161,N_22545);
nor U29052 (N_29052,N_24303,N_22447);
nand U29053 (N_29053,N_24160,N_24114);
and U29054 (N_29054,N_21248,N_20990);
or U29055 (N_29055,N_20790,N_20886);
and U29056 (N_29056,N_21516,N_21197);
nor U29057 (N_29057,N_22542,N_22949);
and U29058 (N_29058,N_21766,N_20025);
nor U29059 (N_29059,N_21778,N_24059);
and U29060 (N_29060,N_23029,N_21395);
nor U29061 (N_29061,N_24941,N_23886);
or U29062 (N_29062,N_22269,N_21700);
nand U29063 (N_29063,N_23586,N_20382);
and U29064 (N_29064,N_23672,N_23548);
and U29065 (N_29065,N_23297,N_24365);
and U29066 (N_29066,N_21926,N_24654);
nand U29067 (N_29067,N_24156,N_21853);
or U29068 (N_29068,N_23082,N_20051);
and U29069 (N_29069,N_20358,N_20563);
xnor U29070 (N_29070,N_21007,N_22712);
xnor U29071 (N_29071,N_20051,N_20493);
nor U29072 (N_29072,N_23669,N_24914);
nand U29073 (N_29073,N_20353,N_20298);
nand U29074 (N_29074,N_24997,N_23077);
nand U29075 (N_29075,N_21390,N_22543);
nand U29076 (N_29076,N_21826,N_20442);
and U29077 (N_29077,N_20768,N_23900);
or U29078 (N_29078,N_20817,N_20007);
nor U29079 (N_29079,N_20858,N_20372);
and U29080 (N_29080,N_21208,N_20506);
nor U29081 (N_29081,N_22074,N_24034);
nand U29082 (N_29082,N_20916,N_22378);
and U29083 (N_29083,N_21719,N_23800);
nand U29084 (N_29084,N_20901,N_23655);
nor U29085 (N_29085,N_22033,N_22509);
nand U29086 (N_29086,N_22635,N_20685);
and U29087 (N_29087,N_21488,N_23790);
xnor U29088 (N_29088,N_20077,N_20920);
or U29089 (N_29089,N_22723,N_21487);
and U29090 (N_29090,N_20426,N_24479);
nand U29091 (N_29091,N_20748,N_21474);
and U29092 (N_29092,N_21079,N_23779);
nor U29093 (N_29093,N_23728,N_24953);
or U29094 (N_29094,N_20060,N_21207);
nand U29095 (N_29095,N_23597,N_23290);
and U29096 (N_29096,N_22552,N_22952);
nor U29097 (N_29097,N_22440,N_20014);
nor U29098 (N_29098,N_20607,N_20922);
xnor U29099 (N_29099,N_23893,N_20033);
nand U29100 (N_29100,N_21608,N_21941);
and U29101 (N_29101,N_22730,N_21604);
or U29102 (N_29102,N_23539,N_23759);
nor U29103 (N_29103,N_22258,N_22318);
nand U29104 (N_29104,N_20751,N_24739);
nand U29105 (N_29105,N_22582,N_20939);
or U29106 (N_29106,N_21017,N_20602);
or U29107 (N_29107,N_23431,N_20301);
nor U29108 (N_29108,N_22358,N_24726);
or U29109 (N_29109,N_24089,N_21496);
nand U29110 (N_29110,N_21044,N_24920);
or U29111 (N_29111,N_24929,N_21689);
and U29112 (N_29112,N_22363,N_21451);
and U29113 (N_29113,N_23005,N_21370);
nand U29114 (N_29114,N_20983,N_24445);
and U29115 (N_29115,N_24998,N_22755);
nand U29116 (N_29116,N_24489,N_21485);
and U29117 (N_29117,N_21563,N_23469);
or U29118 (N_29118,N_23012,N_24735);
nand U29119 (N_29119,N_23626,N_24492);
or U29120 (N_29120,N_23058,N_21336);
or U29121 (N_29121,N_23437,N_22998);
or U29122 (N_29122,N_24174,N_24789);
and U29123 (N_29123,N_22394,N_20296);
and U29124 (N_29124,N_22336,N_22235);
or U29125 (N_29125,N_24799,N_22177);
nand U29126 (N_29126,N_22488,N_21184);
xor U29127 (N_29127,N_21340,N_24428);
nand U29128 (N_29128,N_24179,N_22217);
nand U29129 (N_29129,N_21101,N_21624);
or U29130 (N_29130,N_20846,N_21309);
and U29131 (N_29131,N_24795,N_20494);
and U29132 (N_29132,N_23477,N_20524);
or U29133 (N_29133,N_23444,N_24173);
or U29134 (N_29134,N_22078,N_23083);
and U29135 (N_29135,N_22315,N_24664);
or U29136 (N_29136,N_23193,N_21713);
and U29137 (N_29137,N_22646,N_23168);
nor U29138 (N_29138,N_22113,N_23542);
nor U29139 (N_29139,N_24176,N_21425);
or U29140 (N_29140,N_20384,N_22140);
xor U29141 (N_29141,N_23918,N_20229);
and U29142 (N_29142,N_23411,N_20572);
and U29143 (N_29143,N_24892,N_21010);
nor U29144 (N_29144,N_20536,N_21851);
nand U29145 (N_29145,N_21038,N_24995);
and U29146 (N_29146,N_24373,N_20483);
nor U29147 (N_29147,N_20739,N_22683);
nand U29148 (N_29148,N_23449,N_20871);
and U29149 (N_29149,N_21325,N_21026);
nor U29150 (N_29150,N_24842,N_20490);
and U29151 (N_29151,N_20249,N_20917);
nor U29152 (N_29152,N_24025,N_21937);
and U29153 (N_29153,N_20972,N_23755);
nand U29154 (N_29154,N_22567,N_20645);
nor U29155 (N_29155,N_20285,N_23049);
nand U29156 (N_29156,N_21486,N_23944);
nand U29157 (N_29157,N_22270,N_23464);
and U29158 (N_29158,N_20083,N_20862);
and U29159 (N_29159,N_23489,N_23142);
nor U29160 (N_29160,N_20734,N_21685);
xor U29161 (N_29161,N_21706,N_24319);
nor U29162 (N_29162,N_22788,N_21028);
and U29163 (N_29163,N_21423,N_23224);
nand U29164 (N_29164,N_22053,N_23285);
and U29165 (N_29165,N_22080,N_21400);
and U29166 (N_29166,N_20908,N_21917);
nor U29167 (N_29167,N_23658,N_24460);
and U29168 (N_29168,N_22846,N_22628);
xnor U29169 (N_29169,N_21711,N_22263);
nand U29170 (N_29170,N_21721,N_23890);
or U29171 (N_29171,N_24535,N_22399);
nor U29172 (N_29172,N_22567,N_23349);
nand U29173 (N_29173,N_21463,N_23790);
nand U29174 (N_29174,N_22646,N_20594);
nand U29175 (N_29175,N_23579,N_20275);
or U29176 (N_29176,N_23714,N_22991);
or U29177 (N_29177,N_24883,N_20348);
nor U29178 (N_29178,N_20443,N_23062);
or U29179 (N_29179,N_24699,N_23713);
nand U29180 (N_29180,N_20110,N_24122);
nor U29181 (N_29181,N_21514,N_23605);
or U29182 (N_29182,N_21580,N_21666);
nand U29183 (N_29183,N_21253,N_20481);
nand U29184 (N_29184,N_24297,N_23543);
and U29185 (N_29185,N_23126,N_21548);
or U29186 (N_29186,N_20085,N_21551);
or U29187 (N_29187,N_20977,N_23628);
or U29188 (N_29188,N_20952,N_20533);
and U29189 (N_29189,N_23755,N_20471);
xor U29190 (N_29190,N_21313,N_20361);
or U29191 (N_29191,N_22668,N_24462);
xor U29192 (N_29192,N_21749,N_20600);
or U29193 (N_29193,N_22885,N_23239);
and U29194 (N_29194,N_21535,N_21434);
nand U29195 (N_29195,N_22780,N_24618);
nor U29196 (N_29196,N_22511,N_23463);
xnor U29197 (N_29197,N_24545,N_23659);
and U29198 (N_29198,N_20147,N_22620);
nand U29199 (N_29199,N_24884,N_24927);
nor U29200 (N_29200,N_23556,N_20373);
or U29201 (N_29201,N_23250,N_20371);
nand U29202 (N_29202,N_23877,N_23383);
nand U29203 (N_29203,N_24134,N_21229);
nand U29204 (N_29204,N_23767,N_24192);
nand U29205 (N_29205,N_24641,N_22858);
nand U29206 (N_29206,N_20274,N_23923);
nand U29207 (N_29207,N_21432,N_24214);
or U29208 (N_29208,N_23748,N_20877);
nor U29209 (N_29209,N_24972,N_20506);
nor U29210 (N_29210,N_23169,N_24414);
and U29211 (N_29211,N_22056,N_20942);
nand U29212 (N_29212,N_24439,N_23859);
nor U29213 (N_29213,N_20851,N_24028);
or U29214 (N_29214,N_21669,N_21819);
or U29215 (N_29215,N_23277,N_21384);
xnor U29216 (N_29216,N_23304,N_22899);
or U29217 (N_29217,N_23799,N_21126);
and U29218 (N_29218,N_20705,N_21148);
nand U29219 (N_29219,N_20375,N_24000);
nor U29220 (N_29220,N_20139,N_20058);
and U29221 (N_29221,N_21699,N_20451);
nor U29222 (N_29222,N_22060,N_22394);
nand U29223 (N_29223,N_20806,N_23836);
nand U29224 (N_29224,N_22172,N_20987);
or U29225 (N_29225,N_22631,N_21075);
or U29226 (N_29226,N_23263,N_23639);
nor U29227 (N_29227,N_22684,N_21330);
or U29228 (N_29228,N_23066,N_23546);
and U29229 (N_29229,N_23753,N_23284);
or U29230 (N_29230,N_22121,N_22096);
and U29231 (N_29231,N_22778,N_22997);
nor U29232 (N_29232,N_24310,N_23246);
nor U29233 (N_29233,N_24207,N_23855);
and U29234 (N_29234,N_21809,N_23570);
nand U29235 (N_29235,N_21188,N_23323);
and U29236 (N_29236,N_22880,N_23881);
or U29237 (N_29237,N_23497,N_20922);
and U29238 (N_29238,N_22828,N_21415);
or U29239 (N_29239,N_24081,N_23302);
nand U29240 (N_29240,N_24319,N_24862);
or U29241 (N_29241,N_21060,N_23682);
and U29242 (N_29242,N_24830,N_21328);
or U29243 (N_29243,N_21737,N_24922);
and U29244 (N_29244,N_24054,N_24726);
xnor U29245 (N_29245,N_21267,N_20463);
xor U29246 (N_29246,N_23250,N_21440);
nor U29247 (N_29247,N_22301,N_23462);
and U29248 (N_29248,N_23251,N_21579);
nor U29249 (N_29249,N_24599,N_24641);
and U29250 (N_29250,N_21817,N_23542);
xnor U29251 (N_29251,N_24571,N_21029);
nor U29252 (N_29252,N_24985,N_24504);
nor U29253 (N_29253,N_24170,N_23094);
xnor U29254 (N_29254,N_24956,N_24816);
nand U29255 (N_29255,N_22442,N_21656);
and U29256 (N_29256,N_22887,N_21778);
or U29257 (N_29257,N_24074,N_24171);
nand U29258 (N_29258,N_23673,N_21610);
or U29259 (N_29259,N_20640,N_23831);
nand U29260 (N_29260,N_24325,N_22253);
nor U29261 (N_29261,N_23372,N_24648);
nand U29262 (N_29262,N_22196,N_20508);
and U29263 (N_29263,N_21948,N_20707);
or U29264 (N_29264,N_21319,N_21878);
nor U29265 (N_29265,N_22280,N_23871);
and U29266 (N_29266,N_23724,N_20790);
or U29267 (N_29267,N_23676,N_22944);
nor U29268 (N_29268,N_24350,N_24108);
and U29269 (N_29269,N_20635,N_24274);
and U29270 (N_29270,N_20210,N_20347);
or U29271 (N_29271,N_21707,N_22404);
nand U29272 (N_29272,N_24847,N_24473);
or U29273 (N_29273,N_22856,N_24198);
or U29274 (N_29274,N_22940,N_23398);
nor U29275 (N_29275,N_24052,N_21742);
or U29276 (N_29276,N_23581,N_24029);
nor U29277 (N_29277,N_24491,N_24075);
nor U29278 (N_29278,N_22849,N_21716);
and U29279 (N_29279,N_22415,N_21648);
or U29280 (N_29280,N_24112,N_21234);
nand U29281 (N_29281,N_22601,N_23964);
nor U29282 (N_29282,N_24439,N_22622);
xor U29283 (N_29283,N_22052,N_22861);
nand U29284 (N_29284,N_21267,N_21152);
nor U29285 (N_29285,N_22600,N_24694);
or U29286 (N_29286,N_22081,N_24889);
nor U29287 (N_29287,N_21861,N_22556);
nor U29288 (N_29288,N_22647,N_21529);
and U29289 (N_29289,N_22529,N_23386);
xnor U29290 (N_29290,N_22791,N_24371);
xnor U29291 (N_29291,N_24230,N_20180);
and U29292 (N_29292,N_23282,N_24677);
and U29293 (N_29293,N_23650,N_22808);
nor U29294 (N_29294,N_23723,N_20304);
or U29295 (N_29295,N_20112,N_24669);
and U29296 (N_29296,N_21155,N_21836);
nand U29297 (N_29297,N_22274,N_20704);
and U29298 (N_29298,N_23951,N_24948);
and U29299 (N_29299,N_23997,N_20985);
nor U29300 (N_29300,N_23704,N_24241);
and U29301 (N_29301,N_20751,N_23418);
or U29302 (N_29302,N_21972,N_24678);
or U29303 (N_29303,N_23282,N_22722);
xor U29304 (N_29304,N_20741,N_22126);
nand U29305 (N_29305,N_21355,N_20622);
nand U29306 (N_29306,N_23808,N_21228);
or U29307 (N_29307,N_21368,N_21859);
and U29308 (N_29308,N_24048,N_20298);
or U29309 (N_29309,N_22593,N_20496);
xor U29310 (N_29310,N_22515,N_22923);
or U29311 (N_29311,N_23120,N_20264);
or U29312 (N_29312,N_20907,N_22269);
and U29313 (N_29313,N_20184,N_21061);
and U29314 (N_29314,N_23232,N_20282);
and U29315 (N_29315,N_23460,N_24439);
or U29316 (N_29316,N_21126,N_23083);
nor U29317 (N_29317,N_21149,N_24969);
xnor U29318 (N_29318,N_21879,N_24112);
or U29319 (N_29319,N_22433,N_23863);
and U29320 (N_29320,N_24521,N_23097);
or U29321 (N_29321,N_24179,N_20223);
or U29322 (N_29322,N_20612,N_21201);
nor U29323 (N_29323,N_23404,N_24912);
and U29324 (N_29324,N_23638,N_20039);
and U29325 (N_29325,N_23587,N_24247);
nor U29326 (N_29326,N_20452,N_22235);
nand U29327 (N_29327,N_21901,N_23380);
xor U29328 (N_29328,N_20387,N_22106);
and U29329 (N_29329,N_24985,N_23689);
and U29330 (N_29330,N_24084,N_21106);
or U29331 (N_29331,N_20686,N_20029);
and U29332 (N_29332,N_22919,N_20943);
nor U29333 (N_29333,N_23932,N_23350);
or U29334 (N_29334,N_24179,N_20834);
nor U29335 (N_29335,N_22007,N_22435);
or U29336 (N_29336,N_22821,N_23315);
and U29337 (N_29337,N_24769,N_22920);
nor U29338 (N_29338,N_21704,N_21728);
xnor U29339 (N_29339,N_21763,N_22598);
or U29340 (N_29340,N_24770,N_23598);
and U29341 (N_29341,N_24789,N_21021);
xor U29342 (N_29342,N_24110,N_21784);
and U29343 (N_29343,N_24808,N_24755);
nor U29344 (N_29344,N_20805,N_22417);
and U29345 (N_29345,N_23715,N_24179);
and U29346 (N_29346,N_20669,N_24102);
and U29347 (N_29347,N_20636,N_21422);
xnor U29348 (N_29348,N_24987,N_22876);
nand U29349 (N_29349,N_21629,N_24222);
nand U29350 (N_29350,N_20666,N_22995);
and U29351 (N_29351,N_24194,N_24002);
nand U29352 (N_29352,N_23343,N_23866);
or U29353 (N_29353,N_23638,N_21715);
nand U29354 (N_29354,N_20995,N_24123);
xor U29355 (N_29355,N_22049,N_24100);
nor U29356 (N_29356,N_20016,N_22149);
nand U29357 (N_29357,N_21261,N_22947);
xnor U29358 (N_29358,N_20612,N_21469);
nand U29359 (N_29359,N_23278,N_20290);
nand U29360 (N_29360,N_21607,N_24685);
and U29361 (N_29361,N_23247,N_24429);
nand U29362 (N_29362,N_23361,N_24441);
xor U29363 (N_29363,N_20081,N_20842);
nor U29364 (N_29364,N_22812,N_24320);
or U29365 (N_29365,N_20680,N_20129);
nor U29366 (N_29366,N_22145,N_21239);
nor U29367 (N_29367,N_23157,N_23914);
nand U29368 (N_29368,N_24095,N_23026);
and U29369 (N_29369,N_20512,N_24566);
nor U29370 (N_29370,N_24664,N_23921);
xnor U29371 (N_29371,N_21724,N_20815);
and U29372 (N_29372,N_24653,N_21967);
nor U29373 (N_29373,N_24023,N_23507);
and U29374 (N_29374,N_24894,N_20856);
nand U29375 (N_29375,N_24962,N_21365);
nor U29376 (N_29376,N_22265,N_21558);
or U29377 (N_29377,N_20182,N_23863);
nor U29378 (N_29378,N_23168,N_24167);
or U29379 (N_29379,N_22189,N_24201);
nor U29380 (N_29380,N_24205,N_22153);
or U29381 (N_29381,N_23347,N_24623);
nor U29382 (N_29382,N_21138,N_22311);
nor U29383 (N_29383,N_22969,N_24174);
xor U29384 (N_29384,N_22821,N_24742);
and U29385 (N_29385,N_24338,N_21743);
nor U29386 (N_29386,N_24359,N_20104);
and U29387 (N_29387,N_22306,N_23159);
or U29388 (N_29388,N_22230,N_22783);
nor U29389 (N_29389,N_22150,N_24011);
or U29390 (N_29390,N_24879,N_22288);
or U29391 (N_29391,N_24340,N_21702);
nand U29392 (N_29392,N_20140,N_22619);
nand U29393 (N_29393,N_21039,N_20509);
or U29394 (N_29394,N_24686,N_20686);
or U29395 (N_29395,N_22204,N_24096);
nand U29396 (N_29396,N_20594,N_21694);
nand U29397 (N_29397,N_21823,N_24566);
nand U29398 (N_29398,N_23583,N_20480);
or U29399 (N_29399,N_20300,N_22644);
nand U29400 (N_29400,N_20056,N_21131);
or U29401 (N_29401,N_21738,N_22651);
xnor U29402 (N_29402,N_22162,N_20085);
or U29403 (N_29403,N_21448,N_23006);
or U29404 (N_29404,N_21973,N_22399);
or U29405 (N_29405,N_23224,N_22801);
and U29406 (N_29406,N_20420,N_20920);
xor U29407 (N_29407,N_21043,N_24542);
nor U29408 (N_29408,N_21394,N_20299);
nand U29409 (N_29409,N_20542,N_23121);
nand U29410 (N_29410,N_24988,N_20346);
xor U29411 (N_29411,N_24309,N_21568);
or U29412 (N_29412,N_21166,N_22496);
or U29413 (N_29413,N_22436,N_21694);
and U29414 (N_29414,N_24288,N_23346);
nand U29415 (N_29415,N_23395,N_22885);
nor U29416 (N_29416,N_20243,N_20177);
nand U29417 (N_29417,N_22395,N_24416);
nor U29418 (N_29418,N_20520,N_20467);
nand U29419 (N_29419,N_21846,N_24942);
nand U29420 (N_29420,N_21792,N_23120);
and U29421 (N_29421,N_21689,N_23533);
or U29422 (N_29422,N_21087,N_23764);
nand U29423 (N_29423,N_20842,N_23730);
or U29424 (N_29424,N_20194,N_22706);
nand U29425 (N_29425,N_21786,N_22764);
nor U29426 (N_29426,N_23482,N_21175);
nor U29427 (N_29427,N_23995,N_20523);
or U29428 (N_29428,N_23629,N_21122);
nor U29429 (N_29429,N_24209,N_22389);
or U29430 (N_29430,N_22554,N_22376);
or U29431 (N_29431,N_22267,N_20107);
nor U29432 (N_29432,N_22225,N_22195);
nor U29433 (N_29433,N_23198,N_22251);
and U29434 (N_29434,N_20350,N_22380);
and U29435 (N_29435,N_20527,N_24863);
and U29436 (N_29436,N_23006,N_20806);
or U29437 (N_29437,N_20427,N_24174);
or U29438 (N_29438,N_22299,N_21243);
nand U29439 (N_29439,N_24496,N_23573);
nand U29440 (N_29440,N_21756,N_22452);
nand U29441 (N_29441,N_24640,N_23159);
nor U29442 (N_29442,N_23227,N_21570);
nand U29443 (N_29443,N_21326,N_24648);
xnor U29444 (N_29444,N_24060,N_20498);
or U29445 (N_29445,N_21746,N_23516);
or U29446 (N_29446,N_24557,N_21468);
nor U29447 (N_29447,N_22921,N_20844);
and U29448 (N_29448,N_22688,N_21991);
nor U29449 (N_29449,N_20452,N_20710);
xnor U29450 (N_29450,N_24046,N_20771);
and U29451 (N_29451,N_23911,N_21176);
and U29452 (N_29452,N_23794,N_23326);
or U29453 (N_29453,N_20209,N_20301);
nand U29454 (N_29454,N_20001,N_23294);
and U29455 (N_29455,N_24370,N_21527);
nand U29456 (N_29456,N_24702,N_21682);
or U29457 (N_29457,N_21141,N_22772);
and U29458 (N_29458,N_21605,N_20808);
or U29459 (N_29459,N_23334,N_24535);
or U29460 (N_29460,N_20958,N_22172);
and U29461 (N_29461,N_24326,N_20009);
or U29462 (N_29462,N_21794,N_22016);
nor U29463 (N_29463,N_22114,N_22391);
and U29464 (N_29464,N_24265,N_24033);
and U29465 (N_29465,N_20591,N_22463);
nand U29466 (N_29466,N_24837,N_22310);
nand U29467 (N_29467,N_24849,N_24695);
or U29468 (N_29468,N_23498,N_23869);
and U29469 (N_29469,N_22375,N_20657);
nand U29470 (N_29470,N_23265,N_22280);
nor U29471 (N_29471,N_20170,N_20017);
and U29472 (N_29472,N_23430,N_24726);
nand U29473 (N_29473,N_23833,N_20134);
and U29474 (N_29474,N_22202,N_22921);
or U29475 (N_29475,N_21763,N_24103);
or U29476 (N_29476,N_21111,N_21518);
nand U29477 (N_29477,N_23868,N_21347);
nand U29478 (N_29478,N_20101,N_22610);
or U29479 (N_29479,N_23206,N_23285);
xnor U29480 (N_29480,N_21883,N_23204);
and U29481 (N_29481,N_20246,N_21395);
nor U29482 (N_29482,N_20108,N_20962);
nand U29483 (N_29483,N_21602,N_24698);
xnor U29484 (N_29484,N_23530,N_21199);
and U29485 (N_29485,N_21908,N_23609);
and U29486 (N_29486,N_24818,N_22173);
nor U29487 (N_29487,N_20156,N_22558);
and U29488 (N_29488,N_21808,N_20743);
nand U29489 (N_29489,N_24362,N_21634);
nand U29490 (N_29490,N_20203,N_22587);
nand U29491 (N_29491,N_22306,N_24905);
and U29492 (N_29492,N_24174,N_24682);
and U29493 (N_29493,N_21890,N_21491);
or U29494 (N_29494,N_21675,N_23439);
and U29495 (N_29495,N_23879,N_23848);
and U29496 (N_29496,N_22344,N_24111);
nand U29497 (N_29497,N_21215,N_21650);
nand U29498 (N_29498,N_21297,N_21860);
nand U29499 (N_29499,N_22585,N_22373);
nor U29500 (N_29500,N_20882,N_24897);
nor U29501 (N_29501,N_22489,N_23934);
or U29502 (N_29502,N_22292,N_22617);
nand U29503 (N_29503,N_24167,N_20226);
nor U29504 (N_29504,N_22317,N_21102);
nor U29505 (N_29505,N_21376,N_24014);
and U29506 (N_29506,N_23503,N_21998);
or U29507 (N_29507,N_20092,N_22375);
nand U29508 (N_29508,N_21490,N_23533);
nor U29509 (N_29509,N_21134,N_24027);
or U29510 (N_29510,N_22428,N_21945);
nand U29511 (N_29511,N_20018,N_24542);
nor U29512 (N_29512,N_21882,N_22564);
and U29513 (N_29513,N_21577,N_23789);
nand U29514 (N_29514,N_21606,N_20157);
and U29515 (N_29515,N_22747,N_22310);
or U29516 (N_29516,N_24372,N_20701);
xnor U29517 (N_29517,N_20876,N_21491);
nand U29518 (N_29518,N_20475,N_21379);
and U29519 (N_29519,N_23806,N_21984);
and U29520 (N_29520,N_23378,N_21807);
and U29521 (N_29521,N_20861,N_20748);
nand U29522 (N_29522,N_23839,N_22369);
xor U29523 (N_29523,N_24963,N_21890);
or U29524 (N_29524,N_22301,N_23639);
nand U29525 (N_29525,N_20751,N_24390);
and U29526 (N_29526,N_22553,N_22012);
nor U29527 (N_29527,N_20735,N_24457);
nand U29528 (N_29528,N_21600,N_23986);
or U29529 (N_29529,N_21365,N_22643);
and U29530 (N_29530,N_23585,N_21087);
or U29531 (N_29531,N_23147,N_24078);
nor U29532 (N_29532,N_24794,N_22516);
nor U29533 (N_29533,N_20970,N_24996);
nor U29534 (N_29534,N_21843,N_22089);
xnor U29535 (N_29535,N_22811,N_20642);
and U29536 (N_29536,N_20006,N_22705);
or U29537 (N_29537,N_21123,N_24716);
or U29538 (N_29538,N_21707,N_20999);
and U29539 (N_29539,N_23172,N_22612);
or U29540 (N_29540,N_21700,N_20633);
and U29541 (N_29541,N_20980,N_21418);
nand U29542 (N_29542,N_20513,N_21488);
nand U29543 (N_29543,N_23688,N_22660);
and U29544 (N_29544,N_24476,N_20266);
nand U29545 (N_29545,N_21272,N_21207);
or U29546 (N_29546,N_24081,N_24335);
and U29547 (N_29547,N_20998,N_23734);
or U29548 (N_29548,N_22971,N_20306);
or U29549 (N_29549,N_21975,N_23910);
nand U29550 (N_29550,N_20339,N_24591);
and U29551 (N_29551,N_22712,N_21675);
nor U29552 (N_29552,N_20874,N_24448);
nor U29553 (N_29553,N_20078,N_21941);
and U29554 (N_29554,N_20020,N_23027);
nand U29555 (N_29555,N_20933,N_21707);
nand U29556 (N_29556,N_21076,N_20370);
and U29557 (N_29557,N_21196,N_21905);
and U29558 (N_29558,N_22969,N_24935);
nand U29559 (N_29559,N_23670,N_23322);
nand U29560 (N_29560,N_23709,N_20980);
or U29561 (N_29561,N_24506,N_22884);
nor U29562 (N_29562,N_20738,N_22623);
nor U29563 (N_29563,N_21018,N_23878);
and U29564 (N_29564,N_23032,N_24324);
nor U29565 (N_29565,N_22195,N_21150);
and U29566 (N_29566,N_22459,N_21816);
or U29567 (N_29567,N_22702,N_20111);
or U29568 (N_29568,N_20872,N_23066);
xor U29569 (N_29569,N_20678,N_24147);
or U29570 (N_29570,N_21144,N_22714);
or U29571 (N_29571,N_24814,N_23379);
nor U29572 (N_29572,N_23327,N_20326);
or U29573 (N_29573,N_24641,N_24080);
nor U29574 (N_29574,N_23884,N_23734);
nor U29575 (N_29575,N_24611,N_24854);
nor U29576 (N_29576,N_21626,N_24865);
nor U29577 (N_29577,N_21880,N_21153);
nor U29578 (N_29578,N_21680,N_20334);
xnor U29579 (N_29579,N_20587,N_24135);
nor U29580 (N_29580,N_21082,N_24182);
xor U29581 (N_29581,N_22935,N_20756);
nand U29582 (N_29582,N_24701,N_21924);
nor U29583 (N_29583,N_23286,N_24255);
nor U29584 (N_29584,N_21113,N_24537);
nand U29585 (N_29585,N_20202,N_23026);
nand U29586 (N_29586,N_21842,N_24306);
or U29587 (N_29587,N_21919,N_20394);
and U29588 (N_29588,N_21911,N_21939);
nor U29589 (N_29589,N_20755,N_23810);
and U29590 (N_29590,N_23647,N_22145);
and U29591 (N_29591,N_20375,N_24915);
nand U29592 (N_29592,N_24285,N_21828);
nand U29593 (N_29593,N_22137,N_20434);
and U29594 (N_29594,N_22652,N_21083);
and U29595 (N_29595,N_24142,N_21837);
or U29596 (N_29596,N_24275,N_20659);
nor U29597 (N_29597,N_21292,N_24614);
xnor U29598 (N_29598,N_20462,N_23837);
nor U29599 (N_29599,N_22506,N_22236);
nor U29600 (N_29600,N_23413,N_21202);
nor U29601 (N_29601,N_23942,N_21071);
xor U29602 (N_29602,N_24435,N_21341);
nor U29603 (N_29603,N_21683,N_22975);
or U29604 (N_29604,N_21651,N_20927);
nor U29605 (N_29605,N_22464,N_24785);
nand U29606 (N_29606,N_24948,N_23914);
or U29607 (N_29607,N_20363,N_24934);
nor U29608 (N_29608,N_23659,N_21596);
xnor U29609 (N_29609,N_23179,N_22675);
or U29610 (N_29610,N_23281,N_23758);
nand U29611 (N_29611,N_21586,N_24938);
nand U29612 (N_29612,N_20591,N_23042);
nand U29613 (N_29613,N_24804,N_23579);
and U29614 (N_29614,N_22319,N_24847);
and U29615 (N_29615,N_21284,N_20229);
or U29616 (N_29616,N_22437,N_21658);
xor U29617 (N_29617,N_21817,N_22416);
and U29618 (N_29618,N_20422,N_21559);
and U29619 (N_29619,N_21996,N_20223);
xor U29620 (N_29620,N_22655,N_23364);
or U29621 (N_29621,N_21505,N_21715);
or U29622 (N_29622,N_21225,N_22089);
nor U29623 (N_29623,N_21476,N_22892);
nand U29624 (N_29624,N_23904,N_21485);
or U29625 (N_29625,N_21551,N_24541);
or U29626 (N_29626,N_21132,N_21504);
nor U29627 (N_29627,N_20589,N_24579);
nor U29628 (N_29628,N_23834,N_21921);
and U29629 (N_29629,N_24699,N_20906);
xnor U29630 (N_29630,N_24082,N_22114);
nand U29631 (N_29631,N_20398,N_22065);
nand U29632 (N_29632,N_24498,N_20521);
nand U29633 (N_29633,N_20324,N_23658);
nor U29634 (N_29634,N_24724,N_23001);
nor U29635 (N_29635,N_22360,N_24212);
nor U29636 (N_29636,N_21921,N_20431);
and U29637 (N_29637,N_20277,N_24621);
or U29638 (N_29638,N_20819,N_20873);
and U29639 (N_29639,N_24828,N_23892);
xnor U29640 (N_29640,N_23277,N_24597);
and U29641 (N_29641,N_23491,N_23203);
nor U29642 (N_29642,N_24146,N_20756);
and U29643 (N_29643,N_23536,N_21252);
nor U29644 (N_29644,N_21994,N_24175);
or U29645 (N_29645,N_23238,N_20620);
nand U29646 (N_29646,N_24800,N_24485);
xor U29647 (N_29647,N_22882,N_20170);
and U29648 (N_29648,N_23568,N_24801);
nor U29649 (N_29649,N_20650,N_22479);
xor U29650 (N_29650,N_21447,N_20742);
nand U29651 (N_29651,N_21743,N_24722);
nor U29652 (N_29652,N_24556,N_20843);
nand U29653 (N_29653,N_23489,N_20903);
nand U29654 (N_29654,N_22994,N_20329);
nor U29655 (N_29655,N_22771,N_23752);
and U29656 (N_29656,N_23519,N_20346);
and U29657 (N_29657,N_20416,N_24257);
and U29658 (N_29658,N_22242,N_24913);
and U29659 (N_29659,N_20477,N_22227);
nand U29660 (N_29660,N_22794,N_24012);
or U29661 (N_29661,N_22847,N_24085);
nor U29662 (N_29662,N_20185,N_22337);
nor U29663 (N_29663,N_22246,N_20994);
or U29664 (N_29664,N_21038,N_22048);
xnor U29665 (N_29665,N_23671,N_22964);
or U29666 (N_29666,N_22164,N_24742);
or U29667 (N_29667,N_23114,N_22165);
and U29668 (N_29668,N_20173,N_22283);
and U29669 (N_29669,N_22967,N_22338);
and U29670 (N_29670,N_23997,N_21169);
nand U29671 (N_29671,N_21021,N_22909);
and U29672 (N_29672,N_23062,N_22472);
nand U29673 (N_29673,N_23049,N_21733);
or U29674 (N_29674,N_20209,N_24829);
nor U29675 (N_29675,N_21035,N_24946);
and U29676 (N_29676,N_22946,N_22318);
and U29677 (N_29677,N_22850,N_22403);
nand U29678 (N_29678,N_22096,N_23679);
nor U29679 (N_29679,N_24108,N_24531);
xor U29680 (N_29680,N_24029,N_21123);
nor U29681 (N_29681,N_20957,N_22647);
nand U29682 (N_29682,N_20940,N_21260);
and U29683 (N_29683,N_23777,N_22746);
or U29684 (N_29684,N_22798,N_23949);
and U29685 (N_29685,N_21144,N_22589);
xor U29686 (N_29686,N_22740,N_21837);
nor U29687 (N_29687,N_22460,N_23054);
and U29688 (N_29688,N_22306,N_22668);
nand U29689 (N_29689,N_24873,N_21371);
or U29690 (N_29690,N_22202,N_23350);
xor U29691 (N_29691,N_23244,N_24658);
nor U29692 (N_29692,N_22427,N_23513);
and U29693 (N_29693,N_24824,N_24628);
nand U29694 (N_29694,N_22240,N_23378);
nand U29695 (N_29695,N_23955,N_21911);
xor U29696 (N_29696,N_20986,N_24353);
and U29697 (N_29697,N_22977,N_24981);
nor U29698 (N_29698,N_23010,N_20714);
nand U29699 (N_29699,N_24387,N_20954);
or U29700 (N_29700,N_20892,N_23372);
nand U29701 (N_29701,N_21807,N_23493);
nor U29702 (N_29702,N_23044,N_21543);
or U29703 (N_29703,N_23212,N_20743);
xor U29704 (N_29704,N_23794,N_21720);
and U29705 (N_29705,N_21734,N_20127);
or U29706 (N_29706,N_24203,N_20119);
nand U29707 (N_29707,N_23433,N_24311);
or U29708 (N_29708,N_20796,N_23677);
or U29709 (N_29709,N_24057,N_24443);
or U29710 (N_29710,N_22932,N_20081);
nand U29711 (N_29711,N_23376,N_23055);
nor U29712 (N_29712,N_21161,N_22381);
and U29713 (N_29713,N_20552,N_22457);
nor U29714 (N_29714,N_23871,N_24274);
xor U29715 (N_29715,N_24268,N_21843);
nor U29716 (N_29716,N_21438,N_24429);
xor U29717 (N_29717,N_20987,N_22574);
nand U29718 (N_29718,N_20716,N_21932);
nand U29719 (N_29719,N_24120,N_22018);
xnor U29720 (N_29720,N_23629,N_23006);
nor U29721 (N_29721,N_21586,N_20622);
nand U29722 (N_29722,N_22359,N_24756);
or U29723 (N_29723,N_22318,N_24957);
or U29724 (N_29724,N_24660,N_21602);
nor U29725 (N_29725,N_22200,N_21460);
and U29726 (N_29726,N_23351,N_21270);
and U29727 (N_29727,N_22450,N_23920);
nand U29728 (N_29728,N_20709,N_24141);
or U29729 (N_29729,N_23608,N_21819);
nand U29730 (N_29730,N_22265,N_22651);
or U29731 (N_29731,N_20605,N_20864);
nand U29732 (N_29732,N_21037,N_24553);
nor U29733 (N_29733,N_23686,N_23443);
or U29734 (N_29734,N_23655,N_23078);
or U29735 (N_29735,N_21857,N_21914);
nor U29736 (N_29736,N_22122,N_23939);
and U29737 (N_29737,N_22991,N_20141);
or U29738 (N_29738,N_23159,N_22323);
nor U29739 (N_29739,N_21625,N_24311);
nand U29740 (N_29740,N_21412,N_24091);
nor U29741 (N_29741,N_24246,N_23647);
and U29742 (N_29742,N_23801,N_21584);
nand U29743 (N_29743,N_21777,N_23665);
nor U29744 (N_29744,N_21478,N_23296);
and U29745 (N_29745,N_23724,N_22609);
nand U29746 (N_29746,N_24007,N_23812);
or U29747 (N_29747,N_22189,N_22311);
nor U29748 (N_29748,N_23062,N_24092);
nor U29749 (N_29749,N_20532,N_22022);
and U29750 (N_29750,N_22649,N_22741);
or U29751 (N_29751,N_20272,N_22594);
xor U29752 (N_29752,N_24255,N_22217);
or U29753 (N_29753,N_22906,N_23220);
or U29754 (N_29754,N_21468,N_20812);
nor U29755 (N_29755,N_21264,N_22958);
xor U29756 (N_29756,N_23345,N_23355);
or U29757 (N_29757,N_23889,N_22356);
nor U29758 (N_29758,N_24537,N_20573);
xor U29759 (N_29759,N_23063,N_23930);
nor U29760 (N_29760,N_20358,N_24748);
or U29761 (N_29761,N_23537,N_20512);
nor U29762 (N_29762,N_22047,N_21948);
and U29763 (N_29763,N_23248,N_22344);
nor U29764 (N_29764,N_21670,N_22430);
or U29765 (N_29765,N_23797,N_24742);
xor U29766 (N_29766,N_21935,N_24529);
and U29767 (N_29767,N_23439,N_24913);
nor U29768 (N_29768,N_22755,N_20067);
nor U29769 (N_29769,N_20938,N_21285);
nand U29770 (N_29770,N_22491,N_23549);
xnor U29771 (N_29771,N_23917,N_20168);
and U29772 (N_29772,N_23353,N_20306);
and U29773 (N_29773,N_22736,N_23050);
or U29774 (N_29774,N_24312,N_22102);
or U29775 (N_29775,N_20596,N_24419);
or U29776 (N_29776,N_22489,N_21844);
or U29777 (N_29777,N_23478,N_22206);
nor U29778 (N_29778,N_24632,N_21378);
and U29779 (N_29779,N_20481,N_21516);
xor U29780 (N_29780,N_22136,N_23990);
or U29781 (N_29781,N_24096,N_21914);
nand U29782 (N_29782,N_22057,N_24089);
nor U29783 (N_29783,N_23323,N_24222);
and U29784 (N_29784,N_20978,N_23265);
or U29785 (N_29785,N_21044,N_20003);
or U29786 (N_29786,N_24763,N_22226);
nor U29787 (N_29787,N_23874,N_23445);
xnor U29788 (N_29788,N_24754,N_23138);
xor U29789 (N_29789,N_23595,N_23856);
xor U29790 (N_29790,N_20341,N_23932);
and U29791 (N_29791,N_20362,N_23593);
nor U29792 (N_29792,N_21368,N_24211);
or U29793 (N_29793,N_20592,N_21705);
nor U29794 (N_29794,N_24839,N_24153);
nand U29795 (N_29795,N_21964,N_23561);
nand U29796 (N_29796,N_21145,N_21603);
nor U29797 (N_29797,N_22728,N_22084);
nand U29798 (N_29798,N_22348,N_23031);
nand U29799 (N_29799,N_21926,N_24616);
nor U29800 (N_29800,N_23474,N_21081);
xor U29801 (N_29801,N_22872,N_21251);
nand U29802 (N_29802,N_23907,N_20914);
or U29803 (N_29803,N_22672,N_21739);
or U29804 (N_29804,N_24736,N_21456);
nand U29805 (N_29805,N_23530,N_24725);
nor U29806 (N_29806,N_24632,N_22275);
nor U29807 (N_29807,N_24679,N_24577);
or U29808 (N_29808,N_20556,N_24114);
nand U29809 (N_29809,N_21906,N_24013);
and U29810 (N_29810,N_20598,N_22780);
nor U29811 (N_29811,N_20948,N_22326);
nand U29812 (N_29812,N_21650,N_21470);
or U29813 (N_29813,N_21915,N_20290);
nand U29814 (N_29814,N_24311,N_24457);
nand U29815 (N_29815,N_21422,N_24470);
nor U29816 (N_29816,N_24124,N_21736);
and U29817 (N_29817,N_22298,N_21801);
or U29818 (N_29818,N_23283,N_21557);
nor U29819 (N_29819,N_23086,N_22230);
xnor U29820 (N_29820,N_23934,N_23078);
xnor U29821 (N_29821,N_20054,N_23528);
nor U29822 (N_29822,N_23457,N_24464);
and U29823 (N_29823,N_21611,N_24112);
nor U29824 (N_29824,N_24982,N_22107);
nor U29825 (N_29825,N_21800,N_21950);
nor U29826 (N_29826,N_23691,N_24058);
nor U29827 (N_29827,N_20223,N_22847);
and U29828 (N_29828,N_20084,N_23474);
or U29829 (N_29829,N_22590,N_21136);
nand U29830 (N_29830,N_24739,N_21471);
nor U29831 (N_29831,N_22049,N_21030);
or U29832 (N_29832,N_22893,N_21694);
nor U29833 (N_29833,N_23949,N_23569);
and U29834 (N_29834,N_21529,N_22723);
and U29835 (N_29835,N_24106,N_21483);
nor U29836 (N_29836,N_21785,N_22399);
or U29837 (N_29837,N_21005,N_24781);
or U29838 (N_29838,N_20738,N_20013);
nor U29839 (N_29839,N_20233,N_20221);
nand U29840 (N_29840,N_23817,N_20721);
or U29841 (N_29841,N_22719,N_24059);
or U29842 (N_29842,N_20076,N_22394);
or U29843 (N_29843,N_23943,N_23141);
nand U29844 (N_29844,N_21207,N_24520);
or U29845 (N_29845,N_20211,N_21980);
nand U29846 (N_29846,N_24355,N_21524);
and U29847 (N_29847,N_22031,N_21359);
nand U29848 (N_29848,N_23873,N_21596);
or U29849 (N_29849,N_21998,N_22239);
or U29850 (N_29850,N_20848,N_22861);
and U29851 (N_29851,N_24659,N_23105);
or U29852 (N_29852,N_22689,N_23351);
nand U29853 (N_29853,N_23967,N_23223);
or U29854 (N_29854,N_23948,N_22552);
nand U29855 (N_29855,N_24865,N_21936);
xnor U29856 (N_29856,N_24783,N_23081);
and U29857 (N_29857,N_21916,N_23929);
nand U29858 (N_29858,N_21236,N_20164);
nand U29859 (N_29859,N_24973,N_21817);
nand U29860 (N_29860,N_23618,N_21091);
or U29861 (N_29861,N_23028,N_23622);
nand U29862 (N_29862,N_20552,N_21945);
or U29863 (N_29863,N_21557,N_20216);
nor U29864 (N_29864,N_22273,N_20861);
or U29865 (N_29865,N_22915,N_22493);
or U29866 (N_29866,N_20762,N_23452);
and U29867 (N_29867,N_23149,N_20115);
nand U29868 (N_29868,N_20277,N_22630);
or U29869 (N_29869,N_24133,N_21195);
nor U29870 (N_29870,N_24244,N_23023);
nor U29871 (N_29871,N_21612,N_24072);
nand U29872 (N_29872,N_20707,N_24198);
nor U29873 (N_29873,N_24825,N_24964);
and U29874 (N_29874,N_20773,N_20747);
nand U29875 (N_29875,N_22020,N_24335);
xnor U29876 (N_29876,N_22212,N_22642);
or U29877 (N_29877,N_20512,N_24558);
and U29878 (N_29878,N_23123,N_20892);
or U29879 (N_29879,N_23510,N_24200);
nor U29880 (N_29880,N_23848,N_20017);
and U29881 (N_29881,N_23579,N_20661);
xor U29882 (N_29882,N_20959,N_24191);
nor U29883 (N_29883,N_20381,N_24356);
nor U29884 (N_29884,N_21113,N_21026);
xor U29885 (N_29885,N_22362,N_24732);
xor U29886 (N_29886,N_23897,N_23282);
and U29887 (N_29887,N_23037,N_23383);
nor U29888 (N_29888,N_24814,N_22970);
and U29889 (N_29889,N_24354,N_23143);
or U29890 (N_29890,N_23333,N_20537);
and U29891 (N_29891,N_22194,N_23170);
or U29892 (N_29892,N_23604,N_20815);
nand U29893 (N_29893,N_22820,N_22893);
xor U29894 (N_29894,N_21656,N_23615);
and U29895 (N_29895,N_20635,N_20540);
and U29896 (N_29896,N_24988,N_21955);
and U29897 (N_29897,N_20226,N_21588);
or U29898 (N_29898,N_21683,N_20262);
nand U29899 (N_29899,N_20720,N_21904);
and U29900 (N_29900,N_21236,N_24875);
xor U29901 (N_29901,N_24062,N_22119);
and U29902 (N_29902,N_20540,N_24516);
nand U29903 (N_29903,N_21562,N_22747);
nand U29904 (N_29904,N_23530,N_22315);
nand U29905 (N_29905,N_23093,N_20122);
nor U29906 (N_29906,N_23976,N_20966);
nor U29907 (N_29907,N_24055,N_22131);
nand U29908 (N_29908,N_20286,N_24767);
or U29909 (N_29909,N_21704,N_20349);
xnor U29910 (N_29910,N_23660,N_21217);
xnor U29911 (N_29911,N_24489,N_23184);
nor U29912 (N_29912,N_20717,N_24522);
nor U29913 (N_29913,N_24149,N_22947);
or U29914 (N_29914,N_24480,N_24612);
and U29915 (N_29915,N_23006,N_22044);
nor U29916 (N_29916,N_21703,N_23842);
nand U29917 (N_29917,N_20380,N_22189);
nand U29918 (N_29918,N_23651,N_22733);
or U29919 (N_29919,N_23949,N_23454);
and U29920 (N_29920,N_20634,N_20481);
or U29921 (N_29921,N_21117,N_24040);
xnor U29922 (N_29922,N_21336,N_24632);
nand U29923 (N_29923,N_24301,N_21036);
nand U29924 (N_29924,N_23737,N_21601);
xnor U29925 (N_29925,N_21613,N_20414);
nand U29926 (N_29926,N_21864,N_21768);
nor U29927 (N_29927,N_22604,N_21640);
nor U29928 (N_29928,N_23313,N_20969);
and U29929 (N_29929,N_21736,N_22379);
nand U29930 (N_29930,N_21398,N_24948);
or U29931 (N_29931,N_23500,N_24796);
or U29932 (N_29932,N_22747,N_22725);
nand U29933 (N_29933,N_21979,N_21335);
nand U29934 (N_29934,N_23662,N_22375);
or U29935 (N_29935,N_24768,N_24322);
nand U29936 (N_29936,N_22778,N_24322);
nand U29937 (N_29937,N_24674,N_21254);
and U29938 (N_29938,N_24665,N_22680);
or U29939 (N_29939,N_22425,N_23720);
and U29940 (N_29940,N_22413,N_22280);
or U29941 (N_29941,N_23390,N_24937);
nor U29942 (N_29942,N_21064,N_23277);
xor U29943 (N_29943,N_23559,N_21221);
and U29944 (N_29944,N_20253,N_20414);
nor U29945 (N_29945,N_23536,N_24757);
or U29946 (N_29946,N_21175,N_22424);
xor U29947 (N_29947,N_22188,N_20675);
nand U29948 (N_29948,N_22450,N_20698);
and U29949 (N_29949,N_20617,N_20640);
nand U29950 (N_29950,N_22024,N_22982);
and U29951 (N_29951,N_21941,N_24855);
nor U29952 (N_29952,N_21793,N_23105);
nor U29953 (N_29953,N_24843,N_22744);
nor U29954 (N_29954,N_23945,N_21090);
xor U29955 (N_29955,N_21657,N_22580);
and U29956 (N_29956,N_23021,N_23669);
or U29957 (N_29957,N_23064,N_22080);
nor U29958 (N_29958,N_23768,N_24337);
nand U29959 (N_29959,N_21457,N_23321);
and U29960 (N_29960,N_24572,N_23700);
nor U29961 (N_29961,N_20139,N_20736);
and U29962 (N_29962,N_22696,N_20012);
nor U29963 (N_29963,N_24282,N_23097);
nor U29964 (N_29964,N_22309,N_22264);
xnor U29965 (N_29965,N_21378,N_22249);
nand U29966 (N_29966,N_24012,N_21703);
and U29967 (N_29967,N_24596,N_24510);
or U29968 (N_29968,N_24985,N_24314);
or U29969 (N_29969,N_23750,N_24622);
and U29970 (N_29970,N_23666,N_21510);
or U29971 (N_29971,N_24105,N_22088);
and U29972 (N_29972,N_22493,N_24456);
nor U29973 (N_29973,N_24844,N_24638);
nand U29974 (N_29974,N_23516,N_20315);
nand U29975 (N_29975,N_24067,N_21079);
nor U29976 (N_29976,N_20930,N_22680);
or U29977 (N_29977,N_21236,N_20262);
and U29978 (N_29978,N_23236,N_24795);
or U29979 (N_29979,N_21616,N_22394);
and U29980 (N_29980,N_20026,N_23072);
xnor U29981 (N_29981,N_21061,N_22879);
nand U29982 (N_29982,N_24003,N_24142);
nor U29983 (N_29983,N_23255,N_23327);
and U29984 (N_29984,N_23132,N_23973);
or U29985 (N_29985,N_24408,N_24066);
nor U29986 (N_29986,N_21016,N_20744);
nand U29987 (N_29987,N_20203,N_24698);
nand U29988 (N_29988,N_21917,N_23707);
xnor U29989 (N_29989,N_23328,N_23507);
xnor U29990 (N_29990,N_24240,N_20899);
and U29991 (N_29991,N_24790,N_23938);
nor U29992 (N_29992,N_24793,N_22492);
and U29993 (N_29993,N_24308,N_21327);
nand U29994 (N_29994,N_23564,N_22407);
nor U29995 (N_29995,N_23201,N_24727);
or U29996 (N_29996,N_24403,N_21652);
or U29997 (N_29997,N_24382,N_20472);
nor U29998 (N_29998,N_23523,N_22335);
or U29999 (N_29999,N_21897,N_22837);
nor UO_0 (O_0,N_29662,N_27988);
and UO_1 (O_1,N_27656,N_25741);
nand UO_2 (O_2,N_27922,N_29402);
and UO_3 (O_3,N_28468,N_29442);
and UO_4 (O_4,N_26159,N_29999);
or UO_5 (O_5,N_25112,N_25593);
nand UO_6 (O_6,N_29724,N_25721);
nand UO_7 (O_7,N_27954,N_26845);
or UO_8 (O_8,N_26130,N_27130);
or UO_9 (O_9,N_25638,N_29904);
nand UO_10 (O_10,N_26374,N_26734);
or UO_11 (O_11,N_27859,N_27305);
nand UO_12 (O_12,N_25683,N_29886);
or UO_13 (O_13,N_26501,N_28877);
and UO_14 (O_14,N_29756,N_26471);
and UO_15 (O_15,N_29706,N_29197);
nand UO_16 (O_16,N_25830,N_25273);
or UO_17 (O_17,N_26521,N_29859);
xnor UO_18 (O_18,N_26210,N_27927);
and UO_19 (O_19,N_27022,N_28371);
or UO_20 (O_20,N_25716,N_25911);
xnor UO_21 (O_21,N_29500,N_26138);
nor UO_22 (O_22,N_27473,N_29989);
nand UO_23 (O_23,N_28958,N_29173);
and UO_24 (O_24,N_26476,N_26446);
nand UO_25 (O_25,N_29494,N_27843);
or UO_26 (O_26,N_26444,N_26127);
and UO_27 (O_27,N_26518,N_26408);
or UO_28 (O_28,N_26566,N_26744);
nand UO_29 (O_29,N_28467,N_26601);
xor UO_30 (O_30,N_27402,N_29757);
nand UO_31 (O_31,N_25857,N_26477);
nand UO_32 (O_32,N_29169,N_29217);
nand UO_33 (O_33,N_26083,N_25447);
nor UO_34 (O_34,N_25811,N_25012);
nor UO_35 (O_35,N_27410,N_25434);
and UO_36 (O_36,N_25587,N_28037);
nand UO_37 (O_37,N_25008,N_25933);
nor UO_38 (O_38,N_26202,N_26814);
nand UO_39 (O_39,N_27379,N_29552);
or UO_40 (O_40,N_25757,N_26841);
nor UO_41 (O_41,N_29103,N_29518);
nand UO_42 (O_42,N_25411,N_26665);
nand UO_43 (O_43,N_25069,N_26214);
and UO_44 (O_44,N_29378,N_28179);
and UO_45 (O_45,N_26591,N_29389);
nor UO_46 (O_46,N_27467,N_29791);
or UO_47 (O_47,N_26321,N_27575);
and UO_48 (O_48,N_28053,N_29594);
or UO_49 (O_49,N_29455,N_29079);
and UO_50 (O_50,N_28665,N_29767);
nand UO_51 (O_51,N_25272,N_25771);
or UO_52 (O_52,N_29581,N_27849);
and UO_53 (O_53,N_27340,N_25891);
nand UO_54 (O_54,N_25547,N_25583);
xor UO_55 (O_55,N_28662,N_25235);
nor UO_56 (O_56,N_26807,N_27027);
nand UO_57 (O_57,N_28507,N_28527);
and UO_58 (O_58,N_29208,N_28304);
xnor UO_59 (O_59,N_25499,N_25868);
and UO_60 (O_60,N_28533,N_26515);
and UO_61 (O_61,N_26301,N_28860);
nand UO_62 (O_62,N_27227,N_26910);
nor UO_63 (O_63,N_26342,N_27406);
and UO_64 (O_64,N_29038,N_27049);
nand UO_65 (O_65,N_27011,N_25849);
or UO_66 (O_66,N_25257,N_25739);
nor UO_67 (O_67,N_28157,N_27720);
nand UO_68 (O_68,N_29120,N_29356);
or UO_69 (O_69,N_27142,N_25347);
nor UO_70 (O_70,N_27599,N_26816);
nand UO_71 (O_71,N_28672,N_28350);
and UO_72 (O_72,N_25336,N_27616);
or UO_73 (O_73,N_28504,N_29396);
nor UO_74 (O_74,N_29776,N_28045);
nand UO_75 (O_75,N_26421,N_26035);
nand UO_76 (O_76,N_26672,N_29002);
nand UO_77 (O_77,N_29915,N_25128);
or UO_78 (O_78,N_28586,N_26865);
and UO_79 (O_79,N_25253,N_28992);
nand UO_80 (O_80,N_26215,N_28510);
nand UO_81 (O_81,N_27491,N_25743);
nand UO_82 (O_82,N_29101,N_25668);
nor UO_83 (O_83,N_26324,N_26074);
nor UO_84 (O_84,N_28006,N_25546);
nand UO_85 (O_85,N_29407,N_25774);
nand UO_86 (O_86,N_26454,N_26249);
nor UO_87 (O_87,N_28077,N_29582);
or UO_88 (O_88,N_25221,N_25027);
or UO_89 (O_89,N_29602,N_25642);
nand UO_90 (O_90,N_28039,N_27837);
or UO_91 (O_91,N_29945,N_27053);
nand UO_92 (O_92,N_25091,N_25875);
or UO_93 (O_93,N_26503,N_29109);
xor UO_94 (O_94,N_28286,N_28149);
nor UO_95 (O_95,N_28060,N_26191);
or UO_96 (O_96,N_25533,N_27790);
nor UO_97 (O_97,N_28838,N_27994);
and UO_98 (O_98,N_25985,N_27427);
nand UO_99 (O_99,N_25972,N_28904);
and UO_100 (O_100,N_27945,N_27315);
nor UO_101 (O_101,N_28983,N_25711);
nand UO_102 (O_102,N_25828,N_26493);
and UO_103 (O_103,N_28748,N_27664);
or UO_104 (O_104,N_28397,N_25841);
and UO_105 (O_105,N_26160,N_26611);
xnor UO_106 (O_106,N_25935,N_27594);
nand UO_107 (O_107,N_25775,N_28800);
xnor UO_108 (O_108,N_27505,N_26252);
and UO_109 (O_109,N_26176,N_27546);
and UO_110 (O_110,N_28516,N_29976);
or UO_111 (O_111,N_26802,N_26464);
nand UO_112 (O_112,N_28895,N_25766);
nor UO_113 (O_113,N_25872,N_25964);
or UO_114 (O_114,N_27489,N_28757);
or UO_115 (O_115,N_25368,N_26738);
or UO_116 (O_116,N_28046,N_28688);
or UO_117 (O_117,N_29764,N_27797);
nor UO_118 (O_118,N_29158,N_28754);
xor UO_119 (O_119,N_28383,N_27221);
or UO_120 (O_120,N_26212,N_27885);
or UO_121 (O_121,N_28065,N_28898);
or UO_122 (O_122,N_27151,N_28971);
or UO_123 (O_123,N_25908,N_28148);
and UO_124 (O_124,N_27858,N_28576);
and UO_125 (O_125,N_26415,N_29012);
nor UO_126 (O_126,N_27219,N_26383);
and UO_127 (O_127,N_26375,N_25013);
and UO_128 (O_128,N_25239,N_26288);
nor UO_129 (O_129,N_27152,N_28433);
nand UO_130 (O_130,N_29729,N_27228);
nand UO_131 (O_131,N_29974,N_28613);
nand UO_132 (O_132,N_27218,N_25607);
and UO_133 (O_133,N_29473,N_29577);
or UO_134 (O_134,N_25051,N_25374);
or UO_135 (O_135,N_25586,N_29133);
nor UO_136 (O_136,N_29256,N_26875);
xor UO_137 (O_137,N_25408,N_27289);
and UO_138 (O_138,N_27108,N_25243);
or UO_139 (O_139,N_28851,N_27123);
nor UO_140 (O_140,N_28768,N_25528);
nor UO_141 (O_141,N_27019,N_27112);
nor UO_142 (O_142,N_27171,N_25855);
nor UO_143 (O_143,N_26692,N_29227);
xor UO_144 (O_144,N_28170,N_25287);
xnor UO_145 (O_145,N_26380,N_29631);
nor UO_146 (O_146,N_27192,N_29470);
xor UO_147 (O_147,N_25302,N_26144);
or UO_148 (O_148,N_25529,N_27155);
and UO_149 (O_149,N_29211,N_27765);
and UO_150 (O_150,N_25929,N_29786);
nand UO_151 (O_151,N_28025,N_29635);
nor UO_152 (O_152,N_29045,N_27832);
nor UO_153 (O_153,N_27989,N_27015);
or UO_154 (O_154,N_26676,N_26850);
nor UO_155 (O_155,N_29275,N_26347);
or UO_156 (O_156,N_28685,N_26399);
and UO_157 (O_157,N_26681,N_29875);
nor UO_158 (O_158,N_28677,N_28874);
nand UO_159 (O_159,N_27475,N_27821);
xor UO_160 (O_160,N_27697,N_28044);
nand UO_161 (O_161,N_28028,N_25817);
and UO_162 (O_162,N_29629,N_29474);
or UO_163 (O_163,N_29873,N_26898);
and UO_164 (O_164,N_26156,N_27190);
nand UO_165 (O_165,N_26588,N_26864);
nor UO_166 (O_166,N_25399,N_27908);
or UO_167 (O_167,N_29469,N_25921);
nor UO_168 (O_168,N_29841,N_29434);
nand UO_169 (O_169,N_29740,N_27972);
nor UO_170 (O_170,N_29130,N_27414);
and UO_171 (O_171,N_25264,N_27604);
nor UO_172 (O_172,N_28119,N_26021);
nor UO_173 (O_173,N_27668,N_25691);
nand UO_174 (O_174,N_28325,N_29082);
xor UO_175 (O_175,N_29060,N_28223);
and UO_176 (O_176,N_28731,N_26473);
or UO_177 (O_177,N_28809,N_25108);
or UO_178 (O_178,N_25147,N_28461);
nand UO_179 (O_179,N_25009,N_26360);
nand UO_180 (O_180,N_29210,N_25641);
xnor UO_181 (O_181,N_27609,N_26287);
nand UO_182 (O_182,N_27495,N_27570);
and UO_183 (O_183,N_29921,N_27970);
nand UO_184 (O_184,N_27258,N_26059);
nand UO_185 (O_185,N_25366,N_27671);
xnor UO_186 (O_186,N_28298,N_29897);
or UO_187 (O_187,N_27029,N_27783);
and UO_188 (O_188,N_28808,N_25596);
nor UO_189 (O_189,N_29298,N_26038);
nor UO_190 (O_190,N_26553,N_29182);
and UO_191 (O_191,N_28364,N_26036);
nand UO_192 (O_192,N_28583,N_26517);
nor UO_193 (O_193,N_27685,N_29061);
or UO_194 (O_194,N_29016,N_26479);
and UO_195 (O_195,N_27509,N_29471);
or UO_196 (O_196,N_28084,N_27545);
nor UO_197 (O_197,N_26972,N_25297);
nand UO_198 (O_198,N_27909,N_25920);
xor UO_199 (O_199,N_29331,N_25567);
or UO_200 (O_200,N_26815,N_27349);
nand UO_201 (O_201,N_25390,N_26629);
or UO_202 (O_202,N_27533,N_25669);
and UO_203 (O_203,N_27176,N_26339);
and UO_204 (O_204,N_26549,N_26662);
nor UO_205 (O_205,N_27739,N_26142);
and UO_206 (O_206,N_26872,N_28872);
nor UO_207 (O_207,N_27380,N_26686);
or UO_208 (O_208,N_25573,N_26818);
nand UO_209 (O_209,N_29531,N_26999);
xnor UO_210 (O_210,N_28627,N_26861);
nand UO_211 (O_211,N_25444,N_26235);
nor UO_212 (O_212,N_25248,N_27088);
and UO_213 (O_213,N_29860,N_28994);
xor UO_214 (O_214,N_29144,N_27245);
nor UO_215 (O_215,N_26668,N_26436);
xor UO_216 (O_216,N_29498,N_25196);
or UO_217 (O_217,N_27078,N_29542);
nand UO_218 (O_218,N_26076,N_28790);
xnor UO_219 (O_219,N_27200,N_25667);
and UO_220 (O_220,N_29185,N_29485);
and UO_221 (O_221,N_28753,N_28193);
xnor UO_222 (O_222,N_27198,N_26948);
and UO_223 (O_223,N_29847,N_26704);
nand UO_224 (O_224,N_28332,N_29838);
nor UO_225 (O_225,N_29183,N_29885);
xnor UO_226 (O_226,N_26381,N_27232);
nand UO_227 (O_227,N_27725,N_29328);
xnor UO_228 (O_228,N_29076,N_28712);
or UO_229 (O_229,N_29655,N_26931);
or UO_230 (O_230,N_25658,N_25631);
and UO_231 (O_231,N_28128,N_29159);
nor UO_232 (O_232,N_29647,N_25662);
nand UO_233 (O_233,N_25863,N_29285);
nand UO_234 (O_234,N_26757,N_28645);
and UO_235 (O_235,N_25784,N_26856);
xnor UO_236 (O_236,N_26296,N_27483);
and UO_237 (O_237,N_26979,N_25032);
and UO_238 (O_238,N_27165,N_29321);
nor UO_239 (O_239,N_29078,N_25130);
or UO_240 (O_240,N_25751,N_29327);
or UO_241 (O_241,N_26959,N_27882);
or UO_242 (O_242,N_29284,N_29923);
and UO_243 (O_243,N_29905,N_25513);
nand UO_244 (O_244,N_29353,N_25461);
and UO_245 (O_245,N_28606,N_26732);
xnor UO_246 (O_246,N_25986,N_26741);
xnor UO_247 (O_247,N_25842,N_26178);
or UO_248 (O_248,N_25793,N_26808);
nand UO_249 (O_249,N_26118,N_25099);
nor UO_250 (O_250,N_28144,N_29719);
or UO_251 (O_251,N_25800,N_28866);
or UO_252 (O_252,N_27224,N_26422);
and UO_253 (O_253,N_26325,N_29417);
or UO_254 (O_254,N_25983,N_26294);
nand UO_255 (O_255,N_29937,N_26497);
nand UO_256 (O_256,N_29175,N_26039);
or UO_257 (O_257,N_29449,N_26554);
and UO_258 (O_258,N_26924,N_27413);
nand UO_259 (O_259,N_28854,N_26306);
and UO_260 (O_260,N_25768,N_29845);
nand UO_261 (O_261,N_29004,N_29730);
and UO_262 (O_262,N_26080,N_26590);
xor UO_263 (O_263,N_28916,N_29394);
and UO_264 (O_264,N_27325,N_26196);
or UO_265 (O_265,N_25381,N_25216);
nor UO_266 (O_266,N_29855,N_29626);
nand UO_267 (O_267,N_26777,N_27026);
nor UO_268 (O_268,N_27513,N_27025);
or UO_269 (O_269,N_27910,N_27348);
nor UO_270 (O_270,N_27110,N_28969);
and UO_271 (O_271,N_28787,N_25836);
xnor UO_272 (O_272,N_26812,N_26693);
and UO_273 (O_273,N_27216,N_27378);
nand UO_274 (O_274,N_25370,N_27128);
and UO_275 (O_275,N_27727,N_25704);
and UO_276 (O_276,N_25815,N_29096);
xnor UO_277 (O_277,N_25989,N_27431);
nor UO_278 (O_278,N_28706,N_25489);
nor UO_279 (O_279,N_25672,N_26855);
or UO_280 (O_280,N_29980,N_25378);
xnor UO_281 (O_281,N_28709,N_29545);
or UO_282 (O_282,N_25354,N_29990);
xor UO_283 (O_283,N_25953,N_29461);
nor UO_284 (O_284,N_26869,N_27099);
or UO_285 (O_285,N_28886,N_26172);
nand UO_286 (O_286,N_27566,N_27037);
xnor UO_287 (O_287,N_25457,N_29961);
nor UO_288 (O_288,N_27811,N_27618);
or UO_289 (O_289,N_27181,N_25476);
or UO_290 (O_290,N_25116,N_28490);
and UO_291 (O_291,N_29373,N_27959);
nor UO_292 (O_292,N_27949,N_28051);
or UO_293 (O_293,N_28617,N_27208);
or UO_294 (O_294,N_28208,N_27676);
nand UO_295 (O_295,N_26379,N_26790);
xor UO_296 (O_296,N_28036,N_25288);
nand UO_297 (O_297,N_26207,N_29497);
xor UO_298 (O_298,N_27663,N_26920);
nand UO_299 (O_299,N_27312,N_27752);
nor UO_300 (O_300,N_29432,N_27804);
and UO_301 (O_301,N_25283,N_29352);
nor UO_302 (O_302,N_25560,N_29966);
nor UO_303 (O_303,N_28982,N_25211);
or UO_304 (O_304,N_27653,N_28147);
or UO_305 (O_305,N_28341,N_29777);
and UO_306 (O_306,N_27900,N_27386);
nand UO_307 (O_307,N_27845,N_28532);
and UO_308 (O_308,N_26961,N_28118);
and UO_309 (O_309,N_25572,N_25209);
and UO_310 (O_310,N_27805,N_27809);
or UO_311 (O_311,N_27829,N_29555);
or UO_312 (O_312,N_28375,N_28059);
nor UO_313 (O_313,N_27468,N_27062);
and UO_314 (O_314,N_28218,N_26005);
nor UO_315 (O_315,N_29648,N_26663);
and UO_316 (O_316,N_28684,N_26725);
or UO_317 (O_317,N_25104,N_25997);
nor UO_318 (O_318,N_25639,N_29487);
or UO_319 (O_319,N_25673,N_26007);
nor UO_320 (O_320,N_28360,N_29335);
nor UO_321 (O_321,N_26857,N_25826);
and UO_322 (O_322,N_26579,N_25500);
xnor UO_323 (O_323,N_29639,N_28785);
and UO_324 (O_324,N_27139,N_29883);
nor UO_325 (O_325,N_26671,N_26242);
or UO_326 (O_326,N_28226,N_27309);
nand UO_327 (O_327,N_26615,N_29364);
or UO_328 (O_328,N_28778,N_26830);
and UO_329 (O_329,N_28117,N_25357);
and UO_330 (O_330,N_26519,N_26136);
and UO_331 (O_331,N_28209,N_27240);
and UO_332 (O_332,N_27934,N_25979);
nor UO_333 (O_333,N_27365,N_27412);
xor UO_334 (O_334,N_27282,N_27958);
nor UO_335 (O_335,N_27610,N_25687);
nand UO_336 (O_336,N_28320,N_27646);
and UO_337 (O_337,N_25291,N_26434);
nor UO_338 (O_338,N_28447,N_28500);
nor UO_339 (O_339,N_27887,N_25011);
xor UO_340 (O_340,N_28640,N_28793);
nor UO_341 (O_341,N_26720,N_26394);
nor UO_342 (O_342,N_27124,N_28786);
nor UO_343 (O_343,N_28322,N_26106);
and UO_344 (O_344,N_27666,N_25064);
and UO_345 (O_345,N_25694,N_28242);
xor UO_346 (O_346,N_27700,N_29749);
and UO_347 (O_347,N_26610,N_29170);
nand UO_348 (O_348,N_26733,N_25214);
xor UO_349 (O_349,N_27710,N_28905);
nand UO_350 (O_350,N_29906,N_26753);
nor UO_351 (O_351,N_26146,N_28270);
or UO_352 (O_352,N_28013,N_29132);
nor UO_353 (O_353,N_26862,N_26776);
or UO_354 (O_354,N_26925,N_25615);
and UO_355 (O_355,N_25417,N_26240);
nand UO_356 (O_356,N_27350,N_28828);
nor UO_357 (O_357,N_26149,N_25156);
nor UO_358 (O_358,N_29584,N_29585);
and UO_359 (O_359,N_29772,N_25019);
and UO_360 (O_360,N_27654,N_26811);
nand UO_361 (O_361,N_25821,N_25552);
nor UO_362 (O_362,N_26927,N_27898);
nor UO_363 (O_363,N_28463,N_27641);
and UO_364 (O_364,N_25208,N_29600);
or UO_365 (O_365,N_25309,N_25232);
or UO_366 (O_366,N_27561,N_27488);
and UO_367 (O_367,N_27628,N_25189);
and UO_368 (O_368,N_28911,N_26697);
nor UO_369 (O_369,N_29862,N_29513);
nor UO_370 (O_370,N_28848,N_25846);
nor UO_371 (O_371,N_27631,N_27705);
and UO_372 (O_372,N_26631,N_29931);
nand UO_373 (O_373,N_28530,N_26886);
and UO_374 (O_374,N_25230,N_26922);
nand UO_375 (O_375,N_26594,N_25889);
nand UO_376 (O_376,N_27936,N_29799);
and UO_377 (O_377,N_26973,N_26164);
and UO_378 (O_378,N_28741,N_27106);
nor UO_379 (O_379,N_26455,N_29052);
nand UO_380 (O_380,N_26620,N_28460);
or UO_381 (O_381,N_28862,N_28523);
nand UO_382 (O_382,N_25990,N_25885);
or UO_383 (O_383,N_29059,N_25619);
or UO_384 (O_384,N_26834,N_29548);
and UO_385 (O_385,N_29149,N_29683);
or UO_386 (O_386,N_28580,N_29077);
nor UO_387 (O_387,N_27150,N_27347);
and UO_388 (O_388,N_25165,N_29693);
nor UO_389 (O_389,N_27020,N_26552);
and UO_390 (O_390,N_26227,N_25143);
nand UO_391 (O_391,N_25017,N_29938);
or UO_392 (O_392,N_29111,N_29612);
or UO_393 (O_393,N_29122,N_28374);
or UO_394 (O_394,N_25473,N_28003);
nand UO_395 (O_395,N_27090,N_29954);
nand UO_396 (O_396,N_25135,N_28723);
nand UO_397 (O_397,N_27272,N_25088);
nor UO_398 (O_398,N_26427,N_25851);
and UO_399 (O_399,N_26485,N_26395);
or UO_400 (O_400,N_27313,N_28967);
nor UO_401 (O_401,N_28995,N_25335);
or UO_402 (O_402,N_27180,N_28389);
and UO_403 (O_403,N_29695,N_27574);
and UO_404 (O_404,N_28116,N_29506);
xor UO_405 (O_405,N_25843,N_29710);
and UO_406 (O_406,N_28525,N_29745);
nor UO_407 (O_407,N_29851,N_29229);
or UO_408 (O_408,N_28577,N_25654);
nor UO_409 (O_409,N_25033,N_27985);
and UO_410 (O_410,N_28750,N_28289);
nor UO_411 (O_411,N_29301,N_28570);
and UO_412 (O_412,N_25495,N_28921);
nand UO_413 (O_413,N_29143,N_25423);
and UO_414 (O_414,N_28254,N_25002);
or UO_415 (O_415,N_28413,N_27823);
and UO_416 (O_416,N_29124,N_28975);
nor UO_417 (O_417,N_27731,N_25118);
nor UO_418 (O_418,N_25523,N_26050);
or UO_419 (O_419,N_29563,N_29503);
xnor UO_420 (O_420,N_27136,N_26751);
nor UO_421 (O_421,N_26915,N_25801);
nor UO_422 (O_422,N_26337,N_26402);
or UO_423 (O_423,N_28324,N_28426);
and UO_424 (O_424,N_28108,N_26185);
nand UO_425 (O_425,N_29088,N_28569);
nand UO_426 (O_426,N_25869,N_26425);
and UO_427 (O_427,N_25882,N_25025);
and UO_428 (O_428,N_28942,N_26458);
and UO_429 (O_429,N_27897,N_27399);
or UO_430 (O_430,N_25389,N_29817);
or UO_431 (O_431,N_25176,N_29521);
xnor UO_432 (O_432,N_25824,N_29160);
nor UO_433 (O_433,N_28694,N_25522);
and UO_434 (O_434,N_25710,N_28362);
nand UO_435 (O_435,N_26277,N_28291);
xnor UO_436 (O_436,N_27516,N_25566);
or UO_437 (O_437,N_27612,N_25621);
and UO_438 (O_438,N_27223,N_29462);
nand UO_439 (O_439,N_26357,N_27004);
nand UO_440 (O_440,N_28758,N_27761);
nand UO_441 (O_441,N_28112,N_29747);
xnor UO_442 (O_442,N_27844,N_25145);
or UO_443 (O_443,N_25172,N_26219);
nor UO_444 (O_444,N_27953,N_29559);
nor UO_445 (O_445,N_27598,N_27306);
xnor UO_446 (O_446,N_28336,N_26478);
nand UO_447 (O_447,N_25343,N_26318);
and UO_448 (O_448,N_29362,N_27824);
nand UO_449 (O_449,N_26873,N_25094);
and UO_450 (O_450,N_28598,N_27819);
and UO_451 (O_451,N_27304,N_25175);
nand UO_452 (O_452,N_28603,N_25597);
xor UO_453 (O_453,N_29330,N_27966);
and UO_454 (O_454,N_27450,N_26248);
nor UO_455 (O_455,N_28385,N_25907);
xnor UO_456 (O_456,N_27132,N_26246);
nand UO_457 (O_457,N_28166,N_29688);
nor UO_458 (O_458,N_26891,N_26089);
and UO_459 (O_459,N_28472,N_25379);
nor UO_460 (O_460,N_26452,N_25325);
nand UO_461 (O_461,N_26466,N_27127);
nor UO_462 (O_462,N_28417,N_27270);
nor UO_463 (O_463,N_26070,N_26987);
or UO_464 (O_464,N_25918,N_29075);
nor UO_465 (O_465,N_29231,N_29742);
nor UO_466 (O_466,N_25968,N_26532);
nor UO_467 (O_467,N_26426,N_26859);
nand UO_468 (O_468,N_29161,N_27538);
xnor UO_469 (O_469,N_27686,N_28178);
and UO_470 (O_470,N_28335,N_25556);
xnor UO_471 (O_471,N_26847,N_27153);
nand UO_472 (O_472,N_25747,N_28476);
xor UO_473 (O_473,N_27319,N_29744);
nor UO_474 (O_474,N_27963,N_25722);
nor UO_475 (O_475,N_28777,N_29890);
and UO_476 (O_476,N_26678,N_27524);
and UO_477 (O_477,N_27928,N_25777);
xor UO_478 (O_478,N_26344,N_26783);
xnor UO_479 (O_479,N_28827,N_26507);
xnor UO_480 (O_480,N_28581,N_27238);
nand UO_481 (O_481,N_28092,N_25403);
nor UO_482 (O_482,N_26769,N_25612);
or UO_483 (O_483,N_25823,N_26653);
nor UO_484 (O_484,N_28743,N_29617);
and UO_485 (O_485,N_26389,N_27905);
nand UO_486 (O_486,N_27696,N_28429);
and UO_487 (O_487,N_29977,N_28579);
xnor UO_488 (O_488,N_25630,N_28517);
nor UO_489 (O_489,N_29248,N_28847);
nor UO_490 (O_490,N_25251,N_26871);
nand UO_491 (O_491,N_27292,N_25284);
and UO_492 (O_492,N_29422,N_28479);
or UO_493 (O_493,N_29491,N_25206);
nand UO_494 (O_494,N_27460,N_26205);
or UO_495 (O_495,N_27065,N_27687);
and UO_496 (O_496,N_28977,N_27454);
nand UO_497 (O_497,N_27040,N_26929);
or UO_498 (O_498,N_27603,N_25420);
nand UO_499 (O_499,N_27404,N_27436);
nor UO_500 (O_500,N_29671,N_27358);
and UO_501 (O_501,N_28856,N_29934);
nor UO_502 (O_502,N_26075,N_26409);
or UO_503 (O_503,N_29466,N_27170);
or UO_504 (O_504,N_27457,N_29716);
and UO_505 (O_505,N_25038,N_28772);
nand UO_506 (O_506,N_25778,N_25540);
nor UO_507 (O_507,N_29125,N_25575);
or UO_508 (O_508,N_28363,N_28183);
or UO_509 (O_509,N_25089,N_28871);
nor UO_510 (O_510,N_26026,N_28831);
and UO_511 (O_511,N_27486,N_27342);
or UO_512 (O_512,N_27559,N_29519);
and UO_513 (O_513,N_28326,N_25355);
xor UO_514 (O_514,N_26461,N_26740);
or UO_515 (O_515,N_26696,N_26705);
or UO_516 (O_516,N_25530,N_27759);
nor UO_517 (O_517,N_27816,N_28194);
and UO_518 (O_518,N_25485,N_26030);
xnor UO_519 (O_519,N_29051,N_27742);
or UO_520 (O_520,N_26576,N_28237);
xnor UO_521 (O_521,N_25723,N_25949);
or UO_522 (O_522,N_29315,N_25746);
and UO_523 (O_523,N_29820,N_29272);
or UO_524 (O_524,N_27626,N_26451);
nand UO_525 (O_525,N_25563,N_26688);
nor UO_526 (O_526,N_26524,N_28295);
and UO_527 (O_527,N_25886,N_25396);
nor UO_528 (O_528,N_26268,N_29967);
and UO_529 (O_529,N_29041,N_26555);
and UO_530 (O_530,N_26717,N_26691);
or UO_531 (O_531,N_27881,N_28154);
and UO_532 (O_532,N_26934,N_26121);
xnor UO_533 (O_533,N_28210,N_27149);
nor UO_534 (O_534,N_26599,N_25961);
or UO_535 (O_535,N_29310,N_29543);
or UO_536 (O_536,N_25351,N_25787);
nor UO_537 (O_537,N_28497,N_28806);
and UO_538 (O_538,N_29164,N_27356);
nand UO_539 (O_539,N_25326,N_25876);
nand UO_540 (O_540,N_27504,N_29370);
nand UO_541 (O_541,N_26145,N_29642);
nand UO_542 (O_542,N_27033,N_26571);
and UO_543 (O_543,N_29540,N_29993);
nand UO_544 (O_544,N_26487,N_25439);
and UO_545 (O_545,N_28165,N_28011);
nor UO_546 (O_546,N_25731,N_29254);
or UO_547 (O_547,N_27672,N_29869);
or UO_548 (O_548,N_29006,N_26307);
or UO_549 (O_549,N_28711,N_25950);
xor UO_550 (O_550,N_28852,N_29674);
or UO_551 (O_551,N_27117,N_26974);
and UO_552 (O_552,N_25422,N_27539);
nor UO_553 (O_553,N_27931,N_29427);
nand UO_554 (O_554,N_28355,N_26743);
nor UO_555 (O_555,N_27496,N_28931);
and UO_556 (O_556,N_27455,N_26710);
nor UO_557 (O_557,N_26209,N_27915);
nor UO_558 (O_558,N_28686,N_25418);
and UO_559 (O_559,N_28093,N_25249);
xnor UO_560 (O_560,N_28358,N_27853);
or UO_561 (O_561,N_29685,N_29557);
nor UO_562 (O_562,N_29758,N_26980);
or UO_563 (O_563,N_26768,N_26596);
nand UO_564 (O_564,N_26370,N_25568);
nand UO_565 (O_565,N_25903,N_25034);
nor UO_566 (O_566,N_26286,N_25959);
and UO_567 (O_567,N_28173,N_27762);
nand UO_568 (O_568,N_29445,N_25974);
and UO_569 (O_569,N_29054,N_28064);
nand UO_570 (O_570,N_29805,N_27980);
nor UO_571 (O_571,N_29418,N_27779);
nand UO_572 (O_572,N_27073,N_26255);
nand UO_573 (O_573,N_27400,N_29770);
xor UO_574 (O_574,N_25912,N_27135);
nor UO_575 (O_575,N_28252,N_28557);
xor UO_576 (O_576,N_26109,N_26645);
and UO_577 (O_577,N_29733,N_27109);
nor UO_578 (O_578,N_26622,N_26606);
and UO_579 (O_579,N_28666,N_27063);
nor UO_580 (O_580,N_26535,N_28042);
and UO_581 (O_581,N_29238,N_25977);
xnor UO_582 (O_582,N_29239,N_29286);
and UO_583 (O_583,N_29121,N_26082);
xor UO_584 (O_584,N_28232,N_26529);
xor UO_585 (O_585,N_27331,N_26809);
and UO_586 (O_586,N_25074,N_26708);
and UO_587 (O_587,N_27981,N_26004);
or UO_588 (O_588,N_29233,N_28283);
and UO_589 (O_589,N_26295,N_26982);
xor UO_590 (O_590,N_27706,N_27537);
nor UO_591 (O_591,N_28807,N_25286);
and UO_592 (O_592,N_27973,N_26659);
xnor UO_593 (O_593,N_27254,N_27586);
or UO_594 (O_594,N_27024,N_27755);
and UO_595 (O_595,N_28167,N_26481);
nor UO_596 (O_596,N_25030,N_29388);
nor UO_597 (O_597,N_26706,N_28502);
or UO_598 (O_598,N_28213,N_25678);
nor UO_599 (O_599,N_29459,N_27166);
nand UO_600 (O_600,N_28771,N_27408);
nand UO_601 (O_601,N_26851,N_29854);
xnor UO_602 (O_602,N_26612,N_26025);
nor UO_603 (O_603,N_28765,N_25365);
nor UO_604 (O_604,N_25260,N_26386);
or UO_605 (O_605,N_27148,N_28103);
or UO_606 (O_606,N_29099,N_25186);
and UO_607 (O_607,N_27723,N_27968);
xor UO_608 (O_608,N_25559,N_27810);
and UO_609 (O_609,N_28822,N_27802);
or UO_610 (O_610,N_29050,N_27917);
or UO_611 (O_611,N_28373,N_27536);
and UO_612 (O_612,N_27930,N_28306);
xnor UO_613 (O_613,N_25919,N_29920);
or UO_614 (O_614,N_26304,N_26157);
xor UO_615 (O_615,N_29909,N_25137);
or UO_616 (O_616,N_28230,N_26884);
xor UO_617 (O_617,N_28409,N_25608);
nor UO_618 (O_618,N_29475,N_26220);
and UO_619 (O_619,N_29203,N_25506);
and UO_620 (O_620,N_26562,N_25460);
nand UO_621 (O_621,N_27470,N_29780);
nand UO_622 (O_622,N_29408,N_28996);
nand UO_623 (O_623,N_25761,N_28372);
xnor UO_624 (O_624,N_26411,N_25624);
and UO_625 (O_625,N_27550,N_29661);
nand UO_626 (O_626,N_26058,N_28663);
nor UO_627 (O_627,N_27577,N_25883);
and UO_628 (O_628,N_25707,N_25194);
or UO_629 (O_629,N_29480,N_26954);
and UO_630 (O_630,N_26644,N_29180);
nor UO_631 (O_631,N_28730,N_26966);
nor UO_632 (O_632,N_25109,N_25072);
or UO_633 (O_633,N_29289,N_29981);
nor UO_634 (O_634,N_25850,N_25134);
xnor UO_635 (O_635,N_27952,N_26053);
nor UO_636 (O_636,N_25036,N_27572);
nor UO_637 (O_637,N_25078,N_25190);
and UO_638 (O_638,N_27322,N_28313);
nand UO_639 (O_639,N_25113,N_28553);
and UO_640 (O_640,N_25705,N_25647);
or UO_641 (O_641,N_28899,N_27716);
nand UO_642 (O_642,N_26619,N_26234);
and UO_643 (O_643,N_28721,N_28698);
xnor UO_644 (O_644,N_28707,N_29965);
or UO_645 (O_645,N_25219,N_27321);
nor UO_646 (O_646,N_26204,N_25939);
nor UO_647 (O_647,N_27689,N_27820);
and UO_648 (O_648,N_28587,N_27777);
nand UO_649 (O_649,N_25312,N_29720);
nor UO_650 (O_650,N_29490,N_27440);
or UO_651 (O_651,N_28634,N_29308);
nand UO_652 (O_652,N_28691,N_28094);
nand UO_653 (O_653,N_28334,N_29429);
or UO_654 (O_654,N_28519,N_27114);
nor UO_655 (O_655,N_29984,N_27748);
nor UO_656 (O_656,N_26372,N_28293);
nor UO_657 (O_657,N_27226,N_27487);
or UO_658 (O_658,N_29551,N_25490);
xnor UO_659 (O_659,N_25487,N_26291);
nand UO_660 (O_660,N_26197,N_28498);
and UO_661 (O_661,N_25383,N_27749);
and UO_662 (O_662,N_26918,N_27637);
or UO_663 (O_663,N_25945,N_28797);
and UO_664 (O_664,N_28823,N_27058);
nand UO_665 (O_665,N_26187,N_27042);
nor UO_666 (O_666,N_26336,N_25154);
nand UO_667 (O_667,N_28153,N_28015);
nor UO_668 (O_668,N_29204,N_29236);
and UO_669 (O_669,N_29783,N_29723);
and UO_670 (O_670,N_28623,N_27737);
nor UO_671 (O_671,N_26382,N_27017);
and UO_672 (O_672,N_29241,N_29628);
nand UO_673 (O_673,N_26780,N_29645);
and UO_674 (O_674,N_25465,N_28941);
nand UO_675 (O_675,N_28782,N_29998);
nand UO_676 (O_676,N_27071,N_27634);
and UO_677 (O_677,N_28290,N_29263);
nand UO_678 (O_678,N_28953,N_29499);
or UO_679 (O_679,N_26711,N_28440);
nand UO_680 (O_680,N_25107,N_28382);
nor UO_681 (O_681,N_25660,N_27508);
nand UO_682 (O_682,N_27474,N_27699);
nand UO_683 (O_683,N_28225,N_29354);
and UO_684 (O_684,N_27549,N_29815);
nor UO_685 (O_685,N_25636,N_29995);
nor UO_686 (O_686,N_29971,N_25491);
nand UO_687 (O_687,N_27528,N_26243);
or UO_688 (O_688,N_29220,N_29831);
nor UO_689 (O_689,N_26200,N_29502);
and UO_690 (O_690,N_28631,N_29186);
nand UO_691 (O_691,N_26290,N_27246);
and UO_692 (O_692,N_26516,N_29609);
nor UO_693 (O_693,N_25543,N_27253);
nor UO_694 (O_694,N_26745,N_29514);
or UO_695 (O_695,N_27660,N_28713);
nand UO_696 (O_696,N_27357,N_25991);
or UO_697 (O_697,N_28273,N_25643);
xnor UO_698 (O_698,N_27172,N_25481);
nor UO_699 (O_699,N_25185,N_25159);
and UO_700 (O_700,N_26935,N_25066);
nand UO_701 (O_701,N_25947,N_26015);
or UO_702 (O_702,N_28444,N_27808);
and UO_703 (O_703,N_28281,N_27826);
nand UO_704 (O_704,N_26747,N_28976);
or UO_705 (O_705,N_27395,N_25571);
and UO_706 (O_706,N_25467,N_28067);
and UO_707 (O_707,N_29318,N_26940);
nand UO_708 (O_708,N_27590,N_28764);
xnor UO_709 (O_709,N_25517,N_25114);
nand UO_710 (O_710,N_28927,N_26623);
nand UO_711 (O_711,N_29761,N_28125);
nor UO_712 (O_712,N_25141,N_27387);
nand UO_713 (O_713,N_29667,N_28729);
nor UO_714 (O_714,N_29822,N_29795);
nand UO_715 (O_715,N_25229,N_27923);
nand UO_716 (O_716,N_27522,N_27924);
xnor UO_717 (O_717,N_29014,N_28469);
and UO_718 (O_718,N_25241,N_27996);
or UO_719 (O_719,N_28151,N_26317);
nand UO_720 (O_720,N_28867,N_25521);
or UO_721 (O_721,N_25537,N_25345);
nand UO_722 (O_722,N_25202,N_28308);
xnor UO_723 (O_723,N_26953,N_25737);
or UO_724 (O_724,N_25254,N_25394);
xnor UO_725 (O_725,N_28041,N_26091);
nand UO_726 (O_726,N_26804,N_29871);
nand UO_727 (O_727,N_25661,N_25564);
and UO_728 (O_728,N_27220,N_28675);
nor UO_729 (O_729,N_27690,N_27841);
or UO_730 (O_730,N_29640,N_25925);
or UO_731 (O_731,N_25541,N_27526);
nor UO_732 (O_732,N_26995,N_28288);
nor UO_733 (O_733,N_25498,N_29718);
or UO_734 (O_734,N_28102,N_27568);
or UO_735 (O_735,N_26273,N_29930);
or UO_736 (O_736,N_28404,N_26607);
or UO_737 (O_737,N_26947,N_28485);
or UO_738 (O_738,N_28520,N_25507);
or UO_739 (O_739,N_25398,N_25943);
or UO_740 (O_740,N_25730,N_25584);
or UO_741 (O_741,N_28536,N_29409);
nand UO_742 (O_742,N_29228,N_26244);
nand UO_743 (O_743,N_25097,N_27894);
xnor UO_744 (O_744,N_29214,N_29598);
or UO_745 (O_745,N_28875,N_29305);
or UO_746 (O_746,N_29996,N_27416);
nor UO_747 (O_747,N_26192,N_29881);
xor UO_748 (O_748,N_29493,N_28395);
nor UO_749 (O_749,N_28186,N_27776);
nand UO_750 (O_750,N_26700,N_29530);
nor UO_751 (O_751,N_26759,N_29196);
nand UO_752 (O_752,N_25256,N_29147);
xor UO_753 (O_753,N_29107,N_29168);
nor UO_754 (O_754,N_26604,N_28647);
and UO_755 (O_755,N_26329,N_26721);
nor UO_756 (O_756,N_27567,N_25780);
nand UO_757 (O_757,N_26799,N_25369);
and UO_758 (O_758,N_26313,N_27376);
or UO_759 (O_759,N_27167,N_25428);
or UO_760 (O_760,N_26400,N_29888);
and UO_761 (O_761,N_28541,N_26449);
and UO_762 (O_762,N_25588,N_26945);
or UO_763 (O_763,N_26609,N_28834);
and UO_764 (O_764,N_29827,N_26056);
and UO_765 (O_765,N_25071,N_29884);
nand UO_766 (O_766,N_25277,N_27695);
or UO_767 (O_767,N_27195,N_28217);
nor UO_768 (O_768,N_26880,N_29686);
nor UO_769 (O_769,N_28518,N_28275);
nor UO_770 (O_770,N_29668,N_27979);
nor UO_771 (O_771,N_26616,N_28206);
nor UO_772 (O_772,N_28265,N_29529);
and UO_773 (O_773,N_28279,N_29198);
and UO_774 (O_774,N_28903,N_28136);
and UO_775 (O_775,N_27129,N_28643);
xnor UO_776 (O_776,N_25740,N_27842);
nor UO_777 (O_777,N_27323,N_27381);
and UO_778 (O_778,N_25429,N_26713);
xor UO_779 (O_779,N_27977,N_28515);
or UO_780 (O_780,N_27284,N_25999);
xor UO_781 (O_781,N_25356,N_26168);
and UO_782 (O_782,N_29887,N_27532);
or UO_783 (O_783,N_27974,N_26116);
nand UO_784 (O_784,N_27175,N_26177);
and UO_785 (O_785,N_26009,N_29837);
and UO_786 (O_786,N_25318,N_28593);
xor UO_787 (O_787,N_28138,N_25954);
or UO_788 (O_788,N_28700,N_26573);
and UO_789 (O_789,N_29376,N_25839);
or UO_790 (O_790,N_26237,N_27187);
nor UO_791 (O_791,N_28082,N_29646);
nor UO_792 (O_792,N_29601,N_25781);
and UO_793 (O_793,N_27384,N_28432);
or UO_794 (O_794,N_27875,N_26174);
xnor UO_795 (O_795,N_28115,N_27661);
and UO_796 (O_796,N_27280,N_27836);
nor UO_797 (O_797,N_26642,N_25258);
and UO_798 (O_798,N_26755,N_27008);
or UO_799 (O_799,N_29794,N_29118);
xor UO_800 (O_800,N_28900,N_29800);
or UO_801 (O_801,N_29986,N_28346);
xor UO_802 (O_802,N_29932,N_25063);
or UO_803 (O_803,N_27047,N_27530);
nand UO_804 (O_804,N_26952,N_28303);
and UO_805 (O_805,N_25806,N_27607);
xor UO_806 (O_806,N_26546,N_25577);
nor UO_807 (O_807,N_29424,N_26170);
and UO_808 (O_808,N_26669,N_27461);
and UO_809 (O_809,N_28913,N_29634);
xnor UO_810 (O_810,N_26289,N_28100);
and UO_811 (O_811,N_25609,N_25294);
nand UO_812 (O_812,N_25544,N_29902);
or UO_813 (O_813,N_26198,N_29828);
and UO_814 (O_814,N_25993,N_27390);
nor UO_815 (O_815,N_29049,N_29391);
xor UO_816 (O_816,N_25331,N_28205);
or UO_817 (O_817,N_25077,N_26660);
nand UO_818 (O_818,N_27159,N_27074);
nor UO_819 (O_819,N_26499,N_25735);
nand UO_820 (O_820,N_28892,N_26840);
and UO_821 (O_821,N_26061,N_25679);
or UO_822 (O_822,N_25065,N_26371);
xnor UO_823 (O_823,N_28076,N_26051);
and UO_824 (O_824,N_25070,N_28537);
and UO_825 (O_825,N_28412,N_28269);
and UO_826 (O_826,N_29128,N_28539);
xor UO_827 (O_827,N_25948,N_25204);
nand UO_828 (O_828,N_25453,N_29153);
and UO_829 (O_829,N_28547,N_27828);
or UO_830 (O_830,N_29064,N_28597);
nand UO_831 (O_831,N_26262,N_25819);
nor UO_832 (O_832,N_28376,N_27523);
nor UO_833 (O_833,N_27950,N_29978);
xnor UO_834 (O_834,N_26828,N_25718);
nor UO_835 (O_835,N_26685,N_28555);
and UO_836 (O_836,N_27833,N_25007);
and UO_837 (O_837,N_29830,N_29941);
nand UO_838 (O_838,N_26494,N_26677);
and UO_839 (O_839,N_26763,N_26437);
and UO_840 (O_840,N_28920,N_26133);
nor UO_841 (O_841,N_25814,N_28347);
nor UO_842 (O_842,N_29191,N_29086);
and UO_843 (O_843,N_29568,N_29460);
nor UO_844 (O_844,N_29250,N_27888);
xnor UO_845 (O_845,N_25265,N_28908);
or UO_846 (O_846,N_28737,N_28020);
nand UO_847 (O_847,N_26377,N_28001);
and UO_848 (O_848,N_28380,N_27424);
and UO_849 (O_849,N_28792,N_27271);
nor UO_850 (O_850,N_27497,N_27101);
or UO_851 (O_851,N_26699,N_29398);
nand UO_852 (O_852,N_29065,N_26122);
and UO_853 (O_853,N_25187,N_27863);
nand UO_854 (O_854,N_26716,N_26293);
and UO_855 (O_855,N_28654,N_29033);
or UO_856 (O_856,N_25095,N_25978);
or UO_857 (O_857,N_27298,N_27382);
or UO_858 (O_858,N_26128,N_28396);
xnor UO_859 (O_859,N_25922,N_29801);
nor UO_860 (O_860,N_25173,N_28323);
and UO_861 (O_861,N_29637,N_27638);
nor UO_862 (O_862,N_26701,N_29043);
nand UO_863 (O_863,N_27883,N_28228);
nand UO_864 (O_864,N_25518,N_28491);
nand UO_865 (O_865,N_29561,N_26328);
nor UO_866 (O_866,N_25802,N_26649);
or UO_867 (O_867,N_26635,N_28988);
and UO_868 (O_868,N_25503,N_26592);
and UO_869 (O_869,N_29397,N_29769);
or UO_870 (O_870,N_25702,N_25246);
nor UO_871 (O_871,N_28247,N_25927);
nor UO_872 (O_872,N_29242,N_26100);
or UO_873 (O_873,N_26983,N_28489);
nor UO_874 (O_874,N_29265,N_29292);
nor UO_875 (O_875,N_28177,N_27344);
xor UO_876 (O_876,N_26698,N_29199);
nor UO_877 (O_877,N_25611,N_28240);
or UO_878 (O_878,N_27565,N_28098);
nand UO_879 (O_879,N_29946,N_28919);
and UO_880 (O_880,N_29798,N_25844);
and UO_881 (O_881,N_26636,N_27275);
or UO_882 (O_882,N_27250,N_28620);
xnor UO_883 (O_883,N_27283,N_25380);
nor UO_884 (O_884,N_28804,N_27294);
nand UO_885 (O_885,N_25759,N_29456);
nand UO_886 (O_886,N_26190,N_27182);
nand UO_887 (O_887,N_27632,N_25874);
and UO_888 (O_888,N_27780,N_29380);
or UO_889 (O_889,N_25400,N_29899);
nand UO_890 (O_890,N_27116,N_28763);
and UO_891 (O_891,N_27263,N_29055);
and UO_892 (O_892,N_27362,N_28602);
or UO_893 (O_893,N_26789,N_25942);
nor UO_894 (O_894,N_27617,N_28954);
nand UO_895 (O_895,N_27946,N_25626);
nor UO_896 (O_896,N_26393,N_25152);
nor UO_897 (O_897,N_27693,N_26201);
xor UO_898 (O_898,N_27769,N_26991);
nand UO_899 (O_899,N_29877,N_27499);
or UO_900 (O_900,N_26715,N_28633);
or UO_901 (O_901,N_29656,N_25402);
nor UO_902 (O_902,N_29829,N_28761);
and UO_903 (O_903,N_27589,N_29579);
nor UO_904 (O_904,N_28464,N_28345);
nand UO_905 (O_905,N_29870,N_29243);
and UO_906 (O_906,N_27683,N_26767);
and UO_907 (O_907,N_28985,N_25281);
nand UO_908 (O_908,N_27089,N_27052);
and UO_909 (O_909,N_28239,N_27884);
nor UO_910 (O_910,N_29784,N_29401);
nand UO_911 (O_911,N_26251,N_25340);
and UO_912 (O_912,N_25946,N_29615);
or UO_913 (O_913,N_28524,N_25832);
or UO_914 (O_914,N_28402,N_28738);
nand UO_915 (O_915,N_26105,N_27743);
or UO_916 (O_916,N_25813,N_29093);
and UO_917 (O_917,N_27753,N_26749);
and UO_918 (O_918,N_26526,N_29176);
nand UO_919 (O_919,N_29788,N_27484);
xnor UO_920 (O_920,N_29603,N_26078);
and UO_921 (O_921,N_28058,N_25098);
nand UO_922 (O_922,N_27485,N_28493);
xnor UO_923 (O_923,N_25600,N_27430);
and UO_924 (O_924,N_26326,N_26936);
nand UO_925 (O_925,N_25785,N_28435);
xor UO_926 (O_926,N_27503,N_25364);
nand UO_927 (O_927,N_28853,N_26028);
and UO_928 (O_928,N_25962,N_29202);
xnor UO_929 (O_929,N_25822,N_28486);
nand UO_930 (O_930,N_28251,N_26221);
and UO_931 (O_931,N_29206,N_28180);
or UO_932 (O_932,N_28215,N_29636);
and UO_933 (O_933,N_28826,N_29737);
nor UO_934 (O_934,N_26218,N_28458);
or UO_935 (O_935,N_26731,N_25681);
or UO_936 (O_936,N_26911,N_28732);
xor UO_937 (O_937,N_26771,N_27794);
nand UO_938 (O_938,N_25274,N_25696);
nor UO_939 (O_939,N_26147,N_29910);
nor UO_940 (O_940,N_25057,N_26226);
nor UO_941 (O_941,N_27976,N_27498);
and UO_942 (O_942,N_28531,N_25914);
or UO_943 (O_943,N_29314,N_28095);
and UO_944 (O_944,N_27456,N_25455);
nand UO_945 (O_945,N_27016,N_25080);
and UO_946 (O_946,N_25653,N_29874);
nand UO_947 (O_947,N_28526,N_25791);
xnor UO_948 (O_948,N_28388,N_25697);
and UO_949 (O_949,N_26539,N_25101);
xnor UO_950 (O_950,N_25595,N_29812);
xor UO_951 (O_951,N_29619,N_28113);
or UO_952 (O_952,N_25805,N_29415);
or UO_953 (O_953,N_28987,N_27103);
nand UO_954 (O_954,N_25085,N_29484);
and UO_955 (O_955,N_26259,N_29325);
xnor UO_956 (O_956,N_28424,N_25458);
xnor UO_957 (O_957,N_25073,N_29926);
and UO_958 (O_958,N_25424,N_28337);
nor UO_959 (O_959,N_29246,N_27087);
nand UO_960 (O_960,N_28972,N_27865);
or UO_961 (O_961,N_29097,N_28668);
xor UO_962 (O_962,N_25492,N_28211);
or UO_963 (O_963,N_25745,N_26868);
nor UO_964 (O_964,N_26239,N_25632);
nand UO_965 (O_965,N_27396,N_25726);
and UO_966 (O_966,N_29446,N_25031);
xor UO_967 (O_967,N_27551,N_26254);
nor UO_968 (O_968,N_25384,N_29684);
nand UO_969 (O_969,N_29017,N_29472);
or UO_970 (O_970,N_28249,N_29280);
xnor UO_971 (O_971,N_26544,N_26495);
nor UO_972 (O_972,N_27904,N_29546);
xnor UO_973 (O_973,N_28175,N_27411);
nor UO_974 (O_974,N_25640,N_26964);
and UO_975 (O_975,N_27726,N_29044);
xnor UO_976 (O_976,N_26568,N_26186);
nor UO_977 (O_977,N_28650,N_25628);
nand UO_978 (O_978,N_27009,N_29825);
nand UO_979 (O_979,N_29439,N_28683);
or UO_980 (O_980,N_26189,N_27364);
and UO_981 (O_981,N_28231,N_29056);
nand UO_982 (O_982,N_25125,N_27285);
nor UO_983 (O_983,N_25561,N_27256);
nand UO_984 (O_984,N_25535,N_28068);
nor UO_985 (O_985,N_28073,N_28263);
or UO_986 (O_986,N_25111,N_26852);
and UO_987 (O_987,N_28740,N_28410);
xor UO_988 (O_988,N_25385,N_25050);
xor UO_989 (O_989,N_29095,N_27786);
nor UO_990 (O_990,N_26558,N_28079);
nor UO_991 (O_991,N_25395,N_27629);
or UO_992 (O_992,N_29230,N_25671);
nor UO_993 (O_993,N_27458,N_26598);
nor UO_994 (O_994,N_27453,N_27010);
nand UO_995 (O_995,N_29721,N_28708);
or UO_996 (O_996,N_28105,N_28227);
nor UO_997 (O_997,N_26284,N_29633);
or UO_998 (O_998,N_29988,N_26823);
and UO_999 (O_999,N_25505,N_26309);
nor UO_1000 (O_1000,N_25715,N_27709);
nor UO_1001 (O_1001,N_26893,N_26013);
or UO_1002 (O_1002,N_27048,N_27377);
xor UO_1003 (O_1003,N_26960,N_27942);
and UO_1004 (O_1004,N_26119,N_28089);
and UO_1005 (O_1005,N_28679,N_28829);
and UO_1006 (O_1006,N_27850,N_27156);
or UO_1007 (O_1007,N_25086,N_28607);
nand UO_1008 (O_1008,N_25957,N_25684);
and UO_1009 (O_1009,N_25913,N_28596);
nand UO_1010 (O_1010,N_27595,N_29922);
nor UO_1011 (O_1011,N_28588,N_29858);
nor UO_1012 (O_1012,N_29483,N_27462);
or UO_1013 (O_1013,N_27351,N_29127);
nand UO_1014 (O_1014,N_26090,N_26602);
and UO_1015 (O_1015,N_28075,N_29550);
or UO_1016 (O_1016,N_27901,N_29620);
and UO_1017 (O_1017,N_29085,N_28294);
nor UO_1018 (O_1018,N_27383,N_28034);
and UO_1019 (O_1019,N_26890,N_26042);
nor UO_1020 (O_1020,N_29046,N_26514);
nand UO_1021 (O_1021,N_25853,N_27770);
nor UO_1022 (O_1022,N_29057,N_28870);
and UO_1023 (O_1023,N_29167,N_25923);
or UO_1024 (O_1024,N_25203,N_26842);
nor UO_1025 (O_1025,N_29400,N_26420);
nand UO_1026 (O_1026,N_29255,N_27422);
nor UO_1027 (O_1027,N_26531,N_27121);
nand UO_1028 (O_1028,N_25686,N_26846);
or UO_1029 (O_1029,N_29569,N_26683);
nor UO_1030 (O_1030,N_27838,N_27854);
or UO_1031 (O_1031,N_25084,N_29714);
nor UO_1032 (O_1032,N_29538,N_25878);
and UO_1033 (O_1033,N_25218,N_29312);
and UO_1034 (O_1034,N_25404,N_29525);
nor UO_1035 (O_1035,N_28902,N_29539);
and UO_1036 (O_1036,N_25479,N_26876);
or UO_1037 (O_1037,N_28297,N_25606);
or UO_1038 (O_1038,N_27621,N_26719);
and UO_1039 (O_1039,N_26384,N_27839);
nand UO_1040 (O_1040,N_29413,N_25858);
and UO_1041 (O_1041,N_29614,N_26057);
nand UO_1042 (O_1042,N_29687,N_29578);
nor UO_1043 (O_1043,N_29793,N_25788);
nor UO_1044 (O_1044,N_28818,N_29337);
or UO_1045 (O_1045,N_28392,N_25469);
nand UO_1046 (O_1046,N_29372,N_28885);
and UO_1047 (O_1047,N_25900,N_28563);
and UO_1048 (O_1048,N_27051,N_27619);
xnor UO_1049 (O_1049,N_26534,N_25426);
and UO_1050 (O_1050,N_27162,N_27472);
nor UO_1051 (O_1051,N_25023,N_27092);
or UO_1052 (O_1052,N_26073,N_28897);
and UO_1053 (O_1053,N_28503,N_28416);
nor UO_1054 (O_1054,N_29339,N_29913);
and UO_1055 (O_1055,N_26132,N_28329);
or UO_1056 (O_1056,N_26498,N_26572);
nor UO_1057 (O_1057,N_27418,N_26125);
nand UO_1058 (O_1058,N_25590,N_28863);
nand UO_1059 (O_1059,N_28378,N_26899);
xor UO_1060 (O_1060,N_25005,N_27225);
nor UO_1061 (O_1061,N_29297,N_27788);
and UO_1062 (O_1062,N_27799,N_26391);
nor UO_1063 (O_1063,N_29806,N_25502);
nor UO_1064 (O_1064,N_25693,N_25382);
xor UO_1065 (O_1065,N_25046,N_26718);
and UO_1066 (O_1066,N_28722,N_29701);
and UO_1067 (O_1067,N_28280,N_26457);
nor UO_1068 (O_1068,N_29712,N_25982);
and UO_1069 (O_1069,N_26484,N_27257);
or UO_1070 (O_1070,N_29537,N_28745);
and UO_1071 (O_1071,N_27057,N_26275);
nor UO_1072 (O_1072,N_29306,N_29564);
or UO_1073 (O_1073,N_28459,N_28010);
and UO_1074 (O_1074,N_26756,N_26071);
nand UO_1075 (O_1075,N_29189,N_25237);
xor UO_1076 (O_1076,N_28993,N_29218);
xnor UO_1077 (O_1077,N_25150,N_28312);
nor UO_1078 (O_1078,N_25191,N_29864);
nand UO_1079 (O_1079,N_29916,N_26858);
xnor UO_1080 (O_1080,N_28795,N_29650);
nand UO_1081 (O_1081,N_25322,N_26292);
nand UO_1082 (O_1082,N_28033,N_28947);
nand UO_1083 (O_1083,N_27995,N_28087);
nand UO_1084 (O_1084,N_29606,N_28934);
nand UO_1085 (O_1085,N_28933,N_25551);
or UO_1086 (O_1086,N_28928,N_28612);
nand UO_1087 (O_1087,N_25725,N_26195);
xor UO_1088 (O_1088,N_29673,N_28817);
nor UO_1089 (O_1089,N_27147,N_25896);
xor UO_1090 (O_1090,N_27415,N_28540);
nor UO_1091 (O_1091,N_27948,N_27721);
and UO_1092 (O_1092,N_25388,N_26651);
nand UO_1093 (O_1093,N_28552,N_27429);
and UO_1094 (O_1094,N_27951,N_27987);
nand UO_1095 (O_1095,N_28528,N_25406);
nor UO_1096 (O_1096,N_29754,N_27064);
nand UO_1097 (O_1097,N_26263,N_27956);
and UO_1098 (O_1098,N_29508,N_28803);
or UO_1099 (O_1099,N_29347,N_25808);
and UO_1100 (O_1100,N_28600,N_28929);
nor UO_1101 (O_1101,N_27494,N_28150);
or UO_1102 (O_1102,N_26120,N_28197);
nand UO_1103 (O_1103,N_28739,N_29903);
and UO_1104 (O_1104,N_26008,N_25692);
and UO_1105 (O_1105,N_26739,N_27702);
and UO_1106 (O_1106,N_28122,N_29245);
nand UO_1107 (O_1107,N_28534,N_25799);
and UO_1108 (O_1108,N_29477,N_28635);
or UO_1109 (O_1109,N_28594,N_25767);
or UO_1110 (O_1110,N_26224,N_29129);
and UO_1111 (O_1111,N_26737,N_26955);
nor UO_1112 (O_1112,N_28276,N_29058);
nand UO_1113 (O_1113,N_28879,N_27426);
xnor UO_1114 (O_1114,N_28506,N_26646);
and UO_1115 (O_1115,N_28789,N_28258);
and UO_1116 (O_1116,N_29139,N_28005);
and UO_1117 (O_1117,N_28644,N_29252);
or UO_1118 (O_1118,N_28146,N_28671);
and UO_1119 (O_1119,N_29501,N_28414);
or UO_1120 (O_1120,N_27370,N_26228);
nor UO_1121 (O_1121,N_25106,N_29317);
or UO_1122 (O_1122,N_29283,N_25511);
and UO_1123 (O_1123,N_28484,N_25712);
or UO_1124 (O_1124,N_28751,N_28483);
nor UO_1125 (O_1125,N_28452,N_26766);
xnor UO_1126 (O_1126,N_28695,N_29062);
xor UO_1127 (O_1127,N_25742,N_27625);
nand UO_1128 (O_1128,N_27338,N_26587);
or UO_1129 (O_1129,N_29891,N_28674);
xor UO_1130 (O_1130,N_26002,N_27678);
xnor UO_1131 (O_1131,N_25862,N_28843);
xor UO_1132 (O_1132,N_27814,N_25574);
or UO_1133 (O_1133,N_29404,N_28422);
nor UO_1134 (O_1134,N_26044,N_29430);
nand UO_1135 (O_1135,N_27477,N_26114);
or UO_1136 (O_1136,N_26506,N_26904);
nor UO_1137 (O_1137,N_29809,N_25764);
and UO_1138 (O_1138,N_28687,N_27903);
nand UO_1139 (O_1139,N_25477,N_25213);
nor UO_1140 (O_1140,N_28825,N_29717);
or UO_1141 (O_1141,N_25377,N_29028);
or UO_1142 (O_1142,N_26488,N_26764);
nand UO_1143 (O_1143,N_28788,N_29949);
and UO_1144 (O_1144,N_27929,N_26314);
nand UO_1145 (O_1145,N_25482,N_29541);
or UO_1146 (O_1146,N_27978,N_29092);
or UO_1147 (O_1147,N_27708,N_26250);
nand UO_1148 (O_1148,N_25634,N_28548);
nor UO_1149 (O_1149,N_29102,N_28262);
nand UO_1150 (O_1150,N_26113,N_29678);
or UO_1151 (O_1151,N_28069,N_26041);
xor UO_1152 (O_1152,N_27091,N_28244);
and UO_1153 (O_1153,N_28669,N_26639);
nand UO_1154 (O_1154,N_25315,N_26650);
nor UO_1155 (O_1155,N_27084,N_25934);
nand UO_1156 (O_1156,N_29414,N_28924);
nand UO_1157 (O_1157,N_25685,N_27738);
or UO_1158 (O_1158,N_26154,N_28813);
xor UO_1159 (O_1159,N_25917,N_26447);
and UO_1160 (O_1160,N_25549,N_27314);
or UO_1161 (O_1161,N_26236,N_29833);
nand UO_1162 (O_1162,N_26167,N_25818);
nor UO_1163 (O_1163,N_27855,N_25020);
nand UO_1164 (O_1164,N_29156,N_26536);
nor UO_1165 (O_1165,N_26887,N_26978);
or UO_1166 (O_1166,N_27300,N_26474);
or UO_1167 (O_1167,N_29104,N_29379);
xor UO_1168 (O_1168,N_25153,N_25614);
nand UO_1169 (O_1169,N_27902,N_26340);
nor UO_1170 (O_1170,N_28614,N_28351);
and UO_1171 (O_1171,N_28344,N_25303);
and UO_1172 (O_1172,N_29677,N_28796);
xnor UO_1173 (O_1173,N_27891,N_25397);
xor UO_1174 (O_1174,N_29141,N_26522);
and UO_1175 (O_1175,N_25527,N_27862);
or UO_1176 (O_1176,N_27308,N_26016);
nand UO_1177 (O_1177,N_28833,N_27160);
or UO_1178 (O_1178,N_25236,N_28282);
xor UO_1179 (O_1179,N_28043,N_25803);
nand UO_1180 (O_1180,N_27465,N_26440);
or UO_1181 (O_1181,N_26996,N_25859);
nor UO_1182 (O_1182,N_28835,N_26023);
or UO_1183 (O_1183,N_28492,N_27579);
nand UO_1184 (O_1184,N_28961,N_26266);
xnor UO_1185 (O_1185,N_27251,N_29098);
or UO_1186 (O_1186,N_27501,N_27452);
and UO_1187 (O_1187,N_28880,N_28584);
and UO_1188 (O_1188,N_28384,N_27143);
and UO_1189 (O_1189,N_27449,N_25361);
and UO_1190 (O_1190,N_27448,N_27707);
nor UO_1191 (O_1191,N_28292,N_28488);
nand UO_1192 (O_1192,N_25804,N_28907);
nand UO_1193 (O_1193,N_29219,N_27796);
and UO_1194 (O_1194,N_26993,N_26140);
or UO_1195 (O_1195,N_27330,N_28990);
or UO_1196 (O_1196,N_26282,N_26655);
xor UO_1197 (O_1197,N_25167,N_29835);
nand UO_1198 (O_1198,N_26482,N_25906);
or UO_1199 (O_1199,N_25430,N_28246);
or UO_1200 (O_1200,N_28080,N_29991);
xnor UO_1201 (O_1201,N_27719,N_27199);
nand UO_1202 (O_1202,N_28966,N_25308);
nand UO_1203 (O_1203,N_28348,N_26800);
and UO_1204 (O_1204,N_28925,N_27520);
and UO_1205 (O_1205,N_26303,N_29520);
nand UO_1206 (O_1206,N_29863,N_28123);
and UO_1207 (O_1207,N_29205,N_27202);
xnor UO_1208 (O_1208,N_27847,N_28475);
or UO_1209 (O_1209,N_29013,N_25496);
or UO_1210 (O_1210,N_27421,N_28250);
and UO_1211 (O_1211,N_26867,N_26923);
or UO_1212 (O_1212,N_27077,N_27562);
and UO_1213 (O_1213,N_26115,N_25807);
or UO_1214 (O_1214,N_28453,N_27961);
nand UO_1215 (O_1215,N_27648,N_27346);
and UO_1216 (O_1216,N_27558,N_29009);
or UO_1217 (O_1217,N_29278,N_26261);
and UO_1218 (O_1218,N_27540,N_29063);
or UO_1219 (O_1219,N_29868,N_25796);
and UO_1220 (O_1220,N_26801,N_27803);
nand UO_1221 (O_1221,N_25557,N_25864);
and UO_1222 (O_1222,N_25733,N_25022);
or UO_1223 (O_1223,N_25646,N_29488);
and UO_1224 (O_1224,N_25207,N_29296);
and UO_1225 (O_1225,N_25035,N_26943);
nor UO_1226 (O_1226,N_25014,N_29565);
nor UO_1227 (O_1227,N_28816,N_27812);
nor UO_1228 (O_1228,N_26926,N_27730);
nor UO_1229 (O_1229,N_26971,N_29420);
nand UO_1230 (O_1230,N_29008,N_28038);
nand UO_1231 (O_1231,N_28319,N_27333);
or UO_1232 (O_1232,N_29866,N_25006);
nor UO_1233 (O_1233,N_27353,N_25376);
nand UO_1234 (O_1234,N_29249,N_28023);
and UO_1235 (O_1235,N_29115,N_25504);
and UO_1236 (O_1236,N_29951,N_29290);
nor UO_1237 (O_1237,N_28152,N_25902);
nor UO_1238 (O_1238,N_28465,N_27174);
or UO_1239 (O_1239,N_25895,N_26582);
nand UO_1240 (O_1240,N_28142,N_29032);
nor UO_1241 (O_1241,N_25975,N_28604);
or UO_1242 (O_1242,N_27757,N_29260);
and UO_1243 (O_1243,N_29495,N_26778);
and UO_1244 (O_1244,N_27813,N_27178);
nand UO_1245 (O_1245,N_27066,N_27301);
nand UO_1246 (O_1246,N_26895,N_29468);
nor UO_1247 (O_1247,N_25024,N_25442);
nand UO_1248 (O_1248,N_27869,N_27434);
nor UO_1249 (O_1249,N_28425,N_28858);
or UO_1250 (O_1250,N_25306,N_27234);
nand UO_1251 (O_1251,N_29715,N_28487);
xor UO_1252 (O_1252,N_27476,N_25756);
xor UO_1253 (O_1253,N_27371,N_28703);
nor UO_1254 (O_1254,N_29332,N_28720);
and UO_1255 (O_1255,N_28567,N_26163);
and UO_1256 (O_1256,N_27288,N_29964);
and UO_1257 (O_1257,N_28812,N_25717);
and UO_1258 (O_1258,N_26150,N_29452);
nand UO_1259 (O_1259,N_26280,N_27940);
nor UO_1260 (O_1260,N_27070,N_28690);
nor UO_1261 (O_1261,N_26661,N_28253);
or UO_1262 (O_1262,N_27317,N_25259);
and UO_1263 (O_1263,N_26937,N_27939);
or UO_1264 (O_1264,N_27605,N_26225);
xnor UO_1265 (O_1265,N_28017,N_26990);
nor UO_1266 (O_1266,N_25450,N_25358);
and UO_1267 (O_1267,N_29200,N_28256);
nor UO_1268 (O_1268,N_26152,N_28747);
xnor UO_1269 (O_1269,N_27444,N_29947);
nor UO_1270 (O_1270,N_28421,N_29137);
nor UO_1271 (O_1271,N_26709,N_28605);
nor UO_1272 (O_1272,N_27096,N_25100);
and UO_1273 (O_1273,N_27445,N_29773);
nor UO_1274 (O_1274,N_29768,N_26181);
nand UO_1275 (O_1275,N_29704,N_27235);
nor UO_1276 (O_1276,N_25856,N_27801);
or UO_1277 (O_1277,N_29443,N_27921);
or UO_1278 (O_1278,N_27079,N_29215);
nand UO_1279 (O_1279,N_28004,N_27717);
or UO_1280 (O_1280,N_28340,N_25931);
nor UO_1281 (O_1281,N_28266,N_28169);
nand UO_1282 (O_1282,N_28400,N_29703);
or UO_1283 (O_1283,N_28773,N_29523);
nor UO_1284 (O_1284,N_28204,N_28415);
and UO_1285 (O_1285,N_29660,N_26765);
and UO_1286 (O_1286,N_26967,N_29100);
nor UO_1287 (O_1287,N_28331,N_29572);
or UO_1288 (O_1288,N_26729,N_26878);
or UO_1289 (O_1289,N_28354,N_28680);
or UO_1290 (O_1290,N_28512,N_29154);
nand UO_1291 (O_1291,N_28582,N_27433);
nand UO_1292 (O_1292,N_27527,N_29316);
and UO_1293 (O_1293,N_27553,N_25554);
and UO_1294 (O_1294,N_26048,N_28770);
and UO_1295 (O_1295,N_25180,N_29333);
nand UO_1296 (O_1296,N_26556,N_27701);
nand UO_1297 (O_1297,N_27649,N_25706);
nand UO_1298 (O_1298,N_25620,N_27179);
xor UO_1299 (O_1299,N_27193,N_29392);
nand UO_1300 (O_1300,N_25240,N_29522);
and UO_1301 (O_1301,N_28749,N_26419);
nand UO_1302 (O_1302,N_29975,N_29341);
xnor UO_1303 (O_1303,N_29604,N_26349);
and UO_1304 (O_1304,N_28799,N_28267);
xnor UO_1305 (O_1305,N_25470,N_27912);
nor UO_1306 (O_1306,N_27983,N_28140);
and UO_1307 (O_1307,N_26052,N_28830);
nor UO_1308 (O_1308,N_28648,N_25092);
and UO_1309 (O_1309,N_26703,N_26341);
and UO_1310 (O_1310,N_29985,N_26618);
or UO_1311 (O_1311,N_26017,N_27817);
or UO_1312 (O_1312,N_29901,N_29748);
and UO_1313 (O_1313,N_25432,N_28979);
nor UO_1314 (O_1314,N_29590,N_27597);
and UO_1315 (O_1315,N_28692,N_27601);
or UO_1316 (O_1316,N_29192,N_26513);
nand UO_1317 (O_1317,N_27177,N_25015);
and UO_1318 (O_1318,N_27635,N_29179);
nor UO_1319 (O_1319,N_26969,N_25166);
nor UO_1320 (O_1320,N_29722,N_25837);
nand UO_1321 (O_1321,N_25193,N_28653);
and UO_1322 (O_1322,N_27681,N_29797);
and UO_1323 (O_1323,N_29808,N_26941);
nor UO_1324 (O_1324,N_26435,N_26316);
and UO_1325 (O_1325,N_26269,N_25655);
nor UO_1326 (O_1326,N_27013,N_28317);
or UO_1327 (O_1327,N_29735,N_27201);
xor UO_1328 (O_1328,N_25352,N_27125);
nand UO_1329 (O_1329,N_29270,N_25242);
nor UO_1330 (O_1330,N_26173,N_26441);
nor UO_1331 (O_1331,N_26085,N_25651);
nand UO_1332 (O_1332,N_26533,N_27667);
nand UO_1333 (O_1333,N_26958,N_29665);
nand UO_1334 (O_1334,N_25650,N_29320);
nand UO_1335 (O_1335,N_28767,N_26905);
and UO_1336 (O_1336,N_25797,N_28841);
xor UO_1337 (O_1337,N_27967,N_26362);
or UO_1338 (O_1338,N_25682,N_28717);
nand UO_1339 (O_1339,N_27606,N_29917);
or UO_1340 (O_1340,N_26863,N_26331);
nor UO_1341 (O_1341,N_26343,N_29080);
nand UO_1342 (O_1342,N_27758,N_29853);
and UO_1343 (O_1343,N_28474,N_26003);
or UO_1344 (O_1344,N_25068,N_28632);
xnor UO_1345 (O_1345,N_29755,N_25372);
nor UO_1346 (O_1346,N_28096,N_25998);
or UO_1347 (O_1347,N_27005,N_25689);
nor UO_1348 (O_1348,N_28837,N_27825);
nand UO_1349 (O_1349,N_25337,N_29878);
and UO_1350 (O_1350,N_27417,N_27031);
and UO_1351 (O_1351,N_28930,N_26714);
and UO_1352 (O_1352,N_28805,N_28156);
and UO_1353 (O_1353,N_29736,N_29575);
nor UO_1354 (O_1354,N_29960,N_26055);
nor UO_1355 (O_1355,N_26634,N_28775);
and UO_1356 (O_1356,N_27620,N_26597);
or UO_1357 (O_1357,N_27822,N_28714);
nor UO_1358 (O_1358,N_25594,N_29053);
or UO_1359 (O_1359,N_27893,N_26565);
or UO_1360 (O_1360,N_26203,N_27806);
or UO_1361 (O_1361,N_25285,N_28999);
or UO_1362 (O_1362,N_27584,N_29583);
or UO_1363 (O_1363,N_27492,N_28556);
and UO_1364 (O_1364,N_28243,N_29702);
nor UO_1365 (O_1365,N_26632,N_28109);
nand UO_1366 (O_1366,N_25825,N_28811);
and UO_1367 (O_1367,N_25848,N_27870);
nor UO_1368 (O_1368,N_27800,N_27630);
and UO_1369 (O_1369,N_28259,N_29912);
nand UO_1370 (O_1370,N_27420,N_27339);
or UO_1371 (O_1371,N_28704,N_25250);
or UO_1372 (O_1372,N_26256,N_27943);
and UO_1373 (O_1373,N_26410,N_27368);
nand UO_1374 (O_1374,N_28589,N_28986);
nand UO_1375 (O_1375,N_29087,N_27137);
and UO_1376 (O_1376,N_25371,N_27892);
nor UO_1377 (O_1377,N_28611,N_25738);
and UO_1378 (O_1378,N_26126,N_26917);
nand UO_1379 (O_1379,N_29234,N_26866);
or UO_1380 (O_1380,N_26827,N_27874);
or UO_1381 (O_1381,N_27732,N_26742);
xor UO_1382 (O_1382,N_29844,N_29593);
nand UO_1383 (O_1383,N_29942,N_26826);
and UO_1384 (O_1384,N_26102,N_25293);
xor UO_1385 (O_1385,N_25663,N_28495);
nand UO_1386 (O_1386,N_25576,N_28890);
and UO_1387 (O_1387,N_27432,N_29262);
and UO_1388 (O_1388,N_26527,N_27766);
or UO_1389 (O_1389,N_25324,N_27080);
nand UO_1390 (O_1390,N_27059,N_29135);
or UO_1391 (O_1391,N_26027,N_29431);
or UO_1392 (O_1392,N_25996,N_25436);
and UO_1393 (O_1393,N_26413,N_26135);
nor UO_1394 (O_1394,N_26545,N_27068);
or UO_1395 (O_1395,N_28850,N_26072);
nand UO_1396 (O_1396,N_28909,N_29271);
nand UO_1397 (O_1397,N_28734,N_26946);
and UO_1398 (O_1398,N_28143,N_27502);
or UO_1399 (O_1399,N_29653,N_25234);
nor UO_1400 (O_1400,N_27815,N_28022);
or UO_1401 (O_1401,N_27145,N_25899);
or UO_1402 (O_1402,N_26512,N_26404);
nand UO_1403 (O_1403,N_27679,N_29651);
xor UO_1404 (O_1404,N_29467,N_28542);
and UO_1405 (O_1405,N_27593,N_26468);
and UO_1406 (O_1406,N_29823,N_29482);
xnor UO_1407 (O_1407,N_27778,N_26787);
or UO_1408 (O_1408,N_29348,N_27334);
or UO_1409 (O_1409,N_29625,N_29534);
or UO_1410 (O_1410,N_25110,N_27307);
or UO_1411 (O_1411,N_28626,N_27867);
xor UO_1412 (O_1412,N_25058,N_25182);
and UO_1413 (O_1413,N_27229,N_26045);
nor UO_1414 (O_1414,N_25317,N_28302);
or UO_1415 (O_1415,N_25769,N_27086);
xor UO_1416 (O_1416,N_27471,N_25174);
nand UO_1417 (O_1417,N_28349,N_27925);
or UO_1418 (O_1418,N_26322,N_26854);
nor UO_1419 (O_1419,N_25870,N_26412);
and UO_1420 (O_1420,N_25164,N_29329);
and UO_1421 (O_1421,N_26853,N_29360);
nand UO_1422 (O_1422,N_26901,N_29435);
and UO_1423 (O_1423,N_26475,N_29336);
or UO_1424 (O_1424,N_29872,N_25300);
nand UO_1425 (O_1425,N_29681,N_28781);
nand UO_1426 (O_1426,N_25168,N_25753);
nand UO_1427 (O_1427,N_26392,N_29163);
or UO_1428 (O_1428,N_27295,N_28110);
and UO_1429 (O_1429,N_25183,N_29481);
or UO_1430 (O_1430,N_26467,N_27840);
and UO_1431 (O_1431,N_29839,N_29732);
nand UO_1432 (O_1432,N_28365,N_27286);
nor UO_1433 (O_1433,N_26414,N_29440);
or UO_1434 (O_1434,N_29304,N_28055);
and UO_1435 (O_1435,N_29643,N_29509);
nor UO_1436 (O_1436,N_26260,N_29846);
nor UO_1437 (O_1437,N_27361,N_29935);
nand UO_1438 (O_1438,N_27290,N_26462);
nor UO_1439 (O_1439,N_25464,N_28769);
or UO_1440 (O_1440,N_27864,N_28956);
nand UO_1441 (O_1441,N_28508,N_26216);
and UO_1442 (O_1442,N_25524,N_26907);
nand UO_1443 (O_1443,N_26175,N_26153);
or UO_1444 (O_1444,N_26184,N_26641);
nor UO_1445 (O_1445,N_29925,N_28009);
and UO_1446 (O_1446,N_25275,N_29071);
xor UO_1447 (O_1447,N_25585,N_25138);
nand UO_1448 (O_1448,N_29273,N_29338);
or UO_1449 (O_1449,N_26158,N_26335);
nand UO_1450 (O_1450,N_28214,N_27367);
nand UO_1451 (O_1451,N_25966,N_26069);
xnor UO_1452 (O_1452,N_26773,N_27281);
nor UO_1453 (O_1453,N_26088,N_27784);
or UO_1454 (O_1454,N_25664,N_29892);
xnor UO_1455 (O_1455,N_26297,N_27435);
xor UO_1456 (O_1456,N_28078,N_25510);
and UO_1457 (O_1457,N_25471,N_28328);
nand UO_1458 (O_1458,N_25419,N_26530);
nor UO_1459 (O_1459,N_28387,N_27563);
nor UO_1460 (O_1460,N_26595,N_29011);
or UO_1461 (O_1461,N_25056,N_27425);
nor UO_1462 (O_1462,N_25041,N_28535);
nor UO_1463 (O_1463,N_27023,N_28434);
nor UO_1464 (O_1464,N_29796,N_27140);
nand UO_1465 (O_1465,N_28310,N_29326);
or UO_1466 (O_1466,N_29692,N_29463);
nand UO_1467 (O_1467,N_29190,N_28330);
or UO_1468 (O_1468,N_26416,N_26148);
nor UO_1469 (O_1469,N_27441,N_25860);
xnor UO_1470 (O_1470,N_25360,N_29765);
nor UO_1471 (O_1471,N_28257,N_28245);
or UO_1472 (O_1472,N_25327,N_29155);
nand UO_1473 (O_1473,N_28133,N_28656);
and UO_1474 (O_1474,N_29478,N_25016);
nand UO_1475 (O_1475,N_25427,N_25981);
xnor UO_1476 (O_1476,N_26684,N_26320);
nor UO_1477 (O_1477,N_27655,N_29042);
nor UO_1478 (O_1478,N_29698,N_28088);
xnor UO_1479 (O_1479,N_26014,N_29226);
or UO_1480 (O_1480,N_28912,N_26143);
nand UO_1481 (O_1481,N_25840,N_27189);
and UO_1482 (O_1482,N_25222,N_27781);
nand UO_1483 (O_1483,N_27877,N_26271);
nand UO_1484 (O_1484,N_25531,N_27919);
nor UO_1485 (O_1485,N_29112,N_28681);
nand UO_1486 (O_1486,N_29302,N_29334);
nand UO_1487 (O_1487,N_29760,N_29992);
and UO_1488 (O_1488,N_25494,N_28888);
nor UO_1489 (O_1489,N_29813,N_25987);
and UO_1490 (O_1490,N_29789,N_25096);
or UO_1491 (O_1491,N_28481,N_29562);
xnor UO_1492 (O_1492,N_25897,N_28284);
or UO_1493 (O_1493,N_27588,N_29024);
and UO_1494 (O_1494,N_28855,N_27104);
nand UO_1495 (O_1495,N_27734,N_26912);
and UO_1496 (O_1496,N_26690,N_28521);
and UO_1497 (O_1497,N_25967,N_28938);
xor UO_1498 (O_1498,N_29842,N_27374);
nor UO_1499 (O_1499,N_27388,N_29070);
nand UO_1500 (O_1500,N_28190,N_25054);
and UO_1501 (O_1501,N_27297,N_29779);
or UO_1502 (O_1502,N_26453,N_25463);
nand UO_1503 (O_1503,N_26589,N_25792);
nor UO_1504 (O_1504,N_25026,N_28342);
nor UO_1505 (O_1505,N_26829,N_28274);
and UO_1506 (O_1506,N_25988,N_26608);
nor UO_1507 (O_1507,N_27215,N_25724);
or UO_1508 (O_1508,N_26848,N_29963);
nor UO_1509 (O_1509,N_28431,N_29739);
and UO_1510 (O_1510,N_25867,N_25699);
nand UO_1511 (O_1511,N_26459,N_28455);
nand UO_1512 (O_1512,N_28727,N_26730);
and UO_1513 (O_1513,N_25311,N_25178);
nand UO_1514 (O_1514,N_29365,N_26779);
nand UO_1515 (O_1515,N_29709,N_28070);
or UO_1516 (O_1516,N_28446,N_29345);
and UO_1517 (O_1517,N_27185,N_25622);
nand UO_1518 (O_1518,N_28591,N_28937);
nor UO_1519 (O_1519,N_27518,N_26675);
or UO_1520 (O_1520,N_29595,N_27469);
nor UO_1521 (O_1521,N_27535,N_25083);
and UO_1522 (O_1522,N_27878,N_27555);
nor UO_1523 (O_1523,N_28639,N_25610);
and UO_1524 (O_1524,N_28315,N_26354);
and UO_1525 (O_1525,N_29377,N_29187);
or UO_1526 (O_1526,N_28411,N_25440);
or UO_1527 (O_1527,N_29659,N_29027);
nor UO_1528 (O_1528,N_25043,N_28590);
xor UO_1529 (O_1529,N_26373,N_25040);
nor UO_1530 (O_1530,N_27782,N_29731);
and UO_1531 (O_1531,N_27657,N_29165);
or UO_1532 (O_1532,N_28164,N_28755);
and UO_1533 (O_1533,N_26951,N_27447);
and UO_1534 (O_1534,N_27446,N_25131);
or UO_1535 (O_1535,N_26561,N_27510);
and UO_1536 (O_1536,N_26063,N_26658);
nor UO_1537 (O_1537,N_28224,N_27754);
nor UO_1538 (O_1538,N_26359,N_28922);
or UO_1539 (O_1539,N_25373,N_27442);
nand UO_1540 (O_1540,N_29108,N_26405);
nand UO_1541 (O_1541,N_26310,N_26888);
nand UO_1542 (O_1542,N_27639,N_28366);
nor UO_1543 (O_1543,N_29281,N_29119);
or UO_1544 (O_1544,N_27764,N_27259);
and UO_1545 (O_1545,N_27095,N_28056);
nand UO_1546 (O_1546,N_26319,N_25676);
nor UO_1547 (O_1547,N_28054,N_26758);
nand UO_1548 (O_1548,N_26613,N_29973);
nor UO_1549 (O_1549,N_25703,N_27115);
or UO_1550 (O_1550,N_29142,N_29423);
xor UO_1551 (O_1551,N_25951,N_27937);
nor UO_1552 (O_1552,N_27002,N_25558);
and UO_1553 (O_1553,N_29894,N_25349);
nor UO_1554 (O_1554,N_27437,N_25534);
and UO_1555 (O_1555,N_29157,N_28248);
or UO_1556 (O_1556,N_29882,N_28949);
nor UO_1557 (O_1557,N_25644,N_29599);
nor UO_1558 (O_1558,N_27647,N_28869);
nand UO_1559 (O_1559,N_25238,N_25708);
and UO_1560 (O_1560,N_27787,N_25157);
nand UO_1561 (O_1561,N_29929,N_26000);
nand UO_1562 (O_1562,N_29580,N_27688);
nor UO_1563 (O_1563,N_25148,N_29194);
or UO_1564 (O_1564,N_27260,N_25798);
nand UO_1565 (O_1565,N_27500,N_29679);
nand UO_1566 (O_1566,N_25519,N_28846);
xor UO_1567 (O_1567,N_27138,N_26849);
nand UO_1568 (O_1568,N_27352,N_28819);
nor UO_1569 (O_1569,N_28007,N_28264);
and UO_1570 (O_1570,N_27244,N_26583);
and UO_1571 (O_1571,N_28202,N_26785);
nor UO_1572 (O_1572,N_26463,N_29570);
and UO_1573 (O_1573,N_29670,N_28561);
nand UO_1574 (O_1574,N_28171,N_29616);
or UO_1575 (O_1575,N_26327,N_25695);
nand UO_1576 (O_1576,N_28019,N_25158);
or UO_1577 (O_1577,N_26963,N_27194);
and UO_1578 (O_1578,N_25198,N_25776);
nor UO_1579 (O_1579,N_25892,N_27722);
and UO_1580 (O_1580,N_27525,N_26123);
or UO_1581 (O_1581,N_27665,N_28057);
xor UO_1582 (O_1582,N_27712,N_27918);
and UO_1583 (O_1583,N_29918,N_27327);
or UO_1584 (O_1584,N_29861,N_26465);
xor UO_1585 (O_1585,N_27578,N_25657);
or UO_1586 (O_1586,N_25047,N_28272);
and UO_1587 (O_1587,N_26603,N_28658);
nor UO_1588 (O_1588,N_25127,N_25562);
or UO_1589 (O_1589,N_27213,N_26877);
nand UO_1590 (O_1590,N_28571,N_25719);
nand UO_1591 (O_1591,N_29507,N_28625);
or UO_1592 (O_1592,N_28705,N_26012);
xor UO_1593 (O_1593,N_28097,N_27459);
nor UO_1594 (O_1594,N_27337,N_29368);
or UO_1595 (O_1595,N_27993,N_26011);
or UO_1596 (O_1596,N_28733,N_26064);
nand UO_1597 (O_1597,N_25701,N_28114);
or UO_1598 (O_1598,N_28158,N_28111);
nand UO_1599 (O_1599,N_26584,N_25940);
nand UO_1600 (O_1600,N_26387,N_29323);
nor UO_1601 (O_1601,N_28121,N_29549);
and UO_1602 (O_1602,N_28260,N_29907);
nand UO_1603 (O_1603,N_27935,N_29293);
nand UO_1604 (O_1604,N_27542,N_26695);
and UO_1605 (O_1605,N_27278,N_27997);
and UO_1606 (O_1606,N_28881,N_29034);
or UO_1607 (O_1607,N_27957,N_25969);
and UO_1608 (O_1608,N_27154,N_28948);
and UO_1609 (O_1609,N_28726,N_29623);
nor UO_1610 (O_1610,N_26510,N_27287);
and UO_1611 (O_1611,N_28964,N_28575);
xor UO_1612 (O_1612,N_26874,N_29588);
nor UO_1613 (O_1613,N_27916,N_26431);
and UO_1614 (O_1614,N_29711,N_29802);
nor UO_1615 (O_1615,N_29019,N_26101);
xor UO_1616 (O_1616,N_26824,N_27557);
or UO_1617 (O_1617,N_25227,N_27134);
xnor UO_1618 (O_1618,N_25177,N_29515);
and UO_1619 (O_1619,N_25928,N_28878);
and UO_1620 (O_1620,N_29018,N_28970);
nor UO_1621 (O_1621,N_26355,N_27691);
and UO_1622 (O_1622,N_27880,N_29680);
nand UO_1623 (O_1623,N_26117,N_26833);
xnor UO_1624 (O_1624,N_29259,N_25884);
nand UO_1625 (O_1625,N_29048,N_27242);
and UO_1626 (O_1626,N_25067,N_26223);
and UO_1627 (O_1627,N_28549,N_29369);
and UO_1628 (O_1628,N_25532,N_26786);
nor UO_1629 (O_1629,N_27932,N_29465);
and UO_1630 (O_1630,N_28012,N_25348);
nand UO_1631 (O_1631,N_26111,N_26066);
or UO_1632 (O_1632,N_28407,N_25443);
or UO_1633 (O_1633,N_27633,N_26305);
and UO_1634 (O_1634,N_29106,N_26998);
or UO_1635 (O_1635,N_28035,N_28301);
or UO_1636 (O_1636,N_28935,N_28287);
nor UO_1637 (O_1637,N_25909,N_27792);
nor UO_1638 (O_1638,N_26338,N_28965);
and UO_1639 (O_1639,N_25782,N_25838);
nor UO_1640 (O_1640,N_25199,N_26569);
xor UO_1641 (O_1641,N_26034,N_28160);
nand UO_1642 (O_1642,N_27659,N_25224);
xor UO_1643 (O_1643,N_25061,N_28159);
and UO_1644 (O_1644,N_26624,N_29536);
and UO_1645 (O_1645,N_25790,N_27141);
and UO_1646 (O_1646,N_25028,N_29288);
nor UO_1647 (O_1647,N_27986,N_27868);
nand UO_1648 (O_1648,N_25965,N_29893);
nor UO_1649 (O_1649,N_27389,N_26989);
and UO_1650 (O_1650,N_27146,N_28189);
and UO_1651 (O_1651,N_25210,N_26550);
nand UO_1652 (O_1652,N_28437,N_29571);
and UO_1653 (O_1653,N_25129,N_29138);
nor UO_1654 (O_1654,N_27624,N_25316);
nand UO_1655 (O_1655,N_29387,N_28072);
nor UO_1656 (O_1656,N_28106,N_29895);
xor UO_1657 (O_1657,N_27756,N_29803);
nor UO_1658 (O_1658,N_25613,N_26433);
xor UO_1659 (O_1659,N_26417,N_28876);
xnor UO_1660 (O_1660,N_25472,N_26350);
and UO_1661 (O_1661,N_25865,N_26129);
nor UO_1662 (O_1662,N_26707,N_27733);
xor UO_1663 (O_1663,N_29666,N_26084);
nand UO_1664 (O_1664,N_26502,N_29022);
nor UO_1665 (O_1665,N_26664,N_25616);
nand UO_1666 (O_1666,N_27279,N_29664);
and UO_1667 (O_1667,N_28198,N_29261);
nand UO_1668 (O_1668,N_26838,N_26559);
nor UO_1669 (O_1669,N_28560,N_25748);
nand UO_1670 (O_1670,N_25344,N_27363);
and UO_1671 (O_1671,N_29694,N_29983);
nor UO_1672 (O_1672,N_28960,N_27715);
xnor UO_1673 (O_1673,N_26736,N_26456);
and UO_1674 (O_1674,N_28027,N_25960);
and UO_1675 (O_1675,N_27310,N_29528);
and UO_1676 (O_1676,N_29035,N_26267);
nor UO_1677 (O_1677,N_25339,N_29116);
or UO_1678 (O_1678,N_26365,N_28008);
or UO_1679 (O_1679,N_29357,N_26509);
nor UO_1680 (O_1680,N_29073,N_25126);
xor UO_1681 (O_1681,N_28882,N_29741);
and UO_1682 (O_1682,N_25333,N_25956);
or UO_1683 (O_1683,N_29126,N_26450);
and UO_1684 (O_1684,N_25215,N_28622);
and UO_1685 (O_1685,N_26916,N_27728);
xor UO_1686 (O_1686,N_28974,N_27514);
or UO_1687 (O_1687,N_27392,N_25270);
nand UO_1688 (O_1688,N_27157,N_29174);
xnor UO_1689 (O_1689,N_25192,N_27083);
nor UO_1690 (O_1690,N_25783,N_26657);
nand UO_1691 (O_1691,N_27034,N_28438);
or UO_1692 (O_1692,N_25569,N_28661);
and UO_1693 (O_1693,N_28832,N_25762);
nor UO_1694 (O_1694,N_25905,N_28725);
nand UO_1695 (O_1695,N_29970,N_29279);
and UO_1696 (O_1696,N_28127,N_28423);
and UO_1697 (O_1697,N_25548,N_26754);
xnor UO_1698 (O_1698,N_27670,N_26213);
xor UO_1699 (O_1699,N_26352,N_29311);
or UO_1700 (O_1700,N_27144,N_28719);
and UO_1701 (O_1701,N_27506,N_28176);
and UO_1702 (O_1702,N_25915,N_26788);
or UO_1703 (O_1703,N_27911,N_28255);
nor UO_1704 (O_1704,N_25827,N_25605);
or UO_1705 (O_1705,N_27401,N_28636);
or UO_1706 (O_1706,N_25526,N_26179);
nor UO_1707 (O_1707,N_26570,N_25971);
xnor UO_1708 (O_1708,N_25124,N_26022);
nand UO_1709 (O_1709,N_27273,N_26333);
or UO_1710 (O_1710,N_29188,N_26445);
nand UO_1711 (O_1711,N_25750,N_27303);
nand UO_1712 (O_1712,N_27552,N_28439);
nand UO_1713 (O_1713,N_26981,N_25736);
and UO_1714 (O_1714,N_25944,N_29363);
nor UO_1715 (O_1715,N_27291,N_25179);
or UO_1716 (O_1716,N_27512,N_28652);
nand UO_1717 (O_1717,N_25789,N_26024);
and UO_1718 (O_1718,N_27992,N_25269);
or UO_1719 (O_1719,N_27941,N_27736);
xor UO_1720 (O_1720,N_26276,N_27373);
or UO_1721 (O_1721,N_26836,N_25926);
nor UO_1722 (O_1722,N_29425,N_26628);
or UO_1723 (O_1723,N_25468,N_26099);
nand UO_1724 (O_1724,N_28268,N_29826);
nor UO_1725 (O_1725,N_27120,N_28420);
nor UO_1726 (O_1726,N_25765,N_26881);
or UO_1727 (O_1727,N_27056,N_25105);
or UO_1728 (O_1728,N_26096,N_27113);
xnor UO_1729 (O_1729,N_27964,N_29804);
or UO_1730 (O_1730,N_29117,N_29573);
nor UO_1731 (O_1731,N_29956,N_28529);
and UO_1732 (O_1732,N_27366,N_28185);
or UO_1733 (O_1733,N_29821,N_25021);
or UO_1734 (O_1734,N_28377,N_27602);
or UO_1735 (O_1735,N_28546,N_29751);
xnor UO_1736 (O_1736,N_26928,N_27133);
xnor UO_1737 (O_1737,N_28040,N_29000);
or UO_1738 (O_1738,N_28568,N_27544);
nor UO_1739 (O_1739,N_29763,N_27186);
or UO_1740 (O_1740,N_28394,N_25391);
xnor UO_1741 (O_1741,N_28086,N_25321);
and UO_1742 (O_1742,N_26231,N_27906);
and UO_1743 (O_1743,N_25437,N_29464);
nor UO_1744 (O_1744,N_25924,N_29030);
or UO_1745 (O_1745,N_27583,N_28406);
xor UO_1746 (O_1746,N_26702,N_28408);
or UO_1747 (O_1747,N_26364,N_28914);
or UO_1748 (O_1748,N_28649,N_27131);
and UO_1749 (O_1749,N_26428,N_29774);
and UO_1750 (O_1750,N_28061,N_29867);
or UO_1751 (O_1751,N_29105,N_28564);
or UO_1752 (O_1752,N_26820,N_28784);
or UO_1753 (O_1753,N_27039,N_26018);
nor UO_1754 (O_1754,N_26470,N_26049);
nand UO_1755 (O_1755,N_25598,N_26274);
and UO_1756 (O_1756,N_25984,N_26791);
nand UO_1757 (O_1757,N_26407,N_26448);
nor UO_1758 (O_1758,N_26750,N_29533);
or UO_1759 (O_1759,N_28857,N_28616);
nand UO_1760 (O_1760,N_28451,N_27851);
nand UO_1761 (O_1761,N_27789,N_26563);
or UO_1762 (O_1762,N_25304,N_28021);
xnor UO_1763 (O_1763,N_27658,N_26283);
nand UO_1764 (O_1764,N_25871,N_28168);
or UO_1765 (O_1765,N_26029,N_29608);
nand UO_1766 (O_1766,N_29676,N_29682);
or UO_1767 (O_1767,N_29948,N_26258);
nor UO_1768 (O_1768,N_25217,N_27158);
or UO_1769 (O_1769,N_26079,N_29268);
xnor UO_1770 (O_1770,N_26728,N_26540);
and UO_1771 (O_1771,N_28511,N_26020);
nand UO_1772 (O_1772,N_28047,N_29223);
nor UO_1773 (O_1773,N_29222,N_29454);
and UO_1774 (O_1774,N_29003,N_27674);
and UO_1775 (O_1775,N_28327,N_28810);
nor UO_1776 (O_1776,N_25410,N_27203);
nand UO_1777 (O_1777,N_28131,N_28910);
nor UO_1778 (O_1778,N_26171,N_26183);
nand UO_1779 (O_1779,N_27466,N_25773);
and UO_1780 (O_1780,N_27161,N_28608);
or UO_1781 (O_1781,N_26330,N_29258);
nor UO_1782 (O_1782,N_27791,N_29532);
or UO_1783 (O_1783,N_26805,N_28314);
and UO_1784 (O_1784,N_29811,N_27573);
nand UO_1785 (O_1785,N_28728,N_29889);
and UO_1786 (O_1786,N_26346,N_26977);
and UO_1787 (O_1787,N_29390,N_25509);
nand UO_1788 (O_1788,N_26233,N_25449);
nand UO_1789 (O_1789,N_29924,N_29094);
xnor UO_1790 (O_1790,N_26047,N_27490);
nand UO_1791 (O_1791,N_28545,N_26500);
or UO_1792 (O_1792,N_25904,N_27316);
or UO_1793 (O_1793,N_27889,N_27326);
or UO_1794 (O_1794,N_29726,N_27636);
xnor UO_1795 (O_1795,N_28430,N_27650);
nor UO_1796 (O_1796,N_26956,N_25121);
and UO_1797 (O_1797,N_29567,N_26585);
nand UO_1798 (O_1798,N_28296,N_25280);
and UO_1799 (O_1799,N_26575,N_27798);
or UO_1800 (O_1800,N_29406,N_28889);
and UO_1801 (O_1801,N_25412,N_27955);
and UO_1802 (O_1802,N_29933,N_29201);
nand UO_1803 (O_1803,N_26279,N_29083);
nor UO_1804 (O_1804,N_28129,N_27296);
nand UO_1805 (O_1805,N_26222,N_25001);
or UO_1806 (O_1806,N_29110,N_25578);
and UO_1807 (O_1807,N_26442,N_29450);
nor UO_1808 (O_1808,N_25809,N_29152);
and UO_1809 (O_1809,N_25852,N_27478);
and UO_1810 (O_1810,N_27920,N_28814);
xor UO_1811 (O_1811,N_25414,N_27375);
nand UO_1812 (O_1812,N_26666,N_28780);
nor UO_1813 (O_1813,N_29782,N_27872);
nand UO_1814 (O_1814,N_26680,N_26429);
nor UO_1815 (O_1815,N_29235,N_25629);
and UO_1816 (O_1816,N_25758,N_29927);
nand UO_1817 (O_1817,N_26086,N_29150);
and UO_1818 (O_1818,N_27741,N_26581);
nand UO_1819 (O_1819,N_29426,N_25244);
nor UO_1820 (O_1820,N_29029,N_29900);
nand UO_1821 (O_1821,N_27164,N_29224);
and UO_1822 (O_1822,N_29560,N_28184);
nor UO_1823 (O_1823,N_25589,N_28562);
xor UO_1824 (O_1824,N_26614,N_25305);
or UO_1825 (O_1825,N_28090,N_27328);
and UO_1826 (O_1826,N_29113,N_29346);
or UO_1827 (O_1827,N_28715,N_29382);
nand UO_1828 (O_1828,N_26930,N_27541);
and UO_1829 (O_1829,N_29374,N_28794);
nor UO_1830 (O_1830,N_29856,N_25446);
or UO_1831 (O_1831,N_25873,N_25545);
nor UO_1832 (O_1832,N_29944,N_27640);
and UO_1833 (O_1833,N_28724,N_29696);
or UO_1834 (O_1834,N_26600,N_27615);
or UO_1835 (O_1835,N_26131,N_27831);
or UO_1836 (O_1836,N_28861,N_28873);
nand UO_1837 (O_1837,N_27704,N_27760);
or UO_1838 (O_1838,N_28824,N_29663);
nor UO_1839 (O_1839,N_28951,N_26784);
nand UO_1840 (O_1840,N_27644,N_29240);
nand UO_1841 (O_1841,N_25075,N_25087);
or UO_1842 (O_1842,N_27611,N_29691);
and UO_1843 (O_1843,N_28309,N_26682);
nand UO_1844 (O_1844,N_25754,N_26970);
and UO_1845 (O_1845,N_26774,N_25812);
and UO_1846 (O_1846,N_25656,N_28379);
nor UO_1847 (O_1847,N_29257,N_26537);
nor UO_1848 (O_1848,N_28978,N_29005);
and UO_1849 (O_1849,N_25323,N_29411);
nand UO_1850 (O_1850,N_29516,N_26332);
nand UO_1851 (O_1851,N_27899,N_28624);
nor UO_1852 (O_1852,N_28628,N_29586);
or UO_1853 (O_1853,N_28551,N_29355);
nor UO_1854 (O_1854,N_26542,N_25592);
nor UO_1855 (O_1855,N_28083,N_26798);
nand UO_1856 (O_1856,N_29359,N_28418);
and UO_1857 (O_1857,N_26957,N_26155);
and UO_1858 (O_1858,N_25652,N_29366);
or UO_1859 (O_1859,N_27991,N_27775);
nor UO_1860 (O_1860,N_28621,N_26574);
nand UO_1861 (O_1861,N_27249,N_29652);
nand UO_1862 (O_1862,N_27069,N_29969);
or UO_1863 (O_1863,N_29511,N_28031);
nand UO_1864 (O_1864,N_28543,N_28462);
and UO_1865 (O_1865,N_27879,N_26245);
nor UO_1866 (O_1866,N_28466,N_25245);
nand UO_1867 (O_1867,N_27041,N_28766);
xor UO_1868 (O_1868,N_25980,N_27835);
nor UO_1869 (O_1869,N_28844,N_29807);
nand UO_1870 (O_1870,N_25732,N_29669);
and UO_1871 (O_1871,N_29504,N_26673);
nand UO_1872 (O_1872,N_26230,N_29322);
xor UO_1873 (O_1873,N_27043,N_26810);
nand UO_1874 (O_1874,N_27343,N_25276);
nor UO_1875 (O_1875,N_26031,N_25362);
and UO_1876 (O_1876,N_27293,N_25690);
or UO_1877 (O_1877,N_28370,N_26528);
or UO_1878 (O_1878,N_25452,N_28032);
or UO_1879 (O_1879,N_25093,N_29324);
and UO_1880 (O_1880,N_29558,N_26770);
or UO_1881 (O_1881,N_26472,N_28277);
nand UO_1882 (O_1882,N_29025,N_28066);
or UO_1883 (O_1883,N_25497,N_27669);
xor UO_1884 (O_1884,N_25225,N_29068);
xnor UO_1885 (O_1885,N_28573,N_28124);
nor UO_1886 (O_1886,N_26726,N_25212);
and UO_1887 (O_1887,N_25665,N_25550);
and UO_1888 (O_1888,N_29753,N_25680);
or UO_1889 (O_1889,N_25618,N_27740);
nor UO_1890 (O_1890,N_27231,N_25834);
and UO_1891 (O_1891,N_29010,N_25729);
and UO_1892 (O_1892,N_25149,N_26567);
or UO_1893 (O_1893,N_27608,N_27975);
nor UO_1894 (O_1894,N_29843,N_27359);
nand UO_1895 (O_1895,N_28609,N_25602);
nand UO_1896 (O_1896,N_27211,N_28305);
or UO_1897 (O_1897,N_29383,N_25320);
or UO_1898 (O_1898,N_29069,N_27745);
or UO_1899 (O_1899,N_27354,N_27511);
or UO_1900 (O_1900,N_27463,N_25103);
and UO_1901 (O_1901,N_26062,N_25752);
nor UO_1902 (O_1902,N_27372,N_25880);
xor UO_1903 (O_1903,N_25082,N_25486);
nand UO_1904 (O_1904,N_27729,N_28884);
or UO_1905 (O_1905,N_28989,N_26962);
and UO_1906 (O_1906,N_27944,N_25010);
or UO_1907 (O_1907,N_29195,N_26806);
and UO_1908 (O_1908,N_28710,N_25197);
or UO_1909 (O_1909,N_28655,N_29090);
xor UO_1910 (O_1910,N_28736,N_28191);
or UO_1911 (O_1911,N_29066,N_25582);
and UO_1912 (O_1912,N_26913,N_27311);
or UO_1913 (O_1913,N_27067,N_28145);
nor UO_1914 (O_1914,N_28234,N_28381);
nor UO_1915 (O_1915,N_25670,N_26813);
and UO_1916 (O_1916,N_27163,N_29037);
nor UO_1917 (O_1917,N_26107,N_29950);
nor UO_1918 (O_1918,N_27277,N_26492);
and UO_1919 (O_1919,N_27587,N_25151);
and UO_1920 (O_1920,N_25162,N_27030);
and UO_1921 (O_1921,N_27861,N_27191);
and UO_1922 (O_1922,N_27094,N_26460);
nand UO_1923 (O_1923,N_29381,N_27990);
or UO_1924 (O_1924,N_25580,N_26054);
nor UO_1925 (O_1925,N_26162,N_28181);
or UO_1926 (O_1926,N_27076,N_27206);
and UO_1927 (O_1927,N_27938,N_26092);
nor UO_1928 (O_1928,N_27947,N_25462);
nor UO_1929 (O_1929,N_29972,N_25932);
nor UO_1930 (O_1930,N_29244,N_26369);
nor UO_1931 (O_1931,N_28024,N_29787);
nand UO_1932 (O_1932,N_25604,N_25581);
nand UO_1933 (O_1933,N_26356,N_27857);
or UO_1934 (O_1934,N_25044,N_28756);
nor UO_1935 (O_1935,N_27188,N_27217);
xor UO_1936 (O_1936,N_25474,N_29091);
and UO_1937 (O_1937,N_27493,N_28950);
and UO_1938 (O_1938,N_27724,N_26994);
or UO_1939 (O_1939,N_26879,N_27230);
nor UO_1940 (O_1940,N_25169,N_29857);
nand UO_1941 (O_1941,N_27517,N_29276);
or UO_1942 (O_1942,N_25516,N_28442);
nor UO_1943 (O_1943,N_26161,N_26627);
or UO_1944 (O_1944,N_26689,N_26134);
nand UO_1945 (O_1945,N_25700,N_29607);
or UO_1946 (O_1946,N_29403,N_28637);
nor UO_1947 (O_1947,N_28000,N_28696);
nor UO_1948 (O_1948,N_27871,N_25346);
nand UO_1949 (O_1949,N_27933,N_27100);
xor UO_1950 (O_1950,N_29512,N_26438);
and UO_1951 (O_1951,N_29957,N_25448);
xnor UO_1952 (O_1952,N_25714,N_28991);
nand UO_1953 (O_1953,N_29657,N_28659);
nand UO_1954 (O_1954,N_28802,N_29914);
nor UO_1955 (O_1955,N_29865,N_26942);
and UO_1956 (O_1956,N_28791,N_27652);
nand UO_1957 (O_1957,N_29587,N_28701);
nand UO_1958 (O_1958,N_27332,N_29632);
or UO_1959 (O_1959,N_27168,N_29036);
nor UO_1960 (O_1960,N_26825,N_28238);
nand UO_1961 (O_1961,N_28923,N_29734);
nand UO_1962 (O_1962,N_27097,N_28963);
or UO_1963 (O_1963,N_28505,N_27651);
and UO_1964 (O_1964,N_25633,N_29031);
nor UO_1965 (O_1965,N_27003,N_28945);
nor UO_1966 (O_1966,N_26821,N_28196);
or UO_1967 (O_1967,N_28815,N_29367);
nor UO_1968 (O_1968,N_26169,N_25201);
and UO_1969 (O_1969,N_27684,N_29274);
xnor UO_1970 (O_1970,N_26617,N_29172);
nor UO_1971 (O_1971,N_25786,N_28443);
and UO_1972 (O_1972,N_25266,N_25890);
xnor UO_1973 (O_1973,N_26137,N_29178);
nor UO_1974 (O_1974,N_25508,N_29151);
nor UO_1975 (O_1975,N_25039,N_28842);
and UO_1976 (O_1976,N_29505,N_26298);
or UO_1977 (O_1977,N_25301,N_26578);
nor UO_1978 (O_1978,N_25160,N_29433);
and UO_1979 (O_1979,N_28393,N_28029);
and UO_1980 (O_1980,N_27907,N_29344);
nand UO_1981 (O_1981,N_26803,N_29162);
nand UO_1982 (O_1982,N_26638,N_27896);
nor UO_1983 (O_1983,N_29556,N_27405);
nand UO_1984 (O_1984,N_27044,N_26586);
and UO_1985 (O_1985,N_29896,N_26302);
and UO_1986 (O_1986,N_26199,N_25053);
nor UO_1987 (O_1987,N_29146,N_25625);
nand UO_1988 (O_1988,N_26265,N_28968);
nand UO_1989 (O_1989,N_26194,N_29349);
xor UO_1990 (O_1990,N_27036,N_26323);
or UO_1991 (O_1991,N_25342,N_29416);
nor UO_1992 (O_1992,N_26193,N_26921);
and UO_1993 (O_1993,N_26406,N_26986);
nand UO_1994 (O_1994,N_27394,N_27852);
nor UO_1995 (O_1995,N_26679,N_28448);
nor UO_1996 (O_1996,N_29911,N_26902);
and UO_1997 (O_1997,N_28399,N_29547);
nor UO_1998 (O_1998,N_26892,N_26508);
xnor UO_1999 (O_1999,N_26882,N_29476);
and UO_2000 (O_2000,N_27627,N_27119);
and UO_2001 (O_2001,N_29447,N_25820);
nand UO_2002 (O_2002,N_26480,N_28955);
nor UO_2003 (O_2003,N_28018,N_26491);
nor UO_2004 (O_2004,N_28141,N_29836);
and UO_2005 (O_2005,N_26525,N_27269);
nor UO_2006 (O_2006,N_25278,N_26781);
and UO_2007 (O_2007,N_26094,N_28544);
nand UO_2008 (O_2008,N_29023,N_29269);
and UO_2009 (O_2009,N_25512,N_29384);
and UO_2010 (O_2010,N_26648,N_26835);
nor UO_2011 (O_2011,N_28369,N_25081);
or UO_2012 (O_2012,N_26469,N_26165);
and UO_2013 (O_2013,N_25698,N_28261);
nand UO_2014 (O_2014,N_26217,N_29953);
nand UO_2015 (O_2015,N_25310,N_29778);
nand UO_2016 (O_2016,N_29622,N_26883);
and UO_2017 (O_2017,N_26723,N_27642);
and UO_2018 (O_2018,N_26112,N_27507);
or UO_2019 (O_2019,N_25484,N_25140);
nand UO_2020 (O_2020,N_29428,N_27111);
xnor UO_2021 (O_2021,N_28957,N_26906);
xnor UO_2022 (O_2022,N_26043,N_28318);
or UO_2023 (O_2023,N_29436,N_25295);
xor UO_2024 (O_2024,N_27890,N_28107);
and UO_2025 (O_2025,N_27055,N_29492);
nor UO_2026 (O_2026,N_26397,N_28522);
nand UO_2027 (O_2027,N_26104,N_26976);
nor UO_2028 (O_2028,N_28682,N_27403);
xnor UO_2029 (O_2029,N_25299,N_26760);
or UO_2030 (O_2030,N_26625,N_29627);
or UO_2031 (O_2031,N_27793,N_27126);
nand UO_2032 (O_2032,N_26505,N_29267);
nor UO_2033 (O_2033,N_29554,N_26232);
nor UO_2034 (O_2034,N_25515,N_28161);
xnor UO_2035 (O_2035,N_26633,N_28050);
and UO_2036 (O_2036,N_25117,N_26667);
nand UO_2037 (O_2037,N_27960,N_29880);
and UO_2038 (O_2038,N_25454,N_25603);
nand UO_2039 (O_2039,N_28339,N_29526);
nand UO_2040 (O_2040,N_25330,N_27876);
and UO_2041 (O_2041,N_28311,N_29824);
nand UO_2042 (O_2042,N_27012,N_28845);
nor UO_2043 (O_2043,N_27237,N_25520);
nor UO_2044 (O_2044,N_26361,N_27262);
nand UO_2045 (O_2045,N_26348,N_27576);
xor UO_2046 (O_2046,N_27600,N_28595);
nor UO_2047 (O_2047,N_29613,N_27409);
or UO_2048 (O_2048,N_28906,N_25247);
nor UO_2049 (O_2049,N_25319,N_28558);
nand UO_2050 (O_2050,N_29576,N_29939);
xor UO_2051 (O_2051,N_26694,N_26795);
nor UO_2052 (O_2052,N_26398,N_28946);
and UO_2053 (O_2053,N_29654,N_26794);
nor UO_2054 (O_2054,N_27569,N_27214);
nand UO_2055 (O_2055,N_29943,N_29810);
nor UO_2056 (O_2056,N_26093,N_27692);
xor UO_2057 (O_2057,N_29089,N_28074);
nand UO_2058 (O_2058,N_28718,N_27873);
and UO_2059 (O_2059,N_25090,N_27591);
and UO_2060 (O_2060,N_27102,N_25363);
nand UO_2061 (O_2061,N_26403,N_25170);
nor UO_2062 (O_2062,N_26621,N_29007);
nand UO_2063 (O_2063,N_25480,N_25048);
xnor UO_2064 (O_2064,N_27093,N_28585);
and UO_2065 (O_2065,N_28233,N_26511);
and UO_2066 (O_2066,N_28137,N_25881);
nor UO_2067 (O_2067,N_25648,N_28926);
and UO_2068 (O_2068,N_27329,N_25279);
and UO_2069 (O_2069,N_28565,N_29952);
nand UO_2070 (O_2070,N_28554,N_27393);
and UO_2071 (O_2071,N_29591,N_28014);
and UO_2072 (O_2072,N_25601,N_29134);
xor UO_2073 (O_2073,N_25514,N_25252);
and UO_2074 (O_2074,N_28936,N_28566);
nor UO_2075 (O_2075,N_27000,N_28454);
nand UO_2076 (O_2076,N_25018,N_29775);
or UO_2077 (O_2077,N_28574,N_25415);
xor UO_2078 (O_2078,N_27001,N_26670);
nand UO_2079 (O_2079,N_28132,N_25916);
or UO_2080 (O_2080,N_27682,N_27866);
or UO_2081 (O_2081,N_26108,N_26281);
nor UO_2082 (O_2082,N_28229,N_26037);
and UO_2083 (O_2083,N_28939,N_27747);
or UO_2084 (O_2084,N_26166,N_25421);
or UO_2085 (O_2085,N_27007,N_26180);
nor UO_2086 (O_2086,N_26975,N_28752);
or UO_2087 (O_2087,N_28480,N_27713);
nor UO_2088 (O_2088,N_28893,N_26439);
and UO_2089 (O_2089,N_26897,N_26752);
nand UO_2090 (O_2090,N_26423,N_26312);
nand UO_2091 (O_2091,N_28207,N_28316);
nor UO_2092 (O_2092,N_28760,N_25627);
xnor UO_2093 (O_2093,N_29393,N_29832);
nand UO_2094 (O_2094,N_26822,N_28471);
or UO_2095 (O_2095,N_25059,N_26997);
and UO_2096 (O_2096,N_29212,N_29524);
nand UO_2097 (O_2097,N_29997,N_26772);
or UO_2098 (O_2098,N_26548,N_27673);
and UO_2099 (O_2099,N_25386,N_25475);
or UO_2100 (O_2100,N_26376,N_25350);
nand UO_2101 (O_2101,N_25579,N_27860);
nand UO_2102 (O_2102,N_29247,N_28182);
and UO_2103 (O_2103,N_28052,N_28401);
nand UO_2104 (O_2104,N_29697,N_26264);
nor UO_2105 (O_2105,N_28390,N_29216);
and UO_2106 (O_2106,N_29746,N_28610);
and UO_2107 (O_2107,N_29351,N_27391);
and UO_2108 (O_2108,N_28998,N_26903);
xnor UO_2109 (O_2109,N_28959,N_25226);
nand UO_2110 (O_2110,N_29040,N_28839);
and UO_2111 (O_2111,N_25845,N_28550);
xor UO_2112 (O_2112,N_29294,N_26033);
and UO_2113 (O_2113,N_25425,N_28932);
nand UO_2114 (O_2114,N_25459,N_26345);
or UO_2115 (O_2115,N_29818,N_26860);
or UO_2116 (O_2116,N_25220,N_25894);
or UO_2117 (O_2117,N_25760,N_29145);
xnor UO_2118 (O_2118,N_25290,N_27680);
nor UO_2119 (O_2119,N_29936,N_29566);
nand UO_2120 (O_2120,N_25123,N_26819);
and UO_2121 (O_2121,N_29597,N_29979);
or UO_2122 (O_2122,N_25483,N_25976);
or UO_2123 (O_2123,N_26211,N_27355);
xor UO_2124 (O_2124,N_28299,N_28774);
or UO_2125 (O_2125,N_25688,N_28352);
and UO_2126 (O_2126,N_27360,N_27818);
xnor UO_2127 (O_2127,N_26229,N_27582);
nand UO_2128 (O_2128,N_27543,N_28188);
or UO_2129 (O_2129,N_25755,N_28981);
nand UO_2130 (O_2130,N_28091,N_29437);
nand UO_2131 (O_2131,N_27054,N_25282);
nor UO_2132 (O_2132,N_26378,N_25525);
or UO_2133 (O_2133,N_27236,N_25599);
nor UO_2134 (O_2134,N_26837,N_25938);
nand UO_2135 (O_2135,N_28405,N_28002);
nand UO_2136 (O_2136,N_27592,N_25263);
nand UO_2137 (O_2137,N_26727,N_27407);
or UO_2138 (O_2138,N_27675,N_25262);
nor UO_2139 (O_2139,N_25338,N_28693);
and UO_2140 (O_2140,N_29444,N_28120);
and UO_2141 (O_2141,N_25328,N_27571);
nand UO_2142 (O_2142,N_28470,N_28918);
and UO_2143 (O_2143,N_25833,N_25677);
or UO_2144 (O_2144,N_29928,N_26870);
and UO_2145 (O_2145,N_28367,N_27335);
nor UO_2146 (O_2146,N_29072,N_28984);
and UO_2147 (O_2147,N_29589,N_28278);
or UO_2148 (O_2148,N_29114,N_29136);
nand UO_2149 (O_2149,N_29299,N_25478);
or UO_2150 (O_2150,N_26985,N_26032);
and UO_2151 (O_2151,N_27169,N_29291);
nand UO_2152 (O_2152,N_26247,N_29641);
nor UO_2153 (O_2153,N_26761,N_25994);
and UO_2154 (O_2154,N_27255,N_29959);
and UO_2155 (O_2155,N_29689,N_26272);
nor UO_2156 (O_2156,N_28759,N_25501);
and UO_2157 (O_2157,N_25004,N_29852);
and UO_2158 (O_2158,N_28201,N_26746);
nand UO_2159 (O_2159,N_29713,N_28840);
or UO_2160 (O_2160,N_29987,N_29123);
xnor UO_2161 (O_2161,N_29395,N_25184);
nor UO_2162 (O_2162,N_26564,N_29958);
nand UO_2163 (O_2163,N_29350,N_25296);
nand UO_2164 (O_2164,N_29457,N_29399);
nor UO_2165 (O_2165,N_29725,N_28361);
or UO_2166 (O_2166,N_29081,N_25995);
or UO_2167 (O_2167,N_27965,N_26046);
or UO_2168 (O_2168,N_28798,N_27212);
nor UO_2169 (O_2169,N_28599,N_25431);
or UO_2170 (O_2170,N_26334,N_25144);
xnor UO_2171 (O_2171,N_29727,N_27482);
and UO_2172 (O_2172,N_27613,N_25132);
nor UO_2173 (O_2173,N_27233,N_28699);
nand UO_2174 (O_2174,N_29940,N_26748);
and UO_2175 (O_2175,N_27302,N_26626);
nand UO_2176 (O_2176,N_27423,N_28085);
or UO_2177 (O_2177,N_26368,N_26110);
and UO_2178 (O_2178,N_26366,N_29819);
nand UO_2179 (O_2179,N_28642,N_28618);
xnor UO_2180 (O_2180,N_28357,N_25000);
nand UO_2181 (O_2181,N_27581,N_28572);
and UO_2182 (O_2182,N_29510,N_27369);
nor UO_2183 (O_2183,N_28163,N_28678);
nand UO_2184 (O_2184,N_25375,N_25052);
and UO_2185 (O_2185,N_28126,N_26933);
xor UO_2186 (O_2186,N_27827,N_26520);
nand UO_2187 (O_2187,N_29184,N_28016);
nand UO_2188 (O_2188,N_26992,N_25970);
nand UO_2189 (O_2189,N_29419,N_29618);
or UO_2190 (O_2190,N_27443,N_28646);
nand UO_2191 (O_2191,N_27698,N_25930);
nand UO_2192 (O_2192,N_26687,N_27050);
or UO_2193 (O_2193,N_25553,N_25866);
or UO_2194 (O_2194,N_26593,N_26363);
or UO_2195 (O_2195,N_25228,N_29361);
or UO_2196 (O_2196,N_27830,N_29343);
or UO_2197 (O_2197,N_25332,N_28419);
or UO_2198 (O_2198,N_26040,N_28864);
nor UO_2199 (O_2199,N_29792,N_28071);
or UO_2200 (O_2200,N_27183,N_27018);
or UO_2201 (O_2201,N_29527,N_28062);
xor UO_2202 (O_2202,N_27398,N_26844);
or UO_2203 (O_2203,N_27107,N_27554);
nor UO_2204 (O_2204,N_25744,N_28285);
nor UO_2205 (O_2205,N_25635,N_26735);
and UO_2206 (O_2206,N_27580,N_25816);
or UO_2207 (O_2207,N_27439,N_26241);
nor UO_2208 (O_2208,N_26299,N_27984);
nand UO_2209 (O_2209,N_25055,N_26674);
and UO_2210 (O_2210,N_25433,N_28578);
and UO_2211 (O_2211,N_26722,N_27081);
and UO_2212 (O_2212,N_29644,N_29596);
and UO_2213 (O_2213,N_28449,N_25877);
and UO_2214 (O_2214,N_28221,N_27645);
nor UO_2215 (O_2215,N_26894,N_28220);
or UO_2216 (O_2216,N_29605,N_25307);
xor UO_2217 (O_2217,N_26311,N_29781);
and UO_2218 (O_2218,N_25405,N_25779);
nand UO_2219 (O_2219,N_26001,N_29816);
and UO_2220 (O_2220,N_29814,N_29453);
nor UO_2221 (O_2221,N_28559,N_29876);
nand UO_2222 (O_2222,N_26095,N_29489);
and UO_2223 (O_2223,N_27718,N_27856);
nor UO_2224 (O_2224,N_27767,N_29850);
or UO_2225 (O_2225,N_25794,N_29171);
nor UO_2226 (O_2226,N_29358,N_28333);
nor UO_2227 (O_2227,N_25076,N_29496);
xor UO_2228 (O_2228,N_27480,N_27711);
xnor UO_2229 (O_2229,N_27614,N_28048);
or UO_2230 (O_2230,N_27264,N_28321);
nor UO_2231 (O_2231,N_29412,N_27643);
and UO_2232 (O_2232,N_26388,N_29517);
xnor UO_2233 (O_2233,N_27848,N_25893);
nand UO_2234 (O_2234,N_25910,N_25289);
nand UO_2235 (O_2235,N_27914,N_27556);
or UO_2236 (O_2236,N_26557,N_27210);
xor UO_2237 (O_2237,N_28081,N_27774);
or UO_2238 (O_2238,N_27521,N_26315);
and UO_2239 (O_2239,N_27082,N_28630);
or UO_2240 (O_2240,N_26019,N_27585);
and UO_2241 (O_2241,N_25205,N_29919);
or UO_2242 (O_2242,N_29225,N_27085);
nor UO_2243 (O_2243,N_28702,N_28187);
or UO_2244 (O_2244,N_28134,N_26577);
and UO_2245 (O_2245,N_26551,N_29313);
xnor UO_2246 (O_2246,N_28859,N_26944);
and UO_2247 (O_2247,N_26647,N_27547);
nand UO_2248 (O_2248,N_26401,N_26443);
nand UO_2249 (O_2249,N_28271,N_25223);
and UO_2250 (O_2250,N_27714,N_29020);
nor UO_2251 (O_2251,N_26950,N_29968);
or UO_2252 (O_2252,N_28746,N_25200);
and UO_2253 (O_2253,N_26775,N_28236);
nor UO_2254 (O_2254,N_28509,N_27564);
xor UO_2255 (O_2255,N_29728,N_29592);
and UO_2256 (O_2256,N_27261,N_26885);
xor UO_2257 (O_2257,N_25392,N_25861);
or UO_2258 (O_2258,N_27196,N_28445);
and UO_2259 (O_2259,N_27345,N_27072);
and UO_2260 (O_2260,N_28657,N_27014);
or UO_2261 (O_2261,N_27061,N_28915);
nand UO_2262 (O_2262,N_28049,N_25079);
nor UO_2263 (O_2263,N_28973,N_25659);
nor UO_2264 (O_2264,N_27239,N_25435);
nand UO_2265 (O_2265,N_27299,N_27046);
nand UO_2266 (O_2266,N_25887,N_29067);
and UO_2267 (O_2267,N_28868,N_25879);
or UO_2268 (O_2268,N_29675,N_26656);
xor UO_2269 (O_2269,N_26103,N_28494);
or UO_2270 (O_2270,N_26640,N_29282);
xor UO_2271 (O_2271,N_28359,N_26919);
nand UO_2272 (O_2272,N_27531,N_26914);
and UO_2273 (O_2273,N_27694,N_25267);
nand UO_2274 (O_2274,N_27038,N_29759);
or UO_2275 (O_2275,N_29840,N_25441);
nor UO_2276 (O_2276,N_29908,N_29638);
nand UO_2277 (O_2277,N_29166,N_25810);
and UO_2278 (O_2278,N_27771,N_27428);
and UO_2279 (O_2279,N_29319,N_28776);
nor UO_2280 (O_2280,N_28063,N_25359);
or UO_2281 (O_2281,N_25045,N_25133);
and UO_2282 (O_2282,N_28514,N_26010);
and UO_2283 (O_2283,N_27268,N_28135);
xnor UO_2284 (O_2284,N_27267,N_29448);
nor UO_2285 (O_2285,N_27247,N_28391);
and UO_2286 (O_2286,N_27785,N_27464);
or UO_2287 (O_2287,N_28338,N_27746);
nor UO_2288 (O_2288,N_26541,N_27481);
or UO_2289 (O_2289,N_26643,N_26654);
nor UO_2290 (O_2290,N_28482,N_25155);
nor UO_2291 (O_2291,N_27397,N_28660);
and UO_2292 (O_2292,N_27677,N_26430);
and UO_2293 (O_2293,N_28456,N_27999);
and UO_2294 (O_2294,N_29955,N_26351);
and UO_2295 (O_2295,N_26496,N_27252);
or UO_2296 (O_2296,N_25115,N_25451);
nor UO_2297 (O_2297,N_25623,N_27419);
nand UO_2298 (O_2298,N_29385,N_25847);
nor UO_2299 (O_2299,N_26006,N_25854);
or UO_2300 (O_2300,N_27265,N_28212);
and UO_2301 (O_2301,N_25298,N_25709);
or UO_2302 (O_2302,N_26938,N_29994);
or UO_2303 (O_2303,N_28891,N_25937);
xnor UO_2304 (O_2304,N_28894,N_27276);
xor UO_2305 (O_2305,N_27204,N_26285);
nor UO_2306 (O_2306,N_26065,N_27118);
or UO_2307 (O_2307,N_28222,N_25438);
xnor UO_2308 (O_2308,N_28450,N_29307);
or UO_2309 (O_2309,N_26900,N_28368);
or UO_2310 (O_2310,N_26489,N_25941);
or UO_2311 (O_2311,N_28219,N_29140);
and UO_2312 (O_2312,N_28836,N_29131);
and UO_2313 (O_2313,N_26081,N_29309);
or UO_2314 (O_2314,N_25171,N_26208);
nand UO_2315 (O_2315,N_25936,N_28356);
or UO_2316 (O_2316,N_25122,N_28943);
nor UO_2317 (O_2317,N_26817,N_26432);
nor UO_2318 (O_2318,N_27385,N_29251);
nor UO_2319 (O_2319,N_25539,N_29624);
and UO_2320 (O_2320,N_28697,N_27548);
or UO_2321 (O_2321,N_25407,N_26141);
nor UO_2322 (O_2322,N_28174,N_28952);
and UO_2323 (O_2323,N_26060,N_29750);
or UO_2324 (O_2324,N_28030,N_29410);
and UO_2325 (O_2325,N_25992,N_29771);
nand UO_2326 (O_2326,N_27060,N_28099);
and UO_2327 (O_2327,N_29026,N_25728);
or UO_2328 (O_2328,N_25102,N_26182);
or UO_2329 (O_2329,N_25139,N_28865);
nor UO_2330 (O_2330,N_26270,N_28735);
and UO_2331 (O_2331,N_27438,N_26547);
nand UO_2332 (O_2332,N_27768,N_29708);
nor UO_2333 (O_2333,N_25387,N_28615);
or UO_2334 (O_2334,N_29266,N_25261);
and UO_2335 (O_2335,N_29001,N_28592);
nor UO_2336 (O_2336,N_25255,N_26278);
xor UO_2337 (O_2337,N_26253,N_25367);
and UO_2338 (O_2338,N_25772,N_25120);
nor UO_2339 (O_2339,N_28441,N_26504);
nand UO_2340 (O_2340,N_25973,N_28353);
nand UO_2341 (O_2341,N_29790,N_29300);
or UO_2342 (O_2342,N_28307,N_27529);
nand UO_2343 (O_2343,N_28216,N_26483);
or UO_2344 (O_2344,N_28139,N_26782);
xor UO_2345 (O_2345,N_26968,N_28496);
nand UO_2346 (O_2346,N_28235,N_28162);
nand UO_2347 (O_2347,N_28398,N_29371);
nand UO_2348 (O_2348,N_27006,N_28901);
xor UO_2349 (O_2349,N_26396,N_26889);
nand UO_2350 (O_2350,N_28477,N_27266);
or UO_2351 (O_2351,N_29738,N_29386);
nand UO_2352 (O_2352,N_26793,N_28241);
nand UO_2353 (O_2353,N_25466,N_28104);
nand UO_2354 (O_2354,N_25393,N_26188);
nor UO_2355 (O_2355,N_29486,N_25555);
nor UO_2356 (O_2356,N_29752,N_29287);
and UO_2357 (O_2357,N_26831,N_26486);
or UO_2358 (O_2358,N_29213,N_28619);
or UO_2359 (O_2359,N_29207,N_25119);
and UO_2360 (O_2360,N_26385,N_29743);
xor UO_2361 (O_2361,N_29084,N_29237);
nor UO_2362 (O_2362,N_25231,N_27207);
and UO_2363 (O_2363,N_27962,N_28820);
nor UO_2364 (O_2364,N_25835,N_26067);
nor UO_2365 (O_2365,N_28538,N_28849);
nand UO_2366 (O_2366,N_27703,N_27318);
or UO_2367 (O_2367,N_27324,N_25637);
or UO_2368 (O_2368,N_28427,N_26637);
nand UO_2369 (O_2369,N_29962,N_25958);
and UO_2370 (O_2370,N_28200,N_26424);
and UO_2371 (O_2371,N_25675,N_25749);
and UO_2372 (O_2372,N_26796,N_28457);
or UO_2373 (O_2373,N_27662,N_25570);
and UO_2374 (O_2374,N_28343,N_28130);
or UO_2375 (O_2375,N_26543,N_25271);
nand UO_2376 (O_2376,N_27336,N_26605);
nor UO_2377 (O_2377,N_29834,N_25181);
nor UO_2378 (O_2378,N_25037,N_28917);
nor UO_2379 (O_2379,N_28641,N_28896);
xor UO_2380 (O_2380,N_29177,N_25565);
nor UO_2381 (O_2381,N_29707,N_27744);
and UO_2382 (O_2382,N_29705,N_29074);
and UO_2383 (O_2383,N_28962,N_28601);
nor UO_2384 (O_2384,N_29264,N_28473);
and UO_2385 (O_2385,N_25795,N_25060);
or UO_2386 (O_2386,N_28980,N_25713);
or UO_2387 (O_2387,N_25645,N_29785);
nor UO_2388 (O_2388,N_26490,N_26580);
or UO_2389 (O_2389,N_29458,N_26630);
nor UO_2390 (O_2390,N_27320,N_29441);
and UO_2391 (O_2391,N_27241,N_28195);
or UO_2392 (O_2392,N_29303,N_25538);
and UO_2393 (O_2393,N_27998,N_25591);
xor UO_2394 (O_2394,N_25488,N_29021);
nand UO_2395 (O_2395,N_25952,N_26523);
nand UO_2396 (O_2396,N_26087,N_26949);
and UO_2397 (O_2397,N_28436,N_25831);
and UO_2398 (O_2398,N_29700,N_26538);
and UO_2399 (O_2399,N_28716,N_28499);
or UO_2400 (O_2400,N_27451,N_26792);
or UO_2401 (O_2401,N_29630,N_26560);
nor UO_2402 (O_2402,N_29574,N_29340);
nand UO_2403 (O_2403,N_26712,N_26939);
nor UO_2404 (O_2404,N_27982,N_29649);
nand UO_2405 (O_2405,N_27098,N_26984);
and UO_2406 (O_2406,N_25329,N_25042);
xor UO_2407 (O_2407,N_27122,N_27028);
nor UO_2408 (O_2408,N_28101,N_25617);
and UO_2409 (O_2409,N_25763,N_29181);
nor UO_2410 (O_2410,N_29982,N_27173);
or UO_2411 (O_2411,N_25136,N_26724);
or UO_2412 (O_2412,N_27519,N_25292);
and UO_2413 (O_2413,N_28155,N_26839);
nor UO_2414 (O_2414,N_28997,N_27926);
and UO_2415 (O_2415,N_25413,N_27895);
nor UO_2416 (O_2416,N_29047,N_28403);
nor UO_2417 (O_2417,N_29672,N_27184);
or UO_2418 (O_2418,N_29405,N_27105);
nand UO_2419 (O_2419,N_27243,N_27035);
nor UO_2420 (O_2420,N_26418,N_26300);
and UO_2421 (O_2421,N_28203,N_27886);
or UO_2422 (O_2422,N_26097,N_27807);
or UO_2423 (O_2423,N_27750,N_26652);
nor UO_2424 (O_2424,N_25163,N_25727);
or UO_2425 (O_2425,N_27971,N_25142);
or UO_2426 (O_2426,N_26932,N_27751);
nor UO_2427 (O_2427,N_29553,N_29375);
xnor UO_2428 (O_2428,N_29690,N_26206);
nor UO_2429 (O_2429,N_25666,N_25062);
nand UO_2430 (O_2430,N_27735,N_28026);
nor UO_2431 (O_2431,N_29658,N_26797);
nor UO_2432 (O_2432,N_28944,N_29535);
or UO_2433 (O_2433,N_28667,N_26098);
nand UO_2434 (O_2434,N_26762,N_28501);
and UO_2435 (O_2435,N_27534,N_25674);
nor UO_2436 (O_2436,N_26367,N_29421);
and UO_2437 (O_2437,N_28783,N_27834);
nand UO_2438 (O_2438,N_29253,N_27248);
or UO_2439 (O_2439,N_27075,N_29232);
and UO_2440 (O_2440,N_28629,N_29015);
nor UO_2441 (O_2441,N_25401,N_25341);
nor UO_2442 (O_2442,N_25445,N_28676);
nor UO_2443 (O_2443,N_28689,N_26257);
xnor UO_2444 (O_2444,N_28428,N_29611);
or UO_2445 (O_2445,N_25314,N_27772);
or UO_2446 (O_2446,N_29039,N_25888);
or UO_2447 (O_2447,N_25649,N_26832);
and UO_2448 (O_2448,N_25898,N_28744);
and UO_2449 (O_2449,N_26124,N_28386);
and UO_2450 (O_2450,N_25955,N_25195);
or UO_2451 (O_2451,N_27969,N_29148);
and UO_2452 (O_2452,N_26988,N_25536);
xnor UO_2453 (O_2453,N_29699,N_29762);
xor UO_2454 (O_2454,N_27795,N_27209);
and UO_2455 (O_2455,N_28478,N_26909);
nand UO_2456 (O_2456,N_28887,N_28651);
nand UO_2457 (O_2457,N_28199,N_26843);
nor UO_2458 (O_2458,N_25161,N_27045);
and UO_2459 (O_2459,N_27274,N_29277);
and UO_2460 (O_2460,N_26908,N_25963);
nor UO_2461 (O_2461,N_25542,N_28779);
xor UO_2462 (O_2462,N_27032,N_26238);
nand UO_2463 (O_2463,N_27205,N_28300);
or UO_2464 (O_2464,N_29295,N_28664);
nand UO_2465 (O_2465,N_26139,N_27596);
nor UO_2466 (O_2466,N_28940,N_26068);
nor UO_2467 (O_2467,N_27560,N_27622);
nor UO_2468 (O_2468,N_26353,N_25029);
nor UO_2469 (O_2469,N_29766,N_29221);
nand UO_2470 (O_2470,N_26358,N_29848);
or UO_2471 (O_2471,N_28172,N_27913);
nand UO_2472 (O_2472,N_29898,N_28192);
nand UO_2473 (O_2473,N_25334,N_25049);
xnor UO_2474 (O_2474,N_25409,N_29451);
nand UO_2475 (O_2475,N_26896,N_29544);
and UO_2476 (O_2476,N_27763,N_27773);
nor UO_2477 (O_2477,N_26965,N_25720);
nor UO_2478 (O_2478,N_27222,N_26151);
nand UO_2479 (O_2479,N_28801,N_28821);
or UO_2480 (O_2480,N_25313,N_29438);
and UO_2481 (O_2481,N_27846,N_25233);
or UO_2482 (O_2482,N_25456,N_25770);
nor UO_2483 (O_2483,N_28742,N_25901);
and UO_2484 (O_2484,N_27479,N_28670);
nor UO_2485 (O_2485,N_25416,N_25829);
and UO_2486 (O_2486,N_25146,N_26077);
or UO_2487 (O_2487,N_29342,N_28673);
xor UO_2488 (O_2488,N_25003,N_29849);
and UO_2489 (O_2489,N_25734,N_29610);
or UO_2490 (O_2490,N_26308,N_25268);
nand UO_2491 (O_2491,N_27197,N_25188);
xnor UO_2492 (O_2492,N_28762,N_28513);
or UO_2493 (O_2493,N_29209,N_28883);
or UO_2494 (O_2494,N_28638,N_29479);
and UO_2495 (O_2495,N_27515,N_26390);
and UO_2496 (O_2496,N_27623,N_29193);
nor UO_2497 (O_2497,N_27341,N_25493);
xor UO_2498 (O_2498,N_29879,N_25353);
and UO_2499 (O_2499,N_27021,N_29621);
nor UO_2500 (O_2500,N_26658,N_27071);
nand UO_2501 (O_2501,N_27630,N_26131);
and UO_2502 (O_2502,N_25835,N_27078);
xnor UO_2503 (O_2503,N_29082,N_29053);
or UO_2504 (O_2504,N_29827,N_25169);
or UO_2505 (O_2505,N_27452,N_27491);
and UO_2506 (O_2506,N_26478,N_25240);
nor UO_2507 (O_2507,N_28747,N_28266);
nand UO_2508 (O_2508,N_26240,N_26954);
nor UO_2509 (O_2509,N_28334,N_27161);
nor UO_2510 (O_2510,N_26420,N_26608);
or UO_2511 (O_2511,N_25046,N_26915);
nor UO_2512 (O_2512,N_28735,N_26834);
nor UO_2513 (O_2513,N_27896,N_28633);
nor UO_2514 (O_2514,N_26284,N_26432);
xor UO_2515 (O_2515,N_27215,N_29567);
and UO_2516 (O_2516,N_28865,N_25612);
and UO_2517 (O_2517,N_25795,N_26405);
nand UO_2518 (O_2518,N_26673,N_29038);
or UO_2519 (O_2519,N_29973,N_26841);
nand UO_2520 (O_2520,N_27222,N_27203);
nand UO_2521 (O_2521,N_26313,N_29197);
or UO_2522 (O_2522,N_28002,N_27378);
nand UO_2523 (O_2523,N_25065,N_26245);
nand UO_2524 (O_2524,N_27092,N_29283);
nor UO_2525 (O_2525,N_25004,N_28649);
nor UO_2526 (O_2526,N_26752,N_26800);
and UO_2527 (O_2527,N_25277,N_29518);
or UO_2528 (O_2528,N_28508,N_27271);
or UO_2529 (O_2529,N_25756,N_27923);
and UO_2530 (O_2530,N_26494,N_25277);
nor UO_2531 (O_2531,N_28627,N_26441);
xnor UO_2532 (O_2532,N_26211,N_27335);
nand UO_2533 (O_2533,N_27055,N_29636);
nand UO_2534 (O_2534,N_28550,N_27479);
and UO_2535 (O_2535,N_27863,N_25440);
or UO_2536 (O_2536,N_26142,N_26932);
or UO_2537 (O_2537,N_25351,N_26986);
nor UO_2538 (O_2538,N_29775,N_27615);
or UO_2539 (O_2539,N_25004,N_28464);
and UO_2540 (O_2540,N_28886,N_28320);
and UO_2541 (O_2541,N_26355,N_26927);
and UO_2542 (O_2542,N_25973,N_27276);
or UO_2543 (O_2543,N_27748,N_28213);
nand UO_2544 (O_2544,N_29168,N_25743);
nand UO_2545 (O_2545,N_26809,N_26408);
nor UO_2546 (O_2546,N_26578,N_26013);
nand UO_2547 (O_2547,N_25384,N_27961);
xor UO_2548 (O_2548,N_27907,N_26946);
nand UO_2549 (O_2549,N_25829,N_27347);
or UO_2550 (O_2550,N_26004,N_25116);
nand UO_2551 (O_2551,N_29336,N_26635);
and UO_2552 (O_2552,N_28740,N_27456);
nor UO_2553 (O_2553,N_29854,N_27702);
and UO_2554 (O_2554,N_28037,N_28350);
nor UO_2555 (O_2555,N_28656,N_26370);
xor UO_2556 (O_2556,N_26284,N_26528);
nand UO_2557 (O_2557,N_26767,N_29395);
or UO_2558 (O_2558,N_26514,N_25338);
and UO_2559 (O_2559,N_25473,N_28314);
or UO_2560 (O_2560,N_25075,N_28903);
nand UO_2561 (O_2561,N_28579,N_29702);
xnor UO_2562 (O_2562,N_28324,N_27826);
nor UO_2563 (O_2563,N_27922,N_25425);
and UO_2564 (O_2564,N_29458,N_27199);
or UO_2565 (O_2565,N_25780,N_28775);
nand UO_2566 (O_2566,N_28408,N_29143);
and UO_2567 (O_2567,N_26455,N_28636);
and UO_2568 (O_2568,N_25984,N_26084);
nand UO_2569 (O_2569,N_29946,N_25675);
nand UO_2570 (O_2570,N_26765,N_25706);
nor UO_2571 (O_2571,N_28082,N_26982);
nand UO_2572 (O_2572,N_29402,N_25624);
xor UO_2573 (O_2573,N_28115,N_26503);
nor UO_2574 (O_2574,N_29110,N_25265);
nand UO_2575 (O_2575,N_28705,N_27158);
nand UO_2576 (O_2576,N_26985,N_28528);
xor UO_2577 (O_2577,N_27037,N_27390);
nor UO_2578 (O_2578,N_27578,N_27663);
xnor UO_2579 (O_2579,N_28633,N_28962);
or UO_2580 (O_2580,N_28649,N_25711);
or UO_2581 (O_2581,N_27323,N_25442);
nand UO_2582 (O_2582,N_26972,N_27620);
and UO_2583 (O_2583,N_29119,N_28549);
or UO_2584 (O_2584,N_28365,N_25017);
xor UO_2585 (O_2585,N_28583,N_28294);
nor UO_2586 (O_2586,N_28114,N_29238);
or UO_2587 (O_2587,N_27495,N_29982);
and UO_2588 (O_2588,N_28379,N_29519);
or UO_2589 (O_2589,N_28307,N_26010);
nand UO_2590 (O_2590,N_29464,N_25776);
xor UO_2591 (O_2591,N_27969,N_29360);
or UO_2592 (O_2592,N_25862,N_26793);
nor UO_2593 (O_2593,N_27551,N_27407);
xnor UO_2594 (O_2594,N_27710,N_27089);
or UO_2595 (O_2595,N_26283,N_29401);
or UO_2596 (O_2596,N_29348,N_29894);
nand UO_2597 (O_2597,N_29232,N_26349);
and UO_2598 (O_2598,N_27416,N_25746);
nand UO_2599 (O_2599,N_29321,N_25918);
or UO_2600 (O_2600,N_26734,N_27090);
nor UO_2601 (O_2601,N_28962,N_25734);
nand UO_2602 (O_2602,N_29414,N_28503);
nor UO_2603 (O_2603,N_27681,N_28578);
nor UO_2604 (O_2604,N_26154,N_27024);
or UO_2605 (O_2605,N_25136,N_29780);
or UO_2606 (O_2606,N_29795,N_29467);
or UO_2607 (O_2607,N_29527,N_28920);
nor UO_2608 (O_2608,N_29657,N_28708);
nor UO_2609 (O_2609,N_25502,N_29617);
or UO_2610 (O_2610,N_25353,N_26515);
nand UO_2611 (O_2611,N_27692,N_25711);
and UO_2612 (O_2612,N_26995,N_27065);
nor UO_2613 (O_2613,N_26343,N_27404);
or UO_2614 (O_2614,N_25751,N_26666);
or UO_2615 (O_2615,N_29714,N_27392);
nand UO_2616 (O_2616,N_28519,N_27754);
nand UO_2617 (O_2617,N_29369,N_26530);
and UO_2618 (O_2618,N_28853,N_28984);
nor UO_2619 (O_2619,N_29263,N_25519);
or UO_2620 (O_2620,N_26743,N_25701);
and UO_2621 (O_2621,N_27235,N_25661);
and UO_2622 (O_2622,N_29950,N_26853);
and UO_2623 (O_2623,N_27245,N_28377);
and UO_2624 (O_2624,N_27025,N_27960);
and UO_2625 (O_2625,N_28436,N_29060);
or UO_2626 (O_2626,N_25995,N_27138);
or UO_2627 (O_2627,N_28133,N_27328);
or UO_2628 (O_2628,N_28374,N_27380);
nand UO_2629 (O_2629,N_25794,N_29341);
nor UO_2630 (O_2630,N_25417,N_26636);
nand UO_2631 (O_2631,N_27000,N_29954);
xnor UO_2632 (O_2632,N_28354,N_27295);
and UO_2633 (O_2633,N_28633,N_25640);
or UO_2634 (O_2634,N_27909,N_25767);
and UO_2635 (O_2635,N_25682,N_25098);
or UO_2636 (O_2636,N_25169,N_27257);
xor UO_2637 (O_2637,N_27284,N_27999);
nor UO_2638 (O_2638,N_29234,N_29134);
xnor UO_2639 (O_2639,N_25777,N_26867);
and UO_2640 (O_2640,N_26461,N_28775);
nand UO_2641 (O_2641,N_27128,N_26510);
or UO_2642 (O_2642,N_29788,N_28363);
and UO_2643 (O_2643,N_29270,N_25115);
and UO_2644 (O_2644,N_27572,N_26270);
nor UO_2645 (O_2645,N_27923,N_25140);
nand UO_2646 (O_2646,N_26276,N_26860);
nand UO_2647 (O_2647,N_27764,N_26586);
nor UO_2648 (O_2648,N_28391,N_26462);
nor UO_2649 (O_2649,N_28793,N_28374);
nor UO_2650 (O_2650,N_27689,N_27463);
and UO_2651 (O_2651,N_27512,N_26591);
and UO_2652 (O_2652,N_29795,N_26604);
and UO_2653 (O_2653,N_28784,N_27633);
and UO_2654 (O_2654,N_26461,N_27018);
nor UO_2655 (O_2655,N_26730,N_26018);
nor UO_2656 (O_2656,N_27574,N_29834);
nor UO_2657 (O_2657,N_26238,N_29211);
and UO_2658 (O_2658,N_27471,N_26612);
or UO_2659 (O_2659,N_26283,N_25727);
nand UO_2660 (O_2660,N_27694,N_25284);
nor UO_2661 (O_2661,N_26972,N_27260);
nor UO_2662 (O_2662,N_26589,N_27651);
or UO_2663 (O_2663,N_28028,N_29150);
nand UO_2664 (O_2664,N_29354,N_28806);
nor UO_2665 (O_2665,N_26500,N_25067);
and UO_2666 (O_2666,N_28933,N_25601);
nand UO_2667 (O_2667,N_26030,N_27985);
xnor UO_2668 (O_2668,N_25007,N_25123);
nor UO_2669 (O_2669,N_26578,N_25523);
nand UO_2670 (O_2670,N_29244,N_27896);
nor UO_2671 (O_2671,N_27681,N_27037);
nand UO_2672 (O_2672,N_27040,N_27731);
and UO_2673 (O_2673,N_29948,N_29100);
or UO_2674 (O_2674,N_25325,N_28709);
or UO_2675 (O_2675,N_27135,N_26856);
and UO_2676 (O_2676,N_26586,N_26047);
nand UO_2677 (O_2677,N_25267,N_27023);
nor UO_2678 (O_2678,N_25041,N_26449);
nor UO_2679 (O_2679,N_26563,N_28081);
and UO_2680 (O_2680,N_29271,N_27791);
nor UO_2681 (O_2681,N_28501,N_28335);
nor UO_2682 (O_2682,N_27209,N_25496);
xnor UO_2683 (O_2683,N_25173,N_25347);
and UO_2684 (O_2684,N_25073,N_29066);
nor UO_2685 (O_2685,N_26560,N_28955);
nor UO_2686 (O_2686,N_28215,N_26242);
nor UO_2687 (O_2687,N_29200,N_27001);
nor UO_2688 (O_2688,N_28930,N_29079);
nor UO_2689 (O_2689,N_25958,N_28033);
nor UO_2690 (O_2690,N_25602,N_27980);
nor UO_2691 (O_2691,N_28229,N_28814);
xor UO_2692 (O_2692,N_29222,N_25703);
nor UO_2693 (O_2693,N_27406,N_29918);
nor UO_2694 (O_2694,N_29789,N_29965);
or UO_2695 (O_2695,N_29244,N_29258);
nand UO_2696 (O_2696,N_27454,N_27896);
and UO_2697 (O_2697,N_26921,N_25356);
or UO_2698 (O_2698,N_25497,N_29032);
xor UO_2699 (O_2699,N_29773,N_27809);
and UO_2700 (O_2700,N_25086,N_29278);
or UO_2701 (O_2701,N_27981,N_28795);
nor UO_2702 (O_2702,N_29746,N_28006);
nand UO_2703 (O_2703,N_28171,N_26517);
or UO_2704 (O_2704,N_26262,N_28498);
or UO_2705 (O_2705,N_25245,N_27258);
nand UO_2706 (O_2706,N_29758,N_28320);
nor UO_2707 (O_2707,N_25948,N_27542);
nand UO_2708 (O_2708,N_28940,N_26908);
nand UO_2709 (O_2709,N_26092,N_25200);
nand UO_2710 (O_2710,N_26773,N_27651);
or UO_2711 (O_2711,N_28748,N_25773);
or UO_2712 (O_2712,N_26516,N_26956);
and UO_2713 (O_2713,N_27285,N_26090);
nand UO_2714 (O_2714,N_28712,N_28598);
nor UO_2715 (O_2715,N_27200,N_27730);
nor UO_2716 (O_2716,N_28609,N_28362);
nor UO_2717 (O_2717,N_28899,N_25307);
nand UO_2718 (O_2718,N_28318,N_27531);
nor UO_2719 (O_2719,N_29262,N_28235);
nand UO_2720 (O_2720,N_26097,N_29322);
and UO_2721 (O_2721,N_25588,N_27965);
nor UO_2722 (O_2722,N_27598,N_28371);
and UO_2723 (O_2723,N_28672,N_26190);
nand UO_2724 (O_2724,N_28289,N_27205);
or UO_2725 (O_2725,N_28562,N_29913);
nand UO_2726 (O_2726,N_28993,N_25921);
or UO_2727 (O_2727,N_28133,N_28367);
or UO_2728 (O_2728,N_25207,N_26563);
or UO_2729 (O_2729,N_25284,N_27957);
or UO_2730 (O_2730,N_28374,N_25154);
nand UO_2731 (O_2731,N_25673,N_28324);
xor UO_2732 (O_2732,N_26170,N_25485);
nand UO_2733 (O_2733,N_28262,N_29395);
nor UO_2734 (O_2734,N_29944,N_27306);
nand UO_2735 (O_2735,N_26742,N_26937);
xnor UO_2736 (O_2736,N_26013,N_28179);
and UO_2737 (O_2737,N_28393,N_25648);
or UO_2738 (O_2738,N_25893,N_27763);
nand UO_2739 (O_2739,N_25622,N_28523);
and UO_2740 (O_2740,N_27405,N_29155);
nand UO_2741 (O_2741,N_29454,N_28119);
and UO_2742 (O_2742,N_26737,N_26929);
nand UO_2743 (O_2743,N_28423,N_27938);
or UO_2744 (O_2744,N_26548,N_25727);
or UO_2745 (O_2745,N_27454,N_29911);
xnor UO_2746 (O_2746,N_26569,N_25470);
nor UO_2747 (O_2747,N_25420,N_28754);
nor UO_2748 (O_2748,N_27589,N_26094);
nor UO_2749 (O_2749,N_28437,N_28356);
xor UO_2750 (O_2750,N_25852,N_26674);
or UO_2751 (O_2751,N_26355,N_28170);
or UO_2752 (O_2752,N_27425,N_27842);
or UO_2753 (O_2753,N_28683,N_26544);
and UO_2754 (O_2754,N_26534,N_26474);
nand UO_2755 (O_2755,N_26319,N_29150);
nor UO_2756 (O_2756,N_27664,N_28358);
or UO_2757 (O_2757,N_25888,N_28523);
nand UO_2758 (O_2758,N_29088,N_29067);
nand UO_2759 (O_2759,N_28666,N_27067);
nor UO_2760 (O_2760,N_28828,N_26728);
nand UO_2761 (O_2761,N_27186,N_26041);
and UO_2762 (O_2762,N_28559,N_28232);
and UO_2763 (O_2763,N_28325,N_26289);
nand UO_2764 (O_2764,N_25803,N_26116);
nand UO_2765 (O_2765,N_25163,N_29329);
nor UO_2766 (O_2766,N_25813,N_29788);
nor UO_2767 (O_2767,N_25917,N_26891);
or UO_2768 (O_2768,N_27541,N_26710);
nor UO_2769 (O_2769,N_28107,N_27815);
nand UO_2770 (O_2770,N_28264,N_29574);
or UO_2771 (O_2771,N_25786,N_29349);
or UO_2772 (O_2772,N_29903,N_26888);
and UO_2773 (O_2773,N_28722,N_25088);
nand UO_2774 (O_2774,N_26907,N_27345);
nand UO_2775 (O_2775,N_25520,N_27453);
and UO_2776 (O_2776,N_29982,N_27544);
and UO_2777 (O_2777,N_27107,N_29845);
and UO_2778 (O_2778,N_27982,N_26208);
and UO_2779 (O_2779,N_26662,N_29287);
and UO_2780 (O_2780,N_26917,N_27613);
nor UO_2781 (O_2781,N_27837,N_26821);
or UO_2782 (O_2782,N_25403,N_26744);
nand UO_2783 (O_2783,N_25485,N_27048);
or UO_2784 (O_2784,N_28469,N_29335);
nand UO_2785 (O_2785,N_25306,N_29209);
nor UO_2786 (O_2786,N_29004,N_26655);
or UO_2787 (O_2787,N_29223,N_25190);
or UO_2788 (O_2788,N_29026,N_27074);
nor UO_2789 (O_2789,N_28496,N_29365);
or UO_2790 (O_2790,N_25264,N_27901);
and UO_2791 (O_2791,N_29453,N_27838);
nor UO_2792 (O_2792,N_28697,N_26211);
and UO_2793 (O_2793,N_25384,N_25431);
and UO_2794 (O_2794,N_29433,N_29295);
or UO_2795 (O_2795,N_27556,N_27459);
nand UO_2796 (O_2796,N_26165,N_29132);
nor UO_2797 (O_2797,N_26964,N_29173);
nor UO_2798 (O_2798,N_28258,N_27080);
xor UO_2799 (O_2799,N_27890,N_27658);
nor UO_2800 (O_2800,N_27174,N_29812);
and UO_2801 (O_2801,N_27632,N_29300);
xor UO_2802 (O_2802,N_28214,N_27859);
xor UO_2803 (O_2803,N_29075,N_26631);
nand UO_2804 (O_2804,N_29761,N_27042);
xnor UO_2805 (O_2805,N_27378,N_26271);
xor UO_2806 (O_2806,N_29770,N_28063);
nand UO_2807 (O_2807,N_28201,N_29960);
nand UO_2808 (O_2808,N_25384,N_25129);
and UO_2809 (O_2809,N_25516,N_29937);
xor UO_2810 (O_2810,N_26084,N_28240);
and UO_2811 (O_2811,N_27784,N_27730);
nor UO_2812 (O_2812,N_29903,N_29247);
nor UO_2813 (O_2813,N_25262,N_27421);
and UO_2814 (O_2814,N_25489,N_29597);
and UO_2815 (O_2815,N_29002,N_25331);
or UO_2816 (O_2816,N_26116,N_28364);
or UO_2817 (O_2817,N_25628,N_27593);
xnor UO_2818 (O_2818,N_25347,N_28692);
nor UO_2819 (O_2819,N_28783,N_25311);
nor UO_2820 (O_2820,N_26834,N_27800);
xnor UO_2821 (O_2821,N_25198,N_29404);
nand UO_2822 (O_2822,N_25266,N_27506);
xnor UO_2823 (O_2823,N_27689,N_28360);
and UO_2824 (O_2824,N_27668,N_28918);
nor UO_2825 (O_2825,N_28796,N_29885);
or UO_2826 (O_2826,N_27766,N_26872);
nand UO_2827 (O_2827,N_28928,N_26324);
nor UO_2828 (O_2828,N_26254,N_25839);
nand UO_2829 (O_2829,N_27829,N_25807);
nand UO_2830 (O_2830,N_27378,N_27808);
or UO_2831 (O_2831,N_29068,N_26163);
or UO_2832 (O_2832,N_27541,N_25052);
xnor UO_2833 (O_2833,N_28105,N_28480);
and UO_2834 (O_2834,N_29743,N_29520);
and UO_2835 (O_2835,N_27047,N_27976);
and UO_2836 (O_2836,N_26253,N_26886);
or UO_2837 (O_2837,N_26770,N_29045);
or UO_2838 (O_2838,N_25956,N_27613);
or UO_2839 (O_2839,N_28146,N_28738);
and UO_2840 (O_2840,N_27137,N_28948);
xnor UO_2841 (O_2841,N_26177,N_26950);
and UO_2842 (O_2842,N_25429,N_29627);
or UO_2843 (O_2843,N_26123,N_25936);
nand UO_2844 (O_2844,N_26952,N_27765);
or UO_2845 (O_2845,N_28438,N_28114);
nand UO_2846 (O_2846,N_26657,N_27450);
nand UO_2847 (O_2847,N_28472,N_27750);
and UO_2848 (O_2848,N_25657,N_26479);
and UO_2849 (O_2849,N_27591,N_25008);
nor UO_2850 (O_2850,N_25232,N_27737);
or UO_2851 (O_2851,N_29150,N_26557);
and UO_2852 (O_2852,N_25951,N_28718);
nand UO_2853 (O_2853,N_25697,N_28574);
nand UO_2854 (O_2854,N_27207,N_28957);
and UO_2855 (O_2855,N_28911,N_29352);
or UO_2856 (O_2856,N_28671,N_26871);
xor UO_2857 (O_2857,N_26322,N_26133);
nand UO_2858 (O_2858,N_25911,N_28940);
and UO_2859 (O_2859,N_29286,N_28069);
nor UO_2860 (O_2860,N_29607,N_27969);
nor UO_2861 (O_2861,N_26655,N_29085);
nand UO_2862 (O_2862,N_29852,N_26727);
or UO_2863 (O_2863,N_27450,N_28802);
nand UO_2864 (O_2864,N_26111,N_26186);
or UO_2865 (O_2865,N_27554,N_28755);
xor UO_2866 (O_2866,N_28648,N_27706);
and UO_2867 (O_2867,N_26224,N_26416);
nor UO_2868 (O_2868,N_25809,N_25673);
nand UO_2869 (O_2869,N_28592,N_28141);
and UO_2870 (O_2870,N_26392,N_28181);
nor UO_2871 (O_2871,N_29091,N_25534);
nor UO_2872 (O_2872,N_29652,N_27351);
nor UO_2873 (O_2873,N_28972,N_27343);
and UO_2874 (O_2874,N_25585,N_29143);
or UO_2875 (O_2875,N_25849,N_28906);
nor UO_2876 (O_2876,N_29479,N_27873);
or UO_2877 (O_2877,N_25182,N_28566);
xnor UO_2878 (O_2878,N_28052,N_29373);
nand UO_2879 (O_2879,N_25291,N_29271);
nor UO_2880 (O_2880,N_25491,N_25108);
nand UO_2881 (O_2881,N_25609,N_26157);
nand UO_2882 (O_2882,N_28765,N_27738);
and UO_2883 (O_2883,N_29384,N_26964);
nand UO_2884 (O_2884,N_27512,N_27090);
nand UO_2885 (O_2885,N_28082,N_26692);
nor UO_2886 (O_2886,N_25985,N_25761);
nand UO_2887 (O_2887,N_28542,N_27705);
nand UO_2888 (O_2888,N_28999,N_28727);
nand UO_2889 (O_2889,N_27199,N_29390);
nor UO_2890 (O_2890,N_25002,N_25929);
and UO_2891 (O_2891,N_27701,N_25030);
nand UO_2892 (O_2892,N_27792,N_26277);
and UO_2893 (O_2893,N_25114,N_27459);
or UO_2894 (O_2894,N_25511,N_25720);
or UO_2895 (O_2895,N_28737,N_25906);
nand UO_2896 (O_2896,N_26310,N_25604);
nand UO_2897 (O_2897,N_27914,N_29503);
or UO_2898 (O_2898,N_27124,N_26528);
nor UO_2899 (O_2899,N_27931,N_29876);
nor UO_2900 (O_2900,N_26075,N_25535);
or UO_2901 (O_2901,N_28075,N_29819);
or UO_2902 (O_2902,N_29709,N_25167);
and UO_2903 (O_2903,N_25367,N_28707);
xor UO_2904 (O_2904,N_26095,N_27942);
nand UO_2905 (O_2905,N_27148,N_26006);
xor UO_2906 (O_2906,N_29948,N_25843);
nand UO_2907 (O_2907,N_25457,N_25026);
nand UO_2908 (O_2908,N_26839,N_26827);
and UO_2909 (O_2909,N_26308,N_27537);
or UO_2910 (O_2910,N_25157,N_28928);
and UO_2911 (O_2911,N_28536,N_28994);
nand UO_2912 (O_2912,N_26262,N_29617);
nor UO_2913 (O_2913,N_28170,N_26627);
nor UO_2914 (O_2914,N_27427,N_28043);
or UO_2915 (O_2915,N_26436,N_25762);
nand UO_2916 (O_2916,N_27092,N_29577);
or UO_2917 (O_2917,N_27514,N_29144);
nand UO_2918 (O_2918,N_27727,N_26050);
and UO_2919 (O_2919,N_26140,N_28747);
nand UO_2920 (O_2920,N_26802,N_29359);
nor UO_2921 (O_2921,N_27385,N_27825);
and UO_2922 (O_2922,N_27622,N_29164);
xor UO_2923 (O_2923,N_26641,N_26470);
nand UO_2924 (O_2924,N_27737,N_27601);
xnor UO_2925 (O_2925,N_29541,N_25369);
and UO_2926 (O_2926,N_27556,N_29707);
nor UO_2927 (O_2927,N_27285,N_29495);
nor UO_2928 (O_2928,N_28067,N_29968);
nor UO_2929 (O_2929,N_28384,N_27264);
xor UO_2930 (O_2930,N_29403,N_27210);
and UO_2931 (O_2931,N_25873,N_27964);
and UO_2932 (O_2932,N_27009,N_25800);
nor UO_2933 (O_2933,N_25744,N_25125);
or UO_2934 (O_2934,N_28861,N_29415);
and UO_2935 (O_2935,N_25252,N_27330);
and UO_2936 (O_2936,N_29742,N_26210);
nand UO_2937 (O_2937,N_29057,N_27976);
or UO_2938 (O_2938,N_26580,N_25702);
nand UO_2939 (O_2939,N_27716,N_27450);
nor UO_2940 (O_2940,N_25226,N_26591);
and UO_2941 (O_2941,N_25000,N_26771);
xor UO_2942 (O_2942,N_26160,N_25526);
nand UO_2943 (O_2943,N_28561,N_26121);
xor UO_2944 (O_2944,N_25294,N_26169);
nor UO_2945 (O_2945,N_27258,N_28253);
xor UO_2946 (O_2946,N_27213,N_28034);
nand UO_2947 (O_2947,N_26568,N_27394);
and UO_2948 (O_2948,N_28435,N_26908);
or UO_2949 (O_2949,N_25884,N_25158);
and UO_2950 (O_2950,N_28161,N_25945);
nor UO_2951 (O_2951,N_25603,N_28232);
nor UO_2952 (O_2952,N_28124,N_25516);
nor UO_2953 (O_2953,N_28621,N_25958);
nor UO_2954 (O_2954,N_28476,N_26433);
and UO_2955 (O_2955,N_29346,N_25491);
nor UO_2956 (O_2956,N_25849,N_27324);
or UO_2957 (O_2957,N_25194,N_27502);
or UO_2958 (O_2958,N_26425,N_28236);
and UO_2959 (O_2959,N_27489,N_29677);
or UO_2960 (O_2960,N_26306,N_28708);
or UO_2961 (O_2961,N_25678,N_29463);
nand UO_2962 (O_2962,N_26693,N_29650);
nand UO_2963 (O_2963,N_26407,N_28279);
nor UO_2964 (O_2964,N_26254,N_25366);
nor UO_2965 (O_2965,N_25311,N_27242);
xnor UO_2966 (O_2966,N_27544,N_25298);
nand UO_2967 (O_2967,N_28975,N_25614);
or UO_2968 (O_2968,N_25573,N_28415);
nand UO_2969 (O_2969,N_28107,N_28878);
xor UO_2970 (O_2970,N_27983,N_25130);
nand UO_2971 (O_2971,N_29399,N_27086);
nor UO_2972 (O_2972,N_26053,N_28204);
and UO_2973 (O_2973,N_25110,N_26187);
and UO_2974 (O_2974,N_29435,N_25599);
xor UO_2975 (O_2975,N_29662,N_28059);
and UO_2976 (O_2976,N_29500,N_25778);
nand UO_2977 (O_2977,N_28184,N_29851);
or UO_2978 (O_2978,N_29257,N_27083);
and UO_2979 (O_2979,N_29751,N_28876);
nand UO_2980 (O_2980,N_25004,N_27649);
or UO_2981 (O_2981,N_25195,N_28225);
nor UO_2982 (O_2982,N_25038,N_25983);
xnor UO_2983 (O_2983,N_28017,N_25355);
or UO_2984 (O_2984,N_28971,N_25275);
or UO_2985 (O_2985,N_29727,N_25632);
and UO_2986 (O_2986,N_25895,N_28403);
or UO_2987 (O_2987,N_28751,N_25141);
nand UO_2988 (O_2988,N_25961,N_25874);
and UO_2989 (O_2989,N_29426,N_27969);
nor UO_2990 (O_2990,N_25169,N_25883);
and UO_2991 (O_2991,N_28444,N_26876);
xor UO_2992 (O_2992,N_28214,N_26598);
or UO_2993 (O_2993,N_28081,N_27108);
or UO_2994 (O_2994,N_28160,N_27716);
and UO_2995 (O_2995,N_25753,N_25108);
or UO_2996 (O_2996,N_26789,N_25960);
and UO_2997 (O_2997,N_29588,N_27279);
or UO_2998 (O_2998,N_26236,N_25956);
xor UO_2999 (O_2999,N_29049,N_26051);
xnor UO_3000 (O_3000,N_25370,N_28877);
or UO_3001 (O_3001,N_27979,N_26032);
or UO_3002 (O_3002,N_28605,N_28002);
xnor UO_3003 (O_3003,N_25311,N_26023);
nand UO_3004 (O_3004,N_26767,N_25793);
nor UO_3005 (O_3005,N_28803,N_25438);
nor UO_3006 (O_3006,N_25537,N_29508);
nor UO_3007 (O_3007,N_29784,N_28966);
or UO_3008 (O_3008,N_26808,N_27156);
or UO_3009 (O_3009,N_28352,N_25077);
nand UO_3010 (O_3010,N_28227,N_25166);
and UO_3011 (O_3011,N_25618,N_28536);
or UO_3012 (O_3012,N_28863,N_25821);
or UO_3013 (O_3013,N_28518,N_26598);
or UO_3014 (O_3014,N_28166,N_26840);
nor UO_3015 (O_3015,N_26537,N_29794);
nand UO_3016 (O_3016,N_25166,N_28938);
nor UO_3017 (O_3017,N_26761,N_25877);
xnor UO_3018 (O_3018,N_26380,N_26692);
and UO_3019 (O_3019,N_27770,N_28782);
xnor UO_3020 (O_3020,N_28254,N_28539);
nand UO_3021 (O_3021,N_27902,N_29478);
nor UO_3022 (O_3022,N_27902,N_29134);
or UO_3023 (O_3023,N_25196,N_28295);
nor UO_3024 (O_3024,N_29434,N_25270);
xor UO_3025 (O_3025,N_27554,N_25634);
nor UO_3026 (O_3026,N_26832,N_28914);
nand UO_3027 (O_3027,N_26788,N_28540);
and UO_3028 (O_3028,N_29086,N_27036);
or UO_3029 (O_3029,N_27482,N_25081);
nand UO_3030 (O_3030,N_26655,N_29973);
and UO_3031 (O_3031,N_25744,N_28417);
or UO_3032 (O_3032,N_27379,N_28187);
xnor UO_3033 (O_3033,N_25581,N_29841);
or UO_3034 (O_3034,N_26763,N_27809);
and UO_3035 (O_3035,N_25881,N_25278);
and UO_3036 (O_3036,N_25627,N_29965);
nand UO_3037 (O_3037,N_27617,N_28504);
or UO_3038 (O_3038,N_29239,N_29502);
or UO_3039 (O_3039,N_25673,N_28678);
or UO_3040 (O_3040,N_25887,N_25680);
nor UO_3041 (O_3041,N_25170,N_25745);
or UO_3042 (O_3042,N_25988,N_27686);
or UO_3043 (O_3043,N_28753,N_26568);
and UO_3044 (O_3044,N_26684,N_27858);
or UO_3045 (O_3045,N_28423,N_25780);
nor UO_3046 (O_3046,N_28559,N_28351);
nand UO_3047 (O_3047,N_28555,N_26318);
or UO_3048 (O_3048,N_27095,N_25732);
or UO_3049 (O_3049,N_25012,N_28954);
nand UO_3050 (O_3050,N_25130,N_25098);
and UO_3051 (O_3051,N_28533,N_26123);
or UO_3052 (O_3052,N_26029,N_29727);
nor UO_3053 (O_3053,N_27416,N_26599);
nor UO_3054 (O_3054,N_27963,N_29838);
or UO_3055 (O_3055,N_26546,N_27796);
nand UO_3056 (O_3056,N_27732,N_26227);
and UO_3057 (O_3057,N_27342,N_29550);
nor UO_3058 (O_3058,N_29578,N_26056);
xor UO_3059 (O_3059,N_29858,N_25596);
nand UO_3060 (O_3060,N_27967,N_27255);
nand UO_3061 (O_3061,N_27083,N_29243);
nor UO_3062 (O_3062,N_29875,N_25085);
or UO_3063 (O_3063,N_25406,N_26584);
and UO_3064 (O_3064,N_29589,N_28615);
or UO_3065 (O_3065,N_26947,N_25236);
and UO_3066 (O_3066,N_27525,N_27164);
nand UO_3067 (O_3067,N_29181,N_26237);
nor UO_3068 (O_3068,N_26890,N_27631);
nand UO_3069 (O_3069,N_29180,N_26933);
nor UO_3070 (O_3070,N_26474,N_26460);
nor UO_3071 (O_3071,N_25010,N_26592);
or UO_3072 (O_3072,N_25557,N_29604);
or UO_3073 (O_3073,N_27252,N_29344);
nor UO_3074 (O_3074,N_26831,N_27167);
and UO_3075 (O_3075,N_26031,N_25408);
nor UO_3076 (O_3076,N_26976,N_25928);
nor UO_3077 (O_3077,N_26220,N_28431);
nand UO_3078 (O_3078,N_28403,N_25724);
nand UO_3079 (O_3079,N_28879,N_29222);
nand UO_3080 (O_3080,N_25818,N_26925);
nor UO_3081 (O_3081,N_26318,N_26270);
nand UO_3082 (O_3082,N_26810,N_26303);
or UO_3083 (O_3083,N_29398,N_29788);
or UO_3084 (O_3084,N_27992,N_27604);
nand UO_3085 (O_3085,N_25323,N_27391);
xnor UO_3086 (O_3086,N_26298,N_25961);
nor UO_3087 (O_3087,N_27941,N_25394);
nor UO_3088 (O_3088,N_25041,N_25119);
xor UO_3089 (O_3089,N_29183,N_27502);
or UO_3090 (O_3090,N_26243,N_25165);
and UO_3091 (O_3091,N_26400,N_29872);
nor UO_3092 (O_3092,N_27318,N_26114);
xnor UO_3093 (O_3093,N_29767,N_27385);
or UO_3094 (O_3094,N_29945,N_26957);
nand UO_3095 (O_3095,N_29329,N_28149);
and UO_3096 (O_3096,N_27264,N_29746);
and UO_3097 (O_3097,N_29894,N_25640);
nor UO_3098 (O_3098,N_28845,N_29913);
and UO_3099 (O_3099,N_25231,N_26496);
and UO_3100 (O_3100,N_25050,N_29448);
xor UO_3101 (O_3101,N_28657,N_27826);
nand UO_3102 (O_3102,N_25547,N_27761);
nor UO_3103 (O_3103,N_27003,N_26669);
and UO_3104 (O_3104,N_28040,N_26044);
nor UO_3105 (O_3105,N_28635,N_29431);
or UO_3106 (O_3106,N_28940,N_29408);
nor UO_3107 (O_3107,N_27247,N_25454);
nor UO_3108 (O_3108,N_29860,N_29613);
and UO_3109 (O_3109,N_27207,N_27333);
nand UO_3110 (O_3110,N_27637,N_27139);
and UO_3111 (O_3111,N_28121,N_28509);
or UO_3112 (O_3112,N_26372,N_26620);
nor UO_3113 (O_3113,N_27720,N_27101);
or UO_3114 (O_3114,N_28929,N_27731);
nand UO_3115 (O_3115,N_25995,N_29201);
or UO_3116 (O_3116,N_25572,N_25161);
xnor UO_3117 (O_3117,N_26274,N_26351);
or UO_3118 (O_3118,N_27110,N_29364);
nor UO_3119 (O_3119,N_27431,N_25683);
nor UO_3120 (O_3120,N_28241,N_29086);
nand UO_3121 (O_3121,N_25731,N_27313);
nand UO_3122 (O_3122,N_28398,N_25496);
and UO_3123 (O_3123,N_29968,N_25072);
and UO_3124 (O_3124,N_29301,N_25028);
and UO_3125 (O_3125,N_27220,N_26416);
nand UO_3126 (O_3126,N_26249,N_25415);
and UO_3127 (O_3127,N_29098,N_28024);
nor UO_3128 (O_3128,N_25762,N_29760);
and UO_3129 (O_3129,N_28992,N_28448);
and UO_3130 (O_3130,N_28234,N_27361);
nor UO_3131 (O_3131,N_26492,N_28022);
nand UO_3132 (O_3132,N_27399,N_25149);
nand UO_3133 (O_3133,N_25579,N_29305);
or UO_3134 (O_3134,N_25314,N_29360);
or UO_3135 (O_3135,N_26165,N_27421);
xor UO_3136 (O_3136,N_26854,N_28729);
xor UO_3137 (O_3137,N_29840,N_28869);
nand UO_3138 (O_3138,N_25617,N_25492);
nand UO_3139 (O_3139,N_27252,N_25566);
or UO_3140 (O_3140,N_27439,N_29415);
nor UO_3141 (O_3141,N_26861,N_29681);
nand UO_3142 (O_3142,N_26654,N_29645);
nor UO_3143 (O_3143,N_25616,N_29864);
xor UO_3144 (O_3144,N_26526,N_25391);
or UO_3145 (O_3145,N_28379,N_25855);
or UO_3146 (O_3146,N_29741,N_25016);
and UO_3147 (O_3147,N_25853,N_28215);
nor UO_3148 (O_3148,N_29312,N_29954);
xnor UO_3149 (O_3149,N_26598,N_29263);
xor UO_3150 (O_3150,N_28212,N_28748);
and UO_3151 (O_3151,N_26716,N_25470);
and UO_3152 (O_3152,N_29087,N_28612);
nor UO_3153 (O_3153,N_27063,N_25472);
xnor UO_3154 (O_3154,N_26869,N_29386);
and UO_3155 (O_3155,N_28792,N_25141);
nand UO_3156 (O_3156,N_25521,N_29738);
nor UO_3157 (O_3157,N_28572,N_26870);
and UO_3158 (O_3158,N_25718,N_28450);
or UO_3159 (O_3159,N_28905,N_26210);
xnor UO_3160 (O_3160,N_29933,N_27340);
nor UO_3161 (O_3161,N_29267,N_28241);
and UO_3162 (O_3162,N_28422,N_27991);
or UO_3163 (O_3163,N_29535,N_26417);
or UO_3164 (O_3164,N_25166,N_26748);
and UO_3165 (O_3165,N_27244,N_25427);
or UO_3166 (O_3166,N_29888,N_29875);
or UO_3167 (O_3167,N_25168,N_26443);
nor UO_3168 (O_3168,N_29758,N_25897);
and UO_3169 (O_3169,N_28364,N_27489);
or UO_3170 (O_3170,N_29168,N_26556);
nand UO_3171 (O_3171,N_25590,N_26917);
nor UO_3172 (O_3172,N_29726,N_26099);
nand UO_3173 (O_3173,N_26561,N_27155);
nand UO_3174 (O_3174,N_28095,N_28087);
nand UO_3175 (O_3175,N_29534,N_25459);
nand UO_3176 (O_3176,N_26745,N_25557);
or UO_3177 (O_3177,N_29461,N_27880);
or UO_3178 (O_3178,N_28007,N_29155);
and UO_3179 (O_3179,N_26794,N_26128);
and UO_3180 (O_3180,N_25836,N_29771);
nand UO_3181 (O_3181,N_27688,N_26304);
nor UO_3182 (O_3182,N_28025,N_27975);
and UO_3183 (O_3183,N_25752,N_29040);
nand UO_3184 (O_3184,N_26247,N_25912);
xnor UO_3185 (O_3185,N_25610,N_25820);
or UO_3186 (O_3186,N_29208,N_29754);
nor UO_3187 (O_3187,N_28776,N_28830);
or UO_3188 (O_3188,N_28102,N_26609);
nor UO_3189 (O_3189,N_26371,N_29166);
or UO_3190 (O_3190,N_27115,N_28038);
nand UO_3191 (O_3191,N_28462,N_27711);
and UO_3192 (O_3192,N_28465,N_28922);
nor UO_3193 (O_3193,N_25483,N_26094);
nor UO_3194 (O_3194,N_25120,N_27058);
nand UO_3195 (O_3195,N_28595,N_26345);
or UO_3196 (O_3196,N_25544,N_26580);
nand UO_3197 (O_3197,N_26212,N_29217);
and UO_3198 (O_3198,N_25106,N_25712);
and UO_3199 (O_3199,N_26839,N_25867);
nand UO_3200 (O_3200,N_29177,N_27996);
xor UO_3201 (O_3201,N_29278,N_26648);
nor UO_3202 (O_3202,N_26563,N_26609);
xor UO_3203 (O_3203,N_29124,N_28321);
nand UO_3204 (O_3204,N_27131,N_27669);
nor UO_3205 (O_3205,N_27114,N_28483);
and UO_3206 (O_3206,N_28426,N_26423);
nand UO_3207 (O_3207,N_25936,N_27878);
nand UO_3208 (O_3208,N_27124,N_29056);
nand UO_3209 (O_3209,N_27299,N_26685);
and UO_3210 (O_3210,N_29145,N_29997);
nor UO_3211 (O_3211,N_28391,N_25235);
nand UO_3212 (O_3212,N_27355,N_28155);
or UO_3213 (O_3213,N_26753,N_26729);
nand UO_3214 (O_3214,N_25915,N_26328);
nor UO_3215 (O_3215,N_28312,N_29328);
nor UO_3216 (O_3216,N_29285,N_25539);
nor UO_3217 (O_3217,N_28910,N_29785);
and UO_3218 (O_3218,N_26422,N_29820);
nand UO_3219 (O_3219,N_27411,N_28885);
nor UO_3220 (O_3220,N_25090,N_26283);
and UO_3221 (O_3221,N_27571,N_27748);
and UO_3222 (O_3222,N_29819,N_25579);
and UO_3223 (O_3223,N_28770,N_29517);
or UO_3224 (O_3224,N_28615,N_26468);
and UO_3225 (O_3225,N_29823,N_28992);
nand UO_3226 (O_3226,N_27326,N_26807);
xnor UO_3227 (O_3227,N_27054,N_26903);
and UO_3228 (O_3228,N_29244,N_27328);
or UO_3229 (O_3229,N_26951,N_26583);
nand UO_3230 (O_3230,N_25228,N_26674);
nand UO_3231 (O_3231,N_27388,N_27506);
and UO_3232 (O_3232,N_25888,N_29991);
nand UO_3233 (O_3233,N_29329,N_28953);
nor UO_3234 (O_3234,N_28916,N_27046);
nor UO_3235 (O_3235,N_28224,N_26888);
and UO_3236 (O_3236,N_25928,N_26424);
nor UO_3237 (O_3237,N_26349,N_29074);
xor UO_3238 (O_3238,N_25792,N_25494);
and UO_3239 (O_3239,N_29857,N_26948);
and UO_3240 (O_3240,N_27380,N_28988);
or UO_3241 (O_3241,N_26807,N_29985);
and UO_3242 (O_3242,N_28177,N_28849);
xor UO_3243 (O_3243,N_26127,N_29780);
nand UO_3244 (O_3244,N_26147,N_28232);
nor UO_3245 (O_3245,N_26484,N_27250);
and UO_3246 (O_3246,N_27236,N_26880);
nor UO_3247 (O_3247,N_26164,N_25838);
and UO_3248 (O_3248,N_29267,N_26573);
nand UO_3249 (O_3249,N_26195,N_25353);
nor UO_3250 (O_3250,N_27228,N_25754);
xor UO_3251 (O_3251,N_27750,N_25886);
nand UO_3252 (O_3252,N_28324,N_28762);
nor UO_3253 (O_3253,N_25360,N_28843);
and UO_3254 (O_3254,N_27343,N_25501);
nand UO_3255 (O_3255,N_25816,N_28443);
and UO_3256 (O_3256,N_29270,N_25716);
and UO_3257 (O_3257,N_28261,N_29304);
nand UO_3258 (O_3258,N_28107,N_25739);
nand UO_3259 (O_3259,N_26375,N_27667);
and UO_3260 (O_3260,N_29430,N_28587);
or UO_3261 (O_3261,N_25401,N_28382);
and UO_3262 (O_3262,N_25323,N_25293);
and UO_3263 (O_3263,N_26092,N_26381);
and UO_3264 (O_3264,N_28052,N_27604);
or UO_3265 (O_3265,N_27364,N_26989);
or UO_3266 (O_3266,N_28612,N_27745);
nand UO_3267 (O_3267,N_25999,N_26322);
or UO_3268 (O_3268,N_26944,N_25910);
or UO_3269 (O_3269,N_29369,N_25977);
nand UO_3270 (O_3270,N_26079,N_25017);
and UO_3271 (O_3271,N_25803,N_26148);
and UO_3272 (O_3272,N_29178,N_28363);
nand UO_3273 (O_3273,N_26292,N_26529);
or UO_3274 (O_3274,N_27290,N_27517);
and UO_3275 (O_3275,N_25857,N_26197);
and UO_3276 (O_3276,N_26658,N_29917);
and UO_3277 (O_3277,N_27330,N_26554);
nor UO_3278 (O_3278,N_27224,N_26078);
and UO_3279 (O_3279,N_25525,N_29177);
nand UO_3280 (O_3280,N_27191,N_27344);
and UO_3281 (O_3281,N_25309,N_26548);
or UO_3282 (O_3282,N_27144,N_28936);
and UO_3283 (O_3283,N_29591,N_25267);
and UO_3284 (O_3284,N_29467,N_27190);
xnor UO_3285 (O_3285,N_26684,N_27568);
nand UO_3286 (O_3286,N_25102,N_26977);
and UO_3287 (O_3287,N_26426,N_26645);
nand UO_3288 (O_3288,N_25113,N_29695);
nand UO_3289 (O_3289,N_26166,N_26861);
and UO_3290 (O_3290,N_29432,N_27177);
or UO_3291 (O_3291,N_29082,N_25948);
nand UO_3292 (O_3292,N_26510,N_28353);
nand UO_3293 (O_3293,N_29770,N_29939);
or UO_3294 (O_3294,N_27713,N_28631);
nand UO_3295 (O_3295,N_25561,N_28294);
nand UO_3296 (O_3296,N_25878,N_29121);
or UO_3297 (O_3297,N_25072,N_29856);
or UO_3298 (O_3298,N_28260,N_25960);
nor UO_3299 (O_3299,N_28788,N_27987);
or UO_3300 (O_3300,N_26016,N_27413);
xor UO_3301 (O_3301,N_28590,N_25614);
and UO_3302 (O_3302,N_27118,N_26882);
nand UO_3303 (O_3303,N_26090,N_25590);
nor UO_3304 (O_3304,N_29047,N_27052);
nand UO_3305 (O_3305,N_27625,N_25235);
xnor UO_3306 (O_3306,N_27678,N_28419);
nand UO_3307 (O_3307,N_29412,N_25889);
or UO_3308 (O_3308,N_28427,N_26893);
xor UO_3309 (O_3309,N_28801,N_25609);
or UO_3310 (O_3310,N_29397,N_28624);
nand UO_3311 (O_3311,N_26176,N_25112);
or UO_3312 (O_3312,N_27769,N_29608);
nor UO_3313 (O_3313,N_26637,N_27039);
or UO_3314 (O_3314,N_26133,N_27169);
or UO_3315 (O_3315,N_26391,N_29196);
or UO_3316 (O_3316,N_28401,N_29369);
and UO_3317 (O_3317,N_25955,N_26195);
and UO_3318 (O_3318,N_26007,N_25469);
and UO_3319 (O_3319,N_29681,N_25289);
or UO_3320 (O_3320,N_27418,N_27830);
nand UO_3321 (O_3321,N_26271,N_29476);
nor UO_3322 (O_3322,N_26433,N_26013);
nand UO_3323 (O_3323,N_26418,N_29133);
nor UO_3324 (O_3324,N_27676,N_26235);
or UO_3325 (O_3325,N_29729,N_27888);
and UO_3326 (O_3326,N_28671,N_25691);
nand UO_3327 (O_3327,N_28944,N_26707);
xnor UO_3328 (O_3328,N_29338,N_26003);
nor UO_3329 (O_3329,N_28106,N_26174);
nand UO_3330 (O_3330,N_27154,N_29483);
nand UO_3331 (O_3331,N_29419,N_27684);
or UO_3332 (O_3332,N_26832,N_28161);
or UO_3333 (O_3333,N_29996,N_25206);
and UO_3334 (O_3334,N_29626,N_28430);
and UO_3335 (O_3335,N_26780,N_25155);
and UO_3336 (O_3336,N_25869,N_27858);
or UO_3337 (O_3337,N_29839,N_29951);
nand UO_3338 (O_3338,N_26275,N_29442);
nand UO_3339 (O_3339,N_29574,N_27416);
nand UO_3340 (O_3340,N_29863,N_28370);
or UO_3341 (O_3341,N_29899,N_25165);
and UO_3342 (O_3342,N_29335,N_27573);
nor UO_3343 (O_3343,N_26838,N_28030);
nor UO_3344 (O_3344,N_29438,N_26880);
and UO_3345 (O_3345,N_27513,N_25482);
xnor UO_3346 (O_3346,N_28935,N_29712);
nor UO_3347 (O_3347,N_28984,N_25729);
and UO_3348 (O_3348,N_26259,N_25884);
or UO_3349 (O_3349,N_25923,N_27902);
or UO_3350 (O_3350,N_27786,N_28593);
or UO_3351 (O_3351,N_27668,N_29067);
or UO_3352 (O_3352,N_27041,N_27239);
nand UO_3353 (O_3353,N_29010,N_29909);
xor UO_3354 (O_3354,N_28253,N_25478);
and UO_3355 (O_3355,N_26714,N_26076);
nor UO_3356 (O_3356,N_25460,N_27793);
nand UO_3357 (O_3357,N_29881,N_25902);
nor UO_3358 (O_3358,N_27554,N_26604);
and UO_3359 (O_3359,N_27064,N_28429);
nand UO_3360 (O_3360,N_28836,N_28368);
nand UO_3361 (O_3361,N_26221,N_25870);
nand UO_3362 (O_3362,N_28684,N_25067);
and UO_3363 (O_3363,N_27366,N_26592);
or UO_3364 (O_3364,N_29863,N_26530);
and UO_3365 (O_3365,N_25022,N_26077);
and UO_3366 (O_3366,N_28533,N_28743);
xor UO_3367 (O_3367,N_26964,N_27140);
and UO_3368 (O_3368,N_29460,N_28360);
and UO_3369 (O_3369,N_26642,N_29237);
and UO_3370 (O_3370,N_25999,N_26924);
and UO_3371 (O_3371,N_27955,N_29641);
nand UO_3372 (O_3372,N_28138,N_28098);
nand UO_3373 (O_3373,N_28678,N_25843);
nand UO_3374 (O_3374,N_25726,N_27589);
nand UO_3375 (O_3375,N_27217,N_29166);
xnor UO_3376 (O_3376,N_25535,N_25953);
or UO_3377 (O_3377,N_26302,N_27254);
nand UO_3378 (O_3378,N_26047,N_29157);
xnor UO_3379 (O_3379,N_25592,N_26728);
xor UO_3380 (O_3380,N_28171,N_25728);
and UO_3381 (O_3381,N_27640,N_27079);
nand UO_3382 (O_3382,N_29135,N_26965);
nor UO_3383 (O_3383,N_28939,N_29929);
and UO_3384 (O_3384,N_28586,N_26098);
or UO_3385 (O_3385,N_29691,N_29807);
or UO_3386 (O_3386,N_29054,N_26232);
and UO_3387 (O_3387,N_29000,N_29425);
nand UO_3388 (O_3388,N_29730,N_25959);
nor UO_3389 (O_3389,N_28941,N_28170);
nor UO_3390 (O_3390,N_28791,N_28267);
and UO_3391 (O_3391,N_25648,N_25489);
or UO_3392 (O_3392,N_27158,N_26568);
and UO_3393 (O_3393,N_29117,N_28582);
nor UO_3394 (O_3394,N_26627,N_27469);
nand UO_3395 (O_3395,N_29935,N_29983);
xor UO_3396 (O_3396,N_27935,N_29470);
nand UO_3397 (O_3397,N_25317,N_26097);
nand UO_3398 (O_3398,N_28518,N_26933);
or UO_3399 (O_3399,N_27773,N_29174);
or UO_3400 (O_3400,N_27003,N_27723);
and UO_3401 (O_3401,N_25296,N_28771);
nor UO_3402 (O_3402,N_28012,N_29414);
or UO_3403 (O_3403,N_29864,N_25008);
nand UO_3404 (O_3404,N_25349,N_29174);
and UO_3405 (O_3405,N_26216,N_28351);
or UO_3406 (O_3406,N_28714,N_25764);
nor UO_3407 (O_3407,N_27377,N_25123);
and UO_3408 (O_3408,N_25851,N_28501);
or UO_3409 (O_3409,N_29027,N_29519);
nor UO_3410 (O_3410,N_28122,N_28156);
and UO_3411 (O_3411,N_28927,N_28336);
and UO_3412 (O_3412,N_25504,N_29427);
and UO_3413 (O_3413,N_25015,N_27976);
and UO_3414 (O_3414,N_25500,N_29914);
nand UO_3415 (O_3415,N_28459,N_27852);
nor UO_3416 (O_3416,N_27533,N_29522);
xnor UO_3417 (O_3417,N_26807,N_27764);
nor UO_3418 (O_3418,N_27413,N_29063);
and UO_3419 (O_3419,N_29391,N_28542);
or UO_3420 (O_3420,N_29260,N_25718);
and UO_3421 (O_3421,N_26631,N_28139);
or UO_3422 (O_3422,N_29197,N_26244);
or UO_3423 (O_3423,N_29783,N_27961);
or UO_3424 (O_3424,N_26233,N_27550);
xnor UO_3425 (O_3425,N_27719,N_25173);
nand UO_3426 (O_3426,N_25555,N_27271);
and UO_3427 (O_3427,N_27608,N_28714);
and UO_3428 (O_3428,N_27706,N_27620);
nand UO_3429 (O_3429,N_26634,N_26146);
xor UO_3430 (O_3430,N_29701,N_29391);
nor UO_3431 (O_3431,N_29357,N_29158);
and UO_3432 (O_3432,N_26275,N_28619);
and UO_3433 (O_3433,N_29598,N_28984);
nand UO_3434 (O_3434,N_29054,N_29060);
nor UO_3435 (O_3435,N_28170,N_29353);
nand UO_3436 (O_3436,N_26461,N_25127);
nand UO_3437 (O_3437,N_25415,N_25911);
or UO_3438 (O_3438,N_29969,N_26049);
nand UO_3439 (O_3439,N_26759,N_25777);
or UO_3440 (O_3440,N_26758,N_29055);
xnor UO_3441 (O_3441,N_25818,N_28046);
or UO_3442 (O_3442,N_27656,N_29256);
nor UO_3443 (O_3443,N_27721,N_27618);
or UO_3444 (O_3444,N_25092,N_25284);
nand UO_3445 (O_3445,N_27062,N_26482);
nand UO_3446 (O_3446,N_27640,N_25564);
and UO_3447 (O_3447,N_28271,N_27004);
and UO_3448 (O_3448,N_26601,N_26051);
or UO_3449 (O_3449,N_25724,N_29195);
xnor UO_3450 (O_3450,N_29791,N_29573);
nor UO_3451 (O_3451,N_27586,N_29245);
nand UO_3452 (O_3452,N_26331,N_27007);
and UO_3453 (O_3453,N_28478,N_27194);
nor UO_3454 (O_3454,N_29040,N_28806);
or UO_3455 (O_3455,N_25861,N_29283);
nor UO_3456 (O_3456,N_26058,N_25743);
nand UO_3457 (O_3457,N_27754,N_28960);
or UO_3458 (O_3458,N_26891,N_28696);
or UO_3459 (O_3459,N_29837,N_27817);
nand UO_3460 (O_3460,N_26765,N_29111);
and UO_3461 (O_3461,N_27297,N_29106);
and UO_3462 (O_3462,N_27759,N_25933);
nor UO_3463 (O_3463,N_28193,N_26212);
and UO_3464 (O_3464,N_25588,N_29118);
or UO_3465 (O_3465,N_28512,N_25404);
nor UO_3466 (O_3466,N_29409,N_28868);
nor UO_3467 (O_3467,N_27187,N_26135);
or UO_3468 (O_3468,N_25462,N_27191);
nand UO_3469 (O_3469,N_28216,N_28857);
nand UO_3470 (O_3470,N_26346,N_26156);
and UO_3471 (O_3471,N_27397,N_27962);
nor UO_3472 (O_3472,N_26700,N_28725);
nor UO_3473 (O_3473,N_28221,N_29723);
or UO_3474 (O_3474,N_26787,N_26816);
or UO_3475 (O_3475,N_26576,N_26222);
xnor UO_3476 (O_3476,N_27513,N_25200);
nand UO_3477 (O_3477,N_25050,N_28936);
xnor UO_3478 (O_3478,N_26776,N_29986);
and UO_3479 (O_3479,N_25697,N_28626);
or UO_3480 (O_3480,N_25940,N_28716);
nand UO_3481 (O_3481,N_25197,N_26325);
xnor UO_3482 (O_3482,N_29034,N_26892);
nand UO_3483 (O_3483,N_27988,N_26086);
nor UO_3484 (O_3484,N_29476,N_27561);
nand UO_3485 (O_3485,N_27041,N_28102);
nand UO_3486 (O_3486,N_29368,N_29615);
and UO_3487 (O_3487,N_29248,N_26906);
and UO_3488 (O_3488,N_27083,N_27685);
nand UO_3489 (O_3489,N_27291,N_28187);
nand UO_3490 (O_3490,N_26557,N_26175);
nand UO_3491 (O_3491,N_25614,N_29500);
and UO_3492 (O_3492,N_27645,N_29947);
or UO_3493 (O_3493,N_25595,N_28508);
nand UO_3494 (O_3494,N_28033,N_29426);
nand UO_3495 (O_3495,N_25178,N_29584);
xor UO_3496 (O_3496,N_27189,N_26367);
and UO_3497 (O_3497,N_29141,N_27517);
nor UO_3498 (O_3498,N_26721,N_28847);
and UO_3499 (O_3499,N_25514,N_26898);
endmodule