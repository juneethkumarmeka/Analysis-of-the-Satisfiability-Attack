module basic_2000_20000_2500_4_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_824,In_516);
nand U1 (N_1,In_543,In_1464);
nand U2 (N_2,In_1694,In_836);
nor U3 (N_3,In_754,In_1323);
nor U4 (N_4,In_890,In_581);
or U5 (N_5,In_354,In_613);
and U6 (N_6,In_429,In_1177);
nor U7 (N_7,In_1700,In_1235);
xor U8 (N_8,In_353,In_1359);
or U9 (N_9,In_548,In_1869);
nand U10 (N_10,In_59,In_412);
or U11 (N_11,In_1685,In_1919);
xor U12 (N_12,In_1158,In_1486);
nand U13 (N_13,In_840,In_689);
or U14 (N_14,In_1267,In_1231);
and U15 (N_15,In_1663,In_69);
nor U16 (N_16,In_1073,In_1612);
or U17 (N_17,In_1991,In_1061);
nand U18 (N_18,In_506,In_1266);
nor U19 (N_19,In_1053,In_70);
nor U20 (N_20,In_1760,In_10);
nand U21 (N_21,In_261,In_1664);
and U22 (N_22,In_85,In_787);
nor U23 (N_23,In_1121,In_1480);
and U24 (N_24,In_293,In_1169);
xor U25 (N_25,In_1906,In_515);
and U26 (N_26,In_635,In_1796);
nor U27 (N_27,In_1409,In_327);
nand U28 (N_28,In_956,In_77);
nor U29 (N_29,In_554,In_1490);
and U30 (N_30,In_1154,In_123);
nor U31 (N_31,In_1828,In_1321);
nor U32 (N_32,In_1843,In_1624);
xnor U33 (N_33,In_408,In_1155);
nor U34 (N_34,In_1522,In_1075);
or U35 (N_35,In_1678,In_1008);
nor U36 (N_36,In_99,In_1277);
nor U37 (N_37,In_170,In_1602);
nor U38 (N_38,In_1927,In_111);
xnor U39 (N_39,In_1581,In_181);
xnor U40 (N_40,In_195,In_316);
nor U41 (N_41,In_1866,In_1728);
and U42 (N_42,In_216,In_1106);
nand U43 (N_43,In_1850,In_1093);
nand U44 (N_44,In_1338,In_1912);
and U45 (N_45,In_1199,In_1);
xnor U46 (N_46,In_1766,In_1795);
and U47 (N_47,In_28,In_570);
and U48 (N_48,In_949,In_1576);
or U49 (N_49,In_1201,In_601);
nand U50 (N_50,In_1352,In_1156);
and U51 (N_51,In_1043,In_1849);
xnor U52 (N_52,In_551,In_102);
nor U53 (N_53,In_575,In_1346);
or U54 (N_54,In_1481,In_1249);
nor U55 (N_55,In_419,In_1520);
nand U56 (N_56,In_1269,In_1811);
or U57 (N_57,In_538,In_1608);
nor U58 (N_58,In_1809,In_698);
xnor U59 (N_59,In_1018,In_146);
xnor U60 (N_60,In_734,In_1360);
and U61 (N_61,In_1047,In_12);
nand U62 (N_62,In_1592,In_893);
xnor U63 (N_63,In_1268,In_481);
nor U64 (N_64,In_1897,In_669);
nor U65 (N_65,In_1597,In_1773);
or U66 (N_66,In_376,In_349);
nand U67 (N_67,In_1317,In_631);
nor U68 (N_68,In_1258,In_304);
or U69 (N_69,In_1180,In_1794);
xor U70 (N_70,In_660,In_1119);
xor U71 (N_71,In_873,In_1463);
xnor U72 (N_72,In_646,In_1362);
or U73 (N_73,In_174,In_1288);
nor U74 (N_74,In_121,In_1802);
nand U75 (N_75,In_544,In_112);
or U76 (N_76,In_839,In_550);
nand U77 (N_77,In_64,In_1557);
xnor U78 (N_78,In_1846,In_1752);
nand U79 (N_79,In_1309,In_169);
and U80 (N_80,In_645,In_1790);
and U81 (N_81,In_1250,In_230);
xnor U82 (N_82,In_701,In_866);
xor U83 (N_83,In_396,In_464);
and U84 (N_84,In_943,In_1998);
and U85 (N_85,In_1696,In_571);
nor U86 (N_86,In_1993,In_66);
nor U87 (N_87,In_184,In_572);
nor U88 (N_88,In_1625,In_530);
xor U89 (N_89,In_1152,In_1966);
nor U90 (N_90,In_528,In_517);
and U91 (N_91,In_1675,In_1944);
nor U92 (N_92,In_1071,In_567);
nand U93 (N_93,In_1378,In_1341);
or U94 (N_94,In_1813,In_1764);
nor U95 (N_95,In_1871,In_449);
nor U96 (N_96,In_1745,In_1908);
and U97 (N_97,In_1411,In_876);
nor U98 (N_98,In_724,In_1246);
and U99 (N_99,In_1725,In_1142);
or U100 (N_100,In_1203,In_425);
nor U101 (N_101,In_1689,In_479);
xnor U102 (N_102,In_1916,In_83);
nor U103 (N_103,In_473,In_534);
nand U104 (N_104,In_1355,In_1432);
and U105 (N_105,In_1793,In_1482);
or U106 (N_106,In_510,In_889);
nor U107 (N_107,In_1005,In_305);
and U108 (N_108,In_847,In_302);
and U109 (N_109,In_915,In_526);
and U110 (N_110,In_1070,In_751);
nand U111 (N_111,In_1436,In_225);
xor U112 (N_112,In_206,In_341);
nand U113 (N_113,In_1032,In_1600);
nand U114 (N_114,In_80,In_199);
xor U115 (N_115,In_546,In_1223);
or U116 (N_116,In_332,In_1414);
and U117 (N_117,In_1461,In_1782);
xnor U118 (N_118,In_767,In_829);
xnor U119 (N_119,In_1386,In_1164);
nor U120 (N_120,In_1854,In_1140);
or U121 (N_121,In_124,In_894);
nand U122 (N_122,In_1593,In_1394);
nor U123 (N_123,In_1781,In_553);
and U124 (N_124,In_1303,In_1304);
nand U125 (N_125,In_108,In_1336);
nor U126 (N_126,In_311,In_1650);
xor U127 (N_127,In_1507,In_974);
and U128 (N_128,In_427,In_1619);
and U129 (N_129,In_1589,In_978);
and U130 (N_130,In_907,In_1212);
xnor U131 (N_131,In_706,In_746);
xor U132 (N_132,In_278,In_1108);
or U133 (N_133,In_512,In_789);
or U134 (N_134,In_1647,In_79);
xor U135 (N_135,In_979,In_1731);
nand U136 (N_136,In_151,In_397);
xor U137 (N_137,In_229,In_603);
xnor U138 (N_138,In_968,In_1491);
nor U139 (N_139,In_728,In_1380);
and U140 (N_140,In_1639,In_88);
or U141 (N_141,In_1702,In_1353);
xnor U142 (N_142,In_624,In_461);
or U143 (N_143,In_1296,In_2);
xnor U144 (N_144,In_1928,In_511);
nor U145 (N_145,In_1166,In_1974);
nand U146 (N_146,In_450,In_1420);
nor U147 (N_147,In_1995,In_900);
nand U148 (N_148,In_1348,In_1920);
and U149 (N_149,In_75,In_1157);
nand U150 (N_150,In_1738,In_297);
and U151 (N_151,In_1475,In_1613);
xor U152 (N_152,In_1826,In_292);
xnor U153 (N_153,In_171,In_26);
nand U154 (N_154,In_1049,In_1864);
nand U155 (N_155,In_1146,In_606);
nand U156 (N_156,In_704,In_667);
nand U157 (N_157,In_1272,In_1175);
xor U158 (N_158,In_443,In_987);
and U159 (N_159,In_422,In_1935);
or U160 (N_160,In_458,In_492);
and U161 (N_161,In_1068,In_251);
xor U162 (N_162,In_1375,In_1130);
or U163 (N_163,In_1965,In_1237);
and U164 (N_164,In_918,In_1926);
xnor U165 (N_165,In_1544,In_21);
nor U166 (N_166,In_1545,In_13);
nand U167 (N_167,In_1980,In_1948);
and U168 (N_168,In_621,In_1020);
xnor U169 (N_169,In_1743,In_1384);
xor U170 (N_170,In_457,In_472);
xnor U171 (N_171,In_1449,In_735);
and U172 (N_172,In_952,In_1191);
nand U173 (N_173,In_130,In_1945);
nand U174 (N_174,In_1489,In_1076);
xor U175 (N_175,In_1571,In_508);
and U176 (N_176,In_560,In_1095);
and U177 (N_177,In_535,In_1763);
or U178 (N_178,In_557,In_1709);
nor U179 (N_179,In_1501,In_1282);
nor U180 (N_180,In_17,In_127);
xor U181 (N_181,In_793,In_54);
nor U182 (N_182,In_1051,In_1265);
nor U183 (N_183,In_1462,In_1101);
nor U184 (N_184,In_86,In_218);
nor U185 (N_185,In_1295,In_219);
and U186 (N_186,In_394,In_911);
nor U187 (N_187,In_1335,In_1805);
and U188 (N_188,In_315,In_404);
nor U189 (N_189,In_109,In_858);
nand U190 (N_190,In_1783,In_919);
nand U191 (N_191,In_568,In_60);
nand U192 (N_192,In_659,In_330);
and U193 (N_193,In_1657,In_1318);
nor U194 (N_194,In_737,In_355);
xnor U195 (N_195,In_1088,In_810);
xor U196 (N_196,In_175,In_37);
xnor U197 (N_197,In_145,In_1682);
or U198 (N_198,In_1910,In_973);
xnor U199 (N_199,In_1202,In_1455);
or U200 (N_200,In_418,In_1065);
and U201 (N_201,In_1891,In_844);
and U202 (N_202,In_1454,In_616);
or U203 (N_203,In_401,In_191);
nand U204 (N_204,In_1413,In_1280);
and U205 (N_205,In_1220,In_678);
and U206 (N_206,In_869,In_768);
nor U207 (N_207,In_212,In_33);
nand U208 (N_208,In_1055,In_1564);
nand U209 (N_209,In_266,In_1366);
and U210 (N_210,In_1275,In_1390);
xnor U211 (N_211,In_1772,In_947);
nor U212 (N_212,In_1098,In_202);
and U213 (N_213,In_870,In_1844);
xor U214 (N_214,In_1044,In_371);
or U215 (N_215,In_815,In_565);
and U216 (N_216,In_166,In_1084);
nand U217 (N_217,In_778,In_477);
xnor U218 (N_218,In_605,In_1260);
or U219 (N_219,In_1655,In_465);
and U220 (N_220,In_1648,In_1911);
xnor U221 (N_221,In_1285,In_1913);
nand U222 (N_222,In_1753,In_1503);
and U223 (N_223,In_875,In_856);
and U224 (N_224,In_456,In_811);
nor U225 (N_225,In_61,In_1292);
and U226 (N_226,In_322,In_0);
and U227 (N_227,In_1517,In_990);
nand U228 (N_228,In_1033,In_1615);
nor U229 (N_229,In_298,In_1063);
nor U230 (N_230,In_280,In_154);
xnor U231 (N_231,In_967,In_1604);
nand U232 (N_232,In_1845,In_561);
nand U233 (N_233,In_1858,In_1601);
and U234 (N_234,In_1889,In_756);
nand U235 (N_235,In_361,In_1046);
nor U236 (N_236,In_1392,In_597);
xnor U237 (N_237,In_682,In_1162);
nor U238 (N_238,In_541,In_1042);
xor U239 (N_239,In_1984,In_393);
nand U240 (N_240,In_806,In_1931);
or U241 (N_241,In_932,In_1479);
or U242 (N_242,In_825,In_708);
and U243 (N_243,In_373,In_1968);
xor U244 (N_244,In_1695,In_91);
and U245 (N_245,In_1208,In_1458);
xnor U246 (N_246,In_276,In_820);
or U247 (N_247,In_785,In_309);
and U248 (N_248,In_1013,In_281);
nand U249 (N_249,In_14,In_177);
nand U250 (N_250,In_435,In_1374);
and U251 (N_251,In_1930,In_1605);
or U252 (N_252,In_1372,In_854);
and U253 (N_253,In_470,In_743);
or U254 (N_254,In_1182,In_1456);
or U255 (N_255,In_1561,In_1582);
and U256 (N_256,In_1830,In_1936);
nor U257 (N_257,In_874,In_685);
nor U258 (N_258,In_236,In_922);
or U259 (N_259,In_863,In_1532);
nor U260 (N_260,In_1111,In_1184);
nor U261 (N_261,In_1219,In_1734);
xor U262 (N_262,In_861,In_755);
xor U263 (N_263,In_582,In_49);
xor U264 (N_264,In_58,In_447);
xnor U265 (N_265,In_849,In_1918);
or U266 (N_266,In_1497,In_1513);
or U267 (N_267,In_938,In_1179);
or U268 (N_268,In_1504,In_45);
and U269 (N_269,In_1389,In_929);
and U270 (N_270,In_770,In_1801);
nand U271 (N_271,In_1131,In_1502);
nand U272 (N_272,In_409,In_248);
and U273 (N_273,In_1787,In_804);
and U274 (N_274,In_326,In_1450);
nor U275 (N_275,In_1129,In_1746);
nand U276 (N_276,In_1314,In_1769);
nor U277 (N_277,In_1284,In_1777);
nand U278 (N_278,In_1149,In_1778);
and U279 (N_279,In_1609,In_1631);
xor U280 (N_280,In_116,In_986);
nor U281 (N_281,In_1026,In_1165);
nor U282 (N_282,In_1797,In_1658);
and U283 (N_283,In_1344,In_686);
and U284 (N_284,In_344,In_1634);
nor U285 (N_285,In_204,In_1232);
nor U286 (N_286,In_1057,In_740);
nand U287 (N_287,In_389,In_1468);
or U288 (N_288,In_617,In_1122);
or U289 (N_289,In_395,In_431);
nor U290 (N_290,In_24,In_579);
nor U291 (N_291,In_1147,In_558);
nor U292 (N_292,In_1859,In_1880);
or U293 (N_293,In_1933,In_1672);
xor U294 (N_294,In_365,In_1216);
xor U295 (N_295,In_289,In_463);
xnor U296 (N_296,In_730,In_381);
nor U297 (N_297,In_1459,In_415);
or U298 (N_298,In_1553,In_370);
xor U299 (N_299,In_1904,In_1153);
nor U300 (N_300,In_279,In_1319);
nand U301 (N_301,In_329,In_1516);
nand U302 (N_302,In_1874,In_805);
or U303 (N_303,In_1656,In_1437);
xnor U304 (N_304,In_103,In_1325);
nor U305 (N_305,In_1270,In_823);
xnor U306 (N_306,In_1483,In_303);
or U307 (N_307,In_1925,In_954);
nand U308 (N_308,In_1022,In_380);
xnor U309 (N_309,In_52,In_1890);
xnor U310 (N_310,In_1240,In_703);
nor U311 (N_311,In_1442,In_471);
nand U312 (N_312,In_1271,In_1377);
and U313 (N_313,In_1087,In_1835);
xor U314 (N_314,In_1816,In_1465);
xor U315 (N_315,In_1578,In_1855);
and U316 (N_316,In_995,In_1596);
xnor U317 (N_317,In_883,In_1007);
nor U318 (N_318,In_1715,In_194);
or U319 (N_319,In_1640,In_1331);
or U320 (N_320,In_1946,In_139);
nor U321 (N_321,In_76,In_287);
nor U322 (N_322,In_1248,In_1832);
or U323 (N_323,In_1646,In_378);
xor U324 (N_324,In_991,In_1193);
nand U325 (N_325,In_1626,In_1954);
or U326 (N_326,In_1045,In_690);
nand U327 (N_327,In_542,In_67);
and U328 (N_328,In_228,In_827);
nor U329 (N_329,In_50,In_7);
nor U330 (N_330,In_157,In_1397);
nand U331 (N_331,In_934,In_1329);
and U332 (N_332,In_1707,In_343);
nor U333 (N_333,In_1118,In_1126);
xor U334 (N_334,In_1510,In_1173);
and U335 (N_335,In_484,In_273);
and U336 (N_336,In_1718,In_1211);
nor U337 (N_337,In_1580,In_707);
xor U338 (N_338,In_1938,In_417);
nor U339 (N_339,In_673,In_1168);
and U340 (N_340,In_1780,In_140);
xor U341 (N_341,In_242,In_1577);
xor U342 (N_342,In_1429,In_437);
nand U343 (N_343,In_342,In_1873);
xnor U344 (N_344,In_1825,In_999);
nor U345 (N_345,In_306,In_1264);
and U346 (N_346,In_1286,In_1496);
or U347 (N_347,In_519,In_122);
or U348 (N_348,In_446,In_623);
nor U349 (N_349,In_488,In_133);
xnor U350 (N_350,In_1001,In_834);
nand U351 (N_351,In_93,In_566);
nand U352 (N_352,In_587,In_117);
and U353 (N_353,In_747,In_960);
or U354 (N_354,In_1259,In_71);
or U355 (N_355,In_1395,In_359);
xnor U356 (N_356,In_263,In_586);
and U357 (N_357,In_469,In_1358);
nor U358 (N_358,In_1369,In_504);
nand U359 (N_359,In_36,In_1337);
nand U360 (N_360,In_1457,In_1298);
or U361 (N_361,In_1637,In_1294);
xor U362 (N_362,In_1109,In_383);
xnor U363 (N_363,In_310,In_721);
or U364 (N_364,In_1810,In_286);
xor U365 (N_365,In_1900,In_106);
nor U366 (N_366,In_1401,In_763);
or U367 (N_367,In_1607,In_35);
or U368 (N_368,In_822,In_5);
nor U369 (N_369,In_141,In_1159);
nand U370 (N_370,In_764,In_1868);
or U371 (N_371,In_977,In_441);
xor U372 (N_372,In_1009,In_742);
or U373 (N_373,In_972,In_129);
nor U374 (N_374,In_84,In_1107);
and U375 (N_375,In_857,In_902);
or U376 (N_376,In_485,In_1531);
or U377 (N_377,In_738,In_1200);
xnor U378 (N_378,In_607,In_496);
and U379 (N_379,In_1206,In_1528);
xnor U380 (N_380,In_1887,In_1431);
and U381 (N_381,In_975,In_750);
or U382 (N_382,In_1444,In_1840);
or U383 (N_383,In_137,In_1135);
and U384 (N_384,In_351,In_937);
xor U385 (N_385,In_599,In_244);
xor U386 (N_386,In_402,In_1515);
nand U387 (N_387,In_1909,In_1951);
xnor U388 (N_388,In_665,In_160);
xnor U389 (N_389,In_32,In_1127);
and U390 (N_390,In_615,In_1654);
xor U391 (N_391,In_1410,In_1754);
and U392 (N_392,In_1289,In_436);
xor U393 (N_393,In_628,In_4);
xnor U394 (N_394,In_1163,In_1905);
and U395 (N_395,In_120,In_1566);
and U396 (N_396,In_1116,In_1765);
nor U397 (N_397,In_283,In_1603);
or U398 (N_398,In_1080,In_240);
nand U399 (N_399,In_830,In_769);
nor U400 (N_400,In_209,In_549);
nor U401 (N_401,In_1004,In_537);
and U402 (N_402,In_1803,In_105);
nor U403 (N_403,In_705,In_1804);
xor U404 (N_404,In_399,In_1623);
and U405 (N_405,In_468,In_1960);
or U406 (N_406,In_1245,In_913);
and U407 (N_407,In_1328,In_1824);
or U408 (N_408,In_1565,In_150);
xor U409 (N_409,In_899,In_1856);
or U410 (N_410,In_1614,In_11);
or U411 (N_411,In_656,In_1412);
nand U412 (N_412,In_520,In_1870);
xnor U413 (N_413,In_403,In_1396);
and U414 (N_414,In_803,In_357);
nand U415 (N_415,In_1537,In_1676);
nor U416 (N_416,In_585,In_1030);
or U417 (N_417,In_497,In_927);
and U418 (N_418,In_1083,In_1536);
nand U419 (N_419,In_998,In_720);
or U420 (N_420,In_752,In_1027);
or U421 (N_421,In_580,In_82);
xnor U422 (N_422,In_483,In_110);
nand U423 (N_423,In_906,In_259);
and U424 (N_424,In_1784,In_1741);
xnor U425 (N_425,In_267,In_1276);
and U426 (N_426,In_254,In_1957);
or U427 (N_427,In_1722,In_848);
or U428 (N_428,In_333,In_1590);
or U429 (N_429,In_1956,In_176);
or U430 (N_430,In_1750,In_1067);
or U431 (N_431,In_749,In_1148);
nand U432 (N_432,In_649,In_564);
or U433 (N_433,In_925,In_1453);
or U434 (N_434,In_1899,In_1755);
and U435 (N_435,In_984,In_608);
and U436 (N_436,In_486,In_1903);
and U437 (N_437,In_914,In_159);
nand U438 (N_438,In_1661,In_1751);
xor U439 (N_439,In_997,In_1633);
or U440 (N_440,In_636,In_1985);
nor U441 (N_441,In_1031,In_1535);
nor U442 (N_442,In_1171,In_1440);
and U443 (N_443,In_48,In_1040);
nor U444 (N_444,In_814,In_1981);
and U445 (N_445,In_1990,In_731);
xor U446 (N_446,In_1241,In_247);
nand U447 (N_447,In_38,In_1560);
and U448 (N_448,In_723,In_1761);
or U449 (N_449,In_1921,In_648);
or U450 (N_450,In_1299,In_777);
and U451 (N_451,In_1688,In_148);
and U452 (N_452,In_655,In_459);
nand U453 (N_453,In_319,In_1406);
nand U454 (N_454,In_503,In_1999);
and U455 (N_455,In_1519,In_732);
or U456 (N_456,In_233,In_620);
nor U457 (N_457,In_879,In_1572);
nor U458 (N_458,In_1417,In_1419);
nand U459 (N_459,In_1779,In_523);
and U460 (N_460,In_766,In_1708);
and U461 (N_461,In_107,In_813);
or U462 (N_462,In_43,In_100);
nor U463 (N_463,In_595,In_779);
nand U464 (N_464,In_220,In_197);
and U465 (N_465,In_1518,In_165);
nand U466 (N_466,In_596,In_475);
or U467 (N_467,In_424,In_715);
and U468 (N_468,In_434,In_1651);
or U469 (N_469,In_308,In_982);
and U470 (N_470,In_727,In_1469);
nor U471 (N_471,In_1878,In_518);
nand U472 (N_472,In_1224,In_501);
nand U473 (N_473,In_290,In_1478);
xor U474 (N_474,In_1842,In_1788);
xnor U475 (N_475,In_1949,In_56);
or U476 (N_476,In_313,In_1808);
nand U477 (N_477,In_94,In_187);
xnor U478 (N_478,In_1205,In_363);
nor U479 (N_479,In_1740,In_1922);
and U480 (N_480,In_1703,In_1243);
or U481 (N_481,In_950,In_1196);
or U482 (N_482,In_612,In_135);
xnor U483 (N_483,In_946,In_1941);
nor U484 (N_484,In_772,In_1029);
nor U485 (N_485,In_1534,In_1059);
or U486 (N_486,In_1666,In_98);
or U487 (N_487,In_1915,In_1895);
xor U488 (N_488,In_411,In_1244);
nor U489 (N_489,In_589,In_1218);
nor U490 (N_490,In_22,In_23);
xnor U491 (N_491,In_1161,In_1770);
or U492 (N_492,In_590,In_808);
xnor U493 (N_493,In_1014,In_161);
xor U494 (N_494,In_1143,In_1262);
nor U495 (N_495,In_92,In_299);
nor U496 (N_496,In_657,In_153);
or U497 (N_497,In_800,In_338);
or U498 (N_498,In_324,In_1434);
nand U499 (N_499,In_1423,In_1133);
nand U500 (N_500,In_993,In_1879);
or U501 (N_501,In_563,In_905);
nor U502 (N_502,In_1310,In_1812);
or U503 (N_503,In_574,In_1807);
xnor U504 (N_504,In_182,In_1167);
or U505 (N_505,In_1144,In_1025);
xor U506 (N_506,In_224,In_881);
and U507 (N_507,In_350,In_152);
nor U508 (N_508,In_1488,In_862);
nand U509 (N_509,In_474,In_430);
nand U510 (N_510,In_1428,In_27);
and U511 (N_511,In_1333,In_916);
nor U512 (N_512,In_521,In_936);
nor U513 (N_513,In_1800,In_630);
xnor U514 (N_514,In_51,In_256);
or U515 (N_515,In_666,In_300);
or U516 (N_516,In_1762,In_681);
nand U517 (N_517,In_1509,In_909);
and U518 (N_518,In_795,In_545);
and U519 (N_519,In_578,In_134);
xnor U520 (N_520,In_1701,In_958);
xnor U521 (N_521,In_1884,In_1717);
or U522 (N_522,In_1829,In_1052);
and U523 (N_523,In_1388,In_1552);
xnor U524 (N_524,In_1729,In_833);
xnor U525 (N_525,In_1587,In_692);
and U526 (N_526,In_1710,In_807);
or U527 (N_527,In_442,In_1239);
and U528 (N_528,In_1069,In_1028);
xor U529 (N_529,In_794,In_339);
and U530 (N_530,In_1422,In_1247);
nand U531 (N_531,In_1881,In_1799);
xor U532 (N_532,In_1791,In_183);
xnor U533 (N_533,In_1050,In_257);
nand U534 (N_534,In_1591,In_1937);
nor U535 (N_535,In_1892,In_725);
xor U536 (N_536,In_864,In_356);
nand U537 (N_537,In_1575,In_444);
xnor U538 (N_538,In_1361,In_1399);
or U539 (N_539,In_654,In_239);
xor U540 (N_540,In_697,In_72);
or U541 (N_541,In_696,In_691);
or U542 (N_542,In_1542,In_19);
nand U543 (N_543,In_375,In_1064);
or U544 (N_544,In_1848,In_158);
or U545 (N_545,In_658,In_1477);
xor U546 (N_546,In_1533,In_1283);
nor U547 (N_547,In_1190,In_1967);
and U548 (N_548,In_963,In_1992);
or U549 (N_549,In_726,In_1556);
and U550 (N_550,In_143,In_1445);
xnor U551 (N_551,In_235,In_1228);
and U552 (N_552,In_562,In_1447);
nand U553 (N_553,In_671,In_34);
nand U554 (N_554,In_957,In_799);
nand U555 (N_555,In_367,In_1441);
xor U556 (N_556,In_895,In_260);
or U557 (N_557,In_253,In_1253);
or U558 (N_558,In_1767,In_1588);
nor U559 (N_559,In_221,In_1186);
or U560 (N_560,In_1234,In_629);
xnor U561 (N_561,In_1425,In_1495);
nand U562 (N_562,In_1817,In_641);
and U563 (N_563,In_495,In_1089);
nor U564 (N_564,In_1671,In_1546);
nor U565 (N_565,In_1823,In_1302);
xor U566 (N_566,In_489,In_368);
nand U567 (N_567,In_275,In_1291);
nand U568 (N_568,In_201,In_452);
or U569 (N_569,In_1543,In_20);
nor U570 (N_570,In_1103,In_901);
nand U571 (N_571,In_372,In_672);
and U572 (N_572,In_1078,In_232);
nand U573 (N_573,In_1630,In_1100);
or U574 (N_574,In_416,In_1617);
nor U575 (N_575,In_1538,In_1301);
and U576 (N_576,In_1659,In_1350);
or U577 (N_577,In_238,In_759);
or U578 (N_578,In_817,In_42);
nor U579 (N_579,In_320,In_234);
or U580 (N_580,In_1215,In_1833);
or U581 (N_581,In_1723,In_73);
nor U582 (N_582,In_700,In_268);
nor U583 (N_583,In_1097,In_1549);
nor U584 (N_584,In_505,In_837);
and U585 (N_585,In_192,In_1508);
nor U586 (N_586,In_1628,In_1641);
or U587 (N_587,In_942,In_414);
xor U588 (N_588,In_1622,In_1227);
or U589 (N_589,In_996,In_1470);
and U590 (N_590,In_1019,In_1120);
nor U591 (N_591,In_325,In_1408);
or U592 (N_592,In_207,In_668);
nor U593 (N_593,In_994,In_1077);
or U594 (N_594,In_1896,In_1901);
and U595 (N_595,In_3,In_1867);
and U596 (N_596,In_637,In_53);
nor U597 (N_597,In_712,In_694);
nor U598 (N_598,In_214,In_1485);
xor U599 (N_599,In_1125,In_989);
and U600 (N_600,In_1499,In_1252);
nor U601 (N_601,In_1102,In_384);
nor U602 (N_602,In_912,In_1929);
nand U603 (N_603,In_262,In_1586);
and U604 (N_604,In_614,In_1616);
xor U605 (N_605,In_265,In_812);
nand U606 (N_606,In_1555,In_1415);
xnor U607 (N_607,In_626,In_843);
and U608 (N_608,In_63,In_971);
or U609 (N_609,In_30,In_1527);
xnor U610 (N_610,In_1851,In_1066);
and U611 (N_611,In_1512,In_198);
xor U612 (N_612,In_1932,In_1368);
nor U613 (N_613,In_1815,In_1987);
nor U614 (N_614,In_1514,In_231);
and U615 (N_615,In_1988,In_1382);
nand U616 (N_616,In_1525,In_935);
nand U617 (N_617,In_1923,In_258);
nor U618 (N_618,In_1105,In_1642);
and U619 (N_619,In_142,In_529);
nand U620 (N_620,In_1838,In_1128);
and U621 (N_621,In_850,In_1506);
xnor U622 (N_622,In_1354,In_284);
and U623 (N_623,In_555,In_1345);
nor U624 (N_624,In_871,In_801);
and U625 (N_625,In_1888,In_1194);
xor U626 (N_626,In_1367,In_1978);
and U627 (N_627,In_790,In_1230);
or U628 (N_628,In_1530,In_930);
nand U629 (N_629,In_1000,In_491);
nand U630 (N_630,In_188,In_1448);
nor U631 (N_631,In_1214,In_227);
and U632 (N_632,In_1724,In_410);
or U633 (N_633,In_1385,In_345);
or U634 (N_634,In_1226,In_1343);
and U635 (N_635,In_101,In_962);
xnor U636 (N_636,In_1583,In_1986);
xnor U637 (N_637,In_1058,In_1673);
xnor U638 (N_638,In_1365,In_291);
xor U639 (N_639,In_1340,In_1238);
and U640 (N_640,In_1732,In_1364);
nor U641 (N_641,In_1160,In_1821);
nand U642 (N_642,In_1785,In_969);
or U643 (N_643,In_955,In_642);
nand U644 (N_644,In_1559,In_1569);
nor U645 (N_645,In_1024,In_1357);
nand U646 (N_646,In_1726,In_1834);
nor U647 (N_647,In_115,In_178);
xnor U648 (N_648,In_951,In_885);
nor U649 (N_649,In_1023,In_439);
or U650 (N_650,In_1048,In_1652);
or U651 (N_651,In_1339,In_493);
nor U652 (N_652,In_453,In_1421);
or U653 (N_653,In_1606,In_1983);
or U654 (N_654,In_1472,In_1451);
nor U655 (N_655,In_841,In_592);
or U656 (N_656,In_1426,In_1610);
xnor U657 (N_657,In_1471,In_1822);
nor U658 (N_658,In_1839,In_1320);
and U659 (N_659,In_455,In_1550);
or U660 (N_660,In_215,In_1775);
nor U661 (N_661,In_826,In_771);
nor U662 (N_662,In_57,In_882);
nand U663 (N_663,In_786,In_205);
and U664 (N_664,In_1744,In_953);
or U665 (N_665,In_1197,In_360);
xnor U666 (N_666,In_1759,In_638);
and U667 (N_667,In_783,In_200);
or U668 (N_668,In_331,In_640);
nor U669 (N_669,In_312,In_277);
xnor U670 (N_670,In_203,In_1611);
xnor U671 (N_671,In_1706,In_1841);
or U672 (N_672,In_583,In_1112);
nor U673 (N_673,In_1886,In_1308);
or U674 (N_674,In_136,In_1950);
and U675 (N_675,In_1123,In_189);
nand U676 (N_676,In_1670,In_1727);
xnor U677 (N_677,In_1687,In_1698);
and U678 (N_678,In_719,In_651);
nor U679 (N_679,In_536,In_1082);
or U680 (N_680,In_1771,In_522);
and U681 (N_681,In_1595,In_643);
nand U682 (N_682,In_1021,In_377);
nor U683 (N_683,In_924,In_31);
nand U684 (N_684,In_1526,In_944);
xor U685 (N_685,In_167,In_272);
nand U686 (N_686,In_440,In_1847);
nand U687 (N_687,In_210,In_1997);
nand U688 (N_688,In_965,In_1446);
xor U689 (N_689,In_317,In_838);
or U690 (N_690,In_352,In_285);
or U691 (N_691,In_1584,In_1351);
nand U692 (N_692,In_602,In_379);
xor U693 (N_693,In_1885,In_1882);
xnor U694 (N_694,In_413,In_1287);
nor U695 (N_695,In_1883,In_711);
nor U696 (N_696,In_1758,In_765);
or U697 (N_697,In_1629,In_1872);
xor U698 (N_698,In_831,In_168);
or U699 (N_699,In_855,In_97);
or U700 (N_700,In_1907,In_1187);
or U701 (N_701,In_498,In_1964);
nand U702 (N_702,In_423,In_593);
nor U703 (N_703,In_382,In_540);
or U704 (N_704,In_223,In_1213);
nand U705 (N_705,In_1003,In_1940);
nand U706 (N_706,In_886,In_1668);
or U707 (N_707,In_664,In_964);
nand U708 (N_708,In_1902,In_903);
xor U709 (N_709,In_432,In_981);
nand U710 (N_710,In_1104,In_1242);
or U711 (N_711,In_632,In_387);
and U712 (N_712,In_1714,In_125);
nand U713 (N_713,In_41,In_149);
xnor U714 (N_714,In_1136,In_1170);
nand U715 (N_715,In_1523,In_1493);
or U716 (N_716,In_985,In_1554);
xor U717 (N_717,In_1558,In_74);
xor U718 (N_718,In_1861,In_144);
or U719 (N_719,In_702,In_87);
xnor U720 (N_720,In_1099,In_68);
and U721 (N_721,In_832,In_407);
and U722 (N_722,In_741,In_1347);
nand U723 (N_723,In_328,In_1716);
xor U724 (N_724,In_9,In_1072);
nand U725 (N_725,In_792,In_271);
xnor U726 (N_726,In_1756,In_1977);
nand U727 (N_727,In_784,In_1113);
and U728 (N_728,In_421,In_744);
and U729 (N_729,In_296,In_269);
nor U730 (N_730,In_1862,In_1189);
nand U731 (N_731,In_186,In_920);
xnor U732 (N_732,In_1278,In_1994);
xor U733 (N_733,In_1818,In_1204);
nand U734 (N_734,In_364,In_1085);
nand U735 (N_735,In_1117,In_1090);
nand U736 (N_736,In_509,In_466);
or U737 (N_737,In_1568,In_1017);
xor U738 (N_738,In_193,In_348);
nor U739 (N_739,In_966,In_1683);
nor U740 (N_740,In_722,In_1487);
xnor U741 (N_741,In_369,In_1185);
or U742 (N_742,In_1041,In_1768);
nor U743 (N_743,In_1407,In_1776);
and U744 (N_744,In_745,In_1439);
nand U745 (N_745,In_1521,In_716);
or U746 (N_746,In_513,In_1290);
nor U747 (N_747,In_1383,In_460);
nor U748 (N_748,In_1860,In_531);
and U749 (N_749,In_1034,In_775);
nand U750 (N_750,In_796,In_921);
xnor U751 (N_751,In_718,In_1079);
nand U752 (N_752,In_480,In_533);
xnor U753 (N_753,In_634,In_39);
and U754 (N_754,In_1819,In_1649);
or U755 (N_755,In_1427,In_190);
or U756 (N_756,In_185,In_1371);
nor U757 (N_757,In_25,In_249);
or U758 (N_758,In_1893,In_1209);
nor U759 (N_759,In_448,In_797);
nand U760 (N_760,In_1370,In_1692);
nor U761 (N_761,In_321,In_650);
xnor U762 (N_762,In_1054,In_798);
nand U763 (N_763,In_1474,In_1669);
and U764 (N_764,In_264,In_1012);
xor U765 (N_765,In_1198,In_307);
nand U766 (N_766,In_1183,In_1749);
and U767 (N_767,In_138,In_172);
xnor U768 (N_768,In_1498,In_46);
nor U769 (N_769,In_933,In_761);
xor U770 (N_770,In_1934,In_1500);
and U771 (N_771,In_1494,In_1697);
nor U772 (N_772,In_917,In_878);
xor U773 (N_773,In_1036,In_391);
and U774 (N_774,In_908,In_760);
or U775 (N_775,In_1865,In_252);
and U776 (N_776,In_1621,In_1996);
nor U777 (N_777,In_65,In_693);
nor U778 (N_778,In_1207,In_1225);
or U779 (N_779,In_897,In_104);
nand U780 (N_780,In_1721,In_1548);
and U781 (N_781,In_1680,In_1660);
nor U782 (N_782,In_710,In_406);
xnor U783 (N_783,In_1806,In_762);
nor U784 (N_784,In_1539,In_1210);
xnor U785 (N_785,In_1056,In_1110);
nor U786 (N_786,In_609,In_390);
xor U787 (N_787,In_1969,In_1387);
nand U788 (N_788,In_433,In_598);
nand U789 (N_789,In_788,In_910);
or U790 (N_790,In_1875,In_1814);
xnor U791 (N_791,In_980,In_928);
nand U792 (N_792,In_774,In_1748);
nor U793 (N_793,In_1305,In_222);
nand U794 (N_794,In_1792,In_208);
or U795 (N_795,In_90,In_1334);
xnor U796 (N_796,In_243,In_438);
xor U797 (N_797,In_132,In_217);
nor U798 (N_798,In_1430,In_939);
nand U799 (N_799,In_47,In_1192);
xnor U800 (N_800,In_1233,In_610);
nor U801 (N_801,In_1541,In_81);
or U802 (N_802,In_1363,In_662);
nor U803 (N_803,In_941,In_1342);
nor U804 (N_804,In_1327,In_729);
xnor U805 (N_805,In_1086,In_1975);
and U806 (N_806,In_270,In_1452);
xor U807 (N_807,In_1181,In_1273);
nor U808 (N_808,In_892,In_1405);
xnor U809 (N_809,In_1962,In_576);
xor U810 (N_810,In_539,In_1096);
xor U811 (N_811,In_386,In_44);
xnor U812 (N_812,In_196,In_318);
or U813 (N_813,In_211,In_494);
nand U814 (N_814,In_388,In_366);
and U815 (N_815,In_588,In_226);
and U816 (N_816,In_842,In_845);
nand U817 (N_817,In_618,In_1114);
nand U818 (N_818,In_819,In_1579);
and U819 (N_819,In_1035,In_1433);
xnor U820 (N_820,In_1332,In_714);
and U821 (N_821,In_1958,In_362);
nor U822 (N_822,In_1836,In_334);
nand U823 (N_823,In_1381,In_1145);
and U824 (N_824,In_1955,In_335);
nor U825 (N_825,In_1635,In_155);
and U826 (N_826,In_611,In_336);
or U827 (N_827,In_1443,In_644);
xor U828 (N_828,In_114,In_1662);
nor U829 (N_829,In_1115,In_337);
nand U830 (N_830,In_1857,In_1877);
nand U831 (N_831,In_828,In_1742);
xor U832 (N_832,In_1263,In_1665);
xor U833 (N_833,In_241,In_288);
or U834 (N_834,In_594,In_896);
or U835 (N_835,In_347,In_1973);
xor U836 (N_836,In_1311,In_1492);
or U837 (N_837,In_835,In_250);
and U838 (N_838,In_1403,In_853);
or U839 (N_839,In_1644,In_688);
nor U840 (N_840,In_1959,In_274);
and U841 (N_841,In_1398,In_1677);
or U842 (N_842,In_1691,In_663);
nand U843 (N_843,In_677,In_780);
and U844 (N_844,In_1645,In_346);
and U845 (N_845,In_1466,In_717);
xor U846 (N_846,In_1094,In_1667);
and U847 (N_847,In_1562,In_500);
or U848 (N_848,In_1570,In_676);
nor U849 (N_849,In_809,In_398);
nand U850 (N_850,In_887,In_16);
nand U851 (N_851,In_1257,In_736);
or U852 (N_852,In_18,In_1306);
and U853 (N_853,In_1643,In_95);
and U854 (N_854,In_1006,In_600);
or U855 (N_855,In_1820,In_245);
and U856 (N_856,In_884,In_478);
or U857 (N_857,In_1322,In_400);
or U858 (N_858,In_128,In_1281);
nand U859 (N_859,In_1261,In_1324);
and U860 (N_860,In_791,In_970);
and U861 (N_861,In_1713,In_1894);
nand U862 (N_862,In_1737,In_888);
and U863 (N_863,In_295,In_8);
and U864 (N_864,In_577,In_695);
nor U865 (N_865,In_1598,In_639);
nand U866 (N_866,In_89,In_1141);
or U867 (N_867,In_670,In_992);
nor U868 (N_868,In_591,In_78);
xor U869 (N_869,In_865,In_1699);
or U870 (N_870,In_1674,In_713);
and U871 (N_871,In_1091,In_1632);
nand U872 (N_872,In_476,In_872);
nor U873 (N_873,In_781,In_633);
nor U874 (N_874,In_1831,In_482);
nor U875 (N_875,In_1943,In_405);
and U876 (N_876,In_1989,In_282);
or U877 (N_877,In_162,In_1735);
and U878 (N_878,In_1150,In_1898);
nand U879 (N_879,In_1774,In_1038);
or U880 (N_880,In_680,In_1316);
and U881 (N_881,In_1229,In_818);
xor U882 (N_882,In_1274,In_1594);
nand U883 (N_883,In_776,In_1574);
nand U884 (N_884,In_859,In_451);
nand U885 (N_885,In_1730,In_524);
and U886 (N_886,In_1174,In_1529);
and U887 (N_887,In_1011,In_29);
and U888 (N_888,In_983,In_898);
nor U889 (N_889,In_1524,In_1798);
nand U890 (N_890,In_687,In_428);
and U891 (N_891,In_1074,In_625);
and U892 (N_892,In_499,In_1551);
nor U893 (N_893,In_733,In_1961);
nor U894 (N_894,In_525,In_1297);
xor U895 (N_895,In_1255,In_358);
and U896 (N_896,In_753,In_1953);
xnor U897 (N_897,In_868,In_851);
and U898 (N_898,In_1618,In_487);
or U899 (N_899,In_674,In_547);
nor U900 (N_900,In_880,In_1356);
xor U901 (N_901,In_1736,In_758);
or U902 (N_902,In_1132,In_314);
xnor U903 (N_903,In_1326,In_604);
nand U904 (N_904,In_1638,In_1540);
or U905 (N_905,In_490,In_1015);
nand U906 (N_906,In_1620,In_1236);
or U907 (N_907,In_1684,In_1720);
xor U908 (N_908,In_454,In_1081);
and U909 (N_909,In_709,In_948);
and U910 (N_910,In_1254,In_1221);
nand U911 (N_911,In_584,In_126);
nor U912 (N_912,In_374,In_246);
and U913 (N_913,In_156,In_502);
nor U914 (N_914,In_1653,In_213);
and U915 (N_915,In_1416,In_653);
nor U916 (N_916,In_1719,In_1373);
and U917 (N_917,In_699,In_757);
nand U918 (N_918,In_1982,In_891);
nor U919 (N_919,In_1307,In_255);
nor U920 (N_920,In_6,In_420);
xnor U921 (N_921,In_877,In_661);
nand U922 (N_922,In_1391,In_940);
nor U923 (N_923,In_1679,In_1251);
or U924 (N_924,In_1460,In_340);
xnor U925 (N_925,In_1138,In_988);
nor U926 (N_926,In_1505,In_945);
and U927 (N_927,In_1293,In_1599);
xor U928 (N_928,In_816,In_1376);
nor U929 (N_929,In_1484,In_1424);
and U930 (N_930,In_1134,In_1330);
nand U931 (N_931,In_1852,In_1313);
and U932 (N_932,In_1686,In_1711);
xor U933 (N_933,In_180,In_1972);
or U934 (N_934,In_323,In_1349);
and U935 (N_935,In_1704,In_147);
nor U936 (N_936,In_1627,In_852);
xnor U937 (N_937,In_1172,In_1393);
nand U938 (N_938,In_748,In_462);
and U939 (N_939,In_385,In_164);
nand U940 (N_940,In_619,In_1876);
nand U941 (N_941,In_1789,In_622);
and U942 (N_942,In_1939,In_1300);
and U943 (N_943,In_118,In_802);
xor U944 (N_944,In_1573,In_1188);
and U945 (N_945,In_739,In_867);
nand U946 (N_946,In_62,In_773);
and U947 (N_947,In_1400,In_1681);
xnor U948 (N_948,In_1402,In_426);
nand U949 (N_949,In_926,In_96);
nor U950 (N_950,In_1315,In_445);
nor U951 (N_951,In_1979,In_1547);
and U952 (N_952,In_569,In_163);
and U953 (N_953,In_294,In_113);
nor U954 (N_954,In_1060,In_961);
nand U955 (N_955,In_573,In_652);
nand U956 (N_956,In_1256,In_1693);
and U957 (N_957,In_1585,In_1947);
and U958 (N_958,In_1195,In_532);
and U959 (N_959,In_1467,In_514);
xor U960 (N_960,In_1636,In_119);
xnor U961 (N_961,In_1476,In_860);
nand U962 (N_962,In_679,In_1917);
xnor U963 (N_963,In_1914,In_647);
xnor U964 (N_964,In_1092,In_782);
or U965 (N_965,In_1039,In_1124);
xnor U966 (N_966,In_1137,In_1705);
nor U967 (N_967,In_1002,In_556);
or U968 (N_968,In_1312,In_1976);
nand U969 (N_969,In_467,In_1747);
xnor U970 (N_970,In_1217,In_1970);
xnor U971 (N_971,In_675,In_1151);
and U972 (N_972,In_821,In_559);
nor U973 (N_973,In_1837,In_1010);
or U974 (N_974,In_1176,In_1178);
xor U975 (N_975,In_1379,In_1567);
nor U976 (N_976,In_1827,In_976);
or U977 (N_977,In_527,In_301);
nor U978 (N_978,In_1952,In_131);
or U979 (N_979,In_1924,In_55);
and U980 (N_980,In_904,In_1139);
nand U981 (N_981,In_1473,In_1786);
nand U982 (N_982,In_1712,In_1963);
xnor U983 (N_983,In_959,In_179);
xor U984 (N_984,In_1563,In_1511);
xnor U985 (N_985,In_1435,In_1690);
and U986 (N_986,In_683,In_1739);
nand U987 (N_987,In_1863,In_237);
nand U988 (N_988,In_1853,In_1037);
or U989 (N_989,In_684,In_1942);
and U990 (N_990,In_1404,In_846);
nor U991 (N_991,In_552,In_1279);
nand U992 (N_992,In_1016,In_173);
nand U993 (N_993,In_15,In_1757);
nor U994 (N_994,In_392,In_1438);
and U995 (N_995,In_507,In_627);
or U996 (N_996,In_1418,In_1733);
nor U997 (N_997,In_923,In_1971);
or U998 (N_998,In_931,In_1062);
xnor U999 (N_999,In_1222,In_40);
nor U1000 (N_1000,In_876,In_1274);
nand U1001 (N_1001,In_1702,In_376);
nand U1002 (N_1002,In_1890,In_297);
and U1003 (N_1003,In_1711,In_1701);
or U1004 (N_1004,In_122,In_1005);
nand U1005 (N_1005,In_863,In_837);
or U1006 (N_1006,In_1216,In_1771);
or U1007 (N_1007,In_841,In_1495);
and U1008 (N_1008,In_1969,In_1341);
and U1009 (N_1009,In_699,In_367);
xnor U1010 (N_1010,In_72,In_1597);
and U1011 (N_1011,In_1127,In_192);
xor U1012 (N_1012,In_1098,In_1831);
nor U1013 (N_1013,In_591,In_1554);
nor U1014 (N_1014,In_3,In_67);
and U1015 (N_1015,In_1863,In_302);
or U1016 (N_1016,In_1928,In_1302);
and U1017 (N_1017,In_1608,In_653);
and U1018 (N_1018,In_1105,In_924);
and U1019 (N_1019,In_1665,In_239);
or U1020 (N_1020,In_567,In_1006);
and U1021 (N_1021,In_442,In_1890);
nand U1022 (N_1022,In_1939,In_1794);
nor U1023 (N_1023,In_1972,In_966);
and U1024 (N_1024,In_1524,In_447);
xor U1025 (N_1025,In_1338,In_387);
or U1026 (N_1026,In_166,In_1300);
nor U1027 (N_1027,In_1036,In_215);
nand U1028 (N_1028,In_423,In_387);
nor U1029 (N_1029,In_1367,In_1946);
xnor U1030 (N_1030,In_556,In_1184);
or U1031 (N_1031,In_1553,In_1628);
nor U1032 (N_1032,In_623,In_1550);
or U1033 (N_1033,In_1185,In_350);
or U1034 (N_1034,In_823,In_1810);
nand U1035 (N_1035,In_1947,In_1955);
and U1036 (N_1036,In_114,In_1161);
xnor U1037 (N_1037,In_1057,In_1677);
xor U1038 (N_1038,In_1995,In_1330);
and U1039 (N_1039,In_1939,In_1019);
nand U1040 (N_1040,In_1915,In_995);
nand U1041 (N_1041,In_184,In_234);
or U1042 (N_1042,In_1588,In_580);
nand U1043 (N_1043,In_954,In_151);
xor U1044 (N_1044,In_289,In_1560);
xnor U1045 (N_1045,In_376,In_1803);
or U1046 (N_1046,In_1498,In_1359);
and U1047 (N_1047,In_1585,In_1665);
nor U1048 (N_1048,In_1604,In_430);
nor U1049 (N_1049,In_991,In_85);
xor U1050 (N_1050,In_208,In_1830);
xnor U1051 (N_1051,In_227,In_528);
nor U1052 (N_1052,In_430,In_1536);
xnor U1053 (N_1053,In_206,In_12);
or U1054 (N_1054,In_601,In_733);
xnor U1055 (N_1055,In_408,In_133);
xnor U1056 (N_1056,In_768,In_1048);
nand U1057 (N_1057,In_682,In_792);
nand U1058 (N_1058,In_701,In_1892);
nand U1059 (N_1059,In_1560,In_300);
and U1060 (N_1060,In_1274,In_1331);
or U1061 (N_1061,In_790,In_255);
nand U1062 (N_1062,In_1145,In_958);
or U1063 (N_1063,In_1335,In_267);
nand U1064 (N_1064,In_460,In_138);
nand U1065 (N_1065,In_665,In_291);
and U1066 (N_1066,In_545,In_688);
and U1067 (N_1067,In_360,In_1943);
nand U1068 (N_1068,In_1133,In_1191);
or U1069 (N_1069,In_1716,In_1324);
nor U1070 (N_1070,In_852,In_578);
xnor U1071 (N_1071,In_563,In_1725);
xnor U1072 (N_1072,In_349,In_1090);
xor U1073 (N_1073,In_549,In_1187);
nor U1074 (N_1074,In_550,In_1284);
xnor U1075 (N_1075,In_769,In_542);
xnor U1076 (N_1076,In_953,In_607);
xor U1077 (N_1077,In_432,In_1182);
nor U1078 (N_1078,In_27,In_1585);
nor U1079 (N_1079,In_1228,In_361);
or U1080 (N_1080,In_498,In_344);
nor U1081 (N_1081,In_1892,In_781);
xnor U1082 (N_1082,In_873,In_897);
or U1083 (N_1083,In_642,In_901);
xor U1084 (N_1084,In_1306,In_1377);
nor U1085 (N_1085,In_1513,In_756);
and U1086 (N_1086,In_718,In_1861);
and U1087 (N_1087,In_122,In_1195);
xnor U1088 (N_1088,In_905,In_1573);
nor U1089 (N_1089,In_1486,In_294);
nor U1090 (N_1090,In_432,In_643);
xnor U1091 (N_1091,In_352,In_152);
nand U1092 (N_1092,In_1219,In_863);
nand U1093 (N_1093,In_468,In_1179);
or U1094 (N_1094,In_30,In_1405);
and U1095 (N_1095,In_1349,In_34);
xor U1096 (N_1096,In_581,In_1849);
nor U1097 (N_1097,In_1096,In_1708);
nand U1098 (N_1098,In_913,In_1185);
xnor U1099 (N_1099,In_1966,In_782);
nand U1100 (N_1100,In_103,In_1640);
nor U1101 (N_1101,In_119,In_1842);
or U1102 (N_1102,In_478,In_146);
or U1103 (N_1103,In_1969,In_248);
or U1104 (N_1104,In_1521,In_1630);
nand U1105 (N_1105,In_976,In_829);
nand U1106 (N_1106,In_1551,In_531);
nand U1107 (N_1107,In_1882,In_1279);
nor U1108 (N_1108,In_1526,In_494);
xnor U1109 (N_1109,In_116,In_752);
xnor U1110 (N_1110,In_1901,In_1671);
nand U1111 (N_1111,In_355,In_1071);
nor U1112 (N_1112,In_1199,In_459);
and U1113 (N_1113,In_1174,In_378);
xnor U1114 (N_1114,In_864,In_1642);
nand U1115 (N_1115,In_796,In_164);
xnor U1116 (N_1116,In_1577,In_1558);
and U1117 (N_1117,In_1431,In_1485);
nand U1118 (N_1118,In_611,In_962);
nand U1119 (N_1119,In_1388,In_1428);
xor U1120 (N_1120,In_315,In_1254);
nand U1121 (N_1121,In_1164,In_1683);
nand U1122 (N_1122,In_751,In_1147);
nand U1123 (N_1123,In_1998,In_1679);
and U1124 (N_1124,In_115,In_95);
and U1125 (N_1125,In_1817,In_1947);
xnor U1126 (N_1126,In_1709,In_1984);
and U1127 (N_1127,In_1668,In_1117);
xnor U1128 (N_1128,In_1290,In_1533);
and U1129 (N_1129,In_257,In_1659);
xnor U1130 (N_1130,In_1050,In_1971);
nor U1131 (N_1131,In_550,In_1444);
xnor U1132 (N_1132,In_188,In_44);
and U1133 (N_1133,In_955,In_1171);
or U1134 (N_1134,In_1642,In_1513);
or U1135 (N_1135,In_1140,In_1821);
nor U1136 (N_1136,In_1915,In_1953);
or U1137 (N_1137,In_785,In_1568);
nand U1138 (N_1138,In_1018,In_262);
nor U1139 (N_1139,In_196,In_1780);
and U1140 (N_1140,In_1631,In_1503);
and U1141 (N_1141,In_1363,In_1534);
and U1142 (N_1142,In_51,In_1437);
xnor U1143 (N_1143,In_348,In_1359);
and U1144 (N_1144,In_1704,In_1447);
or U1145 (N_1145,In_1811,In_618);
and U1146 (N_1146,In_1972,In_656);
nor U1147 (N_1147,In_1954,In_841);
nand U1148 (N_1148,In_1388,In_1176);
nor U1149 (N_1149,In_885,In_543);
xor U1150 (N_1150,In_1373,In_1009);
nand U1151 (N_1151,In_1308,In_1559);
nor U1152 (N_1152,In_1072,In_1128);
nor U1153 (N_1153,In_1873,In_885);
nand U1154 (N_1154,In_904,In_1502);
xnor U1155 (N_1155,In_1858,In_486);
nor U1156 (N_1156,In_615,In_1367);
nand U1157 (N_1157,In_387,In_1057);
nand U1158 (N_1158,In_1639,In_1002);
nor U1159 (N_1159,In_1379,In_204);
nand U1160 (N_1160,In_1442,In_807);
and U1161 (N_1161,In_1179,In_93);
nor U1162 (N_1162,In_1316,In_1478);
nand U1163 (N_1163,In_827,In_1208);
and U1164 (N_1164,In_1258,In_1895);
and U1165 (N_1165,In_1523,In_699);
or U1166 (N_1166,In_242,In_1504);
or U1167 (N_1167,In_1554,In_405);
or U1168 (N_1168,In_986,In_965);
xnor U1169 (N_1169,In_471,In_682);
or U1170 (N_1170,In_1187,In_984);
or U1171 (N_1171,In_1907,In_1771);
xnor U1172 (N_1172,In_1692,In_452);
and U1173 (N_1173,In_357,In_844);
and U1174 (N_1174,In_1163,In_728);
and U1175 (N_1175,In_58,In_898);
xnor U1176 (N_1176,In_872,In_843);
and U1177 (N_1177,In_1665,In_1435);
and U1178 (N_1178,In_671,In_1537);
and U1179 (N_1179,In_501,In_1050);
nor U1180 (N_1180,In_1938,In_242);
nor U1181 (N_1181,In_1616,In_1874);
and U1182 (N_1182,In_1790,In_274);
nand U1183 (N_1183,In_196,In_1288);
xnor U1184 (N_1184,In_1515,In_265);
nor U1185 (N_1185,In_1984,In_1130);
and U1186 (N_1186,In_541,In_942);
nor U1187 (N_1187,In_1452,In_882);
or U1188 (N_1188,In_1486,In_1298);
nor U1189 (N_1189,In_1712,In_1942);
or U1190 (N_1190,In_1708,In_607);
or U1191 (N_1191,In_1547,In_177);
or U1192 (N_1192,In_838,In_440);
nand U1193 (N_1193,In_75,In_1505);
nand U1194 (N_1194,In_1556,In_1555);
nand U1195 (N_1195,In_826,In_1337);
or U1196 (N_1196,In_1785,In_1627);
nand U1197 (N_1197,In_1706,In_90);
nor U1198 (N_1198,In_823,In_209);
or U1199 (N_1199,In_1842,In_952);
nand U1200 (N_1200,In_1743,In_1996);
nand U1201 (N_1201,In_476,In_349);
xnor U1202 (N_1202,In_1967,In_901);
and U1203 (N_1203,In_1198,In_1383);
xor U1204 (N_1204,In_1872,In_933);
nand U1205 (N_1205,In_725,In_768);
nand U1206 (N_1206,In_1317,In_864);
xor U1207 (N_1207,In_754,In_640);
nand U1208 (N_1208,In_167,In_1098);
nand U1209 (N_1209,In_1038,In_706);
nand U1210 (N_1210,In_288,In_1925);
nand U1211 (N_1211,In_1230,In_859);
nand U1212 (N_1212,In_468,In_1250);
and U1213 (N_1213,In_1609,In_926);
or U1214 (N_1214,In_609,In_1726);
nor U1215 (N_1215,In_1093,In_1329);
and U1216 (N_1216,In_796,In_126);
and U1217 (N_1217,In_1078,In_735);
xnor U1218 (N_1218,In_1665,In_1831);
or U1219 (N_1219,In_1826,In_1166);
and U1220 (N_1220,In_1406,In_1666);
nand U1221 (N_1221,In_844,In_1283);
xnor U1222 (N_1222,In_1577,In_1833);
nor U1223 (N_1223,In_241,In_536);
xnor U1224 (N_1224,In_216,In_1942);
or U1225 (N_1225,In_925,In_453);
xnor U1226 (N_1226,In_1082,In_1378);
and U1227 (N_1227,In_596,In_164);
nor U1228 (N_1228,In_907,In_1018);
xnor U1229 (N_1229,In_543,In_408);
xor U1230 (N_1230,In_1724,In_454);
xor U1231 (N_1231,In_1074,In_46);
and U1232 (N_1232,In_430,In_234);
nand U1233 (N_1233,In_818,In_895);
nand U1234 (N_1234,In_221,In_1028);
nor U1235 (N_1235,In_1010,In_583);
xnor U1236 (N_1236,In_1970,In_1363);
nor U1237 (N_1237,In_1105,In_889);
or U1238 (N_1238,In_658,In_105);
nand U1239 (N_1239,In_98,In_950);
or U1240 (N_1240,In_1388,In_985);
and U1241 (N_1241,In_1254,In_323);
and U1242 (N_1242,In_1559,In_1208);
xnor U1243 (N_1243,In_107,In_182);
xnor U1244 (N_1244,In_362,In_1481);
nand U1245 (N_1245,In_424,In_123);
or U1246 (N_1246,In_371,In_216);
nor U1247 (N_1247,In_1433,In_419);
or U1248 (N_1248,In_324,In_1750);
and U1249 (N_1249,In_1739,In_1873);
nand U1250 (N_1250,In_1828,In_505);
nor U1251 (N_1251,In_829,In_1513);
or U1252 (N_1252,In_344,In_1166);
and U1253 (N_1253,In_143,In_663);
and U1254 (N_1254,In_1451,In_470);
nor U1255 (N_1255,In_676,In_1419);
xnor U1256 (N_1256,In_1466,In_1684);
nand U1257 (N_1257,In_145,In_1714);
or U1258 (N_1258,In_1493,In_1075);
and U1259 (N_1259,In_840,In_489);
and U1260 (N_1260,In_1770,In_1496);
xor U1261 (N_1261,In_638,In_1909);
xor U1262 (N_1262,In_1074,In_871);
nor U1263 (N_1263,In_1837,In_840);
xnor U1264 (N_1264,In_150,In_867);
and U1265 (N_1265,In_1219,In_568);
and U1266 (N_1266,In_1932,In_1694);
nand U1267 (N_1267,In_650,In_71);
and U1268 (N_1268,In_194,In_1276);
or U1269 (N_1269,In_904,In_1434);
or U1270 (N_1270,In_664,In_678);
and U1271 (N_1271,In_1412,In_1046);
or U1272 (N_1272,In_1995,In_332);
or U1273 (N_1273,In_1033,In_387);
and U1274 (N_1274,In_291,In_1977);
nand U1275 (N_1275,In_1164,In_1087);
and U1276 (N_1276,In_1773,In_1935);
and U1277 (N_1277,In_263,In_1266);
nand U1278 (N_1278,In_740,In_1162);
nor U1279 (N_1279,In_1188,In_1794);
xor U1280 (N_1280,In_1417,In_1211);
or U1281 (N_1281,In_1304,In_1916);
nand U1282 (N_1282,In_1301,In_1589);
nor U1283 (N_1283,In_1373,In_269);
nor U1284 (N_1284,In_1834,In_1191);
and U1285 (N_1285,In_515,In_493);
and U1286 (N_1286,In_1531,In_370);
and U1287 (N_1287,In_130,In_73);
nor U1288 (N_1288,In_247,In_1582);
and U1289 (N_1289,In_1665,In_139);
and U1290 (N_1290,In_1471,In_1228);
nor U1291 (N_1291,In_1139,In_1325);
xor U1292 (N_1292,In_190,In_1782);
or U1293 (N_1293,In_1030,In_1211);
xnor U1294 (N_1294,In_691,In_1181);
nand U1295 (N_1295,In_1644,In_729);
or U1296 (N_1296,In_1534,In_165);
xor U1297 (N_1297,In_1765,In_166);
or U1298 (N_1298,In_838,In_688);
nand U1299 (N_1299,In_1062,In_1628);
and U1300 (N_1300,In_809,In_598);
xnor U1301 (N_1301,In_106,In_429);
or U1302 (N_1302,In_1419,In_1392);
nor U1303 (N_1303,In_332,In_1533);
nor U1304 (N_1304,In_706,In_1007);
nand U1305 (N_1305,In_1922,In_1549);
or U1306 (N_1306,In_704,In_1491);
xnor U1307 (N_1307,In_1634,In_1837);
nor U1308 (N_1308,In_1023,In_687);
or U1309 (N_1309,In_1067,In_1227);
xor U1310 (N_1310,In_451,In_636);
xor U1311 (N_1311,In_1263,In_1456);
or U1312 (N_1312,In_1321,In_865);
nor U1313 (N_1313,In_1440,In_141);
or U1314 (N_1314,In_174,In_1876);
nand U1315 (N_1315,In_1920,In_1074);
and U1316 (N_1316,In_76,In_1815);
nor U1317 (N_1317,In_1930,In_252);
and U1318 (N_1318,In_1700,In_1262);
or U1319 (N_1319,In_1278,In_1545);
nor U1320 (N_1320,In_1314,In_69);
nor U1321 (N_1321,In_1604,In_1099);
xor U1322 (N_1322,In_1471,In_1040);
xor U1323 (N_1323,In_892,In_333);
xor U1324 (N_1324,In_440,In_1546);
and U1325 (N_1325,In_109,In_1001);
or U1326 (N_1326,In_87,In_504);
xor U1327 (N_1327,In_452,In_200);
or U1328 (N_1328,In_1998,In_1055);
xor U1329 (N_1329,In_912,In_785);
nor U1330 (N_1330,In_383,In_1746);
nor U1331 (N_1331,In_1415,In_1263);
nand U1332 (N_1332,In_1728,In_69);
or U1333 (N_1333,In_350,In_794);
or U1334 (N_1334,In_1783,In_1371);
or U1335 (N_1335,In_1351,In_1900);
xnor U1336 (N_1336,In_682,In_614);
xnor U1337 (N_1337,In_1006,In_1163);
or U1338 (N_1338,In_239,In_595);
nand U1339 (N_1339,In_1774,In_901);
nor U1340 (N_1340,In_703,In_197);
nand U1341 (N_1341,In_451,In_1623);
or U1342 (N_1342,In_1479,In_1766);
or U1343 (N_1343,In_1751,In_277);
nor U1344 (N_1344,In_1632,In_1726);
nand U1345 (N_1345,In_713,In_540);
xnor U1346 (N_1346,In_1968,In_783);
and U1347 (N_1347,In_1532,In_592);
nand U1348 (N_1348,In_1833,In_139);
nor U1349 (N_1349,In_424,In_585);
nand U1350 (N_1350,In_45,In_566);
and U1351 (N_1351,In_1627,In_409);
and U1352 (N_1352,In_521,In_513);
and U1353 (N_1353,In_1688,In_1486);
and U1354 (N_1354,In_769,In_468);
nor U1355 (N_1355,In_405,In_189);
and U1356 (N_1356,In_738,In_349);
or U1357 (N_1357,In_1508,In_1561);
and U1358 (N_1358,In_1553,In_550);
or U1359 (N_1359,In_214,In_973);
or U1360 (N_1360,In_829,In_1776);
and U1361 (N_1361,In_61,In_1274);
nand U1362 (N_1362,In_847,In_42);
and U1363 (N_1363,In_314,In_1336);
nor U1364 (N_1364,In_383,In_1353);
xor U1365 (N_1365,In_0,In_744);
nor U1366 (N_1366,In_1271,In_148);
nor U1367 (N_1367,In_626,In_280);
or U1368 (N_1368,In_1564,In_225);
nand U1369 (N_1369,In_29,In_756);
nor U1370 (N_1370,In_1631,In_247);
and U1371 (N_1371,In_1394,In_266);
or U1372 (N_1372,In_715,In_1144);
nor U1373 (N_1373,In_659,In_306);
and U1374 (N_1374,In_1309,In_512);
or U1375 (N_1375,In_1212,In_782);
nand U1376 (N_1376,In_1344,In_478);
nor U1377 (N_1377,In_257,In_1015);
nor U1378 (N_1378,In_157,In_116);
nor U1379 (N_1379,In_1153,In_896);
nor U1380 (N_1380,In_1797,In_1528);
or U1381 (N_1381,In_957,In_735);
xnor U1382 (N_1382,In_1775,In_878);
and U1383 (N_1383,In_1016,In_1855);
xnor U1384 (N_1384,In_1952,In_1439);
or U1385 (N_1385,In_623,In_609);
xnor U1386 (N_1386,In_497,In_143);
nor U1387 (N_1387,In_495,In_1447);
xor U1388 (N_1388,In_450,In_87);
nor U1389 (N_1389,In_1341,In_1948);
or U1390 (N_1390,In_824,In_1893);
nand U1391 (N_1391,In_867,In_526);
nor U1392 (N_1392,In_1158,In_1360);
xor U1393 (N_1393,In_4,In_1143);
xnor U1394 (N_1394,In_649,In_1766);
xnor U1395 (N_1395,In_1377,In_312);
or U1396 (N_1396,In_387,In_1961);
nor U1397 (N_1397,In_26,In_1759);
nor U1398 (N_1398,In_869,In_937);
or U1399 (N_1399,In_1173,In_1142);
nor U1400 (N_1400,In_1584,In_871);
xnor U1401 (N_1401,In_934,In_1947);
nand U1402 (N_1402,In_1948,In_1280);
nand U1403 (N_1403,In_1288,In_757);
and U1404 (N_1404,In_486,In_621);
or U1405 (N_1405,In_98,In_1807);
and U1406 (N_1406,In_882,In_690);
nand U1407 (N_1407,In_806,In_1312);
or U1408 (N_1408,In_525,In_283);
nand U1409 (N_1409,In_160,In_1998);
nand U1410 (N_1410,In_1252,In_1711);
xor U1411 (N_1411,In_635,In_973);
nand U1412 (N_1412,In_1638,In_1547);
or U1413 (N_1413,In_1309,In_1357);
nand U1414 (N_1414,In_734,In_1365);
or U1415 (N_1415,In_145,In_869);
and U1416 (N_1416,In_4,In_233);
and U1417 (N_1417,In_839,In_740);
nor U1418 (N_1418,In_285,In_372);
nand U1419 (N_1419,In_1034,In_864);
xor U1420 (N_1420,In_1579,In_604);
nand U1421 (N_1421,In_160,In_1756);
or U1422 (N_1422,In_11,In_831);
and U1423 (N_1423,In_287,In_1667);
nand U1424 (N_1424,In_1589,In_1204);
and U1425 (N_1425,In_1422,In_1153);
nor U1426 (N_1426,In_1869,In_188);
nor U1427 (N_1427,In_1970,In_1815);
nor U1428 (N_1428,In_1790,In_1005);
nand U1429 (N_1429,In_1525,In_964);
and U1430 (N_1430,In_289,In_832);
and U1431 (N_1431,In_90,In_578);
nand U1432 (N_1432,In_231,In_848);
nor U1433 (N_1433,In_1387,In_1070);
xor U1434 (N_1434,In_775,In_1009);
nor U1435 (N_1435,In_521,In_4);
nor U1436 (N_1436,In_353,In_1617);
and U1437 (N_1437,In_1078,In_437);
nand U1438 (N_1438,In_584,In_1353);
xor U1439 (N_1439,In_1959,In_429);
nor U1440 (N_1440,In_499,In_301);
nand U1441 (N_1441,In_1048,In_543);
nand U1442 (N_1442,In_1398,In_289);
nand U1443 (N_1443,In_508,In_1058);
or U1444 (N_1444,In_607,In_1186);
and U1445 (N_1445,In_1878,In_1530);
nand U1446 (N_1446,In_1208,In_967);
or U1447 (N_1447,In_787,In_102);
nand U1448 (N_1448,In_1027,In_1119);
and U1449 (N_1449,In_1456,In_1583);
nand U1450 (N_1450,In_1817,In_653);
nor U1451 (N_1451,In_397,In_1327);
xor U1452 (N_1452,In_1887,In_1191);
nand U1453 (N_1453,In_1170,In_1908);
xor U1454 (N_1454,In_1143,In_1662);
and U1455 (N_1455,In_929,In_771);
and U1456 (N_1456,In_1777,In_1910);
or U1457 (N_1457,In_1394,In_1951);
xnor U1458 (N_1458,In_1260,In_1732);
or U1459 (N_1459,In_1569,In_165);
nor U1460 (N_1460,In_1685,In_788);
and U1461 (N_1461,In_1939,In_388);
or U1462 (N_1462,In_86,In_682);
or U1463 (N_1463,In_517,In_468);
or U1464 (N_1464,In_820,In_1507);
and U1465 (N_1465,In_249,In_39);
nand U1466 (N_1466,In_1703,In_1629);
and U1467 (N_1467,In_43,In_1324);
or U1468 (N_1468,In_1043,In_1841);
nor U1469 (N_1469,In_1412,In_1289);
or U1470 (N_1470,In_1362,In_934);
or U1471 (N_1471,In_801,In_399);
and U1472 (N_1472,In_1633,In_1282);
nor U1473 (N_1473,In_1136,In_1056);
and U1474 (N_1474,In_519,In_1958);
nand U1475 (N_1475,In_1183,In_1659);
nand U1476 (N_1476,In_228,In_579);
nor U1477 (N_1477,In_1320,In_1960);
nand U1478 (N_1478,In_1171,In_285);
and U1479 (N_1479,In_645,In_1110);
nand U1480 (N_1480,In_143,In_1009);
nand U1481 (N_1481,In_19,In_1144);
xnor U1482 (N_1482,In_1279,In_993);
and U1483 (N_1483,In_1768,In_1904);
or U1484 (N_1484,In_58,In_393);
or U1485 (N_1485,In_618,In_194);
or U1486 (N_1486,In_1973,In_217);
and U1487 (N_1487,In_904,In_1928);
nor U1488 (N_1488,In_1849,In_819);
and U1489 (N_1489,In_1312,In_650);
or U1490 (N_1490,In_1648,In_1930);
nand U1491 (N_1491,In_1606,In_1065);
and U1492 (N_1492,In_1914,In_215);
xnor U1493 (N_1493,In_1778,In_1108);
and U1494 (N_1494,In_1947,In_559);
nor U1495 (N_1495,In_1275,In_32);
nor U1496 (N_1496,In_929,In_339);
xnor U1497 (N_1497,In_1472,In_67);
xnor U1498 (N_1498,In_356,In_47);
nor U1499 (N_1499,In_315,In_1745);
and U1500 (N_1500,In_1076,In_1019);
nand U1501 (N_1501,In_1236,In_115);
and U1502 (N_1502,In_158,In_841);
nor U1503 (N_1503,In_1178,In_1389);
nor U1504 (N_1504,In_870,In_995);
and U1505 (N_1505,In_687,In_1540);
nand U1506 (N_1506,In_190,In_1925);
or U1507 (N_1507,In_121,In_482);
and U1508 (N_1508,In_277,In_222);
and U1509 (N_1509,In_1703,In_961);
xor U1510 (N_1510,In_1348,In_541);
xor U1511 (N_1511,In_1471,In_34);
or U1512 (N_1512,In_1523,In_820);
and U1513 (N_1513,In_730,In_846);
or U1514 (N_1514,In_1668,In_1805);
nor U1515 (N_1515,In_1419,In_662);
xor U1516 (N_1516,In_827,In_1338);
nor U1517 (N_1517,In_977,In_1568);
nand U1518 (N_1518,In_171,In_1073);
nand U1519 (N_1519,In_1521,In_1537);
xnor U1520 (N_1520,In_340,In_194);
nor U1521 (N_1521,In_1886,In_552);
nand U1522 (N_1522,In_864,In_252);
xnor U1523 (N_1523,In_1952,In_1852);
and U1524 (N_1524,In_29,In_868);
nor U1525 (N_1525,In_1718,In_233);
or U1526 (N_1526,In_1297,In_182);
nor U1527 (N_1527,In_220,In_1368);
nor U1528 (N_1528,In_172,In_537);
and U1529 (N_1529,In_1764,In_287);
xnor U1530 (N_1530,In_525,In_1120);
or U1531 (N_1531,In_438,In_1017);
nor U1532 (N_1532,In_671,In_227);
and U1533 (N_1533,In_1108,In_199);
xor U1534 (N_1534,In_1663,In_1678);
xor U1535 (N_1535,In_1287,In_1393);
or U1536 (N_1536,In_742,In_1438);
nand U1537 (N_1537,In_1046,In_1069);
and U1538 (N_1538,In_418,In_1696);
xnor U1539 (N_1539,In_1891,In_162);
or U1540 (N_1540,In_353,In_1656);
and U1541 (N_1541,In_1344,In_1746);
xor U1542 (N_1542,In_1302,In_887);
nand U1543 (N_1543,In_376,In_193);
nand U1544 (N_1544,In_57,In_79);
and U1545 (N_1545,In_1231,In_881);
xnor U1546 (N_1546,In_1006,In_1732);
and U1547 (N_1547,In_1138,In_1196);
or U1548 (N_1548,In_1043,In_653);
xnor U1549 (N_1549,In_288,In_1012);
nor U1550 (N_1550,In_991,In_1100);
and U1551 (N_1551,In_1238,In_1351);
nand U1552 (N_1552,In_1636,In_1043);
or U1553 (N_1553,In_1843,In_1952);
and U1554 (N_1554,In_549,In_1326);
xnor U1555 (N_1555,In_1209,In_75);
and U1556 (N_1556,In_453,In_1075);
xnor U1557 (N_1557,In_636,In_621);
xor U1558 (N_1558,In_1396,In_1750);
xor U1559 (N_1559,In_1157,In_999);
or U1560 (N_1560,In_110,In_149);
xor U1561 (N_1561,In_1215,In_1237);
nor U1562 (N_1562,In_906,In_1737);
nand U1563 (N_1563,In_1295,In_318);
and U1564 (N_1564,In_1697,In_351);
nor U1565 (N_1565,In_795,In_707);
nand U1566 (N_1566,In_1288,In_294);
xor U1567 (N_1567,In_359,In_452);
and U1568 (N_1568,In_721,In_1786);
nand U1569 (N_1569,In_555,In_841);
nor U1570 (N_1570,In_1513,In_1589);
xor U1571 (N_1571,In_1268,In_1954);
or U1572 (N_1572,In_1250,In_1473);
or U1573 (N_1573,In_101,In_1304);
and U1574 (N_1574,In_228,In_200);
or U1575 (N_1575,In_64,In_646);
xor U1576 (N_1576,In_389,In_704);
nor U1577 (N_1577,In_28,In_1163);
or U1578 (N_1578,In_1058,In_756);
xor U1579 (N_1579,In_1815,In_123);
and U1580 (N_1580,In_1641,In_246);
and U1581 (N_1581,In_314,In_412);
nand U1582 (N_1582,In_1184,In_207);
or U1583 (N_1583,In_258,In_1974);
xnor U1584 (N_1584,In_225,In_421);
nor U1585 (N_1585,In_1987,In_1189);
or U1586 (N_1586,In_1767,In_439);
nor U1587 (N_1587,In_1759,In_1203);
or U1588 (N_1588,In_577,In_1669);
xnor U1589 (N_1589,In_1428,In_1762);
xnor U1590 (N_1590,In_1687,In_531);
or U1591 (N_1591,In_629,In_73);
and U1592 (N_1592,In_1574,In_1351);
or U1593 (N_1593,In_1510,In_868);
and U1594 (N_1594,In_1989,In_1021);
nor U1595 (N_1595,In_1918,In_1326);
nor U1596 (N_1596,In_731,In_600);
and U1597 (N_1597,In_1342,In_520);
or U1598 (N_1598,In_143,In_224);
nand U1599 (N_1599,In_1141,In_120);
and U1600 (N_1600,In_1076,In_626);
xnor U1601 (N_1601,In_1486,In_207);
and U1602 (N_1602,In_238,In_1503);
or U1603 (N_1603,In_1215,In_952);
and U1604 (N_1604,In_1262,In_1558);
xor U1605 (N_1605,In_969,In_999);
nand U1606 (N_1606,In_43,In_299);
and U1607 (N_1607,In_753,In_1685);
xnor U1608 (N_1608,In_219,In_357);
or U1609 (N_1609,In_203,In_1291);
or U1610 (N_1610,In_1105,In_1362);
or U1611 (N_1611,In_743,In_1903);
and U1612 (N_1612,In_1087,In_1185);
or U1613 (N_1613,In_1999,In_759);
and U1614 (N_1614,In_948,In_1312);
nor U1615 (N_1615,In_1782,In_5);
or U1616 (N_1616,In_1638,In_66);
or U1617 (N_1617,In_668,In_1167);
and U1618 (N_1618,In_988,In_1930);
nor U1619 (N_1619,In_1110,In_1922);
and U1620 (N_1620,In_455,In_226);
or U1621 (N_1621,In_1881,In_229);
or U1622 (N_1622,In_387,In_1971);
nand U1623 (N_1623,In_873,In_148);
and U1624 (N_1624,In_531,In_31);
or U1625 (N_1625,In_421,In_1741);
nand U1626 (N_1626,In_1281,In_82);
xor U1627 (N_1627,In_1186,In_770);
and U1628 (N_1628,In_247,In_533);
and U1629 (N_1629,In_1856,In_1194);
nand U1630 (N_1630,In_1920,In_1524);
nor U1631 (N_1631,In_1292,In_1396);
xnor U1632 (N_1632,In_1016,In_573);
and U1633 (N_1633,In_144,In_1873);
and U1634 (N_1634,In_1820,In_1450);
and U1635 (N_1635,In_1920,In_1358);
nor U1636 (N_1636,In_1758,In_512);
or U1637 (N_1637,In_712,In_552);
nor U1638 (N_1638,In_809,In_805);
nor U1639 (N_1639,In_1056,In_1606);
nor U1640 (N_1640,In_630,In_1197);
and U1641 (N_1641,In_1647,In_363);
or U1642 (N_1642,In_1310,In_1428);
nor U1643 (N_1643,In_165,In_1236);
nand U1644 (N_1644,In_671,In_346);
nand U1645 (N_1645,In_635,In_715);
nor U1646 (N_1646,In_857,In_1882);
nand U1647 (N_1647,In_378,In_1361);
and U1648 (N_1648,In_1755,In_1771);
nand U1649 (N_1649,In_943,In_592);
and U1650 (N_1650,In_1968,In_455);
nor U1651 (N_1651,In_1914,In_175);
xnor U1652 (N_1652,In_1977,In_1440);
and U1653 (N_1653,In_1414,In_721);
xor U1654 (N_1654,In_1143,In_1020);
and U1655 (N_1655,In_327,In_243);
nand U1656 (N_1656,In_1855,In_1729);
and U1657 (N_1657,In_1486,In_656);
or U1658 (N_1658,In_1624,In_1721);
nor U1659 (N_1659,In_1970,In_175);
nor U1660 (N_1660,In_1358,In_1362);
and U1661 (N_1661,In_472,In_1961);
or U1662 (N_1662,In_749,In_244);
and U1663 (N_1663,In_948,In_1095);
and U1664 (N_1664,In_685,In_245);
nand U1665 (N_1665,In_1704,In_1638);
nand U1666 (N_1666,In_1934,In_1537);
nor U1667 (N_1667,In_434,In_1465);
nand U1668 (N_1668,In_396,In_1070);
or U1669 (N_1669,In_1818,In_1944);
nor U1670 (N_1670,In_1344,In_1618);
nand U1671 (N_1671,In_53,In_1632);
nand U1672 (N_1672,In_1124,In_1380);
nor U1673 (N_1673,In_1797,In_423);
and U1674 (N_1674,In_1400,In_462);
and U1675 (N_1675,In_1339,In_438);
xnor U1676 (N_1676,In_1969,In_177);
xnor U1677 (N_1677,In_1088,In_587);
nand U1678 (N_1678,In_824,In_1145);
xor U1679 (N_1679,In_129,In_1516);
or U1680 (N_1680,In_1381,In_540);
nand U1681 (N_1681,In_36,In_926);
nor U1682 (N_1682,In_1317,In_1292);
and U1683 (N_1683,In_956,In_1794);
and U1684 (N_1684,In_559,In_229);
nor U1685 (N_1685,In_419,In_108);
or U1686 (N_1686,In_1291,In_433);
xor U1687 (N_1687,In_1407,In_615);
or U1688 (N_1688,In_820,In_530);
xor U1689 (N_1689,In_1877,In_741);
nor U1690 (N_1690,In_819,In_1163);
nand U1691 (N_1691,In_1810,In_1160);
xor U1692 (N_1692,In_988,In_1847);
nand U1693 (N_1693,In_1157,In_1462);
xor U1694 (N_1694,In_832,In_1936);
nand U1695 (N_1695,In_1415,In_350);
nor U1696 (N_1696,In_752,In_1970);
or U1697 (N_1697,In_369,In_1289);
nor U1698 (N_1698,In_1805,In_1492);
nor U1699 (N_1699,In_594,In_1429);
and U1700 (N_1700,In_1577,In_344);
or U1701 (N_1701,In_1465,In_172);
nor U1702 (N_1702,In_1237,In_599);
nand U1703 (N_1703,In_1225,In_1937);
xor U1704 (N_1704,In_1446,In_1557);
nor U1705 (N_1705,In_1880,In_1602);
or U1706 (N_1706,In_966,In_1104);
and U1707 (N_1707,In_229,In_267);
or U1708 (N_1708,In_1118,In_352);
nand U1709 (N_1709,In_776,In_412);
xnor U1710 (N_1710,In_1544,In_1109);
nor U1711 (N_1711,In_678,In_1732);
xnor U1712 (N_1712,In_1961,In_866);
or U1713 (N_1713,In_928,In_1032);
and U1714 (N_1714,In_849,In_732);
and U1715 (N_1715,In_1827,In_1953);
or U1716 (N_1716,In_404,In_1154);
xnor U1717 (N_1717,In_1886,In_1048);
xnor U1718 (N_1718,In_1623,In_468);
nor U1719 (N_1719,In_1591,In_1779);
nor U1720 (N_1720,In_34,In_1482);
xnor U1721 (N_1721,In_953,In_783);
xnor U1722 (N_1722,In_887,In_1501);
and U1723 (N_1723,In_171,In_526);
xnor U1724 (N_1724,In_1240,In_496);
and U1725 (N_1725,In_280,In_1536);
or U1726 (N_1726,In_928,In_332);
and U1727 (N_1727,In_1737,In_834);
or U1728 (N_1728,In_920,In_1423);
nand U1729 (N_1729,In_1793,In_73);
nor U1730 (N_1730,In_68,In_278);
or U1731 (N_1731,In_1143,In_1107);
xor U1732 (N_1732,In_1001,In_52);
or U1733 (N_1733,In_1003,In_380);
and U1734 (N_1734,In_782,In_598);
and U1735 (N_1735,In_1230,In_970);
nor U1736 (N_1736,In_619,In_552);
nand U1737 (N_1737,In_726,In_1263);
nor U1738 (N_1738,In_571,In_93);
and U1739 (N_1739,In_755,In_332);
nor U1740 (N_1740,In_1844,In_1407);
xor U1741 (N_1741,In_970,In_1981);
xor U1742 (N_1742,In_1502,In_306);
or U1743 (N_1743,In_377,In_1339);
and U1744 (N_1744,In_204,In_1536);
or U1745 (N_1745,In_673,In_230);
nand U1746 (N_1746,In_159,In_1215);
and U1747 (N_1747,In_15,In_666);
or U1748 (N_1748,In_824,In_864);
nand U1749 (N_1749,In_195,In_384);
nor U1750 (N_1750,In_218,In_32);
nor U1751 (N_1751,In_170,In_584);
xnor U1752 (N_1752,In_347,In_1485);
nor U1753 (N_1753,In_1364,In_938);
nand U1754 (N_1754,In_470,In_1913);
and U1755 (N_1755,In_1192,In_1248);
xnor U1756 (N_1756,In_506,In_281);
and U1757 (N_1757,In_567,In_400);
nor U1758 (N_1758,In_1124,In_1331);
nor U1759 (N_1759,In_912,In_200);
nor U1760 (N_1760,In_1567,In_193);
xnor U1761 (N_1761,In_1793,In_1049);
or U1762 (N_1762,In_1667,In_247);
or U1763 (N_1763,In_1134,In_570);
nand U1764 (N_1764,In_345,In_1020);
xor U1765 (N_1765,In_44,In_247);
xnor U1766 (N_1766,In_395,In_103);
nor U1767 (N_1767,In_171,In_1224);
nand U1768 (N_1768,In_1381,In_197);
nor U1769 (N_1769,In_986,In_157);
xor U1770 (N_1770,In_897,In_1843);
xnor U1771 (N_1771,In_99,In_1281);
nor U1772 (N_1772,In_788,In_1252);
xnor U1773 (N_1773,In_486,In_1759);
and U1774 (N_1774,In_348,In_376);
nand U1775 (N_1775,In_1636,In_1681);
xor U1776 (N_1776,In_741,In_1580);
or U1777 (N_1777,In_854,In_1957);
and U1778 (N_1778,In_54,In_290);
or U1779 (N_1779,In_1586,In_1384);
nor U1780 (N_1780,In_1874,In_781);
or U1781 (N_1781,In_1246,In_1390);
xnor U1782 (N_1782,In_111,In_1067);
nand U1783 (N_1783,In_396,In_1295);
nor U1784 (N_1784,In_439,In_684);
xnor U1785 (N_1785,In_1621,In_1986);
nand U1786 (N_1786,In_1564,In_1793);
or U1787 (N_1787,In_1338,In_1378);
nand U1788 (N_1788,In_157,In_411);
or U1789 (N_1789,In_1135,In_1448);
xnor U1790 (N_1790,In_1695,In_926);
and U1791 (N_1791,In_1814,In_843);
or U1792 (N_1792,In_1528,In_1307);
or U1793 (N_1793,In_1241,In_381);
nand U1794 (N_1794,In_793,In_1376);
nor U1795 (N_1795,In_1623,In_1322);
or U1796 (N_1796,In_1333,In_31);
and U1797 (N_1797,In_853,In_1811);
xnor U1798 (N_1798,In_1595,In_149);
nand U1799 (N_1799,In_615,In_578);
or U1800 (N_1800,In_1292,In_1852);
xor U1801 (N_1801,In_1675,In_745);
or U1802 (N_1802,In_1564,In_1201);
and U1803 (N_1803,In_1079,In_1817);
xnor U1804 (N_1804,In_1298,In_1754);
nand U1805 (N_1805,In_1060,In_697);
xnor U1806 (N_1806,In_412,In_387);
or U1807 (N_1807,In_1226,In_1146);
xnor U1808 (N_1808,In_1398,In_1480);
nor U1809 (N_1809,In_945,In_247);
nand U1810 (N_1810,In_503,In_1701);
nor U1811 (N_1811,In_1090,In_237);
xnor U1812 (N_1812,In_1956,In_33);
or U1813 (N_1813,In_1393,In_1027);
nand U1814 (N_1814,In_1538,In_1164);
xnor U1815 (N_1815,In_412,In_1639);
nor U1816 (N_1816,In_1007,In_879);
xor U1817 (N_1817,In_1194,In_1040);
xor U1818 (N_1818,In_971,In_566);
nor U1819 (N_1819,In_770,In_1174);
nor U1820 (N_1820,In_765,In_527);
nor U1821 (N_1821,In_350,In_1194);
nor U1822 (N_1822,In_1758,In_749);
xnor U1823 (N_1823,In_502,In_991);
and U1824 (N_1824,In_422,In_1332);
nor U1825 (N_1825,In_97,In_637);
nand U1826 (N_1826,In_1093,In_1293);
or U1827 (N_1827,In_1438,In_1284);
nand U1828 (N_1828,In_1189,In_1467);
or U1829 (N_1829,In_155,In_136);
nor U1830 (N_1830,In_1475,In_1389);
or U1831 (N_1831,In_1845,In_1022);
xnor U1832 (N_1832,In_826,In_703);
nand U1833 (N_1833,In_1754,In_1979);
nor U1834 (N_1834,In_57,In_268);
or U1835 (N_1835,In_994,In_166);
or U1836 (N_1836,In_831,In_335);
nor U1837 (N_1837,In_1196,In_1659);
and U1838 (N_1838,In_102,In_72);
xnor U1839 (N_1839,In_1718,In_1675);
nor U1840 (N_1840,In_1161,In_330);
and U1841 (N_1841,In_1809,In_1191);
xnor U1842 (N_1842,In_1519,In_759);
nor U1843 (N_1843,In_967,In_444);
and U1844 (N_1844,In_1693,In_1054);
nor U1845 (N_1845,In_1399,In_903);
and U1846 (N_1846,In_843,In_246);
nor U1847 (N_1847,In_867,In_1693);
or U1848 (N_1848,In_4,In_1127);
nor U1849 (N_1849,In_1384,In_1755);
nor U1850 (N_1850,In_957,In_1530);
xor U1851 (N_1851,In_848,In_383);
or U1852 (N_1852,In_409,In_193);
nand U1853 (N_1853,In_55,In_952);
or U1854 (N_1854,In_1415,In_1206);
nor U1855 (N_1855,In_855,In_1843);
nor U1856 (N_1856,In_1401,In_879);
nor U1857 (N_1857,In_1484,In_502);
nor U1858 (N_1858,In_1139,In_1094);
or U1859 (N_1859,In_1429,In_462);
and U1860 (N_1860,In_1263,In_1168);
xnor U1861 (N_1861,In_280,In_15);
xor U1862 (N_1862,In_404,In_695);
or U1863 (N_1863,In_113,In_168);
nand U1864 (N_1864,In_977,In_1478);
nand U1865 (N_1865,In_636,In_368);
and U1866 (N_1866,In_1497,In_781);
nor U1867 (N_1867,In_1132,In_1553);
xor U1868 (N_1868,In_650,In_1801);
and U1869 (N_1869,In_241,In_1457);
and U1870 (N_1870,In_1332,In_298);
nand U1871 (N_1871,In_1389,In_1293);
xor U1872 (N_1872,In_1220,In_1920);
nor U1873 (N_1873,In_1563,In_639);
or U1874 (N_1874,In_927,In_405);
and U1875 (N_1875,In_182,In_1843);
nand U1876 (N_1876,In_1290,In_1962);
or U1877 (N_1877,In_1057,In_841);
or U1878 (N_1878,In_288,In_1193);
and U1879 (N_1879,In_1331,In_735);
nand U1880 (N_1880,In_1454,In_457);
and U1881 (N_1881,In_1317,In_1669);
or U1882 (N_1882,In_1594,In_449);
or U1883 (N_1883,In_368,In_1995);
xnor U1884 (N_1884,In_64,In_111);
and U1885 (N_1885,In_1522,In_62);
nor U1886 (N_1886,In_121,In_1498);
xnor U1887 (N_1887,In_343,In_45);
xor U1888 (N_1888,In_836,In_309);
xnor U1889 (N_1889,In_1677,In_1993);
nor U1890 (N_1890,In_1941,In_1854);
or U1891 (N_1891,In_701,In_1832);
xor U1892 (N_1892,In_1610,In_468);
xor U1893 (N_1893,In_1583,In_1085);
nor U1894 (N_1894,In_866,In_583);
nor U1895 (N_1895,In_387,In_1425);
and U1896 (N_1896,In_702,In_548);
nor U1897 (N_1897,In_494,In_1684);
xor U1898 (N_1898,In_134,In_1654);
nor U1899 (N_1899,In_309,In_1778);
and U1900 (N_1900,In_1243,In_1472);
nor U1901 (N_1901,In_531,In_595);
xnor U1902 (N_1902,In_843,In_1474);
and U1903 (N_1903,In_1709,In_1692);
nand U1904 (N_1904,In_479,In_1711);
nand U1905 (N_1905,In_1106,In_1155);
nand U1906 (N_1906,In_700,In_175);
or U1907 (N_1907,In_863,In_739);
or U1908 (N_1908,In_411,In_1752);
or U1909 (N_1909,In_262,In_104);
nor U1910 (N_1910,In_992,In_1265);
and U1911 (N_1911,In_1720,In_846);
xor U1912 (N_1912,In_1442,In_1852);
xor U1913 (N_1913,In_1108,In_1627);
or U1914 (N_1914,In_512,In_823);
nand U1915 (N_1915,In_657,In_1359);
nand U1916 (N_1916,In_1618,In_41);
nand U1917 (N_1917,In_933,In_178);
or U1918 (N_1918,In_314,In_319);
xor U1919 (N_1919,In_1167,In_990);
and U1920 (N_1920,In_218,In_354);
nor U1921 (N_1921,In_1956,In_27);
and U1922 (N_1922,In_1363,In_1460);
and U1923 (N_1923,In_1398,In_931);
and U1924 (N_1924,In_1518,In_1172);
nand U1925 (N_1925,In_891,In_721);
nand U1926 (N_1926,In_1387,In_1628);
nor U1927 (N_1927,In_289,In_1715);
nand U1928 (N_1928,In_1072,In_1145);
nor U1929 (N_1929,In_92,In_1873);
and U1930 (N_1930,In_1068,In_932);
or U1931 (N_1931,In_1890,In_500);
nand U1932 (N_1932,In_1615,In_1809);
or U1933 (N_1933,In_1777,In_28);
or U1934 (N_1934,In_652,In_1722);
and U1935 (N_1935,In_91,In_1331);
or U1936 (N_1936,In_278,In_442);
and U1937 (N_1937,In_1448,In_1198);
and U1938 (N_1938,In_396,In_1548);
or U1939 (N_1939,In_1085,In_487);
nand U1940 (N_1940,In_1410,In_514);
nor U1941 (N_1941,In_1215,In_1571);
xor U1942 (N_1942,In_1205,In_746);
xnor U1943 (N_1943,In_1931,In_1889);
nand U1944 (N_1944,In_1063,In_589);
xnor U1945 (N_1945,In_1063,In_1157);
xnor U1946 (N_1946,In_1745,In_1159);
nand U1947 (N_1947,In_1707,In_310);
and U1948 (N_1948,In_857,In_12);
or U1949 (N_1949,In_1419,In_180);
nand U1950 (N_1950,In_1562,In_1269);
and U1951 (N_1951,In_518,In_154);
nor U1952 (N_1952,In_1602,In_204);
nor U1953 (N_1953,In_1936,In_694);
nor U1954 (N_1954,In_431,In_1285);
or U1955 (N_1955,In_363,In_1140);
and U1956 (N_1956,In_816,In_1557);
xor U1957 (N_1957,In_682,In_1259);
and U1958 (N_1958,In_324,In_1453);
xnor U1959 (N_1959,In_267,In_1366);
or U1960 (N_1960,In_1928,In_372);
nor U1961 (N_1961,In_1061,In_665);
and U1962 (N_1962,In_975,In_1475);
or U1963 (N_1963,In_1558,In_1652);
nand U1964 (N_1964,In_164,In_26);
nor U1965 (N_1965,In_882,In_257);
or U1966 (N_1966,In_1911,In_1656);
nand U1967 (N_1967,In_758,In_666);
nor U1968 (N_1968,In_1041,In_1746);
or U1969 (N_1969,In_189,In_1295);
xor U1970 (N_1970,In_1932,In_147);
or U1971 (N_1971,In_1300,In_276);
or U1972 (N_1972,In_1045,In_115);
and U1973 (N_1973,In_1668,In_907);
nand U1974 (N_1974,In_421,In_1934);
or U1975 (N_1975,In_283,In_1488);
nor U1976 (N_1976,In_646,In_315);
nand U1977 (N_1977,In_1523,In_1685);
nand U1978 (N_1978,In_1942,In_844);
nor U1979 (N_1979,In_968,In_1504);
xnor U1980 (N_1980,In_1338,In_1789);
nand U1981 (N_1981,In_822,In_382);
and U1982 (N_1982,In_1832,In_1363);
nor U1983 (N_1983,In_38,In_1421);
nor U1984 (N_1984,In_352,In_180);
or U1985 (N_1985,In_1860,In_1456);
nor U1986 (N_1986,In_751,In_436);
nor U1987 (N_1987,In_1400,In_337);
or U1988 (N_1988,In_1187,In_775);
or U1989 (N_1989,In_1529,In_935);
xnor U1990 (N_1990,In_134,In_1364);
xor U1991 (N_1991,In_15,In_634);
and U1992 (N_1992,In_1683,In_832);
nor U1993 (N_1993,In_1728,In_43);
xnor U1994 (N_1994,In_607,In_1657);
nand U1995 (N_1995,In_1981,In_1326);
nor U1996 (N_1996,In_1456,In_272);
or U1997 (N_1997,In_1696,In_1739);
or U1998 (N_1998,In_1055,In_1748);
nor U1999 (N_1999,In_709,In_1018);
xnor U2000 (N_2000,In_556,In_1946);
nor U2001 (N_2001,In_27,In_1477);
and U2002 (N_2002,In_34,In_401);
or U2003 (N_2003,In_1152,In_497);
or U2004 (N_2004,In_1955,In_231);
nand U2005 (N_2005,In_869,In_1471);
or U2006 (N_2006,In_980,In_1801);
or U2007 (N_2007,In_1698,In_1821);
nand U2008 (N_2008,In_1689,In_1151);
nand U2009 (N_2009,In_663,In_1816);
xnor U2010 (N_2010,In_236,In_437);
xnor U2011 (N_2011,In_511,In_512);
nor U2012 (N_2012,In_1425,In_1786);
nand U2013 (N_2013,In_1139,In_184);
and U2014 (N_2014,In_304,In_553);
or U2015 (N_2015,In_1817,In_1984);
xnor U2016 (N_2016,In_41,In_1306);
nor U2017 (N_2017,In_645,In_1914);
or U2018 (N_2018,In_1991,In_1498);
xnor U2019 (N_2019,In_1514,In_778);
nand U2020 (N_2020,In_1004,In_568);
nand U2021 (N_2021,In_1658,In_1623);
nand U2022 (N_2022,In_1616,In_889);
xnor U2023 (N_2023,In_1163,In_713);
or U2024 (N_2024,In_1699,In_1979);
or U2025 (N_2025,In_1247,In_389);
and U2026 (N_2026,In_1125,In_431);
or U2027 (N_2027,In_1725,In_78);
xnor U2028 (N_2028,In_1485,In_1379);
and U2029 (N_2029,In_637,In_1758);
nor U2030 (N_2030,In_55,In_919);
nand U2031 (N_2031,In_227,In_1088);
xor U2032 (N_2032,In_874,In_61);
nand U2033 (N_2033,In_1860,In_125);
and U2034 (N_2034,In_1178,In_1980);
xnor U2035 (N_2035,In_599,In_992);
nand U2036 (N_2036,In_294,In_1707);
and U2037 (N_2037,In_886,In_200);
and U2038 (N_2038,In_456,In_1338);
xnor U2039 (N_2039,In_1743,In_1651);
or U2040 (N_2040,In_1844,In_1226);
nor U2041 (N_2041,In_602,In_991);
nor U2042 (N_2042,In_596,In_1600);
and U2043 (N_2043,In_994,In_1499);
nor U2044 (N_2044,In_787,In_1111);
xor U2045 (N_2045,In_690,In_410);
and U2046 (N_2046,In_55,In_132);
and U2047 (N_2047,In_489,In_975);
nor U2048 (N_2048,In_1316,In_1802);
nand U2049 (N_2049,In_207,In_1276);
or U2050 (N_2050,In_1225,In_1713);
nor U2051 (N_2051,In_118,In_1940);
nand U2052 (N_2052,In_1013,In_933);
nor U2053 (N_2053,In_890,In_1085);
xnor U2054 (N_2054,In_1987,In_1173);
or U2055 (N_2055,In_195,In_438);
nor U2056 (N_2056,In_135,In_572);
or U2057 (N_2057,In_1798,In_1145);
xor U2058 (N_2058,In_1414,In_284);
nand U2059 (N_2059,In_483,In_80);
and U2060 (N_2060,In_1350,In_1209);
or U2061 (N_2061,In_1843,In_1087);
nand U2062 (N_2062,In_338,In_1053);
nand U2063 (N_2063,In_569,In_1690);
nor U2064 (N_2064,In_1767,In_845);
nand U2065 (N_2065,In_1442,In_1174);
or U2066 (N_2066,In_1664,In_1867);
or U2067 (N_2067,In_547,In_1522);
and U2068 (N_2068,In_1550,In_680);
xnor U2069 (N_2069,In_359,In_1496);
nand U2070 (N_2070,In_612,In_631);
nor U2071 (N_2071,In_1647,In_273);
or U2072 (N_2072,In_1534,In_139);
xnor U2073 (N_2073,In_659,In_439);
and U2074 (N_2074,In_196,In_1819);
or U2075 (N_2075,In_427,In_261);
nor U2076 (N_2076,In_761,In_1839);
or U2077 (N_2077,In_1278,In_1245);
nand U2078 (N_2078,In_339,In_1732);
nor U2079 (N_2079,In_1853,In_1779);
xnor U2080 (N_2080,In_1941,In_1689);
xnor U2081 (N_2081,In_1949,In_1999);
nor U2082 (N_2082,In_1478,In_755);
xor U2083 (N_2083,In_569,In_434);
xnor U2084 (N_2084,In_206,In_298);
and U2085 (N_2085,In_1810,In_1524);
nand U2086 (N_2086,In_241,In_475);
and U2087 (N_2087,In_332,In_1753);
and U2088 (N_2088,In_1293,In_1505);
xor U2089 (N_2089,In_381,In_582);
or U2090 (N_2090,In_1940,In_1407);
xor U2091 (N_2091,In_1370,In_1035);
nand U2092 (N_2092,In_1652,In_338);
nand U2093 (N_2093,In_1102,In_1882);
and U2094 (N_2094,In_599,In_820);
xnor U2095 (N_2095,In_1826,In_1809);
xor U2096 (N_2096,In_1468,In_1279);
xor U2097 (N_2097,In_1284,In_1080);
or U2098 (N_2098,In_549,In_1195);
xnor U2099 (N_2099,In_830,In_1045);
xor U2100 (N_2100,In_656,In_988);
or U2101 (N_2101,In_1741,In_1983);
or U2102 (N_2102,In_74,In_1889);
and U2103 (N_2103,In_281,In_403);
nor U2104 (N_2104,In_1441,In_65);
nor U2105 (N_2105,In_1320,In_157);
and U2106 (N_2106,In_744,In_974);
and U2107 (N_2107,In_177,In_523);
nand U2108 (N_2108,In_1230,In_907);
and U2109 (N_2109,In_1996,In_509);
xor U2110 (N_2110,In_1804,In_1856);
nor U2111 (N_2111,In_1648,In_351);
nor U2112 (N_2112,In_1589,In_1295);
nand U2113 (N_2113,In_845,In_944);
and U2114 (N_2114,In_1803,In_900);
nand U2115 (N_2115,In_1199,In_401);
or U2116 (N_2116,In_943,In_1721);
xor U2117 (N_2117,In_1628,In_969);
and U2118 (N_2118,In_1429,In_1203);
or U2119 (N_2119,In_1861,In_1509);
and U2120 (N_2120,In_1021,In_1669);
xnor U2121 (N_2121,In_1559,In_1741);
xor U2122 (N_2122,In_1614,In_1117);
nand U2123 (N_2123,In_172,In_323);
nor U2124 (N_2124,In_1303,In_503);
xnor U2125 (N_2125,In_1498,In_1762);
xor U2126 (N_2126,In_1341,In_5);
and U2127 (N_2127,In_1032,In_1982);
xnor U2128 (N_2128,In_184,In_1830);
and U2129 (N_2129,In_482,In_283);
or U2130 (N_2130,In_1850,In_241);
or U2131 (N_2131,In_1227,In_551);
nor U2132 (N_2132,In_1574,In_1359);
and U2133 (N_2133,In_1200,In_706);
and U2134 (N_2134,In_252,In_1454);
and U2135 (N_2135,In_883,In_1930);
nor U2136 (N_2136,In_1210,In_1922);
nand U2137 (N_2137,In_938,In_536);
nor U2138 (N_2138,In_749,In_1226);
or U2139 (N_2139,In_981,In_971);
or U2140 (N_2140,In_141,In_688);
nor U2141 (N_2141,In_1081,In_1428);
or U2142 (N_2142,In_612,In_1918);
and U2143 (N_2143,In_407,In_1889);
and U2144 (N_2144,In_336,In_237);
xnor U2145 (N_2145,In_1805,In_1936);
nor U2146 (N_2146,In_1601,In_605);
and U2147 (N_2147,In_1791,In_1851);
xnor U2148 (N_2148,In_1950,In_330);
and U2149 (N_2149,In_1358,In_1838);
nand U2150 (N_2150,In_971,In_1276);
and U2151 (N_2151,In_121,In_2);
xnor U2152 (N_2152,In_889,In_1612);
xnor U2153 (N_2153,In_229,In_1795);
xnor U2154 (N_2154,In_1475,In_870);
xnor U2155 (N_2155,In_1705,In_1479);
xnor U2156 (N_2156,In_1869,In_1458);
nor U2157 (N_2157,In_673,In_700);
or U2158 (N_2158,In_581,In_346);
nand U2159 (N_2159,In_1637,In_452);
nand U2160 (N_2160,In_1086,In_1970);
or U2161 (N_2161,In_1645,In_1695);
nor U2162 (N_2162,In_1981,In_1432);
nor U2163 (N_2163,In_1904,In_1635);
nand U2164 (N_2164,In_194,In_1131);
or U2165 (N_2165,In_1456,In_192);
or U2166 (N_2166,In_1579,In_1183);
nor U2167 (N_2167,In_673,In_642);
nor U2168 (N_2168,In_1841,In_64);
nor U2169 (N_2169,In_350,In_1660);
or U2170 (N_2170,In_1243,In_844);
nand U2171 (N_2171,In_1960,In_336);
xnor U2172 (N_2172,In_458,In_839);
or U2173 (N_2173,In_771,In_1758);
xnor U2174 (N_2174,In_1557,In_975);
and U2175 (N_2175,In_1689,In_1668);
nor U2176 (N_2176,In_1432,In_1657);
xor U2177 (N_2177,In_230,In_1284);
nand U2178 (N_2178,In_1293,In_1435);
xor U2179 (N_2179,In_686,In_1788);
nor U2180 (N_2180,In_147,In_1962);
or U2181 (N_2181,In_579,In_1423);
and U2182 (N_2182,In_405,In_18);
and U2183 (N_2183,In_420,In_1992);
xor U2184 (N_2184,In_1720,In_307);
or U2185 (N_2185,In_89,In_404);
nand U2186 (N_2186,In_735,In_1478);
xor U2187 (N_2187,In_1971,In_496);
or U2188 (N_2188,In_1018,In_1609);
or U2189 (N_2189,In_937,In_1667);
nor U2190 (N_2190,In_1149,In_1270);
or U2191 (N_2191,In_1968,In_204);
and U2192 (N_2192,In_530,In_871);
nand U2193 (N_2193,In_1705,In_959);
or U2194 (N_2194,In_249,In_285);
or U2195 (N_2195,In_1960,In_1707);
and U2196 (N_2196,In_1718,In_1598);
xnor U2197 (N_2197,In_1981,In_587);
nor U2198 (N_2198,In_74,In_507);
nor U2199 (N_2199,In_553,In_1947);
nor U2200 (N_2200,In_1018,In_1772);
and U2201 (N_2201,In_138,In_1218);
xor U2202 (N_2202,In_1443,In_682);
xnor U2203 (N_2203,In_772,In_1172);
and U2204 (N_2204,In_288,In_1908);
and U2205 (N_2205,In_83,In_687);
nor U2206 (N_2206,In_366,In_993);
or U2207 (N_2207,In_514,In_1571);
and U2208 (N_2208,In_600,In_1328);
nand U2209 (N_2209,In_1392,In_869);
xor U2210 (N_2210,In_320,In_1592);
nor U2211 (N_2211,In_506,In_1643);
nor U2212 (N_2212,In_1886,In_1033);
and U2213 (N_2213,In_1090,In_807);
nand U2214 (N_2214,In_1161,In_1237);
or U2215 (N_2215,In_605,In_392);
or U2216 (N_2216,In_1773,In_932);
and U2217 (N_2217,In_1960,In_807);
or U2218 (N_2218,In_606,In_259);
and U2219 (N_2219,In_1327,In_1683);
nor U2220 (N_2220,In_1476,In_474);
or U2221 (N_2221,In_682,In_931);
nand U2222 (N_2222,In_34,In_1976);
and U2223 (N_2223,In_277,In_151);
xor U2224 (N_2224,In_146,In_1919);
or U2225 (N_2225,In_930,In_627);
xor U2226 (N_2226,In_1157,In_1935);
or U2227 (N_2227,In_1013,In_962);
or U2228 (N_2228,In_1715,In_347);
or U2229 (N_2229,In_1999,In_710);
and U2230 (N_2230,In_1449,In_504);
nor U2231 (N_2231,In_1955,In_1734);
nor U2232 (N_2232,In_203,In_703);
or U2233 (N_2233,In_1711,In_413);
xnor U2234 (N_2234,In_1404,In_55);
xor U2235 (N_2235,In_506,In_425);
nand U2236 (N_2236,In_1725,In_217);
nor U2237 (N_2237,In_1197,In_1641);
nand U2238 (N_2238,In_374,In_728);
or U2239 (N_2239,In_1680,In_1037);
nand U2240 (N_2240,In_1348,In_1272);
nor U2241 (N_2241,In_863,In_1235);
nor U2242 (N_2242,In_1303,In_298);
nor U2243 (N_2243,In_625,In_929);
or U2244 (N_2244,In_1982,In_1192);
and U2245 (N_2245,In_1206,In_383);
and U2246 (N_2246,In_463,In_1626);
or U2247 (N_2247,In_952,In_355);
or U2248 (N_2248,In_637,In_738);
or U2249 (N_2249,In_1617,In_836);
nor U2250 (N_2250,In_512,In_1536);
nor U2251 (N_2251,In_199,In_717);
nand U2252 (N_2252,In_1136,In_1974);
or U2253 (N_2253,In_967,In_1748);
nor U2254 (N_2254,In_763,In_496);
xor U2255 (N_2255,In_607,In_1105);
xnor U2256 (N_2256,In_18,In_1199);
or U2257 (N_2257,In_1948,In_917);
or U2258 (N_2258,In_1087,In_1418);
xnor U2259 (N_2259,In_220,In_1238);
or U2260 (N_2260,In_136,In_1722);
or U2261 (N_2261,In_1966,In_1780);
nor U2262 (N_2262,In_374,In_511);
or U2263 (N_2263,In_972,In_1686);
nor U2264 (N_2264,In_1340,In_721);
and U2265 (N_2265,In_1541,In_1940);
nand U2266 (N_2266,In_1080,In_589);
and U2267 (N_2267,In_1383,In_367);
nand U2268 (N_2268,In_436,In_1057);
and U2269 (N_2269,In_1904,In_1908);
or U2270 (N_2270,In_1854,In_119);
xor U2271 (N_2271,In_664,In_1886);
xor U2272 (N_2272,In_719,In_1064);
xnor U2273 (N_2273,In_1467,In_660);
and U2274 (N_2274,In_1760,In_74);
and U2275 (N_2275,In_1950,In_96);
or U2276 (N_2276,In_1199,In_1103);
or U2277 (N_2277,In_1466,In_626);
xnor U2278 (N_2278,In_1791,In_206);
or U2279 (N_2279,In_7,In_735);
and U2280 (N_2280,In_481,In_66);
nand U2281 (N_2281,In_1455,In_666);
and U2282 (N_2282,In_1924,In_1815);
xnor U2283 (N_2283,In_1591,In_859);
and U2284 (N_2284,In_1757,In_45);
nor U2285 (N_2285,In_160,In_583);
or U2286 (N_2286,In_187,In_129);
and U2287 (N_2287,In_1559,In_654);
nand U2288 (N_2288,In_646,In_57);
and U2289 (N_2289,In_392,In_536);
nor U2290 (N_2290,In_1101,In_1803);
and U2291 (N_2291,In_957,In_1595);
nand U2292 (N_2292,In_680,In_160);
and U2293 (N_2293,In_713,In_1950);
nand U2294 (N_2294,In_436,In_1946);
xor U2295 (N_2295,In_97,In_366);
and U2296 (N_2296,In_890,In_414);
nor U2297 (N_2297,In_884,In_1879);
nor U2298 (N_2298,In_1188,In_182);
nor U2299 (N_2299,In_1344,In_1102);
nor U2300 (N_2300,In_1114,In_1811);
nor U2301 (N_2301,In_463,In_1527);
nand U2302 (N_2302,In_1741,In_1308);
or U2303 (N_2303,In_496,In_34);
or U2304 (N_2304,In_1390,In_1552);
or U2305 (N_2305,In_1771,In_1419);
or U2306 (N_2306,In_1749,In_1541);
xor U2307 (N_2307,In_1007,In_785);
nand U2308 (N_2308,In_888,In_774);
nor U2309 (N_2309,In_673,In_1999);
nor U2310 (N_2310,In_188,In_1161);
and U2311 (N_2311,In_665,In_849);
and U2312 (N_2312,In_1519,In_140);
nor U2313 (N_2313,In_806,In_602);
nand U2314 (N_2314,In_519,In_1288);
nor U2315 (N_2315,In_1095,In_1438);
and U2316 (N_2316,In_1338,In_508);
or U2317 (N_2317,In_980,In_1465);
nand U2318 (N_2318,In_1006,In_1418);
xnor U2319 (N_2319,In_1317,In_1935);
or U2320 (N_2320,In_1405,In_1246);
xor U2321 (N_2321,In_1904,In_1711);
nand U2322 (N_2322,In_840,In_317);
nand U2323 (N_2323,In_425,In_1682);
nor U2324 (N_2324,In_476,In_1480);
and U2325 (N_2325,In_607,In_1966);
and U2326 (N_2326,In_484,In_669);
and U2327 (N_2327,In_53,In_1181);
nand U2328 (N_2328,In_1520,In_1507);
xor U2329 (N_2329,In_1418,In_1692);
nand U2330 (N_2330,In_486,In_237);
nor U2331 (N_2331,In_871,In_4);
nand U2332 (N_2332,In_1890,In_44);
nor U2333 (N_2333,In_1480,In_500);
nor U2334 (N_2334,In_434,In_1931);
xnor U2335 (N_2335,In_1122,In_856);
nor U2336 (N_2336,In_558,In_1821);
nand U2337 (N_2337,In_132,In_1320);
and U2338 (N_2338,In_1030,In_832);
nor U2339 (N_2339,In_910,In_1415);
and U2340 (N_2340,In_1039,In_356);
xor U2341 (N_2341,In_1055,In_154);
nand U2342 (N_2342,In_1327,In_809);
and U2343 (N_2343,In_1022,In_1185);
nand U2344 (N_2344,In_468,In_1534);
or U2345 (N_2345,In_1153,In_1048);
xor U2346 (N_2346,In_1088,In_890);
and U2347 (N_2347,In_592,In_78);
and U2348 (N_2348,In_850,In_879);
nor U2349 (N_2349,In_1474,In_1393);
or U2350 (N_2350,In_287,In_460);
xor U2351 (N_2351,In_1238,In_1016);
and U2352 (N_2352,In_1838,In_1948);
xnor U2353 (N_2353,In_1500,In_1228);
nand U2354 (N_2354,In_1016,In_1999);
nor U2355 (N_2355,In_434,In_211);
nor U2356 (N_2356,In_835,In_190);
and U2357 (N_2357,In_1233,In_397);
and U2358 (N_2358,In_867,In_921);
nand U2359 (N_2359,In_1720,In_239);
or U2360 (N_2360,In_1045,In_1921);
and U2361 (N_2361,In_1066,In_395);
nor U2362 (N_2362,In_1346,In_1754);
nand U2363 (N_2363,In_1983,In_1880);
nand U2364 (N_2364,In_664,In_1436);
nor U2365 (N_2365,In_920,In_1160);
nand U2366 (N_2366,In_890,In_525);
or U2367 (N_2367,In_108,In_194);
and U2368 (N_2368,In_236,In_382);
nand U2369 (N_2369,In_1036,In_1910);
nand U2370 (N_2370,In_368,In_1055);
nand U2371 (N_2371,In_1118,In_1173);
and U2372 (N_2372,In_81,In_1242);
nand U2373 (N_2373,In_1869,In_699);
nor U2374 (N_2374,In_1786,In_489);
or U2375 (N_2375,In_1271,In_387);
or U2376 (N_2376,In_676,In_67);
nand U2377 (N_2377,In_1430,In_1509);
nor U2378 (N_2378,In_1682,In_675);
nand U2379 (N_2379,In_1057,In_1511);
xnor U2380 (N_2380,In_122,In_807);
nor U2381 (N_2381,In_209,In_1297);
nor U2382 (N_2382,In_757,In_265);
and U2383 (N_2383,In_946,In_1605);
nand U2384 (N_2384,In_386,In_1047);
nor U2385 (N_2385,In_28,In_1196);
or U2386 (N_2386,In_479,In_1389);
and U2387 (N_2387,In_477,In_1610);
and U2388 (N_2388,In_693,In_434);
and U2389 (N_2389,In_625,In_1500);
nand U2390 (N_2390,In_445,In_572);
nor U2391 (N_2391,In_1251,In_280);
nand U2392 (N_2392,In_1916,In_891);
xnor U2393 (N_2393,In_1827,In_1191);
nand U2394 (N_2394,In_1821,In_220);
nor U2395 (N_2395,In_1129,In_826);
and U2396 (N_2396,In_1512,In_618);
xnor U2397 (N_2397,In_190,In_194);
or U2398 (N_2398,In_422,In_1689);
or U2399 (N_2399,In_1172,In_809);
nor U2400 (N_2400,In_848,In_187);
or U2401 (N_2401,In_1487,In_291);
or U2402 (N_2402,In_1223,In_367);
and U2403 (N_2403,In_1181,In_1399);
and U2404 (N_2404,In_1791,In_1775);
and U2405 (N_2405,In_1526,In_1398);
nor U2406 (N_2406,In_299,In_574);
nor U2407 (N_2407,In_288,In_1460);
nor U2408 (N_2408,In_178,In_1517);
and U2409 (N_2409,In_512,In_1393);
nand U2410 (N_2410,In_1420,In_1913);
or U2411 (N_2411,In_1283,In_994);
nor U2412 (N_2412,In_626,In_855);
and U2413 (N_2413,In_99,In_970);
and U2414 (N_2414,In_263,In_685);
nor U2415 (N_2415,In_699,In_441);
nand U2416 (N_2416,In_1687,In_279);
nor U2417 (N_2417,In_629,In_255);
nor U2418 (N_2418,In_1486,In_1102);
xor U2419 (N_2419,In_678,In_1958);
nand U2420 (N_2420,In_139,In_1702);
or U2421 (N_2421,In_1429,In_1910);
and U2422 (N_2422,In_358,In_118);
or U2423 (N_2423,In_324,In_1019);
or U2424 (N_2424,In_295,In_1195);
and U2425 (N_2425,In_985,In_1639);
nand U2426 (N_2426,In_1832,In_184);
or U2427 (N_2427,In_1955,In_117);
nor U2428 (N_2428,In_664,In_734);
nand U2429 (N_2429,In_199,In_72);
nor U2430 (N_2430,In_1261,In_550);
or U2431 (N_2431,In_1282,In_55);
or U2432 (N_2432,In_130,In_1082);
nand U2433 (N_2433,In_1336,In_572);
xor U2434 (N_2434,In_787,In_781);
and U2435 (N_2435,In_697,In_681);
and U2436 (N_2436,In_1378,In_692);
or U2437 (N_2437,In_51,In_1969);
nand U2438 (N_2438,In_409,In_280);
and U2439 (N_2439,In_335,In_1665);
xnor U2440 (N_2440,In_601,In_1304);
nor U2441 (N_2441,In_1822,In_839);
or U2442 (N_2442,In_174,In_217);
and U2443 (N_2443,In_178,In_1411);
or U2444 (N_2444,In_1580,In_670);
xor U2445 (N_2445,In_1906,In_1359);
nor U2446 (N_2446,In_1354,In_494);
xnor U2447 (N_2447,In_624,In_586);
and U2448 (N_2448,In_1885,In_1387);
and U2449 (N_2449,In_839,In_347);
nand U2450 (N_2450,In_1308,In_1621);
xor U2451 (N_2451,In_1706,In_1891);
xnor U2452 (N_2452,In_1638,In_620);
xor U2453 (N_2453,In_90,In_263);
or U2454 (N_2454,In_1494,In_196);
and U2455 (N_2455,In_82,In_747);
nand U2456 (N_2456,In_374,In_585);
xor U2457 (N_2457,In_944,In_1046);
nand U2458 (N_2458,In_181,In_106);
xnor U2459 (N_2459,In_1349,In_1668);
and U2460 (N_2460,In_1669,In_1385);
nand U2461 (N_2461,In_1607,In_682);
xor U2462 (N_2462,In_107,In_1879);
nand U2463 (N_2463,In_1336,In_1330);
nand U2464 (N_2464,In_903,In_169);
and U2465 (N_2465,In_839,In_1196);
nand U2466 (N_2466,In_1698,In_439);
and U2467 (N_2467,In_910,In_1445);
and U2468 (N_2468,In_505,In_1881);
and U2469 (N_2469,In_629,In_1351);
nand U2470 (N_2470,In_976,In_1938);
nor U2471 (N_2471,In_1231,In_1380);
and U2472 (N_2472,In_775,In_982);
or U2473 (N_2473,In_1129,In_76);
and U2474 (N_2474,In_322,In_263);
xor U2475 (N_2475,In_501,In_817);
and U2476 (N_2476,In_661,In_965);
xnor U2477 (N_2477,In_1837,In_236);
and U2478 (N_2478,In_1292,In_767);
xnor U2479 (N_2479,In_1074,In_1686);
nand U2480 (N_2480,In_736,In_230);
nand U2481 (N_2481,In_1308,In_724);
or U2482 (N_2482,In_1982,In_729);
nand U2483 (N_2483,In_767,In_532);
and U2484 (N_2484,In_950,In_1830);
or U2485 (N_2485,In_655,In_1388);
or U2486 (N_2486,In_171,In_1926);
nand U2487 (N_2487,In_1652,In_46);
and U2488 (N_2488,In_1857,In_303);
or U2489 (N_2489,In_908,In_719);
nor U2490 (N_2490,In_894,In_145);
xor U2491 (N_2491,In_1233,In_1020);
and U2492 (N_2492,In_821,In_369);
nand U2493 (N_2493,In_1536,In_35);
nand U2494 (N_2494,In_565,In_1503);
xor U2495 (N_2495,In_1545,In_747);
nand U2496 (N_2496,In_1908,In_503);
xnor U2497 (N_2497,In_956,In_1839);
nand U2498 (N_2498,In_454,In_1553);
nor U2499 (N_2499,In_1174,In_1547);
or U2500 (N_2500,In_1552,In_1046);
and U2501 (N_2501,In_1773,In_628);
nor U2502 (N_2502,In_1382,In_1838);
xnor U2503 (N_2503,In_1847,In_1326);
nor U2504 (N_2504,In_1298,In_894);
and U2505 (N_2505,In_467,In_1);
xnor U2506 (N_2506,In_787,In_1291);
and U2507 (N_2507,In_179,In_1176);
xnor U2508 (N_2508,In_494,In_498);
nor U2509 (N_2509,In_890,In_1283);
and U2510 (N_2510,In_1346,In_436);
nand U2511 (N_2511,In_1051,In_649);
and U2512 (N_2512,In_70,In_385);
nand U2513 (N_2513,In_169,In_1504);
nand U2514 (N_2514,In_1115,In_1908);
nand U2515 (N_2515,In_662,In_536);
xnor U2516 (N_2516,In_573,In_1230);
and U2517 (N_2517,In_401,In_1075);
nand U2518 (N_2518,In_118,In_1435);
xor U2519 (N_2519,In_1078,In_1433);
or U2520 (N_2520,In_524,In_1670);
nand U2521 (N_2521,In_645,In_1267);
xor U2522 (N_2522,In_1488,In_717);
nor U2523 (N_2523,In_674,In_1344);
or U2524 (N_2524,In_1853,In_531);
xor U2525 (N_2525,In_52,In_244);
xor U2526 (N_2526,In_1554,In_1754);
nor U2527 (N_2527,In_282,In_391);
xnor U2528 (N_2528,In_921,In_1934);
and U2529 (N_2529,In_594,In_1866);
nand U2530 (N_2530,In_515,In_1173);
or U2531 (N_2531,In_1057,In_1394);
or U2532 (N_2532,In_1240,In_789);
xor U2533 (N_2533,In_1447,In_267);
xnor U2534 (N_2534,In_1568,In_1096);
nand U2535 (N_2535,In_860,In_1878);
or U2536 (N_2536,In_1163,In_446);
xnor U2537 (N_2537,In_401,In_1332);
and U2538 (N_2538,In_677,In_1135);
and U2539 (N_2539,In_696,In_1200);
nand U2540 (N_2540,In_1781,In_1817);
and U2541 (N_2541,In_736,In_1957);
nor U2542 (N_2542,In_1078,In_956);
and U2543 (N_2543,In_259,In_662);
nor U2544 (N_2544,In_1695,In_131);
nor U2545 (N_2545,In_1165,In_460);
and U2546 (N_2546,In_1618,In_689);
and U2547 (N_2547,In_589,In_563);
nand U2548 (N_2548,In_1352,In_218);
xor U2549 (N_2549,In_629,In_478);
or U2550 (N_2550,In_413,In_455);
nand U2551 (N_2551,In_242,In_1582);
and U2552 (N_2552,In_1270,In_1342);
nor U2553 (N_2553,In_55,In_1432);
nor U2554 (N_2554,In_1705,In_1149);
xnor U2555 (N_2555,In_634,In_477);
xnor U2556 (N_2556,In_1739,In_1842);
and U2557 (N_2557,In_728,In_383);
or U2558 (N_2558,In_1793,In_57);
xnor U2559 (N_2559,In_730,In_485);
and U2560 (N_2560,In_288,In_604);
and U2561 (N_2561,In_845,In_1820);
xor U2562 (N_2562,In_183,In_1833);
nand U2563 (N_2563,In_1351,In_269);
nand U2564 (N_2564,In_230,In_945);
nand U2565 (N_2565,In_1535,In_1002);
xor U2566 (N_2566,In_1035,In_363);
nand U2567 (N_2567,In_727,In_1588);
and U2568 (N_2568,In_1554,In_697);
nor U2569 (N_2569,In_834,In_378);
nor U2570 (N_2570,In_1332,In_1563);
nand U2571 (N_2571,In_1460,In_1837);
and U2572 (N_2572,In_1625,In_1951);
and U2573 (N_2573,In_933,In_1079);
or U2574 (N_2574,In_1440,In_1164);
and U2575 (N_2575,In_336,In_1511);
xor U2576 (N_2576,In_878,In_1529);
and U2577 (N_2577,In_913,In_1877);
nor U2578 (N_2578,In_30,In_155);
nand U2579 (N_2579,In_391,In_455);
or U2580 (N_2580,In_1567,In_409);
or U2581 (N_2581,In_1907,In_748);
and U2582 (N_2582,In_1536,In_1527);
or U2583 (N_2583,In_1347,In_1268);
nand U2584 (N_2584,In_973,In_587);
xor U2585 (N_2585,In_1758,In_633);
xnor U2586 (N_2586,In_395,In_1075);
nand U2587 (N_2587,In_1110,In_632);
nor U2588 (N_2588,In_902,In_8);
or U2589 (N_2589,In_1389,In_397);
nor U2590 (N_2590,In_575,In_123);
nand U2591 (N_2591,In_395,In_773);
and U2592 (N_2592,In_5,In_1595);
nand U2593 (N_2593,In_1101,In_496);
nand U2594 (N_2594,In_345,In_795);
and U2595 (N_2595,In_629,In_974);
or U2596 (N_2596,In_1729,In_483);
xor U2597 (N_2597,In_348,In_829);
nand U2598 (N_2598,In_1606,In_270);
nand U2599 (N_2599,In_335,In_1943);
or U2600 (N_2600,In_948,In_121);
and U2601 (N_2601,In_1591,In_506);
xnor U2602 (N_2602,In_1080,In_129);
nor U2603 (N_2603,In_580,In_223);
or U2604 (N_2604,In_1384,In_1571);
xnor U2605 (N_2605,In_1222,In_1471);
and U2606 (N_2606,In_203,In_1802);
xor U2607 (N_2607,In_1448,In_1192);
nor U2608 (N_2608,In_1806,In_550);
xnor U2609 (N_2609,In_224,In_500);
nand U2610 (N_2610,In_1735,In_1216);
nand U2611 (N_2611,In_380,In_518);
nand U2612 (N_2612,In_1898,In_703);
xor U2613 (N_2613,In_76,In_1141);
nor U2614 (N_2614,In_1460,In_1288);
and U2615 (N_2615,In_1370,In_117);
nor U2616 (N_2616,In_1165,In_1063);
nand U2617 (N_2617,In_472,In_206);
nand U2618 (N_2618,In_1125,In_1171);
and U2619 (N_2619,In_99,In_1765);
nor U2620 (N_2620,In_1144,In_1408);
or U2621 (N_2621,In_1879,In_25);
xnor U2622 (N_2622,In_1036,In_372);
nand U2623 (N_2623,In_1845,In_171);
or U2624 (N_2624,In_1462,In_1736);
nand U2625 (N_2625,In_360,In_291);
and U2626 (N_2626,In_1006,In_951);
and U2627 (N_2627,In_1294,In_738);
and U2628 (N_2628,In_1541,In_1116);
xor U2629 (N_2629,In_692,In_64);
xnor U2630 (N_2630,In_1090,In_567);
and U2631 (N_2631,In_1997,In_162);
and U2632 (N_2632,In_476,In_1732);
nand U2633 (N_2633,In_865,In_1809);
and U2634 (N_2634,In_216,In_494);
xor U2635 (N_2635,In_81,In_1973);
and U2636 (N_2636,In_157,In_1607);
and U2637 (N_2637,In_782,In_440);
nand U2638 (N_2638,In_797,In_1283);
nand U2639 (N_2639,In_1313,In_417);
xnor U2640 (N_2640,In_661,In_647);
nor U2641 (N_2641,In_1039,In_1763);
nor U2642 (N_2642,In_1443,In_1296);
nor U2643 (N_2643,In_1278,In_598);
and U2644 (N_2644,In_1350,In_414);
nand U2645 (N_2645,In_1108,In_1342);
xor U2646 (N_2646,In_956,In_300);
or U2647 (N_2647,In_1654,In_1517);
and U2648 (N_2648,In_250,In_229);
nor U2649 (N_2649,In_1239,In_1822);
nor U2650 (N_2650,In_1299,In_912);
nor U2651 (N_2651,In_588,In_813);
nand U2652 (N_2652,In_1655,In_318);
and U2653 (N_2653,In_1004,In_1230);
or U2654 (N_2654,In_1020,In_1611);
and U2655 (N_2655,In_1591,In_263);
xnor U2656 (N_2656,In_126,In_1860);
nand U2657 (N_2657,In_139,In_884);
nand U2658 (N_2658,In_515,In_1964);
and U2659 (N_2659,In_915,In_1622);
nor U2660 (N_2660,In_1246,In_1488);
nor U2661 (N_2661,In_1057,In_1411);
nor U2662 (N_2662,In_39,In_1304);
or U2663 (N_2663,In_339,In_391);
and U2664 (N_2664,In_1075,In_1279);
nor U2665 (N_2665,In_882,In_1657);
nand U2666 (N_2666,In_1744,In_1710);
and U2667 (N_2667,In_887,In_1296);
nand U2668 (N_2668,In_1507,In_146);
nor U2669 (N_2669,In_53,In_1438);
xnor U2670 (N_2670,In_1636,In_584);
or U2671 (N_2671,In_1152,In_1964);
and U2672 (N_2672,In_981,In_1940);
xor U2673 (N_2673,In_1572,In_616);
or U2674 (N_2674,In_1492,In_470);
nand U2675 (N_2675,In_671,In_1208);
or U2676 (N_2676,In_1863,In_440);
xor U2677 (N_2677,In_1070,In_94);
nand U2678 (N_2678,In_870,In_1864);
nand U2679 (N_2679,In_235,In_121);
xor U2680 (N_2680,In_411,In_1718);
nand U2681 (N_2681,In_954,In_1506);
and U2682 (N_2682,In_820,In_333);
or U2683 (N_2683,In_406,In_1809);
nor U2684 (N_2684,In_842,In_98);
or U2685 (N_2685,In_124,In_914);
nor U2686 (N_2686,In_1550,In_551);
or U2687 (N_2687,In_1960,In_1689);
nor U2688 (N_2688,In_1365,In_991);
or U2689 (N_2689,In_1223,In_1582);
and U2690 (N_2690,In_1538,In_49);
nor U2691 (N_2691,In_1630,In_760);
xnor U2692 (N_2692,In_1686,In_596);
xnor U2693 (N_2693,In_345,In_543);
or U2694 (N_2694,In_72,In_880);
or U2695 (N_2695,In_1561,In_60);
and U2696 (N_2696,In_1331,In_821);
nand U2697 (N_2697,In_178,In_75);
nor U2698 (N_2698,In_591,In_794);
xor U2699 (N_2699,In_881,In_622);
xnor U2700 (N_2700,In_1712,In_288);
xor U2701 (N_2701,In_162,In_1267);
or U2702 (N_2702,In_1794,In_1842);
and U2703 (N_2703,In_442,In_199);
nor U2704 (N_2704,In_1862,In_646);
nand U2705 (N_2705,In_240,In_1205);
nand U2706 (N_2706,In_1428,In_6);
nand U2707 (N_2707,In_1476,In_331);
or U2708 (N_2708,In_1003,In_1828);
nand U2709 (N_2709,In_1187,In_1887);
xor U2710 (N_2710,In_190,In_1836);
xor U2711 (N_2711,In_922,In_1456);
and U2712 (N_2712,In_302,In_558);
nand U2713 (N_2713,In_564,In_921);
or U2714 (N_2714,In_561,In_1381);
xnor U2715 (N_2715,In_1385,In_1727);
nor U2716 (N_2716,In_1170,In_1019);
nand U2717 (N_2717,In_1853,In_1008);
xor U2718 (N_2718,In_54,In_345);
xnor U2719 (N_2719,In_1916,In_1462);
xor U2720 (N_2720,In_1495,In_632);
nor U2721 (N_2721,In_187,In_1963);
and U2722 (N_2722,In_1338,In_158);
or U2723 (N_2723,In_1297,In_474);
xor U2724 (N_2724,In_342,In_551);
or U2725 (N_2725,In_1406,In_611);
or U2726 (N_2726,In_1938,In_897);
nor U2727 (N_2727,In_1483,In_470);
nor U2728 (N_2728,In_1691,In_410);
or U2729 (N_2729,In_563,In_1260);
nor U2730 (N_2730,In_386,In_1429);
and U2731 (N_2731,In_1657,In_289);
or U2732 (N_2732,In_1865,In_862);
nor U2733 (N_2733,In_437,In_1484);
and U2734 (N_2734,In_1994,In_438);
nand U2735 (N_2735,In_692,In_665);
or U2736 (N_2736,In_1166,In_339);
nand U2737 (N_2737,In_959,In_1845);
or U2738 (N_2738,In_352,In_1575);
xnor U2739 (N_2739,In_1205,In_1895);
and U2740 (N_2740,In_247,In_1026);
nor U2741 (N_2741,In_1360,In_1054);
or U2742 (N_2742,In_819,In_1515);
nand U2743 (N_2743,In_1967,In_1638);
or U2744 (N_2744,In_633,In_624);
or U2745 (N_2745,In_919,In_1554);
or U2746 (N_2746,In_1421,In_684);
xor U2747 (N_2747,In_445,In_637);
xor U2748 (N_2748,In_876,In_1632);
and U2749 (N_2749,In_1864,In_936);
or U2750 (N_2750,In_1329,In_1330);
nor U2751 (N_2751,In_1974,In_1315);
xor U2752 (N_2752,In_1416,In_1059);
and U2753 (N_2753,In_229,In_12);
nor U2754 (N_2754,In_976,In_89);
and U2755 (N_2755,In_989,In_898);
nor U2756 (N_2756,In_456,In_835);
xor U2757 (N_2757,In_638,In_1982);
nor U2758 (N_2758,In_435,In_444);
nand U2759 (N_2759,In_1961,In_1016);
or U2760 (N_2760,In_1944,In_1800);
and U2761 (N_2761,In_921,In_1377);
and U2762 (N_2762,In_1356,In_1243);
and U2763 (N_2763,In_1258,In_394);
and U2764 (N_2764,In_200,In_1923);
or U2765 (N_2765,In_1972,In_738);
or U2766 (N_2766,In_1151,In_1629);
xnor U2767 (N_2767,In_797,In_1435);
nor U2768 (N_2768,In_788,In_1788);
xor U2769 (N_2769,In_1378,In_1957);
xnor U2770 (N_2770,In_1318,In_1950);
xnor U2771 (N_2771,In_1579,In_1487);
and U2772 (N_2772,In_934,In_1390);
or U2773 (N_2773,In_1512,In_1178);
and U2774 (N_2774,In_1037,In_1163);
nor U2775 (N_2775,In_488,In_1795);
and U2776 (N_2776,In_1089,In_560);
nand U2777 (N_2777,In_240,In_1464);
nand U2778 (N_2778,In_587,In_933);
nor U2779 (N_2779,In_1265,In_267);
nor U2780 (N_2780,In_1497,In_1792);
or U2781 (N_2781,In_457,In_1242);
and U2782 (N_2782,In_819,In_329);
nor U2783 (N_2783,In_1094,In_973);
or U2784 (N_2784,In_1032,In_486);
nor U2785 (N_2785,In_1412,In_1727);
and U2786 (N_2786,In_699,In_964);
and U2787 (N_2787,In_1943,In_836);
and U2788 (N_2788,In_669,In_732);
nor U2789 (N_2789,In_201,In_1873);
nand U2790 (N_2790,In_1887,In_1535);
nand U2791 (N_2791,In_793,In_1193);
and U2792 (N_2792,In_275,In_713);
nor U2793 (N_2793,In_147,In_495);
nand U2794 (N_2794,In_1086,In_628);
nor U2795 (N_2795,In_1617,In_1682);
nor U2796 (N_2796,In_1494,In_1618);
and U2797 (N_2797,In_1160,In_378);
or U2798 (N_2798,In_272,In_1533);
xor U2799 (N_2799,In_535,In_1264);
and U2800 (N_2800,In_1109,In_1752);
nor U2801 (N_2801,In_1756,In_971);
or U2802 (N_2802,In_903,In_1473);
and U2803 (N_2803,In_265,In_948);
nand U2804 (N_2804,In_422,In_1039);
and U2805 (N_2805,In_1152,In_1752);
or U2806 (N_2806,In_740,In_718);
nor U2807 (N_2807,In_693,In_1655);
or U2808 (N_2808,In_1928,In_1666);
and U2809 (N_2809,In_444,In_1521);
nand U2810 (N_2810,In_502,In_461);
nor U2811 (N_2811,In_1753,In_1632);
xor U2812 (N_2812,In_1756,In_364);
and U2813 (N_2813,In_557,In_297);
nand U2814 (N_2814,In_458,In_1090);
nor U2815 (N_2815,In_346,In_168);
nand U2816 (N_2816,In_92,In_341);
or U2817 (N_2817,In_1899,In_66);
nor U2818 (N_2818,In_1879,In_462);
nand U2819 (N_2819,In_410,In_504);
xnor U2820 (N_2820,In_497,In_1873);
nand U2821 (N_2821,In_1322,In_1437);
nor U2822 (N_2822,In_1934,In_143);
nand U2823 (N_2823,In_1818,In_1744);
or U2824 (N_2824,In_1870,In_1756);
or U2825 (N_2825,In_1374,In_589);
nand U2826 (N_2826,In_543,In_1766);
xnor U2827 (N_2827,In_534,In_34);
and U2828 (N_2828,In_239,In_1069);
nor U2829 (N_2829,In_1748,In_1174);
and U2830 (N_2830,In_1629,In_1592);
nor U2831 (N_2831,In_1985,In_1257);
nor U2832 (N_2832,In_1041,In_690);
or U2833 (N_2833,In_1542,In_1071);
or U2834 (N_2834,In_1905,In_1411);
xnor U2835 (N_2835,In_1590,In_275);
and U2836 (N_2836,In_1589,In_1281);
nand U2837 (N_2837,In_1790,In_370);
nor U2838 (N_2838,In_447,In_502);
and U2839 (N_2839,In_788,In_1527);
or U2840 (N_2840,In_1190,In_446);
or U2841 (N_2841,In_134,In_437);
xor U2842 (N_2842,In_1176,In_1411);
nor U2843 (N_2843,In_1225,In_303);
nor U2844 (N_2844,In_1568,In_926);
and U2845 (N_2845,In_991,In_1593);
xnor U2846 (N_2846,In_1933,In_847);
nand U2847 (N_2847,In_360,In_480);
nor U2848 (N_2848,In_111,In_1097);
xor U2849 (N_2849,In_531,In_1487);
nand U2850 (N_2850,In_195,In_1997);
nand U2851 (N_2851,In_1397,In_136);
nor U2852 (N_2852,In_1193,In_750);
nand U2853 (N_2853,In_1147,In_372);
xor U2854 (N_2854,In_1083,In_402);
and U2855 (N_2855,In_1970,In_66);
nand U2856 (N_2856,In_352,In_1791);
or U2857 (N_2857,In_1346,In_1192);
nand U2858 (N_2858,In_641,In_690);
nand U2859 (N_2859,In_751,In_1723);
xor U2860 (N_2860,In_603,In_1798);
or U2861 (N_2861,In_236,In_482);
and U2862 (N_2862,In_805,In_1407);
xor U2863 (N_2863,In_177,In_1383);
nor U2864 (N_2864,In_72,In_770);
and U2865 (N_2865,In_1145,In_1787);
xor U2866 (N_2866,In_1918,In_115);
xnor U2867 (N_2867,In_786,In_831);
or U2868 (N_2868,In_613,In_1025);
or U2869 (N_2869,In_1777,In_1339);
nor U2870 (N_2870,In_441,In_1319);
or U2871 (N_2871,In_1505,In_1037);
or U2872 (N_2872,In_1430,In_786);
and U2873 (N_2873,In_1546,In_528);
or U2874 (N_2874,In_1155,In_227);
and U2875 (N_2875,In_49,In_1938);
xor U2876 (N_2876,In_1455,In_1054);
or U2877 (N_2877,In_1401,In_1066);
and U2878 (N_2878,In_878,In_990);
nor U2879 (N_2879,In_112,In_139);
or U2880 (N_2880,In_1386,In_135);
xor U2881 (N_2881,In_1054,In_1528);
or U2882 (N_2882,In_528,In_1495);
xor U2883 (N_2883,In_469,In_1366);
or U2884 (N_2884,In_1327,In_1882);
nand U2885 (N_2885,In_480,In_934);
nor U2886 (N_2886,In_1667,In_952);
and U2887 (N_2887,In_250,In_1170);
or U2888 (N_2888,In_1254,In_1916);
nor U2889 (N_2889,In_715,In_392);
or U2890 (N_2890,In_1797,In_265);
nor U2891 (N_2891,In_1648,In_983);
nand U2892 (N_2892,In_1692,In_1755);
nand U2893 (N_2893,In_161,In_632);
or U2894 (N_2894,In_1248,In_1241);
nand U2895 (N_2895,In_55,In_1314);
and U2896 (N_2896,In_319,In_764);
nand U2897 (N_2897,In_1710,In_596);
or U2898 (N_2898,In_911,In_969);
nor U2899 (N_2899,In_770,In_32);
xnor U2900 (N_2900,In_941,In_825);
and U2901 (N_2901,In_1855,In_337);
and U2902 (N_2902,In_8,In_1649);
nor U2903 (N_2903,In_1447,In_1589);
nor U2904 (N_2904,In_1341,In_816);
nand U2905 (N_2905,In_598,In_1619);
nor U2906 (N_2906,In_949,In_1953);
nand U2907 (N_2907,In_671,In_570);
nand U2908 (N_2908,In_145,In_1117);
and U2909 (N_2909,In_204,In_401);
nor U2910 (N_2910,In_1500,In_458);
nand U2911 (N_2911,In_406,In_969);
and U2912 (N_2912,In_1741,In_1347);
or U2913 (N_2913,In_203,In_1067);
xnor U2914 (N_2914,In_1246,In_1895);
or U2915 (N_2915,In_354,In_838);
nand U2916 (N_2916,In_509,In_1947);
nor U2917 (N_2917,In_527,In_480);
xnor U2918 (N_2918,In_455,In_1408);
nor U2919 (N_2919,In_762,In_367);
or U2920 (N_2920,In_1936,In_808);
nand U2921 (N_2921,In_1259,In_1058);
nor U2922 (N_2922,In_1690,In_21);
and U2923 (N_2923,In_1985,In_999);
nor U2924 (N_2924,In_1819,In_1161);
xor U2925 (N_2925,In_946,In_1454);
xor U2926 (N_2926,In_1667,In_1489);
or U2927 (N_2927,In_1166,In_156);
nand U2928 (N_2928,In_1662,In_666);
and U2929 (N_2929,In_120,In_748);
or U2930 (N_2930,In_1668,In_865);
and U2931 (N_2931,In_653,In_296);
and U2932 (N_2932,In_1719,In_1209);
nor U2933 (N_2933,In_1513,In_1060);
and U2934 (N_2934,In_984,In_607);
nor U2935 (N_2935,In_580,In_1050);
and U2936 (N_2936,In_1234,In_1419);
or U2937 (N_2937,In_1553,In_1033);
nand U2938 (N_2938,In_109,In_30);
nand U2939 (N_2939,In_15,In_1365);
nand U2940 (N_2940,In_984,In_214);
and U2941 (N_2941,In_1989,In_1095);
nor U2942 (N_2942,In_361,In_42);
and U2943 (N_2943,In_1140,In_1544);
and U2944 (N_2944,In_575,In_316);
or U2945 (N_2945,In_1010,In_856);
or U2946 (N_2946,In_877,In_1503);
nor U2947 (N_2947,In_909,In_1710);
xnor U2948 (N_2948,In_1388,In_335);
or U2949 (N_2949,In_805,In_543);
or U2950 (N_2950,In_619,In_1219);
xnor U2951 (N_2951,In_1894,In_1395);
nor U2952 (N_2952,In_1706,In_449);
xor U2953 (N_2953,In_750,In_1718);
nor U2954 (N_2954,In_1979,In_806);
xor U2955 (N_2955,In_1927,In_1590);
or U2956 (N_2956,In_1508,In_793);
and U2957 (N_2957,In_1092,In_76);
nand U2958 (N_2958,In_1622,In_1420);
xor U2959 (N_2959,In_1237,In_1933);
nand U2960 (N_2960,In_1419,In_425);
and U2961 (N_2961,In_1336,In_148);
nor U2962 (N_2962,In_1846,In_439);
and U2963 (N_2963,In_12,In_1283);
nand U2964 (N_2964,In_867,In_958);
xor U2965 (N_2965,In_1299,In_1452);
nor U2966 (N_2966,In_228,In_1911);
or U2967 (N_2967,In_1044,In_1489);
xor U2968 (N_2968,In_1826,In_1026);
and U2969 (N_2969,In_990,In_771);
xnor U2970 (N_2970,In_58,In_1284);
xor U2971 (N_2971,In_613,In_1685);
or U2972 (N_2972,In_780,In_627);
xnor U2973 (N_2973,In_584,In_1205);
nor U2974 (N_2974,In_940,In_1465);
or U2975 (N_2975,In_710,In_1862);
xor U2976 (N_2976,In_191,In_859);
or U2977 (N_2977,In_1653,In_1547);
or U2978 (N_2978,In_1881,In_415);
nand U2979 (N_2979,In_1653,In_56);
xnor U2980 (N_2980,In_576,In_1095);
nand U2981 (N_2981,In_805,In_830);
or U2982 (N_2982,In_1451,In_1621);
nor U2983 (N_2983,In_159,In_1717);
nor U2984 (N_2984,In_503,In_85);
xnor U2985 (N_2985,In_608,In_814);
nand U2986 (N_2986,In_525,In_264);
nor U2987 (N_2987,In_1849,In_441);
or U2988 (N_2988,In_636,In_831);
nor U2989 (N_2989,In_619,In_1790);
nand U2990 (N_2990,In_870,In_394);
nor U2991 (N_2991,In_36,In_1989);
xor U2992 (N_2992,In_957,In_701);
nand U2993 (N_2993,In_404,In_53);
nand U2994 (N_2994,In_312,In_1441);
nand U2995 (N_2995,In_1998,In_1001);
nand U2996 (N_2996,In_356,In_63);
nor U2997 (N_2997,In_332,In_464);
nand U2998 (N_2998,In_961,In_178);
and U2999 (N_2999,In_1676,In_620);
xnor U3000 (N_3000,In_1477,In_22);
xor U3001 (N_3001,In_833,In_92);
xnor U3002 (N_3002,In_1097,In_1795);
nor U3003 (N_3003,In_931,In_1883);
nor U3004 (N_3004,In_1084,In_1005);
or U3005 (N_3005,In_1587,In_1425);
or U3006 (N_3006,In_1327,In_1619);
xnor U3007 (N_3007,In_208,In_1425);
and U3008 (N_3008,In_1402,In_1079);
xnor U3009 (N_3009,In_1024,In_69);
nor U3010 (N_3010,In_1468,In_708);
nor U3011 (N_3011,In_154,In_1128);
nand U3012 (N_3012,In_1354,In_213);
nor U3013 (N_3013,In_1422,In_1209);
or U3014 (N_3014,In_1070,In_1999);
or U3015 (N_3015,In_160,In_473);
or U3016 (N_3016,In_139,In_845);
nand U3017 (N_3017,In_1590,In_612);
nor U3018 (N_3018,In_1978,In_1608);
xor U3019 (N_3019,In_1492,In_1453);
xor U3020 (N_3020,In_269,In_311);
nor U3021 (N_3021,In_243,In_1374);
xor U3022 (N_3022,In_1949,In_305);
nor U3023 (N_3023,In_1511,In_880);
xor U3024 (N_3024,In_1414,In_401);
and U3025 (N_3025,In_1832,In_189);
and U3026 (N_3026,In_1925,In_735);
nor U3027 (N_3027,In_1552,In_1981);
xnor U3028 (N_3028,In_1628,In_287);
or U3029 (N_3029,In_1605,In_1665);
nor U3030 (N_3030,In_1145,In_975);
or U3031 (N_3031,In_1707,In_1615);
xnor U3032 (N_3032,In_1000,In_589);
nor U3033 (N_3033,In_1482,In_1202);
nor U3034 (N_3034,In_773,In_1960);
nor U3035 (N_3035,In_1649,In_475);
or U3036 (N_3036,In_1716,In_7);
nand U3037 (N_3037,In_1963,In_1180);
nor U3038 (N_3038,In_228,In_1054);
xnor U3039 (N_3039,In_1486,In_359);
nand U3040 (N_3040,In_581,In_262);
or U3041 (N_3041,In_1575,In_145);
and U3042 (N_3042,In_1934,In_991);
nor U3043 (N_3043,In_1553,In_130);
xor U3044 (N_3044,In_1211,In_1450);
nor U3045 (N_3045,In_858,In_1989);
or U3046 (N_3046,In_210,In_1714);
and U3047 (N_3047,In_245,In_1057);
nor U3048 (N_3048,In_978,In_649);
and U3049 (N_3049,In_966,In_254);
xor U3050 (N_3050,In_1620,In_258);
nand U3051 (N_3051,In_274,In_1836);
nor U3052 (N_3052,In_1946,In_1705);
nand U3053 (N_3053,In_1946,In_1992);
nand U3054 (N_3054,In_1752,In_1789);
nand U3055 (N_3055,In_1388,In_1917);
xor U3056 (N_3056,In_1207,In_668);
nor U3057 (N_3057,In_178,In_921);
nand U3058 (N_3058,In_1078,In_132);
xnor U3059 (N_3059,In_508,In_1593);
xor U3060 (N_3060,In_1084,In_183);
and U3061 (N_3061,In_759,In_242);
xor U3062 (N_3062,In_1877,In_53);
and U3063 (N_3063,In_1685,In_951);
xnor U3064 (N_3064,In_1909,In_1362);
nand U3065 (N_3065,In_585,In_1299);
nand U3066 (N_3066,In_214,In_1119);
nor U3067 (N_3067,In_825,In_1543);
nor U3068 (N_3068,In_363,In_495);
xor U3069 (N_3069,In_1316,In_1005);
xnor U3070 (N_3070,In_960,In_999);
nor U3071 (N_3071,In_134,In_618);
and U3072 (N_3072,In_1399,In_22);
or U3073 (N_3073,In_929,In_1746);
nor U3074 (N_3074,In_52,In_793);
or U3075 (N_3075,In_1957,In_1175);
nand U3076 (N_3076,In_1963,In_282);
and U3077 (N_3077,In_1673,In_38);
and U3078 (N_3078,In_343,In_512);
nor U3079 (N_3079,In_154,In_1545);
and U3080 (N_3080,In_970,In_1057);
and U3081 (N_3081,In_716,In_585);
nand U3082 (N_3082,In_894,In_852);
or U3083 (N_3083,In_1624,In_892);
nor U3084 (N_3084,In_1212,In_1258);
nor U3085 (N_3085,In_1157,In_391);
nand U3086 (N_3086,In_1760,In_1629);
xor U3087 (N_3087,In_1892,In_580);
and U3088 (N_3088,In_386,In_1665);
and U3089 (N_3089,In_204,In_724);
and U3090 (N_3090,In_152,In_1171);
nand U3091 (N_3091,In_80,In_1463);
and U3092 (N_3092,In_1486,In_1859);
xor U3093 (N_3093,In_275,In_1176);
and U3094 (N_3094,In_1418,In_1510);
nand U3095 (N_3095,In_727,In_1144);
nand U3096 (N_3096,In_1207,In_1677);
or U3097 (N_3097,In_1926,In_785);
or U3098 (N_3098,In_1867,In_115);
xor U3099 (N_3099,In_324,In_18);
and U3100 (N_3100,In_1938,In_632);
nand U3101 (N_3101,In_513,In_510);
and U3102 (N_3102,In_675,In_795);
and U3103 (N_3103,In_1558,In_590);
or U3104 (N_3104,In_454,In_486);
and U3105 (N_3105,In_828,In_1216);
nand U3106 (N_3106,In_1592,In_760);
nand U3107 (N_3107,In_466,In_503);
and U3108 (N_3108,In_1198,In_1000);
nor U3109 (N_3109,In_1166,In_1396);
or U3110 (N_3110,In_710,In_1543);
nor U3111 (N_3111,In_1945,In_1292);
or U3112 (N_3112,In_1293,In_1081);
or U3113 (N_3113,In_1011,In_1977);
nor U3114 (N_3114,In_194,In_1485);
and U3115 (N_3115,In_766,In_1042);
nand U3116 (N_3116,In_1926,In_1476);
or U3117 (N_3117,In_1176,In_1415);
xnor U3118 (N_3118,In_1186,In_537);
xnor U3119 (N_3119,In_89,In_228);
nor U3120 (N_3120,In_1068,In_233);
xnor U3121 (N_3121,In_574,In_1459);
and U3122 (N_3122,In_1779,In_995);
or U3123 (N_3123,In_1007,In_1924);
nand U3124 (N_3124,In_1091,In_538);
and U3125 (N_3125,In_336,In_1657);
nor U3126 (N_3126,In_463,In_388);
nor U3127 (N_3127,In_629,In_580);
xnor U3128 (N_3128,In_1052,In_1645);
nand U3129 (N_3129,In_61,In_1845);
nor U3130 (N_3130,In_1673,In_128);
xnor U3131 (N_3131,In_635,In_1969);
nand U3132 (N_3132,In_274,In_578);
and U3133 (N_3133,In_1529,In_1997);
xnor U3134 (N_3134,In_995,In_389);
nand U3135 (N_3135,In_695,In_179);
xnor U3136 (N_3136,In_1538,In_1485);
xor U3137 (N_3137,In_554,In_1784);
or U3138 (N_3138,In_1041,In_1461);
or U3139 (N_3139,In_1764,In_1542);
or U3140 (N_3140,In_1239,In_1334);
nor U3141 (N_3141,In_334,In_940);
nor U3142 (N_3142,In_201,In_1689);
and U3143 (N_3143,In_1236,In_1990);
xor U3144 (N_3144,In_1452,In_240);
nand U3145 (N_3145,In_237,In_1041);
xnor U3146 (N_3146,In_1697,In_1861);
and U3147 (N_3147,In_1532,In_1527);
and U3148 (N_3148,In_1840,In_1364);
nor U3149 (N_3149,In_1664,In_530);
nand U3150 (N_3150,In_1326,In_399);
and U3151 (N_3151,In_1018,In_746);
or U3152 (N_3152,In_1024,In_1330);
nand U3153 (N_3153,In_1016,In_106);
nand U3154 (N_3154,In_1374,In_1224);
xnor U3155 (N_3155,In_797,In_1580);
nor U3156 (N_3156,In_1133,In_342);
or U3157 (N_3157,In_1608,In_269);
and U3158 (N_3158,In_301,In_794);
nand U3159 (N_3159,In_1477,In_857);
xnor U3160 (N_3160,In_1375,In_843);
xnor U3161 (N_3161,In_60,In_12);
and U3162 (N_3162,In_339,In_1800);
nor U3163 (N_3163,In_874,In_1944);
nor U3164 (N_3164,In_1572,In_658);
nor U3165 (N_3165,In_1423,In_796);
and U3166 (N_3166,In_847,In_1284);
or U3167 (N_3167,In_1764,In_1266);
nand U3168 (N_3168,In_179,In_1894);
and U3169 (N_3169,In_346,In_1216);
nor U3170 (N_3170,In_1240,In_1210);
nor U3171 (N_3171,In_1962,In_1662);
nor U3172 (N_3172,In_1304,In_206);
and U3173 (N_3173,In_1336,In_516);
or U3174 (N_3174,In_494,In_1588);
nor U3175 (N_3175,In_837,In_1164);
nor U3176 (N_3176,In_1029,In_1557);
and U3177 (N_3177,In_1970,In_1504);
nand U3178 (N_3178,In_1643,In_570);
and U3179 (N_3179,In_342,In_206);
nor U3180 (N_3180,In_1917,In_506);
xnor U3181 (N_3181,In_20,In_945);
nand U3182 (N_3182,In_1720,In_1869);
nand U3183 (N_3183,In_1969,In_1630);
or U3184 (N_3184,In_1736,In_655);
and U3185 (N_3185,In_1683,In_245);
nand U3186 (N_3186,In_1074,In_1768);
nor U3187 (N_3187,In_1130,In_1908);
nor U3188 (N_3188,In_1986,In_919);
and U3189 (N_3189,In_1409,In_9);
and U3190 (N_3190,In_523,In_1766);
or U3191 (N_3191,In_639,In_1776);
nor U3192 (N_3192,In_1645,In_1750);
nand U3193 (N_3193,In_26,In_668);
xor U3194 (N_3194,In_86,In_605);
and U3195 (N_3195,In_1774,In_1512);
and U3196 (N_3196,In_132,In_958);
and U3197 (N_3197,In_541,In_31);
nor U3198 (N_3198,In_1977,In_1173);
or U3199 (N_3199,In_1535,In_420);
xor U3200 (N_3200,In_1636,In_1656);
nand U3201 (N_3201,In_1317,In_1947);
xor U3202 (N_3202,In_75,In_1740);
nor U3203 (N_3203,In_737,In_268);
and U3204 (N_3204,In_1749,In_736);
and U3205 (N_3205,In_914,In_181);
or U3206 (N_3206,In_1853,In_432);
nor U3207 (N_3207,In_1285,In_927);
nor U3208 (N_3208,In_605,In_500);
or U3209 (N_3209,In_343,In_612);
nand U3210 (N_3210,In_1349,In_1639);
nand U3211 (N_3211,In_1834,In_1542);
and U3212 (N_3212,In_1676,In_125);
nand U3213 (N_3213,In_1201,In_1925);
or U3214 (N_3214,In_127,In_1008);
nand U3215 (N_3215,In_779,In_1321);
xnor U3216 (N_3216,In_253,In_803);
and U3217 (N_3217,In_1132,In_1262);
and U3218 (N_3218,In_1779,In_411);
nor U3219 (N_3219,In_963,In_1489);
xnor U3220 (N_3220,In_1656,In_1450);
or U3221 (N_3221,In_1192,In_460);
nor U3222 (N_3222,In_1488,In_272);
xor U3223 (N_3223,In_1015,In_1684);
xor U3224 (N_3224,In_1667,In_1689);
nor U3225 (N_3225,In_1964,In_995);
or U3226 (N_3226,In_1816,In_142);
nand U3227 (N_3227,In_1318,In_57);
nor U3228 (N_3228,In_1798,In_856);
nand U3229 (N_3229,In_590,In_1649);
xnor U3230 (N_3230,In_1578,In_1900);
nand U3231 (N_3231,In_1746,In_124);
nand U3232 (N_3232,In_769,In_1139);
nand U3233 (N_3233,In_1876,In_865);
or U3234 (N_3234,In_1083,In_754);
xnor U3235 (N_3235,In_1808,In_424);
nand U3236 (N_3236,In_1936,In_672);
xor U3237 (N_3237,In_366,In_1448);
nor U3238 (N_3238,In_1919,In_1270);
or U3239 (N_3239,In_1069,In_1552);
xor U3240 (N_3240,In_1747,In_693);
and U3241 (N_3241,In_423,In_502);
and U3242 (N_3242,In_1505,In_318);
xnor U3243 (N_3243,In_1095,In_903);
or U3244 (N_3244,In_1279,In_353);
nor U3245 (N_3245,In_561,In_440);
nor U3246 (N_3246,In_379,In_226);
xor U3247 (N_3247,In_1973,In_1244);
or U3248 (N_3248,In_1989,In_1498);
nand U3249 (N_3249,In_902,In_976);
nand U3250 (N_3250,In_1088,In_1862);
nor U3251 (N_3251,In_28,In_239);
and U3252 (N_3252,In_673,In_766);
and U3253 (N_3253,In_271,In_198);
or U3254 (N_3254,In_1836,In_1087);
xnor U3255 (N_3255,In_1749,In_850);
or U3256 (N_3256,In_761,In_1467);
xor U3257 (N_3257,In_39,In_1661);
xnor U3258 (N_3258,In_444,In_1460);
nor U3259 (N_3259,In_1244,In_888);
nor U3260 (N_3260,In_144,In_1447);
and U3261 (N_3261,In_340,In_1549);
nor U3262 (N_3262,In_962,In_1184);
nor U3263 (N_3263,In_1732,In_1248);
and U3264 (N_3264,In_1138,In_1945);
nor U3265 (N_3265,In_917,In_1179);
xnor U3266 (N_3266,In_1288,In_566);
nor U3267 (N_3267,In_1006,In_1171);
nor U3268 (N_3268,In_195,In_1206);
nand U3269 (N_3269,In_1358,In_787);
nor U3270 (N_3270,In_1521,In_45);
and U3271 (N_3271,In_1757,In_1412);
or U3272 (N_3272,In_182,In_1428);
nand U3273 (N_3273,In_734,In_44);
xor U3274 (N_3274,In_303,In_1545);
nand U3275 (N_3275,In_1212,In_1701);
and U3276 (N_3276,In_1075,In_1867);
xor U3277 (N_3277,In_467,In_857);
nor U3278 (N_3278,In_865,In_548);
or U3279 (N_3279,In_639,In_1287);
or U3280 (N_3280,In_975,In_90);
xnor U3281 (N_3281,In_375,In_1539);
nand U3282 (N_3282,In_1116,In_1681);
or U3283 (N_3283,In_1025,In_1135);
and U3284 (N_3284,In_500,In_186);
xnor U3285 (N_3285,In_453,In_587);
xnor U3286 (N_3286,In_185,In_1682);
nor U3287 (N_3287,In_1507,In_1375);
nor U3288 (N_3288,In_749,In_925);
nor U3289 (N_3289,In_347,In_1826);
and U3290 (N_3290,In_737,In_1358);
and U3291 (N_3291,In_730,In_356);
or U3292 (N_3292,In_1987,In_1775);
and U3293 (N_3293,In_505,In_1115);
nand U3294 (N_3294,In_1259,In_771);
nand U3295 (N_3295,In_723,In_283);
nor U3296 (N_3296,In_1598,In_1375);
nor U3297 (N_3297,In_85,In_1733);
xnor U3298 (N_3298,In_995,In_1447);
nor U3299 (N_3299,In_1138,In_1204);
nand U3300 (N_3300,In_94,In_205);
or U3301 (N_3301,In_1149,In_808);
or U3302 (N_3302,In_1354,In_1141);
xnor U3303 (N_3303,In_303,In_657);
and U3304 (N_3304,In_1579,In_994);
xnor U3305 (N_3305,In_1234,In_1012);
nand U3306 (N_3306,In_36,In_1916);
nor U3307 (N_3307,In_523,In_1283);
nand U3308 (N_3308,In_1825,In_329);
nor U3309 (N_3309,In_1021,In_1747);
nor U3310 (N_3310,In_555,In_822);
or U3311 (N_3311,In_1437,In_1498);
nand U3312 (N_3312,In_1121,In_1523);
xor U3313 (N_3313,In_94,In_1461);
and U3314 (N_3314,In_904,In_884);
nor U3315 (N_3315,In_712,In_1786);
nand U3316 (N_3316,In_823,In_32);
xnor U3317 (N_3317,In_543,In_695);
or U3318 (N_3318,In_1195,In_1362);
nor U3319 (N_3319,In_1783,In_1048);
nor U3320 (N_3320,In_959,In_266);
or U3321 (N_3321,In_1507,In_1095);
and U3322 (N_3322,In_1383,In_1736);
and U3323 (N_3323,In_1344,In_1319);
or U3324 (N_3324,In_441,In_176);
nor U3325 (N_3325,In_796,In_19);
xnor U3326 (N_3326,In_550,In_196);
nand U3327 (N_3327,In_904,In_1666);
nor U3328 (N_3328,In_1979,In_665);
or U3329 (N_3329,In_859,In_1729);
xor U3330 (N_3330,In_1794,In_1019);
and U3331 (N_3331,In_1755,In_159);
xor U3332 (N_3332,In_1377,In_1783);
and U3333 (N_3333,In_392,In_1513);
and U3334 (N_3334,In_1357,In_739);
xor U3335 (N_3335,In_528,In_175);
or U3336 (N_3336,In_283,In_1084);
and U3337 (N_3337,In_1528,In_1395);
nor U3338 (N_3338,In_897,In_224);
xor U3339 (N_3339,In_740,In_108);
nand U3340 (N_3340,In_1707,In_1172);
and U3341 (N_3341,In_589,In_1617);
nor U3342 (N_3342,In_216,In_680);
nand U3343 (N_3343,In_1204,In_1585);
nand U3344 (N_3344,In_1661,In_1936);
xor U3345 (N_3345,In_1357,In_1926);
or U3346 (N_3346,In_81,In_1252);
nand U3347 (N_3347,In_930,In_732);
nor U3348 (N_3348,In_1487,In_1080);
xor U3349 (N_3349,In_1438,In_1890);
xor U3350 (N_3350,In_504,In_622);
nor U3351 (N_3351,In_766,In_203);
xnor U3352 (N_3352,In_1378,In_1712);
xnor U3353 (N_3353,In_480,In_10);
or U3354 (N_3354,In_1267,In_991);
xnor U3355 (N_3355,In_133,In_373);
or U3356 (N_3356,In_1767,In_1776);
nor U3357 (N_3357,In_1938,In_1897);
and U3358 (N_3358,In_43,In_1710);
and U3359 (N_3359,In_91,In_730);
xnor U3360 (N_3360,In_1926,In_309);
nand U3361 (N_3361,In_1205,In_998);
nor U3362 (N_3362,In_1926,In_1743);
nor U3363 (N_3363,In_4,In_136);
and U3364 (N_3364,In_1943,In_1106);
xnor U3365 (N_3365,In_1212,In_137);
nor U3366 (N_3366,In_1376,In_827);
nand U3367 (N_3367,In_108,In_595);
xnor U3368 (N_3368,In_31,In_1411);
and U3369 (N_3369,In_312,In_128);
nor U3370 (N_3370,In_1776,In_1913);
xor U3371 (N_3371,In_787,In_1411);
or U3372 (N_3372,In_322,In_1028);
and U3373 (N_3373,In_1538,In_1833);
and U3374 (N_3374,In_169,In_1218);
and U3375 (N_3375,In_349,In_1304);
nor U3376 (N_3376,In_1410,In_1028);
nand U3377 (N_3377,In_901,In_1910);
and U3378 (N_3378,In_964,In_1667);
xor U3379 (N_3379,In_1662,In_471);
nand U3380 (N_3380,In_125,In_592);
xor U3381 (N_3381,In_369,In_882);
xnor U3382 (N_3382,In_832,In_514);
and U3383 (N_3383,In_1642,In_270);
and U3384 (N_3384,In_625,In_407);
nor U3385 (N_3385,In_708,In_1600);
nand U3386 (N_3386,In_1862,In_1975);
and U3387 (N_3387,In_1882,In_1576);
or U3388 (N_3388,In_417,In_768);
nand U3389 (N_3389,In_392,In_1944);
nand U3390 (N_3390,In_645,In_241);
or U3391 (N_3391,In_1137,In_641);
xnor U3392 (N_3392,In_1311,In_1898);
xnor U3393 (N_3393,In_1899,In_1654);
or U3394 (N_3394,In_258,In_1959);
and U3395 (N_3395,In_1859,In_1610);
xnor U3396 (N_3396,In_552,In_228);
nor U3397 (N_3397,In_1496,In_245);
and U3398 (N_3398,In_769,In_1537);
nand U3399 (N_3399,In_643,In_1959);
nand U3400 (N_3400,In_1803,In_997);
and U3401 (N_3401,In_1501,In_244);
and U3402 (N_3402,In_29,In_876);
nor U3403 (N_3403,In_323,In_1333);
nor U3404 (N_3404,In_743,In_692);
and U3405 (N_3405,In_1328,In_671);
or U3406 (N_3406,In_740,In_1229);
and U3407 (N_3407,In_1720,In_1599);
nor U3408 (N_3408,In_962,In_1523);
or U3409 (N_3409,In_675,In_180);
nor U3410 (N_3410,In_1794,In_663);
nand U3411 (N_3411,In_412,In_97);
xnor U3412 (N_3412,In_1311,In_180);
xnor U3413 (N_3413,In_1499,In_1886);
or U3414 (N_3414,In_1290,In_47);
and U3415 (N_3415,In_1750,In_1824);
nand U3416 (N_3416,In_1287,In_300);
xnor U3417 (N_3417,In_91,In_1595);
xor U3418 (N_3418,In_789,In_198);
nand U3419 (N_3419,In_1751,In_1460);
nand U3420 (N_3420,In_959,In_1473);
and U3421 (N_3421,In_1184,In_1723);
xor U3422 (N_3422,In_575,In_396);
or U3423 (N_3423,In_686,In_1954);
or U3424 (N_3424,In_1888,In_90);
or U3425 (N_3425,In_1434,In_277);
and U3426 (N_3426,In_923,In_1636);
xnor U3427 (N_3427,In_1208,In_1369);
nand U3428 (N_3428,In_1325,In_1477);
and U3429 (N_3429,In_1704,In_433);
or U3430 (N_3430,In_1299,In_675);
or U3431 (N_3431,In_1088,In_616);
xor U3432 (N_3432,In_866,In_1459);
xnor U3433 (N_3433,In_726,In_828);
nand U3434 (N_3434,In_1187,In_1157);
nand U3435 (N_3435,In_537,In_1586);
nand U3436 (N_3436,In_1556,In_935);
nand U3437 (N_3437,In_1097,In_179);
nor U3438 (N_3438,In_898,In_165);
or U3439 (N_3439,In_831,In_204);
or U3440 (N_3440,In_72,In_1896);
xor U3441 (N_3441,In_1719,In_303);
xor U3442 (N_3442,In_326,In_1067);
nand U3443 (N_3443,In_872,In_1279);
nand U3444 (N_3444,In_1856,In_371);
nand U3445 (N_3445,In_1541,In_32);
xor U3446 (N_3446,In_1606,In_1667);
and U3447 (N_3447,In_386,In_1168);
xnor U3448 (N_3448,In_1680,In_143);
nand U3449 (N_3449,In_252,In_31);
xnor U3450 (N_3450,In_1929,In_1923);
nand U3451 (N_3451,In_1581,In_1828);
xor U3452 (N_3452,In_906,In_1523);
xor U3453 (N_3453,In_1683,In_1620);
or U3454 (N_3454,In_1076,In_1487);
nor U3455 (N_3455,In_54,In_1223);
nand U3456 (N_3456,In_1677,In_1546);
and U3457 (N_3457,In_406,In_1678);
nand U3458 (N_3458,In_1145,In_1961);
xor U3459 (N_3459,In_1683,In_1667);
and U3460 (N_3460,In_1842,In_241);
and U3461 (N_3461,In_1211,In_1923);
nand U3462 (N_3462,In_787,In_638);
xnor U3463 (N_3463,In_123,In_914);
xor U3464 (N_3464,In_879,In_1258);
nand U3465 (N_3465,In_1302,In_51);
or U3466 (N_3466,In_1919,In_1532);
and U3467 (N_3467,In_403,In_1596);
xnor U3468 (N_3468,In_188,In_647);
or U3469 (N_3469,In_861,In_34);
nor U3470 (N_3470,In_1638,In_347);
or U3471 (N_3471,In_1032,In_1891);
or U3472 (N_3472,In_1312,In_1549);
and U3473 (N_3473,In_44,In_434);
nand U3474 (N_3474,In_1672,In_1486);
nor U3475 (N_3475,In_479,In_1275);
nor U3476 (N_3476,In_1267,In_1065);
and U3477 (N_3477,In_630,In_42);
xnor U3478 (N_3478,In_268,In_812);
xor U3479 (N_3479,In_747,In_1073);
nor U3480 (N_3480,In_1987,In_1703);
xor U3481 (N_3481,In_1587,In_1215);
nor U3482 (N_3482,In_1133,In_1609);
nor U3483 (N_3483,In_115,In_329);
and U3484 (N_3484,In_1180,In_1808);
or U3485 (N_3485,In_1925,In_1553);
or U3486 (N_3486,In_419,In_521);
nor U3487 (N_3487,In_1740,In_1060);
or U3488 (N_3488,In_588,In_1461);
and U3489 (N_3489,In_102,In_1631);
and U3490 (N_3490,In_1715,In_1663);
or U3491 (N_3491,In_97,In_1575);
xnor U3492 (N_3492,In_1444,In_858);
and U3493 (N_3493,In_941,In_651);
nor U3494 (N_3494,In_1670,In_1519);
nand U3495 (N_3495,In_609,In_716);
and U3496 (N_3496,In_1846,In_387);
or U3497 (N_3497,In_100,In_1036);
nor U3498 (N_3498,In_749,In_921);
nand U3499 (N_3499,In_1496,In_442);
and U3500 (N_3500,In_557,In_1921);
xor U3501 (N_3501,In_937,In_1013);
xor U3502 (N_3502,In_519,In_571);
nand U3503 (N_3503,In_1721,In_1447);
nor U3504 (N_3504,In_350,In_1037);
and U3505 (N_3505,In_1707,In_694);
nand U3506 (N_3506,In_1699,In_157);
or U3507 (N_3507,In_1141,In_1163);
nand U3508 (N_3508,In_1869,In_463);
xnor U3509 (N_3509,In_529,In_683);
nor U3510 (N_3510,In_1542,In_801);
and U3511 (N_3511,In_1079,In_1619);
xnor U3512 (N_3512,In_809,In_1197);
xnor U3513 (N_3513,In_494,In_383);
xor U3514 (N_3514,In_1495,In_1195);
nand U3515 (N_3515,In_1399,In_1199);
nand U3516 (N_3516,In_854,In_402);
nor U3517 (N_3517,In_1960,In_759);
nand U3518 (N_3518,In_519,In_373);
nor U3519 (N_3519,In_1414,In_1448);
and U3520 (N_3520,In_901,In_1318);
xnor U3521 (N_3521,In_1,In_495);
nor U3522 (N_3522,In_291,In_1501);
and U3523 (N_3523,In_1331,In_567);
nand U3524 (N_3524,In_1171,In_1554);
xnor U3525 (N_3525,In_141,In_1347);
and U3526 (N_3526,In_769,In_651);
or U3527 (N_3527,In_274,In_1594);
nand U3528 (N_3528,In_2,In_1240);
or U3529 (N_3529,In_910,In_1473);
and U3530 (N_3530,In_1605,In_445);
nand U3531 (N_3531,In_275,In_579);
or U3532 (N_3532,In_30,In_1757);
and U3533 (N_3533,In_679,In_244);
or U3534 (N_3534,In_704,In_1507);
nor U3535 (N_3535,In_775,In_154);
nor U3536 (N_3536,In_1779,In_1493);
nand U3537 (N_3537,In_91,In_255);
and U3538 (N_3538,In_1635,In_1859);
or U3539 (N_3539,In_1234,In_1409);
nand U3540 (N_3540,In_1491,In_1465);
nand U3541 (N_3541,In_1134,In_99);
nor U3542 (N_3542,In_1643,In_1284);
xor U3543 (N_3543,In_1474,In_1770);
nor U3544 (N_3544,In_1721,In_125);
nand U3545 (N_3545,In_1739,In_1408);
and U3546 (N_3546,In_63,In_474);
or U3547 (N_3547,In_1337,In_16);
or U3548 (N_3548,In_1748,In_1263);
nor U3549 (N_3549,In_278,In_1176);
nor U3550 (N_3550,In_730,In_501);
and U3551 (N_3551,In_1979,In_617);
nor U3552 (N_3552,In_225,In_355);
xor U3553 (N_3553,In_1905,In_160);
xnor U3554 (N_3554,In_1397,In_1528);
or U3555 (N_3555,In_1529,In_438);
and U3556 (N_3556,In_633,In_1807);
xnor U3557 (N_3557,In_238,In_1037);
nor U3558 (N_3558,In_923,In_423);
or U3559 (N_3559,In_1634,In_788);
nand U3560 (N_3560,In_63,In_537);
xnor U3561 (N_3561,In_1514,In_990);
xnor U3562 (N_3562,In_1818,In_246);
xnor U3563 (N_3563,In_218,In_1225);
nand U3564 (N_3564,In_1275,In_1473);
or U3565 (N_3565,In_1791,In_1871);
or U3566 (N_3566,In_1994,In_1122);
and U3567 (N_3567,In_153,In_174);
or U3568 (N_3568,In_209,In_1733);
nor U3569 (N_3569,In_894,In_1536);
and U3570 (N_3570,In_1622,In_851);
nor U3571 (N_3571,In_420,In_561);
nor U3572 (N_3572,In_782,In_747);
or U3573 (N_3573,In_431,In_1361);
or U3574 (N_3574,In_326,In_1069);
nand U3575 (N_3575,In_788,In_0);
or U3576 (N_3576,In_238,In_598);
xnor U3577 (N_3577,In_1242,In_1773);
xor U3578 (N_3578,In_637,In_1906);
nand U3579 (N_3579,In_791,In_1215);
or U3580 (N_3580,In_1490,In_343);
or U3581 (N_3581,In_1047,In_1701);
and U3582 (N_3582,In_1027,In_796);
xnor U3583 (N_3583,In_584,In_1446);
or U3584 (N_3584,In_1389,In_1180);
or U3585 (N_3585,In_311,In_1268);
nor U3586 (N_3586,In_1828,In_597);
xnor U3587 (N_3587,In_1789,In_1910);
nor U3588 (N_3588,In_1253,In_1105);
nand U3589 (N_3589,In_467,In_1620);
nor U3590 (N_3590,In_1041,In_6);
xor U3591 (N_3591,In_1809,In_441);
xor U3592 (N_3592,In_1668,In_533);
nor U3593 (N_3593,In_42,In_880);
and U3594 (N_3594,In_1274,In_293);
and U3595 (N_3595,In_1864,In_897);
nor U3596 (N_3596,In_1825,In_1447);
and U3597 (N_3597,In_1803,In_1926);
nand U3598 (N_3598,In_1203,In_298);
and U3599 (N_3599,In_665,In_1834);
or U3600 (N_3600,In_1107,In_572);
or U3601 (N_3601,In_863,In_1173);
and U3602 (N_3602,In_1575,In_23);
xnor U3603 (N_3603,In_986,In_1082);
nor U3604 (N_3604,In_461,In_1368);
xor U3605 (N_3605,In_192,In_1461);
xor U3606 (N_3606,In_96,In_1073);
nand U3607 (N_3607,In_1023,In_308);
or U3608 (N_3608,In_478,In_343);
nor U3609 (N_3609,In_622,In_593);
and U3610 (N_3610,In_972,In_1921);
nand U3611 (N_3611,In_660,In_701);
nand U3612 (N_3612,In_1832,In_236);
xor U3613 (N_3613,In_769,In_456);
nand U3614 (N_3614,In_1816,In_21);
or U3615 (N_3615,In_1197,In_495);
nor U3616 (N_3616,In_813,In_379);
and U3617 (N_3617,In_1812,In_1263);
and U3618 (N_3618,In_380,In_1407);
nor U3619 (N_3619,In_884,In_422);
nand U3620 (N_3620,In_379,In_375);
or U3621 (N_3621,In_789,In_1924);
nor U3622 (N_3622,In_400,In_258);
nor U3623 (N_3623,In_543,In_1425);
or U3624 (N_3624,In_22,In_1498);
nor U3625 (N_3625,In_1392,In_1474);
nor U3626 (N_3626,In_754,In_1450);
and U3627 (N_3627,In_749,In_134);
and U3628 (N_3628,In_1208,In_1980);
nor U3629 (N_3629,In_443,In_730);
nor U3630 (N_3630,In_730,In_336);
or U3631 (N_3631,In_753,In_43);
xor U3632 (N_3632,In_168,In_624);
or U3633 (N_3633,In_543,In_1220);
nand U3634 (N_3634,In_888,In_1798);
and U3635 (N_3635,In_301,In_362);
and U3636 (N_3636,In_1111,In_1685);
nand U3637 (N_3637,In_709,In_94);
nor U3638 (N_3638,In_93,In_1229);
or U3639 (N_3639,In_781,In_1278);
and U3640 (N_3640,In_551,In_682);
nor U3641 (N_3641,In_197,In_842);
or U3642 (N_3642,In_1813,In_596);
nor U3643 (N_3643,In_324,In_1117);
nor U3644 (N_3644,In_1603,In_407);
and U3645 (N_3645,In_348,In_1753);
or U3646 (N_3646,In_913,In_140);
xnor U3647 (N_3647,In_1322,In_1332);
and U3648 (N_3648,In_29,In_1314);
or U3649 (N_3649,In_1827,In_157);
nor U3650 (N_3650,In_1228,In_1016);
nor U3651 (N_3651,In_950,In_676);
or U3652 (N_3652,In_150,In_1268);
nor U3653 (N_3653,In_991,In_1316);
or U3654 (N_3654,In_1576,In_1620);
and U3655 (N_3655,In_1857,In_351);
xnor U3656 (N_3656,In_974,In_1090);
nor U3657 (N_3657,In_960,In_498);
nor U3658 (N_3658,In_924,In_385);
nand U3659 (N_3659,In_1297,In_1764);
and U3660 (N_3660,In_566,In_1929);
nand U3661 (N_3661,In_1092,In_1790);
or U3662 (N_3662,In_1156,In_1628);
xor U3663 (N_3663,In_698,In_1958);
nand U3664 (N_3664,In_340,In_1397);
nor U3665 (N_3665,In_203,In_417);
xnor U3666 (N_3666,In_1129,In_1303);
and U3667 (N_3667,In_1054,In_1518);
xor U3668 (N_3668,In_342,In_810);
nand U3669 (N_3669,In_1932,In_581);
and U3670 (N_3670,In_1734,In_1682);
nand U3671 (N_3671,In_1073,In_1645);
or U3672 (N_3672,In_1854,In_544);
or U3673 (N_3673,In_1842,In_157);
xor U3674 (N_3674,In_1926,In_444);
nor U3675 (N_3675,In_1506,In_414);
xnor U3676 (N_3676,In_1529,In_1795);
or U3677 (N_3677,In_673,In_1528);
or U3678 (N_3678,In_1397,In_361);
or U3679 (N_3679,In_255,In_1548);
nand U3680 (N_3680,In_579,In_1409);
and U3681 (N_3681,In_718,In_914);
nand U3682 (N_3682,In_1983,In_1008);
and U3683 (N_3683,In_1727,In_713);
nand U3684 (N_3684,In_709,In_732);
and U3685 (N_3685,In_86,In_434);
nand U3686 (N_3686,In_746,In_1172);
or U3687 (N_3687,In_1138,In_1287);
or U3688 (N_3688,In_86,In_1415);
nand U3689 (N_3689,In_146,In_1646);
nor U3690 (N_3690,In_1585,In_1870);
or U3691 (N_3691,In_1889,In_1935);
nor U3692 (N_3692,In_1734,In_7);
nor U3693 (N_3693,In_1079,In_1325);
or U3694 (N_3694,In_544,In_1043);
nor U3695 (N_3695,In_805,In_1877);
and U3696 (N_3696,In_1014,In_234);
or U3697 (N_3697,In_1950,In_1792);
nand U3698 (N_3698,In_1393,In_261);
or U3699 (N_3699,In_1656,In_112);
and U3700 (N_3700,In_1920,In_1249);
nand U3701 (N_3701,In_140,In_1273);
nand U3702 (N_3702,In_908,In_1543);
xnor U3703 (N_3703,In_501,In_340);
nor U3704 (N_3704,In_1192,In_1271);
and U3705 (N_3705,In_68,In_31);
nor U3706 (N_3706,In_1092,In_1675);
xnor U3707 (N_3707,In_830,In_630);
or U3708 (N_3708,In_3,In_1984);
xnor U3709 (N_3709,In_316,In_1962);
nand U3710 (N_3710,In_537,In_117);
or U3711 (N_3711,In_1942,In_1711);
and U3712 (N_3712,In_744,In_1981);
or U3713 (N_3713,In_1026,In_1219);
and U3714 (N_3714,In_537,In_1773);
or U3715 (N_3715,In_367,In_1283);
or U3716 (N_3716,In_1272,In_569);
nor U3717 (N_3717,In_1827,In_1868);
nor U3718 (N_3718,In_729,In_697);
nor U3719 (N_3719,In_145,In_1430);
nor U3720 (N_3720,In_113,In_1342);
and U3721 (N_3721,In_661,In_573);
xor U3722 (N_3722,In_1201,In_1070);
nand U3723 (N_3723,In_1379,In_1309);
and U3724 (N_3724,In_1686,In_732);
nor U3725 (N_3725,In_119,In_455);
nand U3726 (N_3726,In_1692,In_276);
xor U3727 (N_3727,In_978,In_1170);
and U3728 (N_3728,In_1707,In_1971);
and U3729 (N_3729,In_603,In_188);
nand U3730 (N_3730,In_961,In_364);
and U3731 (N_3731,In_1317,In_541);
and U3732 (N_3732,In_66,In_732);
and U3733 (N_3733,In_106,In_1582);
xor U3734 (N_3734,In_1402,In_1336);
nor U3735 (N_3735,In_146,In_1324);
xor U3736 (N_3736,In_629,In_955);
or U3737 (N_3737,In_992,In_1722);
xnor U3738 (N_3738,In_303,In_163);
nor U3739 (N_3739,In_103,In_1686);
xnor U3740 (N_3740,In_230,In_147);
nor U3741 (N_3741,In_1028,In_572);
xnor U3742 (N_3742,In_238,In_1472);
xor U3743 (N_3743,In_1506,In_581);
xor U3744 (N_3744,In_309,In_1189);
nor U3745 (N_3745,In_1334,In_720);
and U3746 (N_3746,In_304,In_157);
nor U3747 (N_3747,In_399,In_871);
xnor U3748 (N_3748,In_107,In_922);
or U3749 (N_3749,In_386,In_96);
or U3750 (N_3750,In_784,In_1819);
nor U3751 (N_3751,In_1209,In_1372);
and U3752 (N_3752,In_1378,In_452);
nand U3753 (N_3753,In_1144,In_176);
nand U3754 (N_3754,In_1911,In_934);
nand U3755 (N_3755,In_155,In_1779);
nand U3756 (N_3756,In_223,In_123);
nand U3757 (N_3757,In_1856,In_1005);
or U3758 (N_3758,In_1726,In_1335);
and U3759 (N_3759,In_972,In_1771);
nand U3760 (N_3760,In_551,In_143);
xnor U3761 (N_3761,In_1324,In_800);
nand U3762 (N_3762,In_973,In_1390);
and U3763 (N_3763,In_451,In_1673);
nor U3764 (N_3764,In_1130,In_396);
or U3765 (N_3765,In_1728,In_1627);
nor U3766 (N_3766,In_1592,In_1999);
or U3767 (N_3767,In_464,In_24);
xor U3768 (N_3768,In_619,In_1070);
xnor U3769 (N_3769,In_1519,In_925);
nor U3770 (N_3770,In_1537,In_1701);
or U3771 (N_3771,In_34,In_175);
nand U3772 (N_3772,In_296,In_849);
nand U3773 (N_3773,In_1887,In_1294);
nor U3774 (N_3774,In_767,In_756);
xnor U3775 (N_3775,In_702,In_1163);
or U3776 (N_3776,In_968,In_1889);
nand U3777 (N_3777,In_790,In_154);
xnor U3778 (N_3778,In_656,In_1420);
and U3779 (N_3779,In_1320,In_1883);
and U3780 (N_3780,In_1500,In_473);
or U3781 (N_3781,In_918,In_434);
nor U3782 (N_3782,In_592,In_230);
nor U3783 (N_3783,In_138,In_1554);
and U3784 (N_3784,In_38,In_380);
nor U3785 (N_3785,In_790,In_39);
xnor U3786 (N_3786,In_1324,In_583);
or U3787 (N_3787,In_814,In_994);
xor U3788 (N_3788,In_1719,In_1586);
nor U3789 (N_3789,In_1818,In_859);
nor U3790 (N_3790,In_1913,In_1849);
nor U3791 (N_3791,In_1662,In_1572);
xor U3792 (N_3792,In_1952,In_1632);
or U3793 (N_3793,In_1118,In_280);
nor U3794 (N_3794,In_66,In_1596);
nand U3795 (N_3795,In_1587,In_1030);
xor U3796 (N_3796,In_653,In_1582);
and U3797 (N_3797,In_1094,In_537);
nand U3798 (N_3798,In_437,In_1131);
nand U3799 (N_3799,In_1017,In_1761);
and U3800 (N_3800,In_1285,In_104);
xnor U3801 (N_3801,In_1136,In_422);
or U3802 (N_3802,In_1675,In_1248);
xnor U3803 (N_3803,In_800,In_1441);
nor U3804 (N_3804,In_1805,In_1814);
nor U3805 (N_3805,In_739,In_59);
nand U3806 (N_3806,In_963,In_1822);
and U3807 (N_3807,In_321,In_1389);
nand U3808 (N_3808,In_1123,In_77);
xor U3809 (N_3809,In_231,In_29);
xnor U3810 (N_3810,In_414,In_1041);
nand U3811 (N_3811,In_1237,In_1219);
and U3812 (N_3812,In_1934,In_85);
xnor U3813 (N_3813,In_110,In_1324);
and U3814 (N_3814,In_1145,In_1310);
and U3815 (N_3815,In_479,In_388);
xnor U3816 (N_3816,In_567,In_1400);
and U3817 (N_3817,In_75,In_420);
nor U3818 (N_3818,In_1930,In_621);
xor U3819 (N_3819,In_1177,In_725);
xnor U3820 (N_3820,In_605,In_1550);
xnor U3821 (N_3821,In_407,In_1756);
nor U3822 (N_3822,In_592,In_654);
nor U3823 (N_3823,In_1847,In_1007);
xnor U3824 (N_3824,In_322,In_1321);
or U3825 (N_3825,In_759,In_678);
xnor U3826 (N_3826,In_1634,In_1058);
nor U3827 (N_3827,In_886,In_1427);
and U3828 (N_3828,In_763,In_1343);
xor U3829 (N_3829,In_1539,In_706);
and U3830 (N_3830,In_541,In_437);
nand U3831 (N_3831,In_1395,In_927);
or U3832 (N_3832,In_1698,In_1174);
and U3833 (N_3833,In_1136,In_1202);
nor U3834 (N_3834,In_1010,In_1809);
or U3835 (N_3835,In_715,In_1895);
nor U3836 (N_3836,In_127,In_440);
nor U3837 (N_3837,In_734,In_1527);
xnor U3838 (N_3838,In_670,In_1716);
nor U3839 (N_3839,In_1726,In_420);
nand U3840 (N_3840,In_316,In_887);
nor U3841 (N_3841,In_1025,In_1488);
nand U3842 (N_3842,In_1304,In_973);
nor U3843 (N_3843,In_1193,In_998);
xor U3844 (N_3844,In_1400,In_164);
and U3845 (N_3845,In_1607,In_718);
nand U3846 (N_3846,In_429,In_638);
or U3847 (N_3847,In_1436,In_249);
and U3848 (N_3848,In_1460,In_521);
or U3849 (N_3849,In_1305,In_1151);
xnor U3850 (N_3850,In_904,In_248);
and U3851 (N_3851,In_1558,In_1798);
and U3852 (N_3852,In_1719,In_1837);
nand U3853 (N_3853,In_14,In_892);
nand U3854 (N_3854,In_558,In_645);
nand U3855 (N_3855,In_135,In_1320);
and U3856 (N_3856,In_266,In_317);
nor U3857 (N_3857,In_740,In_982);
and U3858 (N_3858,In_1278,In_1427);
nand U3859 (N_3859,In_1497,In_82);
xor U3860 (N_3860,In_1867,In_424);
and U3861 (N_3861,In_1705,In_713);
or U3862 (N_3862,In_2,In_765);
or U3863 (N_3863,In_477,In_938);
and U3864 (N_3864,In_1417,In_1156);
or U3865 (N_3865,In_644,In_1009);
nand U3866 (N_3866,In_1056,In_1289);
nor U3867 (N_3867,In_1458,In_1463);
and U3868 (N_3868,In_1367,In_1974);
nand U3869 (N_3869,In_514,In_1834);
or U3870 (N_3870,In_358,In_642);
xnor U3871 (N_3871,In_795,In_423);
and U3872 (N_3872,In_755,In_1440);
nor U3873 (N_3873,In_1469,In_1189);
xnor U3874 (N_3874,In_449,In_783);
or U3875 (N_3875,In_1579,In_1168);
nor U3876 (N_3876,In_687,In_999);
xor U3877 (N_3877,In_710,In_1613);
nand U3878 (N_3878,In_1483,In_647);
and U3879 (N_3879,In_1174,In_1991);
xnor U3880 (N_3880,In_1901,In_41);
nand U3881 (N_3881,In_892,In_242);
xor U3882 (N_3882,In_26,In_1172);
xor U3883 (N_3883,In_1705,In_1123);
nand U3884 (N_3884,In_1202,In_1281);
nand U3885 (N_3885,In_1097,In_158);
xor U3886 (N_3886,In_1121,In_503);
and U3887 (N_3887,In_1065,In_1203);
xnor U3888 (N_3888,In_1725,In_127);
xor U3889 (N_3889,In_1967,In_714);
or U3890 (N_3890,In_1403,In_991);
xor U3891 (N_3891,In_1621,In_1217);
xnor U3892 (N_3892,In_650,In_758);
nor U3893 (N_3893,In_1775,In_1271);
xnor U3894 (N_3894,In_764,In_1138);
nand U3895 (N_3895,In_103,In_361);
and U3896 (N_3896,In_224,In_1967);
nand U3897 (N_3897,In_1831,In_1796);
nor U3898 (N_3898,In_353,In_923);
nor U3899 (N_3899,In_274,In_1298);
xnor U3900 (N_3900,In_62,In_1565);
xnor U3901 (N_3901,In_1439,In_709);
xor U3902 (N_3902,In_1343,In_998);
or U3903 (N_3903,In_724,In_915);
nand U3904 (N_3904,In_1957,In_1736);
nand U3905 (N_3905,In_1664,In_215);
nand U3906 (N_3906,In_801,In_747);
and U3907 (N_3907,In_910,In_1103);
or U3908 (N_3908,In_1333,In_921);
nor U3909 (N_3909,In_624,In_529);
nor U3910 (N_3910,In_470,In_900);
nand U3911 (N_3911,In_332,In_505);
nand U3912 (N_3912,In_1198,In_1021);
nor U3913 (N_3913,In_854,In_518);
and U3914 (N_3914,In_1506,In_293);
nand U3915 (N_3915,In_1941,In_997);
and U3916 (N_3916,In_1063,In_1209);
nor U3917 (N_3917,In_1381,In_1347);
nor U3918 (N_3918,In_1518,In_157);
xor U3919 (N_3919,In_738,In_194);
nand U3920 (N_3920,In_1362,In_50);
nand U3921 (N_3921,In_705,In_743);
nor U3922 (N_3922,In_739,In_1934);
or U3923 (N_3923,In_1907,In_1806);
xor U3924 (N_3924,In_374,In_901);
or U3925 (N_3925,In_662,In_640);
xnor U3926 (N_3926,In_417,In_326);
xor U3927 (N_3927,In_1122,In_764);
nor U3928 (N_3928,In_1028,In_81);
xnor U3929 (N_3929,In_344,In_763);
nor U3930 (N_3930,In_456,In_1921);
and U3931 (N_3931,In_936,In_849);
xnor U3932 (N_3932,In_1215,In_1727);
xnor U3933 (N_3933,In_859,In_1209);
nand U3934 (N_3934,In_313,In_1992);
xnor U3935 (N_3935,In_88,In_1381);
or U3936 (N_3936,In_1137,In_816);
nand U3937 (N_3937,In_564,In_1438);
or U3938 (N_3938,In_1902,In_1736);
nand U3939 (N_3939,In_1202,In_1609);
or U3940 (N_3940,In_1957,In_1556);
and U3941 (N_3941,In_80,In_651);
nand U3942 (N_3942,In_324,In_1409);
xor U3943 (N_3943,In_1341,In_870);
or U3944 (N_3944,In_1329,In_183);
xnor U3945 (N_3945,In_860,In_1916);
xor U3946 (N_3946,In_629,In_1074);
and U3947 (N_3947,In_200,In_1101);
nand U3948 (N_3948,In_517,In_609);
xor U3949 (N_3949,In_1412,In_894);
xnor U3950 (N_3950,In_240,In_756);
and U3951 (N_3951,In_615,In_944);
nor U3952 (N_3952,In_336,In_586);
nor U3953 (N_3953,In_1082,In_154);
nor U3954 (N_3954,In_1087,In_742);
nand U3955 (N_3955,In_1701,In_395);
xor U3956 (N_3956,In_646,In_1144);
or U3957 (N_3957,In_1696,In_150);
xnor U3958 (N_3958,In_1805,In_382);
xor U3959 (N_3959,In_383,In_1894);
and U3960 (N_3960,In_1668,In_274);
xor U3961 (N_3961,In_131,In_1928);
xor U3962 (N_3962,In_885,In_1329);
xnor U3963 (N_3963,In_1276,In_139);
nor U3964 (N_3964,In_675,In_1037);
and U3965 (N_3965,In_639,In_1661);
nand U3966 (N_3966,In_1802,In_1293);
or U3967 (N_3967,In_730,In_1833);
xor U3968 (N_3968,In_1894,In_562);
or U3969 (N_3969,In_408,In_1675);
xnor U3970 (N_3970,In_897,In_27);
xnor U3971 (N_3971,In_461,In_542);
or U3972 (N_3972,In_1266,In_1288);
xnor U3973 (N_3973,In_1427,In_1894);
or U3974 (N_3974,In_981,In_1444);
or U3975 (N_3975,In_882,In_347);
nor U3976 (N_3976,In_126,In_161);
nor U3977 (N_3977,In_1987,In_1718);
nor U3978 (N_3978,In_188,In_1107);
or U3979 (N_3979,In_899,In_320);
or U3980 (N_3980,In_1565,In_1974);
and U3981 (N_3981,In_933,In_630);
or U3982 (N_3982,In_792,In_1448);
xor U3983 (N_3983,In_588,In_1085);
or U3984 (N_3984,In_134,In_1804);
nor U3985 (N_3985,In_1456,In_1959);
nand U3986 (N_3986,In_120,In_1505);
xor U3987 (N_3987,In_990,In_138);
or U3988 (N_3988,In_60,In_1150);
and U3989 (N_3989,In_1632,In_497);
and U3990 (N_3990,In_1873,In_1206);
or U3991 (N_3991,In_1997,In_644);
or U3992 (N_3992,In_137,In_1714);
or U3993 (N_3993,In_549,In_630);
or U3994 (N_3994,In_1131,In_1620);
nand U3995 (N_3995,In_1609,In_411);
or U3996 (N_3996,In_244,In_1516);
nor U3997 (N_3997,In_659,In_1555);
or U3998 (N_3998,In_285,In_1861);
nand U3999 (N_3999,In_1765,In_951);
xor U4000 (N_4000,In_1389,In_217);
and U4001 (N_4001,In_1772,In_931);
and U4002 (N_4002,In_744,In_1866);
and U4003 (N_4003,In_653,In_224);
nor U4004 (N_4004,In_1955,In_1913);
or U4005 (N_4005,In_450,In_125);
or U4006 (N_4006,In_1912,In_1734);
or U4007 (N_4007,In_1597,In_1593);
xor U4008 (N_4008,In_1055,In_683);
and U4009 (N_4009,In_417,In_1434);
nand U4010 (N_4010,In_1082,In_1956);
xnor U4011 (N_4011,In_1985,In_52);
and U4012 (N_4012,In_1199,In_1299);
or U4013 (N_4013,In_384,In_1643);
and U4014 (N_4014,In_416,In_75);
xnor U4015 (N_4015,In_1682,In_1861);
nor U4016 (N_4016,In_1325,In_1067);
or U4017 (N_4017,In_234,In_1928);
or U4018 (N_4018,In_1232,In_1933);
or U4019 (N_4019,In_1474,In_1454);
nor U4020 (N_4020,In_1977,In_930);
nor U4021 (N_4021,In_110,In_321);
xnor U4022 (N_4022,In_156,In_126);
xor U4023 (N_4023,In_1901,In_1062);
nor U4024 (N_4024,In_1508,In_1289);
xor U4025 (N_4025,In_1473,In_695);
and U4026 (N_4026,In_933,In_1068);
nor U4027 (N_4027,In_1947,In_951);
nand U4028 (N_4028,In_53,In_656);
or U4029 (N_4029,In_1220,In_1950);
nand U4030 (N_4030,In_444,In_120);
nand U4031 (N_4031,In_410,In_225);
nand U4032 (N_4032,In_993,In_425);
nor U4033 (N_4033,In_669,In_795);
nand U4034 (N_4034,In_1850,In_822);
xnor U4035 (N_4035,In_20,In_37);
nor U4036 (N_4036,In_596,In_1066);
nand U4037 (N_4037,In_3,In_1790);
or U4038 (N_4038,In_858,In_265);
xor U4039 (N_4039,In_1336,In_428);
xnor U4040 (N_4040,In_646,In_738);
or U4041 (N_4041,In_515,In_765);
and U4042 (N_4042,In_297,In_578);
nor U4043 (N_4043,In_411,In_702);
xor U4044 (N_4044,In_1369,In_295);
or U4045 (N_4045,In_53,In_601);
nor U4046 (N_4046,In_246,In_1438);
nand U4047 (N_4047,In_1944,In_489);
or U4048 (N_4048,In_1085,In_83);
xor U4049 (N_4049,In_572,In_1481);
xnor U4050 (N_4050,In_1023,In_1162);
or U4051 (N_4051,In_864,In_1119);
nand U4052 (N_4052,In_1247,In_1467);
nand U4053 (N_4053,In_1775,In_1627);
xor U4054 (N_4054,In_1477,In_1724);
nor U4055 (N_4055,In_1990,In_749);
nand U4056 (N_4056,In_708,In_240);
nor U4057 (N_4057,In_448,In_1897);
and U4058 (N_4058,In_1940,In_1620);
nor U4059 (N_4059,In_1732,In_1274);
xnor U4060 (N_4060,In_489,In_738);
nand U4061 (N_4061,In_515,In_324);
or U4062 (N_4062,In_251,In_980);
or U4063 (N_4063,In_804,In_1465);
xor U4064 (N_4064,In_780,In_1554);
and U4065 (N_4065,In_1214,In_849);
nand U4066 (N_4066,In_1141,In_927);
xor U4067 (N_4067,In_1232,In_1550);
nor U4068 (N_4068,In_1966,In_1105);
or U4069 (N_4069,In_52,In_1775);
nand U4070 (N_4070,In_1272,In_1129);
nand U4071 (N_4071,In_1876,In_141);
or U4072 (N_4072,In_1736,In_135);
nand U4073 (N_4073,In_1484,In_670);
and U4074 (N_4074,In_904,In_410);
nor U4075 (N_4075,In_734,In_940);
and U4076 (N_4076,In_1626,In_1485);
nand U4077 (N_4077,In_855,In_1002);
xnor U4078 (N_4078,In_1284,In_1084);
nor U4079 (N_4079,In_1824,In_1466);
and U4080 (N_4080,In_1187,In_1783);
or U4081 (N_4081,In_1219,In_177);
and U4082 (N_4082,In_1591,In_260);
nand U4083 (N_4083,In_133,In_1050);
nand U4084 (N_4084,In_115,In_1670);
nor U4085 (N_4085,In_937,In_133);
nand U4086 (N_4086,In_48,In_1999);
xor U4087 (N_4087,In_338,In_548);
or U4088 (N_4088,In_1812,In_756);
or U4089 (N_4089,In_1161,In_1053);
nand U4090 (N_4090,In_206,In_1578);
nor U4091 (N_4091,In_97,In_1097);
and U4092 (N_4092,In_1976,In_1919);
nor U4093 (N_4093,In_130,In_524);
xnor U4094 (N_4094,In_1157,In_762);
nand U4095 (N_4095,In_155,In_284);
xnor U4096 (N_4096,In_1894,In_1997);
nand U4097 (N_4097,In_687,In_54);
xor U4098 (N_4098,In_1549,In_216);
xnor U4099 (N_4099,In_479,In_966);
xnor U4100 (N_4100,In_1484,In_1892);
xor U4101 (N_4101,In_1164,In_1722);
nor U4102 (N_4102,In_958,In_1806);
xor U4103 (N_4103,In_1559,In_914);
and U4104 (N_4104,In_738,In_23);
xnor U4105 (N_4105,In_1531,In_1822);
or U4106 (N_4106,In_55,In_639);
xnor U4107 (N_4107,In_1809,In_1893);
and U4108 (N_4108,In_1304,In_937);
xor U4109 (N_4109,In_1633,In_346);
nand U4110 (N_4110,In_655,In_584);
and U4111 (N_4111,In_1640,In_1001);
xor U4112 (N_4112,In_1134,In_1534);
nand U4113 (N_4113,In_1621,In_1583);
or U4114 (N_4114,In_1120,In_1889);
nor U4115 (N_4115,In_1678,In_1417);
xnor U4116 (N_4116,In_1283,In_1694);
or U4117 (N_4117,In_1097,In_1611);
nor U4118 (N_4118,In_1604,In_932);
or U4119 (N_4119,In_71,In_1791);
nand U4120 (N_4120,In_642,In_1043);
nand U4121 (N_4121,In_203,In_1538);
and U4122 (N_4122,In_1637,In_1415);
nor U4123 (N_4123,In_1936,In_530);
nand U4124 (N_4124,In_613,In_297);
or U4125 (N_4125,In_1404,In_1752);
or U4126 (N_4126,In_1106,In_993);
xnor U4127 (N_4127,In_1658,In_290);
nand U4128 (N_4128,In_342,In_641);
nand U4129 (N_4129,In_156,In_49);
and U4130 (N_4130,In_821,In_787);
and U4131 (N_4131,In_1244,In_1266);
or U4132 (N_4132,In_68,In_1607);
nand U4133 (N_4133,In_1253,In_604);
nand U4134 (N_4134,In_481,In_1150);
nor U4135 (N_4135,In_256,In_1000);
xnor U4136 (N_4136,In_182,In_1085);
nor U4137 (N_4137,In_1592,In_1958);
nor U4138 (N_4138,In_1195,In_425);
or U4139 (N_4139,In_384,In_478);
nor U4140 (N_4140,In_1059,In_86);
nand U4141 (N_4141,In_781,In_43);
nor U4142 (N_4142,In_1875,In_1748);
nor U4143 (N_4143,In_813,In_1277);
xnor U4144 (N_4144,In_836,In_917);
and U4145 (N_4145,In_515,In_26);
xnor U4146 (N_4146,In_242,In_956);
or U4147 (N_4147,In_261,In_1659);
xnor U4148 (N_4148,In_422,In_589);
nand U4149 (N_4149,In_1420,In_1451);
nor U4150 (N_4150,In_385,In_437);
xnor U4151 (N_4151,In_1049,In_1625);
and U4152 (N_4152,In_42,In_1522);
nor U4153 (N_4153,In_556,In_596);
nor U4154 (N_4154,In_1981,In_1606);
nor U4155 (N_4155,In_31,In_1226);
nand U4156 (N_4156,In_1155,In_1978);
nor U4157 (N_4157,In_1568,In_141);
and U4158 (N_4158,In_201,In_1072);
nor U4159 (N_4159,In_1849,In_1642);
and U4160 (N_4160,In_797,In_1566);
or U4161 (N_4161,In_936,In_1111);
and U4162 (N_4162,In_813,In_1276);
or U4163 (N_4163,In_362,In_407);
xor U4164 (N_4164,In_1717,In_1668);
nand U4165 (N_4165,In_1074,In_1246);
nor U4166 (N_4166,In_205,In_1796);
nand U4167 (N_4167,In_1001,In_646);
or U4168 (N_4168,In_538,In_326);
or U4169 (N_4169,In_1369,In_194);
nand U4170 (N_4170,In_69,In_222);
or U4171 (N_4171,In_50,In_1987);
xnor U4172 (N_4172,In_1272,In_1992);
or U4173 (N_4173,In_401,In_499);
nor U4174 (N_4174,In_1857,In_1730);
and U4175 (N_4175,In_1709,In_48);
xor U4176 (N_4176,In_118,In_1483);
nor U4177 (N_4177,In_880,In_938);
nand U4178 (N_4178,In_1365,In_1284);
nand U4179 (N_4179,In_357,In_1554);
nor U4180 (N_4180,In_1040,In_560);
and U4181 (N_4181,In_1245,In_544);
nand U4182 (N_4182,In_1554,In_1067);
nor U4183 (N_4183,In_636,In_883);
and U4184 (N_4184,In_1354,In_543);
and U4185 (N_4185,In_1631,In_965);
or U4186 (N_4186,In_828,In_223);
xor U4187 (N_4187,In_1150,In_1074);
nor U4188 (N_4188,In_476,In_423);
nor U4189 (N_4189,In_1463,In_1572);
nand U4190 (N_4190,In_1126,In_263);
xnor U4191 (N_4191,In_837,In_503);
and U4192 (N_4192,In_513,In_487);
xor U4193 (N_4193,In_1539,In_1523);
and U4194 (N_4194,In_743,In_449);
nor U4195 (N_4195,In_1104,In_973);
nor U4196 (N_4196,In_876,In_402);
or U4197 (N_4197,In_817,In_1458);
nand U4198 (N_4198,In_321,In_307);
nor U4199 (N_4199,In_263,In_1794);
and U4200 (N_4200,In_15,In_1840);
xor U4201 (N_4201,In_288,In_234);
nor U4202 (N_4202,In_581,In_1745);
nand U4203 (N_4203,In_525,In_613);
nor U4204 (N_4204,In_269,In_1698);
nand U4205 (N_4205,In_196,In_208);
nor U4206 (N_4206,In_1264,In_487);
or U4207 (N_4207,In_332,In_1104);
or U4208 (N_4208,In_105,In_646);
xnor U4209 (N_4209,In_1558,In_55);
nor U4210 (N_4210,In_556,In_1542);
xor U4211 (N_4211,In_672,In_429);
and U4212 (N_4212,In_1556,In_382);
xor U4213 (N_4213,In_817,In_1021);
nor U4214 (N_4214,In_438,In_1573);
xnor U4215 (N_4215,In_1023,In_134);
xor U4216 (N_4216,In_73,In_1858);
xnor U4217 (N_4217,In_235,In_1244);
nor U4218 (N_4218,In_1134,In_83);
and U4219 (N_4219,In_1947,In_229);
nand U4220 (N_4220,In_1581,In_1874);
nor U4221 (N_4221,In_473,In_186);
nor U4222 (N_4222,In_1950,In_159);
and U4223 (N_4223,In_555,In_476);
xor U4224 (N_4224,In_1968,In_38);
xor U4225 (N_4225,In_90,In_1251);
nand U4226 (N_4226,In_344,In_120);
and U4227 (N_4227,In_1445,In_479);
nand U4228 (N_4228,In_915,In_612);
and U4229 (N_4229,In_889,In_695);
and U4230 (N_4230,In_464,In_383);
nand U4231 (N_4231,In_933,In_1635);
nand U4232 (N_4232,In_674,In_417);
and U4233 (N_4233,In_364,In_1721);
xnor U4234 (N_4234,In_1912,In_0);
nand U4235 (N_4235,In_1104,In_410);
xor U4236 (N_4236,In_210,In_1342);
and U4237 (N_4237,In_1872,In_1531);
xor U4238 (N_4238,In_1325,In_331);
or U4239 (N_4239,In_545,In_771);
xor U4240 (N_4240,In_1992,In_941);
or U4241 (N_4241,In_791,In_233);
nand U4242 (N_4242,In_883,In_791);
xnor U4243 (N_4243,In_427,In_1372);
nor U4244 (N_4244,In_1561,In_1424);
or U4245 (N_4245,In_917,In_1055);
or U4246 (N_4246,In_1678,In_407);
or U4247 (N_4247,In_81,In_1283);
and U4248 (N_4248,In_1813,In_516);
xnor U4249 (N_4249,In_646,In_1374);
nor U4250 (N_4250,In_1629,In_1336);
xnor U4251 (N_4251,In_839,In_358);
or U4252 (N_4252,In_773,In_768);
nor U4253 (N_4253,In_1587,In_719);
and U4254 (N_4254,In_918,In_1846);
xnor U4255 (N_4255,In_654,In_842);
xnor U4256 (N_4256,In_953,In_447);
nand U4257 (N_4257,In_1490,In_873);
xor U4258 (N_4258,In_1583,In_710);
and U4259 (N_4259,In_583,In_1400);
nor U4260 (N_4260,In_337,In_1223);
nor U4261 (N_4261,In_200,In_1491);
nor U4262 (N_4262,In_1752,In_635);
xnor U4263 (N_4263,In_622,In_897);
or U4264 (N_4264,In_1275,In_391);
nand U4265 (N_4265,In_1126,In_480);
or U4266 (N_4266,In_942,In_1139);
nand U4267 (N_4267,In_1355,In_76);
nor U4268 (N_4268,In_1640,In_1795);
nand U4269 (N_4269,In_206,In_569);
nand U4270 (N_4270,In_851,In_1689);
and U4271 (N_4271,In_413,In_353);
and U4272 (N_4272,In_1241,In_541);
nor U4273 (N_4273,In_1596,In_232);
nor U4274 (N_4274,In_1868,In_1211);
xnor U4275 (N_4275,In_745,In_1785);
xor U4276 (N_4276,In_923,In_1419);
nor U4277 (N_4277,In_1971,In_28);
and U4278 (N_4278,In_750,In_961);
nand U4279 (N_4279,In_60,In_137);
xor U4280 (N_4280,In_1564,In_948);
and U4281 (N_4281,In_755,In_1135);
nand U4282 (N_4282,In_587,In_1374);
nand U4283 (N_4283,In_1169,In_569);
nand U4284 (N_4284,In_1630,In_1717);
nor U4285 (N_4285,In_718,In_1747);
nor U4286 (N_4286,In_1968,In_1972);
nand U4287 (N_4287,In_717,In_492);
nand U4288 (N_4288,In_1247,In_1635);
nor U4289 (N_4289,In_1443,In_1562);
or U4290 (N_4290,In_1287,In_1070);
xnor U4291 (N_4291,In_456,In_707);
or U4292 (N_4292,In_1155,In_1561);
xnor U4293 (N_4293,In_1657,In_63);
nand U4294 (N_4294,In_933,In_798);
and U4295 (N_4295,In_939,In_687);
nor U4296 (N_4296,In_646,In_1054);
nor U4297 (N_4297,In_1727,In_565);
xnor U4298 (N_4298,In_1046,In_1239);
nand U4299 (N_4299,In_1295,In_1640);
nor U4300 (N_4300,In_1235,In_972);
nor U4301 (N_4301,In_216,In_964);
nand U4302 (N_4302,In_652,In_1525);
or U4303 (N_4303,In_1212,In_385);
nand U4304 (N_4304,In_139,In_1796);
and U4305 (N_4305,In_1054,In_1050);
and U4306 (N_4306,In_348,In_1614);
or U4307 (N_4307,In_1817,In_2);
nor U4308 (N_4308,In_1798,In_91);
and U4309 (N_4309,In_1213,In_1090);
nor U4310 (N_4310,In_1937,In_1173);
and U4311 (N_4311,In_460,In_178);
nor U4312 (N_4312,In_283,In_538);
and U4313 (N_4313,In_990,In_584);
and U4314 (N_4314,In_104,In_726);
or U4315 (N_4315,In_1729,In_1663);
or U4316 (N_4316,In_1247,In_203);
nor U4317 (N_4317,In_387,In_1182);
nand U4318 (N_4318,In_1411,In_1497);
or U4319 (N_4319,In_454,In_1992);
xnor U4320 (N_4320,In_938,In_1027);
xor U4321 (N_4321,In_1339,In_872);
and U4322 (N_4322,In_129,In_854);
xor U4323 (N_4323,In_161,In_1035);
nand U4324 (N_4324,In_1360,In_244);
nor U4325 (N_4325,In_87,In_1313);
or U4326 (N_4326,In_298,In_1955);
and U4327 (N_4327,In_897,In_1300);
xnor U4328 (N_4328,In_1712,In_1547);
nand U4329 (N_4329,In_1279,In_439);
nor U4330 (N_4330,In_687,In_347);
nand U4331 (N_4331,In_168,In_1647);
and U4332 (N_4332,In_856,In_210);
or U4333 (N_4333,In_1802,In_487);
nand U4334 (N_4334,In_329,In_1475);
and U4335 (N_4335,In_109,In_1328);
nor U4336 (N_4336,In_1712,In_655);
xnor U4337 (N_4337,In_1222,In_1954);
and U4338 (N_4338,In_379,In_395);
xnor U4339 (N_4339,In_1181,In_261);
xor U4340 (N_4340,In_605,In_1894);
or U4341 (N_4341,In_1288,In_625);
nand U4342 (N_4342,In_1035,In_649);
xor U4343 (N_4343,In_282,In_731);
nor U4344 (N_4344,In_1591,In_197);
and U4345 (N_4345,In_1875,In_997);
or U4346 (N_4346,In_21,In_129);
and U4347 (N_4347,In_278,In_1736);
or U4348 (N_4348,In_211,In_1782);
and U4349 (N_4349,In_1714,In_1631);
nand U4350 (N_4350,In_1771,In_1941);
nand U4351 (N_4351,In_965,In_1756);
nor U4352 (N_4352,In_1366,In_1780);
nand U4353 (N_4353,In_63,In_1033);
nand U4354 (N_4354,In_1445,In_1303);
or U4355 (N_4355,In_32,In_1056);
nor U4356 (N_4356,In_1439,In_359);
nand U4357 (N_4357,In_575,In_233);
nor U4358 (N_4358,In_1683,In_463);
and U4359 (N_4359,In_1575,In_1047);
xor U4360 (N_4360,In_1717,In_440);
or U4361 (N_4361,In_1610,In_226);
and U4362 (N_4362,In_391,In_1628);
xnor U4363 (N_4363,In_1971,In_816);
nand U4364 (N_4364,In_848,In_1132);
nand U4365 (N_4365,In_1014,In_1104);
and U4366 (N_4366,In_163,In_574);
nand U4367 (N_4367,In_844,In_487);
nor U4368 (N_4368,In_799,In_174);
nor U4369 (N_4369,In_521,In_727);
nor U4370 (N_4370,In_1667,In_654);
nor U4371 (N_4371,In_1109,In_1331);
nor U4372 (N_4372,In_31,In_139);
or U4373 (N_4373,In_1444,In_685);
nor U4374 (N_4374,In_1102,In_1389);
nand U4375 (N_4375,In_1668,In_254);
and U4376 (N_4376,In_1111,In_1153);
xnor U4377 (N_4377,In_356,In_80);
nor U4378 (N_4378,In_901,In_576);
and U4379 (N_4379,In_512,In_519);
and U4380 (N_4380,In_1590,In_198);
nand U4381 (N_4381,In_1740,In_393);
nor U4382 (N_4382,In_1937,In_274);
or U4383 (N_4383,In_1031,In_1004);
and U4384 (N_4384,In_836,In_248);
nand U4385 (N_4385,In_1902,In_611);
or U4386 (N_4386,In_208,In_932);
nand U4387 (N_4387,In_1960,In_739);
nand U4388 (N_4388,In_1926,In_415);
xor U4389 (N_4389,In_1969,In_1364);
xnor U4390 (N_4390,In_1800,In_1523);
and U4391 (N_4391,In_1994,In_971);
xor U4392 (N_4392,In_1312,In_750);
or U4393 (N_4393,In_902,In_495);
nor U4394 (N_4394,In_1121,In_1654);
xnor U4395 (N_4395,In_591,In_1202);
nand U4396 (N_4396,In_1936,In_39);
nor U4397 (N_4397,In_738,In_363);
and U4398 (N_4398,In_1569,In_1437);
xnor U4399 (N_4399,In_64,In_222);
or U4400 (N_4400,In_1711,In_1910);
and U4401 (N_4401,In_1507,In_93);
or U4402 (N_4402,In_520,In_1103);
nand U4403 (N_4403,In_1967,In_870);
nor U4404 (N_4404,In_1482,In_714);
xor U4405 (N_4405,In_1805,In_602);
and U4406 (N_4406,In_960,In_1573);
nand U4407 (N_4407,In_310,In_980);
xor U4408 (N_4408,In_1725,In_1238);
nand U4409 (N_4409,In_523,In_441);
nand U4410 (N_4410,In_997,In_246);
nand U4411 (N_4411,In_13,In_1323);
and U4412 (N_4412,In_475,In_1352);
xor U4413 (N_4413,In_1451,In_1808);
nand U4414 (N_4414,In_521,In_1704);
nor U4415 (N_4415,In_337,In_1396);
nor U4416 (N_4416,In_1700,In_1896);
nand U4417 (N_4417,In_1867,In_1106);
and U4418 (N_4418,In_122,In_1907);
and U4419 (N_4419,In_1310,In_1711);
and U4420 (N_4420,In_1303,In_1759);
or U4421 (N_4421,In_1455,In_307);
nor U4422 (N_4422,In_706,In_626);
or U4423 (N_4423,In_1132,In_1934);
nor U4424 (N_4424,In_1927,In_927);
xor U4425 (N_4425,In_329,In_540);
nor U4426 (N_4426,In_1428,In_627);
and U4427 (N_4427,In_1993,In_938);
nand U4428 (N_4428,In_1165,In_1715);
nor U4429 (N_4429,In_1686,In_1702);
nor U4430 (N_4430,In_831,In_23);
xor U4431 (N_4431,In_1781,In_452);
xor U4432 (N_4432,In_729,In_42);
or U4433 (N_4433,In_794,In_1308);
or U4434 (N_4434,In_952,In_651);
nor U4435 (N_4435,In_1633,In_1450);
nand U4436 (N_4436,In_1459,In_1231);
xnor U4437 (N_4437,In_1182,In_1681);
nand U4438 (N_4438,In_1778,In_133);
xor U4439 (N_4439,In_424,In_1435);
nand U4440 (N_4440,In_1751,In_410);
nor U4441 (N_4441,In_7,In_306);
and U4442 (N_4442,In_37,In_478);
nand U4443 (N_4443,In_847,In_1911);
xnor U4444 (N_4444,In_924,In_723);
or U4445 (N_4445,In_1518,In_1181);
or U4446 (N_4446,In_984,In_943);
or U4447 (N_4447,In_969,In_307);
xnor U4448 (N_4448,In_1471,In_1049);
nor U4449 (N_4449,In_1440,In_1625);
or U4450 (N_4450,In_332,In_719);
nor U4451 (N_4451,In_1876,In_628);
xor U4452 (N_4452,In_1114,In_1882);
or U4453 (N_4453,In_1517,In_1751);
xor U4454 (N_4454,In_1903,In_59);
xnor U4455 (N_4455,In_1025,In_1095);
xor U4456 (N_4456,In_606,In_1498);
or U4457 (N_4457,In_1610,In_1362);
and U4458 (N_4458,In_1207,In_761);
xor U4459 (N_4459,In_1561,In_1905);
nor U4460 (N_4460,In_1007,In_716);
and U4461 (N_4461,In_1595,In_1342);
and U4462 (N_4462,In_1703,In_1675);
xor U4463 (N_4463,In_150,In_670);
nand U4464 (N_4464,In_1960,In_1498);
or U4465 (N_4465,In_1127,In_1678);
nor U4466 (N_4466,In_715,In_1496);
and U4467 (N_4467,In_1271,In_1908);
or U4468 (N_4468,In_562,In_615);
nor U4469 (N_4469,In_1989,In_346);
or U4470 (N_4470,In_1936,In_992);
and U4471 (N_4471,In_791,In_1124);
and U4472 (N_4472,In_1916,In_890);
nand U4473 (N_4473,In_1328,In_1181);
or U4474 (N_4474,In_266,In_1888);
or U4475 (N_4475,In_1637,In_1511);
xnor U4476 (N_4476,In_1964,In_174);
xnor U4477 (N_4477,In_1587,In_1791);
and U4478 (N_4478,In_698,In_1520);
xor U4479 (N_4479,In_1862,In_1043);
and U4480 (N_4480,In_1073,In_1293);
nand U4481 (N_4481,In_1020,In_1069);
nand U4482 (N_4482,In_644,In_1844);
nor U4483 (N_4483,In_474,In_35);
nand U4484 (N_4484,In_1888,In_552);
nor U4485 (N_4485,In_278,In_1618);
nand U4486 (N_4486,In_811,In_1270);
xnor U4487 (N_4487,In_1499,In_1244);
nor U4488 (N_4488,In_1447,In_754);
xnor U4489 (N_4489,In_1541,In_1240);
and U4490 (N_4490,In_896,In_1090);
or U4491 (N_4491,In_1580,In_632);
nor U4492 (N_4492,In_573,In_1579);
xnor U4493 (N_4493,In_1294,In_1971);
nor U4494 (N_4494,In_710,In_967);
nor U4495 (N_4495,In_1999,In_618);
nor U4496 (N_4496,In_28,In_349);
and U4497 (N_4497,In_1881,In_1125);
or U4498 (N_4498,In_1324,In_449);
nor U4499 (N_4499,In_1941,In_1999);
and U4500 (N_4500,In_616,In_1388);
xor U4501 (N_4501,In_1862,In_222);
or U4502 (N_4502,In_711,In_590);
xor U4503 (N_4503,In_1298,In_1893);
nor U4504 (N_4504,In_703,In_944);
nor U4505 (N_4505,In_1404,In_1132);
xor U4506 (N_4506,In_1055,In_1450);
nor U4507 (N_4507,In_98,In_115);
and U4508 (N_4508,In_1926,In_152);
xnor U4509 (N_4509,In_998,In_731);
nor U4510 (N_4510,In_1279,In_1914);
and U4511 (N_4511,In_938,In_1679);
or U4512 (N_4512,In_268,In_1448);
nand U4513 (N_4513,In_1992,In_1110);
nand U4514 (N_4514,In_544,In_758);
nor U4515 (N_4515,In_712,In_679);
xor U4516 (N_4516,In_1491,In_989);
nand U4517 (N_4517,In_591,In_64);
or U4518 (N_4518,In_1020,In_1695);
or U4519 (N_4519,In_1792,In_481);
xor U4520 (N_4520,In_936,In_1343);
nor U4521 (N_4521,In_1425,In_556);
xnor U4522 (N_4522,In_927,In_212);
nor U4523 (N_4523,In_1591,In_1674);
nand U4524 (N_4524,In_646,In_1212);
nor U4525 (N_4525,In_1820,In_1231);
nor U4526 (N_4526,In_1813,In_115);
or U4527 (N_4527,In_923,In_1732);
nand U4528 (N_4528,In_332,In_108);
xnor U4529 (N_4529,In_1348,In_830);
xor U4530 (N_4530,In_1304,In_1832);
nor U4531 (N_4531,In_576,In_520);
xnor U4532 (N_4532,In_590,In_756);
and U4533 (N_4533,In_1581,In_378);
nand U4534 (N_4534,In_750,In_239);
nand U4535 (N_4535,In_1914,In_1522);
nand U4536 (N_4536,In_934,In_108);
xor U4537 (N_4537,In_381,In_1495);
and U4538 (N_4538,In_1609,In_1178);
xor U4539 (N_4539,In_1891,In_1345);
and U4540 (N_4540,In_1335,In_999);
and U4541 (N_4541,In_1203,In_799);
or U4542 (N_4542,In_1145,In_134);
or U4543 (N_4543,In_451,In_277);
and U4544 (N_4544,In_1519,In_943);
and U4545 (N_4545,In_269,In_1099);
and U4546 (N_4546,In_1513,In_995);
xor U4547 (N_4547,In_1628,In_1017);
and U4548 (N_4548,In_424,In_611);
nand U4549 (N_4549,In_292,In_873);
nor U4550 (N_4550,In_1327,In_555);
or U4551 (N_4551,In_37,In_564);
or U4552 (N_4552,In_488,In_936);
nor U4553 (N_4553,In_1718,In_271);
nand U4554 (N_4554,In_49,In_1042);
and U4555 (N_4555,In_196,In_1169);
xnor U4556 (N_4556,In_996,In_879);
xor U4557 (N_4557,In_1403,In_1352);
and U4558 (N_4558,In_1546,In_1950);
or U4559 (N_4559,In_1843,In_1524);
nand U4560 (N_4560,In_1242,In_1016);
and U4561 (N_4561,In_1477,In_1814);
nor U4562 (N_4562,In_1221,In_1413);
and U4563 (N_4563,In_1604,In_864);
xnor U4564 (N_4564,In_1970,In_664);
or U4565 (N_4565,In_1433,In_392);
and U4566 (N_4566,In_878,In_3);
nand U4567 (N_4567,In_1944,In_1102);
nor U4568 (N_4568,In_678,In_1105);
or U4569 (N_4569,In_1710,In_825);
nand U4570 (N_4570,In_1297,In_1592);
and U4571 (N_4571,In_1752,In_1855);
nand U4572 (N_4572,In_1743,In_1982);
or U4573 (N_4573,In_850,In_396);
nor U4574 (N_4574,In_931,In_840);
and U4575 (N_4575,In_1892,In_1183);
and U4576 (N_4576,In_26,In_1327);
nand U4577 (N_4577,In_1776,In_1641);
nand U4578 (N_4578,In_1786,In_1774);
and U4579 (N_4579,In_429,In_39);
xor U4580 (N_4580,In_1562,In_466);
nor U4581 (N_4581,In_1119,In_1756);
nor U4582 (N_4582,In_1262,In_671);
or U4583 (N_4583,In_685,In_736);
nand U4584 (N_4584,In_1409,In_1218);
and U4585 (N_4585,In_1578,In_345);
or U4586 (N_4586,In_780,In_1855);
xnor U4587 (N_4587,In_1753,In_35);
nor U4588 (N_4588,In_1538,In_5);
nand U4589 (N_4589,In_1978,In_549);
nand U4590 (N_4590,In_76,In_257);
or U4591 (N_4591,In_1109,In_1604);
or U4592 (N_4592,In_154,In_1219);
or U4593 (N_4593,In_24,In_1135);
or U4594 (N_4594,In_663,In_599);
nor U4595 (N_4595,In_1463,In_896);
nand U4596 (N_4596,In_1828,In_526);
nor U4597 (N_4597,In_130,In_1518);
nand U4598 (N_4598,In_1104,In_1871);
nand U4599 (N_4599,In_1204,In_990);
or U4600 (N_4600,In_1773,In_145);
and U4601 (N_4601,In_520,In_1146);
xor U4602 (N_4602,In_1032,In_1182);
or U4603 (N_4603,In_1163,In_243);
nor U4604 (N_4604,In_790,In_611);
and U4605 (N_4605,In_226,In_1074);
nor U4606 (N_4606,In_1956,In_1508);
nand U4607 (N_4607,In_1136,In_1282);
or U4608 (N_4608,In_1532,In_190);
nor U4609 (N_4609,In_1133,In_1103);
nor U4610 (N_4610,In_1024,In_979);
or U4611 (N_4611,In_1788,In_1002);
xor U4612 (N_4612,In_937,In_840);
and U4613 (N_4613,In_79,In_1452);
or U4614 (N_4614,In_1445,In_1887);
nor U4615 (N_4615,In_556,In_740);
xor U4616 (N_4616,In_1112,In_406);
or U4617 (N_4617,In_161,In_82);
nand U4618 (N_4618,In_1753,In_486);
nand U4619 (N_4619,In_1103,In_758);
xor U4620 (N_4620,In_1664,In_343);
nor U4621 (N_4621,In_1865,In_733);
nor U4622 (N_4622,In_1069,In_298);
nand U4623 (N_4623,In_823,In_1822);
and U4624 (N_4624,In_1905,In_119);
nor U4625 (N_4625,In_518,In_1541);
nand U4626 (N_4626,In_1080,In_1861);
nand U4627 (N_4627,In_1826,In_381);
and U4628 (N_4628,In_909,In_1565);
nor U4629 (N_4629,In_462,In_358);
and U4630 (N_4630,In_259,In_1865);
and U4631 (N_4631,In_589,In_504);
nor U4632 (N_4632,In_954,In_1149);
or U4633 (N_4633,In_1962,In_425);
or U4634 (N_4634,In_1442,In_1074);
nor U4635 (N_4635,In_1187,In_149);
xor U4636 (N_4636,In_1723,In_1292);
or U4637 (N_4637,In_1319,In_372);
or U4638 (N_4638,In_228,In_1282);
and U4639 (N_4639,In_1235,In_1834);
or U4640 (N_4640,In_1254,In_989);
or U4641 (N_4641,In_313,In_88);
nand U4642 (N_4642,In_1851,In_1361);
nor U4643 (N_4643,In_1611,In_330);
or U4644 (N_4644,In_675,In_1472);
nand U4645 (N_4645,In_1584,In_467);
or U4646 (N_4646,In_646,In_191);
nor U4647 (N_4647,In_354,In_312);
or U4648 (N_4648,In_14,In_1572);
nand U4649 (N_4649,In_502,In_715);
nand U4650 (N_4650,In_1173,In_115);
nand U4651 (N_4651,In_1999,In_469);
nand U4652 (N_4652,In_77,In_1208);
nor U4653 (N_4653,In_1648,In_804);
or U4654 (N_4654,In_1783,In_1869);
or U4655 (N_4655,In_1484,In_1573);
nor U4656 (N_4656,In_472,In_1329);
or U4657 (N_4657,In_548,In_363);
nor U4658 (N_4658,In_1694,In_1552);
or U4659 (N_4659,In_1527,In_240);
nor U4660 (N_4660,In_282,In_1602);
or U4661 (N_4661,In_241,In_1699);
or U4662 (N_4662,In_241,In_1270);
nor U4663 (N_4663,In_161,In_54);
nor U4664 (N_4664,In_1262,In_1644);
or U4665 (N_4665,In_1609,In_712);
nor U4666 (N_4666,In_1879,In_18);
nor U4667 (N_4667,In_1264,In_918);
nand U4668 (N_4668,In_1599,In_54);
nand U4669 (N_4669,In_561,In_796);
nand U4670 (N_4670,In_780,In_756);
xor U4671 (N_4671,In_1662,In_954);
or U4672 (N_4672,In_1475,In_937);
or U4673 (N_4673,In_1380,In_40);
and U4674 (N_4674,In_1939,In_1183);
xnor U4675 (N_4675,In_68,In_1027);
or U4676 (N_4676,In_875,In_1834);
nor U4677 (N_4677,In_960,In_23);
xnor U4678 (N_4678,In_956,In_388);
nor U4679 (N_4679,In_306,In_1028);
xnor U4680 (N_4680,In_1660,In_798);
nor U4681 (N_4681,In_288,In_1492);
and U4682 (N_4682,In_1331,In_1598);
or U4683 (N_4683,In_688,In_1952);
xnor U4684 (N_4684,In_911,In_73);
nor U4685 (N_4685,In_1412,In_528);
xor U4686 (N_4686,In_1476,In_1205);
xor U4687 (N_4687,In_327,In_1430);
xor U4688 (N_4688,In_224,In_1619);
nand U4689 (N_4689,In_1100,In_524);
nor U4690 (N_4690,In_1355,In_1873);
nand U4691 (N_4691,In_470,In_1261);
or U4692 (N_4692,In_1586,In_1129);
xor U4693 (N_4693,In_671,In_943);
nor U4694 (N_4694,In_80,In_1955);
nor U4695 (N_4695,In_935,In_451);
or U4696 (N_4696,In_1852,In_1098);
and U4697 (N_4697,In_98,In_37);
or U4698 (N_4698,In_660,In_220);
xor U4699 (N_4699,In_1382,In_1477);
nand U4700 (N_4700,In_636,In_1997);
or U4701 (N_4701,In_697,In_711);
and U4702 (N_4702,In_1097,In_65);
or U4703 (N_4703,In_1646,In_1528);
nand U4704 (N_4704,In_1353,In_556);
xor U4705 (N_4705,In_233,In_1278);
and U4706 (N_4706,In_1409,In_1969);
xnor U4707 (N_4707,In_249,In_849);
nand U4708 (N_4708,In_1339,In_1213);
nor U4709 (N_4709,In_722,In_972);
and U4710 (N_4710,In_718,In_1755);
and U4711 (N_4711,In_687,In_1844);
nand U4712 (N_4712,In_380,In_1899);
and U4713 (N_4713,In_1545,In_936);
and U4714 (N_4714,In_849,In_221);
nor U4715 (N_4715,In_1099,In_612);
or U4716 (N_4716,In_544,In_1686);
nand U4717 (N_4717,In_1200,In_885);
nand U4718 (N_4718,In_494,In_1523);
nor U4719 (N_4719,In_388,In_1755);
xor U4720 (N_4720,In_1835,In_1203);
or U4721 (N_4721,In_1960,In_79);
nand U4722 (N_4722,In_1046,In_686);
and U4723 (N_4723,In_219,In_1952);
or U4724 (N_4724,In_341,In_1471);
nor U4725 (N_4725,In_267,In_1828);
xnor U4726 (N_4726,In_762,In_1055);
and U4727 (N_4727,In_686,In_872);
and U4728 (N_4728,In_480,In_1076);
nand U4729 (N_4729,In_9,In_272);
and U4730 (N_4730,In_1158,In_586);
or U4731 (N_4731,In_1756,In_1121);
nor U4732 (N_4732,In_101,In_427);
and U4733 (N_4733,In_1112,In_89);
or U4734 (N_4734,In_1152,In_1861);
nor U4735 (N_4735,In_1570,In_240);
or U4736 (N_4736,In_1318,In_685);
or U4737 (N_4737,In_530,In_1488);
xnor U4738 (N_4738,In_901,In_21);
and U4739 (N_4739,In_1720,In_590);
and U4740 (N_4740,In_391,In_1481);
nand U4741 (N_4741,In_795,In_152);
nand U4742 (N_4742,In_1496,In_352);
nor U4743 (N_4743,In_923,In_94);
nor U4744 (N_4744,In_1316,In_1200);
nor U4745 (N_4745,In_1616,In_1293);
or U4746 (N_4746,In_1534,In_144);
nand U4747 (N_4747,In_1352,In_499);
and U4748 (N_4748,In_1414,In_1544);
xor U4749 (N_4749,In_1654,In_510);
nand U4750 (N_4750,In_1033,In_396);
nor U4751 (N_4751,In_974,In_133);
and U4752 (N_4752,In_297,In_270);
or U4753 (N_4753,In_944,In_127);
nand U4754 (N_4754,In_1062,In_347);
or U4755 (N_4755,In_1664,In_1933);
and U4756 (N_4756,In_871,In_1435);
and U4757 (N_4757,In_69,In_1956);
and U4758 (N_4758,In_1981,In_1214);
and U4759 (N_4759,In_261,In_715);
and U4760 (N_4760,In_1564,In_1679);
or U4761 (N_4761,In_1394,In_310);
nor U4762 (N_4762,In_298,In_1588);
nor U4763 (N_4763,In_938,In_1581);
xnor U4764 (N_4764,In_1287,In_35);
or U4765 (N_4765,In_179,In_38);
and U4766 (N_4766,In_421,In_1642);
and U4767 (N_4767,In_1181,In_1550);
xor U4768 (N_4768,In_1996,In_1936);
nor U4769 (N_4769,In_444,In_265);
xor U4770 (N_4770,In_713,In_805);
or U4771 (N_4771,In_1139,In_244);
nor U4772 (N_4772,In_1138,In_957);
xnor U4773 (N_4773,In_566,In_1259);
nor U4774 (N_4774,In_685,In_1218);
and U4775 (N_4775,In_1362,In_1380);
nand U4776 (N_4776,In_720,In_1401);
nand U4777 (N_4777,In_325,In_1187);
and U4778 (N_4778,In_651,In_850);
nor U4779 (N_4779,In_1190,In_1318);
nor U4780 (N_4780,In_1901,In_724);
or U4781 (N_4781,In_1492,In_550);
or U4782 (N_4782,In_1875,In_24);
nand U4783 (N_4783,In_561,In_484);
nor U4784 (N_4784,In_872,In_534);
nor U4785 (N_4785,In_1093,In_583);
nor U4786 (N_4786,In_1387,In_588);
or U4787 (N_4787,In_1042,In_573);
or U4788 (N_4788,In_1019,In_1061);
nand U4789 (N_4789,In_1241,In_811);
and U4790 (N_4790,In_1587,In_1605);
and U4791 (N_4791,In_604,In_1691);
nand U4792 (N_4792,In_1816,In_832);
and U4793 (N_4793,In_529,In_1686);
nand U4794 (N_4794,In_924,In_1169);
or U4795 (N_4795,In_264,In_1613);
xor U4796 (N_4796,In_1363,In_1710);
nor U4797 (N_4797,In_1510,In_900);
xnor U4798 (N_4798,In_980,In_463);
nand U4799 (N_4799,In_300,In_446);
nand U4800 (N_4800,In_1289,In_988);
or U4801 (N_4801,In_555,In_1127);
and U4802 (N_4802,In_1374,In_50);
or U4803 (N_4803,In_652,In_1937);
nand U4804 (N_4804,In_1062,In_1810);
nand U4805 (N_4805,In_124,In_1728);
xor U4806 (N_4806,In_1889,In_908);
nor U4807 (N_4807,In_988,In_754);
and U4808 (N_4808,In_1693,In_1062);
nor U4809 (N_4809,In_46,In_137);
nor U4810 (N_4810,In_1490,In_1158);
nand U4811 (N_4811,In_1462,In_183);
or U4812 (N_4812,In_1741,In_216);
xnor U4813 (N_4813,In_600,In_1884);
xnor U4814 (N_4814,In_39,In_1461);
or U4815 (N_4815,In_1135,In_1185);
and U4816 (N_4816,In_1114,In_688);
nor U4817 (N_4817,In_785,In_385);
nor U4818 (N_4818,In_398,In_707);
xnor U4819 (N_4819,In_604,In_1289);
or U4820 (N_4820,In_1036,In_607);
and U4821 (N_4821,In_1489,In_1016);
and U4822 (N_4822,In_370,In_540);
nor U4823 (N_4823,In_1054,In_233);
or U4824 (N_4824,In_1464,In_1989);
or U4825 (N_4825,In_446,In_659);
nor U4826 (N_4826,In_1156,In_485);
nor U4827 (N_4827,In_44,In_1300);
and U4828 (N_4828,In_812,In_229);
xor U4829 (N_4829,In_437,In_587);
nor U4830 (N_4830,In_891,In_1377);
nor U4831 (N_4831,In_438,In_1561);
or U4832 (N_4832,In_1678,In_1818);
or U4833 (N_4833,In_1786,In_1781);
nand U4834 (N_4834,In_1013,In_1736);
nor U4835 (N_4835,In_814,In_414);
nor U4836 (N_4836,In_706,In_17);
nand U4837 (N_4837,In_916,In_1872);
or U4838 (N_4838,In_1810,In_1577);
and U4839 (N_4839,In_1303,In_281);
xnor U4840 (N_4840,In_990,In_941);
or U4841 (N_4841,In_686,In_467);
xnor U4842 (N_4842,In_944,In_1318);
and U4843 (N_4843,In_871,In_599);
or U4844 (N_4844,In_1416,In_565);
or U4845 (N_4845,In_168,In_1068);
nand U4846 (N_4846,In_577,In_646);
and U4847 (N_4847,In_5,In_1322);
or U4848 (N_4848,In_1993,In_402);
nand U4849 (N_4849,In_1975,In_1139);
xnor U4850 (N_4850,In_1570,In_362);
and U4851 (N_4851,In_530,In_1749);
nand U4852 (N_4852,In_847,In_1267);
or U4853 (N_4853,In_1507,In_1762);
xnor U4854 (N_4854,In_1884,In_1082);
xnor U4855 (N_4855,In_181,In_1261);
nor U4856 (N_4856,In_1923,In_611);
xnor U4857 (N_4857,In_17,In_1619);
xor U4858 (N_4858,In_16,In_682);
and U4859 (N_4859,In_91,In_395);
and U4860 (N_4860,In_499,In_1138);
nor U4861 (N_4861,In_1916,In_833);
nor U4862 (N_4862,In_1940,In_1747);
nor U4863 (N_4863,In_1111,In_130);
xnor U4864 (N_4864,In_499,In_1358);
and U4865 (N_4865,In_1838,In_1109);
or U4866 (N_4866,In_959,In_32);
xor U4867 (N_4867,In_599,In_292);
and U4868 (N_4868,In_24,In_1688);
xnor U4869 (N_4869,In_1012,In_1171);
nor U4870 (N_4870,In_710,In_326);
nor U4871 (N_4871,In_1782,In_1372);
nand U4872 (N_4872,In_1672,In_1107);
or U4873 (N_4873,In_1577,In_137);
nand U4874 (N_4874,In_590,In_295);
or U4875 (N_4875,In_1589,In_231);
nor U4876 (N_4876,In_526,In_1614);
or U4877 (N_4877,In_1842,In_1481);
or U4878 (N_4878,In_902,In_1087);
nor U4879 (N_4879,In_920,In_402);
nor U4880 (N_4880,In_849,In_937);
and U4881 (N_4881,In_1972,In_1930);
and U4882 (N_4882,In_1566,In_855);
and U4883 (N_4883,In_1956,In_1040);
nor U4884 (N_4884,In_1994,In_298);
xor U4885 (N_4885,In_977,In_28);
or U4886 (N_4886,In_971,In_1306);
nand U4887 (N_4887,In_1329,In_1341);
nand U4888 (N_4888,In_1817,In_1991);
or U4889 (N_4889,In_74,In_897);
nor U4890 (N_4890,In_1691,In_1812);
nand U4891 (N_4891,In_968,In_373);
xor U4892 (N_4892,In_1523,In_130);
or U4893 (N_4893,In_1481,In_1684);
or U4894 (N_4894,In_1322,In_1091);
nor U4895 (N_4895,In_1262,In_1030);
or U4896 (N_4896,In_1898,In_273);
nor U4897 (N_4897,In_1167,In_691);
and U4898 (N_4898,In_1208,In_1775);
or U4899 (N_4899,In_718,In_1024);
nand U4900 (N_4900,In_706,In_1743);
nor U4901 (N_4901,In_871,In_355);
xor U4902 (N_4902,In_146,In_573);
and U4903 (N_4903,In_1151,In_1833);
nor U4904 (N_4904,In_1175,In_1430);
xnor U4905 (N_4905,In_636,In_647);
xnor U4906 (N_4906,In_523,In_734);
or U4907 (N_4907,In_640,In_582);
nand U4908 (N_4908,In_173,In_938);
xnor U4909 (N_4909,In_1537,In_1695);
nand U4910 (N_4910,In_841,In_807);
nand U4911 (N_4911,In_1266,In_1319);
or U4912 (N_4912,In_1999,In_1486);
nand U4913 (N_4913,In_1392,In_279);
and U4914 (N_4914,In_742,In_343);
and U4915 (N_4915,In_674,In_459);
and U4916 (N_4916,In_1946,In_94);
nand U4917 (N_4917,In_1125,In_510);
nand U4918 (N_4918,In_1991,In_1495);
xor U4919 (N_4919,In_1623,In_1821);
nand U4920 (N_4920,In_243,In_1214);
nand U4921 (N_4921,In_1915,In_1558);
and U4922 (N_4922,In_1857,In_1074);
nand U4923 (N_4923,In_1746,In_736);
and U4924 (N_4924,In_727,In_1057);
and U4925 (N_4925,In_1477,In_1875);
nor U4926 (N_4926,In_1654,In_1129);
nor U4927 (N_4927,In_1573,In_425);
xnor U4928 (N_4928,In_1612,In_38);
xnor U4929 (N_4929,In_1455,In_2);
nand U4930 (N_4930,In_628,In_1614);
and U4931 (N_4931,In_1202,In_723);
nand U4932 (N_4932,In_633,In_1645);
xnor U4933 (N_4933,In_1118,In_857);
or U4934 (N_4934,In_565,In_1025);
nor U4935 (N_4935,In_1301,In_1193);
nor U4936 (N_4936,In_1178,In_745);
nand U4937 (N_4937,In_179,In_801);
and U4938 (N_4938,In_1851,In_558);
and U4939 (N_4939,In_232,In_189);
or U4940 (N_4940,In_1512,In_1386);
or U4941 (N_4941,In_1376,In_627);
nand U4942 (N_4942,In_803,In_317);
and U4943 (N_4943,In_1820,In_1962);
xnor U4944 (N_4944,In_1047,In_610);
nor U4945 (N_4945,In_1247,In_809);
and U4946 (N_4946,In_576,In_1707);
xnor U4947 (N_4947,In_607,In_798);
nand U4948 (N_4948,In_576,In_755);
or U4949 (N_4949,In_1336,In_1384);
nand U4950 (N_4950,In_1746,In_935);
or U4951 (N_4951,In_468,In_226);
nor U4952 (N_4952,In_608,In_175);
xnor U4953 (N_4953,In_399,In_1239);
nand U4954 (N_4954,In_291,In_1207);
and U4955 (N_4955,In_1983,In_1939);
and U4956 (N_4956,In_55,In_1281);
or U4957 (N_4957,In_1151,In_1766);
and U4958 (N_4958,In_736,In_1158);
nor U4959 (N_4959,In_943,In_123);
and U4960 (N_4960,In_332,In_363);
or U4961 (N_4961,In_885,In_1483);
and U4962 (N_4962,In_945,In_1180);
nand U4963 (N_4963,In_968,In_1391);
nand U4964 (N_4964,In_1410,In_198);
nor U4965 (N_4965,In_116,In_1163);
nand U4966 (N_4966,In_1277,In_42);
or U4967 (N_4967,In_1228,In_1062);
and U4968 (N_4968,In_1310,In_1775);
and U4969 (N_4969,In_1591,In_1848);
xor U4970 (N_4970,In_765,In_1039);
and U4971 (N_4971,In_223,In_750);
or U4972 (N_4972,In_978,In_661);
nor U4973 (N_4973,In_1320,In_1964);
or U4974 (N_4974,In_195,In_630);
nor U4975 (N_4975,In_600,In_1090);
nand U4976 (N_4976,In_241,In_95);
nor U4977 (N_4977,In_122,In_344);
nor U4978 (N_4978,In_1830,In_192);
and U4979 (N_4979,In_14,In_1962);
and U4980 (N_4980,In_1622,In_740);
nand U4981 (N_4981,In_1596,In_154);
or U4982 (N_4982,In_622,In_183);
nor U4983 (N_4983,In_516,In_158);
xnor U4984 (N_4984,In_1312,In_668);
nor U4985 (N_4985,In_856,In_884);
or U4986 (N_4986,In_1829,In_702);
xnor U4987 (N_4987,In_1926,In_1987);
nor U4988 (N_4988,In_938,In_870);
nor U4989 (N_4989,In_1464,In_54);
nor U4990 (N_4990,In_1310,In_1334);
nand U4991 (N_4991,In_441,In_1811);
and U4992 (N_4992,In_1344,In_1487);
nor U4993 (N_4993,In_1023,In_765);
xnor U4994 (N_4994,In_1784,In_95);
nand U4995 (N_4995,In_353,In_446);
and U4996 (N_4996,In_1845,In_719);
nand U4997 (N_4997,In_1741,In_868);
nor U4998 (N_4998,In_1175,In_806);
xnor U4999 (N_4999,In_751,In_203);
xor U5000 (N_5000,N_1087,N_520);
nand U5001 (N_5001,N_4947,N_503);
nand U5002 (N_5002,N_1362,N_3510);
nand U5003 (N_5003,N_2450,N_181);
or U5004 (N_5004,N_2164,N_1863);
nand U5005 (N_5005,N_3082,N_4586);
nor U5006 (N_5006,N_235,N_187);
and U5007 (N_5007,N_204,N_366);
and U5008 (N_5008,N_4897,N_3518);
xor U5009 (N_5009,N_2386,N_1343);
and U5010 (N_5010,N_4913,N_1556);
nand U5011 (N_5011,N_1305,N_494);
xnor U5012 (N_5012,N_2491,N_2374);
and U5013 (N_5013,N_4290,N_3059);
and U5014 (N_5014,N_2738,N_1553);
and U5015 (N_5015,N_357,N_4090);
nor U5016 (N_5016,N_3598,N_1478);
nor U5017 (N_5017,N_1283,N_2588);
or U5018 (N_5018,N_1552,N_226);
or U5019 (N_5019,N_1729,N_4860);
nand U5020 (N_5020,N_3571,N_3079);
or U5021 (N_5021,N_895,N_837);
nand U5022 (N_5022,N_3291,N_564);
xor U5023 (N_5023,N_4332,N_2595);
nand U5024 (N_5024,N_3227,N_1319);
and U5025 (N_5025,N_1223,N_1370);
and U5026 (N_5026,N_1050,N_3270);
or U5027 (N_5027,N_4142,N_4401);
nand U5028 (N_5028,N_3791,N_3566);
xnor U5029 (N_5029,N_2831,N_3494);
nand U5030 (N_5030,N_97,N_1213);
nand U5031 (N_5031,N_2140,N_4354);
or U5032 (N_5032,N_4920,N_1616);
or U5033 (N_5033,N_3938,N_3233);
nor U5034 (N_5034,N_4210,N_3253);
nand U5035 (N_5035,N_1228,N_3524);
xnor U5036 (N_5036,N_2189,N_1134);
nand U5037 (N_5037,N_2949,N_3184);
or U5038 (N_5038,N_2070,N_2004);
nand U5039 (N_5039,N_2321,N_4239);
and U5040 (N_5040,N_3287,N_935);
xor U5041 (N_5041,N_651,N_2313);
nor U5042 (N_5042,N_931,N_1458);
and U5043 (N_5043,N_756,N_2965);
xnor U5044 (N_5044,N_1809,N_495);
nand U5045 (N_5045,N_2151,N_3765);
or U5046 (N_5046,N_166,N_439);
nor U5047 (N_5047,N_1926,N_4640);
xor U5048 (N_5048,N_3289,N_3353);
or U5049 (N_5049,N_4956,N_1379);
nand U5050 (N_5050,N_3318,N_472);
xor U5051 (N_5051,N_1566,N_1197);
or U5052 (N_5052,N_2184,N_269);
nor U5053 (N_5053,N_2011,N_4540);
nor U5054 (N_5054,N_227,N_2293);
nor U5055 (N_5055,N_3495,N_3280);
xnor U5056 (N_5056,N_4594,N_1234);
nand U5057 (N_5057,N_1650,N_4682);
xor U5058 (N_5058,N_2631,N_1535);
and U5059 (N_5059,N_3626,N_2224);
nor U5060 (N_5060,N_1452,N_2360);
and U5061 (N_5061,N_3503,N_2812);
or U5062 (N_5062,N_448,N_3385);
nand U5063 (N_5063,N_459,N_553);
and U5064 (N_5064,N_4637,N_1732);
and U5065 (N_5065,N_3007,N_3700);
nand U5066 (N_5066,N_1963,N_201);
xor U5067 (N_5067,N_157,N_1514);
xor U5068 (N_5068,N_2780,N_876);
or U5069 (N_5069,N_0,N_4365);
nand U5070 (N_5070,N_2461,N_3941);
nor U5071 (N_5071,N_4843,N_3367);
and U5072 (N_5072,N_4716,N_4882);
nor U5073 (N_5073,N_2594,N_4267);
xnor U5074 (N_5074,N_4978,N_2923);
nor U5075 (N_5075,N_4722,N_4954);
and U5076 (N_5076,N_513,N_1992);
or U5077 (N_5077,N_1090,N_1911);
and U5078 (N_5078,N_991,N_2798);
nor U5079 (N_5079,N_555,N_4160);
nand U5080 (N_5080,N_2128,N_4538);
nor U5081 (N_5081,N_875,N_1310);
nor U5082 (N_5082,N_2410,N_754);
nor U5083 (N_5083,N_2706,N_2833);
or U5084 (N_5084,N_2768,N_2983);
and U5085 (N_5085,N_289,N_3914);
xnor U5086 (N_5086,N_2922,N_2481);
nand U5087 (N_5087,N_2921,N_2357);
or U5088 (N_5088,N_2159,N_3905);
or U5089 (N_5089,N_3612,N_1568);
nor U5090 (N_5090,N_854,N_3131);
and U5091 (N_5091,N_276,N_690);
nand U5092 (N_5092,N_2396,N_4970);
and U5093 (N_5093,N_4434,N_947);
nand U5094 (N_5094,N_285,N_4742);
xnor U5095 (N_5095,N_208,N_3274);
and U5096 (N_5096,N_3067,N_2085);
and U5097 (N_5097,N_163,N_3559);
and U5098 (N_5098,N_3927,N_4576);
nand U5099 (N_5099,N_2757,N_2333);
nand U5100 (N_5100,N_4685,N_4271);
and U5101 (N_5101,N_3561,N_627);
or U5102 (N_5102,N_4322,N_3207);
nand U5103 (N_5103,N_1372,N_2094);
xnor U5104 (N_5104,N_1152,N_3530);
nand U5105 (N_5105,N_2205,N_3871);
or U5106 (N_5106,N_4299,N_2528);
xnor U5107 (N_5107,N_4135,N_4318);
or U5108 (N_5108,N_440,N_1254);
nor U5109 (N_5109,N_4754,N_147);
xnor U5110 (N_5110,N_698,N_1089);
nor U5111 (N_5111,N_2551,N_2846);
or U5112 (N_5112,N_3256,N_2659);
and U5113 (N_5113,N_1112,N_1107);
or U5114 (N_5114,N_3642,N_504);
xnor U5115 (N_5115,N_3349,N_4406);
and U5116 (N_5116,N_863,N_2581);
or U5117 (N_5117,N_1690,N_22);
xnor U5118 (N_5118,N_3666,N_1576);
and U5119 (N_5119,N_4720,N_582);
nor U5120 (N_5120,N_1925,N_1292);
and U5121 (N_5121,N_524,N_1313);
or U5122 (N_5122,N_3712,N_2653);
or U5123 (N_5123,N_4861,N_2955);
and U5124 (N_5124,N_4687,N_1339);
xnor U5125 (N_5125,N_2220,N_3752);
xor U5126 (N_5126,N_2329,N_1888);
nor U5127 (N_5127,N_1561,N_2580);
or U5128 (N_5128,N_4775,N_4427);
nand U5129 (N_5129,N_2380,N_3931);
and U5130 (N_5130,N_3934,N_2275);
nor U5131 (N_5131,N_3847,N_675);
or U5132 (N_5132,N_3872,N_2815);
nor U5133 (N_5133,N_156,N_842);
nand U5134 (N_5134,N_343,N_4283);
or U5135 (N_5135,N_3687,N_4200);
or U5136 (N_5136,N_447,N_3877);
nor U5137 (N_5137,N_3010,N_2123);
or U5138 (N_5138,N_4512,N_3188);
xnor U5139 (N_5139,N_3133,N_2839);
xor U5140 (N_5140,N_2473,N_4292);
or U5141 (N_5141,N_919,N_4460);
xor U5142 (N_5142,N_4565,N_1233);
nand U5143 (N_5143,N_491,N_430);
or U5144 (N_5144,N_333,N_4987);
and U5145 (N_5145,N_261,N_4389);
and U5146 (N_5146,N_3865,N_244);
nand U5147 (N_5147,N_2935,N_2507);
nand U5148 (N_5148,N_3462,N_3108);
nand U5149 (N_5149,N_1814,N_4645);
xor U5150 (N_5150,N_402,N_4407);
nand U5151 (N_5151,N_1894,N_4070);
or U5152 (N_5152,N_838,N_3011);
nand U5153 (N_5153,N_2435,N_2578);
or U5154 (N_5154,N_1147,N_1676);
xor U5155 (N_5155,N_1536,N_4238);
and U5156 (N_5156,N_714,N_2861);
and U5157 (N_5157,N_3311,N_1666);
xnor U5158 (N_5158,N_4827,N_3266);
nand U5159 (N_5159,N_396,N_3595);
or U5160 (N_5160,N_3102,N_660);
nand U5161 (N_5161,N_3220,N_893);
and U5162 (N_5162,N_580,N_2060);
nor U5163 (N_5163,N_1591,N_1889);
nand U5164 (N_5164,N_4976,N_3599);
or U5165 (N_5165,N_464,N_936);
xnor U5166 (N_5166,N_2139,N_4990);
nand U5167 (N_5167,N_3812,N_358);
and U5168 (N_5168,N_3107,N_1918);
nor U5169 (N_5169,N_2945,N_1739);
xnor U5170 (N_5170,N_2550,N_3751);
nor U5171 (N_5171,N_260,N_2233);
xor U5172 (N_5172,N_3878,N_2840);
xnor U5173 (N_5173,N_1121,N_844);
nand U5174 (N_5174,N_4361,N_3917);
xnor U5175 (N_5175,N_2206,N_4744);
and U5176 (N_5176,N_1180,N_2740);
xnor U5177 (N_5177,N_2250,N_2288);
and U5178 (N_5178,N_571,N_1772);
nor U5179 (N_5179,N_4713,N_2804);
nor U5180 (N_5180,N_2197,N_197);
and U5181 (N_5181,N_903,N_1707);
and U5182 (N_5182,N_4963,N_2195);
or U5183 (N_5183,N_2315,N_1126);
nand U5184 (N_5184,N_1852,N_3630);
nand U5185 (N_5185,N_4485,N_3424);
xor U5186 (N_5186,N_836,N_275);
and U5187 (N_5187,N_3838,N_3166);
xnor U5188 (N_5188,N_173,N_4062);
or U5189 (N_5189,N_231,N_2673);
and U5190 (N_5190,N_508,N_2456);
nand U5191 (N_5191,N_3602,N_1430);
nand U5192 (N_5192,N_2514,N_2548);
xnor U5193 (N_5193,N_3068,N_2889);
nor U5194 (N_5194,N_310,N_2806);
nor U5195 (N_5195,N_199,N_3532);
xnor U5196 (N_5196,N_605,N_3628);
or U5197 (N_5197,N_336,N_4693);
and U5198 (N_5198,N_4523,N_24);
nand U5199 (N_5199,N_4045,N_4579);
and U5200 (N_5200,N_3758,N_3379);
and U5201 (N_5201,N_1462,N_3641);
or U5202 (N_5202,N_2379,N_1636);
nand U5203 (N_5203,N_3577,N_4648);
nor U5204 (N_5204,N_4680,N_770);
xor U5205 (N_5205,N_3043,N_1076);
xor U5206 (N_5206,N_2193,N_1193);
or U5207 (N_5207,N_2444,N_3484);
and U5208 (N_5208,N_1906,N_2970);
xnor U5209 (N_5209,N_1848,N_2503);
or U5210 (N_5210,N_4139,N_4181);
xor U5211 (N_5211,N_758,N_4317);
or U5212 (N_5212,N_2733,N_3189);
xnor U5213 (N_5213,N_1723,N_15);
and U5214 (N_5214,N_708,N_4047);
nand U5215 (N_5215,N_2084,N_2200);
xor U5216 (N_5216,N_3552,N_843);
or U5217 (N_5217,N_3918,N_2340);
nand U5218 (N_5218,N_1450,N_3924);
or U5219 (N_5219,N_1981,N_4337);
nand U5220 (N_5220,N_1725,N_1455);
nand U5221 (N_5221,N_4166,N_3675);
nor U5222 (N_5222,N_663,N_3065);
or U5223 (N_5223,N_1189,N_4457);
xor U5224 (N_5224,N_2388,N_2196);
and U5225 (N_5225,N_2873,N_3903);
xnor U5226 (N_5226,N_4125,N_2743);
or U5227 (N_5227,N_450,N_3395);
or U5228 (N_5228,N_3716,N_4691);
and U5229 (N_5229,N_1151,N_2901);
nand U5230 (N_5230,N_1727,N_2287);
nor U5231 (N_5231,N_534,N_799);
nand U5232 (N_5232,N_2353,N_145);
nor U5233 (N_5233,N_4076,N_4399);
or U5234 (N_5234,N_1329,N_924);
nor U5235 (N_5235,N_2549,N_1106);
nand U5236 (N_5236,N_1761,N_2492);
nor U5237 (N_5237,N_855,N_4205);
xnor U5238 (N_5238,N_2681,N_469);
nand U5239 (N_5239,N_2942,N_1869);
nand U5240 (N_5240,N_4898,N_2585);
or U5241 (N_5241,N_1923,N_1186);
and U5242 (N_5242,N_3048,N_3117);
and U5243 (N_5243,N_3348,N_3155);
nand U5244 (N_5244,N_409,N_943);
or U5245 (N_5245,N_1860,N_397);
or U5246 (N_5246,N_3608,N_2991);
nor U5247 (N_5247,N_415,N_2056);
xor U5248 (N_5248,N_878,N_3899);
and U5249 (N_5249,N_4279,N_3778);
nor U5250 (N_5250,N_4146,N_3025);
and U5251 (N_5251,N_1083,N_4018);
xnor U5252 (N_5252,N_2782,N_2536);
or U5253 (N_5253,N_2712,N_891);
and U5254 (N_5254,N_4721,N_1807);
nor U5255 (N_5255,N_1079,N_589);
nand U5256 (N_5256,N_1038,N_3913);
and U5257 (N_5257,N_3140,N_590);
and U5258 (N_5258,N_3841,N_602);
and U5259 (N_5259,N_1491,N_108);
or U5260 (N_5260,N_725,N_3964);
or U5261 (N_5261,N_2041,N_3928);
and U5262 (N_5262,N_1903,N_1104);
nand U5263 (N_5263,N_3590,N_1510);
and U5264 (N_5264,N_203,N_1742);
or U5265 (N_5265,N_545,N_2553);
nand U5266 (N_5266,N_1977,N_4305);
or U5267 (N_5267,N_3717,N_4081);
nand U5268 (N_5268,N_2166,N_598);
xor U5269 (N_5269,N_3638,N_576);
nor U5270 (N_5270,N_386,N_1784);
nor U5271 (N_5271,N_870,N_1476);
nor U5272 (N_5272,N_64,N_2941);
or U5273 (N_5273,N_1039,N_2677);
and U5274 (N_5274,N_3968,N_1013);
nand U5275 (N_5275,N_3257,N_2530);
or U5276 (N_5276,N_1482,N_4785);
xnor U5277 (N_5277,N_1779,N_1944);
xor U5278 (N_5278,N_3498,N_248);
and U5279 (N_5279,N_4169,N_2939);
nor U5280 (N_5280,N_4592,N_3830);
and U5281 (N_5281,N_2446,N_2217);
or U5282 (N_5282,N_2411,N_1530);
nor U5283 (N_5283,N_3673,N_819);
nand U5284 (N_5284,N_1543,N_4184);
and U5285 (N_5285,N_1181,N_1564);
and U5286 (N_5286,N_2218,N_793);
xnor U5287 (N_5287,N_1970,N_2517);
nand U5288 (N_5288,N_523,N_320);
nand U5289 (N_5289,N_3769,N_2073);
xnor U5290 (N_5290,N_4593,N_4063);
and U5291 (N_5291,N_3859,N_3784);
nor U5292 (N_5292,N_4084,N_2149);
nand U5293 (N_5293,N_3091,N_4451);
or U5294 (N_5294,N_4935,N_4327);
nor U5295 (N_5295,N_2537,N_4331);
or U5296 (N_5296,N_300,N_4017);
nor U5297 (N_5297,N_2480,N_255);
or U5298 (N_5298,N_1939,N_1961);
xor U5299 (N_5299,N_992,N_2709);
nor U5300 (N_5300,N_2323,N_2883);
nand U5301 (N_5301,N_2558,N_3464);
nand U5302 (N_5302,N_76,N_2442);
xor U5303 (N_5303,N_2539,N_1494);
nand U5304 (N_5304,N_1984,N_4188);
and U5305 (N_5305,N_3795,N_4826);
nor U5306 (N_5306,N_2124,N_4649);
xnor U5307 (N_5307,N_2427,N_597);
nand U5308 (N_5308,N_3659,N_3900);
nand U5309 (N_5309,N_982,N_2547);
and U5310 (N_5310,N_2478,N_420);
nand U5311 (N_5311,N_1615,N_3226);
xor U5312 (N_5312,N_3975,N_840);
or U5313 (N_5313,N_4581,N_4929);
and U5314 (N_5314,N_60,N_4470);
or U5315 (N_5315,N_1808,N_3083);
nand U5316 (N_5316,N_2613,N_2393);
nor U5317 (N_5317,N_2805,N_1851);
nand U5318 (N_5318,N_1055,N_2968);
nand U5319 (N_5319,N_4053,N_3430);
nor U5320 (N_5320,N_2061,N_2752);
or U5321 (N_5321,N_4270,N_1133);
nand U5322 (N_5322,N_2420,N_127);
or U5323 (N_5323,N_4250,N_405);
nor U5324 (N_5324,N_1855,N_1644);
nand U5325 (N_5325,N_1098,N_3465);
xor U5326 (N_5326,N_1737,N_1628);
and U5327 (N_5327,N_3062,N_3493);
nand U5328 (N_5328,N_2108,N_1278);
xor U5329 (N_5329,N_2776,N_3990);
and U5330 (N_5330,N_591,N_1559);
and U5331 (N_5331,N_2796,N_1651);
or U5332 (N_5332,N_3665,N_2207);
nand U5333 (N_5333,N_4962,N_3589);
or U5334 (N_5334,N_2531,N_3668);
and U5335 (N_5335,N_4993,N_2009);
xnor U5336 (N_5336,N_1453,N_2399);
nor U5337 (N_5337,N_3036,N_2314);
and U5338 (N_5338,N_480,N_507);
xnor U5339 (N_5339,N_7,N_2020);
and U5340 (N_5340,N_3962,N_850);
and U5341 (N_5341,N_4625,N_1298);
or U5342 (N_5342,N_3639,N_406);
nor U5343 (N_5343,N_4817,N_1082);
xnor U5344 (N_5344,N_2756,N_1877);
and U5345 (N_5345,N_2038,N_1901);
nor U5346 (N_5346,N_3325,N_1592);
or U5347 (N_5347,N_1804,N_2552);
xnor U5348 (N_5348,N_1957,N_2135);
and U5349 (N_5349,N_2244,N_162);
nand U5350 (N_5350,N_4289,N_874);
nand U5351 (N_5351,N_3960,N_4025);
xor U5352 (N_5352,N_3926,N_4934);
or U5353 (N_5353,N_1694,N_4120);
xnor U5354 (N_5354,N_4425,N_2182);
nor U5355 (N_5355,N_1032,N_2979);
or U5356 (N_5356,N_2685,N_3790);
and U5357 (N_5357,N_592,N_777);
or U5358 (N_5358,N_311,N_69);
nand U5359 (N_5359,N_3759,N_1070);
and U5360 (N_5360,N_4002,N_3413);
nand U5361 (N_5361,N_4464,N_2557);
and U5362 (N_5362,N_404,N_3525);
and U5363 (N_5363,N_3643,N_138);
nor U5364 (N_5364,N_609,N_4644);
nor U5365 (N_5365,N_210,N_3709);
nor U5366 (N_5366,N_1678,N_3168);
nor U5367 (N_5367,N_3569,N_4975);
nand U5368 (N_5368,N_4772,N_3662);
nor U5369 (N_5369,N_4830,N_1008);
and U5370 (N_5370,N_1847,N_718);
xor U5371 (N_5371,N_1780,N_4122);
and U5372 (N_5372,N_2302,N_1002);
xor U5373 (N_5373,N_23,N_1640);
nor U5374 (N_5374,N_556,N_2919);
nor U5375 (N_5375,N_729,N_3652);
xnor U5376 (N_5376,N_1115,N_4859);
xnor U5377 (N_5377,N_1352,N_3112);
nor U5378 (N_5378,N_677,N_1012);
and U5379 (N_5379,N_955,N_3714);
and U5380 (N_5380,N_3815,N_786);
and U5381 (N_5381,N_4613,N_3301);
nand U5382 (N_5382,N_4751,N_3647);
nand U5383 (N_5383,N_2817,N_4651);
or U5384 (N_5384,N_2748,N_4621);
and U5385 (N_5385,N_4953,N_4659);
nand U5386 (N_5386,N_2285,N_4177);
nand U5387 (N_5387,N_379,N_2168);
nand U5388 (N_5388,N_636,N_4253);
or U5389 (N_5389,N_196,N_4266);
xor U5390 (N_5390,N_1364,N_1388);
or U5391 (N_5391,N_4450,N_533);
xor U5392 (N_5392,N_4842,N_2728);
nand U5393 (N_5393,N_2746,N_3582);
nand U5394 (N_5394,N_1417,N_4156);
xor U5395 (N_5395,N_4027,N_4286);
and U5396 (N_5396,N_2764,N_4884);
xor U5397 (N_5397,N_1569,N_2064);
or U5398 (N_5398,N_3425,N_1881);
nor U5399 (N_5399,N_1786,N_780);
or U5400 (N_5400,N_1331,N_3583);
and U5401 (N_5401,N_1327,N_1353);
nor U5402 (N_5402,N_1975,N_4941);
and U5403 (N_5403,N_4012,N_3515);
xor U5404 (N_5404,N_3943,N_4663);
or U5405 (N_5405,N_3617,N_215);
xnor U5406 (N_5406,N_2346,N_4487);
or U5407 (N_5407,N_3298,N_2008);
and U5408 (N_5408,N_3012,N_3435);
xor U5409 (N_5409,N_3978,N_2649);
nor U5410 (N_5410,N_2515,N_2930);
or U5411 (N_5411,N_65,N_2663);
and U5412 (N_5412,N_3111,N_3743);
and U5413 (N_5413,N_364,N_4875);
nor U5414 (N_5414,N_263,N_4308);
nor U5415 (N_5415,N_3149,N_3760);
nor U5416 (N_5416,N_1398,N_2384);
nand U5417 (N_5417,N_1525,N_3050);
nor U5418 (N_5418,N_3998,N_1326);
xor U5419 (N_5419,N_4341,N_798);
xor U5420 (N_5420,N_1401,N_1465);
or U5421 (N_5421,N_2660,N_4569);
xnor U5422 (N_5422,N_1935,N_1685);
or U5423 (N_5423,N_2633,N_411);
and U5424 (N_5424,N_2433,N_3340);
and U5425 (N_5425,N_179,N_3753);
xor U5426 (N_5426,N_3267,N_962);
or U5427 (N_5427,N_2079,N_1574);
nor U5428 (N_5428,N_1657,N_2429);
nand U5429 (N_5429,N_692,N_3119);
and U5430 (N_5430,N_2511,N_1230);
xnor U5431 (N_5431,N_2457,N_3061);
nand U5432 (N_5432,N_899,N_3027);
nand U5433 (N_5433,N_3969,N_1674);
nor U5434 (N_5434,N_3183,N_4165);
nor U5435 (N_5435,N_3084,N_542);
and U5436 (N_5436,N_4521,N_4151);
nor U5437 (N_5437,N_435,N_4840);
nand U5438 (N_5438,N_2255,N_87);
xor U5439 (N_5439,N_463,N_1281);
nand U5440 (N_5440,N_2499,N_4071);
nor U5441 (N_5441,N_4473,N_1743);
xor U5442 (N_5442,N_1639,N_647);
or U5443 (N_5443,N_730,N_2697);
nand U5444 (N_5444,N_1195,N_1160);
nand U5445 (N_5445,N_154,N_2306);
xor U5446 (N_5446,N_3203,N_2987);
xnor U5447 (N_5447,N_2679,N_2607);
nor U5448 (N_5448,N_1065,N_573);
nor U5449 (N_5449,N_2417,N_3200);
or U5450 (N_5450,N_3688,N_4757);
xor U5451 (N_5451,N_1257,N_4522);
and U5452 (N_5452,N_3755,N_1787);
and U5453 (N_5453,N_2785,N_679);
xnor U5454 (N_5454,N_1066,N_350);
nand U5455 (N_5455,N_334,N_1423);
and U5456 (N_5456,N_4553,N_1167);
and U5457 (N_5457,N_3970,N_1893);
or U5458 (N_5458,N_3676,N_1258);
nor U5459 (N_5459,N_1222,N_1184);
and U5460 (N_5460,N_86,N_2148);
xnor U5461 (N_5461,N_2230,N_237);
xor U5462 (N_5462,N_2973,N_4703);
and U5463 (N_5463,N_81,N_3777);
xnor U5464 (N_5464,N_1471,N_916);
or U5465 (N_5465,N_2467,N_2522);
nand U5466 (N_5466,N_1294,N_2645);
xor U5467 (N_5467,N_1041,N_3953);
nand U5468 (N_5468,N_1857,N_3002);
nand U5469 (N_5469,N_4708,N_4541);
nand U5470 (N_5470,N_4458,N_2146);
nor U5471 (N_5471,N_3281,N_1256);
xor U5472 (N_5472,N_4356,N_313);
xor U5473 (N_5473,N_1500,N_4482);
nor U5474 (N_5474,N_1501,N_2811);
xor U5475 (N_5475,N_4971,N_3077);
xor U5476 (N_5476,N_3146,N_252);
and U5477 (N_5477,N_4433,N_2342);
and U5478 (N_5478,N_2715,N_1998);
xor U5479 (N_5479,N_2228,N_641);
or U5480 (N_5480,N_652,N_862);
or U5481 (N_5481,N_4995,N_3763);
nand U5482 (N_5482,N_3141,N_2801);
xor U5483 (N_5483,N_4611,N_2489);
nor U5484 (N_5484,N_266,N_98);
xnor U5485 (N_5485,N_775,N_2927);
and U5486 (N_5486,N_3368,N_3883);
or U5487 (N_5487,N_4723,N_387);
nor U5488 (N_5488,N_1048,N_2894);
xor U5489 (N_5489,N_4204,N_1266);
xnor U5490 (N_5490,N_4686,N_281);
nor U5491 (N_5491,N_2176,N_1381);
xor U5492 (N_5492,N_858,N_4259);
xnor U5493 (N_5493,N_3159,N_678);
nand U5494 (N_5494,N_1156,N_2251);
nand U5495 (N_5495,N_2412,N_4622);
or U5496 (N_5496,N_4101,N_1360);
or U5497 (N_5497,N_4710,N_2072);
nor U5498 (N_5498,N_381,N_3995);
xnor U5499 (N_5499,N_2283,N_3819);
and U5500 (N_5500,N_3750,N_1908);
nor U5501 (N_5501,N_1753,N_3147);
xnor U5502 (N_5502,N_417,N_4903);
nand U5503 (N_5503,N_1336,N_4009);
or U5504 (N_5504,N_2376,N_1795);
and U5505 (N_5505,N_1007,N_4961);
nand U5506 (N_5506,N_3210,N_3591);
or U5507 (N_5507,N_2236,N_2995);
xor U5508 (N_5508,N_1764,N_4787);
xor U5509 (N_5509,N_517,N_3129);
xnor U5510 (N_5510,N_2111,N_2837);
nand U5511 (N_5511,N_42,N_1366);
xor U5512 (N_5512,N_929,N_2373);
xor U5513 (N_5513,N_1240,N_3981);
xor U5514 (N_5514,N_2870,N_1031);
nor U5515 (N_5515,N_222,N_4150);
nor U5516 (N_5516,N_1858,N_3263);
or U5517 (N_5517,N_912,N_2001);
and U5518 (N_5518,N_3442,N_314);
nand U5519 (N_5519,N_3805,N_4642);
nor U5520 (N_5520,N_2828,N_2154);
xor U5521 (N_5521,N_806,N_1188);
or U5522 (N_5522,N_67,N_4832);
nor U5523 (N_5523,N_3772,N_2065);
nor U5524 (N_5524,N_2934,N_3240);
nand U5525 (N_5525,N_2221,N_3771);
xor U5526 (N_5526,N_1297,N_4542);
nor U5527 (N_5527,N_1788,N_1390);
and U5528 (N_5528,N_2929,N_1363);
and U5529 (N_5529,N_4983,N_11);
xor U5530 (N_5530,N_319,N_1709);
or U5531 (N_5531,N_242,N_2896);
nand U5532 (N_5532,N_2322,N_1157);
nand U5533 (N_5533,N_1198,N_458);
xnor U5534 (N_5534,N_4255,N_3034);
xor U5535 (N_5535,N_4379,N_4351);
nor U5536 (N_5536,N_3891,N_3126);
nor U5537 (N_5537,N_3640,N_431);
or U5538 (N_5538,N_374,N_4706);
or U5539 (N_5539,N_2643,N_1068);
and U5540 (N_5540,N_3669,N_4702);
and U5541 (N_5541,N_4319,N_2269);
nand U5542 (N_5542,N_3324,N_4635);
or U5543 (N_5543,N_72,N_1194);
nor U5544 (N_5544,N_851,N_483);
and U5545 (N_5545,N_1598,N_3259);
nand U5546 (N_5546,N_4666,N_3575);
nor U5547 (N_5547,N_905,N_1077);
xor U5548 (N_5548,N_2783,N_809);
xnor U5549 (N_5549,N_4841,N_2017);
xnor U5550 (N_5550,N_4097,N_4363);
or U5551 (N_5551,N_4634,N_3912);
and U5552 (N_5552,N_1611,N_2847);
nor U5553 (N_5553,N_3078,N_824);
and U5554 (N_5554,N_3033,N_141);
nor U5555 (N_5555,N_2795,N_1744);
or U5556 (N_5556,N_993,N_3362);
and U5557 (N_5557,N_3094,N_805);
xnor U5558 (N_5558,N_152,N_3152);
nand U5559 (N_5559,N_4164,N_2647);
nor U5560 (N_5560,N_613,N_1477);
xnor U5561 (N_5561,N_1922,N_1021);
xnor U5562 (N_5562,N_2526,N_4065);
or U5563 (N_5563,N_4874,N_2284);
or U5564 (N_5564,N_327,N_1322);
xnor U5565 (N_5565,N_3670,N_1614);
xnor U5566 (N_5566,N_372,N_3729);
nor U5567 (N_5567,N_3528,N_2591);
nor U5568 (N_5568,N_441,N_3966);
nor U5569 (N_5569,N_1128,N_768);
or U5570 (N_5570,N_2246,N_236);
or U5571 (N_5571,N_1443,N_853);
and U5572 (N_5572,N_3619,N_3764);
nand U5573 (N_5573,N_1016,N_1308);
nor U5574 (N_5574,N_4763,N_4272);
and U5575 (N_5575,N_772,N_1789);
xnor U5576 (N_5576,N_4753,N_2249);
xnor U5577 (N_5577,N_2210,N_2114);
and U5578 (N_5578,N_1108,N_3021);
nor U5579 (N_5579,N_2996,N_2152);
xor U5580 (N_5580,N_4631,N_129);
and U5581 (N_5581,N_890,N_1006);
and U5582 (N_5582,N_3625,N_2863);
nor U5583 (N_5583,N_3046,N_4739);
and U5584 (N_5584,N_332,N_3864);
nor U5585 (N_5585,N_2848,N_630);
or U5586 (N_5586,N_2270,N_3313);
xnor U5587 (N_5587,N_622,N_1005);
nand U5588 (N_5588,N_4917,N_634);
nand U5589 (N_5589,N_1053,N_1612);
and U5590 (N_5590,N_2238,N_645);
nor U5591 (N_5591,N_1051,N_849);
and U5592 (N_5592,N_839,N_4506);
and U5593 (N_5593,N_4886,N_831);
xnor U5594 (N_5594,N_28,N_161);
nand U5595 (N_5595,N_2147,N_2695);
or U5596 (N_5596,N_394,N_3610);
and U5597 (N_5597,N_1052,N_3315);
or U5598 (N_5598,N_1120,N_4802);
or U5599 (N_5599,N_3370,N_3333);
or U5600 (N_5600,N_1527,N_2505);
nand U5601 (N_5601,N_1365,N_1192);
or U5602 (N_5602,N_3861,N_2183);
or U5603 (N_5603,N_2120,N_3955);
nand U5604 (N_5604,N_3215,N_1432);
nand U5605 (N_5605,N_4342,N_3715);
xor U5606 (N_5606,N_2907,N_1127);
xor U5607 (N_5607,N_3344,N_1839);
and U5608 (N_5608,N_3605,N_618);
and U5609 (N_5609,N_4823,N_3609);
xor U5610 (N_5610,N_2802,N_4430);
nor U5611 (N_5611,N_1659,N_2532);
nand U5612 (N_5612,N_4246,N_885);
and U5613 (N_5613,N_776,N_1361);
xor U5614 (N_5614,N_3519,N_2316);
xnor U5615 (N_5615,N_2933,N_2854);
nor U5616 (N_5616,N_3099,N_1868);
xnor U5617 (N_5617,N_3169,N_3833);
and U5618 (N_5618,N_2024,N_2104);
nor U5619 (N_5619,N_4157,N_4347);
nor U5620 (N_5620,N_2932,N_511);
nand U5621 (N_5621,N_4452,N_4877);
nand U5622 (N_5622,N_4050,N_2771);
and U5623 (N_5623,N_1951,N_693);
xnor U5624 (N_5624,N_2243,N_2068);
and U5625 (N_5625,N_3150,N_1660);
xor U5626 (N_5626,N_3658,N_4497);
nor U5627 (N_5627,N_4026,N_4310);
or U5628 (N_5628,N_2402,N_1806);
nor U5629 (N_5629,N_360,N_4872);
or U5630 (N_5630,N_14,N_4815);
nand U5631 (N_5631,N_4623,N_4468);
xnor U5632 (N_5632,N_980,N_585);
nand U5633 (N_5633,N_2686,N_1778);
xnor U5634 (N_5634,N_2666,N_1677);
or U5635 (N_5635,N_4519,N_2431);
or U5636 (N_5636,N_1320,N_2000);
nor U5637 (N_5637,N_51,N_412);
or U5638 (N_5638,N_3,N_2957);
nand U5639 (N_5639,N_3661,N_3466);
nand U5640 (N_5640,N_1447,N_4924);
and U5641 (N_5641,N_4226,N_2610);
nand U5642 (N_5642,N_1647,N_2775);
nor U5643 (N_5643,N_2787,N_1509);
nor U5644 (N_5644,N_950,N_3517);
or U5645 (N_5645,N_4459,N_4366);
nor U5646 (N_5646,N_234,N_3456);
xnor U5647 (N_5647,N_543,N_2301);
nand U5648 (N_5648,N_134,N_2562);
or U5649 (N_5649,N_3680,N_1905);
xnor U5650 (N_5650,N_3798,N_1837);
or U5651 (N_5651,N_4677,N_1745);
or U5652 (N_5652,N_1846,N_1526);
or U5653 (N_5653,N_3038,N_4424);
and U5654 (N_5654,N_3109,N_1267);
nand U5655 (N_5655,N_4449,N_2330);
nand U5656 (N_5656,N_981,N_1956);
and U5657 (N_5657,N_3134,N_642);
xor U5658 (N_5658,N_4853,N_4306);
xnor U5659 (N_5659,N_4902,N_2116);
xor U5660 (N_5660,N_2022,N_723);
and U5661 (N_5661,N_1554,N_3303);
xnor U5662 (N_5662,N_2824,N_2403);
or U5663 (N_5663,N_697,N_1796);
nor U5664 (N_5664,N_2328,N_3306);
xnor U5665 (N_5665,N_525,N_1733);
nand U5666 (N_5666,N_3418,N_4825);
or U5667 (N_5667,N_673,N_682);
or U5668 (N_5668,N_262,N_2192);
nor U5669 (N_5669,N_4215,N_1248);
nor U5670 (N_5670,N_4489,N_2289);
nand U5671 (N_5671,N_4894,N_710);
nand U5672 (N_5672,N_3984,N_2361);
nand U5673 (N_5673,N_3706,N_3317);
nor U5674 (N_5674,N_3410,N_481);
nor U5675 (N_5675,N_4483,N_4086);
or U5676 (N_5676,N_3522,N_497);
or U5677 (N_5677,N_4106,N_3218);
nor U5678 (N_5678,N_3735,N_873);
nor U5679 (N_5679,N_1886,N_2136);
nor U5680 (N_5680,N_1580,N_3983);
and U5681 (N_5681,N_4137,N_8);
xor U5682 (N_5682,N_735,N_745);
xor U5683 (N_5683,N_351,N_325);
nand U5684 (N_5684,N_2982,N_1004);
or U5685 (N_5685,N_2618,N_1930);
and U5686 (N_5686,N_3906,N_4111);
nor U5687 (N_5687,N_2033,N_2239);
and U5688 (N_5688,N_4382,N_1890);
or U5689 (N_5689,N_1272,N_4790);
nor U5690 (N_5690,N_1289,N_4245);
and U5691 (N_5691,N_4024,N_1867);
nor U5692 (N_5692,N_661,N_3307);
nand U5693 (N_5693,N_4221,N_140);
and U5694 (N_5694,N_3592,N_4577);
nor U5695 (N_5695,N_1200,N_4807);
nand U5696 (N_5696,N_1208,N_54);
xnor U5697 (N_5697,N_427,N_2119);
nand U5698 (N_5698,N_4813,N_4414);
or U5699 (N_5699,N_974,N_2261);
nand U5700 (N_5700,N_4000,N_4570);
or U5701 (N_5701,N_2753,N_45);
xnor U5702 (N_5702,N_1499,N_1976);
nand U5703 (N_5703,N_2040,N_1876);
and U5704 (N_5704,N_1864,N_4999);
or U5705 (N_5705,N_2039,N_4241);
and U5706 (N_5706,N_1987,N_2107);
and U5707 (N_5707,N_3796,N_4764);
nor U5708 (N_5708,N_3825,N_4636);
or U5709 (N_5709,N_3161,N_4948);
and U5710 (N_5710,N_3300,N_1776);
and U5711 (N_5711,N_4108,N_4749);
and U5712 (N_5712,N_1756,N_3069);
and U5713 (N_5713,N_3378,N_4130);
xor U5714 (N_5714,N_1301,N_3288);
nor U5715 (N_5715,N_519,N_3949);
nor U5716 (N_5716,N_4964,N_3904);
xor U5717 (N_5717,N_1503,N_1734);
and U5718 (N_5718,N_367,N_2509);
and U5719 (N_5719,N_2772,N_2750);
xor U5720 (N_5720,N_4662,N_4854);
or U5721 (N_5721,N_2372,N_1392);
nor U5722 (N_5722,N_1351,N_2884);
nand U5723 (N_5723,N_2542,N_493);
xor U5724 (N_5724,N_2584,N_3472);
or U5725 (N_5725,N_1375,N_4079);
and U5726 (N_5726,N_183,N_1475);
nor U5727 (N_5727,N_983,N_880);
and U5728 (N_5728,N_792,N_2813);
nor U5729 (N_5729,N_3620,N_4011);
and U5730 (N_5730,N_2692,N_1703);
xor U5731 (N_5731,N_1914,N_1697);
or U5732 (N_5732,N_4881,N_59);
or U5733 (N_5733,N_715,N_6);
or U5734 (N_5734,N_1946,N_3674);
and U5735 (N_5735,N_377,N_4056);
xor U5736 (N_5736,N_3521,N_1285);
and U5737 (N_5737,N_2445,N_4296);
nand U5738 (N_5738,N_137,N_3740);
or U5739 (N_5739,N_2842,N_1461);
nand U5740 (N_5740,N_620,N_4624);
nor U5741 (N_5741,N_1708,N_2304);
nor U5742 (N_5742,N_649,N_4865);
and U5743 (N_5743,N_789,N_1367);
nor U5744 (N_5744,N_2986,N_2834);
or U5745 (N_5745,N_3415,N_2476);
and U5746 (N_5746,N_3113,N_1355);
xnor U5747 (N_5747,N_1168,N_2118);
nand U5748 (N_5748,N_359,N_1766);
or U5749 (N_5749,N_438,N_988);
and U5750 (N_5750,N_4243,N_1142);
nor U5751 (N_5751,N_4016,N_4591);
xor U5752 (N_5752,N_2703,N_4170);
nand U5753 (N_5753,N_1175,N_1751);
and U5754 (N_5754,N_521,N_4211);
and U5755 (N_5755,N_815,N_1531);
and U5756 (N_5756,N_3001,N_2281);
nor U5757 (N_5757,N_4746,N_2096);
xor U5758 (N_5758,N_2098,N_4316);
xnor U5759 (N_5759,N_3463,N_4237);
nand U5760 (N_5760,N_1311,N_4737);
nor U5761 (N_5761,N_1988,N_2415);
or U5762 (N_5762,N_3008,N_3622);
nand U5763 (N_5763,N_1701,N_347);
nand U5764 (N_5764,N_3449,N_579);
nor U5765 (N_5765,N_3390,N_4689);
xor U5766 (N_5766,N_1815,N_3567);
or U5767 (N_5767,N_4123,N_3100);
xor U5768 (N_5768,N_4143,N_4049);
nor U5769 (N_5769,N_2142,N_3660);
nand U5770 (N_5770,N_1316,N_3081);
nor U5771 (N_5771,N_4615,N_2900);
xor U5772 (N_5772,N_3060,N_1693);
and U5773 (N_5773,N_2012,N_2906);
or U5774 (N_5774,N_4819,N_451);
xnor U5775 (N_5775,N_1489,N_1196);
nor U5776 (N_5776,N_4391,N_2555);
nor U5777 (N_5777,N_2370,N_330);
nand U5778 (N_5778,N_4060,N_1551);
or U5779 (N_5779,N_2669,N_3779);
nand U5780 (N_5780,N_2758,N_1103);
or U5781 (N_5781,N_4740,N_2484);
or U5782 (N_5782,N_633,N_4371);
nand U5783 (N_5783,N_2611,N_1898);
xnor U5784 (N_5784,N_3097,N_4584);
or U5785 (N_5785,N_3890,N_5);
nand U5786 (N_5786,N_4030,N_2577);
and U5787 (N_5787,N_4350,N_720);
or U5788 (N_5788,N_2028,N_4377);
xor U5789 (N_5789,N_1209,N_4550);
nor U5790 (N_5790,N_3369,N_3523);
and U5791 (N_5791,N_4946,N_34);
or U5792 (N_5792,N_1148,N_413);
and U5793 (N_5793,N_2759,N_646);
and U5794 (N_5794,N_2063,N_4131);
or U5795 (N_5795,N_2946,N_3824);
nand U5796 (N_5796,N_932,N_375);
nand U5797 (N_5797,N_4042,N_3241);
nor U5798 (N_5798,N_1318,N_2416);
xor U5799 (N_5799,N_188,N_574);
xnor U5800 (N_5800,N_4498,N_4236);
and U5801 (N_5801,N_1720,N_1412);
nor U5802 (N_5802,N_3244,N_4779);
or U5803 (N_5803,N_2590,N_501);
nand U5804 (N_5804,N_4203,N_2966);
xor U5805 (N_5805,N_4066,N_2762);
nand U5806 (N_5806,N_1231,N_4148);
xor U5807 (N_5807,N_4838,N_986);
xor U5808 (N_5808,N_4275,N_85);
xnor U5809 (N_5809,N_4658,N_1811);
xnor U5810 (N_5810,N_3730,N_3437);
xnor U5811 (N_5811,N_3540,N_2134);
and U5812 (N_5812,N_2575,N_2366);
nor U5813 (N_5813,N_2770,N_4748);
xor U5814 (N_5814,N_610,N_3252);
and U5815 (N_5815,N_1637,N_4769);
xnor U5816 (N_5816,N_1162,N_4102);
or U5817 (N_5817,N_1210,N_4911);
nand U5818 (N_5818,N_1966,N_4809);
nor U5819 (N_5819,N_3187,N_3238);
and U5820 (N_5820,N_1581,N_2716);
xor U5821 (N_5821,N_1479,N_2394);
or U5822 (N_5822,N_2364,N_3794);
or U5823 (N_5823,N_2449,N_4778);
or U5824 (N_5824,N_3401,N_4511);
and U5825 (N_5825,N_3585,N_691);
nor U5826 (N_5826,N_1934,N_4750);
and U5827 (N_5827,N_4679,N_4213);
nor U5828 (N_5828,N_2338,N_1822);
xor U5829 (N_5829,N_2439,N_1680);
xnor U5830 (N_5830,N_1073,N_2137);
nand U5831 (N_5831,N_1825,N_205);
nand U5832 (N_5832,N_3118,N_2887);
or U5833 (N_5833,N_4194,N_1540);
nand U5834 (N_5834,N_3910,N_4501);
xor U5835 (N_5835,N_2027,N_3022);
nand U5836 (N_5836,N_1862,N_4251);
or U5837 (N_5837,N_341,N_1508);
or U5838 (N_5838,N_3803,N_2820);
nor U5839 (N_5839,N_3138,N_1309);
xor U5840 (N_5840,N_3549,N_4848);
nand U5841 (N_5841,N_2761,N_1404);
nor U5842 (N_5842,N_3556,N_3976);
xnor U5843 (N_5843,N_2803,N_2007);
nand U5844 (N_5844,N_2241,N_4869);
or U5845 (N_5845,N_1940,N_2639);
nand U5846 (N_5846,N_4132,N_1279);
or U5847 (N_5847,N_3480,N_3965);
nor U5848 (N_5848,N_1123,N_934);
xor U5849 (N_5849,N_774,N_596);
nor U5850 (N_5850,N_4810,N_668);
nand U5851 (N_5851,N_2272,N_923);
and U5852 (N_5852,N_3848,N_2763);
xnor U5853 (N_5853,N_1356,N_10);
or U5854 (N_5854,N_4507,N_475);
nand U5855 (N_5855,N_4657,N_3326);
xor U5856 (N_5856,N_3783,N_1245);
nor U5857 (N_5857,N_3698,N_4099);
xor U5858 (N_5858,N_3616,N_4733);
nor U5859 (N_5859,N_2726,N_4952);
or U5860 (N_5860,N_4831,N_3488);
nand U5861 (N_5861,N_1880,N_4057);
or U5862 (N_5862,N_3358,N_2956);
or U5863 (N_5863,N_4339,N_1028);
and U5864 (N_5864,N_4762,N_1227);
xor U5865 (N_5865,N_3852,N_499);
nor U5866 (N_5866,N_2133,N_4923);
xnor U5867 (N_5867,N_2886,N_2076);
xnor U5868 (N_5868,N_4171,N_1422);
and U5869 (N_5869,N_4656,N_4549);
or U5870 (N_5870,N_1534,N_4735);
and U5871 (N_5871,N_1904,N_392);
or U5872 (N_5872,N_3725,N_3935);
or U5873 (N_5873,N_133,N_1681);
or U5874 (N_5874,N_1632,N_342);
nor U5875 (N_5875,N_670,N_328);
nand U5876 (N_5876,N_3940,N_3332);
and U5877 (N_5877,N_3121,N_3345);
or U5878 (N_5878,N_4105,N_4940);
or U5879 (N_5879,N_2455,N_1989);
and U5880 (N_5880,N_3299,N_473);
nand U5881 (N_5881,N_418,N_3030);
xnor U5882 (N_5882,N_3328,N_2615);
or U5883 (N_5883,N_2992,N_4159);
nor U5884 (N_5884,N_89,N_2308);
nand U5885 (N_5885,N_632,N_2208);
nand U5886 (N_5886,N_3343,N_1042);
or U5887 (N_5887,N_1810,N_2972);
nand U5888 (N_5888,N_1656,N_2365);
nand U5889 (N_5889,N_3204,N_1280);
nor U5890 (N_5890,N_897,N_2566);
and U5891 (N_5891,N_268,N_93);
nand U5892 (N_5892,N_1626,N_2240);
xor U5893 (N_5893,N_1859,N_1902);
xnor U5894 (N_5894,N_1029,N_4835);
nand U5895 (N_5895,N_4515,N_302);
and U5896 (N_5896,N_2665,N_794);
nor U5897 (N_5897,N_4641,N_1757);
nand U5898 (N_5898,N_4544,N_1349);
xor U5899 (N_5899,N_790,N_3654);
and U5900 (N_5900,N_3432,N_3882);
xor U5901 (N_5901,N_3202,N_561);
and U5902 (N_5902,N_2628,N_778);
and U5903 (N_5903,N_4600,N_202);
and U5904 (N_5904,N_2256,N_566);
and U5905 (N_5905,N_638,N_195);
or U5906 (N_5906,N_4218,N_1516);
nor U5907 (N_5907,N_2010,N_2616);
and U5908 (N_5908,N_766,N_742);
nor U5909 (N_5909,N_1296,N_2789);
nor U5910 (N_5910,N_4466,N_2153);
and U5911 (N_5911,N_3357,N_4728);
or U5912 (N_5912,N_114,N_233);
nand U5913 (N_5913,N_2866,N_128);
xnor U5914 (N_5914,N_101,N_767);
and U5915 (N_5915,N_149,N_4352);
or U5916 (N_5916,N_841,N_4578);
nand U5917 (N_5917,N_1777,N_1533);
nor U5918 (N_5918,N_4385,N_4374);
nor U5919 (N_5919,N_4095,N_1139);
nor U5920 (N_5920,N_1118,N_1384);
and U5921 (N_5921,N_70,N_2458);
and U5922 (N_5922,N_2109,N_2495);
nand U5923 (N_5923,N_3230,N_2967);
nor U5924 (N_5924,N_1716,N_2614);
nor U5925 (N_5925,N_2075,N_3405);
xor U5926 (N_5926,N_2527,N_33);
or U5927 (N_5927,N_4073,N_3921);
nand U5928 (N_5928,N_4627,N_4358);
or U5929 (N_5929,N_490,N_352);
nand U5930 (N_5930,N_3105,N_3982);
and U5931 (N_5931,N_4847,N_1921);
and U5932 (N_5932,N_416,N_2334);
and U5933 (N_5933,N_4281,N_2650);
and U5934 (N_5934,N_3421,N_2624);
or U5935 (N_5935,N_4103,N_1464);
or U5936 (N_5936,N_4260,N_4933);
and U5937 (N_5937,N_3431,N_3360);
xor U5938 (N_5938,N_1746,N_3748);
or U5939 (N_5939,N_2490,N_3075);
nor U5940 (N_5940,N_4395,N_1173);
or U5941 (N_5941,N_2276,N_739);
and U5942 (N_5942,N_487,N_3320);
or U5943 (N_5943,N_1573,N_3074);
nand U5944 (N_5944,N_3071,N_4359);
nand U5945 (N_5945,N_4514,N_4996);
and U5946 (N_5946,N_1183,N_4905);
and U5947 (N_5947,N_3810,N_3251);
xor U5948 (N_5948,N_1995,N_2592);
nor U5949 (N_5949,N_2036,N_2424);
and U5950 (N_5950,N_835,N_3234);
nand U5951 (N_5951,N_4214,N_2398);
nand U5952 (N_5952,N_3636,N_904);
xor U5953 (N_5953,N_2943,N_2617);
nand U5954 (N_5954,N_3853,N_2454);
xnor U5955 (N_5955,N_1731,N_948);
nor U5956 (N_5956,N_1515,N_4313);
xor U5957 (N_5957,N_1698,N_2844);
and U5958 (N_5958,N_2097,N_4738);
or U5959 (N_5959,N_1263,N_1150);
or U5960 (N_5960,N_3776,N_2735);
nor U5961 (N_5961,N_4258,N_4456);
xor U5962 (N_5962,N_2729,N_324);
xnor U5963 (N_5963,N_3808,N_1608);
xnor U5964 (N_5964,N_2898,N_2265);
xnor U5965 (N_5965,N_3880,N_699);
nor U5966 (N_5966,N_577,N_4334);
nand U5967 (N_5967,N_3741,N_951);
or U5968 (N_5968,N_79,N_3689);
nor U5969 (N_5969,N_4518,N_1061);
xor U5970 (N_5970,N_1523,N_3047);
or U5971 (N_5971,N_1261,N_95);
or U5972 (N_5972,N_4558,N_3015);
xor U5973 (N_5973,N_3692,N_1074);
and U5974 (N_5974,N_2506,N_4647);
and U5975 (N_5975,N_3606,N_1802);
xnor U5976 (N_5976,N_160,N_4094);
nor U5977 (N_5977,N_881,N_804);
and U5978 (N_5978,N_4638,N_4755);
or U5979 (N_5979,N_3225,N_3208);
xnor U5980 (N_5980,N_985,N_4437);
nand U5981 (N_5981,N_4179,N_4078);
or U5982 (N_5982,N_1040,N_3568);
nand U5983 (N_5983,N_1110,N_1333);
or U5984 (N_5984,N_3158,N_1440);
xor U5985 (N_5985,N_2680,N_2938);
or U5986 (N_5986,N_665,N_606);
or U5987 (N_5987,N_631,N_2603);
or U5988 (N_5988,N_1132,N_3911);
and U5989 (N_5989,N_4714,N_2311);
and U5990 (N_5990,N_175,N_4698);
or U5991 (N_5991,N_4390,N_2683);
nor U5992 (N_5992,N_4818,N_4416);
or U5993 (N_5993,N_1302,N_2019);
nor U5994 (N_5994,N_1419,N_2404);
nand U5995 (N_5995,N_444,N_1633);
and U5996 (N_5996,N_150,N_373);
or U5997 (N_5997,N_398,N_3802);
nand U5998 (N_5998,N_198,N_1149);
nand U5999 (N_5999,N_3491,N_3271);
or U6000 (N_6000,N_4020,N_4909);
and U6001 (N_6001,N_3898,N_4117);
or U6002 (N_6002,N_4571,N_3785);
xnor U6003 (N_6003,N_256,N_3135);
nand U6004 (N_6004,N_3356,N_4616);
and U6005 (N_6005,N_4950,N_1084);
xnor U6006 (N_6006,N_3446,N_528);
and U6007 (N_6007,N_2100,N_2300);
nand U6008 (N_6008,N_3531,N_4463);
xnor U6009 (N_6009,N_1057,N_3618);
or U6010 (N_6010,N_4404,N_1577);
xnor U6011 (N_6011,N_2623,N_4994);
xnor U6012 (N_6012,N_1024,N_3250);
xnor U6013 (N_6013,N_2620,N_4029);
nand U6014 (N_6014,N_3986,N_2985);
nor U6015 (N_6015,N_1781,N_4727);
nand U6016 (N_6016,N_2843,N_4985);
or U6017 (N_6017,N_3933,N_2382);
or U6018 (N_6018,N_2830,N_1122);
and U6019 (N_6019,N_748,N_4293);
nand U6020 (N_6020,N_303,N_4672);
and U6021 (N_6021,N_457,N_1672);
nand U6022 (N_6022,N_3663,N_1378);
nand U6023 (N_6023,N_158,N_2621);
nand U6024 (N_6024,N_685,N_4134);
or U6025 (N_6025,N_3579,N_1145);
xor U6026 (N_6026,N_4646,N_2318);
xnor U6027 (N_6027,N_1290,N_2529);
and U6028 (N_6028,N_1332,N_1974);
nand U6029 (N_6029,N_3704,N_2725);
or U6030 (N_6030,N_3952,N_3681);
xnor U6031 (N_6031,N_321,N_2540);
nand U6032 (N_6032,N_3219,N_68);
nand U6033 (N_6033,N_2179,N_3557);
nor U6034 (N_6034,N_1023,N_3026);
xor U6035 (N_6035,N_1036,N_2541);
xnor U6036 (N_6036,N_3514,N_2807);
xor U6037 (N_6037,N_4626,N_2786);
or U6038 (N_6038,N_278,N_2819);
and U6039 (N_6039,N_3376,N_2368);
xnor U6040 (N_6040,N_4383,N_3889);
or U6041 (N_6041,N_1037,N_4098);
nand U6042 (N_6042,N_2245,N_3723);
and U6043 (N_6043,N_1448,N_2664);
nand U6044 (N_6044,N_4141,N_346);
nand U6045 (N_6045,N_3364,N_2400);
and U6046 (N_6046,N_2419,N_4866);
nand U6047 (N_6047,N_3902,N_2286);
nor U6048 (N_6048,N_623,N_3058);
xor U6049 (N_6049,N_318,N_1932);
and U6050 (N_6050,N_1817,N_1250);
nand U6051 (N_6051,N_3901,N_4925);
or U6052 (N_6052,N_1942,N_3414);
and U6053 (N_6053,N_3507,N_3322);
xor U6054 (N_6054,N_3402,N_3341);
and U6055 (N_6055,N_4336,N_3767);
and U6056 (N_6056,N_2773,N_1402);
and U6057 (N_6057,N_4230,N_3879);
xor U6058 (N_6058,N_4771,N_4858);
nor U6059 (N_6059,N_3457,N_3972);
nor U6060 (N_6060,N_1243,N_4088);
nor U6061 (N_6061,N_2998,N_1861);
xnor U6062 (N_6062,N_3637,N_378);
nand U6063 (N_6063,N_4384,N_522);
xnor U6064 (N_6064,N_2051,N_2962);
nand U6065 (N_6065,N_4465,N_3993);
xor U6066 (N_6066,N_4907,N_4077);
or U6067 (N_6067,N_3977,N_1759);
nor U6068 (N_6068,N_2407,N_884);
and U6069 (N_6069,N_4852,N_672);
nand U6070 (N_6070,N_2661,N_3504);
nand U6071 (N_6071,N_369,N_119);
nand U6072 (N_6072,N_4247,N_4263);
nand U6073 (N_6073,N_4119,N_274);
or U6074 (N_6074,N_3835,N_1505);
xor U6075 (N_6075,N_1293,N_2648);
or U6076 (N_6076,N_4697,N_2500);
or U6077 (N_6077,N_2778,N_4873);
or U6078 (N_6078,N_3708,N_1799);
or U6079 (N_6079,N_4431,N_2053);
xor U6080 (N_6080,N_737,N_1260);
and U6081 (N_6081,N_3842,N_3875);
nand U6082 (N_6082,N_3999,N_2989);
xor U6083 (N_6083,N_2701,N_2081);
and U6084 (N_6084,N_3086,N_3601);
nor U6085 (N_6085,N_3334,N_719);
or U6086 (N_6086,N_4568,N_4836);
nand U6087 (N_6087,N_3042,N_4447);
xor U6088 (N_6088,N_3506,N_2999);
xnor U6089 (N_6089,N_2341,N_2132);
nand U6090 (N_6090,N_2700,N_4186);
or U6091 (N_6091,N_4796,N_139);
or U6092 (N_6092,N_3738,N_3988);
nor U6093 (N_6093,N_1790,N_4864);
nor U6094 (N_6094,N_1131,N_1853);
xnor U6095 (N_6095,N_1749,N_3384);
nand U6096 (N_6096,N_3221,N_846);
xnor U6097 (N_6097,N_734,N_4196);
and U6098 (N_6098,N_4265,N_1410);
nand U6099 (N_6099,N_2799,N_2755);
and U6100 (N_6100,N_2874,N_921);
nand U6101 (N_6101,N_1415,N_1692);
xor U6102 (N_6102,N_2343,N_112);
and U6103 (N_6103,N_400,N_2044);
xnor U6104 (N_6104,N_2414,N_860);
and U6105 (N_6105,N_4610,N_593);
and U6106 (N_6106,N_2739,N_4107);
xor U6107 (N_6107,N_1643,N_1470);
nand U6108 (N_6108,N_3678,N_1529);
and U6109 (N_6109,N_3453,N_2047);
or U6110 (N_6110,N_4022,N_4747);
nor U6111 (N_6111,N_2519,N_4583);
nor U6112 (N_6112,N_2635,N_4904);
nand U6113 (N_6113,N_4770,N_2917);
xor U6114 (N_6114,N_1836,N_3656);
and U6115 (N_6115,N_1557,N_1035);
and U6116 (N_6116,N_3485,N_107);
xor U6117 (N_6117,N_2131,N_1718);
or U6118 (N_6118,N_1871,N_621);
nand U6119 (N_6119,N_3683,N_2169);
or U6120 (N_6120,N_4277,N_4223);
nor U6121 (N_6121,N_3217,N_4183);
nor U6122 (N_6122,N_1174,N_1011);
or U6123 (N_6123,N_2093,N_2337);
or U6124 (N_6124,N_2899,N_4467);
or U6125 (N_6125,N_4632,N_4916);
nor U6126 (N_6126,N_1119,N_172);
or U6127 (N_6127,N_446,N_761);
or U6128 (N_6128,N_3849,N_4329);
nor U6129 (N_6129,N_2413,N_4133);
or U6130 (N_6130,N_2605,N_937);
xnor U6131 (N_6131,N_1049,N_2749);
nor U6132 (N_6132,N_279,N_1030);
and U6133 (N_6133,N_2976,N_4582);
or U6134 (N_6134,N_2103,N_2918);
or U6135 (N_6135,N_4249,N_3224);
xnor U6136 (N_6136,N_595,N_3460);
xnor U6137 (N_6137,N_4997,N_3951);
or U6138 (N_6138,N_4759,N_1405);
nand U6139 (N_6139,N_1085,N_434);
xor U6140 (N_6140,N_3728,N_712);
or U6141 (N_6141,N_286,N_1748);
and U6142 (N_6142,N_1600,N_2494);
and U6143 (N_6143,N_3749,N_848);
nand U6144 (N_6144,N_664,N_2298);
and U6145 (N_6145,N_527,N_1344);
or U6146 (N_6146,N_1563,N_4309);
nor U6147 (N_6147,N_532,N_2702);
xnor U6148 (N_6148,N_2162,N_4394);
xnor U6149 (N_6149,N_3035,N_1441);
nand U6150 (N_6150,N_2466,N_4503);
xor U6151 (N_6151,N_111,N_782);
xor U6152 (N_6152,N_214,N_27);
and U6153 (N_6153,N_4888,N_1834);
nor U6154 (N_6154,N_1418,N_177);
nand U6155 (N_6155,N_889,N_219);
and U6156 (N_6156,N_2814,N_1182);
nor U6157 (N_6157,N_433,N_1317);
nor U6158 (N_6158,N_830,N_2698);
xor U6159 (N_6159,N_4734,N_2425);
xnor U6160 (N_6160,N_1205,N_3125);
or U6161 (N_6161,N_1587,N_4019);
or U6162 (N_6162,N_2423,N_4788);
xnor U6163 (N_6163,N_3766,N_1324);
or U6164 (N_6164,N_4618,N_2908);
nor U6165 (N_6165,N_4798,N_945);
or U6166 (N_6166,N_3236,N_1783);
nand U6167 (N_6167,N_4529,N_1971);
nor U6168 (N_6168,N_383,N_4562);
nor U6169 (N_6169,N_3747,N_1958);
xor U6170 (N_6170,N_2627,N_365);
nor U6171 (N_6171,N_1816,N_220);
nor U6172 (N_6172,N_4067,N_2369);
and U6173 (N_6173,N_4367,N_1621);
or U6174 (N_6174,N_2371,N_3587);
nor U6175 (N_6175,N_1154,N_3544);
nand U6176 (N_6176,N_2794,N_3153);
or U6177 (N_6177,N_4797,N_3165);
xor U6178 (N_6178,N_456,N_113);
and U6179 (N_6179,N_1299,N_2825);
nand U6180 (N_6180,N_4231,N_1714);
or U6181 (N_6181,N_4761,N_4783);
xor U6182 (N_6182,N_1069,N_395);
xnor U6183 (N_6183,N_245,N_3696);
xnor U6184 (N_6184,N_3178,N_4474);
and U6185 (N_6185,N_1705,N_2129);
nand U6186 (N_6186,N_1387,N_1067);
and U6187 (N_6187,N_2836,N_2851);
nand U6188 (N_6188,N_2651,N_4893);
or U6189 (N_6189,N_995,N_2247);
nand U6190 (N_6190,N_323,N_1683);
xnor U6191 (N_6191,N_1704,N_2688);
nor U6192 (N_6192,N_4426,N_2751);
nand U6193 (N_6193,N_1201,N_1507);
or U6194 (N_6194,N_2479,N_779);
or U6195 (N_6195,N_3576,N_814);
and U6196 (N_6196,N_4353,N_3426);
xor U6197 (N_6197,N_118,N_3459);
xor U6198 (N_6198,N_612,N_705);
nand U6199 (N_6199,N_90,N_1702);
nand U6200 (N_6200,N_1102,N_1828);
and U6201 (N_6201,N_871,N_2031);
nand U6202 (N_6202,N_2980,N_63);
or U6203 (N_6203,N_4942,N_2145);
xnor U6204 (N_6204,N_4782,N_3468);
and U6205 (N_6205,N_2203,N_2252);
xnor U6206 (N_6206,N_628,N_569);
or U6207 (N_6207,N_4793,N_1831);
nand U6208 (N_6208,N_2048,N_4013);
or U6209 (N_6209,N_2630,N_3264);
xor U6210 (N_6210,N_1190,N_1377);
xor U6211 (N_6211,N_3775,N_2668);
xor U6212 (N_6212,N_422,N_4112);
xor U6213 (N_6213,N_2608,N_4603);
nand U6214 (N_6214,N_2676,N_4745);
nor U6215 (N_6215,N_2268,N_2730);
nor U6216 (N_6216,N_2015,N_4335);
nor U6217 (N_6217,N_3013,N_315);
xnor U6218 (N_6218,N_746,N_1125);
nand U6219 (N_6219,N_4709,N_2292);
nand U6220 (N_6220,N_732,N_3868);
or U6221 (N_6221,N_1770,N_666);
nand U6222 (N_6222,N_3375,N_1224);
and U6223 (N_6223,N_3249,N_1498);
and U6224 (N_6224,N_2564,N_1140);
or U6225 (N_6225,N_1474,N_3192);
nand U6226 (N_6226,N_4725,N_4208);
or U6227 (N_6227,N_2211,N_3648);
and U6228 (N_6228,N_3080,N_3811);
nor U6229 (N_6229,N_4007,N_689);
nand U6230 (N_6230,N_2774,N_4694);
nor U6231 (N_6231,N_1682,N_4321);
nand U6232 (N_6232,N_2173,N_4595);
or U6233 (N_6233,N_1282,N_4901);
nand U6234 (N_6234,N_2320,N_1086);
xor U6235 (N_6235,N_2872,N_4052);
xnor U6236 (N_6236,N_607,N_3354);
and U6237 (N_6237,N_1575,N_626);
or U6238 (N_6238,N_4082,N_3098);
and U6239 (N_6239,N_1654,N_1627);
nor U6240 (N_6240,N_4115,N_785);
nand U6241 (N_6241,N_3272,N_4442);
or U6242 (N_6242,N_316,N_2586);
nor U6243 (N_6243,N_1490,N_1872);
nor U6244 (N_6244,N_3265,N_1347);
and U6245 (N_6245,N_3434,N_4291);
or U6246 (N_6246,N_4392,N_3603);
or U6247 (N_6247,N_4199,N_3031);
xor U6248 (N_6248,N_3211,N_2699);
xnor U6249 (N_6249,N_3245,N_3422);
xor U6250 (N_6250,N_264,N_41);
nand U6251 (N_6251,N_2099,N_505);
and U6252 (N_6252,N_3684,N_3623);
or U6253 (N_6253,N_977,N_4977);
nor U6254 (N_6254,N_4191,N_688);
or U6255 (N_6255,N_223,N_4182);
xor U6256 (N_6256,N_3937,N_1159);
or U6257 (N_6257,N_4162,N_3292);
or U6258 (N_6258,N_1929,N_265);
xnor U6259 (N_6259,N_3041,N_3403);
nand U6260 (N_6260,N_3130,N_243);
xor U6261 (N_6261,N_2928,N_821);
or U6262 (N_6262,N_3014,N_136);
nor U6263 (N_6263,N_3746,N_502);
nand U6264 (N_6264,N_16,N_283);
nand U6265 (N_6265,N_3672,N_1947);
nor U6266 (N_6266,N_4552,N_1584);
or U6267 (N_6267,N_4046,N_1850);
nand U6268 (N_6268,N_654,N_4765);
nand U6269 (N_6269,N_3055,N_3191);
and U6270 (N_6270,N_1826,N_2058);
and U6271 (N_6271,N_2877,N_3167);
nand U6272 (N_6272,N_2150,N_253);
nand U6273 (N_6273,N_2387,N_1913);
xnor U6274 (N_6274,N_2777,N_4412);
xor U6275 (N_6275,N_2606,N_2359);
or U6276 (N_6276,N_4014,N_2559);
nor U6277 (N_6277,N_4958,N_4378);
nand U6278 (N_6278,N_3836,N_2326);
or U6279 (N_6279,N_9,N_4890);
nand U6280 (N_6280,N_567,N_2144);
xnor U6281 (N_6281,N_1350,N_1264);
and U6282 (N_6282,N_1456,N_3172);
nand U6283 (N_6283,N_4572,N_1071);
xor U6284 (N_6284,N_3726,N_3475);
nand U6285 (N_6285,N_629,N_4304);
nor U6286 (N_6286,N_2034,N_1199);
and U6287 (N_6287,N_2397,N_3451);
xnor U6288 (N_6288,N_2002,N_2652);
nand U6289 (N_6289,N_3773,N_3737);
nand U6290 (N_6290,N_1619,N_2862);
or U6291 (N_6291,N_2428,N_1953);
and U6292 (N_6292,N_3520,N_4534);
nor U6293 (N_6293,N_4089,N_2654);
xnor U6294 (N_6294,N_4234,N_2282);
or U6295 (N_6295,N_3733,N_105);
nor U6296 (N_6296,N_3818,N_4699);
or U6297 (N_6297,N_1100,N_2430);
nand U6298 (N_6298,N_4348,N_4091);
nand U6299 (N_6299,N_3285,N_1058);
xnor U6300 (N_6300,N_1715,N_4396);
nand U6301 (N_6301,N_2678,N_2296);
xor U6302 (N_6302,N_3386,N_3452);
and U6303 (N_6303,N_1371,N_3053);
nor U6304 (N_6304,N_4839,N_2731);
or U6305 (N_6305,N_1991,N_246);
xnor U6306 (N_6306,N_706,N_3867);
and U6307 (N_6307,N_3283,N_4789);
xor U6308 (N_6308,N_1541,N_3615);
or U6309 (N_6309,N_2167,N_312);
and U6310 (N_6310,N_1750,N_2226);
and U6311 (N_6311,N_1312,N_3985);
nor U6312 (N_6312,N_4563,N_795);
and U6313 (N_6313,N_384,N_538);
nor U6314 (N_6314,N_1585,N_4889);
nor U6315 (N_6315,N_2486,N_1446);
or U6316 (N_6316,N_2487,N_3547);
nand U6317 (N_6317,N_1945,N_3679);
or U6318 (N_6318,N_3087,N_2234);
and U6319 (N_6319,N_1093,N_4989);
or U6320 (N_6320,N_1710,N_4876);
xor U6321 (N_6321,N_1158,N_864);
and U6322 (N_6322,N_4153,N_3885);
or U6323 (N_6323,N_4387,N_4811);
and U6324 (N_6324,N_4871,N_1229);
xor U6325 (N_6325,N_1330,N_2465);
nand U6326 (N_6326,N_4044,N_2194);
nand U6327 (N_6327,N_259,N_18);
xnor U6328 (N_6328,N_2214,N_960);
xor U6329 (N_6329,N_4420,N_100);
nand U6330 (N_6330,N_4537,N_293);
and U6331 (N_6331,N_1130,N_2110);
and U6332 (N_6332,N_944,N_4717);
nand U6333 (N_6333,N_2383,N_4774);
nor U6334 (N_6334,N_2317,N_3581);
and U6335 (N_6335,N_1425,N_4918);
and U6336 (N_6336,N_4031,N_2727);
xor U6337 (N_6337,N_2609,N_2470);
and U6338 (N_6338,N_3054,N_2460);
xnor U6339 (N_6339,N_3339,N_4981);
xnor U6340 (N_6340,N_957,N_2784);
xor U6341 (N_6341,N_4212,N_3563);
nand U6342 (N_6342,N_1687,N_1675);
xor U6343 (N_6343,N_4349,N_4421);
and U6344 (N_6344,N_1740,N_572);
or U6345 (N_6345,N_4055,N_1897);
and U6346 (N_6346,N_4167,N_4303);
or U6347 (N_6347,N_752,N_3056);
nand U6348 (N_6348,N_4455,N_2160);
nand U6349 (N_6349,N_796,N_407);
or U6350 (N_6350,N_3176,N_1968);
nand U6351 (N_6351,N_731,N_1135);
xnor U6352 (N_6352,N_2822,N_1374);
or U6353 (N_6353,N_4566,N_2497);
xnor U6354 (N_6354,N_998,N_695);
nand U6355 (N_6355,N_1524,N_368);
xnor U6356 (N_6356,N_4743,N_594);
xor U6357 (N_6357,N_2571,N_3377);
and U6358 (N_6358,N_4033,N_492);
and U6359 (N_6359,N_1427,N_3193);
nand U6360 (N_6360,N_1284,N_1835);
xor U6361 (N_6361,N_2587,N_4092);
or U6362 (N_6362,N_2046,N_1630);
nand U6363 (N_6363,N_1618,N_2290);
nor U6364 (N_6364,N_971,N_186);
nand U6365 (N_6365,N_356,N_662);
xnor U6366 (N_6366,N_1117,N_3374);
or U6367 (N_6367,N_975,N_4054);
or U6368 (N_6368,N_4795,N_2800);
nand U6369 (N_6369,N_3284,N_1891);
nand U6370 (N_6370,N_2174,N_1517);
nand U6371 (N_6371,N_3543,N_329);
nand U6372 (N_6372,N_1688,N_1646);
nor U6373 (N_6373,N_2568,N_1560);
nand U6374 (N_6374,N_4254,N_2310);
or U6375 (N_6375,N_1176,N_292);
or U6376 (N_6376,N_1844,N_1765);
xnor U6377 (N_6377,N_1025,N_3209);
and U6378 (N_6378,N_892,N_38);
nor U6379 (N_6379,N_170,N_807);
and U6380 (N_6380,N_859,N_1463);
nand U6381 (N_6381,N_681,N_3732);
nand U6382 (N_6382,N_1635,N_568);
nor U6383 (N_6383,N_1393,N_2674);
or U6384 (N_6384,N_1920,N_2978);
nand U6385 (N_6385,N_471,N_4532);
nor U6386 (N_6386,N_4664,N_2262);
or U6387 (N_6387,N_1593,N_4988);
xnor U6388 (N_6388,N_659,N_3718);
and U6389 (N_6389,N_3956,N_3246);
nor U6390 (N_6390,N_3018,N_1512);
or U6391 (N_6391,N_1933,N_4147);
nor U6392 (N_6392,N_3247,N_3350);
nor U6393 (N_6393,N_4021,N_1386);
xor U6394 (N_6394,N_4791,N_3063);
or U6395 (N_6395,N_2818,N_2035);
xor U6396 (N_6396,N_1095,N_2190);
or U6397 (N_6397,N_917,N_2920);
nor U6398 (N_6398,N_143,N_966);
and U6399 (N_6399,N_2438,N_362);
xnor U6400 (N_6400,N_4596,N_2030);
or U6401 (N_6401,N_83,N_1634);
and U6402 (N_6402,N_996,N_1544);
or U6403 (N_6403,N_740,N_4435);
and U6404 (N_6404,N_3657,N_2880);
xor U6405 (N_6405,N_4520,N_2582);
and U6406 (N_6406,N_3655,N_442);
nand U6407 (N_6407,N_4343,N_1549);
nand U6408 (N_6408,N_182,N_3862);
or U6409 (N_6409,N_4661,N_1798);
or U6410 (N_6410,N_240,N_3101);
or U6411 (N_6411,N_2597,N_271);
xor U6412 (N_6412,N_1391,N_3445);
or U6413 (N_6413,N_973,N_3858);
nand U6414 (N_6414,N_4439,N_4730);
nand U6415 (N_6415,N_4195,N_1141);
nor U6416 (N_6416,N_554,N_4973);
or U6417 (N_6417,N_2636,N_4992);
nand U6418 (N_6418,N_1275,N_3967);
and U6419 (N_6419,N_349,N_2963);
xor U6420 (N_6420,N_2389,N_1113);
nor U6421 (N_6421,N_4931,N_3382);
nor U6422 (N_6422,N_2377,N_1286);
and U6423 (N_6423,N_2037,N_3734);
nand U6424 (N_6424,N_2508,N_3243);
nand U6425 (N_6425,N_4516,N_3973);
xor U6426 (N_6426,N_295,N_2180);
xor U6427 (N_6427,N_3148,N_1548);
and U6428 (N_6428,N_2850,N_4654);
and U6429 (N_6429,N_4040,N_907);
nor U6430 (N_6430,N_2790,N_747);
xor U6431 (N_6431,N_3997,N_2325);
nand U6432 (N_6432,N_1328,N_2845);
and U6433 (N_6433,N_4287,N_1437);
xor U6434 (N_6434,N_4295,N_2498);
nor U6435 (N_6435,N_1129,N_1917);
nand U6436 (N_6436,N_2087,N_3455);
nand U6437 (N_6437,N_3359,N_4417);
and U6438 (N_6438,N_180,N_3309);
and U6439 (N_6439,N_3974,N_4919);
nor U6440 (N_6440,N_4711,N_4315);
and U6441 (N_6441,N_1907,N_4149);
nor U6442 (N_6442,N_1034,N_4939);
xnor U6443 (N_6443,N_1407,N_2744);
or U6444 (N_6444,N_1962,N_4494);
and U6445 (N_6445,N_1225,N_2948);
and U6446 (N_6446,N_3458,N_3686);
nand U6447 (N_6447,N_531,N_1255);
or U6448 (N_6448,N_2077,N_4960);
nand U6449 (N_6449,N_452,N_3305);
nand U6450 (N_6450,N_4294,N_4554);
nand U6451 (N_6451,N_2102,N_4928);
nor U6452 (N_6452,N_3450,N_2375);
xor U6453 (N_6453,N_2827,N_1596);
or U6454 (N_6454,N_2175,N_4794);
and U6455 (N_6455,N_1638,N_4462);
xnor U6456 (N_6456,N_3162,N_4273);
nor U6457 (N_6457,N_4780,N_3383);
and U6458 (N_6458,N_2441,N_2488);
nor U6459 (N_6459,N_3505,N_2050);
nor U6460 (N_6460,N_148,N_1303);
and U6461 (N_6461,N_4991,N_1662);
nand U6462 (N_6462,N_3550,N_2258);
nand U6463 (N_6463,N_1232,N_1124);
nor U6464 (N_6464,N_856,N_1062);
xor U6465 (N_6465,N_3177,N_1421);
nor U6466 (N_6466,N_176,N_2622);
nand U6467 (N_6467,N_4486,N_4235);
or U6468 (N_6468,N_1572,N_4608);
nand U6469 (N_6469,N_1435,N_3770);
and U6470 (N_6470,N_1819,N_74);
nor U6471 (N_6471,N_2378,N_3242);
xor U6472 (N_6472,N_294,N_117);
xnor U6473 (N_6473,N_353,N_743);
or U6474 (N_6474,N_3103,N_3276);
nor U6475 (N_6475,N_103,N_2625);
or U6476 (N_6476,N_1775,N_3782);
nand U6477 (N_6477,N_738,N_4927);
xor U6478 (N_6478,N_4478,N_2266);
xnor U6479 (N_6479,N_4206,N_4480);
or U6480 (N_6480,N_2723,N_1792);
nand U6481 (N_6481,N_3908,N_3855);
nor U6482 (N_6482,N_4851,N_49);
and U6483 (N_6483,N_1931,N_4786);
or U6484 (N_6484,N_604,N_3477);
or U6485 (N_6485,N_4724,N_4965);
nor U6486 (N_6486,N_4093,N_3073);
and U6487 (N_6487,N_3304,N_3003);
nor U6488 (N_6488,N_852,N_4908);
or U6489 (N_6489,N_1457,N_3677);
or U6490 (N_6490,N_4441,N_75);
nor U6491 (N_6491,N_4756,N_1924);
or U6492 (N_6492,N_1,N_1741);
xor U6493 (N_6493,N_73,N_445);
nor U6494 (N_6494,N_4850,N_3070);
nand U6495 (N_6495,N_2684,N_3533);
xnor U6496 (N_6496,N_3578,N_818);
nand U6497 (N_6497,N_1426,N_939);
or U6498 (N_6498,N_3553,N_3722);
xnor U6499 (N_6499,N_3394,N_2523);
xnor U6500 (N_6500,N_2178,N_2821);
xor U6501 (N_6501,N_3720,N_2732);
nand U6502 (N_6502,N_1722,N_1724);
nor U6503 (N_6503,N_1949,N_526);
nor U6504 (N_6504,N_1824,N_701);
nor U6505 (N_6505,N_3948,N_3308);
xnor U6506 (N_6506,N_4261,N_4614);
nor U6507 (N_6507,N_3255,N_4799);
or U6508 (N_6508,N_280,N_625);
xnor U6509 (N_6509,N_4801,N_454);
nand U6510 (N_6510,N_2227,N_4004);
xor U6511 (N_6511,N_1774,N_3886);
and U6512 (N_6512,N_3142,N_120);
or U6513 (N_6513,N_4590,N_2483);
xnor U6514 (N_6514,N_3511,N_4862);
nor U6515 (N_6515,N_2912,N_4718);
or U6516 (N_6516,N_1794,N_4681);
or U6517 (N_6517,N_3020,N_2348);
nor U6518 (N_6518,N_2710,N_4372);
and U6519 (N_6519,N_4891,N_2879);
nor U6520 (N_6520,N_4660,N_1221);
or U6521 (N_6521,N_2324,N_1689);
xor U6522 (N_6522,N_541,N_1091);
or U6523 (N_6523,N_656,N_4244);
xor U6524 (N_6524,N_4499,N_2857);
xor U6525 (N_6525,N_4346,N_1064);
xor U6526 (N_6526,N_3939,N_3693);
nand U6527 (N_6527,N_1506,N_2049);
xnor U6528 (N_6528,N_1782,N_1056);
and U6529 (N_6529,N_4732,N_4805);
nand U6530 (N_6530,N_1054,N_1954);
or U6531 (N_6531,N_676,N_4559);
or U6532 (N_6532,N_1445,N_4914);
and U6533 (N_6533,N_3508,N_640);
and U6534 (N_6534,N_3919,N_1166);
xnor U6535 (N_6535,N_1487,N_1978);
xnor U6536 (N_6536,N_2573,N_1996);
nand U6537 (N_6537,N_802,N_2754);
nor U6538 (N_6538,N_217,N_3502);
and U6539 (N_6539,N_1429,N_1578);
and U6540 (N_6540,N_812,N_2127);
nand U6541 (N_6541,N_2926,N_3930);
or U6542 (N_6542,N_3372,N_2215);
nor U6543 (N_6543,N_2524,N_1138);
xnor U6544 (N_6544,N_2890,N_4580);
and U6545 (N_6545,N_35,N_2569);
or U6546 (N_6546,N_4910,N_4445);
and U6547 (N_6547,N_2598,N_4136);
nor U6548 (N_6548,N_4193,N_1396);
nor U6549 (N_6549,N_4075,N_2670);
nor U6550 (N_6550,N_3478,N_2903);
xnor U6551 (N_6551,N_482,N_537);
and U6552 (N_6552,N_506,N_3961);
and U6553 (N_6553,N_3781,N_4792);
nor U6554 (N_6554,N_3586,N_3439);
nor U6555 (N_6555,N_3039,N_4707);
or U6556 (N_6556,N_978,N_4418);
xor U6557 (N_6557,N_2451,N_4344);
nor U6558 (N_6558,N_2657,N_1220);
and U6559 (N_6559,N_1045,N_1583);
nand U6560 (N_6560,N_2062,N_1604);
and U6561 (N_6561,N_1597,N_3040);
xnor U6562 (N_6562,N_4227,N_1408);
and U6563 (N_6563,N_1060,N_3448);
xor U6564 (N_6564,N_66,N_130);
nor U6565 (N_6565,N_2997,N_4829);
xnor U6566 (N_6566,N_2717,N_4892);
nand U6567 (N_6567,N_3807,N_2219);
xnor U6568 (N_6568,N_4599,N_694);
nand U6569 (N_6569,N_963,N_3104);
nor U6570 (N_6570,N_3090,N_4301);
nor U6571 (N_6571,N_4551,N_50);
nor U6572 (N_6572,N_3839,N_102);
nor U6573 (N_6573,N_3388,N_3006);
nor U6574 (N_6574,N_164,N_3916);
nor U6575 (N_6575,N_1164,N_2339);
nand U6576 (N_6576,N_185,N_3361);
nor U6577 (N_6577,N_4849,N_52);
xnor U6578 (N_6578,N_611,N_1768);
nand U6579 (N_6579,N_2826,N_3144);
and U6580 (N_6580,N_4536,N_80);
or U6581 (N_6581,N_4240,N_3412);
nand U6582 (N_6582,N_540,N_4476);
or U6583 (N_6583,N_2779,N_3929);
nor U6584 (N_6584,N_2747,N_4784);
nor U6585 (N_6585,N_801,N_1983);
and U6586 (N_6586,N_879,N_1821);
and U6587 (N_6587,N_4152,N_4264);
nand U6588 (N_6588,N_1009,N_2307);
nand U6589 (N_6589,N_4370,N_1001);
xnor U6590 (N_6590,N_3173,N_3408);
nand U6591 (N_6591,N_47,N_4633);
or U6592 (N_6592,N_4868,N_2408);
nor U6593 (N_6593,N_2868,N_4116);
xor U6594 (N_6594,N_1424,N_722);
nor U6595 (N_6595,N_669,N_4752);
xnor U6596 (N_6596,N_2512,N_2080);
or U6597 (N_6597,N_4715,N_1856);
nor U6598 (N_6598,N_1840,N_2305);
xnor U6599 (N_6599,N_4643,N_467);
or U6600 (N_6600,N_911,N_2257);
or U6601 (N_6601,N_1265,N_1161);
nor U6602 (N_6602,N_4216,N_3690);
nand U6603 (N_6603,N_317,N_1357);
or U6604 (N_6604,N_918,N_3727);
nand U6605 (N_6605,N_3897,N_956);
or U6606 (N_6606,N_4678,N_191);
nor U6607 (N_6607,N_4492,N_3461);
xnor U6608 (N_6608,N_3793,N_2069);
nand U6609 (N_6609,N_1207,N_4087);
or U6610 (N_6610,N_2299,N_2960);
nor U6611 (N_6611,N_2638,N_4495);
nor U6612 (N_6612,N_1137,N_168);
nor U6613 (N_6613,N_4588,N_615);
xor U6614 (N_6614,N_1555,N_4684);
nor U6615 (N_6615,N_4129,N_1493);
nand U6616 (N_6616,N_2278,N_4601);
xor U6617 (N_6617,N_2115,N_3329);
nor U6618 (N_6618,N_2525,N_4118);
and U6619 (N_6619,N_4719,N_211);
or U6620 (N_6620,N_4665,N_680);
xor U6621 (N_6621,N_2721,N_3237);
nor U6622 (N_6622,N_2719,N_4945);
and U6623 (N_6623,N_1420,N_144);
or U6624 (N_6624,N_755,N_1937);
and U6625 (N_6625,N_3154,N_4484);
nand U6626 (N_6626,N_3139,N_4023);
nand U6627 (N_6627,N_2395,N_1252);
xnor U6628 (N_6628,N_4423,N_1624);
nand U6629 (N_6629,N_4690,N_2809);
nor U6630 (N_6630,N_1185,N_2808);
or U6631 (N_6631,N_509,N_3438);
and U6632 (N_6632,N_608,N_2520);
nand U6633 (N_6633,N_348,N_4454);
or U6634 (N_6634,N_4982,N_764);
or U6635 (N_6635,N_4320,N_3228);
and U6636 (N_6636,N_165,N_700);
and U6637 (N_6637,N_1338,N_933);
and U6638 (N_6638,N_4140,N_3979);
nor U6639 (N_6639,N_1300,N_2856);
xor U6640 (N_6640,N_3580,N_787);
nor U6641 (N_6641,N_4479,N_1295);
and U6642 (N_6642,N_2113,N_3023);
xnor U6643 (N_6643,N_4932,N_443);
or U6644 (N_6644,N_3497,N_2535);
or U6645 (N_6645,N_586,N_3613);
nand U6646 (N_6646,N_2468,N_1879);
or U6647 (N_6647,N_4127,N_717);
or U6648 (N_6648,N_2838,N_4446);
nor U6649 (N_6649,N_1485,N_4393);
and U6650 (N_6650,N_3721,N_2947);
nor U6651 (N_6651,N_4508,N_4006);
nand U6652 (N_6652,N_4936,N_1486);
xor U6653 (N_6653,N_479,N_1874);
xor U6654 (N_6654,N_1547,N_2855);
nor U6655 (N_6655,N_4256,N_3947);
and U6656 (N_6656,N_2871,N_1843);
nand U6657 (N_6657,N_2434,N_867);
nand U6658 (N_6658,N_3156,N_1841);
nor U6659 (N_6659,N_3893,N_2462);
nand U6660 (N_6660,N_4912,N_3614);
nand U6661 (N_6661,N_3170,N_2356);
nor U6662 (N_6662,N_3420,N_3476);
or U6663 (N_6663,N_3923,N_551);
or U6664 (N_6664,N_4185,N_560);
or U6665 (N_6665,N_3106,N_2074);
and U6666 (N_6666,N_2122,N_2708);
xor U6667 (N_6667,N_2816,N_4083);
nand U6668 (N_6668,N_914,N_250);
or U6669 (N_6669,N_4980,N_2691);
and U6670 (N_6670,N_46,N_3992);
nor U6671 (N_6671,N_91,N_1323);
and U6672 (N_6672,N_2951,N_3596);
xor U6673 (N_6673,N_1217,N_4144);
xnor U6674 (N_6674,N_4252,N_3799);
and U6675 (N_6675,N_3145,N_335);
nor U6676 (N_6676,N_393,N_2765);
nor U6677 (N_6677,N_2213,N_810);
xor U6678 (N_6678,N_3143,N_126);
and U6679 (N_6679,N_2924,N_3009);
or U6680 (N_6680,N_3286,N_1146);
or U6681 (N_6681,N_4403,N_388);
xnor U6682 (N_6682,N_1969,N_760);
nor U6683 (N_6683,N_1885,N_4915);
xor U6684 (N_6684,N_1046,N_1340);
nor U6685 (N_6685,N_2931,N_4161);
or U6686 (N_6686,N_3537,N_4609);
nand U6687 (N_6687,N_510,N_4369);
xnor U6688 (N_6688,N_2574,N_3397);
nor U6689 (N_6689,N_1380,N_2675);
and U6690 (N_6690,N_757,N_868);
xor U6691 (N_6691,N_570,N_40);
or U6692 (N_6692,N_3653,N_4555);
or U6693 (N_6693,N_4419,N_2482);
nand U6694 (N_6694,N_3963,N_4598);
nor U6695 (N_6695,N_3821,N_2271);
nand U6696 (N_6696,N_460,N_3500);
nand U6697 (N_6697,N_4502,N_291);
nor U6698 (N_6698,N_4587,N_4505);
nand U6699 (N_6699,N_3273,N_671);
and U6700 (N_6700,N_3724,N_4967);
or U6701 (N_6701,N_55,N_3876);
nand U6702 (N_6702,N_2576,N_3454);
nand U6703 (N_6703,N_2543,N_1214);
or U6704 (N_6704,N_3347,N_2092);
nor U6705 (N_6705,N_3925,N_239);
xor U6706 (N_6706,N_1955,N_4409);
and U6707 (N_6707,N_4712,N_309);
nor U6708 (N_6708,N_894,N_4398);
xnor U6709 (N_6709,N_4878,N_3136);
nand U6710 (N_6710,N_4477,N_4804);
and U6711 (N_6711,N_4539,N_563);
or U6712 (N_6712,N_3710,N_2570);
nor U6713 (N_6713,N_122,N_3342);
or U6714 (N_6714,N_4547,N_4068);
nor U6715 (N_6715,N_4921,N_882);
xnor U6716 (N_6716,N_3195,N_2656);
xor U6717 (N_6717,N_4059,N_4617);
nor U6718 (N_6718,N_877,N_3469);
or U6719 (N_6719,N_4885,N_1735);
nand U6720 (N_6720,N_3216,N_4051);
nand U6721 (N_6721,N_3443,N_2502);
or U6722 (N_6722,N_3633,N_2143);
nand U6723 (N_6723,N_3797,N_2521);
nand U6724 (N_6724,N_1986,N_1253);
nor U6725 (N_6725,N_4197,N_4814);
nor U6726 (N_6726,N_99,N_1661);
and U6727 (N_6727,N_3826,N_3828);
xor U6728 (N_6728,N_4189,N_4174);
nand U6729 (N_6729,N_1019,N_1653);
nor U6730 (N_6730,N_21,N_3573);
and U6731 (N_6731,N_2969,N_1700);
and U6732 (N_6732,N_724,N_1017);
and U6733 (N_6733,N_225,N_3164);
or U6734 (N_6734,N_1673,N_423);
or U6735 (N_6735,N_2057,N_2327);
xnor U6736 (N_6736,N_4373,N_2126);
or U6737 (N_6737,N_1812,N_3474);
nor U6738 (N_6738,N_2974,N_1545);
or U6739 (N_6739,N_2687,N_326);
xor U6740 (N_6740,N_4064,N_1712);
nand U6741 (N_6741,N_2629,N_1521);
and U6742 (N_6742,N_4015,N_2667);
nand U6743 (N_6743,N_920,N_43);
nor U6744 (N_6744,N_1063,N_4528);
nand U6745 (N_6745,N_3996,N_1273);
nor U6746 (N_6746,N_3650,N_2600);
nor U6747 (N_6747,N_1818,N_3096);
xnor U6748 (N_6748,N_1726,N_2915);
and U6749 (N_6749,N_3631,N_3554);
xnor U6750 (N_6750,N_1246,N_1187);
nor U6751 (N_6751,N_1291,N_1652);
or U6752 (N_6752,N_2724,N_2170);
xnor U6753 (N_6753,N_135,N_773);
or U6754 (N_6754,N_910,N_4629);
nor U6755 (N_6755,N_1179,N_1400);
nand U6756 (N_6756,N_2117,N_426);
xnor U6757 (N_6757,N_1606,N_3991);
nand U6758 (N_6758,N_36,N_2696);
nand U6759 (N_6759,N_1980,N_845);
nand U6760 (N_6760,N_1916,N_2936);
or U6761 (N_6761,N_2705,N_3293);
nand U6762 (N_6762,N_94,N_1882);
nand U6763 (N_6763,N_2501,N_728);
xnor U6764 (N_6764,N_2349,N_3163);
xor U6765 (N_6765,N_32,N_376);
nand U6766 (N_6766,N_2994,N_2472);
nand U6767 (N_6767,N_4217,N_184);
nor U6768 (N_6768,N_3122,N_331);
xnor U6769 (N_6769,N_3363,N_2882);
xnor U6770 (N_6770,N_1562,N_4630);
and U6771 (N_6771,N_3541,N_653);
nor U6772 (N_6772,N_3827,N_1609);
and U6773 (N_6773,N_2171,N_1511);
nand U6774 (N_6774,N_408,N_304);
xnor U6775 (N_6775,N_4440,N_3697);
xor U6776 (N_6776,N_928,N_762);
xnor U6777 (N_6777,N_828,N_616);
nor U6778 (N_6778,N_530,N_4490);
or U6779 (N_6779,N_2841,N_3479);
nand U6780 (N_6780,N_4180,N_4803);
xnor U6781 (N_6781,N_2767,N_2319);
xor U6782 (N_6782,N_4080,N_1985);
nand U6783 (N_6783,N_2952,N_3171);
nand U6784 (N_6784,N_2640,N_953);
nor U6785 (N_6785,N_4201,N_4109);
or U6786 (N_6786,N_3604,N_4517);
and U6787 (N_6787,N_4037,N_4415);
nor U6788 (N_6788,N_1307,N_4777);
nor U6789 (N_6789,N_3407,N_3888);
and U6790 (N_6790,N_3338,N_2016);
nand U6791 (N_6791,N_3373,N_4944);
and U6792 (N_6792,N_3447,N_648);
or U6793 (N_6793,N_536,N_488);
nand U6794 (N_6794,N_3806,N_2849);
nor U6795 (N_6795,N_1538,N_4178);
xnor U6796 (N_6796,N_4155,N_2913);
or U6797 (N_6797,N_711,N_1565);
xnor U6798 (N_6798,N_498,N_940);
nor U6799 (N_6799,N_1385,N_1833);
nor U6800 (N_6800,N_1999,N_833);
nor U6801 (N_6801,N_1325,N_3594);
xnor U6802 (N_6802,N_4620,N_3319);
and U6803 (N_6803,N_3831,N_4955);
and U6804 (N_6804,N_771,N_2066);
nand U6805 (N_6805,N_229,N_146);
or U6806 (N_6806,N_1875,N_1805);
nand U6807 (N_6807,N_3789,N_3757);
and U6808 (N_6808,N_4493,N_1368);
nor U6809 (N_6809,N_4806,N_1919);
xor U6810 (N_6810,N_3157,N_385);
or U6811 (N_6811,N_3120,N_1570);
nand U6812 (N_6812,N_4979,N_2362);
or U6813 (N_6813,N_424,N_425);
nand U6814 (N_6814,N_949,N_4121);
or U6815 (N_6815,N_1080,N_3942);
nor U6816 (N_6816,N_703,N_3232);
nor U6817 (N_6817,N_2572,N_3181);
and U6818 (N_6818,N_428,N_4606);
nor U6819 (N_6819,N_1785,N_3085);
xnor U6820 (N_6820,N_3774,N_559);
and U6821 (N_6821,N_1579,N_769);
or U6822 (N_6822,N_3275,N_1736);
nor U6823 (N_6823,N_4219,N_2155);
xor U6824 (N_6824,N_3400,N_4085);
and U6825 (N_6825,N_1143,N_3817);
nand U6826 (N_6826,N_2201,N_3239);
or U6827 (N_6827,N_4844,N_3936);
xnor U6828 (N_6828,N_2619,N_4984);
xnor U6829 (N_6829,N_3089,N_4701);
nand U6830 (N_6830,N_4173,N_4300);
and U6831 (N_6831,N_2954,N_938);
and U6832 (N_6832,N_2940,N_2722);
or U6833 (N_6833,N_544,N_3268);
xnor U6834 (N_6834,N_3016,N_4324);
nor U6835 (N_6835,N_927,N_1241);
and U6836 (N_6836,N_468,N_3486);
and U6837 (N_6837,N_1271,N_1755);
nor U6838 (N_6838,N_3958,N_1348);
or U6839 (N_6839,N_1358,N_4328);
nand U6840 (N_6840,N_4276,N_4061);
nand U6841 (N_6841,N_696,N_3744);
or U6842 (N_6842,N_3703,N_3909);
nor U6843 (N_6843,N_4074,N_2279);
xor U6844 (N_6844,N_1438,N_1892);
nand U6845 (N_6845,N_1249,N_4870);
xnor U6846 (N_6846,N_19,N_1622);
nor U6847 (N_6847,N_4639,N_230);
nand U6848 (N_6848,N_3572,N_2538);
nor U6849 (N_6849,N_4986,N_4202);
xnor U6850 (N_6850,N_4422,N_684);
nor U6851 (N_6851,N_3866,N_3346);
or U6852 (N_6852,N_2693,N_1466);
nor U6853 (N_6853,N_549,N_2071);
nand U6854 (N_6854,N_3896,N_3482);
nor U6855 (N_6855,N_3915,N_2993);
xor U6856 (N_6856,N_1468,N_288);
nor U6857 (N_6857,N_1670,N_3611);
nor U6858 (N_6858,N_529,N_1883);
nor U6859 (N_6859,N_2003,N_3551);
xnor U6860 (N_6860,N_2544,N_3261);
nand U6861 (N_6861,N_2471,N_1537);
nand U6862 (N_6862,N_4653,N_3719);
nand U6863 (N_6863,N_1760,N_687);
xnor U6864 (N_6864,N_2658,N_4274);
xor U6865 (N_6865,N_3399,N_4526);
nor U6866 (N_6866,N_1696,N_3548);
nand U6867 (N_6867,N_1620,N_3804);
nor U6868 (N_6868,N_1170,N_716);
nand U6869 (N_6869,N_552,N_4124);
nand U6870 (N_6870,N_4513,N_287);
nor U6871 (N_6871,N_3417,N_3922);
and U6872 (N_6872,N_2599,N_1439);
xnor U6873 (N_6873,N_2199,N_3945);
and U6874 (N_6874,N_990,N_3856);
and U6875 (N_6875,N_657,N_4428);
nor U6876 (N_6876,N_820,N_2026);
nor U6877 (N_6877,N_3496,N_2914);
or U6878 (N_6878,N_1873,N_2766);
nand U6879 (N_6879,N_4311,N_2637);
nor U6880 (N_6880,N_4278,N_3194);
xnor U6881 (N_6881,N_1383,N_390);
nor U6882 (N_6882,N_251,N_1695);
and U6883 (N_6883,N_3380,N_485);
and U6884 (N_6884,N_84,N_1094);
and U6885 (N_6885,N_721,N_614);
or U6886 (N_6886,N_2565,N_2707);
or U6887 (N_6887,N_1314,N_639);
or U6888 (N_6888,N_1259,N_1738);
or U6889 (N_6889,N_1936,N_1216);
or U6890 (N_6890,N_994,N_3231);
or U6891 (N_6891,N_1406,N_4781);
and U6892 (N_6892,N_3801,N_2905);
and U6893 (N_6893,N_13,N_2742);
nor U6894 (N_6894,N_2925,N_3545);
or U6895 (N_6895,N_3331,N_744);
or U6896 (N_6896,N_2042,N_3895);
nand U6897 (N_6897,N_603,N_547);
and U6898 (N_6898,N_4163,N_886);
nand U6899 (N_6899,N_1315,N_363);
or U6900 (N_6900,N_3222,N_2632);
or U6901 (N_6901,N_1219,N_1191);
nand U6902 (N_6902,N_4822,N_2381);
or U6903 (N_6903,N_3780,N_1304);
nand U6904 (N_6904,N_958,N_2988);
nand U6905 (N_6905,N_4368,N_25);
nand U6906 (N_6906,N_3201,N_2810);
and U6907 (N_6907,N_53,N_959);
and U6908 (N_6908,N_371,N_1397);
xor U6909 (N_6909,N_193,N_221);
nand U6910 (N_6910,N_1251,N_3546);
or U6911 (N_6911,N_548,N_4411);
nor U6912 (N_6912,N_2448,N_4314);
and U6913 (N_6913,N_826,N_153);
or U6914 (N_6914,N_2295,N_4557);
nand U6915 (N_6915,N_4879,N_3691);
or U6916 (N_6916,N_1342,N_3651);
and U6917 (N_6917,N_1613,N_3756);
nor U6918 (N_6918,N_3248,N_4209);
nor U6919 (N_6919,N_2352,N_3671);
xor U6920 (N_6920,N_4269,N_550);
nand U6921 (N_6921,N_2694,N_1026);
nor U6922 (N_6922,N_247,N_3269);
nand U6923 (N_6923,N_2185,N_104);
nand U6924 (N_6924,N_3644,N_3731);
xor U6925 (N_6925,N_1625,N_1442);
nand U6926 (N_6926,N_4906,N_2351);
and U6927 (N_6927,N_3212,N_1262);
xnor U6928 (N_6928,N_3294,N_1532);
nand U6929 (N_6929,N_2453,N_3892);
xor U6930 (N_6930,N_968,N_3312);
nor U6931 (N_6931,N_3512,N_209);
nor U6932 (N_6932,N_340,N_399);
and U6933 (N_6933,N_228,N_3920);
and U6934 (N_6934,N_3032,N_282);
or U6935 (N_6935,N_4381,N_3980);
and U6936 (N_6936,N_861,N_1972);
nor U6937 (N_6937,N_4543,N_3185);
or U6938 (N_6938,N_4731,N_3095);
and U6939 (N_6939,N_4602,N_1096);
nand U6940 (N_6940,N_1668,N_4758);
and U6941 (N_6941,N_414,N_2209);
xor U6942 (N_6942,N_1335,N_3127);
or U6943 (N_6943,N_4225,N_1044);
and U6944 (N_6944,N_4766,N_4604);
xnor U6945 (N_6945,N_4951,N_3471);
or U6946 (N_6946,N_3057,N_3685);
nand U6947 (N_6947,N_2089,N_1451);
and U6948 (N_6948,N_987,N_3473);
nor U6949 (N_6949,N_4041,N_1484);
nor U6950 (N_6950,N_57,N_88);
xnor U6951 (N_6951,N_2452,N_20);
nand U6952 (N_6952,N_3754,N_3884);
nand U6953 (N_6953,N_2734,N_62);
nand U6954 (N_6954,N_898,N_1899);
nand U6955 (N_6955,N_2392,N_2242);
nand U6956 (N_6956,N_1268,N_401);
and U6957 (N_6957,N_4670,N_4038);
and U6958 (N_6958,N_4949,N_4767);
and U6959 (N_6959,N_3132,N_4048);
nor U6960 (N_6960,N_3214,N_1713);
xnor U6961 (N_6961,N_4773,N_1153);
or U6962 (N_6962,N_1849,N_1480);
nand U6963 (N_6963,N_4338,N_644);
xor U6964 (N_6964,N_2713,N_3840);
xnor U6965 (N_6965,N_2792,N_4028);
or U6966 (N_6966,N_380,N_4704);
and U6967 (N_6967,N_2005,N_1215);
xor U6968 (N_6968,N_3393,N_2025);
nand U6969 (N_6969,N_238,N_3160);
and U6970 (N_6970,N_4667,N_3411);
xor U6971 (N_6971,N_3337,N_751);
or U6972 (N_6972,N_2561,N_4567);
or U6973 (N_6973,N_922,N_2823);
nor U6974 (N_6974,N_515,N_3820);
nor U6975 (N_6975,N_1436,N_4110);
nand U6976 (N_6976,N_4612,N_4548);
nor U6977 (N_6977,N_3584,N_658);
and U6978 (N_6978,N_4380,N_967);
nor U6979 (N_6979,N_1389,N_3565);
nand U6980 (N_6980,N_82,N_4302);
nor U6981 (N_6981,N_3123,N_3352);
and U6982 (N_6982,N_115,N_2032);
nor U6983 (N_6983,N_2138,N_575);
nand U6984 (N_6984,N_3535,N_1730);
or U6985 (N_6985,N_322,N_643);
nand U6986 (N_6986,N_3051,N_713);
and U6987 (N_6987,N_4533,N_2303);
nand U6988 (N_6988,N_4036,N_216);
nand U6989 (N_6989,N_3713,N_3282);
or U6990 (N_6990,N_3695,N_3705);
or U6991 (N_6991,N_3316,N_1496);
and U6992 (N_6992,N_2253,N_2975);
nor U6993 (N_6993,N_2067,N_3371);
xnor U6994 (N_6994,N_4655,N_1403);
nand U6995 (N_6995,N_277,N_4069);
nor U6996 (N_6996,N_3501,N_2971);
or U6997 (N_6997,N_2704,N_1373);
or U6998 (N_6998,N_1965,N_2604);
nor U6999 (N_6999,N_1431,N_2682);
nor U7000 (N_7000,N_1203,N_477);
nor U7001 (N_7001,N_2534,N_3562);
nor U7002 (N_7002,N_2596,N_3870);
nor U7003 (N_7003,N_4705,N_453);
xor U7004 (N_7004,N_2130,N_3004);
and U7005 (N_7005,N_1097,N_1960);
or U7006 (N_7006,N_1047,N_4605);
and U7007 (N_7007,N_2981,N_979);
nand U7008 (N_7008,N_2464,N_1589);
xor U7009 (N_7009,N_110,N_3539);
or U7010 (N_7010,N_3088,N_1433);
or U7011 (N_7011,N_432,N_3045);
and U7012 (N_7012,N_901,N_3786);
and U7013 (N_7013,N_2477,N_1144);
nand U7014 (N_7014,N_2229,N_4900);
and U7015 (N_7015,N_1202,N_109);
or U7016 (N_7016,N_3198,N_2513);
nor U7017 (N_7017,N_1813,N_2964);
or U7018 (N_7018,N_2105,N_4207);
nor U7019 (N_7019,N_3335,N_1359);
nand U7020 (N_7020,N_3182,N_3197);
or U7021 (N_7021,N_1842,N_3837);
nand U7022 (N_7022,N_2237,N_4957);
nand U7023 (N_7023,N_1270,N_169);
nor U7024 (N_7024,N_3444,N_3429);
xnor U7025 (N_7025,N_2459,N_1483);
nand U7026 (N_7026,N_3436,N_2655);
nand U7027 (N_7027,N_1762,N_3296);
and U7028 (N_7028,N_4510,N_4628);
nor U7029 (N_7029,N_4696,N_4736);
nand U7030 (N_7030,N_4126,N_1473);
nand U7031 (N_7031,N_4472,N_4362);
nor U7032 (N_7032,N_389,N_2892);
nor U7033 (N_7033,N_4500,N_1269);
xnor U7034 (N_7034,N_370,N_3509);
and U7035 (N_7035,N_56,N_298);
nand U7036 (N_7036,N_3526,N_2560);
nor U7037 (N_7037,N_1414,N_3702);
or U7038 (N_7038,N_3682,N_207);
and U7039 (N_7039,N_1492,N_382);
nand U7040 (N_7040,N_2741,N_1699);
or U7041 (N_7041,N_4674,N_1033);
and U7042 (N_7042,N_2231,N_3538);
and U7043 (N_7043,N_3114,N_4937);
and U7044 (N_7044,N_3645,N_961);
or U7045 (N_7045,N_4700,N_4509);
nor U7046 (N_7046,N_3396,N_4671);
and U7047 (N_7047,N_449,N_2222);
nand U7048 (N_7048,N_1000,N_297);
xnor U7049 (N_7049,N_4010,N_3555);
xnor U7050 (N_7050,N_2082,N_4676);
xor U7051 (N_7051,N_224,N_2793);
or U7052 (N_7052,N_4355,N_2769);
nor U7053 (N_7053,N_2018,N_2563);
xnor U7054 (N_7054,N_2091,N_4695);
and U7055 (N_7055,N_781,N_1459);
and U7056 (N_7056,N_3186,N_2309);
nand U7057 (N_7057,N_3323,N_2);
xor U7058 (N_7058,N_3419,N_2781);
xnor U7059 (N_7059,N_2187,N_344);
xnor U7060 (N_7060,N_1244,N_3409);
nand U7061 (N_7061,N_2406,N_1594);
nor U7062 (N_7062,N_514,N_4357);
or U7063 (N_7063,N_3260,N_4545);
and U7064 (N_7064,N_984,N_1706);
nor U7065 (N_7065,N_1247,N_4364);
nand U7066 (N_7066,N_3711,N_2294);
or U7067 (N_7067,N_4867,N_2440);
or U7068 (N_7068,N_1603,N_273);
and U7069 (N_7069,N_4585,N_2593);
or U7070 (N_7070,N_3534,N_2626);
or U7071 (N_7071,N_3632,N_516);
and U7072 (N_7072,N_4969,N_92);
or U7073 (N_7073,N_969,N_2437);
nor U7074 (N_7074,N_1990,N_2852);
nand U7075 (N_7075,N_1938,N_4895);
xnor U7076 (N_7076,N_1602,N_1912);
nor U7077 (N_7077,N_3440,N_4436);
or U7078 (N_7078,N_419,N_1003);
or U7079 (N_7079,N_194,N_2014);
nand U7080 (N_7080,N_562,N_4453);
or U7081 (N_7081,N_2204,N_2474);
nand U7082 (N_7082,N_2401,N_2043);
or U7083 (N_7083,N_3787,N_1092);
nor U7084 (N_7084,N_1664,N_2897);
nand U7085 (N_7085,N_3017,N_1546);
or U7086 (N_7086,N_4228,N_3180);
xnor U7087 (N_7087,N_4008,N_925);
xor U7088 (N_7088,N_1010,N_4488);
nor U7089 (N_7089,N_1550,N_1728);
or U7090 (N_7090,N_3205,N_3607);
xor U7091 (N_7091,N_3297,N_952);
or U7092 (N_7092,N_4899,N_1022);
xor U7093 (N_7093,N_2612,N_218);
nand U7094 (N_7094,N_1686,N_1667);
nand U7095 (N_7095,N_2953,N_1416);
nand U7096 (N_7096,N_1884,N_829);
xor U7097 (N_7097,N_1382,N_2690);
and U7098 (N_7098,N_759,N_3542);
and U7099 (N_7099,N_4650,N_704);
xnor U7100 (N_7100,N_2881,N_2260);
nor U7101 (N_7101,N_2791,N_1081);
xor U7102 (N_7102,N_189,N_1648);
xnor U7103 (N_7103,N_667,N_213);
nor U7104 (N_7104,N_4330,N_3854);
xnor U7105 (N_7105,N_2895,N_797);
or U7106 (N_7106,N_3851,N_308);
nand U7107 (N_7107,N_257,N_2367);
xnor U7108 (N_7108,N_2385,N_2867);
nor U7109 (N_7109,N_3834,N_3199);
nor U7110 (N_7110,N_558,N_290);
xor U7111 (N_7111,N_3850,N_587);
or U7112 (N_7112,N_2760,N_791);
or U7113 (N_7113,N_4005,N_4443);
xor U7114 (N_7114,N_1413,N_4531);
xor U7115 (N_7115,N_1211,N_1747);
xor U7116 (N_7116,N_1169,N_3029);
nor U7117 (N_7117,N_2909,N_3860);
xnor U7118 (N_7118,N_2345,N_866);
or U7119 (N_7119,N_822,N_3629);
or U7120 (N_7120,N_1337,N_1504);
nand U7121 (N_7121,N_2737,N_2432);
and U7122 (N_7122,N_2714,N_999);
and U7123 (N_7123,N_3742,N_518);
xor U7124 (N_7124,N_3843,N_155);
or U7125 (N_7125,N_2191,N_2358);
and U7126 (N_7126,N_4326,N_3351);
and U7127 (N_7127,N_1595,N_159);
and U7128 (N_7128,N_2644,N_267);
nand U7129 (N_7129,N_1018,N_470);
nand U7130 (N_7130,N_3768,N_2436);
nand U7131 (N_7131,N_2885,N_106);
or U7132 (N_7132,N_3005,N_1691);
nand U7133 (N_7133,N_301,N_2165);
xnor U7134 (N_7134,N_1964,N_1866);
xor U7135 (N_7135,N_3190,N_4224);
nand U7136 (N_7136,N_3707,N_2344);
nor U7137 (N_7137,N_3588,N_3072);
nor U7138 (N_7138,N_4285,N_3404);
xnor U7139 (N_7139,N_4113,N_1467);
xor U7140 (N_7140,N_1236,N_535);
or U7141 (N_7141,N_1519,N_3355);
or U7142 (N_7142,N_4242,N_1927);
nand U7143 (N_7143,N_4966,N_1941);
or U7144 (N_7144,N_2297,N_4233);
and U7145 (N_7145,N_1239,N_913);
xnor U7146 (N_7146,N_3365,N_784);
nor U7147 (N_7147,N_4388,N_4345);
xor U7148 (N_7148,N_601,N_965);
nand U7149 (N_7149,N_455,N_2083);
nor U7150 (N_7150,N_4375,N_3558);
and U7151 (N_7151,N_3389,N_2485);
and U7152 (N_7152,N_4192,N_4683);
or U7153 (N_7153,N_3037,N_4574);
or U7154 (N_7154,N_2177,N_3290);
nand U7155 (N_7155,N_2426,N_3416);
xnor U7156 (N_7156,N_2029,N_500);
xor U7157 (N_7157,N_3950,N_1717);
nand U7158 (N_7158,N_2006,N_474);
nor U7159 (N_7159,N_650,N_2463);
nand U7160 (N_7160,N_131,N_2893);
or U7161 (N_7161,N_1321,N_249);
nand U7162 (N_7162,N_4834,N_726);
xnor U7163 (N_7163,N_1994,N_869);
nor U7164 (N_7164,N_1287,N_2672);
nor U7165 (N_7165,N_436,N_2545);
nand U7166 (N_7166,N_232,N_2172);
nor U7167 (N_7167,N_4145,N_578);
or U7168 (N_7168,N_484,N_1539);
or U7169 (N_7169,N_4974,N_2916);
xor U7170 (N_7170,N_391,N_1020);
xor U7171 (N_7171,N_3649,N_2835);
xor U7172 (N_7172,N_4096,N_1631);
nand U7173 (N_7173,N_4288,N_1495);
or U7174 (N_7174,N_686,N_2720);
nand U7175 (N_7175,N_44,N_2350);
nand U7176 (N_7176,N_3701,N_4232);
nand U7177 (N_7177,N_4828,N_1155);
nor U7178 (N_7178,N_2510,N_3391);
and U7179 (N_7179,N_2950,N_3470);
nor U7180 (N_7180,N_3739,N_1528);
xor U7181 (N_7181,N_1109,N_121);
and U7182 (N_7182,N_2961,N_3989);
xnor U7183 (N_7183,N_1767,N_4535);
and U7184 (N_7184,N_2990,N_2504);
and U7185 (N_7185,N_4104,N_4400);
and U7186 (N_7186,N_2641,N_4808);
xor U7187 (N_7187,N_1395,N_307);
xnor U7188 (N_7188,N_3957,N_3823);
xnor U7189 (N_7189,N_733,N_2662);
or U7190 (N_7190,N_2493,N_4114);
xnor U7191 (N_7191,N_1663,N_1334);
nand U7192 (N_7192,N_4001,N_4222);
nor U7193 (N_7193,N_2355,N_2876);
and U7194 (N_7194,N_17,N_3492);
nand U7195 (N_7195,N_3621,N_3536);
xor U7196 (N_7196,N_707,N_1428);
or U7197 (N_7197,N_410,N_2788);
nand U7198 (N_7198,N_3327,N_4857);
and U7199 (N_7199,N_900,N_2332);
and U7200 (N_7200,N_2671,N_478);
and U7201 (N_7201,N_4058,N_1434);
and U7202 (N_7202,N_4034,N_946);
and U7203 (N_7203,N_4190,N_617);
xor U7204 (N_7204,N_1027,N_4972);
xnor U7205 (N_7205,N_896,N_808);
xnor U7206 (N_7206,N_4527,N_1623);
and U7207 (N_7207,N_3481,N_403);
nor U7208 (N_7208,N_171,N_3846);
nand U7209 (N_7209,N_116,N_2248);
or U7210 (N_7210,N_1910,N_3044);
xnor U7211 (N_7211,N_2125,N_1177);
nand U7212 (N_7212,N_496,N_1679);
and U7213 (N_7213,N_3278,N_765);
xor U7214 (N_7214,N_2235,N_930);
nor U7215 (N_7215,N_2745,N_2163);
xnor U7216 (N_7216,N_3028,N_3115);
or U7217 (N_7217,N_2977,N_4726);
nor U7218 (N_7218,N_1075,N_29);
nand U7219 (N_7219,N_3932,N_3406);
and U7220 (N_7220,N_872,N_2944);
and U7221 (N_7221,N_3574,N_2496);
xor U7222 (N_7222,N_2911,N_1165);
or U7223 (N_7223,N_887,N_3627);
xnor U7224 (N_7224,N_1832,N_1341);
and U7225 (N_7225,N_123,N_3487);
xor U7226 (N_7226,N_3869,N_1590);
or U7227 (N_7227,N_2711,N_2589);
or U7228 (N_7228,N_2567,N_254);
nor U7229 (N_7229,N_972,N_2556);
nor U7230 (N_7230,N_48,N_976);
or U7231 (N_7231,N_2891,N_3093);
or U7232 (N_7232,N_1218,N_2601);
or U7233 (N_7233,N_3994,N_2331);
xnor U7234 (N_7234,N_1518,N_1915);
nand U7235 (N_7235,N_4546,N_4652);
xor U7236 (N_7236,N_4530,N_4496);
and U7237 (N_7237,N_4816,N_3635);
and U7238 (N_7238,N_306,N_339);
and U7239 (N_7239,N_2642,N_3792);
or U7240 (N_7240,N_3064,N_486);
xnor U7241 (N_7241,N_1642,N_270);
nand U7242 (N_7242,N_2875,N_1820);
nand U7243 (N_7243,N_811,N_1567);
nand U7244 (N_7244,N_753,N_989);
nor U7245 (N_7245,N_1900,N_2013);
nand U7246 (N_7246,N_1276,N_1605);
or U7247 (N_7247,N_2188,N_4172);
nor U7248 (N_7248,N_4360,N_2689);
or U7249 (N_7249,N_2390,N_883);
xor U7250 (N_7250,N_2646,N_3092);
xnor U7251 (N_7251,N_1078,N_655);
and U7252 (N_7252,N_4504,N_4168);
xor U7253 (N_7253,N_4998,N_1641);
xnor U7254 (N_7254,N_4692,N_741);
xor U7255 (N_7255,N_2141,N_3213);
or U7256 (N_7256,N_1171,N_3971);
or U7257 (N_7257,N_1658,N_258);
xor U7258 (N_7258,N_635,N_2516);
xnor U7259 (N_7259,N_489,N_3829);
nand U7260 (N_7260,N_2254,N_1754);
xor U7261 (N_7261,N_1306,N_2347);
xnor U7262 (N_7262,N_1481,N_2023);
or U7263 (N_7263,N_3788,N_3560);
nand U7264 (N_7264,N_816,N_3024);
xor U7265 (N_7265,N_3646,N_4187);
xnor U7266 (N_7266,N_1982,N_3196);
or U7267 (N_7267,N_3254,N_2335);
nor U7268 (N_7268,N_2859,N_1649);
xor U7269 (N_7269,N_1454,N_1655);
or U7270 (N_7270,N_3570,N_1967);
and U7271 (N_7271,N_2121,N_3427);
and U7272 (N_7272,N_3873,N_4597);
xnor U7273 (N_7273,N_1163,N_637);
or U7274 (N_7274,N_4741,N_926);
nor U7275 (N_7275,N_3762,N_3174);
and U7276 (N_7276,N_3513,N_200);
xor U7277 (N_7277,N_3019,N_3593);
nand U7278 (N_7278,N_3235,N_1950);
nor U7279 (N_7279,N_3489,N_2829);
nand U7280 (N_7280,N_3959,N_3527);
xor U7281 (N_7281,N_2223,N_4176);
and U7282 (N_7282,N_1793,N_1409);
or U7283 (N_7283,N_241,N_827);
nor U7284 (N_7284,N_71,N_2937);
nor U7285 (N_7285,N_1072,N_3624);
nand U7286 (N_7286,N_1277,N_865);
and U7287 (N_7287,N_4138,N_3944);
nand U7288 (N_7288,N_3467,N_2409);
nand U7289 (N_7289,N_788,N_3423);
or U7290 (N_7290,N_1979,N_997);
and U7291 (N_7291,N_3295,N_4408);
nand U7292 (N_7292,N_462,N_1830);
xor U7293 (N_7293,N_3128,N_1354);
nand U7294 (N_7294,N_1346,N_1111);
xor U7295 (N_7295,N_1800,N_212);
nand U7296 (N_7296,N_354,N_599);
nand U7297 (N_7297,N_1345,N_3664);
or U7298 (N_7298,N_800,N_763);
or U7299 (N_7299,N_4930,N_30);
or U7300 (N_7300,N_4800,N_4556);
and U7301 (N_7301,N_476,N_4475);
or U7302 (N_7302,N_3302,N_4833);
xor U7303 (N_7303,N_1488,N_4376);
xor U7304 (N_7304,N_4297,N_823);
xnor U7305 (N_7305,N_26,N_813);
xor U7306 (N_7306,N_2583,N_4429);
xnor U7307 (N_7307,N_2958,N_1088);
nand U7308 (N_7308,N_2447,N_4675);
or U7309 (N_7309,N_4323,N_1645);
or U7310 (N_7310,N_151,N_736);
xnor U7311 (N_7311,N_1558,N_1235);
or U7312 (N_7312,N_847,N_4032);
nor U7313 (N_7313,N_2045,N_4589);
xor U7314 (N_7314,N_3433,N_2277);
nor U7315 (N_7315,N_3076,N_4003);
xnor U7316 (N_7316,N_1752,N_4922);
and U7317 (N_7317,N_2090,N_4880);
xor U7318 (N_7318,N_2078,N_3954);
xnor U7319 (N_7319,N_1571,N_124);
xnor U7320 (N_7320,N_1238,N_1449);
and U7321 (N_7321,N_3175,N_4820);
xnor U7322 (N_7322,N_465,N_3398);
xor U7323 (N_7323,N_1059,N_3381);
nand U7324 (N_7324,N_674,N_4856);
and U7325 (N_7325,N_1399,N_4812);
nand U7326 (N_7326,N_2469,N_4284);
xnor U7327 (N_7327,N_1719,N_2312);
nor U7328 (N_7328,N_421,N_1610);
nand U7329 (N_7329,N_1114,N_2198);
nand U7330 (N_7330,N_206,N_2267);
nor U7331 (N_7331,N_2443,N_1993);
nor U7332 (N_7332,N_4760,N_4198);
xnor U7333 (N_7333,N_4471,N_3845);
xnor U7334 (N_7334,N_1607,N_1015);
or U7335 (N_7335,N_964,N_3366);
nor U7336 (N_7336,N_3816,N_178);
nor U7337 (N_7337,N_2984,N_1617);
nand U7338 (N_7338,N_3832,N_4968);
nand U7339 (N_7339,N_4402,N_1586);
and U7340 (N_7340,N_4481,N_3321);
nand U7341 (N_7341,N_2181,N_1973);
xor U7342 (N_7342,N_1870,N_437);
nand U7343 (N_7343,N_345,N_2421);
nor U7344 (N_7344,N_4887,N_77);
nor U7345 (N_7345,N_749,N_2853);
nor U7346 (N_7346,N_3800,N_1909);
or U7347 (N_7347,N_619,N_3863);
or U7348 (N_7348,N_2832,N_3597);
nand U7349 (N_7349,N_132,N_4039);
nor U7350 (N_7350,N_583,N_1803);
nand U7351 (N_7351,N_702,N_2422);
nor U7352 (N_7352,N_727,N_1014);
and U7353 (N_7353,N_2052,N_888);
or U7354 (N_7354,N_1513,N_1791);
or U7355 (N_7355,N_4340,N_3179);
nand U7356 (N_7356,N_3330,N_909);
xnor U7357 (N_7357,N_3887,N_2086);
nand U7358 (N_7358,N_3600,N_4837);
xor U7359 (N_7359,N_1895,N_1629);
xnor U7360 (N_7360,N_557,N_2112);
nand U7361 (N_7361,N_461,N_3844);
nand U7362 (N_7362,N_2259,N_3490);
nand U7363 (N_7363,N_2101,N_4668);
nor U7364 (N_7364,N_2634,N_683);
or U7365 (N_7365,N_2158,N_299);
or U7366 (N_7366,N_783,N_1599);
nand U7367 (N_7367,N_4154,N_1769);
and U7368 (N_7368,N_305,N_588);
xor U7369 (N_7369,N_3736,N_1711);
nor U7370 (N_7370,N_4397,N_584);
nand U7371 (N_7371,N_2546,N_834);
nand U7372 (N_7372,N_970,N_624);
or U7373 (N_7373,N_2354,N_1178);
nor U7374 (N_7374,N_3667,N_466);
xnor U7375 (N_7375,N_2418,N_3387);
or U7376 (N_7376,N_2888,N_3110);
or U7377 (N_7377,N_4262,N_4432);
nor U7378 (N_7378,N_1823,N_825);
and U7379 (N_7379,N_2106,N_3000);
nand U7380 (N_7380,N_4410,N_546);
xnor U7381 (N_7381,N_174,N_1829);
nor U7382 (N_7382,N_3814,N_4257);
xnor U7383 (N_7383,N_3258,N_4043);
xor U7384 (N_7384,N_2186,N_2336);
or U7385 (N_7385,N_3813,N_2860);
nor U7386 (N_7386,N_3516,N_78);
nor U7387 (N_7387,N_1878,N_12);
xnor U7388 (N_7388,N_1206,N_3745);
and U7389 (N_7389,N_4100,N_4035);
or U7390 (N_7390,N_709,N_2865);
and U7391 (N_7391,N_3499,N_4560);
nand U7392 (N_7392,N_1865,N_3314);
and U7393 (N_7393,N_4938,N_1472);
or U7394 (N_7394,N_1943,N_3907);
nand U7395 (N_7395,N_167,N_338);
and U7396 (N_7396,N_4268,N_4);
or U7397 (N_7397,N_4072,N_3279);
xor U7398 (N_7398,N_4220,N_600);
and U7399 (N_7399,N_539,N_908);
xor U7400 (N_7400,N_3049,N_3116);
nor U7401 (N_7401,N_3229,N_3694);
and U7402 (N_7402,N_2263,N_1172);
xnor U7403 (N_7403,N_2718,N_1101);
nand U7404 (N_7404,N_1845,N_4229);
and U7405 (N_7405,N_1588,N_1242);
and U7406 (N_7406,N_2161,N_4883);
and U7407 (N_7407,N_1444,N_4564);
nand U7408 (N_7408,N_3277,N_2202);
and U7409 (N_7409,N_857,N_2212);
nor U7410 (N_7410,N_1928,N_1797);
nor U7411 (N_7411,N_337,N_4525);
and U7412 (N_7412,N_2273,N_4688);
nor U7413 (N_7413,N_361,N_296);
nor U7414 (N_7414,N_1684,N_2858);
nand U7415 (N_7415,N_4575,N_3874);
nor U7416 (N_7416,N_1460,N_2602);
xnor U7417 (N_7417,N_190,N_3894);
xnor U7418 (N_7418,N_4386,N_1542);
nand U7419 (N_7419,N_2902,N_58);
nand U7420 (N_7420,N_4673,N_1469);
xor U7421 (N_7421,N_1376,N_1854);
and U7422 (N_7422,N_3262,N_3761);
or U7423 (N_7423,N_1274,N_581);
or U7424 (N_7424,N_61,N_2059);
or U7425 (N_7425,N_4128,N_4444);
or U7426 (N_7426,N_272,N_1582);
xnor U7427 (N_7427,N_3428,N_1116);
xor U7428 (N_7428,N_3857,N_1105);
xnor U7429 (N_7429,N_125,N_2264);
and U7430 (N_7430,N_4405,N_2405);
nand U7431 (N_7431,N_4943,N_1763);
and U7432 (N_7432,N_1601,N_4926);
nor U7433 (N_7433,N_4312,N_1952);
xor U7434 (N_7434,N_1502,N_1288);
and U7435 (N_7435,N_1522,N_4413);
or U7436 (N_7436,N_2910,N_1043);
xnor U7437 (N_7437,N_565,N_1369);
and U7438 (N_7438,N_2736,N_4845);
and U7439 (N_7439,N_1520,N_1827);
xor U7440 (N_7440,N_429,N_284);
and U7441 (N_7441,N_954,N_4298);
xnor U7442 (N_7442,N_96,N_4669);
nor U7443 (N_7443,N_4619,N_2579);
xor U7444 (N_7444,N_1237,N_4824);
nor U7445 (N_7445,N_3987,N_4561);
and U7446 (N_7446,N_4896,N_1773);
nor U7447 (N_7447,N_2959,N_1497);
nand U7448 (N_7448,N_902,N_1838);
and U7449 (N_7449,N_942,N_1226);
nor U7450 (N_7450,N_3483,N_2391);
nand U7451 (N_7451,N_2518,N_31);
or U7452 (N_7452,N_4491,N_1204);
or U7453 (N_7453,N_906,N_2225);
nand U7454 (N_7454,N_3124,N_3946);
nor U7455 (N_7455,N_1959,N_4448);
nand U7456 (N_7456,N_4855,N_3881);
or U7457 (N_7457,N_2021,N_915);
and U7458 (N_7458,N_1997,N_2904);
nor U7459 (N_7459,N_1948,N_4333);
xor U7460 (N_7460,N_39,N_4768);
nor U7461 (N_7461,N_4821,N_4846);
nand U7462 (N_7462,N_2291,N_4863);
nor U7463 (N_7463,N_1721,N_1887);
nand U7464 (N_7464,N_3564,N_2554);
and U7465 (N_7465,N_1669,N_1665);
nor U7466 (N_7466,N_1212,N_3310);
or U7467 (N_7467,N_4175,N_2363);
xnor U7468 (N_7468,N_4280,N_4307);
and U7469 (N_7469,N_4524,N_4607);
xnor U7470 (N_7470,N_2232,N_3137);
or U7471 (N_7471,N_3529,N_3151);
nor U7472 (N_7472,N_1394,N_355);
nor U7473 (N_7473,N_3052,N_4776);
xnor U7474 (N_7474,N_4248,N_1771);
xor U7475 (N_7475,N_832,N_512);
xor U7476 (N_7476,N_4469,N_1671);
nand U7477 (N_7477,N_2533,N_2216);
xnor U7478 (N_7478,N_2475,N_4729);
nand U7479 (N_7479,N_1136,N_2797);
xor U7480 (N_7480,N_2869,N_1801);
xor U7481 (N_7481,N_1411,N_2156);
nand U7482 (N_7482,N_3822,N_817);
nor U7483 (N_7483,N_803,N_2878);
nor U7484 (N_7484,N_4959,N_2280);
nor U7485 (N_7485,N_192,N_2157);
xnor U7486 (N_7486,N_3066,N_2274);
and U7487 (N_7487,N_3634,N_2864);
nor U7488 (N_7488,N_1896,N_1758);
xor U7489 (N_7489,N_4282,N_2055);
and U7490 (N_7490,N_4325,N_3206);
and U7491 (N_7491,N_3336,N_3392);
and U7492 (N_7492,N_142,N_2054);
nand U7493 (N_7493,N_3441,N_4461);
nor U7494 (N_7494,N_37,N_3809);
nand U7495 (N_7495,N_4573,N_2088);
nor U7496 (N_7496,N_1099,N_2095);
xnor U7497 (N_7497,N_750,N_3699);
xnor U7498 (N_7498,N_4158,N_4438);
xnor U7499 (N_7499,N_3223,N_941);
nand U7500 (N_7500,N_4848,N_2593);
and U7501 (N_7501,N_3199,N_2237);
xor U7502 (N_7502,N_681,N_4316);
nor U7503 (N_7503,N_1305,N_411);
nor U7504 (N_7504,N_1214,N_1051);
and U7505 (N_7505,N_606,N_4810);
and U7506 (N_7506,N_4152,N_599);
nor U7507 (N_7507,N_1550,N_1389);
nor U7508 (N_7508,N_375,N_666);
nor U7509 (N_7509,N_3620,N_422);
nor U7510 (N_7510,N_388,N_2684);
nor U7511 (N_7511,N_1594,N_936);
nor U7512 (N_7512,N_1563,N_4238);
or U7513 (N_7513,N_4540,N_4155);
nor U7514 (N_7514,N_2182,N_4327);
nand U7515 (N_7515,N_844,N_3074);
nor U7516 (N_7516,N_4722,N_237);
xor U7517 (N_7517,N_4544,N_1504);
or U7518 (N_7518,N_508,N_4596);
nor U7519 (N_7519,N_3743,N_4044);
and U7520 (N_7520,N_2388,N_4761);
xnor U7521 (N_7521,N_4243,N_223);
nor U7522 (N_7522,N_898,N_4949);
and U7523 (N_7523,N_3649,N_1811);
and U7524 (N_7524,N_122,N_2631);
and U7525 (N_7525,N_3041,N_3096);
nand U7526 (N_7526,N_3743,N_889);
nor U7527 (N_7527,N_4414,N_2750);
and U7528 (N_7528,N_1561,N_2569);
or U7529 (N_7529,N_1201,N_245);
xnor U7530 (N_7530,N_3932,N_3588);
nor U7531 (N_7531,N_1914,N_1442);
or U7532 (N_7532,N_4061,N_4187);
nor U7533 (N_7533,N_4819,N_4743);
and U7534 (N_7534,N_906,N_1719);
and U7535 (N_7535,N_187,N_4697);
and U7536 (N_7536,N_3877,N_3120);
and U7537 (N_7537,N_1081,N_401);
and U7538 (N_7538,N_2190,N_216);
nand U7539 (N_7539,N_2657,N_2862);
xnor U7540 (N_7540,N_1038,N_2824);
nor U7541 (N_7541,N_2692,N_1786);
nand U7542 (N_7542,N_2961,N_679);
xnor U7543 (N_7543,N_4730,N_3809);
nor U7544 (N_7544,N_2863,N_477);
nor U7545 (N_7545,N_1313,N_1013);
xor U7546 (N_7546,N_2824,N_3204);
or U7547 (N_7547,N_3651,N_1259);
nand U7548 (N_7548,N_4097,N_3698);
xnor U7549 (N_7549,N_4696,N_2309);
or U7550 (N_7550,N_2091,N_2439);
and U7551 (N_7551,N_4332,N_3151);
nand U7552 (N_7552,N_3621,N_3490);
xnor U7553 (N_7553,N_2017,N_1747);
and U7554 (N_7554,N_3081,N_3060);
nor U7555 (N_7555,N_898,N_1275);
and U7556 (N_7556,N_3204,N_2739);
nand U7557 (N_7557,N_4562,N_1903);
and U7558 (N_7558,N_3351,N_4133);
xnor U7559 (N_7559,N_1910,N_2078);
nand U7560 (N_7560,N_2319,N_2618);
nand U7561 (N_7561,N_4649,N_1785);
nand U7562 (N_7562,N_4468,N_3877);
nand U7563 (N_7563,N_3157,N_1133);
xor U7564 (N_7564,N_18,N_57);
xnor U7565 (N_7565,N_2591,N_1214);
xor U7566 (N_7566,N_972,N_780);
and U7567 (N_7567,N_4676,N_3275);
nand U7568 (N_7568,N_3980,N_3294);
xnor U7569 (N_7569,N_4123,N_1325);
nor U7570 (N_7570,N_3292,N_3025);
xor U7571 (N_7571,N_2260,N_4584);
nand U7572 (N_7572,N_1473,N_4164);
or U7573 (N_7573,N_3046,N_165);
and U7574 (N_7574,N_2626,N_4708);
nor U7575 (N_7575,N_4753,N_570);
or U7576 (N_7576,N_1717,N_136);
xnor U7577 (N_7577,N_2020,N_1011);
or U7578 (N_7578,N_2655,N_1183);
nor U7579 (N_7579,N_2137,N_4986);
and U7580 (N_7580,N_1556,N_4375);
xor U7581 (N_7581,N_3264,N_1463);
xnor U7582 (N_7582,N_4942,N_2646);
and U7583 (N_7583,N_1994,N_1683);
nor U7584 (N_7584,N_359,N_586);
or U7585 (N_7585,N_2002,N_2470);
nor U7586 (N_7586,N_2050,N_2240);
nor U7587 (N_7587,N_2038,N_3754);
xor U7588 (N_7588,N_3227,N_3245);
or U7589 (N_7589,N_3474,N_3407);
and U7590 (N_7590,N_3417,N_2694);
or U7591 (N_7591,N_1585,N_1902);
and U7592 (N_7592,N_3816,N_598);
or U7593 (N_7593,N_3824,N_4745);
nor U7594 (N_7594,N_3356,N_110);
xnor U7595 (N_7595,N_3508,N_968);
xnor U7596 (N_7596,N_2834,N_2431);
nand U7597 (N_7597,N_3935,N_4603);
or U7598 (N_7598,N_4691,N_3031);
xnor U7599 (N_7599,N_2731,N_3323);
nor U7600 (N_7600,N_3400,N_4836);
or U7601 (N_7601,N_3329,N_4472);
and U7602 (N_7602,N_2398,N_3806);
nand U7603 (N_7603,N_3582,N_2296);
and U7604 (N_7604,N_487,N_2069);
or U7605 (N_7605,N_2580,N_2997);
xor U7606 (N_7606,N_2729,N_4665);
xnor U7607 (N_7607,N_1347,N_1584);
nor U7608 (N_7608,N_1465,N_4179);
nor U7609 (N_7609,N_3760,N_1992);
and U7610 (N_7610,N_638,N_4429);
and U7611 (N_7611,N_2253,N_3269);
nand U7612 (N_7612,N_2079,N_1469);
xor U7613 (N_7613,N_3279,N_619);
nand U7614 (N_7614,N_4481,N_4747);
nand U7615 (N_7615,N_2899,N_4625);
nand U7616 (N_7616,N_1297,N_4427);
nand U7617 (N_7617,N_1310,N_141);
nand U7618 (N_7618,N_4600,N_1926);
nor U7619 (N_7619,N_154,N_2968);
xnor U7620 (N_7620,N_1903,N_2792);
and U7621 (N_7621,N_4196,N_4217);
xor U7622 (N_7622,N_4449,N_94);
or U7623 (N_7623,N_2357,N_4822);
or U7624 (N_7624,N_1157,N_2955);
xor U7625 (N_7625,N_2344,N_3197);
or U7626 (N_7626,N_4038,N_2917);
nor U7627 (N_7627,N_4150,N_973);
xnor U7628 (N_7628,N_3697,N_2150);
and U7629 (N_7629,N_3287,N_1050);
xnor U7630 (N_7630,N_624,N_544);
or U7631 (N_7631,N_3697,N_4443);
nand U7632 (N_7632,N_945,N_3079);
nor U7633 (N_7633,N_2798,N_3572);
nor U7634 (N_7634,N_368,N_1147);
nor U7635 (N_7635,N_1039,N_1707);
nor U7636 (N_7636,N_767,N_839);
nor U7637 (N_7637,N_81,N_1965);
or U7638 (N_7638,N_806,N_2500);
nand U7639 (N_7639,N_3737,N_3192);
or U7640 (N_7640,N_2768,N_3671);
nand U7641 (N_7641,N_1060,N_3307);
or U7642 (N_7642,N_993,N_1255);
and U7643 (N_7643,N_762,N_3514);
xnor U7644 (N_7644,N_2839,N_4890);
nand U7645 (N_7645,N_3221,N_1120);
and U7646 (N_7646,N_4536,N_4223);
xnor U7647 (N_7647,N_820,N_454);
and U7648 (N_7648,N_3060,N_3772);
and U7649 (N_7649,N_1749,N_4357);
nor U7650 (N_7650,N_1807,N_2393);
xor U7651 (N_7651,N_3402,N_1323);
nor U7652 (N_7652,N_508,N_2914);
and U7653 (N_7653,N_2424,N_511);
nand U7654 (N_7654,N_782,N_1447);
and U7655 (N_7655,N_3887,N_1729);
nand U7656 (N_7656,N_1545,N_4584);
xor U7657 (N_7657,N_4965,N_136);
nand U7658 (N_7658,N_3303,N_1851);
nand U7659 (N_7659,N_3809,N_1982);
nor U7660 (N_7660,N_92,N_138);
nor U7661 (N_7661,N_3140,N_1398);
nor U7662 (N_7662,N_4299,N_1247);
nor U7663 (N_7663,N_4500,N_894);
xor U7664 (N_7664,N_1357,N_3615);
or U7665 (N_7665,N_1435,N_1045);
xnor U7666 (N_7666,N_3039,N_94);
and U7667 (N_7667,N_2550,N_4125);
nor U7668 (N_7668,N_4607,N_4139);
xor U7669 (N_7669,N_2160,N_3161);
xor U7670 (N_7670,N_3527,N_2495);
nor U7671 (N_7671,N_382,N_1905);
nor U7672 (N_7672,N_102,N_342);
or U7673 (N_7673,N_2303,N_2962);
xnor U7674 (N_7674,N_879,N_2868);
xor U7675 (N_7675,N_847,N_1001);
nor U7676 (N_7676,N_2031,N_3971);
nand U7677 (N_7677,N_1438,N_3209);
xor U7678 (N_7678,N_2519,N_3439);
xnor U7679 (N_7679,N_4753,N_3725);
xor U7680 (N_7680,N_3824,N_1725);
nor U7681 (N_7681,N_1494,N_2802);
nand U7682 (N_7682,N_1464,N_142);
nor U7683 (N_7683,N_2963,N_2422);
and U7684 (N_7684,N_4615,N_3799);
and U7685 (N_7685,N_4717,N_4608);
xnor U7686 (N_7686,N_503,N_2340);
nor U7687 (N_7687,N_360,N_4284);
nand U7688 (N_7688,N_2917,N_3579);
or U7689 (N_7689,N_578,N_2902);
xnor U7690 (N_7690,N_4758,N_1723);
or U7691 (N_7691,N_1248,N_2753);
nand U7692 (N_7692,N_2601,N_3158);
xor U7693 (N_7693,N_128,N_194);
nor U7694 (N_7694,N_1610,N_937);
xnor U7695 (N_7695,N_1030,N_1728);
or U7696 (N_7696,N_4401,N_1851);
nand U7697 (N_7697,N_1500,N_36);
or U7698 (N_7698,N_3006,N_3980);
nand U7699 (N_7699,N_2863,N_4399);
nor U7700 (N_7700,N_2750,N_2721);
xor U7701 (N_7701,N_2627,N_4992);
nand U7702 (N_7702,N_3917,N_3735);
xnor U7703 (N_7703,N_1490,N_3471);
nand U7704 (N_7704,N_1070,N_1488);
nor U7705 (N_7705,N_3271,N_432);
xor U7706 (N_7706,N_1860,N_4232);
or U7707 (N_7707,N_4755,N_336);
or U7708 (N_7708,N_3642,N_2284);
or U7709 (N_7709,N_2323,N_1906);
nor U7710 (N_7710,N_2807,N_3541);
or U7711 (N_7711,N_4495,N_3077);
nor U7712 (N_7712,N_1160,N_1905);
and U7713 (N_7713,N_754,N_224);
nand U7714 (N_7714,N_4435,N_1594);
nand U7715 (N_7715,N_2698,N_1599);
nor U7716 (N_7716,N_4197,N_3577);
nor U7717 (N_7717,N_4366,N_2432);
and U7718 (N_7718,N_997,N_1679);
nor U7719 (N_7719,N_3006,N_636);
nor U7720 (N_7720,N_2094,N_1683);
nand U7721 (N_7721,N_2040,N_465);
xnor U7722 (N_7722,N_334,N_3555);
nand U7723 (N_7723,N_4152,N_3122);
and U7724 (N_7724,N_527,N_1798);
xnor U7725 (N_7725,N_1972,N_3356);
or U7726 (N_7726,N_3906,N_1991);
nand U7727 (N_7727,N_1285,N_3030);
or U7728 (N_7728,N_2715,N_4205);
nand U7729 (N_7729,N_2697,N_2044);
nor U7730 (N_7730,N_662,N_2658);
nor U7731 (N_7731,N_1000,N_1804);
or U7732 (N_7732,N_2204,N_4019);
xor U7733 (N_7733,N_2393,N_466);
xnor U7734 (N_7734,N_3635,N_2315);
nand U7735 (N_7735,N_1099,N_1288);
or U7736 (N_7736,N_166,N_167);
or U7737 (N_7737,N_4502,N_3268);
and U7738 (N_7738,N_1771,N_113);
nand U7739 (N_7739,N_3130,N_2815);
or U7740 (N_7740,N_274,N_970);
nor U7741 (N_7741,N_3375,N_1614);
or U7742 (N_7742,N_4215,N_1005);
and U7743 (N_7743,N_1122,N_2121);
nor U7744 (N_7744,N_2489,N_3996);
and U7745 (N_7745,N_3996,N_4511);
nand U7746 (N_7746,N_4484,N_201);
nor U7747 (N_7747,N_4140,N_2769);
or U7748 (N_7748,N_4695,N_448);
xnor U7749 (N_7749,N_2216,N_107);
nor U7750 (N_7750,N_2056,N_601);
xor U7751 (N_7751,N_3439,N_1983);
xor U7752 (N_7752,N_1359,N_2253);
xnor U7753 (N_7753,N_392,N_2755);
nor U7754 (N_7754,N_1195,N_1000);
xor U7755 (N_7755,N_4832,N_3086);
nor U7756 (N_7756,N_3582,N_2229);
nor U7757 (N_7757,N_1446,N_970);
xor U7758 (N_7758,N_2500,N_4816);
xor U7759 (N_7759,N_90,N_1787);
xor U7760 (N_7760,N_77,N_2356);
and U7761 (N_7761,N_4993,N_3359);
xor U7762 (N_7762,N_326,N_2548);
nand U7763 (N_7763,N_2271,N_2528);
nand U7764 (N_7764,N_2692,N_2532);
or U7765 (N_7765,N_2042,N_371);
xnor U7766 (N_7766,N_1670,N_2962);
or U7767 (N_7767,N_400,N_3580);
or U7768 (N_7768,N_1700,N_3761);
nor U7769 (N_7769,N_4917,N_422);
nor U7770 (N_7770,N_2699,N_3038);
xnor U7771 (N_7771,N_665,N_124);
nand U7772 (N_7772,N_2598,N_4896);
and U7773 (N_7773,N_4272,N_2450);
nand U7774 (N_7774,N_4702,N_514);
nand U7775 (N_7775,N_4978,N_2854);
and U7776 (N_7776,N_4250,N_4119);
xor U7777 (N_7777,N_2987,N_2253);
nor U7778 (N_7778,N_332,N_176);
xnor U7779 (N_7779,N_4064,N_2964);
xor U7780 (N_7780,N_3119,N_2910);
nand U7781 (N_7781,N_3706,N_1471);
nand U7782 (N_7782,N_4278,N_520);
nand U7783 (N_7783,N_1316,N_1790);
or U7784 (N_7784,N_838,N_1529);
nand U7785 (N_7785,N_3018,N_2434);
xnor U7786 (N_7786,N_1915,N_1023);
nand U7787 (N_7787,N_53,N_941);
nor U7788 (N_7788,N_1614,N_2433);
or U7789 (N_7789,N_1780,N_1289);
and U7790 (N_7790,N_737,N_3901);
and U7791 (N_7791,N_2390,N_3013);
and U7792 (N_7792,N_3109,N_3516);
and U7793 (N_7793,N_1078,N_3933);
nand U7794 (N_7794,N_2251,N_13);
and U7795 (N_7795,N_4182,N_4920);
xor U7796 (N_7796,N_183,N_67);
xor U7797 (N_7797,N_2183,N_3759);
nor U7798 (N_7798,N_1566,N_1653);
or U7799 (N_7799,N_2124,N_4873);
nor U7800 (N_7800,N_3147,N_3482);
and U7801 (N_7801,N_3371,N_2380);
xor U7802 (N_7802,N_2541,N_4020);
or U7803 (N_7803,N_4181,N_2695);
or U7804 (N_7804,N_2924,N_4138);
nor U7805 (N_7805,N_1057,N_2862);
nand U7806 (N_7806,N_544,N_474);
and U7807 (N_7807,N_3817,N_4500);
xnor U7808 (N_7808,N_2027,N_458);
xor U7809 (N_7809,N_326,N_4477);
nor U7810 (N_7810,N_2181,N_3735);
and U7811 (N_7811,N_4305,N_4039);
nor U7812 (N_7812,N_2737,N_2503);
or U7813 (N_7813,N_4606,N_2678);
and U7814 (N_7814,N_327,N_1810);
nor U7815 (N_7815,N_1499,N_2449);
xnor U7816 (N_7816,N_781,N_684);
nor U7817 (N_7817,N_4555,N_3349);
or U7818 (N_7818,N_3036,N_2074);
and U7819 (N_7819,N_4118,N_2332);
nor U7820 (N_7820,N_569,N_460);
xnor U7821 (N_7821,N_3961,N_3543);
xor U7822 (N_7822,N_1666,N_4627);
or U7823 (N_7823,N_480,N_2057);
or U7824 (N_7824,N_2576,N_387);
or U7825 (N_7825,N_1886,N_4393);
or U7826 (N_7826,N_190,N_4583);
nand U7827 (N_7827,N_1790,N_870);
or U7828 (N_7828,N_4074,N_2278);
nand U7829 (N_7829,N_3787,N_3872);
nand U7830 (N_7830,N_2715,N_330);
nand U7831 (N_7831,N_1225,N_1117);
nor U7832 (N_7832,N_660,N_4045);
or U7833 (N_7833,N_3699,N_1277);
and U7834 (N_7834,N_204,N_1952);
and U7835 (N_7835,N_2902,N_1803);
or U7836 (N_7836,N_2559,N_784);
nand U7837 (N_7837,N_872,N_3407);
nor U7838 (N_7838,N_4271,N_3221);
or U7839 (N_7839,N_1730,N_2946);
nor U7840 (N_7840,N_1831,N_1139);
xor U7841 (N_7841,N_908,N_958);
xor U7842 (N_7842,N_2588,N_1773);
nor U7843 (N_7843,N_2078,N_4219);
and U7844 (N_7844,N_1671,N_369);
nor U7845 (N_7845,N_439,N_2463);
or U7846 (N_7846,N_3966,N_2749);
or U7847 (N_7847,N_4939,N_3684);
xnor U7848 (N_7848,N_2135,N_2927);
nand U7849 (N_7849,N_4753,N_72);
nor U7850 (N_7850,N_2357,N_4039);
or U7851 (N_7851,N_2979,N_2358);
or U7852 (N_7852,N_3734,N_1486);
or U7853 (N_7853,N_3269,N_1694);
and U7854 (N_7854,N_4984,N_4084);
or U7855 (N_7855,N_3717,N_1688);
and U7856 (N_7856,N_1545,N_440);
xor U7857 (N_7857,N_3411,N_3175);
xor U7858 (N_7858,N_4731,N_1218);
nand U7859 (N_7859,N_3178,N_2727);
nor U7860 (N_7860,N_2014,N_3675);
and U7861 (N_7861,N_4531,N_4391);
or U7862 (N_7862,N_3935,N_636);
or U7863 (N_7863,N_4901,N_2997);
nand U7864 (N_7864,N_1638,N_226);
nand U7865 (N_7865,N_2648,N_1033);
nor U7866 (N_7866,N_4956,N_865);
nand U7867 (N_7867,N_1319,N_4611);
xnor U7868 (N_7868,N_179,N_2110);
and U7869 (N_7869,N_4451,N_4301);
and U7870 (N_7870,N_285,N_2535);
and U7871 (N_7871,N_2928,N_854);
nand U7872 (N_7872,N_2661,N_1391);
nor U7873 (N_7873,N_2602,N_32);
nor U7874 (N_7874,N_3194,N_1537);
xnor U7875 (N_7875,N_3826,N_1739);
xor U7876 (N_7876,N_3352,N_3764);
and U7877 (N_7877,N_4560,N_38);
or U7878 (N_7878,N_266,N_1322);
xnor U7879 (N_7879,N_4423,N_3065);
nand U7880 (N_7880,N_4683,N_2660);
nor U7881 (N_7881,N_690,N_2206);
nor U7882 (N_7882,N_914,N_972);
xor U7883 (N_7883,N_2041,N_1003);
nor U7884 (N_7884,N_456,N_503);
or U7885 (N_7885,N_2780,N_1450);
nor U7886 (N_7886,N_4022,N_216);
nor U7887 (N_7887,N_514,N_3622);
nand U7888 (N_7888,N_745,N_1983);
and U7889 (N_7889,N_1349,N_405);
nor U7890 (N_7890,N_4047,N_4071);
xor U7891 (N_7891,N_2106,N_2150);
and U7892 (N_7892,N_2990,N_2037);
xor U7893 (N_7893,N_643,N_3129);
and U7894 (N_7894,N_3793,N_88);
nand U7895 (N_7895,N_2549,N_1139);
or U7896 (N_7896,N_1743,N_523);
nand U7897 (N_7897,N_1030,N_973);
nor U7898 (N_7898,N_3637,N_556);
nor U7899 (N_7899,N_4886,N_3550);
xor U7900 (N_7900,N_2798,N_4490);
xor U7901 (N_7901,N_3496,N_181);
and U7902 (N_7902,N_3137,N_1598);
and U7903 (N_7903,N_296,N_3936);
xnor U7904 (N_7904,N_4394,N_725);
or U7905 (N_7905,N_151,N_2798);
or U7906 (N_7906,N_3582,N_1757);
nor U7907 (N_7907,N_3170,N_122);
nand U7908 (N_7908,N_3337,N_1794);
xnor U7909 (N_7909,N_3559,N_2583);
nor U7910 (N_7910,N_264,N_2072);
xor U7911 (N_7911,N_2079,N_4902);
xor U7912 (N_7912,N_960,N_4249);
nand U7913 (N_7913,N_1559,N_3423);
or U7914 (N_7914,N_727,N_3969);
nor U7915 (N_7915,N_2407,N_3008);
nor U7916 (N_7916,N_348,N_2442);
or U7917 (N_7917,N_71,N_3320);
or U7918 (N_7918,N_4615,N_1287);
and U7919 (N_7919,N_3238,N_2277);
and U7920 (N_7920,N_4296,N_3332);
nor U7921 (N_7921,N_4340,N_4526);
nor U7922 (N_7922,N_679,N_4052);
xor U7923 (N_7923,N_1227,N_3730);
or U7924 (N_7924,N_372,N_2161);
and U7925 (N_7925,N_398,N_4480);
nand U7926 (N_7926,N_451,N_3390);
or U7927 (N_7927,N_1331,N_3012);
xor U7928 (N_7928,N_1905,N_1893);
xnor U7929 (N_7929,N_1755,N_3176);
xor U7930 (N_7930,N_84,N_3221);
or U7931 (N_7931,N_808,N_4558);
and U7932 (N_7932,N_44,N_3773);
nand U7933 (N_7933,N_393,N_3874);
nand U7934 (N_7934,N_3949,N_3853);
and U7935 (N_7935,N_2302,N_381);
xor U7936 (N_7936,N_3389,N_2685);
and U7937 (N_7937,N_4998,N_1193);
xor U7938 (N_7938,N_2519,N_259);
nand U7939 (N_7939,N_2292,N_3662);
nand U7940 (N_7940,N_2768,N_2118);
or U7941 (N_7941,N_4988,N_1747);
xnor U7942 (N_7942,N_2900,N_1579);
or U7943 (N_7943,N_603,N_1282);
nand U7944 (N_7944,N_856,N_4974);
or U7945 (N_7945,N_3173,N_1557);
xnor U7946 (N_7946,N_3044,N_859);
nand U7947 (N_7947,N_2755,N_4253);
and U7948 (N_7948,N_2741,N_1036);
nand U7949 (N_7949,N_1061,N_4993);
nand U7950 (N_7950,N_1182,N_52);
xnor U7951 (N_7951,N_4957,N_446);
nor U7952 (N_7952,N_2014,N_1662);
nand U7953 (N_7953,N_2389,N_4782);
nor U7954 (N_7954,N_3908,N_514);
nand U7955 (N_7955,N_3646,N_4926);
nor U7956 (N_7956,N_3922,N_2787);
or U7957 (N_7957,N_1246,N_3648);
xnor U7958 (N_7958,N_1124,N_4814);
nand U7959 (N_7959,N_3715,N_3228);
xor U7960 (N_7960,N_1681,N_3783);
or U7961 (N_7961,N_3743,N_4249);
and U7962 (N_7962,N_3992,N_3486);
and U7963 (N_7963,N_4785,N_4692);
nor U7964 (N_7964,N_4237,N_568);
nor U7965 (N_7965,N_4256,N_2284);
nor U7966 (N_7966,N_1926,N_1120);
nor U7967 (N_7967,N_4146,N_885);
nand U7968 (N_7968,N_134,N_4076);
xnor U7969 (N_7969,N_4491,N_1074);
xor U7970 (N_7970,N_4810,N_2918);
or U7971 (N_7971,N_2311,N_1295);
and U7972 (N_7972,N_3105,N_2937);
xor U7973 (N_7973,N_2991,N_4199);
nor U7974 (N_7974,N_4250,N_3757);
and U7975 (N_7975,N_1882,N_4281);
nor U7976 (N_7976,N_819,N_622);
or U7977 (N_7977,N_578,N_116);
or U7978 (N_7978,N_4338,N_200);
and U7979 (N_7979,N_3060,N_4559);
and U7980 (N_7980,N_4906,N_1039);
or U7981 (N_7981,N_170,N_3295);
nor U7982 (N_7982,N_1195,N_2745);
xor U7983 (N_7983,N_1628,N_777);
xor U7984 (N_7984,N_4080,N_1514);
or U7985 (N_7985,N_1240,N_4117);
nand U7986 (N_7986,N_2676,N_898);
and U7987 (N_7987,N_2648,N_1778);
nand U7988 (N_7988,N_907,N_1234);
nor U7989 (N_7989,N_3071,N_1749);
or U7990 (N_7990,N_4479,N_1130);
xnor U7991 (N_7991,N_1695,N_3659);
nand U7992 (N_7992,N_4029,N_3713);
xnor U7993 (N_7993,N_3705,N_2897);
or U7994 (N_7994,N_1680,N_4742);
xnor U7995 (N_7995,N_2983,N_1390);
or U7996 (N_7996,N_4610,N_1025);
xnor U7997 (N_7997,N_3779,N_3104);
nor U7998 (N_7998,N_4550,N_2486);
xor U7999 (N_7999,N_2272,N_3792);
nand U8000 (N_8000,N_3110,N_4657);
nor U8001 (N_8001,N_290,N_3399);
and U8002 (N_8002,N_1857,N_1818);
nor U8003 (N_8003,N_134,N_4481);
xor U8004 (N_8004,N_4193,N_4957);
nor U8005 (N_8005,N_1985,N_2819);
or U8006 (N_8006,N_2383,N_4821);
nand U8007 (N_8007,N_3931,N_1290);
or U8008 (N_8008,N_1126,N_1140);
and U8009 (N_8009,N_4344,N_3837);
nand U8010 (N_8010,N_1305,N_3209);
and U8011 (N_8011,N_98,N_311);
and U8012 (N_8012,N_323,N_2993);
nor U8013 (N_8013,N_2063,N_1649);
or U8014 (N_8014,N_156,N_1057);
and U8015 (N_8015,N_2138,N_1728);
nand U8016 (N_8016,N_4789,N_4238);
nor U8017 (N_8017,N_1994,N_3123);
nor U8018 (N_8018,N_3046,N_3889);
nor U8019 (N_8019,N_1775,N_268);
xor U8020 (N_8020,N_1261,N_2657);
or U8021 (N_8021,N_4912,N_3182);
nor U8022 (N_8022,N_2273,N_3012);
xnor U8023 (N_8023,N_989,N_451);
nor U8024 (N_8024,N_3550,N_2929);
nor U8025 (N_8025,N_3585,N_3070);
or U8026 (N_8026,N_2089,N_2973);
nand U8027 (N_8027,N_3325,N_1886);
nand U8028 (N_8028,N_1504,N_4987);
or U8029 (N_8029,N_2620,N_2612);
or U8030 (N_8030,N_2844,N_3613);
nand U8031 (N_8031,N_175,N_3405);
or U8032 (N_8032,N_4729,N_796);
nor U8033 (N_8033,N_76,N_2474);
or U8034 (N_8034,N_112,N_2428);
and U8035 (N_8035,N_2123,N_2770);
xor U8036 (N_8036,N_2200,N_2693);
nand U8037 (N_8037,N_3612,N_4836);
nand U8038 (N_8038,N_4608,N_1840);
nor U8039 (N_8039,N_4087,N_1521);
nand U8040 (N_8040,N_538,N_4695);
and U8041 (N_8041,N_156,N_1901);
and U8042 (N_8042,N_3536,N_487);
and U8043 (N_8043,N_1244,N_4661);
xnor U8044 (N_8044,N_29,N_2869);
and U8045 (N_8045,N_4011,N_2252);
nor U8046 (N_8046,N_3549,N_4882);
nor U8047 (N_8047,N_4752,N_3838);
nor U8048 (N_8048,N_4274,N_4511);
xor U8049 (N_8049,N_2913,N_2242);
xnor U8050 (N_8050,N_3517,N_1442);
nand U8051 (N_8051,N_3464,N_2786);
xnor U8052 (N_8052,N_1355,N_2712);
nor U8053 (N_8053,N_515,N_1833);
and U8054 (N_8054,N_2785,N_1156);
or U8055 (N_8055,N_3800,N_1010);
or U8056 (N_8056,N_4157,N_2971);
xor U8057 (N_8057,N_2461,N_278);
nand U8058 (N_8058,N_317,N_121);
nor U8059 (N_8059,N_4278,N_2318);
xnor U8060 (N_8060,N_407,N_2988);
or U8061 (N_8061,N_2016,N_2236);
and U8062 (N_8062,N_276,N_410);
or U8063 (N_8063,N_2922,N_3936);
or U8064 (N_8064,N_1231,N_1271);
xor U8065 (N_8065,N_333,N_2393);
or U8066 (N_8066,N_2123,N_1334);
and U8067 (N_8067,N_723,N_4353);
nor U8068 (N_8068,N_4720,N_2500);
xor U8069 (N_8069,N_799,N_3355);
nand U8070 (N_8070,N_4959,N_1978);
and U8071 (N_8071,N_2342,N_809);
and U8072 (N_8072,N_1697,N_577);
xnor U8073 (N_8073,N_889,N_920);
xor U8074 (N_8074,N_2194,N_3789);
or U8075 (N_8075,N_76,N_65);
or U8076 (N_8076,N_2393,N_729);
nand U8077 (N_8077,N_4124,N_1745);
and U8078 (N_8078,N_1523,N_4449);
nor U8079 (N_8079,N_1689,N_1572);
nor U8080 (N_8080,N_2082,N_4472);
xor U8081 (N_8081,N_4490,N_485);
nand U8082 (N_8082,N_2858,N_757);
nand U8083 (N_8083,N_3083,N_3598);
xor U8084 (N_8084,N_3579,N_3156);
or U8085 (N_8085,N_4216,N_174);
xor U8086 (N_8086,N_2692,N_2379);
nand U8087 (N_8087,N_589,N_1597);
nand U8088 (N_8088,N_429,N_3044);
nor U8089 (N_8089,N_4481,N_3516);
xnor U8090 (N_8090,N_2981,N_1898);
nand U8091 (N_8091,N_682,N_4206);
and U8092 (N_8092,N_678,N_19);
xnor U8093 (N_8093,N_645,N_4007);
nand U8094 (N_8094,N_1873,N_531);
and U8095 (N_8095,N_367,N_2779);
xnor U8096 (N_8096,N_359,N_3033);
nand U8097 (N_8097,N_4316,N_2402);
or U8098 (N_8098,N_793,N_4858);
xnor U8099 (N_8099,N_2154,N_2722);
xnor U8100 (N_8100,N_1439,N_4343);
and U8101 (N_8101,N_2480,N_2349);
nand U8102 (N_8102,N_1852,N_4479);
or U8103 (N_8103,N_1878,N_3699);
nor U8104 (N_8104,N_3090,N_1246);
nor U8105 (N_8105,N_943,N_4274);
nand U8106 (N_8106,N_2279,N_2726);
nand U8107 (N_8107,N_3639,N_2049);
xor U8108 (N_8108,N_2039,N_977);
or U8109 (N_8109,N_2370,N_4308);
xnor U8110 (N_8110,N_3696,N_2772);
nor U8111 (N_8111,N_4969,N_4897);
or U8112 (N_8112,N_692,N_1694);
and U8113 (N_8113,N_2359,N_3564);
and U8114 (N_8114,N_3742,N_113);
or U8115 (N_8115,N_26,N_1441);
and U8116 (N_8116,N_1825,N_3544);
nor U8117 (N_8117,N_3923,N_2868);
nand U8118 (N_8118,N_4012,N_3961);
nor U8119 (N_8119,N_4983,N_529);
nand U8120 (N_8120,N_4944,N_18);
nor U8121 (N_8121,N_4174,N_1036);
nand U8122 (N_8122,N_3420,N_583);
nor U8123 (N_8123,N_4661,N_94);
xor U8124 (N_8124,N_3615,N_4188);
nand U8125 (N_8125,N_1336,N_2281);
xnor U8126 (N_8126,N_2683,N_4384);
and U8127 (N_8127,N_2685,N_2734);
and U8128 (N_8128,N_739,N_768);
nor U8129 (N_8129,N_1706,N_4432);
nor U8130 (N_8130,N_410,N_4729);
xor U8131 (N_8131,N_4901,N_3579);
xnor U8132 (N_8132,N_758,N_4544);
nor U8133 (N_8133,N_2088,N_1579);
nor U8134 (N_8134,N_1301,N_2249);
xnor U8135 (N_8135,N_4579,N_974);
xor U8136 (N_8136,N_2009,N_3303);
xor U8137 (N_8137,N_2250,N_2625);
nor U8138 (N_8138,N_4375,N_4685);
and U8139 (N_8139,N_3062,N_253);
nor U8140 (N_8140,N_1066,N_1254);
or U8141 (N_8141,N_3321,N_2363);
and U8142 (N_8142,N_1103,N_2454);
xor U8143 (N_8143,N_2415,N_1408);
xnor U8144 (N_8144,N_4114,N_4174);
nor U8145 (N_8145,N_2477,N_3949);
nor U8146 (N_8146,N_2600,N_2255);
nand U8147 (N_8147,N_759,N_2751);
xor U8148 (N_8148,N_4243,N_234);
and U8149 (N_8149,N_2764,N_2053);
or U8150 (N_8150,N_4100,N_516);
xor U8151 (N_8151,N_1080,N_4484);
and U8152 (N_8152,N_2773,N_2953);
nand U8153 (N_8153,N_1970,N_356);
nand U8154 (N_8154,N_71,N_4039);
nor U8155 (N_8155,N_4342,N_1190);
xor U8156 (N_8156,N_3882,N_2755);
xnor U8157 (N_8157,N_3025,N_1611);
and U8158 (N_8158,N_272,N_3240);
nor U8159 (N_8159,N_4633,N_2072);
xnor U8160 (N_8160,N_218,N_377);
or U8161 (N_8161,N_2849,N_21);
and U8162 (N_8162,N_1957,N_3156);
xnor U8163 (N_8163,N_3388,N_4817);
xnor U8164 (N_8164,N_4867,N_763);
nor U8165 (N_8165,N_2180,N_2715);
and U8166 (N_8166,N_3059,N_764);
and U8167 (N_8167,N_4150,N_692);
nor U8168 (N_8168,N_4763,N_3983);
or U8169 (N_8169,N_945,N_4061);
and U8170 (N_8170,N_4230,N_1653);
xor U8171 (N_8171,N_24,N_3227);
xor U8172 (N_8172,N_4880,N_4064);
nand U8173 (N_8173,N_3374,N_369);
xor U8174 (N_8174,N_1459,N_1572);
nor U8175 (N_8175,N_2635,N_2991);
and U8176 (N_8176,N_3421,N_3898);
or U8177 (N_8177,N_3877,N_4201);
nor U8178 (N_8178,N_1175,N_3291);
or U8179 (N_8179,N_1038,N_1481);
or U8180 (N_8180,N_483,N_782);
nor U8181 (N_8181,N_721,N_2369);
nor U8182 (N_8182,N_2699,N_4105);
xnor U8183 (N_8183,N_2267,N_3677);
xor U8184 (N_8184,N_1188,N_2002);
nand U8185 (N_8185,N_1973,N_3261);
nor U8186 (N_8186,N_4430,N_1788);
xnor U8187 (N_8187,N_2141,N_3972);
or U8188 (N_8188,N_946,N_3065);
nand U8189 (N_8189,N_1724,N_2370);
nand U8190 (N_8190,N_3266,N_1479);
nand U8191 (N_8191,N_1967,N_3411);
nand U8192 (N_8192,N_3852,N_638);
or U8193 (N_8193,N_2636,N_3347);
or U8194 (N_8194,N_1270,N_781);
xor U8195 (N_8195,N_2028,N_584);
or U8196 (N_8196,N_1628,N_1670);
nor U8197 (N_8197,N_3613,N_3274);
nand U8198 (N_8198,N_3288,N_3006);
nand U8199 (N_8199,N_483,N_4861);
nand U8200 (N_8200,N_252,N_3);
xnor U8201 (N_8201,N_4709,N_691);
nand U8202 (N_8202,N_2237,N_240);
nor U8203 (N_8203,N_1129,N_2838);
and U8204 (N_8204,N_4383,N_1662);
nand U8205 (N_8205,N_2198,N_3069);
or U8206 (N_8206,N_2001,N_4029);
nand U8207 (N_8207,N_1538,N_2175);
or U8208 (N_8208,N_4332,N_2235);
xnor U8209 (N_8209,N_1597,N_253);
nand U8210 (N_8210,N_4550,N_4586);
nand U8211 (N_8211,N_2687,N_162);
xor U8212 (N_8212,N_1215,N_4313);
xor U8213 (N_8213,N_1731,N_294);
nand U8214 (N_8214,N_358,N_4817);
nor U8215 (N_8215,N_4471,N_4971);
nand U8216 (N_8216,N_1323,N_3890);
and U8217 (N_8217,N_1126,N_4123);
and U8218 (N_8218,N_4678,N_1603);
or U8219 (N_8219,N_3257,N_3710);
and U8220 (N_8220,N_1018,N_2506);
nand U8221 (N_8221,N_5,N_1252);
and U8222 (N_8222,N_4146,N_4086);
and U8223 (N_8223,N_74,N_4961);
or U8224 (N_8224,N_1572,N_1540);
and U8225 (N_8225,N_3792,N_3393);
nand U8226 (N_8226,N_4775,N_4296);
nand U8227 (N_8227,N_3375,N_2221);
nand U8228 (N_8228,N_4074,N_2538);
nand U8229 (N_8229,N_690,N_2922);
nor U8230 (N_8230,N_2063,N_710);
nor U8231 (N_8231,N_1818,N_4389);
nor U8232 (N_8232,N_4358,N_3715);
nand U8233 (N_8233,N_828,N_371);
nor U8234 (N_8234,N_4302,N_585);
nor U8235 (N_8235,N_4565,N_1996);
nor U8236 (N_8236,N_918,N_4430);
and U8237 (N_8237,N_2714,N_616);
or U8238 (N_8238,N_2773,N_2035);
and U8239 (N_8239,N_4799,N_2970);
or U8240 (N_8240,N_2347,N_1535);
or U8241 (N_8241,N_2659,N_2646);
or U8242 (N_8242,N_1520,N_2501);
nand U8243 (N_8243,N_1164,N_2986);
or U8244 (N_8244,N_4659,N_4807);
or U8245 (N_8245,N_1277,N_1135);
nor U8246 (N_8246,N_4661,N_1077);
nor U8247 (N_8247,N_2296,N_293);
xnor U8248 (N_8248,N_4885,N_3000);
nor U8249 (N_8249,N_4154,N_2184);
nand U8250 (N_8250,N_3907,N_597);
or U8251 (N_8251,N_3903,N_1498);
and U8252 (N_8252,N_4950,N_4598);
nor U8253 (N_8253,N_3465,N_1900);
nand U8254 (N_8254,N_3272,N_1048);
nor U8255 (N_8255,N_1258,N_3028);
or U8256 (N_8256,N_4078,N_2748);
nor U8257 (N_8257,N_2037,N_4896);
and U8258 (N_8258,N_4700,N_3346);
xnor U8259 (N_8259,N_3506,N_4962);
or U8260 (N_8260,N_3510,N_1748);
and U8261 (N_8261,N_1566,N_2690);
nor U8262 (N_8262,N_4006,N_577);
nand U8263 (N_8263,N_902,N_78);
nand U8264 (N_8264,N_182,N_3205);
nand U8265 (N_8265,N_4946,N_2590);
xor U8266 (N_8266,N_4742,N_1424);
nand U8267 (N_8267,N_4762,N_3304);
and U8268 (N_8268,N_875,N_3539);
nor U8269 (N_8269,N_3378,N_261);
and U8270 (N_8270,N_1096,N_4734);
or U8271 (N_8271,N_3926,N_4245);
xor U8272 (N_8272,N_4184,N_4558);
nand U8273 (N_8273,N_2953,N_4389);
xor U8274 (N_8274,N_2103,N_2447);
and U8275 (N_8275,N_4542,N_1270);
and U8276 (N_8276,N_210,N_1887);
xor U8277 (N_8277,N_2127,N_2564);
nor U8278 (N_8278,N_3110,N_43);
and U8279 (N_8279,N_1975,N_4671);
nand U8280 (N_8280,N_2854,N_2846);
xnor U8281 (N_8281,N_320,N_3609);
xnor U8282 (N_8282,N_3032,N_4479);
or U8283 (N_8283,N_396,N_934);
and U8284 (N_8284,N_1587,N_4452);
nand U8285 (N_8285,N_620,N_3513);
xor U8286 (N_8286,N_411,N_1604);
or U8287 (N_8287,N_218,N_1627);
or U8288 (N_8288,N_4107,N_2407);
and U8289 (N_8289,N_2349,N_3572);
nand U8290 (N_8290,N_2512,N_4330);
xor U8291 (N_8291,N_3643,N_2633);
nor U8292 (N_8292,N_516,N_1141);
nand U8293 (N_8293,N_2378,N_1938);
nor U8294 (N_8294,N_3241,N_3858);
nand U8295 (N_8295,N_3310,N_3400);
and U8296 (N_8296,N_1448,N_4369);
and U8297 (N_8297,N_3338,N_2972);
and U8298 (N_8298,N_4984,N_3011);
nand U8299 (N_8299,N_2059,N_4719);
or U8300 (N_8300,N_3186,N_569);
nor U8301 (N_8301,N_3565,N_3810);
or U8302 (N_8302,N_2967,N_4479);
or U8303 (N_8303,N_3488,N_3245);
xor U8304 (N_8304,N_4344,N_1683);
nor U8305 (N_8305,N_4423,N_3078);
and U8306 (N_8306,N_3170,N_4021);
nand U8307 (N_8307,N_119,N_2425);
nand U8308 (N_8308,N_3370,N_3881);
nand U8309 (N_8309,N_360,N_641);
nand U8310 (N_8310,N_1266,N_1349);
nor U8311 (N_8311,N_4687,N_1064);
xor U8312 (N_8312,N_2688,N_2922);
or U8313 (N_8313,N_4717,N_2902);
nor U8314 (N_8314,N_2285,N_3920);
or U8315 (N_8315,N_2819,N_4637);
nand U8316 (N_8316,N_1448,N_1219);
and U8317 (N_8317,N_1228,N_1811);
xnor U8318 (N_8318,N_76,N_1509);
xor U8319 (N_8319,N_4004,N_2322);
nor U8320 (N_8320,N_4568,N_695);
nor U8321 (N_8321,N_1585,N_3582);
and U8322 (N_8322,N_243,N_3298);
nor U8323 (N_8323,N_2589,N_3114);
and U8324 (N_8324,N_3295,N_208);
xor U8325 (N_8325,N_1557,N_1656);
and U8326 (N_8326,N_3367,N_1591);
or U8327 (N_8327,N_2202,N_4764);
and U8328 (N_8328,N_3877,N_2172);
or U8329 (N_8329,N_2180,N_2845);
nor U8330 (N_8330,N_3108,N_1393);
and U8331 (N_8331,N_1538,N_4076);
nand U8332 (N_8332,N_4091,N_1984);
nor U8333 (N_8333,N_1925,N_2259);
xor U8334 (N_8334,N_1978,N_1152);
xnor U8335 (N_8335,N_4208,N_162);
nor U8336 (N_8336,N_2328,N_4161);
nand U8337 (N_8337,N_947,N_3594);
nand U8338 (N_8338,N_3933,N_2354);
or U8339 (N_8339,N_4310,N_415);
nand U8340 (N_8340,N_958,N_3699);
xnor U8341 (N_8341,N_4654,N_123);
nor U8342 (N_8342,N_1602,N_1174);
nor U8343 (N_8343,N_3634,N_3);
nand U8344 (N_8344,N_16,N_4360);
nand U8345 (N_8345,N_1945,N_263);
nor U8346 (N_8346,N_2460,N_3279);
nand U8347 (N_8347,N_1355,N_1769);
nor U8348 (N_8348,N_4989,N_4188);
nor U8349 (N_8349,N_927,N_2229);
xnor U8350 (N_8350,N_412,N_3188);
or U8351 (N_8351,N_4899,N_3714);
nand U8352 (N_8352,N_458,N_1187);
nor U8353 (N_8353,N_1855,N_3918);
or U8354 (N_8354,N_4980,N_4096);
xnor U8355 (N_8355,N_1685,N_1992);
nor U8356 (N_8356,N_1126,N_626);
or U8357 (N_8357,N_4798,N_1158);
nand U8358 (N_8358,N_1816,N_4290);
xnor U8359 (N_8359,N_621,N_4396);
and U8360 (N_8360,N_503,N_3465);
and U8361 (N_8361,N_4977,N_2197);
or U8362 (N_8362,N_4843,N_3769);
xor U8363 (N_8363,N_797,N_1555);
or U8364 (N_8364,N_4180,N_1666);
xor U8365 (N_8365,N_2015,N_352);
xnor U8366 (N_8366,N_2540,N_1321);
and U8367 (N_8367,N_2225,N_2476);
and U8368 (N_8368,N_438,N_4712);
or U8369 (N_8369,N_2128,N_710);
nand U8370 (N_8370,N_1102,N_3119);
and U8371 (N_8371,N_4621,N_3543);
xnor U8372 (N_8372,N_2204,N_4376);
xor U8373 (N_8373,N_1610,N_335);
xor U8374 (N_8374,N_1315,N_3851);
xnor U8375 (N_8375,N_2510,N_2484);
or U8376 (N_8376,N_521,N_1906);
and U8377 (N_8377,N_1101,N_4161);
and U8378 (N_8378,N_655,N_1728);
xnor U8379 (N_8379,N_4454,N_3877);
or U8380 (N_8380,N_3786,N_4158);
nor U8381 (N_8381,N_2723,N_4774);
and U8382 (N_8382,N_413,N_60);
or U8383 (N_8383,N_1847,N_933);
xnor U8384 (N_8384,N_122,N_2675);
xor U8385 (N_8385,N_1715,N_2504);
and U8386 (N_8386,N_3433,N_368);
nor U8387 (N_8387,N_237,N_3723);
nand U8388 (N_8388,N_2496,N_4087);
or U8389 (N_8389,N_1150,N_4461);
or U8390 (N_8390,N_2137,N_3736);
or U8391 (N_8391,N_4755,N_94);
or U8392 (N_8392,N_1385,N_2323);
xor U8393 (N_8393,N_4788,N_686);
nand U8394 (N_8394,N_4073,N_4199);
nand U8395 (N_8395,N_1396,N_1044);
nor U8396 (N_8396,N_632,N_4667);
nand U8397 (N_8397,N_4845,N_4104);
and U8398 (N_8398,N_4394,N_2233);
or U8399 (N_8399,N_3608,N_4568);
or U8400 (N_8400,N_1062,N_2666);
nor U8401 (N_8401,N_1995,N_1059);
or U8402 (N_8402,N_4810,N_3011);
xor U8403 (N_8403,N_1874,N_1293);
xnor U8404 (N_8404,N_4143,N_4638);
and U8405 (N_8405,N_3895,N_1927);
xnor U8406 (N_8406,N_3754,N_3037);
nor U8407 (N_8407,N_2176,N_3963);
xnor U8408 (N_8408,N_4895,N_3300);
xor U8409 (N_8409,N_2934,N_3811);
xor U8410 (N_8410,N_4312,N_1286);
or U8411 (N_8411,N_4262,N_471);
xor U8412 (N_8412,N_2955,N_1274);
nand U8413 (N_8413,N_3173,N_843);
xnor U8414 (N_8414,N_3199,N_3072);
nand U8415 (N_8415,N_3159,N_1744);
nand U8416 (N_8416,N_4107,N_3171);
xor U8417 (N_8417,N_4553,N_2421);
nand U8418 (N_8418,N_1081,N_3300);
xnor U8419 (N_8419,N_3199,N_2582);
xor U8420 (N_8420,N_693,N_1884);
and U8421 (N_8421,N_1320,N_2616);
xnor U8422 (N_8422,N_2766,N_4458);
or U8423 (N_8423,N_4832,N_1882);
nand U8424 (N_8424,N_3814,N_58);
nand U8425 (N_8425,N_2353,N_1353);
nor U8426 (N_8426,N_819,N_3259);
or U8427 (N_8427,N_816,N_3360);
nor U8428 (N_8428,N_476,N_4608);
and U8429 (N_8429,N_3913,N_3916);
or U8430 (N_8430,N_1934,N_2209);
nand U8431 (N_8431,N_1256,N_1381);
xor U8432 (N_8432,N_951,N_4556);
nor U8433 (N_8433,N_3982,N_354);
nor U8434 (N_8434,N_1248,N_3971);
nand U8435 (N_8435,N_1496,N_477);
or U8436 (N_8436,N_4994,N_3105);
xnor U8437 (N_8437,N_3573,N_2979);
and U8438 (N_8438,N_3545,N_1401);
nor U8439 (N_8439,N_1131,N_2081);
and U8440 (N_8440,N_2285,N_3828);
xnor U8441 (N_8441,N_4988,N_4313);
xor U8442 (N_8442,N_2608,N_81);
nand U8443 (N_8443,N_249,N_464);
and U8444 (N_8444,N_4962,N_4245);
nor U8445 (N_8445,N_1357,N_3689);
and U8446 (N_8446,N_4702,N_1169);
nor U8447 (N_8447,N_1394,N_3586);
nor U8448 (N_8448,N_4688,N_10);
and U8449 (N_8449,N_2895,N_22);
nand U8450 (N_8450,N_2422,N_4947);
nor U8451 (N_8451,N_2874,N_4630);
nor U8452 (N_8452,N_4617,N_4505);
xor U8453 (N_8453,N_4561,N_1380);
xnor U8454 (N_8454,N_892,N_3190);
nand U8455 (N_8455,N_249,N_2500);
nor U8456 (N_8456,N_69,N_1728);
nor U8457 (N_8457,N_1561,N_1332);
xor U8458 (N_8458,N_185,N_4959);
nor U8459 (N_8459,N_4806,N_713);
nor U8460 (N_8460,N_2357,N_4552);
nand U8461 (N_8461,N_2696,N_1532);
xnor U8462 (N_8462,N_685,N_4139);
and U8463 (N_8463,N_2814,N_4410);
and U8464 (N_8464,N_1184,N_1937);
nand U8465 (N_8465,N_4200,N_4358);
and U8466 (N_8466,N_1115,N_2519);
xnor U8467 (N_8467,N_839,N_464);
or U8468 (N_8468,N_964,N_4133);
nor U8469 (N_8469,N_1193,N_3342);
nand U8470 (N_8470,N_547,N_3042);
xnor U8471 (N_8471,N_3201,N_1397);
nand U8472 (N_8472,N_2095,N_493);
nand U8473 (N_8473,N_1078,N_2169);
or U8474 (N_8474,N_2163,N_4345);
nand U8475 (N_8475,N_4245,N_2682);
or U8476 (N_8476,N_3030,N_1184);
xor U8477 (N_8477,N_3994,N_2496);
xor U8478 (N_8478,N_2544,N_4819);
or U8479 (N_8479,N_611,N_1591);
nor U8480 (N_8480,N_2566,N_3758);
and U8481 (N_8481,N_4915,N_1706);
or U8482 (N_8482,N_1037,N_2712);
and U8483 (N_8483,N_655,N_436);
or U8484 (N_8484,N_289,N_1822);
nor U8485 (N_8485,N_3215,N_1356);
and U8486 (N_8486,N_3088,N_1086);
nor U8487 (N_8487,N_778,N_2840);
nor U8488 (N_8488,N_3941,N_4538);
xnor U8489 (N_8489,N_1547,N_1575);
nor U8490 (N_8490,N_478,N_2361);
nor U8491 (N_8491,N_2032,N_2059);
nor U8492 (N_8492,N_4622,N_3075);
or U8493 (N_8493,N_796,N_1465);
nor U8494 (N_8494,N_2215,N_2254);
or U8495 (N_8495,N_757,N_3221);
nor U8496 (N_8496,N_904,N_4546);
nand U8497 (N_8497,N_117,N_401);
nand U8498 (N_8498,N_2554,N_3440);
xnor U8499 (N_8499,N_3175,N_337);
xor U8500 (N_8500,N_955,N_4607);
nand U8501 (N_8501,N_398,N_2994);
xor U8502 (N_8502,N_1387,N_1498);
xor U8503 (N_8503,N_447,N_3684);
nand U8504 (N_8504,N_152,N_2011);
nand U8505 (N_8505,N_727,N_3557);
xnor U8506 (N_8506,N_1673,N_1762);
or U8507 (N_8507,N_1055,N_2620);
or U8508 (N_8508,N_2874,N_259);
and U8509 (N_8509,N_352,N_3905);
and U8510 (N_8510,N_3591,N_1183);
or U8511 (N_8511,N_3134,N_4134);
and U8512 (N_8512,N_1129,N_729);
and U8513 (N_8513,N_2949,N_3859);
xor U8514 (N_8514,N_2938,N_4106);
or U8515 (N_8515,N_2995,N_4691);
nor U8516 (N_8516,N_2682,N_760);
xor U8517 (N_8517,N_4134,N_4637);
nor U8518 (N_8518,N_1461,N_1729);
or U8519 (N_8519,N_2696,N_3707);
nand U8520 (N_8520,N_41,N_473);
nand U8521 (N_8521,N_1934,N_4085);
and U8522 (N_8522,N_1438,N_3761);
and U8523 (N_8523,N_4687,N_855);
nand U8524 (N_8524,N_2096,N_4242);
xnor U8525 (N_8525,N_4531,N_2847);
nand U8526 (N_8526,N_3858,N_3124);
and U8527 (N_8527,N_3548,N_2871);
nor U8528 (N_8528,N_3430,N_73);
nor U8529 (N_8529,N_2731,N_1793);
xnor U8530 (N_8530,N_3024,N_1224);
and U8531 (N_8531,N_4228,N_4170);
nor U8532 (N_8532,N_934,N_4879);
nand U8533 (N_8533,N_3554,N_4001);
xor U8534 (N_8534,N_1486,N_2718);
xor U8535 (N_8535,N_3203,N_4903);
and U8536 (N_8536,N_3589,N_124);
xor U8537 (N_8537,N_2766,N_1292);
and U8538 (N_8538,N_4349,N_704);
and U8539 (N_8539,N_98,N_930);
and U8540 (N_8540,N_2200,N_1474);
nor U8541 (N_8541,N_4748,N_2062);
and U8542 (N_8542,N_2379,N_1998);
xor U8543 (N_8543,N_1990,N_3615);
and U8544 (N_8544,N_3495,N_4289);
nor U8545 (N_8545,N_1168,N_3229);
nor U8546 (N_8546,N_2292,N_2820);
xor U8547 (N_8547,N_678,N_4054);
nor U8548 (N_8548,N_94,N_977);
and U8549 (N_8549,N_2137,N_614);
or U8550 (N_8550,N_4463,N_3016);
nor U8551 (N_8551,N_2559,N_2465);
or U8552 (N_8552,N_3993,N_3995);
nand U8553 (N_8553,N_2541,N_421);
nor U8554 (N_8554,N_206,N_2054);
nand U8555 (N_8555,N_4504,N_1084);
nand U8556 (N_8556,N_242,N_1603);
xor U8557 (N_8557,N_4649,N_3730);
nor U8558 (N_8558,N_900,N_1650);
or U8559 (N_8559,N_2833,N_4605);
or U8560 (N_8560,N_117,N_3304);
xnor U8561 (N_8561,N_3403,N_4709);
or U8562 (N_8562,N_3732,N_4813);
nor U8563 (N_8563,N_2583,N_2574);
nand U8564 (N_8564,N_3953,N_2939);
and U8565 (N_8565,N_3968,N_236);
and U8566 (N_8566,N_3118,N_2292);
or U8567 (N_8567,N_2019,N_3729);
or U8568 (N_8568,N_4268,N_4587);
nor U8569 (N_8569,N_1003,N_4254);
nand U8570 (N_8570,N_2546,N_899);
nand U8571 (N_8571,N_817,N_986);
and U8572 (N_8572,N_1219,N_4011);
nand U8573 (N_8573,N_4630,N_289);
xor U8574 (N_8574,N_2287,N_1357);
and U8575 (N_8575,N_4065,N_2560);
or U8576 (N_8576,N_2960,N_3944);
nor U8577 (N_8577,N_3522,N_3561);
nand U8578 (N_8578,N_4006,N_3730);
nor U8579 (N_8579,N_3809,N_3876);
nand U8580 (N_8580,N_4592,N_402);
nand U8581 (N_8581,N_2283,N_3039);
xnor U8582 (N_8582,N_72,N_4870);
or U8583 (N_8583,N_4026,N_995);
nand U8584 (N_8584,N_1539,N_3076);
xnor U8585 (N_8585,N_1024,N_3223);
and U8586 (N_8586,N_864,N_2959);
nor U8587 (N_8587,N_1796,N_4865);
or U8588 (N_8588,N_4773,N_4301);
nor U8589 (N_8589,N_3068,N_295);
or U8590 (N_8590,N_429,N_772);
nand U8591 (N_8591,N_1918,N_2365);
xnor U8592 (N_8592,N_1717,N_3258);
nor U8593 (N_8593,N_932,N_1527);
xor U8594 (N_8594,N_4662,N_1868);
and U8595 (N_8595,N_202,N_4829);
nand U8596 (N_8596,N_1371,N_4680);
nor U8597 (N_8597,N_2818,N_4776);
nor U8598 (N_8598,N_504,N_3107);
nor U8599 (N_8599,N_1829,N_2);
or U8600 (N_8600,N_708,N_2727);
xor U8601 (N_8601,N_3593,N_3714);
nand U8602 (N_8602,N_3457,N_3812);
and U8603 (N_8603,N_3182,N_3433);
xor U8604 (N_8604,N_467,N_2850);
nand U8605 (N_8605,N_4246,N_1129);
nand U8606 (N_8606,N_1999,N_4795);
nand U8607 (N_8607,N_199,N_3574);
xor U8608 (N_8608,N_2453,N_4548);
and U8609 (N_8609,N_1699,N_3702);
nor U8610 (N_8610,N_1911,N_2139);
and U8611 (N_8611,N_4940,N_2531);
xnor U8612 (N_8612,N_2007,N_4996);
or U8613 (N_8613,N_78,N_2000);
nand U8614 (N_8614,N_4705,N_3178);
and U8615 (N_8615,N_37,N_937);
or U8616 (N_8616,N_4507,N_2398);
nor U8617 (N_8617,N_2844,N_3071);
xnor U8618 (N_8618,N_334,N_3135);
and U8619 (N_8619,N_2181,N_3936);
nor U8620 (N_8620,N_4601,N_3057);
nand U8621 (N_8621,N_594,N_3749);
and U8622 (N_8622,N_147,N_2950);
or U8623 (N_8623,N_2576,N_1760);
and U8624 (N_8624,N_996,N_3489);
and U8625 (N_8625,N_1432,N_2684);
nor U8626 (N_8626,N_4200,N_4800);
nor U8627 (N_8627,N_106,N_1254);
nor U8628 (N_8628,N_2210,N_4084);
and U8629 (N_8629,N_2708,N_3005);
xnor U8630 (N_8630,N_297,N_3359);
or U8631 (N_8631,N_1270,N_4696);
nand U8632 (N_8632,N_3220,N_794);
and U8633 (N_8633,N_2701,N_2540);
nand U8634 (N_8634,N_177,N_3773);
nand U8635 (N_8635,N_2122,N_774);
nand U8636 (N_8636,N_3500,N_4674);
or U8637 (N_8637,N_4899,N_477);
nand U8638 (N_8638,N_3465,N_3730);
and U8639 (N_8639,N_1346,N_3736);
and U8640 (N_8640,N_2424,N_2961);
nand U8641 (N_8641,N_4960,N_1174);
nor U8642 (N_8642,N_2294,N_2796);
nor U8643 (N_8643,N_145,N_3777);
nor U8644 (N_8644,N_314,N_2796);
nor U8645 (N_8645,N_4019,N_2963);
nor U8646 (N_8646,N_803,N_3986);
nand U8647 (N_8647,N_1963,N_2703);
nand U8648 (N_8648,N_2909,N_131);
nor U8649 (N_8649,N_2940,N_1185);
nand U8650 (N_8650,N_4066,N_1906);
nand U8651 (N_8651,N_4321,N_1656);
xor U8652 (N_8652,N_354,N_2235);
and U8653 (N_8653,N_591,N_4618);
or U8654 (N_8654,N_2681,N_3028);
and U8655 (N_8655,N_4522,N_3290);
or U8656 (N_8656,N_3107,N_4076);
xnor U8657 (N_8657,N_2687,N_2556);
or U8658 (N_8658,N_392,N_3097);
xnor U8659 (N_8659,N_4137,N_3904);
xnor U8660 (N_8660,N_3989,N_3346);
nand U8661 (N_8661,N_4016,N_3965);
and U8662 (N_8662,N_3173,N_3142);
xor U8663 (N_8663,N_52,N_4468);
nor U8664 (N_8664,N_3929,N_2719);
or U8665 (N_8665,N_4299,N_915);
xor U8666 (N_8666,N_4429,N_1313);
and U8667 (N_8667,N_4173,N_3270);
and U8668 (N_8668,N_2921,N_847);
and U8669 (N_8669,N_1440,N_3914);
and U8670 (N_8670,N_2041,N_2185);
and U8671 (N_8671,N_4550,N_1310);
and U8672 (N_8672,N_1817,N_839);
nand U8673 (N_8673,N_1030,N_326);
or U8674 (N_8674,N_624,N_2884);
and U8675 (N_8675,N_22,N_624);
nor U8676 (N_8676,N_3561,N_126);
or U8677 (N_8677,N_79,N_3801);
nand U8678 (N_8678,N_3983,N_3787);
and U8679 (N_8679,N_811,N_2105);
and U8680 (N_8680,N_437,N_4356);
and U8681 (N_8681,N_649,N_3057);
and U8682 (N_8682,N_2300,N_189);
xnor U8683 (N_8683,N_2496,N_3891);
nand U8684 (N_8684,N_2136,N_4928);
or U8685 (N_8685,N_1228,N_2192);
or U8686 (N_8686,N_1569,N_1085);
xnor U8687 (N_8687,N_3214,N_1820);
nand U8688 (N_8688,N_3718,N_4331);
or U8689 (N_8689,N_1267,N_4036);
or U8690 (N_8690,N_3939,N_4284);
xor U8691 (N_8691,N_709,N_2026);
and U8692 (N_8692,N_2796,N_3167);
and U8693 (N_8693,N_4739,N_3806);
nand U8694 (N_8694,N_3076,N_4669);
and U8695 (N_8695,N_1919,N_2216);
xor U8696 (N_8696,N_40,N_1163);
xor U8697 (N_8697,N_1312,N_4594);
or U8698 (N_8698,N_2911,N_2188);
nor U8699 (N_8699,N_4896,N_4061);
nor U8700 (N_8700,N_385,N_2662);
nor U8701 (N_8701,N_193,N_274);
nand U8702 (N_8702,N_4607,N_4260);
nor U8703 (N_8703,N_1923,N_318);
nor U8704 (N_8704,N_3606,N_313);
xnor U8705 (N_8705,N_1431,N_4080);
nor U8706 (N_8706,N_3723,N_685);
nand U8707 (N_8707,N_57,N_3851);
nor U8708 (N_8708,N_3218,N_1145);
or U8709 (N_8709,N_1943,N_3164);
and U8710 (N_8710,N_2823,N_1354);
or U8711 (N_8711,N_4937,N_511);
nor U8712 (N_8712,N_3097,N_3548);
or U8713 (N_8713,N_2380,N_615);
or U8714 (N_8714,N_2867,N_4577);
or U8715 (N_8715,N_894,N_4871);
nand U8716 (N_8716,N_4463,N_4081);
or U8717 (N_8717,N_4267,N_2035);
or U8718 (N_8718,N_3203,N_470);
nor U8719 (N_8719,N_1638,N_3517);
and U8720 (N_8720,N_2381,N_3152);
nand U8721 (N_8721,N_3496,N_4402);
nor U8722 (N_8722,N_1785,N_697);
or U8723 (N_8723,N_247,N_803);
nor U8724 (N_8724,N_1731,N_4348);
nand U8725 (N_8725,N_351,N_4842);
nor U8726 (N_8726,N_66,N_2061);
nand U8727 (N_8727,N_756,N_2416);
nor U8728 (N_8728,N_105,N_308);
xor U8729 (N_8729,N_4966,N_3091);
nor U8730 (N_8730,N_4194,N_1617);
nor U8731 (N_8731,N_341,N_2270);
xor U8732 (N_8732,N_720,N_4714);
and U8733 (N_8733,N_633,N_3567);
nor U8734 (N_8734,N_1855,N_4734);
or U8735 (N_8735,N_1049,N_118);
and U8736 (N_8736,N_3823,N_89);
or U8737 (N_8737,N_1788,N_4201);
or U8738 (N_8738,N_114,N_1429);
and U8739 (N_8739,N_3054,N_3510);
or U8740 (N_8740,N_3280,N_4615);
and U8741 (N_8741,N_693,N_869);
nor U8742 (N_8742,N_3232,N_2882);
or U8743 (N_8743,N_667,N_3870);
and U8744 (N_8744,N_1112,N_3009);
nor U8745 (N_8745,N_4050,N_4058);
xnor U8746 (N_8746,N_4229,N_1650);
xnor U8747 (N_8747,N_2787,N_4305);
and U8748 (N_8748,N_4253,N_1571);
nor U8749 (N_8749,N_3840,N_4217);
or U8750 (N_8750,N_957,N_1327);
or U8751 (N_8751,N_2187,N_4041);
or U8752 (N_8752,N_3166,N_4815);
and U8753 (N_8753,N_4253,N_4946);
xor U8754 (N_8754,N_2928,N_3676);
and U8755 (N_8755,N_608,N_583);
nand U8756 (N_8756,N_844,N_2384);
nand U8757 (N_8757,N_1451,N_3528);
nand U8758 (N_8758,N_152,N_3738);
nand U8759 (N_8759,N_2738,N_2442);
and U8760 (N_8760,N_4716,N_4999);
or U8761 (N_8761,N_4009,N_2944);
nand U8762 (N_8762,N_2782,N_1730);
nand U8763 (N_8763,N_2625,N_2055);
nor U8764 (N_8764,N_737,N_4021);
nand U8765 (N_8765,N_3278,N_4663);
and U8766 (N_8766,N_407,N_896);
or U8767 (N_8767,N_2881,N_2354);
and U8768 (N_8768,N_3544,N_1098);
nor U8769 (N_8769,N_2854,N_1695);
xor U8770 (N_8770,N_4523,N_4905);
or U8771 (N_8771,N_2796,N_4151);
or U8772 (N_8772,N_1347,N_3367);
nand U8773 (N_8773,N_991,N_3062);
nand U8774 (N_8774,N_3152,N_1797);
nand U8775 (N_8775,N_1900,N_2280);
and U8776 (N_8776,N_2778,N_2058);
xor U8777 (N_8777,N_4655,N_4507);
nand U8778 (N_8778,N_912,N_3533);
and U8779 (N_8779,N_2611,N_1553);
nand U8780 (N_8780,N_4526,N_2291);
nor U8781 (N_8781,N_248,N_4267);
nor U8782 (N_8782,N_2058,N_1297);
xnor U8783 (N_8783,N_383,N_4925);
xor U8784 (N_8784,N_4316,N_789);
or U8785 (N_8785,N_2322,N_4295);
nor U8786 (N_8786,N_672,N_3421);
and U8787 (N_8787,N_4033,N_3048);
nand U8788 (N_8788,N_1426,N_1549);
xnor U8789 (N_8789,N_4745,N_551);
or U8790 (N_8790,N_2975,N_699);
nor U8791 (N_8791,N_1929,N_3137);
and U8792 (N_8792,N_3840,N_3235);
and U8793 (N_8793,N_4496,N_3859);
or U8794 (N_8794,N_4966,N_1203);
and U8795 (N_8795,N_2913,N_127);
nor U8796 (N_8796,N_2866,N_1481);
and U8797 (N_8797,N_4161,N_2423);
or U8798 (N_8798,N_3093,N_4107);
and U8799 (N_8799,N_1202,N_3645);
nand U8800 (N_8800,N_1881,N_768);
nor U8801 (N_8801,N_1776,N_1536);
nand U8802 (N_8802,N_2640,N_460);
nor U8803 (N_8803,N_168,N_4745);
nor U8804 (N_8804,N_4284,N_2187);
nor U8805 (N_8805,N_3500,N_4000);
and U8806 (N_8806,N_4348,N_1647);
nor U8807 (N_8807,N_314,N_4577);
nor U8808 (N_8808,N_2129,N_511);
or U8809 (N_8809,N_1354,N_1324);
and U8810 (N_8810,N_1210,N_1175);
and U8811 (N_8811,N_121,N_1574);
xor U8812 (N_8812,N_1698,N_4958);
xnor U8813 (N_8813,N_4600,N_3971);
and U8814 (N_8814,N_4401,N_3190);
nand U8815 (N_8815,N_1149,N_1189);
nor U8816 (N_8816,N_4719,N_1435);
or U8817 (N_8817,N_1170,N_2907);
and U8818 (N_8818,N_4037,N_4294);
xor U8819 (N_8819,N_2098,N_173);
nor U8820 (N_8820,N_1802,N_3134);
xnor U8821 (N_8821,N_2900,N_1280);
nor U8822 (N_8822,N_3349,N_3421);
or U8823 (N_8823,N_2280,N_2516);
or U8824 (N_8824,N_666,N_1295);
nand U8825 (N_8825,N_1133,N_2264);
nand U8826 (N_8826,N_823,N_969);
nor U8827 (N_8827,N_1857,N_1232);
xor U8828 (N_8828,N_714,N_1012);
nand U8829 (N_8829,N_2390,N_2572);
xnor U8830 (N_8830,N_4854,N_2227);
xor U8831 (N_8831,N_2082,N_1864);
or U8832 (N_8832,N_1262,N_3847);
nor U8833 (N_8833,N_4537,N_3062);
nand U8834 (N_8834,N_4660,N_422);
nand U8835 (N_8835,N_4736,N_3732);
xor U8836 (N_8836,N_2309,N_735);
and U8837 (N_8837,N_1583,N_2208);
nor U8838 (N_8838,N_79,N_961);
and U8839 (N_8839,N_196,N_1485);
xor U8840 (N_8840,N_298,N_3583);
and U8841 (N_8841,N_2697,N_1020);
and U8842 (N_8842,N_1875,N_2912);
or U8843 (N_8843,N_4416,N_2289);
xor U8844 (N_8844,N_2412,N_3998);
nand U8845 (N_8845,N_4805,N_2080);
and U8846 (N_8846,N_3204,N_2639);
nand U8847 (N_8847,N_3754,N_3816);
xnor U8848 (N_8848,N_312,N_1535);
or U8849 (N_8849,N_4536,N_1027);
nand U8850 (N_8850,N_996,N_2874);
nand U8851 (N_8851,N_2755,N_4178);
and U8852 (N_8852,N_4276,N_1663);
nor U8853 (N_8853,N_192,N_4285);
or U8854 (N_8854,N_3636,N_4908);
and U8855 (N_8855,N_3144,N_3859);
nand U8856 (N_8856,N_2110,N_1021);
xnor U8857 (N_8857,N_1550,N_1877);
nand U8858 (N_8858,N_3739,N_4245);
nand U8859 (N_8859,N_3306,N_4835);
xnor U8860 (N_8860,N_3119,N_3670);
and U8861 (N_8861,N_1229,N_4756);
xnor U8862 (N_8862,N_1514,N_2171);
or U8863 (N_8863,N_235,N_912);
nand U8864 (N_8864,N_1920,N_2854);
nor U8865 (N_8865,N_4658,N_4630);
and U8866 (N_8866,N_1024,N_1178);
and U8867 (N_8867,N_152,N_2039);
nor U8868 (N_8868,N_3009,N_4649);
nand U8869 (N_8869,N_3394,N_2129);
nand U8870 (N_8870,N_2983,N_3967);
or U8871 (N_8871,N_3645,N_1312);
or U8872 (N_8872,N_1495,N_4053);
nand U8873 (N_8873,N_936,N_1688);
nand U8874 (N_8874,N_4929,N_993);
xnor U8875 (N_8875,N_4550,N_1239);
xnor U8876 (N_8876,N_1554,N_201);
nor U8877 (N_8877,N_442,N_3050);
xnor U8878 (N_8878,N_2970,N_2856);
and U8879 (N_8879,N_1021,N_3449);
and U8880 (N_8880,N_4938,N_392);
and U8881 (N_8881,N_2309,N_2712);
nor U8882 (N_8882,N_2228,N_2973);
or U8883 (N_8883,N_2110,N_2941);
or U8884 (N_8884,N_2991,N_2472);
or U8885 (N_8885,N_2757,N_2699);
or U8886 (N_8886,N_2988,N_1993);
nand U8887 (N_8887,N_3468,N_3668);
nand U8888 (N_8888,N_3751,N_3045);
nor U8889 (N_8889,N_1465,N_591);
xor U8890 (N_8890,N_297,N_4390);
or U8891 (N_8891,N_3132,N_4691);
nor U8892 (N_8892,N_3680,N_654);
xnor U8893 (N_8893,N_2173,N_4810);
xnor U8894 (N_8894,N_2982,N_3415);
xnor U8895 (N_8895,N_15,N_1710);
xor U8896 (N_8896,N_3691,N_546);
xor U8897 (N_8897,N_813,N_1053);
nor U8898 (N_8898,N_3226,N_2280);
and U8899 (N_8899,N_2446,N_3361);
xor U8900 (N_8900,N_2773,N_4116);
xor U8901 (N_8901,N_1953,N_4278);
or U8902 (N_8902,N_4226,N_4840);
and U8903 (N_8903,N_3209,N_822);
or U8904 (N_8904,N_4925,N_3598);
or U8905 (N_8905,N_4758,N_4140);
and U8906 (N_8906,N_1112,N_4825);
and U8907 (N_8907,N_3806,N_3687);
nand U8908 (N_8908,N_3369,N_2694);
nor U8909 (N_8909,N_690,N_3000);
xor U8910 (N_8910,N_3902,N_3912);
nor U8911 (N_8911,N_2667,N_147);
nand U8912 (N_8912,N_2339,N_4929);
and U8913 (N_8913,N_2319,N_4870);
and U8914 (N_8914,N_1221,N_1883);
nand U8915 (N_8915,N_2307,N_4310);
and U8916 (N_8916,N_106,N_9);
nor U8917 (N_8917,N_2052,N_4629);
or U8918 (N_8918,N_622,N_3485);
nor U8919 (N_8919,N_4213,N_4361);
and U8920 (N_8920,N_4222,N_1695);
and U8921 (N_8921,N_4454,N_125);
nor U8922 (N_8922,N_722,N_1965);
and U8923 (N_8923,N_3717,N_2027);
and U8924 (N_8924,N_1765,N_4186);
xnor U8925 (N_8925,N_4753,N_462);
and U8926 (N_8926,N_1768,N_504);
and U8927 (N_8927,N_3748,N_942);
xnor U8928 (N_8928,N_4892,N_4631);
xor U8929 (N_8929,N_1991,N_2011);
or U8930 (N_8930,N_4050,N_547);
nand U8931 (N_8931,N_3306,N_4167);
nand U8932 (N_8932,N_418,N_457);
xnor U8933 (N_8933,N_1810,N_2602);
and U8934 (N_8934,N_547,N_4045);
or U8935 (N_8935,N_533,N_4536);
or U8936 (N_8936,N_1666,N_2497);
and U8937 (N_8937,N_1104,N_703);
nand U8938 (N_8938,N_1958,N_2117);
nand U8939 (N_8939,N_2900,N_3675);
nand U8940 (N_8940,N_3125,N_3639);
or U8941 (N_8941,N_4160,N_4654);
or U8942 (N_8942,N_3022,N_4157);
xnor U8943 (N_8943,N_3778,N_4650);
or U8944 (N_8944,N_1371,N_1351);
nor U8945 (N_8945,N_1063,N_3404);
nor U8946 (N_8946,N_4098,N_3369);
or U8947 (N_8947,N_213,N_1445);
nand U8948 (N_8948,N_3722,N_4657);
xnor U8949 (N_8949,N_4896,N_4279);
or U8950 (N_8950,N_3071,N_2405);
or U8951 (N_8951,N_3494,N_3300);
or U8952 (N_8952,N_2819,N_1689);
or U8953 (N_8953,N_1411,N_738);
or U8954 (N_8954,N_4050,N_430);
and U8955 (N_8955,N_1609,N_740);
and U8956 (N_8956,N_2136,N_3229);
nand U8957 (N_8957,N_944,N_3057);
xnor U8958 (N_8958,N_4606,N_4008);
nand U8959 (N_8959,N_417,N_3691);
nor U8960 (N_8960,N_4092,N_1991);
or U8961 (N_8961,N_2146,N_4877);
xor U8962 (N_8962,N_2580,N_4858);
nor U8963 (N_8963,N_2252,N_4974);
or U8964 (N_8964,N_4284,N_1594);
nand U8965 (N_8965,N_1501,N_401);
nand U8966 (N_8966,N_595,N_1137);
and U8967 (N_8967,N_4846,N_1516);
nor U8968 (N_8968,N_659,N_1267);
and U8969 (N_8969,N_4322,N_1138);
or U8970 (N_8970,N_1576,N_3940);
nand U8971 (N_8971,N_1295,N_628);
nor U8972 (N_8972,N_2807,N_867);
xor U8973 (N_8973,N_2330,N_4423);
xnor U8974 (N_8974,N_3433,N_1736);
nand U8975 (N_8975,N_4796,N_1085);
nand U8976 (N_8976,N_669,N_1068);
xnor U8977 (N_8977,N_3000,N_2295);
xnor U8978 (N_8978,N_248,N_646);
nand U8979 (N_8979,N_2674,N_3123);
and U8980 (N_8980,N_3443,N_1999);
and U8981 (N_8981,N_4233,N_4930);
and U8982 (N_8982,N_4079,N_2869);
or U8983 (N_8983,N_763,N_1610);
xnor U8984 (N_8984,N_1070,N_1917);
nor U8985 (N_8985,N_3343,N_3920);
and U8986 (N_8986,N_4400,N_2307);
and U8987 (N_8987,N_2862,N_1323);
xnor U8988 (N_8988,N_3282,N_3951);
nand U8989 (N_8989,N_1401,N_4560);
and U8990 (N_8990,N_40,N_4777);
and U8991 (N_8991,N_3888,N_3166);
xnor U8992 (N_8992,N_4457,N_608);
nor U8993 (N_8993,N_1315,N_4181);
xnor U8994 (N_8994,N_1269,N_3913);
or U8995 (N_8995,N_4181,N_3985);
nand U8996 (N_8996,N_3892,N_3729);
and U8997 (N_8997,N_793,N_385);
xor U8998 (N_8998,N_791,N_561);
nor U8999 (N_8999,N_1146,N_207);
nor U9000 (N_9000,N_2799,N_687);
or U9001 (N_9001,N_1799,N_1009);
nand U9002 (N_9002,N_72,N_34);
or U9003 (N_9003,N_3372,N_4753);
and U9004 (N_9004,N_4883,N_3258);
and U9005 (N_9005,N_1438,N_3536);
nor U9006 (N_9006,N_2447,N_912);
xor U9007 (N_9007,N_195,N_4807);
nand U9008 (N_9008,N_2630,N_2924);
or U9009 (N_9009,N_366,N_1551);
or U9010 (N_9010,N_390,N_1960);
and U9011 (N_9011,N_2768,N_1829);
nor U9012 (N_9012,N_3731,N_3241);
nor U9013 (N_9013,N_3565,N_3207);
and U9014 (N_9014,N_2621,N_1138);
or U9015 (N_9015,N_3606,N_3668);
xor U9016 (N_9016,N_3007,N_1127);
or U9017 (N_9017,N_461,N_229);
and U9018 (N_9018,N_268,N_955);
or U9019 (N_9019,N_1243,N_4577);
or U9020 (N_9020,N_4250,N_3403);
xor U9021 (N_9021,N_1590,N_1275);
or U9022 (N_9022,N_4682,N_2009);
nor U9023 (N_9023,N_821,N_142);
nor U9024 (N_9024,N_1994,N_3763);
or U9025 (N_9025,N_4768,N_4276);
xnor U9026 (N_9026,N_3070,N_4975);
nand U9027 (N_9027,N_961,N_3065);
xor U9028 (N_9028,N_4967,N_4414);
or U9029 (N_9029,N_3215,N_1056);
nand U9030 (N_9030,N_1689,N_2033);
and U9031 (N_9031,N_4217,N_497);
xnor U9032 (N_9032,N_2912,N_4702);
or U9033 (N_9033,N_1185,N_4204);
xor U9034 (N_9034,N_3705,N_2698);
nand U9035 (N_9035,N_4157,N_1698);
nor U9036 (N_9036,N_3663,N_1025);
and U9037 (N_9037,N_2411,N_3979);
and U9038 (N_9038,N_475,N_396);
nand U9039 (N_9039,N_367,N_1911);
and U9040 (N_9040,N_3399,N_1953);
xnor U9041 (N_9041,N_4635,N_294);
and U9042 (N_9042,N_2121,N_4149);
or U9043 (N_9043,N_4622,N_4294);
nand U9044 (N_9044,N_56,N_4894);
xnor U9045 (N_9045,N_3205,N_2007);
xor U9046 (N_9046,N_3355,N_2742);
nor U9047 (N_9047,N_733,N_2948);
nand U9048 (N_9048,N_545,N_355);
nand U9049 (N_9049,N_2470,N_4640);
nand U9050 (N_9050,N_2145,N_2701);
xor U9051 (N_9051,N_4861,N_4771);
or U9052 (N_9052,N_2327,N_355);
or U9053 (N_9053,N_2004,N_341);
nand U9054 (N_9054,N_4099,N_4811);
or U9055 (N_9055,N_2089,N_2272);
or U9056 (N_9056,N_3903,N_1603);
nor U9057 (N_9057,N_4717,N_2291);
xnor U9058 (N_9058,N_2296,N_1512);
or U9059 (N_9059,N_2234,N_4914);
xnor U9060 (N_9060,N_4077,N_1801);
or U9061 (N_9061,N_562,N_1118);
or U9062 (N_9062,N_575,N_3195);
and U9063 (N_9063,N_4825,N_4804);
nand U9064 (N_9064,N_2938,N_4552);
or U9065 (N_9065,N_1477,N_3333);
or U9066 (N_9066,N_4742,N_4061);
and U9067 (N_9067,N_1955,N_1783);
and U9068 (N_9068,N_1758,N_3927);
nor U9069 (N_9069,N_240,N_611);
xnor U9070 (N_9070,N_3346,N_3106);
nor U9071 (N_9071,N_2538,N_3502);
xor U9072 (N_9072,N_4478,N_1231);
xnor U9073 (N_9073,N_3645,N_3012);
and U9074 (N_9074,N_1310,N_4774);
and U9075 (N_9075,N_2946,N_3788);
and U9076 (N_9076,N_99,N_1507);
nand U9077 (N_9077,N_2514,N_1732);
nand U9078 (N_9078,N_2516,N_1094);
nand U9079 (N_9079,N_91,N_4614);
and U9080 (N_9080,N_3283,N_1341);
nor U9081 (N_9081,N_2451,N_2107);
xor U9082 (N_9082,N_3195,N_1566);
nand U9083 (N_9083,N_1231,N_239);
xnor U9084 (N_9084,N_3833,N_1107);
nand U9085 (N_9085,N_2177,N_1474);
xor U9086 (N_9086,N_3541,N_1428);
nand U9087 (N_9087,N_398,N_3397);
or U9088 (N_9088,N_794,N_4801);
xor U9089 (N_9089,N_3087,N_4909);
and U9090 (N_9090,N_4301,N_1546);
nor U9091 (N_9091,N_4117,N_2030);
or U9092 (N_9092,N_3954,N_4511);
nand U9093 (N_9093,N_525,N_2415);
nor U9094 (N_9094,N_3675,N_4234);
nand U9095 (N_9095,N_2258,N_1841);
nand U9096 (N_9096,N_687,N_296);
nand U9097 (N_9097,N_4813,N_219);
nor U9098 (N_9098,N_3047,N_3346);
xnor U9099 (N_9099,N_2360,N_859);
nand U9100 (N_9100,N_3982,N_2769);
xor U9101 (N_9101,N_2583,N_116);
nor U9102 (N_9102,N_3096,N_4125);
xnor U9103 (N_9103,N_70,N_748);
nand U9104 (N_9104,N_1572,N_3693);
xnor U9105 (N_9105,N_3051,N_4664);
nand U9106 (N_9106,N_1607,N_4479);
or U9107 (N_9107,N_3344,N_372);
nor U9108 (N_9108,N_3852,N_109);
xor U9109 (N_9109,N_3420,N_4724);
and U9110 (N_9110,N_3481,N_3166);
nand U9111 (N_9111,N_1195,N_2345);
and U9112 (N_9112,N_4841,N_4082);
or U9113 (N_9113,N_779,N_3582);
or U9114 (N_9114,N_3054,N_4111);
and U9115 (N_9115,N_1450,N_4777);
and U9116 (N_9116,N_79,N_987);
xnor U9117 (N_9117,N_2370,N_322);
xor U9118 (N_9118,N_2516,N_3531);
nand U9119 (N_9119,N_128,N_571);
nor U9120 (N_9120,N_994,N_2282);
xor U9121 (N_9121,N_3233,N_3092);
or U9122 (N_9122,N_4917,N_1350);
xor U9123 (N_9123,N_352,N_3475);
xor U9124 (N_9124,N_910,N_4617);
nor U9125 (N_9125,N_424,N_3507);
xor U9126 (N_9126,N_4514,N_1350);
or U9127 (N_9127,N_1282,N_3927);
nand U9128 (N_9128,N_2296,N_3777);
xnor U9129 (N_9129,N_1171,N_1887);
or U9130 (N_9130,N_4724,N_3820);
nor U9131 (N_9131,N_1663,N_959);
xor U9132 (N_9132,N_4074,N_1024);
nor U9133 (N_9133,N_4523,N_1300);
nand U9134 (N_9134,N_3277,N_3573);
nor U9135 (N_9135,N_709,N_3362);
and U9136 (N_9136,N_149,N_4162);
xnor U9137 (N_9137,N_2829,N_4283);
and U9138 (N_9138,N_342,N_931);
and U9139 (N_9139,N_2479,N_3719);
nor U9140 (N_9140,N_2545,N_3853);
xor U9141 (N_9141,N_4923,N_526);
nor U9142 (N_9142,N_1945,N_849);
nand U9143 (N_9143,N_1182,N_4274);
nor U9144 (N_9144,N_994,N_224);
or U9145 (N_9145,N_3388,N_4578);
nand U9146 (N_9146,N_170,N_3813);
nor U9147 (N_9147,N_4835,N_2991);
nor U9148 (N_9148,N_3964,N_2540);
nand U9149 (N_9149,N_1624,N_233);
nor U9150 (N_9150,N_4890,N_3297);
xor U9151 (N_9151,N_1632,N_888);
and U9152 (N_9152,N_834,N_3738);
nor U9153 (N_9153,N_833,N_2083);
nand U9154 (N_9154,N_4773,N_4120);
xor U9155 (N_9155,N_2776,N_4236);
and U9156 (N_9156,N_4473,N_2512);
xnor U9157 (N_9157,N_2323,N_3155);
nand U9158 (N_9158,N_4681,N_3029);
nand U9159 (N_9159,N_3976,N_1264);
nand U9160 (N_9160,N_2671,N_1048);
xor U9161 (N_9161,N_3702,N_1671);
nor U9162 (N_9162,N_4801,N_2198);
xor U9163 (N_9163,N_2692,N_2482);
and U9164 (N_9164,N_1266,N_4531);
and U9165 (N_9165,N_4969,N_375);
and U9166 (N_9166,N_3615,N_1885);
and U9167 (N_9167,N_1243,N_2534);
nand U9168 (N_9168,N_4247,N_2244);
and U9169 (N_9169,N_3742,N_1705);
nor U9170 (N_9170,N_1757,N_961);
or U9171 (N_9171,N_3111,N_1388);
nor U9172 (N_9172,N_2609,N_4280);
xnor U9173 (N_9173,N_4901,N_2667);
nand U9174 (N_9174,N_1305,N_1465);
nand U9175 (N_9175,N_1704,N_770);
xor U9176 (N_9176,N_491,N_4406);
and U9177 (N_9177,N_707,N_1724);
or U9178 (N_9178,N_1254,N_4641);
or U9179 (N_9179,N_3837,N_1882);
xnor U9180 (N_9180,N_3682,N_2761);
nand U9181 (N_9181,N_3461,N_4561);
and U9182 (N_9182,N_2110,N_4305);
and U9183 (N_9183,N_1242,N_1912);
xnor U9184 (N_9184,N_4389,N_2359);
or U9185 (N_9185,N_2051,N_4904);
and U9186 (N_9186,N_3385,N_1590);
and U9187 (N_9187,N_2715,N_3311);
and U9188 (N_9188,N_2724,N_2667);
nor U9189 (N_9189,N_754,N_62);
nor U9190 (N_9190,N_3402,N_3813);
and U9191 (N_9191,N_1948,N_3278);
nand U9192 (N_9192,N_2974,N_1569);
xor U9193 (N_9193,N_3377,N_1525);
nor U9194 (N_9194,N_1099,N_4913);
xnor U9195 (N_9195,N_3490,N_136);
and U9196 (N_9196,N_4587,N_3665);
nor U9197 (N_9197,N_3893,N_4157);
nor U9198 (N_9198,N_365,N_3387);
xnor U9199 (N_9199,N_1601,N_680);
nand U9200 (N_9200,N_4899,N_1057);
and U9201 (N_9201,N_2925,N_3760);
and U9202 (N_9202,N_928,N_954);
and U9203 (N_9203,N_4829,N_4474);
nand U9204 (N_9204,N_3895,N_4990);
xnor U9205 (N_9205,N_2825,N_3887);
and U9206 (N_9206,N_2728,N_1814);
nand U9207 (N_9207,N_2280,N_3556);
nand U9208 (N_9208,N_216,N_2129);
nor U9209 (N_9209,N_2564,N_4129);
and U9210 (N_9210,N_4820,N_1776);
nor U9211 (N_9211,N_141,N_842);
or U9212 (N_9212,N_848,N_3960);
nor U9213 (N_9213,N_3660,N_3260);
nand U9214 (N_9214,N_2852,N_4539);
xor U9215 (N_9215,N_931,N_3404);
or U9216 (N_9216,N_1767,N_433);
nor U9217 (N_9217,N_2727,N_240);
xor U9218 (N_9218,N_970,N_2292);
and U9219 (N_9219,N_2756,N_930);
nand U9220 (N_9220,N_2757,N_1173);
or U9221 (N_9221,N_3146,N_3880);
or U9222 (N_9222,N_4835,N_2085);
nor U9223 (N_9223,N_2069,N_2107);
and U9224 (N_9224,N_1828,N_1918);
nand U9225 (N_9225,N_4599,N_3596);
and U9226 (N_9226,N_4597,N_1601);
xnor U9227 (N_9227,N_3826,N_3303);
or U9228 (N_9228,N_3344,N_1560);
nor U9229 (N_9229,N_4112,N_3098);
nand U9230 (N_9230,N_2617,N_3811);
nor U9231 (N_9231,N_1175,N_2685);
xnor U9232 (N_9232,N_3168,N_4267);
nand U9233 (N_9233,N_1781,N_2907);
nand U9234 (N_9234,N_3218,N_2090);
xnor U9235 (N_9235,N_3209,N_4295);
nor U9236 (N_9236,N_4047,N_4511);
nor U9237 (N_9237,N_264,N_3638);
nand U9238 (N_9238,N_1351,N_432);
and U9239 (N_9239,N_1265,N_206);
nor U9240 (N_9240,N_1429,N_474);
nand U9241 (N_9241,N_596,N_2417);
and U9242 (N_9242,N_1471,N_4796);
xnor U9243 (N_9243,N_2075,N_231);
nand U9244 (N_9244,N_1383,N_4870);
or U9245 (N_9245,N_2170,N_3958);
nor U9246 (N_9246,N_2788,N_2584);
xnor U9247 (N_9247,N_562,N_759);
nand U9248 (N_9248,N_1333,N_4419);
xor U9249 (N_9249,N_1958,N_4592);
and U9250 (N_9250,N_3360,N_1718);
xnor U9251 (N_9251,N_199,N_193);
or U9252 (N_9252,N_4842,N_2546);
xor U9253 (N_9253,N_2513,N_3597);
xor U9254 (N_9254,N_2386,N_4562);
or U9255 (N_9255,N_62,N_4993);
xnor U9256 (N_9256,N_703,N_4168);
or U9257 (N_9257,N_2319,N_3770);
xor U9258 (N_9258,N_3255,N_2140);
nand U9259 (N_9259,N_3486,N_97);
and U9260 (N_9260,N_4270,N_378);
xnor U9261 (N_9261,N_1595,N_4153);
nand U9262 (N_9262,N_4710,N_1305);
and U9263 (N_9263,N_1303,N_2533);
nor U9264 (N_9264,N_4891,N_273);
xor U9265 (N_9265,N_3778,N_1861);
nor U9266 (N_9266,N_2161,N_4597);
nand U9267 (N_9267,N_1480,N_3471);
and U9268 (N_9268,N_2450,N_3348);
xor U9269 (N_9269,N_3276,N_4495);
nor U9270 (N_9270,N_2204,N_2119);
and U9271 (N_9271,N_3403,N_3167);
nor U9272 (N_9272,N_2701,N_1366);
nor U9273 (N_9273,N_2214,N_3451);
or U9274 (N_9274,N_3439,N_331);
or U9275 (N_9275,N_2673,N_1391);
and U9276 (N_9276,N_2218,N_4380);
nor U9277 (N_9277,N_4456,N_2591);
nor U9278 (N_9278,N_966,N_1699);
and U9279 (N_9279,N_943,N_2863);
or U9280 (N_9280,N_1683,N_2181);
and U9281 (N_9281,N_2362,N_1323);
nor U9282 (N_9282,N_2303,N_954);
and U9283 (N_9283,N_167,N_186);
nand U9284 (N_9284,N_3097,N_2875);
and U9285 (N_9285,N_3024,N_1120);
or U9286 (N_9286,N_365,N_1152);
or U9287 (N_9287,N_3044,N_4887);
xnor U9288 (N_9288,N_4264,N_4128);
nand U9289 (N_9289,N_3884,N_2867);
nand U9290 (N_9290,N_3050,N_3594);
xor U9291 (N_9291,N_511,N_2106);
or U9292 (N_9292,N_4769,N_3952);
or U9293 (N_9293,N_379,N_3381);
and U9294 (N_9294,N_329,N_393);
and U9295 (N_9295,N_2829,N_116);
xnor U9296 (N_9296,N_4009,N_3119);
nor U9297 (N_9297,N_528,N_3600);
xor U9298 (N_9298,N_3539,N_1505);
or U9299 (N_9299,N_1238,N_4639);
or U9300 (N_9300,N_4882,N_261);
nor U9301 (N_9301,N_1527,N_4122);
nor U9302 (N_9302,N_0,N_572);
nand U9303 (N_9303,N_2792,N_3389);
nand U9304 (N_9304,N_2161,N_3592);
xnor U9305 (N_9305,N_1255,N_2281);
and U9306 (N_9306,N_1322,N_1669);
xnor U9307 (N_9307,N_2796,N_4086);
nor U9308 (N_9308,N_673,N_4940);
nand U9309 (N_9309,N_2422,N_1186);
xor U9310 (N_9310,N_3975,N_2291);
xnor U9311 (N_9311,N_63,N_825);
or U9312 (N_9312,N_3929,N_4038);
nor U9313 (N_9313,N_4084,N_2874);
or U9314 (N_9314,N_2689,N_3763);
nand U9315 (N_9315,N_33,N_3855);
or U9316 (N_9316,N_1195,N_2663);
nor U9317 (N_9317,N_2842,N_3808);
or U9318 (N_9318,N_3897,N_2775);
or U9319 (N_9319,N_200,N_4926);
xnor U9320 (N_9320,N_2282,N_3801);
and U9321 (N_9321,N_601,N_4121);
nand U9322 (N_9322,N_4947,N_1525);
nand U9323 (N_9323,N_4829,N_623);
nand U9324 (N_9324,N_2193,N_1642);
and U9325 (N_9325,N_672,N_1855);
xor U9326 (N_9326,N_1263,N_1464);
nand U9327 (N_9327,N_1241,N_960);
xnor U9328 (N_9328,N_3545,N_2431);
and U9329 (N_9329,N_3894,N_873);
and U9330 (N_9330,N_128,N_4072);
and U9331 (N_9331,N_665,N_2504);
or U9332 (N_9332,N_1711,N_3940);
and U9333 (N_9333,N_1354,N_2441);
or U9334 (N_9334,N_3463,N_2290);
or U9335 (N_9335,N_1837,N_1961);
or U9336 (N_9336,N_2599,N_3345);
and U9337 (N_9337,N_188,N_1222);
nor U9338 (N_9338,N_66,N_1479);
nor U9339 (N_9339,N_1202,N_4495);
xor U9340 (N_9340,N_2435,N_4747);
and U9341 (N_9341,N_4456,N_1301);
nor U9342 (N_9342,N_2184,N_2482);
or U9343 (N_9343,N_2693,N_2959);
nand U9344 (N_9344,N_1292,N_3874);
nor U9345 (N_9345,N_3471,N_1987);
nand U9346 (N_9346,N_713,N_4758);
xor U9347 (N_9347,N_4958,N_4531);
nand U9348 (N_9348,N_3777,N_979);
xor U9349 (N_9349,N_1106,N_568);
and U9350 (N_9350,N_4641,N_387);
and U9351 (N_9351,N_4952,N_1134);
nand U9352 (N_9352,N_3709,N_3042);
xnor U9353 (N_9353,N_1524,N_4962);
nand U9354 (N_9354,N_4403,N_551);
or U9355 (N_9355,N_3893,N_510);
nor U9356 (N_9356,N_3610,N_4721);
and U9357 (N_9357,N_4466,N_3269);
and U9358 (N_9358,N_415,N_3578);
nor U9359 (N_9359,N_3720,N_2037);
or U9360 (N_9360,N_1140,N_4403);
or U9361 (N_9361,N_372,N_4513);
nor U9362 (N_9362,N_2241,N_4295);
and U9363 (N_9363,N_4887,N_2604);
and U9364 (N_9364,N_1858,N_3371);
or U9365 (N_9365,N_2857,N_1140);
or U9366 (N_9366,N_1100,N_4636);
and U9367 (N_9367,N_830,N_2900);
and U9368 (N_9368,N_4613,N_3889);
nor U9369 (N_9369,N_625,N_4253);
or U9370 (N_9370,N_1924,N_3348);
nor U9371 (N_9371,N_611,N_4647);
or U9372 (N_9372,N_1097,N_2700);
or U9373 (N_9373,N_836,N_4493);
nor U9374 (N_9374,N_3830,N_858);
nor U9375 (N_9375,N_4469,N_3819);
and U9376 (N_9376,N_4650,N_2833);
nor U9377 (N_9377,N_1695,N_2816);
and U9378 (N_9378,N_3558,N_2531);
or U9379 (N_9379,N_9,N_1717);
nand U9380 (N_9380,N_555,N_439);
and U9381 (N_9381,N_16,N_3514);
or U9382 (N_9382,N_4332,N_1450);
or U9383 (N_9383,N_4733,N_1019);
nor U9384 (N_9384,N_4618,N_3774);
xor U9385 (N_9385,N_769,N_2378);
and U9386 (N_9386,N_2935,N_2702);
xor U9387 (N_9387,N_4926,N_2513);
xor U9388 (N_9388,N_2662,N_4282);
and U9389 (N_9389,N_3713,N_4857);
xnor U9390 (N_9390,N_2769,N_962);
xor U9391 (N_9391,N_2731,N_2643);
xnor U9392 (N_9392,N_3383,N_1941);
nor U9393 (N_9393,N_1308,N_380);
or U9394 (N_9394,N_3357,N_968);
nand U9395 (N_9395,N_4291,N_3314);
and U9396 (N_9396,N_1330,N_3617);
nor U9397 (N_9397,N_142,N_2949);
nor U9398 (N_9398,N_1165,N_4947);
or U9399 (N_9399,N_2028,N_964);
xor U9400 (N_9400,N_1031,N_4536);
nand U9401 (N_9401,N_4344,N_3023);
and U9402 (N_9402,N_4141,N_3521);
nand U9403 (N_9403,N_2222,N_4834);
nand U9404 (N_9404,N_1745,N_4358);
nor U9405 (N_9405,N_695,N_1253);
or U9406 (N_9406,N_4268,N_1792);
and U9407 (N_9407,N_2216,N_733);
nand U9408 (N_9408,N_3979,N_1382);
xor U9409 (N_9409,N_2897,N_4026);
xor U9410 (N_9410,N_3982,N_3185);
nor U9411 (N_9411,N_978,N_4530);
nand U9412 (N_9412,N_3182,N_4779);
and U9413 (N_9413,N_2708,N_4207);
nand U9414 (N_9414,N_2718,N_2425);
or U9415 (N_9415,N_626,N_4633);
or U9416 (N_9416,N_3329,N_2370);
xnor U9417 (N_9417,N_4359,N_1636);
nor U9418 (N_9418,N_874,N_4760);
xor U9419 (N_9419,N_3880,N_4629);
nor U9420 (N_9420,N_502,N_771);
nor U9421 (N_9421,N_3496,N_4032);
nor U9422 (N_9422,N_1533,N_1236);
nand U9423 (N_9423,N_442,N_291);
or U9424 (N_9424,N_233,N_1197);
nand U9425 (N_9425,N_1982,N_83);
nand U9426 (N_9426,N_3071,N_910);
nand U9427 (N_9427,N_3575,N_61);
xnor U9428 (N_9428,N_4875,N_649);
or U9429 (N_9429,N_952,N_2191);
nor U9430 (N_9430,N_4553,N_619);
xor U9431 (N_9431,N_2262,N_3588);
or U9432 (N_9432,N_1685,N_3700);
nand U9433 (N_9433,N_4400,N_2674);
xnor U9434 (N_9434,N_2324,N_4541);
or U9435 (N_9435,N_2189,N_2259);
nand U9436 (N_9436,N_775,N_1122);
nand U9437 (N_9437,N_26,N_388);
nand U9438 (N_9438,N_1469,N_2670);
or U9439 (N_9439,N_1803,N_3034);
and U9440 (N_9440,N_3334,N_1295);
and U9441 (N_9441,N_1969,N_574);
and U9442 (N_9442,N_1545,N_1166);
and U9443 (N_9443,N_4498,N_4329);
and U9444 (N_9444,N_2415,N_3286);
nor U9445 (N_9445,N_4088,N_747);
xor U9446 (N_9446,N_3501,N_3704);
and U9447 (N_9447,N_3972,N_963);
nor U9448 (N_9448,N_4113,N_1045);
xnor U9449 (N_9449,N_395,N_3522);
or U9450 (N_9450,N_2411,N_2871);
nand U9451 (N_9451,N_2978,N_1469);
or U9452 (N_9452,N_4405,N_3044);
nand U9453 (N_9453,N_3531,N_1976);
nand U9454 (N_9454,N_3695,N_3552);
nor U9455 (N_9455,N_4025,N_2077);
or U9456 (N_9456,N_806,N_473);
nor U9457 (N_9457,N_1942,N_4256);
nor U9458 (N_9458,N_1577,N_1840);
or U9459 (N_9459,N_3927,N_3226);
or U9460 (N_9460,N_3469,N_1453);
and U9461 (N_9461,N_4830,N_321);
and U9462 (N_9462,N_4426,N_1927);
or U9463 (N_9463,N_4479,N_2346);
nor U9464 (N_9464,N_1959,N_4489);
nor U9465 (N_9465,N_1778,N_1427);
and U9466 (N_9466,N_1751,N_1421);
and U9467 (N_9467,N_2830,N_4688);
nor U9468 (N_9468,N_519,N_1769);
or U9469 (N_9469,N_2221,N_3654);
nand U9470 (N_9470,N_3825,N_875);
nand U9471 (N_9471,N_2654,N_3407);
nor U9472 (N_9472,N_1030,N_3509);
and U9473 (N_9473,N_3667,N_726);
and U9474 (N_9474,N_4214,N_2272);
nor U9475 (N_9475,N_2763,N_3940);
xnor U9476 (N_9476,N_4509,N_3183);
nor U9477 (N_9477,N_1657,N_4257);
or U9478 (N_9478,N_1335,N_1372);
nor U9479 (N_9479,N_4343,N_4633);
nor U9480 (N_9480,N_2544,N_4555);
nand U9481 (N_9481,N_236,N_984);
nand U9482 (N_9482,N_3042,N_1321);
xor U9483 (N_9483,N_1199,N_3353);
or U9484 (N_9484,N_506,N_4343);
xor U9485 (N_9485,N_4281,N_2372);
and U9486 (N_9486,N_3541,N_2758);
xor U9487 (N_9487,N_4180,N_1020);
or U9488 (N_9488,N_1581,N_1452);
nor U9489 (N_9489,N_1932,N_3615);
and U9490 (N_9490,N_2135,N_1822);
nor U9491 (N_9491,N_3840,N_955);
nor U9492 (N_9492,N_4264,N_1598);
and U9493 (N_9493,N_1026,N_2446);
xor U9494 (N_9494,N_1216,N_4695);
or U9495 (N_9495,N_1045,N_107);
nor U9496 (N_9496,N_3092,N_3531);
nand U9497 (N_9497,N_3285,N_1063);
or U9498 (N_9498,N_1189,N_2556);
and U9499 (N_9499,N_4515,N_3605);
xor U9500 (N_9500,N_650,N_1016);
nor U9501 (N_9501,N_3091,N_2889);
nand U9502 (N_9502,N_2604,N_442);
nand U9503 (N_9503,N_656,N_1168);
nand U9504 (N_9504,N_391,N_1828);
or U9505 (N_9505,N_4558,N_4553);
nor U9506 (N_9506,N_4592,N_2506);
and U9507 (N_9507,N_3275,N_830);
and U9508 (N_9508,N_649,N_3056);
nor U9509 (N_9509,N_4790,N_1923);
nor U9510 (N_9510,N_1625,N_1391);
or U9511 (N_9511,N_3934,N_2961);
nor U9512 (N_9512,N_581,N_481);
nand U9513 (N_9513,N_3676,N_414);
or U9514 (N_9514,N_4853,N_565);
and U9515 (N_9515,N_4113,N_3607);
or U9516 (N_9516,N_1513,N_260);
or U9517 (N_9517,N_4286,N_367);
xnor U9518 (N_9518,N_3458,N_4574);
nand U9519 (N_9519,N_3797,N_875);
nor U9520 (N_9520,N_635,N_237);
and U9521 (N_9521,N_4636,N_4556);
and U9522 (N_9522,N_4516,N_4381);
xnor U9523 (N_9523,N_1289,N_846);
nor U9524 (N_9524,N_758,N_4244);
and U9525 (N_9525,N_1122,N_2218);
nand U9526 (N_9526,N_1694,N_805);
or U9527 (N_9527,N_1940,N_4280);
nand U9528 (N_9528,N_2043,N_999);
and U9529 (N_9529,N_3148,N_2592);
nor U9530 (N_9530,N_3227,N_3537);
nor U9531 (N_9531,N_4021,N_2681);
and U9532 (N_9532,N_383,N_1277);
and U9533 (N_9533,N_2884,N_2573);
and U9534 (N_9534,N_1666,N_726);
nand U9535 (N_9535,N_2521,N_3188);
xor U9536 (N_9536,N_3677,N_16);
or U9537 (N_9537,N_1238,N_4408);
nand U9538 (N_9538,N_1627,N_204);
nand U9539 (N_9539,N_823,N_2387);
nor U9540 (N_9540,N_1142,N_3207);
and U9541 (N_9541,N_2122,N_4000);
nor U9542 (N_9542,N_3196,N_348);
nor U9543 (N_9543,N_177,N_4326);
xnor U9544 (N_9544,N_1663,N_992);
xnor U9545 (N_9545,N_3924,N_4847);
xor U9546 (N_9546,N_3857,N_402);
nand U9547 (N_9547,N_3698,N_3843);
and U9548 (N_9548,N_3469,N_4450);
or U9549 (N_9549,N_1783,N_4580);
and U9550 (N_9550,N_2697,N_4226);
nand U9551 (N_9551,N_2702,N_3921);
nor U9552 (N_9552,N_3654,N_3908);
nand U9553 (N_9553,N_2559,N_1970);
and U9554 (N_9554,N_2300,N_1975);
and U9555 (N_9555,N_1633,N_1905);
or U9556 (N_9556,N_990,N_2704);
nand U9557 (N_9557,N_2193,N_1872);
xnor U9558 (N_9558,N_3088,N_4528);
nand U9559 (N_9559,N_3965,N_2686);
nor U9560 (N_9560,N_1238,N_3794);
nor U9561 (N_9561,N_2689,N_3131);
or U9562 (N_9562,N_952,N_1420);
and U9563 (N_9563,N_2824,N_208);
and U9564 (N_9564,N_4249,N_3067);
and U9565 (N_9565,N_1036,N_3071);
nor U9566 (N_9566,N_2710,N_1845);
xnor U9567 (N_9567,N_2856,N_4816);
nor U9568 (N_9568,N_1971,N_2530);
xnor U9569 (N_9569,N_3874,N_4678);
and U9570 (N_9570,N_1224,N_1687);
nand U9571 (N_9571,N_3928,N_585);
xnor U9572 (N_9572,N_4749,N_1074);
nor U9573 (N_9573,N_3021,N_3399);
and U9574 (N_9574,N_3594,N_4211);
xor U9575 (N_9575,N_1775,N_3862);
nand U9576 (N_9576,N_18,N_3202);
or U9577 (N_9577,N_4731,N_167);
and U9578 (N_9578,N_4067,N_980);
xor U9579 (N_9579,N_9,N_4865);
and U9580 (N_9580,N_211,N_4);
xor U9581 (N_9581,N_4184,N_3926);
or U9582 (N_9582,N_3236,N_2957);
or U9583 (N_9583,N_2532,N_566);
and U9584 (N_9584,N_3565,N_3032);
nor U9585 (N_9585,N_491,N_4171);
and U9586 (N_9586,N_782,N_4444);
xor U9587 (N_9587,N_1225,N_433);
or U9588 (N_9588,N_1154,N_1974);
nand U9589 (N_9589,N_872,N_2344);
nand U9590 (N_9590,N_961,N_3088);
nor U9591 (N_9591,N_1372,N_1019);
nand U9592 (N_9592,N_3025,N_2702);
nand U9593 (N_9593,N_4628,N_765);
xnor U9594 (N_9594,N_4476,N_740);
nor U9595 (N_9595,N_1294,N_2107);
xor U9596 (N_9596,N_387,N_1277);
xnor U9597 (N_9597,N_3134,N_2104);
nand U9598 (N_9598,N_399,N_4963);
and U9599 (N_9599,N_531,N_922);
nor U9600 (N_9600,N_4014,N_4472);
nand U9601 (N_9601,N_298,N_1213);
and U9602 (N_9602,N_2151,N_3397);
nand U9603 (N_9603,N_29,N_68);
nor U9604 (N_9604,N_1337,N_2474);
and U9605 (N_9605,N_1632,N_4388);
nor U9606 (N_9606,N_1262,N_4206);
or U9607 (N_9607,N_1985,N_394);
or U9608 (N_9608,N_189,N_1654);
nor U9609 (N_9609,N_3452,N_3165);
nor U9610 (N_9610,N_2910,N_2296);
and U9611 (N_9611,N_4838,N_1103);
or U9612 (N_9612,N_3913,N_4473);
xor U9613 (N_9613,N_730,N_2105);
and U9614 (N_9614,N_629,N_517);
and U9615 (N_9615,N_3837,N_2713);
nand U9616 (N_9616,N_3518,N_4148);
xor U9617 (N_9617,N_2877,N_3005);
nor U9618 (N_9618,N_4956,N_4802);
xor U9619 (N_9619,N_1722,N_3039);
nor U9620 (N_9620,N_2587,N_1692);
xor U9621 (N_9621,N_1266,N_3799);
or U9622 (N_9622,N_1102,N_4979);
xnor U9623 (N_9623,N_4816,N_4717);
xnor U9624 (N_9624,N_3688,N_673);
xor U9625 (N_9625,N_1688,N_2161);
xnor U9626 (N_9626,N_3000,N_2043);
and U9627 (N_9627,N_1993,N_4163);
or U9628 (N_9628,N_80,N_2969);
and U9629 (N_9629,N_87,N_3183);
xnor U9630 (N_9630,N_2032,N_2871);
or U9631 (N_9631,N_2719,N_2534);
nand U9632 (N_9632,N_1786,N_1029);
nor U9633 (N_9633,N_2668,N_1184);
and U9634 (N_9634,N_4145,N_4481);
xnor U9635 (N_9635,N_2299,N_896);
or U9636 (N_9636,N_236,N_2316);
nand U9637 (N_9637,N_4800,N_2085);
nor U9638 (N_9638,N_907,N_4100);
nand U9639 (N_9639,N_4696,N_3681);
and U9640 (N_9640,N_1396,N_4677);
and U9641 (N_9641,N_2998,N_728);
or U9642 (N_9642,N_4538,N_3791);
and U9643 (N_9643,N_1087,N_1526);
nand U9644 (N_9644,N_3189,N_3630);
xnor U9645 (N_9645,N_559,N_201);
or U9646 (N_9646,N_3343,N_4172);
nor U9647 (N_9647,N_3506,N_4299);
xnor U9648 (N_9648,N_2815,N_1147);
nand U9649 (N_9649,N_849,N_617);
nor U9650 (N_9650,N_2375,N_3692);
and U9651 (N_9651,N_639,N_1912);
nand U9652 (N_9652,N_4589,N_3207);
nor U9653 (N_9653,N_4110,N_3395);
and U9654 (N_9654,N_893,N_4898);
or U9655 (N_9655,N_3153,N_1506);
xnor U9656 (N_9656,N_2860,N_2374);
and U9657 (N_9657,N_3259,N_2898);
xor U9658 (N_9658,N_668,N_1984);
xnor U9659 (N_9659,N_632,N_1965);
xnor U9660 (N_9660,N_351,N_36);
xor U9661 (N_9661,N_3313,N_4491);
and U9662 (N_9662,N_1791,N_2567);
xor U9663 (N_9663,N_1206,N_4286);
and U9664 (N_9664,N_1455,N_1841);
or U9665 (N_9665,N_3572,N_332);
nor U9666 (N_9666,N_578,N_1398);
nand U9667 (N_9667,N_3280,N_4029);
nor U9668 (N_9668,N_4200,N_750);
xor U9669 (N_9669,N_4055,N_3884);
and U9670 (N_9670,N_541,N_4753);
nand U9671 (N_9671,N_4610,N_705);
and U9672 (N_9672,N_278,N_69);
and U9673 (N_9673,N_280,N_1581);
nor U9674 (N_9674,N_1533,N_30);
nand U9675 (N_9675,N_2513,N_1285);
nand U9676 (N_9676,N_654,N_4305);
or U9677 (N_9677,N_1137,N_698);
and U9678 (N_9678,N_3978,N_3210);
nand U9679 (N_9679,N_4317,N_3246);
and U9680 (N_9680,N_4366,N_3363);
nor U9681 (N_9681,N_2481,N_1841);
nor U9682 (N_9682,N_2779,N_907);
nor U9683 (N_9683,N_560,N_4222);
xnor U9684 (N_9684,N_2528,N_3063);
nor U9685 (N_9685,N_716,N_3376);
nand U9686 (N_9686,N_2982,N_1241);
and U9687 (N_9687,N_1395,N_4871);
nor U9688 (N_9688,N_907,N_3949);
nor U9689 (N_9689,N_1909,N_3353);
nor U9690 (N_9690,N_931,N_4875);
or U9691 (N_9691,N_189,N_1962);
and U9692 (N_9692,N_4073,N_2508);
nand U9693 (N_9693,N_3113,N_2217);
xnor U9694 (N_9694,N_1515,N_1837);
nand U9695 (N_9695,N_177,N_3435);
nor U9696 (N_9696,N_1023,N_189);
nor U9697 (N_9697,N_1484,N_4281);
xor U9698 (N_9698,N_3596,N_1660);
or U9699 (N_9699,N_4595,N_3919);
xor U9700 (N_9700,N_2164,N_2830);
nor U9701 (N_9701,N_4404,N_2153);
and U9702 (N_9702,N_3674,N_665);
xor U9703 (N_9703,N_4821,N_3167);
and U9704 (N_9704,N_1077,N_2104);
nor U9705 (N_9705,N_4975,N_2635);
xor U9706 (N_9706,N_1793,N_193);
or U9707 (N_9707,N_2219,N_4788);
xor U9708 (N_9708,N_4278,N_2938);
and U9709 (N_9709,N_3840,N_1441);
nand U9710 (N_9710,N_3549,N_4352);
and U9711 (N_9711,N_1649,N_4501);
nor U9712 (N_9712,N_668,N_1060);
xnor U9713 (N_9713,N_4528,N_2202);
nand U9714 (N_9714,N_4858,N_939);
and U9715 (N_9715,N_4301,N_1740);
and U9716 (N_9716,N_1308,N_1682);
and U9717 (N_9717,N_4807,N_1408);
xor U9718 (N_9718,N_627,N_3593);
xnor U9719 (N_9719,N_755,N_3540);
nor U9720 (N_9720,N_2105,N_711);
xor U9721 (N_9721,N_4726,N_3171);
xnor U9722 (N_9722,N_3115,N_1802);
xor U9723 (N_9723,N_3605,N_759);
nor U9724 (N_9724,N_3491,N_2043);
nand U9725 (N_9725,N_2637,N_4852);
nor U9726 (N_9726,N_1865,N_2778);
and U9727 (N_9727,N_2551,N_2754);
or U9728 (N_9728,N_1597,N_907);
xnor U9729 (N_9729,N_1315,N_1907);
and U9730 (N_9730,N_1269,N_3086);
or U9731 (N_9731,N_2000,N_4180);
nor U9732 (N_9732,N_2203,N_4328);
nand U9733 (N_9733,N_4457,N_4024);
xnor U9734 (N_9734,N_3654,N_2705);
or U9735 (N_9735,N_2630,N_2678);
xor U9736 (N_9736,N_1845,N_369);
nand U9737 (N_9737,N_2570,N_4861);
xor U9738 (N_9738,N_4445,N_4517);
nor U9739 (N_9739,N_2262,N_2234);
nor U9740 (N_9740,N_1769,N_1245);
xor U9741 (N_9741,N_4299,N_2230);
or U9742 (N_9742,N_4829,N_1634);
xor U9743 (N_9743,N_579,N_2423);
nor U9744 (N_9744,N_2067,N_871);
and U9745 (N_9745,N_3456,N_128);
or U9746 (N_9746,N_3425,N_262);
and U9747 (N_9747,N_3221,N_1787);
and U9748 (N_9748,N_3785,N_273);
nand U9749 (N_9749,N_4624,N_1597);
nand U9750 (N_9750,N_4373,N_4287);
nand U9751 (N_9751,N_2567,N_4);
nor U9752 (N_9752,N_4075,N_1448);
xor U9753 (N_9753,N_4087,N_3751);
xor U9754 (N_9754,N_4195,N_1118);
or U9755 (N_9755,N_3908,N_988);
and U9756 (N_9756,N_1956,N_3386);
nand U9757 (N_9757,N_1648,N_2837);
nor U9758 (N_9758,N_662,N_1147);
xor U9759 (N_9759,N_4553,N_1157);
xor U9760 (N_9760,N_1850,N_4678);
or U9761 (N_9761,N_16,N_3548);
or U9762 (N_9762,N_552,N_3164);
or U9763 (N_9763,N_4550,N_2965);
nand U9764 (N_9764,N_4754,N_2217);
xnor U9765 (N_9765,N_4396,N_1282);
or U9766 (N_9766,N_1723,N_1553);
nand U9767 (N_9767,N_4822,N_53);
or U9768 (N_9768,N_2043,N_2739);
nor U9769 (N_9769,N_3819,N_1649);
xnor U9770 (N_9770,N_2811,N_1574);
or U9771 (N_9771,N_3143,N_1899);
xor U9772 (N_9772,N_513,N_2039);
nor U9773 (N_9773,N_4698,N_1170);
nor U9774 (N_9774,N_3668,N_1932);
xor U9775 (N_9775,N_299,N_1277);
nand U9776 (N_9776,N_4324,N_3131);
and U9777 (N_9777,N_2927,N_3272);
and U9778 (N_9778,N_4722,N_2423);
xor U9779 (N_9779,N_4085,N_1600);
nand U9780 (N_9780,N_3624,N_3103);
and U9781 (N_9781,N_2293,N_4503);
and U9782 (N_9782,N_3904,N_497);
xnor U9783 (N_9783,N_3571,N_2747);
xnor U9784 (N_9784,N_712,N_4972);
and U9785 (N_9785,N_2578,N_1511);
or U9786 (N_9786,N_4356,N_2245);
xnor U9787 (N_9787,N_1092,N_629);
xnor U9788 (N_9788,N_4141,N_899);
and U9789 (N_9789,N_367,N_4519);
or U9790 (N_9790,N_754,N_3811);
xor U9791 (N_9791,N_794,N_3593);
or U9792 (N_9792,N_3711,N_4047);
or U9793 (N_9793,N_1954,N_4063);
and U9794 (N_9794,N_4226,N_175);
xor U9795 (N_9795,N_382,N_3678);
nand U9796 (N_9796,N_1393,N_1125);
nand U9797 (N_9797,N_693,N_4823);
nor U9798 (N_9798,N_2228,N_4108);
and U9799 (N_9799,N_1954,N_504);
nor U9800 (N_9800,N_2259,N_4378);
nand U9801 (N_9801,N_724,N_122);
nor U9802 (N_9802,N_4908,N_3064);
and U9803 (N_9803,N_1353,N_3475);
nor U9804 (N_9804,N_3045,N_3757);
xor U9805 (N_9805,N_2472,N_4173);
or U9806 (N_9806,N_2451,N_2324);
and U9807 (N_9807,N_4821,N_2208);
or U9808 (N_9808,N_2678,N_1977);
xor U9809 (N_9809,N_1502,N_2097);
nor U9810 (N_9810,N_519,N_4308);
nand U9811 (N_9811,N_264,N_254);
nor U9812 (N_9812,N_4831,N_2577);
nor U9813 (N_9813,N_1470,N_889);
or U9814 (N_9814,N_722,N_4254);
and U9815 (N_9815,N_2144,N_2706);
nand U9816 (N_9816,N_3211,N_861);
nand U9817 (N_9817,N_866,N_1572);
and U9818 (N_9818,N_2597,N_4824);
xnor U9819 (N_9819,N_4984,N_2625);
nor U9820 (N_9820,N_2285,N_3444);
and U9821 (N_9821,N_149,N_1487);
or U9822 (N_9822,N_4956,N_3307);
and U9823 (N_9823,N_53,N_1968);
xnor U9824 (N_9824,N_1046,N_500);
or U9825 (N_9825,N_3442,N_4612);
xnor U9826 (N_9826,N_3758,N_1881);
xnor U9827 (N_9827,N_705,N_3841);
and U9828 (N_9828,N_547,N_118);
or U9829 (N_9829,N_850,N_2577);
and U9830 (N_9830,N_1553,N_2478);
nand U9831 (N_9831,N_2029,N_3320);
and U9832 (N_9832,N_4547,N_140);
nor U9833 (N_9833,N_898,N_2318);
and U9834 (N_9834,N_2570,N_3400);
xor U9835 (N_9835,N_1630,N_4627);
xor U9836 (N_9836,N_1867,N_4471);
and U9837 (N_9837,N_1036,N_2407);
nor U9838 (N_9838,N_2215,N_2479);
or U9839 (N_9839,N_3920,N_3992);
nand U9840 (N_9840,N_4624,N_2752);
nor U9841 (N_9841,N_1965,N_2193);
or U9842 (N_9842,N_3843,N_579);
or U9843 (N_9843,N_1067,N_3148);
xnor U9844 (N_9844,N_1657,N_141);
xnor U9845 (N_9845,N_3798,N_115);
xnor U9846 (N_9846,N_552,N_539);
nor U9847 (N_9847,N_2194,N_1490);
and U9848 (N_9848,N_664,N_1905);
nand U9849 (N_9849,N_4625,N_2144);
xnor U9850 (N_9850,N_1498,N_885);
xnor U9851 (N_9851,N_1217,N_2);
nand U9852 (N_9852,N_2767,N_4969);
and U9853 (N_9853,N_4852,N_979);
or U9854 (N_9854,N_3134,N_4731);
or U9855 (N_9855,N_4695,N_3850);
nor U9856 (N_9856,N_3003,N_1689);
nand U9857 (N_9857,N_3272,N_3767);
or U9858 (N_9858,N_2112,N_858);
and U9859 (N_9859,N_555,N_1379);
nand U9860 (N_9860,N_1216,N_440);
and U9861 (N_9861,N_3890,N_2354);
nor U9862 (N_9862,N_1596,N_4269);
and U9863 (N_9863,N_4526,N_1034);
or U9864 (N_9864,N_2935,N_1435);
and U9865 (N_9865,N_1759,N_1479);
or U9866 (N_9866,N_2499,N_1524);
or U9867 (N_9867,N_1170,N_3121);
or U9868 (N_9868,N_1514,N_472);
and U9869 (N_9869,N_3772,N_415);
nor U9870 (N_9870,N_676,N_2495);
and U9871 (N_9871,N_516,N_4838);
nand U9872 (N_9872,N_4001,N_1140);
nor U9873 (N_9873,N_3556,N_3085);
and U9874 (N_9874,N_2083,N_4846);
xnor U9875 (N_9875,N_4451,N_308);
xor U9876 (N_9876,N_1263,N_2537);
and U9877 (N_9877,N_1165,N_52);
or U9878 (N_9878,N_1551,N_427);
and U9879 (N_9879,N_334,N_1808);
nor U9880 (N_9880,N_1635,N_4549);
xnor U9881 (N_9881,N_2109,N_459);
nand U9882 (N_9882,N_3958,N_997);
or U9883 (N_9883,N_3264,N_4360);
nand U9884 (N_9884,N_1769,N_4362);
nor U9885 (N_9885,N_4984,N_1160);
xnor U9886 (N_9886,N_38,N_940);
xor U9887 (N_9887,N_3434,N_3356);
nand U9888 (N_9888,N_3514,N_3026);
nor U9889 (N_9889,N_375,N_450);
or U9890 (N_9890,N_2214,N_4635);
nand U9891 (N_9891,N_4918,N_2016);
or U9892 (N_9892,N_4419,N_140);
and U9893 (N_9893,N_768,N_3886);
nand U9894 (N_9894,N_3108,N_2261);
nor U9895 (N_9895,N_135,N_2896);
nor U9896 (N_9896,N_4487,N_4414);
and U9897 (N_9897,N_2812,N_1613);
nor U9898 (N_9898,N_4451,N_3121);
xnor U9899 (N_9899,N_1055,N_3280);
or U9900 (N_9900,N_3145,N_1787);
and U9901 (N_9901,N_2775,N_919);
nand U9902 (N_9902,N_2369,N_4459);
xor U9903 (N_9903,N_3041,N_2917);
xnor U9904 (N_9904,N_4580,N_1638);
nand U9905 (N_9905,N_2476,N_377);
nor U9906 (N_9906,N_4128,N_2458);
xor U9907 (N_9907,N_2966,N_3028);
nand U9908 (N_9908,N_1735,N_3370);
xor U9909 (N_9909,N_125,N_2735);
nor U9910 (N_9910,N_2310,N_521);
and U9911 (N_9911,N_4852,N_1927);
xnor U9912 (N_9912,N_671,N_2531);
or U9913 (N_9913,N_2965,N_1132);
or U9914 (N_9914,N_65,N_3866);
or U9915 (N_9915,N_2975,N_2178);
or U9916 (N_9916,N_3279,N_1906);
nor U9917 (N_9917,N_4191,N_1331);
or U9918 (N_9918,N_4342,N_3636);
nand U9919 (N_9919,N_3044,N_3359);
xnor U9920 (N_9920,N_316,N_1609);
or U9921 (N_9921,N_3130,N_2538);
nor U9922 (N_9922,N_1410,N_1193);
and U9923 (N_9923,N_3344,N_2064);
nor U9924 (N_9924,N_1465,N_3697);
xor U9925 (N_9925,N_320,N_232);
nor U9926 (N_9926,N_784,N_3723);
xnor U9927 (N_9927,N_242,N_2076);
nor U9928 (N_9928,N_3794,N_1484);
xnor U9929 (N_9929,N_3545,N_4700);
and U9930 (N_9930,N_3568,N_3454);
or U9931 (N_9931,N_2253,N_966);
and U9932 (N_9932,N_628,N_2096);
xor U9933 (N_9933,N_756,N_4629);
or U9934 (N_9934,N_3643,N_2203);
or U9935 (N_9935,N_1081,N_4259);
or U9936 (N_9936,N_1172,N_2675);
nor U9937 (N_9937,N_2950,N_3949);
xnor U9938 (N_9938,N_4594,N_2576);
xor U9939 (N_9939,N_323,N_2405);
xnor U9940 (N_9940,N_4661,N_2911);
xnor U9941 (N_9941,N_4663,N_3253);
or U9942 (N_9942,N_1504,N_210);
nor U9943 (N_9943,N_3051,N_4372);
or U9944 (N_9944,N_3802,N_4962);
or U9945 (N_9945,N_2459,N_2326);
or U9946 (N_9946,N_2809,N_4484);
nand U9947 (N_9947,N_4230,N_4049);
nor U9948 (N_9948,N_251,N_2643);
nor U9949 (N_9949,N_2111,N_3440);
xor U9950 (N_9950,N_2994,N_4177);
nor U9951 (N_9951,N_3883,N_3768);
and U9952 (N_9952,N_3377,N_2298);
and U9953 (N_9953,N_4058,N_4388);
nand U9954 (N_9954,N_1917,N_1596);
and U9955 (N_9955,N_4913,N_182);
xor U9956 (N_9956,N_1788,N_2760);
nand U9957 (N_9957,N_170,N_427);
xor U9958 (N_9958,N_415,N_1460);
nand U9959 (N_9959,N_1406,N_4284);
nand U9960 (N_9960,N_1436,N_3255);
nor U9961 (N_9961,N_406,N_484);
and U9962 (N_9962,N_935,N_1429);
nor U9963 (N_9963,N_4782,N_4448);
nand U9964 (N_9964,N_4823,N_4518);
and U9965 (N_9965,N_1364,N_1492);
or U9966 (N_9966,N_78,N_3038);
nor U9967 (N_9967,N_779,N_1129);
xnor U9968 (N_9968,N_1362,N_3457);
nand U9969 (N_9969,N_889,N_4826);
nand U9970 (N_9970,N_1663,N_4041);
nand U9971 (N_9971,N_3558,N_3592);
xor U9972 (N_9972,N_443,N_4229);
or U9973 (N_9973,N_919,N_3426);
nor U9974 (N_9974,N_3526,N_1145);
xor U9975 (N_9975,N_4257,N_1681);
nand U9976 (N_9976,N_3953,N_2248);
nand U9977 (N_9977,N_2467,N_2343);
nand U9978 (N_9978,N_2301,N_4896);
xnor U9979 (N_9979,N_3063,N_3793);
or U9980 (N_9980,N_889,N_4791);
xnor U9981 (N_9981,N_4216,N_2572);
and U9982 (N_9982,N_3967,N_1278);
and U9983 (N_9983,N_1581,N_3540);
or U9984 (N_9984,N_942,N_1837);
or U9985 (N_9985,N_113,N_4363);
nand U9986 (N_9986,N_450,N_366);
xor U9987 (N_9987,N_3793,N_668);
and U9988 (N_9988,N_576,N_4512);
nor U9989 (N_9989,N_746,N_3834);
xnor U9990 (N_9990,N_162,N_1019);
or U9991 (N_9991,N_1743,N_2264);
nand U9992 (N_9992,N_2588,N_3213);
or U9993 (N_9993,N_207,N_2076);
nor U9994 (N_9994,N_950,N_1586);
xor U9995 (N_9995,N_485,N_4893);
xnor U9996 (N_9996,N_4843,N_3145);
and U9997 (N_9997,N_1208,N_1377);
and U9998 (N_9998,N_937,N_2849);
nand U9999 (N_9999,N_683,N_3367);
nor U10000 (N_10000,N_8380,N_6840);
xnor U10001 (N_10001,N_8790,N_8822);
nor U10002 (N_10002,N_5770,N_7548);
xnor U10003 (N_10003,N_5208,N_7907);
or U10004 (N_10004,N_8053,N_9992);
nor U10005 (N_10005,N_6888,N_7282);
xor U10006 (N_10006,N_7817,N_5954);
nor U10007 (N_10007,N_6619,N_5532);
or U10008 (N_10008,N_8404,N_7797);
nand U10009 (N_10009,N_9418,N_6300);
nand U10010 (N_10010,N_8757,N_8217);
xnor U10011 (N_10011,N_6392,N_6009);
or U10012 (N_10012,N_6088,N_6360);
and U10013 (N_10013,N_9402,N_8664);
or U10014 (N_10014,N_8670,N_8958);
or U10015 (N_10015,N_5299,N_5167);
nand U10016 (N_10016,N_9535,N_6509);
xnor U10017 (N_10017,N_5408,N_7026);
and U10018 (N_10018,N_8525,N_8538);
nor U10019 (N_10019,N_9729,N_7179);
xnor U10020 (N_10020,N_6158,N_8581);
xnor U10021 (N_10021,N_8470,N_9682);
xnor U10022 (N_10022,N_5572,N_5022);
nand U10023 (N_10023,N_6689,N_5336);
nand U10024 (N_10024,N_5628,N_9398);
xor U10025 (N_10025,N_5907,N_8554);
or U10026 (N_10026,N_9605,N_7618);
xor U10027 (N_10027,N_6257,N_7075);
or U10028 (N_10028,N_7219,N_8441);
nand U10029 (N_10029,N_8916,N_8335);
or U10030 (N_10030,N_9561,N_9886);
xnor U10031 (N_10031,N_7284,N_9872);
or U10032 (N_10032,N_7128,N_8620);
and U10033 (N_10033,N_9056,N_6377);
nand U10034 (N_10034,N_8704,N_9028);
nand U10035 (N_10035,N_5874,N_5079);
nand U10036 (N_10036,N_9227,N_9728);
xor U10037 (N_10037,N_9599,N_9437);
or U10038 (N_10038,N_8980,N_5311);
nor U10039 (N_10039,N_8678,N_5718);
or U10040 (N_10040,N_9410,N_8370);
or U10041 (N_10041,N_8676,N_5287);
nand U10042 (N_10042,N_9249,N_8329);
xor U10043 (N_10043,N_7714,N_5065);
nor U10044 (N_10044,N_5788,N_8289);
nand U10045 (N_10045,N_5465,N_6708);
and U10046 (N_10046,N_8641,N_8383);
and U10047 (N_10047,N_5649,N_7207);
or U10048 (N_10048,N_7815,N_9280);
and U10049 (N_10049,N_5577,N_6670);
or U10050 (N_10050,N_5966,N_6780);
nand U10051 (N_10051,N_6108,N_8523);
or U10052 (N_10052,N_5400,N_6215);
or U10053 (N_10053,N_7793,N_9826);
xor U10054 (N_10054,N_5710,N_8096);
nor U10055 (N_10055,N_6900,N_8362);
and U10056 (N_10056,N_7305,N_5075);
or U10057 (N_10057,N_6191,N_5840);
nand U10058 (N_10058,N_7098,N_6250);
xnor U10059 (N_10059,N_9669,N_7007);
nand U10060 (N_10060,N_6731,N_9295);
xnor U10061 (N_10061,N_8331,N_6967);
nor U10062 (N_10062,N_5895,N_9604);
nand U10063 (N_10063,N_8020,N_5187);
and U10064 (N_10064,N_6289,N_7575);
and U10065 (N_10065,N_7978,N_5963);
or U10066 (N_10066,N_9825,N_9404);
and U10067 (N_10067,N_8386,N_6334);
nor U10068 (N_10068,N_9797,N_6928);
nor U10069 (N_10069,N_6415,N_5561);
and U10070 (N_10070,N_6968,N_7140);
nand U10071 (N_10071,N_5137,N_7346);
xnor U10072 (N_10072,N_7250,N_8048);
xnor U10073 (N_10073,N_8593,N_7807);
and U10074 (N_10074,N_8268,N_9470);
nor U10075 (N_10075,N_9222,N_6362);
and U10076 (N_10076,N_7821,N_5391);
nor U10077 (N_10077,N_7615,N_7393);
nand U10078 (N_10078,N_5986,N_7425);
xnor U10079 (N_10079,N_9548,N_9677);
nand U10080 (N_10080,N_5251,N_6342);
and U10081 (N_10081,N_8439,N_5571);
xnor U10082 (N_10082,N_7735,N_5358);
nand U10083 (N_10083,N_9043,N_5588);
xor U10084 (N_10084,N_9676,N_9247);
and U10085 (N_10085,N_9477,N_6638);
or U10086 (N_10086,N_6839,N_5162);
nor U10087 (N_10087,N_5712,N_5598);
nor U10088 (N_10088,N_9897,N_6806);
xor U10089 (N_10089,N_8662,N_7625);
nand U10090 (N_10090,N_5186,N_9325);
and U10091 (N_10091,N_8208,N_5270);
xor U10092 (N_10092,N_6858,N_8011);
and U10093 (N_10093,N_7656,N_8021);
or U10094 (N_10094,N_9187,N_6917);
nor U10095 (N_10095,N_7660,N_8953);
nand U10096 (N_10096,N_5988,N_9721);
and U10097 (N_10097,N_5846,N_5460);
nor U10098 (N_10098,N_9851,N_8865);
and U10099 (N_10099,N_9357,N_8827);
and U10100 (N_10100,N_9817,N_9667);
and U10101 (N_10101,N_5584,N_5979);
or U10102 (N_10102,N_9920,N_5488);
xnor U10103 (N_10103,N_6425,N_8834);
and U10104 (N_10104,N_9626,N_7016);
xnor U10105 (N_10105,N_7668,N_6786);
or U10106 (N_10106,N_5158,N_5139);
and U10107 (N_10107,N_9930,N_7171);
xor U10108 (N_10108,N_6869,N_9313);
nor U10109 (N_10109,N_9756,N_9948);
and U10110 (N_10110,N_7164,N_7791);
or U10111 (N_10111,N_5323,N_7475);
nor U10112 (N_10112,N_5604,N_7780);
or U10113 (N_10113,N_9552,N_9146);
nand U10114 (N_10114,N_9838,N_8241);
nand U10115 (N_10115,N_7205,N_9617);
xnor U10116 (N_10116,N_5884,N_9068);
and U10117 (N_10117,N_6284,N_5789);
and U10118 (N_10118,N_5906,N_8852);
nor U10119 (N_10119,N_7375,N_8438);
xnor U10120 (N_10120,N_7311,N_7972);
xor U10121 (N_10121,N_7199,N_7535);
nor U10122 (N_10122,N_8556,N_7161);
nor U10123 (N_10123,N_6441,N_9935);
nor U10124 (N_10124,N_5790,N_9931);
or U10125 (N_10125,N_9478,N_9686);
nor U10126 (N_10126,N_8680,N_8218);
or U10127 (N_10127,N_6700,N_7872);
xnor U10128 (N_10128,N_6402,N_6676);
nand U10129 (N_10129,N_7921,N_9842);
and U10130 (N_10130,N_8823,N_8326);
or U10131 (N_10131,N_9607,N_5839);
xnor U10132 (N_10132,N_9451,N_8826);
or U10133 (N_10133,N_9815,N_5175);
and U10134 (N_10134,N_9081,N_6624);
or U10135 (N_10135,N_9377,N_8191);
nor U10136 (N_10136,N_9112,N_6678);
nor U10137 (N_10137,N_5854,N_8759);
nand U10138 (N_10138,N_8901,N_7290);
xor U10139 (N_10139,N_5934,N_5672);
nand U10140 (N_10140,N_9957,N_5084);
or U10141 (N_10141,N_5289,N_7953);
nor U10142 (N_10142,N_7019,N_6397);
nand U10143 (N_10143,N_9009,N_6329);
nand U10144 (N_10144,N_6593,N_8687);
or U10145 (N_10145,N_8754,N_7722);
xnor U10146 (N_10146,N_5638,N_8491);
xor U10147 (N_10147,N_6372,N_9016);
and U10148 (N_10148,N_5953,N_7035);
and U10149 (N_10149,N_9782,N_5001);
xor U10150 (N_10150,N_7958,N_5977);
and U10151 (N_10151,N_6517,N_9228);
or U10152 (N_10152,N_7810,N_6081);
and U10153 (N_10153,N_7686,N_7530);
or U10154 (N_10154,N_5087,N_6683);
nand U10155 (N_10155,N_5544,N_7288);
and U10156 (N_10156,N_8600,N_9496);
nor U10157 (N_10157,N_5467,N_5096);
xor U10158 (N_10158,N_5616,N_5030);
nor U10159 (N_10159,N_9840,N_7312);
nor U10160 (N_10160,N_7915,N_5292);
nor U10161 (N_10161,N_5935,N_7983);
and U10162 (N_10162,N_7929,N_9964);
and U10163 (N_10163,N_5601,N_8044);
xnor U10164 (N_10164,N_6395,N_9621);
nand U10165 (N_10165,N_9196,N_9639);
or U10166 (N_10166,N_8084,N_6757);
nor U10167 (N_10167,N_9987,N_9201);
or U10168 (N_10168,N_9271,N_5700);
and U10169 (N_10169,N_9002,N_6137);
and U10170 (N_10170,N_8494,N_8574);
nand U10171 (N_10171,N_9775,N_5782);
and U10172 (N_10172,N_5837,N_8057);
or U10173 (N_10173,N_6396,N_6281);
nor U10174 (N_10174,N_7144,N_9902);
or U10175 (N_10175,N_7976,N_5395);
xnor U10176 (N_10176,N_6063,N_8774);
or U10177 (N_10177,N_8213,N_7188);
nor U10178 (N_10178,N_5719,N_6556);
or U10179 (N_10179,N_5160,N_8462);
nand U10180 (N_10180,N_9681,N_5181);
nor U10181 (N_10181,N_6115,N_6553);
nand U10182 (N_10182,N_8292,N_5836);
nand U10183 (N_10183,N_7471,N_8710);
or U10184 (N_10184,N_6829,N_9864);
and U10185 (N_10185,N_9951,N_5301);
nor U10186 (N_10186,N_6138,N_7294);
nand U10187 (N_10187,N_6304,N_5249);
or U10188 (N_10188,N_6253,N_7458);
nand U10189 (N_10189,N_8016,N_5842);
and U10190 (N_10190,N_5855,N_7707);
or U10191 (N_10191,N_7020,N_8226);
nand U10192 (N_10192,N_6637,N_5606);
or U10193 (N_10193,N_7120,N_7598);
or U10194 (N_10194,N_5178,N_9556);
and U10195 (N_10195,N_9571,N_7118);
xnor U10196 (N_10196,N_9356,N_6561);
nor U10197 (N_10197,N_8260,N_6594);
nor U10198 (N_10198,N_6419,N_9905);
and U10199 (N_10199,N_6958,N_9481);
nor U10200 (N_10200,N_5548,N_9113);
and U10201 (N_10201,N_5123,N_8863);
nor U10202 (N_10202,N_8925,N_6827);
and U10203 (N_10203,N_7671,N_8755);
nand U10204 (N_10204,N_7524,N_7998);
or U10205 (N_10205,N_6587,N_7452);
nor U10206 (N_10206,N_9743,N_7612);
nor U10207 (N_10207,N_9455,N_5576);
xnor U10208 (N_10208,N_9395,N_5747);
nor U10209 (N_10209,N_7884,N_7110);
and U10210 (N_10210,N_8460,N_6429);
nand U10211 (N_10211,N_7741,N_8220);
or U10212 (N_10212,N_5316,N_8327);
xnor U10213 (N_10213,N_9171,N_7012);
and U10214 (N_10214,N_8839,N_9521);
xor U10215 (N_10215,N_8584,N_8536);
nor U10216 (N_10216,N_8406,N_8747);
nor U10217 (N_10217,N_9968,N_8229);
nand U10218 (N_10218,N_5511,N_8874);
or U10219 (N_10219,N_9433,N_6243);
nand U10220 (N_10220,N_5558,N_7163);
nand U10221 (N_10221,N_9877,N_9204);
nand U10222 (N_10222,N_7608,N_7562);
and U10223 (N_10223,N_8291,N_5482);
and U10224 (N_10224,N_6686,N_5889);
nand U10225 (N_10225,N_7003,N_9869);
nor U10226 (N_10226,N_6764,N_8777);
nand U10227 (N_10227,N_8199,N_8959);
nand U10228 (N_10228,N_7627,N_8847);
xor U10229 (N_10229,N_5148,N_8789);
or U10230 (N_10230,N_5019,N_5680);
xnor U10231 (N_10231,N_7057,N_9709);
xor U10232 (N_10232,N_8845,N_6297);
xnor U10233 (N_10233,N_9543,N_7119);
or U10234 (N_10234,N_6992,N_9381);
nand U10235 (N_10235,N_5063,N_6994);
xor U10236 (N_10236,N_8635,N_7935);
xor U10237 (N_10237,N_5784,N_9760);
nor U10238 (N_10238,N_7034,N_9727);
nand U10239 (N_10239,N_9367,N_6262);
xnor U10240 (N_10240,N_8436,N_5626);
nand U10241 (N_10241,N_5157,N_7240);
nand U10242 (N_10242,N_6655,N_5695);
nor U10243 (N_10243,N_6142,N_8012);
or U10244 (N_10244,N_6523,N_7400);
and U10245 (N_10245,N_9324,N_9053);
and U10246 (N_10246,N_8764,N_5972);
xor U10247 (N_10247,N_5248,N_9576);
nand U10248 (N_10248,N_6633,N_5361);
and U10249 (N_10249,N_6707,N_6622);
and U10250 (N_10250,N_8187,N_6332);
and U10251 (N_10251,N_5430,N_5639);
nor U10252 (N_10252,N_7637,N_8806);
xnor U10253 (N_10253,N_6811,N_6971);
and U10254 (N_10254,N_6046,N_7088);
nor U10255 (N_10255,N_8809,N_7512);
or U10256 (N_10256,N_5283,N_7537);
and U10257 (N_10257,N_6939,N_7977);
or U10258 (N_10258,N_6251,N_9730);
nor U10259 (N_10259,N_9716,N_6812);
and U10260 (N_10260,N_6563,N_7480);
and U10261 (N_10261,N_8745,N_7715);
nand U10262 (N_10262,N_5863,N_9278);
xnor U10263 (N_10263,N_7508,N_7158);
nor U10264 (N_10264,N_6154,N_6493);
nor U10265 (N_10265,N_7823,N_8989);
nand U10266 (N_10266,N_7439,N_8132);
nor U10267 (N_10267,N_5504,N_9189);
nor U10268 (N_10268,N_8749,N_7669);
or U10269 (N_10269,N_6628,N_6436);
xnor U10270 (N_10270,N_8587,N_5374);
nor U10271 (N_10271,N_5827,N_6223);
xor U10272 (N_10272,N_7401,N_8591);
nor U10273 (N_10273,N_7518,N_5013);
or U10274 (N_10274,N_7385,N_8829);
and U10275 (N_10275,N_8937,N_7261);
nor U10276 (N_10276,N_9944,N_5468);
nand U10277 (N_10277,N_6100,N_7061);
nor U10278 (N_10278,N_9579,N_8379);
nor U10279 (N_10279,N_7028,N_9061);
and U10280 (N_10280,N_9966,N_9591);
or U10281 (N_10281,N_5521,N_5915);
nor U10282 (N_10282,N_8243,N_9215);
or U10283 (N_10283,N_6354,N_6501);
nand U10284 (N_10284,N_9906,N_7619);
nor U10285 (N_10285,N_9005,N_9103);
nor U10286 (N_10286,N_7113,N_6042);
nand U10287 (N_10287,N_9630,N_6179);
and U10288 (N_10288,N_8571,N_8624);
xor U10289 (N_10289,N_5871,N_6011);
nor U10290 (N_10290,N_8776,N_9387);
or U10291 (N_10291,N_5797,N_8286);
or U10292 (N_10292,N_6428,N_8008);
nand U10293 (N_10293,N_8341,N_8803);
or U10294 (N_10294,N_5097,N_8899);
xnor U10295 (N_10295,N_7853,N_7310);
or U10296 (N_10296,N_7990,N_9823);
nor U10297 (N_10297,N_9658,N_6082);
or U10298 (N_10298,N_7326,N_5480);
nor U10299 (N_10299,N_9441,N_8089);
nor U10300 (N_10300,N_9491,N_7071);
nand U10301 (N_10301,N_8186,N_7177);
nor U10302 (N_10302,N_9703,N_9965);
or U10303 (N_10303,N_8824,N_7336);
nand U10304 (N_10304,N_7325,N_8878);
and U10305 (N_10305,N_5851,N_9394);
nor U10306 (N_10306,N_5849,N_7556);
or U10307 (N_10307,N_5968,N_6296);
or U10308 (N_10308,N_9655,N_7916);
and U10309 (N_10309,N_5918,N_5241);
xnor U10310 (N_10310,N_8079,N_7763);
and U10311 (N_10311,N_6386,N_6791);
and U10312 (N_10312,N_5751,N_5763);
and U10313 (N_10313,N_9495,N_8318);
or U10314 (N_10314,N_5004,N_5727);
and U10315 (N_10315,N_5082,N_6906);
and U10316 (N_10316,N_9391,N_7804);
xnor U10317 (N_10317,N_9693,N_9542);
or U10318 (N_10318,N_9058,N_5039);
or U10319 (N_10319,N_9925,N_9546);
nand U10320 (N_10320,N_6538,N_7221);
xnor U10321 (N_10321,N_7526,N_6631);
nand U10322 (N_10322,N_7355,N_6452);
xor U10323 (N_10323,N_7868,N_9408);
or U10324 (N_10324,N_8009,N_7382);
xnor U10325 (N_10325,N_9590,N_9265);
nor U10326 (N_10326,N_6815,N_7504);
nand U10327 (N_10327,N_8744,N_9534);
nor U10328 (N_10328,N_8760,N_5742);
nor U10329 (N_10329,N_7755,N_8039);
and U10330 (N_10330,N_6564,N_6673);
nand U10331 (N_10331,N_9134,N_9997);
nand U10332 (N_10332,N_8434,N_8312);
nand U10333 (N_10333,N_9035,N_8139);
nand U10334 (N_10334,N_9190,N_9638);
and U10335 (N_10335,N_8631,N_5144);
xor U10336 (N_10336,N_9123,N_8511);
nor U10337 (N_10337,N_8787,N_8842);
and U10338 (N_10338,N_8940,N_9124);
and U10339 (N_10339,N_6210,N_9326);
xor U10340 (N_10340,N_5134,N_6615);
and U10341 (N_10341,N_9973,N_5565);
or U10342 (N_10342,N_9240,N_9268);
and U10343 (N_10343,N_6865,N_7431);
xor U10344 (N_10344,N_5961,N_6636);
and U10345 (N_10345,N_5666,N_9528);
and U10346 (N_10346,N_8604,N_5103);
nand U10347 (N_10347,N_5335,N_9142);
xnor U10348 (N_10348,N_8815,N_6008);
and U10349 (N_10349,N_5982,N_6677);
nor U10350 (N_10350,N_7954,N_6504);
nand U10351 (N_10351,N_9233,N_5886);
and U10352 (N_10352,N_5017,N_7022);
and U10353 (N_10353,N_8773,N_5586);
and U10354 (N_10354,N_9132,N_8973);
nand U10355 (N_10355,N_7209,N_8515);
nand U10356 (N_10356,N_9878,N_9798);
or U10357 (N_10357,N_6028,N_8877);
or U10358 (N_10358,N_5791,N_9555);
nor U10359 (N_10359,N_6241,N_5706);
or U10360 (N_10360,N_8282,N_5517);
xnor U10361 (N_10361,N_6198,N_8814);
and U10362 (N_10362,N_9487,N_7636);
xor U10363 (N_10363,N_9656,N_6902);
or U10364 (N_10364,N_7457,N_7067);
and U10365 (N_10365,N_7383,N_5232);
or U10366 (N_10366,N_8168,N_9619);
and U10367 (N_10367,N_5984,N_7441);
nor U10368 (N_10368,N_9919,N_8982);
nand U10369 (N_10369,N_9041,N_7453);
or U10370 (N_10370,N_9095,N_8443);
nor U10371 (N_10371,N_6111,N_8337);
xnor U10372 (N_10372,N_5707,N_6398);
or U10373 (N_10373,N_5636,N_5414);
nand U10374 (N_10374,N_9629,N_5766);
and U10375 (N_10375,N_9346,N_7011);
or U10376 (N_10376,N_9067,N_6098);
nor U10377 (N_10377,N_5050,N_8231);
nand U10378 (N_10378,N_6752,N_5403);
nor U10379 (N_10379,N_9033,N_7850);
and U10380 (N_10380,N_7278,N_6792);
xnor U10381 (N_10381,N_8601,N_7581);
and U10382 (N_10382,N_5833,N_8529);
and U10383 (N_10383,N_6454,N_5266);
nand U10384 (N_10384,N_5673,N_9400);
or U10385 (N_10385,N_5624,N_9500);
xor U10386 (N_10386,N_6139,N_9810);
or U10387 (N_10387,N_8553,N_6176);
or U10388 (N_10388,N_5217,N_8647);
xnor U10389 (N_10389,N_6560,N_8728);
nand U10390 (N_10390,N_7690,N_9744);
nand U10391 (N_10391,N_6592,N_5225);
or U10392 (N_10392,N_5860,N_5904);
xor U10393 (N_10393,N_6531,N_5685);
nand U10394 (N_10394,N_7952,N_9014);
xor U10395 (N_10395,N_5177,N_8461);
nor U10396 (N_10396,N_7316,N_5101);
xnor U10397 (N_10397,N_9623,N_5730);
xnor U10398 (N_10398,N_9642,N_5545);
or U10399 (N_10399,N_9585,N_8446);
nor U10400 (N_10400,N_6189,N_9737);
and U10401 (N_10401,N_7839,N_6227);
xnor U10402 (N_10402,N_8724,N_8017);
nor U10403 (N_10403,N_7046,N_8128);
or U10404 (N_10404,N_5112,N_7376);
nand U10405 (N_10405,N_8851,N_5912);
xor U10406 (N_10406,N_9209,N_8264);
or U10407 (N_10407,N_5092,N_8224);
or U10408 (N_10408,N_7031,N_7942);
nand U10409 (N_10409,N_8705,N_8146);
nor U10410 (N_10410,N_8873,N_8975);
nand U10411 (N_10411,N_9996,N_5411);
or U10412 (N_10412,N_8393,N_8120);
xor U10413 (N_10413,N_9723,N_8875);
nor U10414 (N_10414,N_5002,N_7579);
nor U10415 (N_10415,N_6263,N_6051);
xor U10416 (N_10416,N_6199,N_7354);
xnor U10417 (N_10417,N_5524,N_7476);
nand U10418 (N_10418,N_7647,N_7111);
and U10419 (N_10419,N_9694,N_8907);
or U10420 (N_10420,N_8816,N_8590);
nor U10421 (N_10421,N_5776,N_6303);
nand U10422 (N_10422,N_6266,N_8746);
nor U10423 (N_10423,N_9051,N_7837);
nand U10424 (N_10424,N_5526,N_5145);
nor U10425 (N_10425,N_5992,N_6864);
nor U10426 (N_10426,N_8317,N_9490);
xor U10427 (N_10427,N_9958,N_7744);
nor U10428 (N_10428,N_7474,N_8950);
and U10429 (N_10429,N_6554,N_9045);
nor U10430 (N_10430,N_6382,N_6358);
and U10431 (N_10431,N_6846,N_5007);
nor U10432 (N_10432,N_9863,N_7836);
and U10433 (N_10433,N_5332,N_5568);
nand U10434 (N_10434,N_6106,N_9494);
nand U10435 (N_10435,N_8606,N_8636);
nor U10436 (N_10436,N_7591,N_7115);
nor U10437 (N_10437,N_6935,N_6848);
and U10438 (N_10438,N_5341,N_8459);
or U10439 (N_10439,N_6077,N_9547);
nand U10440 (N_10440,N_7352,N_9763);
xor U10441 (N_10441,N_6724,N_6110);
and U10442 (N_10442,N_7033,N_5748);
and U10443 (N_10443,N_5683,N_6370);
nor U10444 (N_10444,N_8962,N_5542);
or U10445 (N_10445,N_6907,N_8941);
xor U10446 (N_10446,N_5515,N_6188);
nor U10447 (N_10447,N_8495,N_7831);
or U10448 (N_10448,N_6163,N_9953);
or U10449 (N_10449,N_8963,N_8643);
and U10450 (N_10450,N_6671,N_5473);
xor U10451 (N_10451,N_6129,N_7249);
and U10452 (N_10452,N_6357,N_7693);
nand U10453 (N_10453,N_8285,N_7613);
xor U10454 (N_10454,N_6299,N_6507);
nor U10455 (N_10455,N_9019,N_7961);
or U10456 (N_10456,N_8060,N_9509);
or U10457 (N_10457,N_5057,N_5888);
xnor U10458 (N_10458,N_8463,N_8752);
xnor U10459 (N_10459,N_8732,N_9063);
or U10460 (N_10460,N_7538,N_8129);
and U10461 (N_10461,N_6173,N_5893);
and U10462 (N_10462,N_9211,N_6799);
and U10463 (N_10463,N_7975,N_9169);
xor U10464 (N_10464,N_8485,N_8274);
nor U10465 (N_10465,N_8788,N_8293);
nor U10466 (N_10466,N_5668,N_5599);
nor U10467 (N_10467,N_5061,N_6252);
xor U10468 (N_10468,N_7795,N_6793);
nor U10469 (N_10469,N_5099,N_9162);
and U10470 (N_10470,N_7265,N_8930);
nor U10471 (N_10471,N_8339,N_7877);
nand U10472 (N_10472,N_6889,N_6713);
nand U10473 (N_10473,N_9801,N_8180);
xnor U10474 (N_10474,N_8345,N_9382);
nor U10475 (N_10475,N_7677,N_9978);
nor U10476 (N_10476,N_6659,N_5294);
nor U10477 (N_10477,N_8683,N_5136);
and U10478 (N_10478,N_9786,N_9753);
xor U10479 (N_10479,N_9833,N_8792);
nor U10480 (N_10480,N_5664,N_5218);
or U10481 (N_10481,N_6908,N_8482);
or U10482 (N_10482,N_8425,N_9334);
xnor U10483 (N_10483,N_5792,N_7396);
or U10484 (N_10484,N_6978,N_7074);
or U10485 (N_10485,N_7124,N_5607);
and U10486 (N_10486,N_5052,N_8905);
nand U10487 (N_10487,N_5416,N_9632);
and U10488 (N_10488,N_5901,N_7014);
xnor U10489 (N_10489,N_6852,N_8548);
xor U10490 (N_10490,N_9595,N_5350);
and U10491 (N_10491,N_7967,N_6083);
xor U10492 (N_10492,N_6071,N_9237);
xor U10493 (N_10493,N_5987,N_7883);
and U10494 (N_10494,N_8052,N_6144);
nor U10495 (N_10495,N_6784,N_6998);
xnor U10496 (N_10496,N_6438,N_8104);
nor U10497 (N_10497,N_8521,N_7230);
nor U10498 (N_10498,N_6127,N_9331);
or U10499 (N_10499,N_6503,N_6738);
or U10500 (N_10500,N_6762,N_5941);
and U10501 (N_10501,N_7748,N_5040);
nand U10502 (N_10502,N_8691,N_6647);
nor U10503 (N_10503,N_7679,N_6414);
nand U10504 (N_10504,N_9572,N_8546);
nor U10505 (N_10505,N_7800,N_5042);
nand U10506 (N_10506,N_7648,N_5786);
nor U10507 (N_10507,N_5062,N_7938);
and U10508 (N_10508,N_6001,N_6514);
nand U10509 (N_10509,N_8219,N_7782);
or U10510 (N_10510,N_6751,N_6663);
nand U10511 (N_10511,N_5366,N_9484);
nor U10512 (N_10512,N_5298,N_9274);
nor U10513 (N_10513,N_6794,N_7826);
nand U10514 (N_10514,N_8568,N_7495);
or U10515 (N_10515,N_7469,N_6043);
nor U10516 (N_10516,N_7085,N_8420);
or U10517 (N_10517,N_5243,N_7814);
nor U10518 (N_10518,N_9865,N_7281);
nor U10519 (N_10519,N_7805,N_8684);
xnor U10520 (N_10520,N_9940,N_8682);
nand U10521 (N_10521,N_5194,N_5307);
xnor U10522 (N_10522,N_6055,N_5155);
and U10523 (N_10523,N_9154,N_6817);
xor U10524 (N_10524,N_5739,N_5206);
xor U10525 (N_10525,N_7835,N_9119);
and U10526 (N_10526,N_9309,N_5894);
xor U10527 (N_10527,N_8265,N_8444);
xnor U10528 (N_10528,N_5592,N_6448);
xor U10529 (N_10529,N_6838,N_8184);
xnor U10530 (N_10530,N_7890,N_9868);
nor U10531 (N_10531,N_5031,N_6851);
or U10532 (N_10532,N_5005,N_5920);
nor U10533 (N_10533,N_7684,N_9554);
or U10534 (N_10534,N_6029,N_7180);
nor U10535 (N_10535,N_6006,N_6416);
nand U10536 (N_10536,N_8209,N_8621);
nand U10537 (N_10537,N_7499,N_6091);
xnor U10538 (N_10538,N_5993,N_8701);
and U10539 (N_10539,N_8313,N_6513);
and U10540 (N_10540,N_9994,N_9910);
nand U10541 (N_10541,N_6828,N_6373);
nor U10542 (N_10542,N_6172,N_6349);
nor U10543 (N_10543,N_9017,N_7747);
xor U10544 (N_10544,N_6524,N_9185);
nand U10545 (N_10545,N_6875,N_9164);
nor U10546 (N_10546,N_9194,N_6720);
nand U10547 (N_10547,N_8835,N_5246);
nand U10548 (N_10548,N_7030,N_9022);
xnor U10549 (N_10549,N_7824,N_9615);
xnor U10550 (N_10550,N_7298,N_6528);
or U10551 (N_10551,N_5463,N_5320);
or U10552 (N_10552,N_5038,N_7910);
or U10553 (N_10553,N_8758,N_6401);
nor U10554 (N_10554,N_6393,N_5487);
nand U10555 (N_10555,N_5367,N_5098);
nor U10556 (N_10556,N_6213,N_9533);
or U10557 (N_10557,N_6455,N_7332);
xnor U10558 (N_10558,N_5975,N_5753);
or U10559 (N_10559,N_6474,N_9421);
or U10560 (N_10560,N_6087,N_6976);
and U10561 (N_10561,N_7214,N_6116);
and U10562 (N_10562,N_7198,N_8185);
and U10563 (N_10563,N_9405,N_6430);
nor U10564 (N_10564,N_5852,N_7367);
xnor U10565 (N_10565,N_9255,N_7979);
or U10566 (N_10566,N_5254,N_7216);
nand U10567 (N_10567,N_9225,N_9903);
nor U10568 (N_10568,N_6383,N_5551);
nor U10569 (N_10569,N_8879,N_8113);
nor U10570 (N_10570,N_8500,N_6599);
and U10571 (N_10571,N_6530,N_6291);
xor U10572 (N_10572,N_7699,N_8440);
or U10573 (N_10573,N_7750,N_6337);
and U10574 (N_10574,N_6118,N_8967);
and U10575 (N_10575,N_6535,N_9999);
or U10576 (N_10576,N_6874,N_5365);
nor U10577 (N_10577,N_5094,N_7484);
and U10578 (N_10578,N_8435,N_9202);
nand U10579 (N_10579,N_7918,N_5612);
xor U10580 (N_10580,N_5522,N_6672);
and U10581 (N_10581,N_6178,N_7479);
or U10582 (N_10582,N_9483,N_9724);
nand U10583 (N_10583,N_5552,N_8942);
and U10584 (N_10584,N_9597,N_7387);
nor U10585 (N_10585,N_5644,N_5581);
xnor U10586 (N_10586,N_7503,N_9462);
and U10587 (N_10587,N_6201,N_6771);
nor U10588 (N_10588,N_7082,N_8427);
nor U10589 (N_10589,N_9269,N_7516);
or U10590 (N_10590,N_7949,N_8706);
xnor U10591 (N_10591,N_7399,N_7462);
and U10592 (N_10592,N_8614,N_6944);
and U10593 (N_10593,N_8449,N_8262);
nor U10594 (N_10594,N_9922,N_5856);
nand U10595 (N_10595,N_6305,N_6748);
and U10596 (N_10596,N_8333,N_9963);
or U10597 (N_10597,N_9563,N_6855);
and U10598 (N_10598,N_5227,N_9795);
or U10599 (N_10599,N_8657,N_7010);
and U10600 (N_10600,N_8041,N_5962);
or U10601 (N_10601,N_7673,N_7483);
or U10602 (N_10602,N_6997,N_9811);
nor U10603 (N_10603,N_7076,N_8650);
nand U10604 (N_10604,N_9504,N_6461);
xnor U10605 (N_10605,N_7774,N_8098);
or U10606 (N_10606,N_7752,N_5441);
nor U10607 (N_10607,N_5721,N_7390);
or U10608 (N_10608,N_8848,N_6192);
nor U10609 (N_10609,N_9784,N_8530);
and U10610 (N_10610,N_5076,N_8368);
or U10611 (N_10611,N_7342,N_6140);
nor U10612 (N_10612,N_5969,N_7463);
and U10613 (N_10613,N_7299,N_5267);
and U10614 (N_10614,N_7606,N_9666);
xor U10615 (N_10615,N_9976,N_5322);
xnor U10616 (N_10616,N_9401,N_5209);
or U10617 (N_10617,N_7689,N_9086);
or U10618 (N_10618,N_5890,N_8711);
nor U10619 (N_10619,N_5694,N_8025);
nand U10620 (N_10620,N_9807,N_6407);
or U10621 (N_10621,N_6058,N_5449);
nand U10622 (N_10622,N_9970,N_5413);
xor U10623 (N_10623,N_7225,N_7172);
and U10624 (N_10624,N_5173,N_9511);
and U10625 (N_10625,N_8429,N_6457);
and U10626 (N_10626,N_6076,N_7928);
nand U10627 (N_10627,N_8325,N_6760);
nand U10628 (N_10628,N_8917,N_6809);
xnor U10629 (N_10629,N_6702,N_7196);
nand U10630 (N_10630,N_7721,N_7042);
nand U10631 (N_10631,N_8539,N_5529);
xor U10632 (N_10632,N_6883,N_5179);
or U10633 (N_10633,N_9310,N_7306);
nor U10634 (N_10634,N_8197,N_5191);
or U10635 (N_10635,N_5525,N_8204);
xnor U10636 (N_10636,N_7705,N_8314);
xor U10637 (N_10637,N_6940,N_8712);
xor U10638 (N_10638,N_5240,N_7639);
nand U10639 (N_10639,N_7825,N_8658);
or U10640 (N_10640,N_9172,N_8277);
xor U10641 (N_10641,N_7926,N_7343);
and U10642 (N_10642,N_6444,N_5857);
or U10643 (N_10643,N_8890,N_5027);
nand U10644 (N_10644,N_8142,N_5202);
nand U10645 (N_10645,N_9705,N_5974);
or U10646 (N_10646,N_5653,N_5952);
nor U10647 (N_10647,N_9792,N_6613);
xor U10648 (N_10648,N_9250,N_5798);
or U10649 (N_10649,N_7670,N_9386);
nand U10650 (N_10650,N_9388,N_9457);
or U10651 (N_10651,N_8497,N_6701);
nand U10652 (N_10652,N_7829,N_6970);
nor U10653 (N_10653,N_8862,N_5439);
and U10654 (N_10654,N_9101,N_8300);
or U10655 (N_10655,N_5337,N_8212);
xnor U10656 (N_10656,N_8344,N_7626);
xor U10657 (N_10657,N_9429,N_9715);
nand U10658 (N_10658,N_7909,N_8182);
xnor U10659 (N_10659,N_6056,N_6682);
nand U10660 (N_10660,N_5508,N_9008);
nor U10661 (N_10661,N_7851,N_8987);
and U10662 (N_10662,N_5902,N_5492);
nor U10663 (N_10663,N_6977,N_9908);
and U10664 (N_10664,N_6017,N_8252);
nand U10665 (N_10665,N_7571,N_5271);
xnor U10666 (N_10666,N_7960,N_5885);
and U10667 (N_10667,N_5991,N_5729);
and U10668 (N_10668,N_8259,N_5650);
nand U10669 (N_10669,N_7783,N_6824);
or U10670 (N_10670,N_8929,N_9736);
and U10671 (N_10671,N_8031,N_7681);
nand U10672 (N_10672,N_6200,N_6394);
xnor U10673 (N_10673,N_6065,N_5386);
or U10674 (N_10674,N_7008,N_8944);
and U10675 (N_10675,N_6552,N_5865);
nand U10676 (N_10676,N_7017,N_7448);
nor U10677 (N_10677,N_7380,N_9912);
xnor U10678 (N_10678,N_9849,N_6351);
and U10679 (N_10679,N_7716,N_6920);
xnor U10680 (N_10680,N_6258,N_5611);
nor U10681 (N_10681,N_7374,N_8232);
or U10682 (N_10682,N_6239,N_5779);
or U10683 (N_10683,N_9649,N_8002);
and U10684 (N_10684,N_7593,N_5355);
and U10685 (N_10685,N_7945,N_7894);
and U10686 (N_10686,N_7794,N_6664);
nand U10687 (N_10687,N_5603,N_5417);
or U10688 (N_10688,N_9159,N_6459);
xor U10689 (N_10689,N_8334,N_5371);
and U10690 (N_10690,N_9796,N_6030);
nor U10691 (N_10691,N_6277,N_7210);
and U10692 (N_10692,N_6196,N_5569);
nand U10693 (N_10693,N_7047,N_7065);
xnor U10694 (N_10694,N_5822,N_9096);
xnor U10695 (N_10695,N_7239,N_8022);
nand U10696 (N_10696,N_5072,N_8299);
nand U10697 (N_10697,N_5686,N_7181);
or U10698 (N_10698,N_5339,N_9323);
or U10699 (N_10699,N_6094,N_7539);
and U10700 (N_10700,N_8622,N_5214);
xor U10701 (N_10701,N_6668,N_8694);
nand U10702 (N_10702,N_6335,N_9659);
nor U10703 (N_10703,N_5458,N_5171);
xor U10704 (N_10704,N_8388,N_6316);
xor U10705 (N_10705,N_9559,N_9048);
xnor U10706 (N_10706,N_8514,N_6711);
and U10707 (N_10707,N_8884,N_9170);
nand U10708 (N_10708,N_5238,N_8607);
or U10709 (N_10709,N_7854,N_6276);
and U10710 (N_10710,N_7134,N_7371);
xor U10711 (N_10711,N_8993,N_7139);
xor U10712 (N_10712,N_6877,N_6912);
xor U10713 (N_10713,N_6274,N_8637);
and U10714 (N_10714,N_7145,N_7244);
or U10715 (N_10715,N_5436,N_6242);
nand U10716 (N_10716,N_6703,N_9683);
and U10717 (N_10717,N_7569,N_5943);
xor U10718 (N_10718,N_5850,N_7971);
nor U10719 (N_10719,N_5679,N_9393);
or U10720 (N_10720,N_7414,N_6064);
nor U10721 (N_10721,N_6779,N_6500);
xor U10722 (N_10722,N_8111,N_8592);
nor U10723 (N_10723,N_6479,N_8707);
xor U10724 (N_10724,N_6153,N_8551);
xnor U10725 (N_10725,N_9507,N_7424);
or U10726 (N_10726,N_6275,N_5272);
xor U10727 (N_10727,N_6315,N_6709);
xnor U10728 (N_10728,N_8949,N_8088);
or U10729 (N_10729,N_9719,N_8405);
or U10730 (N_10730,N_8086,N_6069);
xnor U10731 (N_10731,N_5696,N_8811);
or U10732 (N_10732,N_7208,N_6778);
xnor U10733 (N_10733,N_5083,N_6319);
xnor U10734 (N_10734,N_6675,N_6966);
xor U10735 (N_10735,N_6341,N_6898);
nor U10736 (N_10736,N_8387,N_7117);
xor U10737 (N_10737,N_8068,N_6466);
nor U10738 (N_10738,N_8223,N_7522);
xnor U10739 (N_10739,N_5388,N_5928);
and U10740 (N_10740,N_8075,N_8070);
xnor U10741 (N_10741,N_9365,N_8585);
or U10742 (N_10742,N_5691,N_7698);
xor U10743 (N_10743,N_8107,N_7986);
nand U10744 (N_10744,N_9913,N_9624);
xnor U10745 (N_10745,N_5239,N_9746);
xor U10746 (N_10746,N_7919,N_9275);
nand U10747 (N_10747,N_9224,N_6626);
nor U10748 (N_10748,N_8550,N_9915);
or U10749 (N_10749,N_5190,N_8513);
xor U10750 (N_10750,N_8544,N_5051);
or U10751 (N_10751,N_5701,N_7190);
or U10752 (N_10752,N_8305,N_7621);
or U10753 (N_10753,N_8353,N_5872);
nand U10754 (N_10754,N_6630,N_8058);
or U10755 (N_10755,N_8097,N_6272);
and U10756 (N_10756,N_9139,N_5709);
nor U10757 (N_10757,N_9253,N_8072);
and U10758 (N_10758,N_6447,N_5226);
xor U10759 (N_10759,N_5553,N_6821);
xor U10760 (N_10760,N_6955,N_9955);
xnor U10761 (N_10761,N_9809,N_9062);
or U10762 (N_10762,N_6497,N_7687);
xnor U10763 (N_10763,N_5967,N_7129);
and U10764 (N_10764,N_5470,N_6542);
xor U10765 (N_10765,N_6228,N_9235);
and U10766 (N_10766,N_5765,N_5959);
nand U10767 (N_10767,N_5280,N_7072);
nand U10768 (N_10768,N_9896,N_6268);
and U10769 (N_10769,N_5338,N_9584);
or U10770 (N_10770,N_9882,N_5253);
or U10771 (N_10771,N_5914,N_6369);
nor U10772 (N_10772,N_8103,N_7599);
nor U10773 (N_10773,N_9806,N_9581);
or U10774 (N_10774,N_7514,N_7445);
nand U10775 (N_10775,N_5921,N_8156);
nand U10776 (N_10776,N_9023,N_8253);
nor U10777 (N_10777,N_7734,N_9980);
and U10778 (N_10778,N_5622,N_7195);
xor U10779 (N_10779,N_7174,N_6439);
nor U10780 (N_10780,N_8769,N_9895);
or U10781 (N_10781,N_9979,N_8432);
nor U10782 (N_10782,N_5333,N_9117);
and U10783 (N_10783,N_6773,N_9879);
xor U10784 (N_10784,N_6010,N_7645);
xor U10785 (N_10785,N_7116,N_7361);
nand U10786 (N_10786,N_9596,N_9532);
nor U10787 (N_10787,N_5261,N_6984);
nand U10788 (N_10788,N_5602,N_9328);
nor U10789 (N_10789,N_8819,N_9273);
nor U10790 (N_10790,N_6117,N_6737);
and U10791 (N_10791,N_6399,N_6472);
and U10792 (N_10792,N_8964,N_5635);
and U10793 (N_10793,N_9742,N_9881);
nand U10794 (N_10794,N_5507,N_7097);
or U10795 (N_10795,N_6317,N_9468);
xor U10796 (N_10796,N_7130,N_8066);
nor U10797 (N_10797,N_8866,N_8569);
xnor U10798 (N_10798,N_7274,N_5870);
xor U10799 (N_10799,N_5141,N_8403);
nand U10800 (N_10800,N_6410,N_9937);
nand U10801 (N_10801,N_9464,N_9651);
or U10802 (N_10802,N_9486,N_6344);
xnor U10803 (N_10803,N_9439,N_9195);
nor U10804 (N_10804,N_6471,N_9531);
or U10805 (N_10805,N_9813,N_9647);
and U10806 (N_10806,N_6680,N_5368);
and U10807 (N_10807,N_8063,N_6209);
nand U10808 (N_10808,N_9588,N_9983);
xor U10809 (N_10809,N_9266,N_8382);
xnor U10810 (N_10810,N_9772,N_5347);
nand U10811 (N_10811,N_5018,N_9777);
xnor U10812 (N_10812,N_7889,N_7830);
xor U10813 (N_10813,N_5938,N_8727);
nor U10814 (N_10814,N_7855,N_5302);
nand U10815 (N_10815,N_5594,N_7368);
or U10816 (N_10816,N_9089,N_9779);
nand U10817 (N_10817,N_5297,N_6632);
nand U10818 (N_10818,N_6491,N_7304);
and U10819 (N_10819,N_6581,N_9578);
nor U10820 (N_10820,N_5089,N_6314);
nor U10821 (N_10821,N_7796,N_5859);
xnor U10822 (N_10822,N_9337,N_8653);
nand U10823 (N_10823,N_6582,N_5461);
xor U10824 (N_10824,N_6057,N_7271);
nor U10825 (N_10825,N_8563,N_6788);
and U10826 (N_10826,N_8400,N_9168);
nand U10827 (N_10827,N_7863,N_5329);
nand U10828 (N_10828,N_7597,N_7691);
or U10829 (N_10829,N_9368,N_6347);
nand U10830 (N_10830,N_7862,N_8784);
nor U10831 (N_10831,N_9414,N_5768);
and U10832 (N_10832,N_8783,N_8840);
or U10833 (N_10833,N_9722,N_8242);
xor U10834 (N_10834,N_6532,N_5501);
nor U10835 (N_10835,N_6577,N_5810);
or U10836 (N_10836,N_9436,N_8122);
nand U10837 (N_10837,N_5121,N_9911);
and U10838 (N_10838,N_9945,N_9702);
or U10839 (N_10839,N_9467,N_7761);
or U10840 (N_10840,N_7405,N_8033);
xnor U10841 (N_10841,N_6384,N_7703);
nand U10842 (N_10842,N_7491,N_7090);
or U10843 (N_10843,N_6206,N_5117);
nor U10844 (N_10844,N_6202,N_6927);
nor U10845 (N_10845,N_8818,N_6131);
nand U10846 (N_10846,N_8480,N_9463);
or U10847 (N_10847,N_6956,N_7202);
xnor U10848 (N_10848,N_5161,N_5396);
nand U10849 (N_10849,N_7878,N_6482);
xnor U10850 (N_10850,N_7218,N_9967);
xnor U10851 (N_10851,N_6768,N_9270);
or U10852 (N_10852,N_8900,N_7435);
xnor U10853 (N_10853,N_7931,N_8081);
nand U10854 (N_10854,N_6913,N_7148);
nand U10855 (N_10855,N_8796,N_5043);
nand U10856 (N_10856,N_7149,N_5757);
xnor U10857 (N_10857,N_6166,N_5549);
nor U10858 (N_10858,N_7908,N_9306);
and U10859 (N_10859,N_5824,N_8100);
xnor U10860 (N_10860,N_8872,N_8794);
xor U10861 (N_10861,N_7009,N_6027);
or U10862 (N_10862,N_8675,N_6568);
and U10863 (N_10863,N_9927,N_5896);
nor U10864 (N_10864,N_6343,N_8027);
nand U10865 (N_10865,N_8699,N_5012);
or U10866 (N_10866,N_9412,N_6887);
xor U10867 (N_10867,N_5377,N_8739);
nand U10868 (N_10868,N_6943,N_7466);
and U10869 (N_10869,N_6433,N_6207);
xor U10870 (N_10870,N_8178,N_6654);
or U10871 (N_10871,N_6586,N_8507);
nor U10872 (N_10872,N_5264,N_8889);
xnor U10873 (N_10873,N_7162,N_8040);
or U10874 (N_10874,N_9602,N_9352);
xnor U10875 (N_10875,N_8205,N_9459);
nand U10876 (N_10876,N_8588,N_5379);
nor U10877 (N_10877,N_7041,N_7678);
nand U10878 (N_10878,N_6124,N_7674);
nand U10879 (N_10879,N_5223,N_5415);
or U10880 (N_10880,N_7654,N_9787);
nor U10881 (N_10881,N_6002,N_5150);
nand U10882 (N_10882,N_9926,N_5224);
or U10883 (N_10883,N_5858,N_7280);
and U10884 (N_10884,N_9179,N_8927);
or U10885 (N_10885,N_5801,N_6957);
and U10886 (N_10886,N_5956,N_7874);
xnor U10887 (N_10887,N_9411,N_6557);
nand U10888 (N_10888,N_9029,N_5783);
or U10889 (N_10889,N_8102,N_7092);
xnor U10890 (N_10890,N_7443,N_9918);
or U10891 (N_10891,N_8234,N_8376);
nand U10892 (N_10892,N_7025,N_9648);
nand U10893 (N_10893,N_5314,N_9285);
nand U10894 (N_10894,N_9432,N_8343);
xor U10895 (N_10895,N_6290,N_5781);
nor U10896 (N_10896,N_9450,N_7506);
xor U10897 (N_10897,N_7340,N_5394);
nor U10898 (N_10898,N_6653,N_5423);
nand U10899 (N_10899,N_8576,N_6361);
and U10900 (N_10900,N_5404,N_7364);
nand U10901 (N_10901,N_9141,N_5862);
nor U10902 (N_10902,N_9026,N_7482);
or U10903 (N_10903,N_5957,N_7557);
nor U10904 (N_10904,N_9923,N_6034);
xor U10905 (N_10905,N_9111,N_7987);
xnor U10906 (N_10906,N_5029,N_9884);
xor U10907 (N_10907,N_6981,N_5445);
and U10908 (N_10908,N_5596,N_7604);
nand U10909 (N_10909,N_6061,N_8985);
nand U10910 (N_10910,N_8830,N_6805);
or U10911 (N_10911,N_8860,N_8562);
nand U10912 (N_10912,N_5973,N_6462);
xor U10913 (N_10913,N_6285,N_8808);
xor U10914 (N_10914,N_6214,N_7069);
nor U10915 (N_10915,N_9031,N_6505);
nand U10916 (N_10916,N_5085,N_7211);
or U10917 (N_10917,N_8898,N_6492);
nor U10918 (N_10918,N_9476,N_8913);
nor U10919 (N_10919,N_8437,N_7676);
xor U10920 (N_10920,N_6311,N_6721);
or U10921 (N_10921,N_7185,N_9774);
nand U10922 (N_10922,N_7039,N_9866);
nor U10923 (N_10923,N_5831,N_9589);
nor U10924 (N_10924,N_6974,N_8304);
xnor U10925 (N_10925,N_6128,N_9601);
or U10926 (N_10926,N_9116,N_7001);
and U10927 (N_10927,N_5213,N_9472);
and U10928 (N_10928,N_7941,N_7245);
nor U10929 (N_10929,N_7643,N_7966);
nand U10930 (N_10930,N_7220,N_5651);
and U10931 (N_10931,N_5047,N_6674);
xor U10932 (N_10932,N_5740,N_7948);
or U10933 (N_10933,N_6408,N_5868);
nand U10934 (N_10934,N_8517,N_7309);
and U10935 (N_10935,N_7329,N_9660);
and U10936 (N_10936,N_6104,N_5154);
xnor U10937 (N_10937,N_6736,N_9633);
and U10938 (N_10938,N_7859,N_7446);
and U10939 (N_10939,N_9519,N_6739);
nand U10940 (N_10940,N_6941,N_6264);
and U10941 (N_10941,N_9105,N_7260);
nor U10942 (N_10942,N_8648,N_9246);
nand U10943 (N_10943,N_8408,N_7974);
xnor U10944 (N_10944,N_9540,N_9264);
and U10945 (N_10945,N_6575,N_5234);
and U10946 (N_10946,N_9359,N_6159);
xor U10947 (N_10947,N_5325,N_9248);
or U10948 (N_10948,N_5496,N_6245);
xor U10949 (N_10949,N_5512,N_5590);
and U10950 (N_10950,N_7718,N_8580);
and U10951 (N_10951,N_7024,N_7246);
and U10952 (N_10952,N_6580,N_6661);
xor U10953 (N_10953,N_5091,N_8239);
nand U10954 (N_10954,N_6508,N_8189);
nor U10955 (N_10955,N_7560,N_8328);
or U10956 (N_10956,N_7372,N_7417);
or U10957 (N_10957,N_7470,N_7644);
or U10958 (N_10958,N_5211,N_6318);
nand U10959 (N_10959,N_5448,N_5233);
and U10960 (N_10960,N_6951,N_9832);
xor U10961 (N_10961,N_7565,N_5960);
xnor U10962 (N_10962,N_5220,N_9767);
xor U10963 (N_10963,N_7062,N_9989);
nand U10964 (N_10964,N_5033,N_6555);
nor U10965 (N_10965,N_9586,N_5613);
nand U10966 (N_10966,N_7176,N_6789);
nor U10967 (N_10967,N_8512,N_9197);
nor U10968 (N_10968,N_6987,N_5021);
nor U10969 (N_10969,N_8603,N_7628);
or U10970 (N_10970,N_7769,N_9582);
and U10971 (N_10971,N_5523,N_7672);
nor U10972 (N_10972,N_7588,N_5848);
or U10973 (N_10973,N_7438,N_6446);
nand U10974 (N_10974,N_6544,N_6511);
and U10975 (N_10975,N_9843,N_8258);
and U10976 (N_10976,N_5153,N_8032);
xor U10977 (N_10977,N_8935,N_5699);
xnor U10978 (N_10978,N_6310,N_7711);
nor U10979 (N_10979,N_9696,N_9192);
nor U10980 (N_10980,N_8652,N_8004);
nand U10981 (N_10981,N_9672,N_6255);
nor U10982 (N_10982,N_7525,N_8123);
nand U10983 (N_10983,N_6929,N_9959);
nand U10984 (N_10984,N_7541,N_8997);
xnor U10985 (N_10985,N_6456,N_6125);
nand U10986 (N_10986,N_6312,N_5055);
and U10987 (N_10987,N_8373,N_5873);
and U10988 (N_10988,N_6717,N_7086);
or U10989 (N_10989,N_5736,N_9652);
xnor U10990 (N_10990,N_8612,N_5344);
and U10991 (N_10991,N_8255,N_5861);
nand U10992 (N_10992,N_6453,N_8735);
and U10993 (N_10993,N_7616,N_8019);
nor U10994 (N_10994,N_8369,N_8602);
nand U10995 (N_10995,N_7930,N_6604);
and U10996 (N_10996,N_9888,N_9383);
or U10997 (N_10997,N_9173,N_8876);
nand U10998 (N_10998,N_6969,N_8595);
nor U10999 (N_10999,N_5715,N_9322);
nand U11000 (N_11000,N_7513,N_7192);
xor U11001 (N_11001,N_9972,N_6234);
xor U11002 (N_11002,N_8516,N_8155);
or U11003 (N_11003,N_9871,N_6714);
nand U11004 (N_11004,N_5869,N_5071);
and U11005 (N_11005,N_9938,N_6237);
nand U11006 (N_11006,N_8561,N_8430);
nand U11007 (N_11007,N_6878,N_6292);
nand U11008 (N_11008,N_5317,N_5406);
nor U11009 (N_11009,N_7551,N_8140);
nand U11010 (N_11010,N_9289,N_8922);
and U11011 (N_11011,N_7704,N_5746);
xnor U11012 (N_11012,N_6143,N_5399);
and U11013 (N_11013,N_9946,N_5376);
nand U11014 (N_11014,N_7970,N_5505);
xor U11015 (N_11015,N_9845,N_8756);
and U11016 (N_11016,N_6464,N_9680);
nor U11017 (N_11017,N_8173,N_7903);
and U11018 (N_11018,N_7213,N_6583);
and U11019 (N_11019,N_6259,N_8348);
nor U11020 (N_11020,N_6774,N_6417);
nor U11021 (N_11021,N_8654,N_6420);
nand U11022 (N_11022,N_9634,N_9526);
nand U11023 (N_11023,N_8671,N_9135);
nor U11024 (N_11024,N_8868,N_5362);
nor U11025 (N_11025,N_9422,N_9283);
and U11026 (N_11026,N_9785,N_7440);
xor U11027 (N_11027,N_6093,N_9673);
and U11028 (N_11028,N_5937,N_7269);
or U11029 (N_11029,N_7276,N_5663);
xor U11030 (N_11030,N_8833,N_8582);
xnor U11031 (N_11031,N_7315,N_6766);
and U11032 (N_11032,N_7620,N_9206);
nor U11033 (N_11033,N_8026,N_7150);
xor U11034 (N_11034,N_6911,N_5479);
and U11035 (N_11035,N_8813,N_9565);
nand U11036 (N_11036,N_8729,N_6070);
or U11037 (N_11037,N_8535,N_6236);
and U11038 (N_11038,N_9714,N_8389);
nand U11039 (N_11039,N_9692,N_8275);
or U11040 (N_11040,N_5809,N_8802);
and U11041 (N_11041,N_9407,N_9662);
xor U11042 (N_11042,N_6603,N_5228);
and U11043 (N_11043,N_5431,N_9287);
and U11044 (N_11044,N_9538,N_9397);
nor U11045 (N_11045,N_6595,N_6204);
nand U11046 (N_11046,N_7509,N_9093);
nor U11047 (N_11047,N_8433,N_6876);
nor U11048 (N_11048,N_5474,N_9166);
nand U11049 (N_11049,N_6922,N_7667);
xnor U11050 (N_11050,N_9403,N_7083);
nor U11051 (N_11051,N_8352,N_5380);
nor U11052 (N_11052,N_9343,N_7848);
or U11053 (N_11053,N_7770,N_5129);
and U11054 (N_11054,N_8882,N_5919);
or U11055 (N_11055,N_9090,N_5354);
xnor U11056 (N_11056,N_5046,N_5964);
and U11057 (N_11057,N_9988,N_7126);
nand U11058 (N_11058,N_7520,N_9091);
xnor U11059 (N_11059,N_6468,N_7996);
and U11060 (N_11060,N_9267,N_8203);
xor U11061 (N_11061,N_8279,N_5589);
xnor U11062 (N_11062,N_7963,N_8467);
or U11063 (N_11063,N_5499,N_6726);
nor U11064 (N_11064,N_9193,N_7764);
and U11065 (N_11065,N_7856,N_6868);
nor U11066 (N_11066,N_6933,N_9148);
or U11067 (N_11067,N_5188,N_7911);
or U11068 (N_11068,N_6012,N_6313);
nor U11069 (N_11069,N_5382,N_6147);
or U11070 (N_11070,N_5958,N_9575);
xor U11071 (N_11071,N_9220,N_9998);
nor U11072 (N_11072,N_7322,N_8524);
nand U11073 (N_11073,N_6406,N_8361);
and U11074 (N_11074,N_6837,N_7049);
nand U11075 (N_11075,N_8947,N_5996);
nand U11076 (N_11076,N_9300,N_7472);
or U11077 (N_11077,N_8251,N_9064);
and U11078 (N_11078,N_9577,N_8116);
nor U11079 (N_11079,N_5303,N_5494);
or U11080 (N_11080,N_5044,N_7858);
or U11081 (N_11081,N_6465,N_7924);
xnor U11082 (N_11082,N_8235,N_5210);
and U11083 (N_11083,N_9217,N_6804);
and U11084 (N_11084,N_7580,N_9303);
nor U11085 (N_11085,N_5630,N_7232);
or U11086 (N_11086,N_9071,N_5014);
xor U11087 (N_11087,N_5370,N_7460);
or U11088 (N_11088,N_5315,N_7054);
nand U11089 (N_11089,N_7301,N_5102);
and U11090 (N_11090,N_9857,N_8254);
nor U11091 (N_11091,N_7223,N_5762);
or U11092 (N_11092,N_8034,N_9376);
nand U11093 (N_11093,N_6232,N_8496);
nor U11094 (N_11094,N_6695,N_5269);
nand U11095 (N_11095,N_5434,N_6836);
nor U11096 (N_11096,N_8478,N_8067);
or U11097 (N_11097,N_8319,N_9473);
nand U11098 (N_11098,N_7132,N_7461);
nor U11099 (N_11099,N_7992,N_9769);
nor U11100 (N_11100,N_6363,N_9688);
nand U11101 (N_11101,N_6066,N_5288);
xor U11102 (N_11102,N_6325,N_6427);
xnor U11103 (N_11103,N_9374,N_5876);
or U11104 (N_11104,N_7543,N_7108);
nand U11105 (N_11105,N_9668,N_9277);
nand U11106 (N_11106,N_8779,N_6923);
nor U11107 (N_11107,N_8895,N_9153);
or U11108 (N_11108,N_5205,N_9241);
xor U11109 (N_11109,N_9445,N_9670);
nor U11110 (N_11110,N_5484,N_5090);
nand U11111 (N_11111,N_6480,N_8896);
nand U11112 (N_11112,N_6991,N_7842);
and U11113 (N_11113,N_6418,N_9102);
or U11114 (N_11114,N_6477,N_5980);
nand U11115 (N_11115,N_7142,N_8492);
and U11116 (N_11116,N_8237,N_5880);
xnor U11117 (N_11117,N_7403,N_9261);
xor U11118 (N_11118,N_6801,N_5446);
or U11119 (N_11119,N_7802,N_8594);
or U11120 (N_11120,N_8457,N_6072);
and U11121 (N_11121,N_9426,N_9942);
and U11122 (N_11122,N_5260,N_6324);
xnor U11123 (N_11123,N_6919,N_9952);
nand U11124 (N_11124,N_9847,N_5113);
xnor U11125 (N_11125,N_5811,N_7564);
xnor U11126 (N_11126,N_5939,N_5477);
xor U11127 (N_11127,N_9305,N_9078);
or U11128 (N_11128,N_9315,N_8346);
nand U11129 (N_11129,N_7529,N_8915);
nand U11130 (N_11130,N_9149,N_9380);
and U11131 (N_11131,N_6016,N_5255);
and U11132 (N_11132,N_8817,N_7338);
xor U11133 (N_11133,N_8153,N_5070);
or U11134 (N_11134,N_9515,N_5024);
nor U11135 (N_11135,N_9413,N_9735);
nand U11136 (N_11136,N_6565,N_6719);
and U11137 (N_11137,N_6345,N_6959);
nor U11138 (N_11138,N_8630,N_5308);
xnor U11139 (N_11139,N_7507,N_9829);
xnor U11140 (N_11140,N_7631,N_7861);
or U11141 (N_11141,N_9522,N_5881);
or U11142 (N_11142,N_7087,N_5257);
xnor U11143 (N_11143,N_5095,N_7756);
xor U11144 (N_11144,N_7496,N_9636);
and U11145 (N_11145,N_9213,N_6336);
xnor U11146 (N_11146,N_9934,N_7321);
and U11147 (N_11147,N_8415,N_5830);
xnor U11148 (N_11148,N_9114,N_8484);
nor U11149 (N_11149,N_5720,N_7318);
xnor U11150 (N_11150,N_8596,N_8564);
and U11151 (N_11151,N_5587,N_9314);
and U11152 (N_11152,N_8445,N_8054);
nor U11153 (N_11153,N_5231,N_6591);
or U11154 (N_11154,N_9569,N_9867);
xor U11155 (N_11155,N_9040,N_9151);
nand U11156 (N_11156,N_5456,N_5737);
nand U11157 (N_11157,N_5752,N_6328);
nand U11158 (N_11158,N_9941,N_8547);
nor U11159 (N_11159,N_6740,N_9508);
or U11160 (N_11160,N_9345,N_6606);
nand U11161 (N_11161,N_5647,N_8549);
or U11162 (N_11162,N_9517,N_7167);
xor U11163 (N_11163,N_6600,N_7159);
or U11164 (N_11164,N_6496,N_9990);
and U11165 (N_11165,N_8109,N_6271);
nand U11166 (N_11166,N_5621,N_9831);
or U11167 (N_11167,N_7865,N_5771);
xor U11168 (N_11168,N_9650,N_5389);
or U11169 (N_11169,N_6233,N_9697);
nand U11170 (N_11170,N_7767,N_9982);
xor U11171 (N_11171,N_6905,N_5026);
or U11172 (N_11172,N_6270,N_6389);
xnor U11173 (N_11173,N_8765,N_8984);
or U11174 (N_11174,N_5662,N_5131);
nor U11175 (N_11175,N_7697,N_5088);
xnor U11176 (N_11176,N_7423,N_6463);
or U11177 (N_11177,N_8555,N_7291);
and U11178 (N_11178,N_9471,N_7359);
xnor U11179 (N_11179,N_8781,N_7477);
nor U11180 (N_11180,N_9018,N_6949);
or U11181 (N_11181,N_7197,N_7812);
or U11182 (N_11182,N_5067,N_7004);
and U11183 (N_11183,N_9768,N_6759);
nor U11184 (N_11184,N_6007,N_7093);
xnor U11185 (N_11185,N_8196,N_7253);
and U11186 (N_11186,N_8364,N_6095);
xor U11187 (N_11187,N_5435,N_5422);
and U11188 (N_11188,N_5997,N_7454);
nand U11189 (N_11189,N_7642,N_7459);
nand U11190 (N_11190,N_6379,N_6135);
nand U11191 (N_11191,N_8447,N_5506);
or U11192 (N_11192,N_8175,N_7745);
nand U11193 (N_11193,N_6822,N_8342);
or U11194 (N_11194,N_5713,N_5946);
xnor U11195 (N_11195,N_6924,N_7155);
or U11196 (N_11196,N_6450,N_6385);
nand U11197 (N_11197,N_5778,N_8365);
xnor U11198 (N_11198,N_5169,N_5166);
or U11199 (N_11199,N_5471,N_9419);
or U11200 (N_11200,N_8035,N_5035);
and U11201 (N_11201,N_9695,N_8108);
or U11202 (N_11202,N_7073,N_5128);
and U11203 (N_11203,N_9317,N_6451);
or U11204 (N_11204,N_5151,N_8939);
or U11205 (N_11205,N_7360,N_5717);
or U11206 (N_11206,N_6097,N_6642);
xnor U11207 (N_11207,N_8303,N_8451);
and U11208 (N_11208,N_5556,N_8308);
nor U11209 (N_11209,N_9977,N_6763);
or U11210 (N_11210,N_9618,N_9311);
and U11211 (N_11211,N_6527,N_9510);
nand U11212 (N_11212,N_7655,N_7296);
nand U11213 (N_11213,N_5398,N_9808);
or U11214 (N_11214,N_8810,N_5764);
or U11215 (N_11215,N_7358,N_7021);
nor U11216 (N_11216,N_7640,N_7398);
nor U11217 (N_11217,N_6570,N_8481);
and U11218 (N_11218,N_8198,N_7337);
nor U11219 (N_11219,N_5476,N_6965);
nand U11220 (N_11220,N_5125,N_6842);
xnor U11221 (N_11221,N_6529,N_9284);
nand U11222 (N_11222,N_6261,N_9389);
nand U11223 (N_11223,N_5493,N_9765);
nand U11224 (N_11224,N_5769,N_6862);
and U11225 (N_11225,N_9870,N_5640);
nand U11226 (N_11226,N_9125,N_8135);
and U11227 (N_11227,N_9435,N_6525);
nor U11228 (N_11228,N_5844,N_9711);
and U11229 (N_11229,N_8288,N_7389);
or U11230 (N_11230,N_9004,N_5853);
nand U11231 (N_11231,N_5048,N_6019);
or U11232 (N_11232,N_7415,N_9859);
nand U11233 (N_11233,N_7379,N_8483);
xor U11234 (N_11234,N_6867,N_7553);
nand U11235 (N_11235,N_7969,N_7064);
xnor U11236 (N_11236,N_5905,N_6571);
and U11237 (N_11237,N_6182,N_5081);
or U11238 (N_11238,N_9663,N_6854);
and U11239 (N_11239,N_5372,N_7044);
nand U11240 (N_11240,N_5252,N_6164);
nand U11241 (N_11241,N_6963,N_6013);
and U11242 (N_11242,N_9032,N_6470);
or U11243 (N_11243,N_5393,N_5221);
nor U11244 (N_11244,N_9158,N_6126);
nand U11245 (N_11245,N_6495,N_5767);
and U11246 (N_11246,N_8545,N_5054);
and U11247 (N_11247,N_8608,N_5312);
nand U11248 (N_11248,N_8431,N_5978);
or U11249 (N_11249,N_7289,N_6080);
or U11250 (N_11250,N_6884,N_5697);
and U11251 (N_11251,N_8211,N_6899);
nor U11252 (N_11252,N_5826,N_8003);
or U11253 (N_11253,N_5949,N_5787);
nor U11254 (N_11254,N_5897,N_5567);
and U11255 (N_11255,N_7077,N_6499);
xor U11256 (N_11256,N_5485,N_9321);
or U11257 (N_11257,N_7731,N_9104);
nor U11258 (N_11258,N_6551,N_6267);
or U11259 (N_11259,N_6942,N_6132);
or U11260 (N_11260,N_7779,N_8946);
nor U11261 (N_11261,N_7661,N_9921);
nor U11262 (N_11262,N_5304,N_9620);
nor U11263 (N_11263,N_6937,N_9891);
nand U11264 (N_11264,N_5073,N_7602);
nor U11265 (N_11265,N_5454,N_7927);
and U11266 (N_11266,N_9687,N_7153);
nand U11267 (N_11267,N_6813,N_8024);
or U11268 (N_11268,N_8397,N_6308);
and U11269 (N_11269,N_6148,N_9800);
or U11270 (N_11270,N_9443,N_5360);
and U11271 (N_11271,N_7594,N_5989);
or U11272 (N_11272,N_9007,N_9330);
nor U11273 (N_11273,N_7277,N_6932);
xor U11274 (N_11274,N_6639,N_7141);
nor U11275 (N_11275,N_5412,N_5619);
nand U11276 (N_11276,N_9299,N_5421);
nand U11277 (N_11277,N_8297,N_5760);
nand U11278 (N_11278,N_7279,N_6426);
or U11279 (N_11279,N_8726,N_6936);
and U11280 (N_11280,N_8933,N_8176);
and U11281 (N_11281,N_6286,N_8409);
or U11282 (N_11282,N_5538,N_6914);
and U11283 (N_11283,N_5658,N_7742);
and U11284 (N_11284,N_7241,N_7968);
nor U11285 (N_11285,N_5059,N_8780);
xor U11286 (N_11286,N_7614,N_5560);
xor U11287 (N_11287,N_9603,N_8634);
nor U11288 (N_11288,N_9136,N_7946);
and U11289 (N_11289,N_9901,N_9855);
nand U11290 (N_11290,N_7568,N_7206);
and U11291 (N_11291,N_5533,N_7534);
or U11292 (N_11292,N_5263,N_5564);
or U11293 (N_11293,N_9598,N_5313);
xnor U11294 (N_11294,N_9788,N_7237);
xnor U11295 (N_11295,N_6618,N_9385);
and U11296 (N_11296,N_7081,N_7410);
nand U11297 (N_11297,N_8970,N_5111);
nand U11298 (N_11298,N_5409,N_7091);
xnor U11299 (N_11299,N_9954,N_9707);
nor U11300 (N_11300,N_8960,N_6145);
or U11301 (N_11301,N_9904,N_9373);
and U11302 (N_11302,N_7485,N_7898);
xor U11303 (N_11303,N_9208,N_9933);
and U11304 (N_11304,N_8509,N_5146);
or U11305 (N_11305,N_5490,N_7595);
xnor U11306 (N_11306,N_9059,N_9049);
nor U11307 (N_11307,N_8166,N_5427);
nor U11308 (N_11308,N_8573,N_8990);
or U11309 (N_11309,N_6666,N_9764);
xnor U11310 (N_11310,N_7060,N_8978);
nand U11311 (N_11311,N_5929,N_6000);
and U11312 (N_11312,N_5318,N_7416);
or U11313 (N_11313,N_7106,N_8499);
nor U11314 (N_11314,N_9643,N_9244);
nor U11315 (N_11315,N_6288,N_8301);
or U11316 (N_11316,N_8801,N_8565);
nor U11317 (N_11317,N_6693,N_9748);
and U11318 (N_11318,N_7999,N_9862);
nand U11319 (N_11319,N_9341,N_5660);
nand U11320 (N_11320,N_8394,N_8805);
and U11321 (N_11321,N_6562,N_5582);
nand U11322 (N_11322,N_9425,N_7068);
or U11323 (N_11323,N_6607,N_9720);
nand U11324 (N_11324,N_6247,N_7959);
xor U11325 (N_11325,N_6885,N_5591);
xor U11326 (N_11326,N_9070,N_5585);
and U11327 (N_11327,N_9434,N_7950);
nand U11328 (N_11328,N_9312,N_6376);
nand U11329 (N_11329,N_7582,N_7662);
or U11330 (N_11330,N_8466,N_8493);
or U11331 (N_11331,N_7719,N_6089);
or U11332 (N_11332,N_7447,N_7353);
nor U11333 (N_11333,N_6841,N_6844);
nand U11334 (N_11334,N_6953,N_8422);
and U11335 (N_11335,N_6694,N_6295);
nand U11336 (N_11336,N_8708,N_6814);
or U11337 (N_11337,N_8307,N_8502);
or U11338 (N_11338,N_5692,N_5418);
or U11339 (N_11339,N_5106,N_8278);
nand U11340 (N_11340,N_6785,N_8533);
nand U11341 (N_11341,N_9899,N_7554);
or U11342 (N_11342,N_6890,N_5180);
xor U11343 (N_11343,N_6861,N_8177);
nor U11344 (N_11344,N_7015,N_5149);
nand U11345 (N_11345,N_8246,N_5813);
nor U11346 (N_11346,N_7345,N_7492);
and U11347 (N_11347,N_5539,N_5794);
or U11348 (N_11348,N_6205,N_5077);
or U11349 (N_11349,N_9366,N_8062);
and U11350 (N_11350,N_7572,N_9335);
xnor U11351 (N_11351,N_8472,N_7137);
nand U11352 (N_11352,N_7465,N_9415);
and U11353 (N_11353,N_7037,N_7880);
nor U11354 (N_11354,N_5428,N_8014);
nand U11355 (N_11355,N_7896,N_8723);
xnor U11356 (N_11356,N_8290,N_9025);
and U11357 (N_11357,N_7228,N_7601);
and U11358 (N_11358,N_7897,N_8283);
or U11359 (N_11359,N_9147,N_8138);
and U11360 (N_11360,N_5498,N_8519);
nor U11361 (N_11361,N_5475,N_9200);
nand U11362 (N_11362,N_9088,N_9446);
nand U11363 (N_11363,N_8276,N_5773);
or U11364 (N_11364,N_5631,N_6339);
nand U11365 (N_11365,N_8391,N_9553);
nor U11366 (N_11366,N_7881,N_7292);
and U11367 (N_11367,N_9044,N_9747);
and U11368 (N_11368,N_5277,N_7985);
or U11369 (N_11369,N_9319,N_8679);
xor U11370 (N_11370,N_6733,N_5610);
nor U11371 (N_11371,N_6706,N_5528);
and U11372 (N_11372,N_8669,N_6816);
xor U11373 (N_11373,N_7922,N_7576);
nor U11374 (N_11374,N_6045,N_8677);
xor U11375 (N_11375,N_7273,N_7303);
and U11376 (N_11376,N_5164,N_5931);
and U11377 (N_11377,N_6346,N_7109);
nor U11378 (N_11378,N_7544,N_6352);
or U11379 (N_11379,N_6894,N_9611);
nand U11380 (N_11380,N_8761,N_7408);
or U11381 (N_11381,N_9492,N_9329);
nor U11382 (N_11382,N_7559,N_6423);
and U11383 (N_11383,N_8087,N_5459);
or U11384 (N_11384,N_9505,N_8804);
nand U11385 (N_11385,N_6038,N_5645);
nand U11386 (N_11386,N_5927,N_5309);
nor U11387 (N_11387,N_5530,N_6723);
nor U11388 (N_11388,N_5219,N_8398);
or U11389 (N_11389,N_8626,N_8270);
xnor U11390 (N_11390,N_7314,N_6753);
nor U11391 (N_11391,N_7838,N_6368);
xor U11392 (N_11392,N_6486,N_8336);
xnor U11393 (N_11393,N_8413,N_7388);
nand U11394 (N_11394,N_7409,N_8721);
xnor U11395 (N_11395,N_8775,N_8280);
and U11396 (N_11396,N_9308,N_6996);
xnor U11397 (N_11397,N_7362,N_7107);
nor U11398 (N_11398,N_9828,N_9163);
xnor U11399 (N_11399,N_6950,N_8991);
nand U11400 (N_11400,N_6915,N_9399);
or U11401 (N_11401,N_7738,N_9001);
nand U11402 (N_11402,N_8617,N_7402);
nand U11403 (N_11403,N_5728,N_9791);
or U11404 (N_11404,N_5447,N_8583);
xnor U11405 (N_11405,N_5738,N_5899);
nor U11406 (N_11406,N_7867,N_6248);
and U11407 (N_11407,N_6728,N_6067);
or U11408 (N_11408,N_5573,N_7776);
or U11409 (N_11409,N_7973,N_5045);
nand U11410 (N_11410,N_6515,N_9363);
nor U11411 (N_11411,N_6366,N_5583);
xor U11412 (N_11412,N_6460,N_8221);
nor U11413 (N_11413,N_6850,N_5265);
or U11414 (N_11414,N_7078,N_8085);
and U11415 (N_11415,N_9251,N_6475);
and U11416 (N_11416,N_7549,N_7567);
nor U11417 (N_11417,N_9566,N_9725);
and U11418 (N_11418,N_6374,N_5275);
or U11419 (N_11419,N_8473,N_5068);
and U11420 (N_11420,N_9221,N_9818);
nand U11421 (N_11421,N_5204,N_7775);
or U11422 (N_11422,N_7803,N_6435);
and U11423 (N_11423,N_7266,N_9950);
xnor U11424 (N_11424,N_6712,N_8250);
nand U11425 (N_11425,N_6547,N_7762);
xnor U11426 (N_11426,N_8716,N_8753);
nor U11427 (N_11427,N_6168,N_5950);
xor U11428 (N_11428,N_9036,N_5216);
xor U11429 (N_11429,N_9024,N_8458);
xnor U11430 (N_11430,N_8210,N_9749);
or U11431 (N_11431,N_6767,N_5385);
xor U11432 (N_11432,N_9369,N_5455);
xor U11433 (N_11433,N_5433,N_7957);
xor U11434 (N_11434,N_8725,N_7070);
xnor U11435 (N_11435,N_5903,N_7489);
nor U11436 (N_11436,N_7955,N_9844);
and U11437 (N_11437,N_6167,N_7590);
and U11438 (N_11438,N_6783,N_8486);
xor U11439 (N_11439,N_5273,N_6692);
nor U11440 (N_11440,N_8508,N_8870);
nor U11441 (N_11441,N_9358,N_9645);
and U11442 (N_11442,N_7833,N_5671);
xnor U11443 (N_11443,N_9778,N_9156);
or U11444 (N_11444,N_9298,N_9440);
and U11445 (N_11445,N_9424,N_9524);
xnor U11446 (N_11446,N_8488,N_6035);
or U11447 (N_11447,N_5469,N_7166);
and U11448 (N_11448,N_9292,N_7664);
nor U11449 (N_11449,N_5725,N_6895);
or U11450 (N_11450,N_8972,N_9293);
and U11451 (N_11451,N_7357,N_5923);
xor U11452 (N_11452,N_7323,N_8885);
and U11453 (N_11453,N_5159,N_6825);
xnor U11454 (N_11454,N_5641,N_5754);
nor U11455 (N_11455,N_8423,N_7203);
or U11456 (N_11456,N_8296,N_9199);
nor U11457 (N_11457,N_5497,N_7624);
nand U11458 (N_11458,N_8202,N_9087);
and U11459 (N_11459,N_7892,N_9852);
nor U11460 (N_11460,N_8695,N_7227);
and U11461 (N_11461,N_5351,N_8642);
and U11462 (N_11462,N_7665,N_9006);
or U11463 (N_11463,N_8534,N_6146);
and U11464 (N_11464,N_5693,N_6323);
and U11465 (N_11465,N_6225,N_6218);
or U11466 (N_11466,N_6353,N_7630);
and U11467 (N_11467,N_8910,N_5675);
or U11468 (N_11468,N_8570,N_6078);
or U11469 (N_11469,N_8455,N_7251);
nor U11470 (N_11470,N_8552,N_5242);
and U11471 (N_11471,N_7766,N_6597);
nor U11472 (N_11472,N_7444,N_9075);
nand U11473 (N_11473,N_9745,N_7029);
nor U11474 (N_11474,N_7937,N_7555);
nand U11475 (N_11475,N_6573,N_7993);
and U11476 (N_11476,N_5168,N_5331);
nand U11477 (N_11477,N_7349,N_8245);
xor U11478 (N_11478,N_6015,N_7832);
nor U11479 (N_11479,N_5425,N_9155);
and U11480 (N_11480,N_5796,N_9127);
xnor U11481 (N_11481,N_7521,N_9361);
xor U11482 (N_11482,N_9065,N_5620);
or U11483 (N_11483,N_8090,N_7753);
or U11484 (N_11484,N_8453,N_9165);
nor U11485 (N_11485,N_8741,N_7493);
xor U11486 (N_11486,N_7133,N_9350);
nand U11487 (N_11487,N_5008,N_8831);
or U11488 (N_11488,N_9092,N_8479);
nor U11489 (N_11489,N_8999,N_5212);
xnor U11490 (N_11490,N_8605,N_5828);
and U11491 (N_11491,N_6109,N_7131);
or U11492 (N_11492,N_7324,N_6934);
nand U11493 (N_11493,N_7740,N_8018);
or U11494 (N_11494,N_8720,N_9641);
or U11495 (N_11495,N_5678,N_5369);
nor U11496 (N_11496,N_7103,N_6567);
nor U11497 (N_11497,N_8050,N_8504);
xnor U11498 (N_11498,N_6031,N_9375);
xnor U11499 (N_11499,N_6979,N_8159);
nor U11500 (N_11500,N_7169,N_6037);
nand U11501 (N_11501,N_9097,N_7600);
xnor U11502 (N_11502,N_5259,N_8030);
nor U11503 (N_11503,N_7519,N_6644);
nor U11504 (N_11504,N_9138,N_5543);
nand U11505 (N_11505,N_8037,N_5879);
nor U11506 (N_11506,N_9654,N_9790);
nor U11507 (N_11507,N_7659,N_5514);
nor U11508 (N_11508,N_6130,N_6381);
nand U11509 (N_11509,N_9420,N_9257);
or U11510 (N_11510,N_7427,N_7989);
xnor U11511 (N_11511,N_7849,N_8281);
xor U11512 (N_11512,N_6134,N_7191);
nand U11513 (N_11513,N_6074,N_5891);
nand U11514 (N_11514,N_9130,N_6302);
and U11515 (N_11515,N_9106,N_6024);
xor U11516 (N_11516,N_6047,N_5559);
and U11517 (N_11517,N_5808,N_9574);
and U11518 (N_11518,N_7102,N_9076);
xor U11519 (N_11519,N_5817,N_7589);
nand U11520 (N_11520,N_6916,N_6186);
and U11521 (N_11521,N_7187,N_8532);
or U11522 (N_11522,N_9536,N_8385);
xnor U11523 (N_11523,N_7852,N_5812);
and U11524 (N_11524,N_7048,N_6152);
xor U11525 (N_11525,N_5384,N_8489);
xnor U11526 (N_11526,N_6539,N_5163);
xnor U11527 (N_11527,N_9969,N_7658);
nor U11528 (N_11528,N_9294,N_6171);
nand U11529 (N_11529,N_8371,N_7105);
or U11530 (N_11530,N_7988,N_8646);
or U11531 (N_11531,N_7547,N_5804);
nor U11532 (N_11532,N_8257,N_9837);
or U11533 (N_11533,N_6589,N_9157);
and U11534 (N_11534,N_5945,N_5203);
and U11535 (N_11535,N_9050,N_8101);
or U11536 (N_11536,N_6307,N_7799);
nor U11537 (N_11537,N_5143,N_9115);
and U11538 (N_11538,N_6136,N_8700);
nor U11539 (N_11539,N_7900,N_8743);
and U11540 (N_11540,N_9430,N_9084);
nor U11541 (N_11541,N_7418,N_8632);
nor U11542 (N_11542,N_8738,N_8194);
xnor U11543 (N_11543,N_9129,N_5438);
and U11544 (N_11544,N_7657,N_6826);
or U11545 (N_11545,N_6120,N_9256);
nor U11546 (N_11546,N_6584,N_9012);
nor U11547 (N_11547,N_5334,N_5909);
xor U11548 (N_11548,N_8995,N_9152);
nor U11549 (N_11549,N_8038,N_5429);
nand U11550 (N_11550,N_5170,N_7450);
nor U11551 (N_11551,N_5780,N_6004);
and U11552 (N_11552,N_5306,N_7412);
or U11553 (N_11553,N_8751,N_8846);
nor U11554 (N_11554,N_5116,N_9302);
or U11555 (N_11555,N_8144,N_6776);
nor U11556 (N_11556,N_9514,N_8238);
nor U11557 (N_11557,N_9503,N_6375);
nand U11558 (N_11558,N_6404,N_9527);
nand U11559 (N_11559,N_9501,N_7820);
and U11560 (N_11560,N_7222,N_6980);
or U11561 (N_11561,N_8766,N_5327);
nor U11562 (N_11562,N_7307,N_8133);
and U11563 (N_11563,N_8986,N_5520);
nor U11564 (N_11564,N_8071,N_7611);
nor U11565 (N_11565,N_8688,N_5705);
or U11566 (N_11566,N_9762,N_7573);
and U11567 (N_11567,N_8540,N_8843);
or U11568 (N_11568,N_5478,N_5744);
nor U11569 (N_11569,N_8124,N_5595);
xnor U11570 (N_11570,N_7653,N_6185);
nand U11571 (N_11571,N_5247,N_7494);
and U11572 (N_11572,N_7254,N_8799);
or U11573 (N_11573,N_9438,N_7760);
or U11574 (N_11574,N_7032,N_7729);
xor U11575 (N_11575,N_7561,N_7442);
or U11576 (N_11576,N_9562,N_7860);
xnor U11577 (N_11577,N_9537,N_6643);
and U11578 (N_11578,N_8906,N_7165);
and U11579 (N_11579,N_9301,N_7666);
or U11580 (N_11580,N_8762,N_6975);
or U11581 (N_11581,N_5838,N_8271);
and U11582 (N_11582,N_9176,N_8417);
nand U11583 (N_11583,N_8503,N_9047);
xor U11584 (N_11584,N_9351,N_7951);
nand U11585 (N_11585,N_7991,N_8010);
or U11586 (N_11586,N_5285,N_7888);
xor U11587 (N_11587,N_5003,N_5402);
and U11588 (N_11588,N_5877,N_7151);
or U11589 (N_11589,N_7947,N_9530);
and U11590 (N_11590,N_9506,N_5745);
or U11591 (N_11591,N_7696,N_7727);
and U11592 (N_11592,N_5684,N_8126);
xnor U11593 (N_11593,N_6330,N_9986);
nor U11594 (N_11594,N_6747,N_5726);
and U11595 (N_11595,N_6810,N_9841);
nor U11596 (N_11596,N_7125,N_8537);
and U11597 (N_11597,N_6744,N_6246);
xor U11598 (N_11598,N_7871,N_5078);
nand U11599 (N_11599,N_6278,N_5010);
xor U11600 (N_11600,N_6220,N_8195);
or U11601 (N_11601,N_6921,N_8316);
nor U11602 (N_11602,N_8029,N_9281);
xor U11603 (N_11603,N_5462,N_8206);
nor U11604 (N_11604,N_5495,N_8923);
nor U11605 (N_11605,N_8660,N_7433);
nand U11606 (N_11606,N_6490,N_6645);
or U11607 (N_11607,N_7789,N_5892);
and U11608 (N_11608,N_5407,N_9370);
and U11609 (N_11609,N_7638,N_7772);
nand U11610 (N_11610,N_9929,N_8131);
nor U11611 (N_11611,N_6735,N_9493);
and U11612 (N_11612,N_8748,N_8531);
nand U11613 (N_11613,N_6170,N_9836);
and U11614 (N_11614,N_6881,N_5803);
xnor U11615 (N_11615,N_5537,N_9916);
nand U11616 (N_11616,N_7574,N_9214);
and U11617 (N_11617,N_7702,N_5733);
nand U11618 (N_11618,N_6665,N_8092);
and U11619 (N_11619,N_8828,N_7694);
nand U11620 (N_11620,N_5392,N_7809);
nand U11621 (N_11621,N_8106,N_8410);
xor U11622 (N_11622,N_9254,N_5642);
nor U11623 (N_11623,N_9038,N_7728);
or U11624 (N_11624,N_7341,N_7587);
xnor U11625 (N_11625,N_8968,N_5681);
nor U11626 (N_11626,N_9210,N_8448);
or U11627 (N_11627,N_6280,N_9011);
nor U11628 (N_11628,N_9887,N_5940);
or U11629 (N_11629,N_7381,N_7238);
nor U11630 (N_11630,N_8673,N_6985);
nor U11631 (N_11631,N_7170,N_7464);
or U11632 (N_11632,N_9835,N_9625);
nor U11633 (N_11633,N_5908,N_8698);
xnor U11634 (N_11634,N_9333,N_7663);
or U11635 (N_11635,N_7840,N_8424);
xnor U11636 (N_11636,N_7455,N_7397);
or U11637 (N_11637,N_5922,N_6802);
nand U11638 (N_11638,N_6309,N_9488);
nor U11639 (N_11639,N_8161,N_7885);
and U11640 (N_11640,N_6612,N_8157);
nor U11641 (N_11641,N_9947,N_9327);
or U11642 (N_11642,N_5086,N_8527);
nand U11643 (N_11643,N_9848,N_7051);
and U11644 (N_11644,N_6833,N_8115);
nor U11645 (N_11645,N_8154,N_9789);
or U11646 (N_11646,N_8689,N_8043);
nand U11647 (N_11647,N_8454,N_5948);
and U11648 (N_11648,N_6745,N_8426);
nand U11649 (N_11649,N_5531,N_7096);
nor U11650 (N_11650,N_9150,N_7490);
or U11651 (N_11651,N_6879,N_5016);
nor U11652 (N_11652,N_6320,N_5999);
nor U11653 (N_11653,N_8786,N_5732);
and U11654 (N_11654,N_8505,N_5990);
and U11655 (N_11655,N_8702,N_9875);
or U11656 (N_11656,N_7430,N_6092);
xnor U11657 (N_11657,N_5513,N_6960);
and U11658 (N_11658,N_6540,N_8772);
xor U11659 (N_11659,N_9015,N_6391);
and U11660 (N_11660,N_9128,N_9131);
nor U11661 (N_11661,N_9108,N_7194);
or U11662 (N_11662,N_6298,N_7710);
nor U11663 (N_11663,N_9580,N_9854);
and U11664 (N_11664,N_9557,N_8036);
or U11665 (N_11665,N_6390,N_5793);
xnor U11666 (N_11666,N_8924,N_5550);
nand U11667 (N_11667,N_9489,N_6122);
and U11668 (N_11668,N_6442,N_7905);
xnor U11669 (N_11669,N_8474,N_5110);
nor U11670 (N_11670,N_7432,N_8399);
xnor U11671 (N_11671,N_7136,N_7184);
xnor U11672 (N_11672,N_9600,N_7053);
and U11673 (N_11673,N_8891,N_8215);
or U11674 (N_11674,N_9133,N_9458);
nor U11675 (N_11675,N_7365,N_8619);
nand U11676 (N_11676,N_9042,N_9260);
xnor U11677 (N_11677,N_9627,N_6590);
nand U11678 (N_11678,N_5284,N_7570);
and U11679 (N_11679,N_6512,N_9349);
and U11680 (N_11680,N_7622,N_6018);
and U11681 (N_11681,N_8998,N_8768);
or U11682 (N_11682,N_5655,N_6772);
xor U11683 (N_11683,N_9207,N_5994);
nand U11684 (N_11684,N_5749,N_5126);
xor U11685 (N_11685,N_9573,N_9653);
nand U11686 (N_11686,N_7331,N_8686);
nor U11687 (N_11687,N_7904,N_8390);
xnor U11688 (N_11688,N_5363,N_5795);
and U11689 (N_11689,N_8850,N_7886);
or U11690 (N_11690,N_5064,N_8042);
and U11691 (N_11691,N_9479,N_9174);
nor U11692 (N_11692,N_6293,N_9416);
and U11693 (N_11693,N_9766,N_9282);
or U11694 (N_11694,N_9917,N_9447);
nand U11695 (N_11695,N_6422,N_6169);
nand U11696 (N_11696,N_7456,N_7531);
nor U11697 (N_11697,N_8674,N_8858);
or U11698 (N_11698,N_6962,N_6033);
xnor U11699 (N_11699,N_5774,N_8351);
nor U11700 (N_11700,N_7685,N_8931);
xor U11701 (N_11701,N_7114,N_8077);
nand U11702 (N_11702,N_7449,N_6690);
nor U11703 (N_11703,N_8360,N_8356);
xnor U11704 (N_11704,N_9932,N_5625);
nand U11705 (N_11705,N_7084,N_6729);
nor U11706 (N_11706,N_7726,N_8273);
nand U11707 (N_11707,N_5115,N_7348);
or U11708 (N_11708,N_9717,N_9182);
xnor U11709 (N_11709,N_6871,N_5133);
nand U11710 (N_11710,N_7730,N_7533);
xor U11711 (N_11711,N_9258,N_9080);
nor U11712 (N_11712,N_7334,N_8528);
or U11713 (N_11713,N_6743,N_9461);
nand U11714 (N_11714,N_9740,N_7788);
or U11715 (N_11715,N_9614,N_7822);
or U11716 (N_11716,N_9332,N_8566);
or U11717 (N_11717,N_7018,N_7778);
xor U11718 (N_11718,N_8321,N_6610);
or U11719 (N_11719,N_5932,N_5516);
nand U11720 (N_11720,N_5703,N_5688);
or U11721 (N_11721,N_9167,N_6983);
nand U11722 (N_11722,N_7327,N_6123);
xor U11723 (N_11723,N_6952,N_6287);
nor U11724 (N_11724,N_9803,N_9512);
nor U11725 (N_11725,N_7175,N_8421);
nor U11726 (N_11726,N_6903,N_6445);
or U11727 (N_11727,N_9616,N_6190);
or U11728 (N_11728,N_9644,N_7540);
and U11729 (N_11729,N_9761,N_9236);
xnor U11730 (N_11730,N_5825,N_7006);
or U11731 (N_11731,N_8623,N_7147);
nor U11732 (N_11732,N_8864,N_6800);
or U11733 (N_11733,N_7089,N_8214);
xor U11734 (N_11734,N_7585,N_9824);
nor U11735 (N_11735,N_7386,N_8023);
nand U11736 (N_11736,N_6180,N_5807);
xnor U11737 (N_11737,N_9502,N_9894);
or U11738 (N_11738,N_7980,N_8475);
nand U11739 (N_11739,N_5633,N_9610);
xnor U11740 (N_11740,N_8112,N_5489);
and U11741 (N_11741,N_6265,N_7746);
nand U11742 (N_11742,N_6947,N_8837);
nor U11743 (N_11743,N_7394,N_7421);
nand U11744 (N_11744,N_9713,N_5916);
xnor U11745 (N_11745,N_6754,N_8943);
nand U11746 (N_11746,N_9340,N_6301);
or U11747 (N_11747,N_5690,N_5670);
xnor U11748 (N_11748,N_6782,N_8061);
nor U11749 (N_11749,N_5823,N_9819);
xnor U11750 (N_11750,N_8192,N_8793);
or U11751 (N_11751,N_7286,N_8134);
xor U11752 (N_11752,N_6614,N_7577);
or U11753 (N_11753,N_6079,N_5172);
nor U11754 (N_11754,N_5200,N_6102);
nand U11755 (N_11755,N_7233,N_8883);
or U11756 (N_11756,N_7406,N_6646);
nand U11757 (N_11757,N_8559,N_5147);
or U11758 (N_11758,N_7295,N_9137);
xor U11759 (N_11759,N_9698,N_9820);
and U11760 (N_11760,N_9880,N_6602);
xnor U11761 (N_11761,N_5036,N_5623);
nor U11762 (N_11762,N_5900,N_8881);
and U11763 (N_11763,N_8979,N_8428);
xnor U11764 (N_11764,N_5185,N_5609);
nor U11765 (N_11765,N_8867,N_5245);
nand U11766 (N_11766,N_8936,N_5676);
xor U11767 (N_11767,N_5820,N_9606);
and U11768 (N_11768,N_6183,N_7268);
and U11769 (N_11769,N_6831,N_5708);
and U11770 (N_11770,N_6948,N_9793);
nand U11771 (N_11771,N_5785,N_7200);
nand U11772 (N_11772,N_9608,N_7899);
nand U11773 (N_11773,N_8001,N_6283);
and U11774 (N_11774,N_9183,N_9960);
or U11775 (N_11775,N_6795,N_8000);
or U11776 (N_11776,N_8655,N_6548);
nand U11777 (N_11777,N_9100,N_6437);
and U11778 (N_11778,N_8926,N_7505);
xor U11779 (N_11779,N_8190,N_8080);
xor U11780 (N_11780,N_6750,N_8961);
and U11781 (N_11781,N_9516,N_5724);
nand U11782 (N_11782,N_5230,N_6625);
xor U11783 (N_11783,N_6371,N_6660);
nor U11784 (N_11784,N_7558,N_7675);
nand U11785 (N_11785,N_6526,N_5410);
and U11786 (N_11786,N_6174,N_9587);
nand U11787 (N_11787,N_6697,N_6857);
and U11788 (N_11788,N_8082,N_8167);
xor U11789 (N_11789,N_6151,N_9219);
xor U11790 (N_11790,N_6574,N_5659);
or U11791 (N_11791,N_5397,N_5777);
and U11792 (N_11792,N_5657,N_9936);
nand U11793 (N_11793,N_6601,N_6579);
and U11794 (N_11794,N_7713,N_8506);
or U11795 (N_11795,N_6101,N_6326);
nor U11796 (N_11796,N_6350,N_7650);
nor U11797 (N_11797,N_5236,N_8616);
and U11798 (N_11798,N_9498,N_8733);
or U11799 (N_11799,N_5654,N_8892);
nor U11800 (N_11800,N_7712,N_9684);
nand U11801 (N_11801,N_5503,N_9892);
nor U11802 (N_11802,N_5755,N_8920);
xor U11803 (N_11803,N_5634,N_7419);
xor U11804 (N_11804,N_7347,N_8767);
nand U11805 (N_11805,N_7104,N_8230);
xnor U11806 (N_11806,N_6938,N_9234);
nand U11807 (N_11807,N_7781,N_6469);
nor U11808 (N_11808,N_5069,N_5562);
or U11809 (N_11809,N_8894,N_5843);
and U11810 (N_11810,N_6543,N_8598);
xnor U11811 (N_11811,N_9549,N_5281);
or U11812 (N_11812,N_5256,N_8464);
and U11813 (N_11813,N_8609,N_5887);
nand U11814 (N_11814,N_5829,N_5278);
or U11815 (N_11815,N_7013,N_7000);
and U11816 (N_11816,N_8731,N_7864);
nor U11817 (N_11817,N_6181,N_8685);
xnor U11818 (N_11818,N_8118,N_7275);
or U11819 (N_11819,N_6409,N_9010);
nor U11820 (N_11820,N_8164,N_9592);
xnor U11821 (N_11821,N_8542,N_6880);
nand U11822 (N_11822,N_8143,N_9545);
xnor U11823 (N_11823,N_6832,N_9485);
nand U11824 (N_11824,N_6449,N_5472);
xor U11825 (N_11825,N_5983,N_5119);
nor U11826 (N_11826,N_7932,N_9279);
and U11827 (N_11827,N_6620,N_8355);
xor U11828 (N_11828,N_9320,N_9812);
or U11829 (N_11829,N_5056,N_8880);
xnor U11830 (N_11830,N_8165,N_5237);
xor U11831 (N_11831,N_5104,N_6333);
nor U11832 (N_11832,N_8469,N_9456);
nand U11833 (N_11833,N_5124,N_7870);
and U11834 (N_11834,N_5917,N_8233);
nor U11835 (N_11835,N_5955,N_5037);
nor U11836 (N_11836,N_6930,N_9985);
or U11837 (N_11837,N_6627,N_5970);
or U11838 (N_11838,N_7370,N_8952);
and U11839 (N_11839,N_5674,N_8222);
xor U11840 (N_11840,N_9362,N_9551);
nand U11841 (N_11841,N_8350,N_6866);
or U11842 (N_11842,N_5120,N_9850);
or U11843 (N_11843,N_8374,N_8064);
nor U11844 (N_11844,N_9003,N_8628);
and U11845 (N_11845,N_5100,N_5882);
or U11846 (N_11846,N_6090,N_6681);
and U11847 (N_11847,N_9118,N_8181);
nor U11848 (N_11848,N_8560,N_9186);
nor U11849 (N_11849,N_5866,N_9354);
nand U11850 (N_11850,N_7816,N_8841);
nor U11851 (N_11851,N_8709,N_5328);
nand U11852 (N_11852,N_6648,N_7420);
nand U11853 (N_11853,N_7819,N_7183);
xnor U11854 (N_11854,N_5518,N_8577);
or U11855 (N_11855,N_6790,N_8791);
xnor U11856 (N_11856,N_9082,N_5176);
or U11857 (N_11857,N_8069,N_9712);
or U11858 (N_11858,N_5440,N_5818);
xnor U11859 (N_11859,N_9939,N_9739);
nand U11860 (N_11860,N_6378,N_7646);
xor U11861 (N_11861,N_7256,N_9396);
or U11862 (N_11862,N_5383,N_9428);
nand U11863 (N_11863,N_6679,N_5364);
nor U11864 (N_11864,N_6756,N_6005);
xor U11865 (N_11865,N_5020,N_8158);
xnor U11866 (N_11866,N_5130,N_5451);
xnor U11867 (N_11867,N_7038,N_8869);
nand U11868 (N_11868,N_5875,N_6863);
or U11869 (N_11869,N_6440,N_6014);
and U11870 (N_11870,N_6502,N_7723);
nand U11871 (N_11871,N_9069,N_5378);
nand U11872 (N_11872,N_5390,N_9474);
xor U11873 (N_11873,N_5546,N_6306);
xor U11874 (N_11874,N_5643,N_7578);
nand U11875 (N_11875,N_9700,N_5058);
and U11876 (N_11876,N_5981,N_7536);
or U11877 (N_11877,N_7500,N_7050);
or U11878 (N_11878,N_5011,N_7792);
nand U11879 (N_11879,N_9291,N_9161);
or U11880 (N_11880,N_8888,N_8656);
or U11881 (N_11881,N_8649,N_8188);
nand U11882 (N_11882,N_5023,N_9731);
and U11883 (N_11883,N_9560,N_8315);
or U11884 (N_11884,N_7801,N_7563);
xor U11885 (N_11885,N_5805,N_7052);
nand U11886 (N_11886,N_6458,N_5450);
or U11887 (N_11887,N_6688,N_6781);
and U11888 (N_11888,N_7841,N_8543);
nor U11889 (N_11889,N_9816,N_9523);
or U11890 (N_11890,N_6432,N_5759);
nand U11891 (N_11891,N_9750,N_7293);
and U11892 (N_11892,N_7215,N_7391);
nand U11893 (N_11893,N_6545,N_5060);
and U11894 (N_11894,N_6053,N_8381);
or U11895 (N_11895,N_5716,N_8179);
nand U11896 (N_11896,N_8955,N_8859);
or U11897 (N_11897,N_6184,N_6662);
nand U11898 (N_11898,N_5936,N_6687);
nor U11899 (N_11899,N_9353,N_7407);
and U11900 (N_11900,N_9000,N_9145);
xor U11901 (N_11901,N_9956,N_6103);
nand U11902 (N_11902,N_6062,N_8045);
and U11903 (N_11903,N_8418,N_9475);
and U11904 (N_11904,N_8059,N_9296);
or U11905 (N_11905,N_9699,N_7623);
xnor U11906 (N_11906,N_8125,N_7193);
nand U11907 (N_11907,N_5262,N_9218);
or U11908 (N_11908,N_6797,N_8836);
nor U11909 (N_11909,N_5142,N_9690);
xnor U11910 (N_11910,N_5502,N_6238);
xnor U11911 (N_11911,N_9344,N_9122);
and U11912 (N_11912,N_6073,N_9873);
or U11913 (N_11913,N_7683,N_9770);
nand U11914 (N_11914,N_7609,N_6084);
nand U11915 (N_11915,N_9679,N_7765);
nand U11916 (N_11916,N_9238,N_7451);
nand U11917 (N_11917,N_5132,N_7940);
nor U11918 (N_11918,N_8298,N_5197);
nand U11919 (N_11919,N_6993,N_7285);
or U11920 (N_11920,N_9066,N_6279);
nand U11921 (N_11921,N_8719,N_5105);
xnor U11922 (N_11922,N_7808,N_8227);
nor U11923 (N_11923,N_9191,N_6710);
nor U11924 (N_11924,N_7468,N_9961);
xor U11925 (N_11925,N_6725,N_8147);
nor U11926 (N_11926,N_6498,N_5570);
nand U11927 (N_11927,N_8207,N_9962);
or U11928 (N_11928,N_8800,N_6961);
or U11929 (N_11929,N_9876,N_9372);
nand U11930 (N_11930,N_8091,N_5575);
nor U11931 (N_11931,N_7426,N_8638);
or U11932 (N_11932,N_6476,N_8073);
nand U11933 (N_11933,N_5182,N_8971);
xnor U11934 (N_11934,N_5207,N_6229);
nand U11935 (N_11935,N_7895,N_6141);
nor U11936 (N_11936,N_9243,N_5535);
and U11937 (N_11937,N_6219,N_5985);
xnor U11938 (N_11938,N_7866,N_8579);
nand U11939 (N_11939,N_6777,N_7247);
xor U11940 (N_11940,N_5279,N_8575);
xor U11941 (N_11941,N_7827,N_9583);
nand U11942 (N_11942,N_7502,N_5557);
and U11943 (N_11943,N_5250,N_8951);
xnor U11944 (N_11944,N_6160,N_7178);
nand U11945 (N_11945,N_6367,N_5534);
nor U11946 (N_11946,N_6769,N_7845);
nor U11947 (N_11947,N_6434,N_6026);
nor U11948 (N_11948,N_9567,N_5648);
nand U11949 (N_11949,N_5802,N_6704);
and U11950 (N_11950,N_8522,N_6669);
nor U11951 (N_11951,N_6926,N_6605);
and U11952 (N_11952,N_9678,N_7725);
nand U11953 (N_11953,N_7692,N_6060);
nor U11954 (N_11954,N_7634,N_7411);
and U11955 (N_11955,N_7962,N_6897);
or U11956 (N_11956,N_9781,N_9757);
nand U11957 (N_11957,N_9121,N_8248);
nor U11958 (N_11958,N_5291,N_5373);
nand U11959 (N_11959,N_5566,N_6796);
and U11960 (N_11960,N_5319,N_9710);
xor U11961 (N_11961,N_9637,N_7201);
and U11962 (N_11962,N_6023,N_8965);
nor U11963 (N_11963,N_8722,N_5348);
nand U11964 (N_11964,N_9733,N_9360);
nand U11965 (N_11965,N_8366,N_5215);
and U11966 (N_11966,N_8742,N_5183);
xor U11967 (N_11967,N_5832,N_9804);
nand U11968 (N_11968,N_6112,N_7027);
or U11969 (N_11969,N_6696,N_8412);
and U11970 (N_11970,N_6973,N_7243);
nand U11971 (N_11971,N_8487,N_6506);
xor U11972 (N_11972,N_6585,N_8615);
xnor U11973 (N_11973,N_6208,N_5971);
and U11974 (N_11974,N_9252,N_5555);
nor U11975 (N_11975,N_6807,N_5761);
and U11976 (N_11976,N_7487,N_9390);
and U11977 (N_11977,N_7135,N_7708);
xor U11978 (N_11978,N_5910,N_7736);
nor U11979 (N_11979,N_9444,N_5466);
and U11980 (N_11980,N_6521,N_5835);
nor U11981 (N_11981,N_7234,N_8782);
or U11982 (N_11982,N_6845,N_7392);
nand U11983 (N_11983,N_5053,N_8750);
or U11984 (N_11984,N_5519,N_8263);
nor U11985 (N_11985,N_8919,N_9856);
and U11986 (N_11986,N_7055,N_6484);
and U11987 (N_11987,N_8659,N_6830);
xor U11988 (N_11988,N_6157,N_8854);
and U11989 (N_11989,N_6684,N_8613);
and U11990 (N_11990,N_7784,N_7121);
and U11991 (N_11991,N_6569,N_6273);
xnor U11992 (N_11992,N_8396,N_7063);
and U11993 (N_11993,N_6348,N_7160);
nor U11994 (N_11994,N_7404,N_6039);
and U11995 (N_11995,N_9631,N_6044);
nor U11996 (N_11996,N_8228,N_7583);
and U11997 (N_11997,N_8148,N_7739);
xnor U11998 (N_11998,N_7510,N_6294);
nand U11999 (N_11999,N_8338,N_9890);
or U12000 (N_12000,N_5375,N_8825);
nor U12001 (N_12001,N_8904,N_5652);
or U12002 (N_12002,N_5093,N_8908);
and U12003 (N_12003,N_5140,N_6413);
xnor U12004 (N_12004,N_6641,N_6036);
xnor U12005 (N_12005,N_6705,N_9160);
and U12006 (N_12006,N_6616,N_5258);
xor U12007 (N_12007,N_7043,N_9452);
xnor U12008 (N_12008,N_8714,N_6716);
and U12009 (N_12009,N_8618,N_5834);
xor U12010 (N_12010,N_9180,N_7944);
or U12011 (N_12011,N_7542,N_7641);
and U12012 (N_12012,N_9525,N_5500);
nor U12013 (N_12013,N_9077,N_6909);
and U12014 (N_12014,N_6588,N_7552);
and U12015 (N_12015,N_8309,N_7857);
nand U12016 (N_12016,N_7488,N_7226);
or U12017 (N_12017,N_5735,N_9057);
nand U12018 (N_12018,N_8093,N_7633);
xor U12019 (N_12019,N_8994,N_7242);
nand U12020 (N_12020,N_5637,N_5593);
xnor U12021 (N_12021,N_6520,N_8110);
nor U12022 (N_12022,N_7384,N_7701);
nor U12023 (N_12023,N_6356,N_9635);
nor U12024 (N_12024,N_9318,N_5646);
nor U12025 (N_12025,N_9691,N_5453);
nor U12026 (N_12026,N_9827,N_5066);
nor U12027 (N_12027,N_9304,N_9054);
and U12028 (N_12028,N_8586,N_5976);
and U12029 (N_12029,N_6651,N_5687);
nand U12030 (N_12030,N_8367,N_8853);
nor U12031 (N_12031,N_9231,N_7768);
nand U12032 (N_12032,N_7997,N_8151);
nand U12033 (N_12033,N_7906,N_6380);
and U12034 (N_12034,N_6365,N_8977);
xor U12035 (N_12035,N_9229,N_5924);
nand U12036 (N_12036,N_9466,N_8402);
nand U12037 (N_12037,N_5540,N_8807);
nor U12038 (N_12038,N_9943,N_9544);
and U12039 (N_12039,N_6734,N_6558);
nand U12040 (N_12040,N_8171,N_9993);
xnor U12041 (N_12041,N_6431,N_6550);
xor U12042 (N_12042,N_6893,N_6068);
and U12043 (N_12043,N_7328,N_6989);
or U12044 (N_12044,N_5627,N_7617);
and U12045 (N_12045,N_9924,N_7607);
nand U12046 (N_12046,N_5578,N_9039);
nand U12047 (N_12047,N_7811,N_5419);
nor U12048 (N_12048,N_7378,N_7157);
and U12049 (N_12049,N_8988,N_7566);
nor U12050 (N_12050,N_8145,N_6510);
xor U12051 (N_12051,N_8886,N_7605);
nor U12052 (N_12052,N_6572,N_8284);
or U12053 (N_12053,N_8897,N_7749);
xor U12054 (N_12054,N_6715,N_8249);
xor U12055 (N_12055,N_5864,N_9384);
nor U12056 (N_12056,N_6032,N_7122);
xor U12057 (N_12057,N_8359,N_6598);
nor U12058 (N_12058,N_9907,N_6834);
and U12059 (N_12059,N_7917,N_9701);
or U12060 (N_12060,N_5734,N_6541);
or U12061 (N_12061,N_7173,N_8193);
xor U12062 (N_12062,N_8572,N_7486);
nor U12063 (N_12063,N_6755,N_7743);
or U12064 (N_12064,N_8065,N_7267);
nand U12065 (N_12065,N_8375,N_6650);
nor U12066 (N_12066,N_6578,N_5282);
or U12067 (N_12067,N_7876,N_9734);
or U12068 (N_12068,N_8713,N_9203);
nand U12069 (N_12069,N_5669,N_6156);
or U12070 (N_12070,N_6085,N_7724);
or U12071 (N_12071,N_5704,N_7413);
nor U12072 (N_12072,N_5743,N_8610);
nand U12073 (N_12073,N_5464,N_7335);
and U12074 (N_12074,N_7377,N_8174);
or U12075 (N_12075,N_5032,N_9107);
xnor U12076 (N_12076,N_5345,N_5925);
nor U12077 (N_12077,N_8633,N_7936);
xor U12078 (N_12078,N_5457,N_7204);
and U12079 (N_12079,N_7528,N_8974);
and U12080 (N_12080,N_5878,N_7709);
nand U12081 (N_12081,N_6048,N_9675);
nor U12082 (N_12082,N_8450,N_6105);
or U12083 (N_12083,N_8152,N_7939);
and U12084 (N_12084,N_6133,N_6177);
nand U12085 (N_12085,N_6487,N_9286);
or U12086 (N_12086,N_8785,N_6041);
nor U12087 (N_12087,N_7270,N_7255);
or U12088 (N_12088,N_6658,N_9055);
nand U12089 (N_12089,N_9928,N_8644);
xor U12090 (N_12090,N_7434,N_7635);
nand U12091 (N_12091,N_9783,N_9098);
nor U12092 (N_12092,N_6096,N_6155);
and U12093 (N_12093,N_7428,N_8049);
nand U12094 (N_12094,N_6412,N_5541);
and U12095 (N_12095,N_5443,N_8055);
nand U12096 (N_12096,N_6576,N_8627);
nor U12097 (N_12097,N_9364,N_5509);
nand U12098 (N_12098,N_7283,N_6260);
nand U12099 (N_12099,N_6107,N_7344);
nor U12100 (N_12100,N_9120,N_8005);
nand U12101 (N_12101,N_6623,N_7981);
and U12102 (N_12102,N_5799,N_7497);
or U12103 (N_12103,N_8320,N_6478);
nand U12104 (N_12104,N_5702,N_5841);
nand U12105 (N_12105,N_7146,N_8272);
nor U12106 (N_12106,N_9409,N_8672);
nand U12107 (N_12107,N_6040,N_8392);
and U12108 (N_12108,N_8969,N_5357);
and U12109 (N_12109,N_5222,N_7369);
nand U12110 (N_12110,N_5656,N_5352);
and U12111 (N_12111,N_7893,N_6231);
or U12112 (N_12112,N_9355,N_5723);
nand U12113 (N_12113,N_7257,N_7517);
and U12114 (N_12114,N_7844,N_8557);
xnor U12115 (N_12115,N_6488,N_7545);
xnor U12116 (N_12116,N_5296,N_6765);
xor U12117 (N_12117,N_8737,N_6732);
or U12118 (N_12118,N_9949,N_8736);
nor U12119 (N_12119,N_6860,N_6049);
or U12120 (N_12120,N_9613,N_9755);
nand U12121 (N_12121,N_7356,N_8015);
and U12122 (N_12122,N_9689,N_6699);
or U12123 (N_12123,N_8578,N_5806);
nor U12124 (N_12124,N_9073,N_9520);
and U12125 (N_12125,N_5346,N_7751);
or U12126 (N_12126,N_7777,N_7515);
nand U12127 (N_12127,N_9568,N_7036);
and U12128 (N_12128,N_8442,N_8911);
or U12129 (N_12129,N_8340,N_7023);
and U12130 (N_12130,N_8795,N_6194);
xor U12131 (N_12131,N_8844,N_9259);
nand U12132 (N_12132,N_6149,N_7914);
or U12133 (N_12133,N_6522,N_6211);
xnor U12134 (N_12134,N_8734,N_9822);
and U12135 (N_12135,N_5293,N_7366);
nand U12136 (N_12136,N_8956,N_5617);
nor U12137 (N_12137,N_7229,N_7263);
or U12138 (N_12138,N_9021,N_9288);
nand U12139 (N_12139,N_5122,N_8310);
nand U12140 (N_12140,N_7732,N_5527);
nand U12141 (N_12141,N_8094,N_9499);
nand U12142 (N_12142,N_5845,N_7156);
and U12143 (N_12143,N_6021,N_8013);
and U12144 (N_12144,N_5321,N_7287);
xor U12145 (N_12145,N_9423,N_7422);
nor U12146 (N_12146,N_6212,N_9140);
or U12147 (N_12147,N_6467,N_8476);
or U12148 (N_12148,N_6421,N_6003);
or U12149 (N_12149,N_7737,N_8240);
xnor U12150 (N_12150,N_8693,N_7099);
nor U12151 (N_12151,N_9297,N_7100);
nor U12152 (N_12152,N_8893,N_6999);
and U12153 (N_12153,N_5947,N_7350);
nand U12154 (N_12154,N_9482,N_9060);
or U12155 (N_12155,N_8992,N_8006);
or U12156 (N_12156,N_8076,N_7834);
or U12157 (N_12157,N_6891,N_5156);
xnor U12158 (N_12158,N_5359,N_7154);
and U12159 (N_12159,N_7901,N_9336);
and U12160 (N_12160,N_5006,N_9622);
nand U12161 (N_12161,N_8095,N_7308);
and U12162 (N_12162,N_5998,N_5025);
nand U12163 (N_12163,N_5483,N_8141);
nand U12164 (N_12164,N_5015,N_7339);
nor U12165 (N_12165,N_9465,N_6494);
nand U12166 (N_12166,N_5198,N_8247);
xnor U12167 (N_12167,N_7258,N_9759);
and U12168 (N_12168,N_8130,N_8541);
nand U12169 (N_12169,N_8696,N_5580);
nand U12170 (N_12170,N_8983,N_9242);
or U12171 (N_12171,N_8162,N_5547);
nor U12172 (N_12172,N_9830,N_5486);
nand U12173 (N_12173,N_9657,N_7059);
or U12174 (N_12174,N_9628,N_5199);
xor U12175 (N_12175,N_8105,N_9513);
and U12176 (N_12176,N_9674,N_5286);
xnor U12177 (N_12177,N_5201,N_9594);
nand U12178 (N_12178,N_8651,N_5632);
xnor U12179 (N_12179,N_7523,N_6910);
or U12180 (N_12180,N_5114,N_9846);
nor U12181 (N_12181,N_7351,N_6162);
nand U12182 (N_12182,N_8119,N_6657);
xor U12183 (N_12183,N_6244,N_8976);
nand U12184 (N_12184,N_7773,N_5944);
xnor U12185 (N_12185,N_6656,N_7632);
xnor U12186 (N_12186,N_6203,N_6820);
and U12187 (N_12187,N_6823,N_8114);
and U12188 (N_12188,N_6787,N_7806);
and U12189 (N_12189,N_8306,N_9262);
nor U12190 (N_12190,N_9834,N_9216);
nor U12191 (N_12191,N_8074,N_5821);
nor U12192 (N_12192,N_8354,N_6282);
and U12193 (N_12193,N_7787,N_6025);
nand U12194 (N_12194,N_5452,N_9671);
nor U12195 (N_12195,N_5193,N_7873);
nand U12196 (N_12196,N_9893,N_5310);
or U12197 (N_12197,N_5300,N_7437);
xor U12198 (N_12198,N_9685,N_7467);
nor U12199 (N_12199,N_9072,N_7550);
nor U12200 (N_12200,N_8611,N_5244);
and U12201 (N_12201,N_6559,N_8099);
nor U12202 (N_12202,N_6235,N_8416);
or U12203 (N_12203,N_7040,N_6519);
nand U12204 (N_12204,N_7498,N_9027);
xor U12205 (N_12205,N_6617,N_5195);
and U12206 (N_12206,N_7395,N_7101);
xnor U12207 (N_12207,N_7123,N_7610);
nor U12208 (N_12208,N_6901,N_7231);
nand U12209 (N_12209,N_8244,N_6843);
nor U12210 (N_12210,N_8668,N_9469);
nand U12211 (N_12211,N_9971,N_9885);
nor U12212 (N_12212,N_8912,N_9347);
xor U12213 (N_12213,N_5405,N_7891);
nor U12214 (N_12214,N_8172,N_9914);
or U12215 (N_12215,N_7652,N_8861);
and U12216 (N_12216,N_7984,N_7700);
or U12217 (N_12217,N_7798,N_6400);
nor U12218 (N_12218,N_8857,N_7527);
nand U12219 (N_12219,N_7473,N_5192);
nand U12220 (N_12220,N_9392,N_7688);
xor U12221 (N_12221,N_8932,N_9307);
nor U12222 (N_12222,N_5926,N_7436);
and U12223 (N_12223,N_5330,N_9052);
xor U12224 (N_12224,N_6691,N_7879);
or U12225 (N_12225,N_6113,N_7481);
or U12226 (N_12226,N_6161,N_9981);
or U12227 (N_12227,N_8163,N_8945);
or U12228 (N_12228,N_8730,N_7302);
or U12229 (N_12229,N_6114,N_7649);
and U12230 (N_12230,N_7217,N_8771);
and U12231 (N_12231,N_5049,N_7143);
or U12232 (N_12232,N_6882,N_8200);
nor U12233 (N_12233,N_5274,N_8510);
nor U12234 (N_12234,N_9181,N_8718);
nor U12235 (N_12235,N_5563,N_9178);
nand U12236 (N_12236,N_7511,N_8948);
nand U12237 (N_12237,N_5536,N_8832);
nand U12238 (N_12238,N_6611,N_6249);
nor U12239 (N_12239,N_7875,N_7546);
xnor U12240 (N_12240,N_9708,N_6269);
and U12241 (N_12241,N_5442,N_7317);
nor U12242 (N_12242,N_7847,N_7252);
nor U12243 (N_12243,N_9379,N_6746);
nor U12244 (N_12244,N_6629,N_5667);
nand U12245 (N_12245,N_5343,N_5800);
nand U12246 (N_12246,N_7964,N_8216);
nand U12247 (N_12247,N_9442,N_9776);
nor U12248 (N_12248,N_8028,N_7828);
and U12249 (N_12249,N_9706,N_7733);
nand U12250 (N_12250,N_6338,N_8294);
or U12251 (N_12251,N_7045,N_8856);
nor U12252 (N_12252,N_6230,N_5756);
xor U12253 (N_12253,N_9223,N_6388);
or U12254 (N_12254,N_9780,N_8665);
nand U12255 (N_12255,N_8717,N_8456);
nand U12256 (N_12256,N_8938,N_6988);
nand U12257 (N_12257,N_7603,N_9984);
xor U12258 (N_12258,N_8871,N_8083);
and U12259 (N_12259,N_8295,N_6256);
xor U12260 (N_12260,N_7152,N_6364);
nor U12261 (N_12261,N_5229,N_8269);
nand U12262 (N_12262,N_9752,N_9529);
nand U12263 (N_12263,N_6086,N_7259);
nor U12264 (N_12264,N_9773,N_8902);
or U12265 (N_12265,N_5189,N_9900);
xnor U12266 (N_12266,N_6896,N_7079);
nor U12267 (N_12267,N_8266,N_9741);
nand U12268 (N_12268,N_9758,N_7912);
xnor U12269 (N_12269,N_6892,N_8477);
and U12270 (N_12270,N_9460,N_9316);
and U12271 (N_12271,N_7695,N_9612);
and U12272 (N_12272,N_5775,N_9661);
nor U12273 (N_12273,N_8703,N_8357);
xnor U12274 (N_12274,N_9898,N_7373);
nand U12275 (N_12275,N_7212,N_6847);
xnor U12276 (N_12276,N_8378,N_6873);
nor U12277 (N_12277,N_6516,N_6698);
nand U12278 (N_12278,N_9883,N_7790);
or U12279 (N_12279,N_8821,N_8287);
nand U12280 (N_12280,N_8372,N_6945);
or U12281 (N_12281,N_8311,N_9083);
nand U12282 (N_12282,N_8407,N_7005);
nand U12283 (N_12283,N_5324,N_8661);
nand U12284 (N_12284,N_8667,N_6443);
and U12285 (N_12285,N_9290,N_5605);
nor U12286 (N_12286,N_8236,N_7682);
nor U12287 (N_12287,N_6331,N_8377);
nor U12288 (N_12288,N_8419,N_7759);
xnor U12289 (N_12289,N_8589,N_6982);
nand U12290 (N_12290,N_7235,N_6403);
and U12291 (N_12291,N_9609,N_9874);
nor U12292 (N_12292,N_5108,N_7333);
nand U12293 (N_12293,N_6849,N_6609);
and U12294 (N_12294,N_5118,N_5614);
nor U12295 (N_12295,N_7994,N_7717);
nand U12296 (N_12296,N_9276,N_8150);
and U12297 (N_12297,N_9889,N_6165);
nor U12298 (N_12298,N_7592,N_9718);
nand U12299 (N_12299,N_7887,N_8160);
nand U12300 (N_12300,N_6534,N_8256);
and U12301 (N_12301,N_6485,N_8411);
and U12302 (N_12302,N_5268,N_8498);
nand U12303 (N_12303,N_7813,N_7186);
or U12304 (N_12304,N_9079,N_8645);
nand U12305 (N_12305,N_6621,N_8518);
and U12306 (N_12306,N_9378,N_5184);
nand U12307 (N_12307,N_6099,N_9541);
nor U12308 (N_12308,N_9570,N_8597);
or U12309 (N_12309,N_8914,N_6649);
nor U12310 (N_12310,N_8697,N_6818);
nand U12311 (N_12311,N_5933,N_6195);
xor U12312 (N_12312,N_9230,N_7002);
xor U12313 (N_12313,N_9726,N_6546);
and U12314 (N_12314,N_6483,N_8046);
nand U12315 (N_12315,N_9239,N_7934);
nand U12316 (N_12316,N_8996,N_5165);
or U12317 (N_12317,N_8465,N_5682);
and U12318 (N_12318,N_9558,N_6946);
nand U12319 (N_12319,N_9794,N_9030);
and U12320 (N_12320,N_6972,N_6226);
xor U12321 (N_12321,N_8358,N_5600);
nor U12322 (N_12322,N_8349,N_7923);
and U12323 (N_12323,N_5554,N_8401);
and U12324 (N_12324,N_6322,N_6872);
nor U12325 (N_12325,N_5235,N_8629);
xnor U12326 (N_12326,N_7754,N_9732);
and U12327 (N_12327,N_9406,N_8526);
and U12328 (N_12328,N_9272,N_6175);
or U12329 (N_12329,N_8056,N_7882);
nand U12330 (N_12330,N_9427,N_5847);
and U12331 (N_12331,N_9738,N_6931);
xor U12332 (N_12332,N_7330,N_7785);
or U12333 (N_12333,N_9640,N_9046);
xnor U12334 (N_12334,N_7262,N_9371);
nor U12335 (N_12335,N_8855,N_9417);
or U12336 (N_12336,N_7429,N_7300);
nand U12337 (N_12337,N_5276,N_5883);
xnor U12338 (N_12338,N_9348,N_5965);
and U12339 (N_12339,N_7182,N_8201);
nor U12340 (N_12340,N_6187,N_7189);
and U12341 (N_12341,N_6730,N_6518);
and U12342 (N_12342,N_6222,N_8330);
xnor U12343 (N_12343,N_9449,N_9037);
or U12344 (N_12344,N_5290,N_8490);
nor U12345 (N_12345,N_9144,N_6537);
nand U12346 (N_12346,N_6405,N_6536);
xnor U12347 (N_12347,N_8136,N_5772);
and U12348 (N_12348,N_5152,N_8225);
or U12349 (N_12349,N_7272,N_6803);
and U12350 (N_12350,N_6859,N_6424);
nor U12351 (N_12351,N_8149,N_5661);
and U12352 (N_12352,N_9754,N_8599);
xor U12353 (N_12353,N_8820,N_6075);
or U12354 (N_12354,N_9074,N_6640);
nand U12355 (N_12355,N_7501,N_5424);
and U12356 (N_12356,N_6221,N_6835);
nand U12357 (N_12357,N_8567,N_6150);
nor U12358 (N_12358,N_9212,N_9339);
or U12359 (N_12359,N_6473,N_6886);
and U12360 (N_12360,N_9860,N_7995);
xor U12361 (N_12361,N_9974,N_9198);
nand U12362 (N_12362,N_8838,N_9991);
xnor U12363 (N_12363,N_5689,N_6770);
xnor U12364 (N_12364,N_5714,N_9799);
or U12365 (N_12365,N_6197,N_9226);
xnor U12366 (N_12366,N_5491,N_5815);
xor U12367 (N_12367,N_5615,N_9704);
and U12368 (N_12368,N_6327,N_5898);
nor U12369 (N_12369,N_9126,N_7771);
or U12370 (N_12370,N_9995,N_6596);
nand U12371 (N_12371,N_9771,N_6718);
or U12372 (N_12372,N_5481,N_8966);
xnor U12373 (N_12373,N_5080,N_9263);
nor U12374 (N_12374,N_7651,N_6749);
or U12375 (N_12375,N_8770,N_6481);
or U12376 (N_12376,N_7933,N_6954);
and U12377 (N_12377,N_6722,N_8798);
xnor U12378 (N_12378,N_8849,N_6742);
xnor U12379 (N_12379,N_8639,N_6549);
nand U12380 (N_12380,N_5034,N_8169);
and U12381 (N_12381,N_7138,N_8981);
nand U12382 (N_12382,N_7236,N_7313);
nand U12383 (N_12383,N_9814,N_9184);
or U12384 (N_12384,N_5107,N_9480);
and U12385 (N_12385,N_7248,N_6856);
or U12386 (N_12386,N_9751,N_5041);
nor U12387 (N_12387,N_5381,N_5349);
nor U12388 (N_12388,N_8520,N_8928);
nor U12389 (N_12389,N_7965,N_9177);
nand U12390 (N_12390,N_9805,N_9839);
or U12391 (N_12391,N_6240,N_8183);
nor U12392 (N_12392,N_8137,N_5109);
and U12393 (N_12393,N_5000,N_8954);
and U12394 (N_12394,N_8121,N_6533);
nor U12395 (N_12395,N_9821,N_7264);
xnor U12396 (N_12396,N_8007,N_9143);
and U12397 (N_12397,N_8934,N_7680);
nor U12398 (N_12398,N_8267,N_7080);
nand U12399 (N_12399,N_5432,N_7818);
and U12400 (N_12400,N_5426,N_7066);
or U12401 (N_12401,N_7757,N_6119);
xnor U12402 (N_12402,N_8452,N_7629);
nand U12403 (N_12403,N_5356,N_8332);
nand U12404 (N_12404,N_6652,N_6254);
and U12405 (N_12405,N_9454,N_9085);
nor U12406 (N_12406,N_9564,N_5305);
xor U12407 (N_12407,N_5814,N_6918);
xor U12408 (N_12408,N_7058,N_9205);
nor U12409 (N_12409,N_7869,N_5608);
or U12410 (N_12410,N_8640,N_5074);
nand U12411 (N_12411,N_8903,N_6761);
nand U12412 (N_12412,N_6727,N_6489);
nor U12413 (N_12413,N_7758,N_6870);
or U12414 (N_12414,N_5816,N_5913);
or U12415 (N_12415,N_6819,N_8692);
and U12416 (N_12416,N_5009,N_9497);
or U12417 (N_12417,N_9188,N_7297);
nand U12418 (N_12418,N_6808,N_6667);
and U12419 (N_12419,N_8322,N_7706);
nand U12420 (N_12420,N_6387,N_5731);
nand U12421 (N_12421,N_5326,N_5353);
or U12422 (N_12422,N_7095,N_7112);
or U12423 (N_12423,N_9861,N_8763);
and U12424 (N_12424,N_5911,N_7843);
and U12425 (N_12425,N_6775,N_7320);
and U12426 (N_12426,N_7094,N_7319);
nand U12427 (N_12427,N_5951,N_5340);
or U12428 (N_12428,N_9453,N_8078);
nor U12429 (N_12429,N_8047,N_9245);
nand U12430 (N_12430,N_8127,N_5867);
nand U12431 (N_12431,N_9020,N_5174);
or U12432 (N_12432,N_8117,N_6904);
or U12433 (N_12433,N_5942,N_8471);
xor U12434 (N_12434,N_5574,N_6990);
or U12435 (N_12435,N_9099,N_7478);
xnor U12436 (N_12436,N_8323,N_6052);
nand U12437 (N_12437,N_9338,N_9034);
xnor U12438 (N_12438,N_5135,N_9646);
nor U12439 (N_12439,N_8715,N_5196);
and U12440 (N_12440,N_6224,N_5995);
nand U12441 (N_12441,N_7956,N_6758);
nand U12442 (N_12442,N_6217,N_8384);
nor U12443 (N_12443,N_5401,N_5665);
nor U12444 (N_12444,N_9550,N_7056);
and U12445 (N_12445,N_6216,N_5618);
nor U12446 (N_12446,N_5510,N_8395);
nand U12447 (N_12447,N_5579,N_5420);
xnor U12448 (N_12448,N_5127,N_9448);
or U12449 (N_12449,N_5741,N_6359);
nor U12450 (N_12450,N_8740,N_6121);
xor U12451 (N_12451,N_5028,N_6995);
xor U12452 (N_12452,N_6340,N_9342);
nand U12453 (N_12453,N_8625,N_6925);
nand U12454 (N_12454,N_5437,N_5819);
nor U12455 (N_12455,N_8501,N_7846);
nand U12456 (N_12456,N_8051,N_7902);
or U12457 (N_12457,N_7920,N_6634);
xnor U12458 (N_12458,N_9232,N_6741);
nor U12459 (N_12459,N_5629,N_9013);
or U12460 (N_12460,N_8797,N_5295);
nand U12461 (N_12461,N_7943,N_8918);
or U12462 (N_12462,N_6355,N_8887);
xnor U12463 (N_12463,N_8261,N_7168);
nand U12464 (N_12464,N_8347,N_9110);
nand U12465 (N_12465,N_6059,N_7127);
and U12466 (N_12466,N_9665,N_6685);
nand U12467 (N_12467,N_5711,N_9518);
and U12468 (N_12468,N_9109,N_9802);
or U12469 (N_12469,N_6635,N_8666);
xnor U12470 (N_12470,N_7982,N_5444);
xor U12471 (N_12471,N_8468,N_9853);
and U12472 (N_12472,N_9175,N_5597);
and U12473 (N_12473,N_9431,N_6566);
xnor U12474 (N_12474,N_5342,N_6050);
and U12475 (N_12475,N_5387,N_9094);
and U12476 (N_12476,N_8812,N_5677);
xnor U12477 (N_12477,N_9909,N_5698);
or U12478 (N_12478,N_6193,N_7584);
and U12479 (N_12479,N_7224,N_9539);
nor U12480 (N_12480,N_7913,N_6020);
and U12481 (N_12481,N_8663,N_6411);
nor U12482 (N_12482,N_7925,N_6054);
nand U12483 (N_12483,N_8909,N_8957);
or U12484 (N_12484,N_6853,N_7596);
and U12485 (N_12485,N_8363,N_5930);
nand U12486 (N_12486,N_8921,N_6608);
nand U12487 (N_12487,N_9975,N_8414);
and U12488 (N_12488,N_5758,N_7786);
xor U12489 (N_12489,N_6964,N_8302);
or U12490 (N_12490,N_8558,N_7720);
or U12491 (N_12491,N_7532,N_9593);
nor U12492 (N_12492,N_7586,N_6022);
or U12493 (N_12493,N_8681,N_8170);
or U12494 (N_12494,N_5750,N_8778);
and U12495 (N_12495,N_8324,N_5138);
and U12496 (N_12496,N_8690,N_9858);
nand U12497 (N_12497,N_6986,N_6798);
nand U12498 (N_12498,N_5722,N_9664);
and U12499 (N_12499,N_7363,N_6321);
xnor U12500 (N_12500,N_5783,N_6197);
xnor U12501 (N_12501,N_8670,N_7412);
xnor U12502 (N_12502,N_7732,N_6431);
xor U12503 (N_12503,N_6231,N_7233);
xnor U12504 (N_12504,N_6262,N_7109);
xnor U12505 (N_12505,N_5226,N_5409);
or U12506 (N_12506,N_9746,N_7219);
nand U12507 (N_12507,N_7807,N_5155);
xor U12508 (N_12508,N_9137,N_7032);
xor U12509 (N_12509,N_8633,N_9679);
or U12510 (N_12510,N_8928,N_8876);
xnor U12511 (N_12511,N_8964,N_8186);
nand U12512 (N_12512,N_8795,N_7270);
and U12513 (N_12513,N_7687,N_6906);
xor U12514 (N_12514,N_9463,N_8744);
nor U12515 (N_12515,N_9291,N_8295);
xnor U12516 (N_12516,N_9278,N_6958);
and U12517 (N_12517,N_5813,N_8885);
nor U12518 (N_12518,N_9525,N_7073);
nor U12519 (N_12519,N_7223,N_5631);
or U12520 (N_12520,N_9533,N_7243);
and U12521 (N_12521,N_6421,N_9869);
xor U12522 (N_12522,N_7813,N_7880);
xor U12523 (N_12523,N_6138,N_6410);
and U12524 (N_12524,N_6070,N_9973);
or U12525 (N_12525,N_5357,N_8857);
nor U12526 (N_12526,N_7852,N_5539);
xor U12527 (N_12527,N_9308,N_9604);
and U12528 (N_12528,N_6841,N_5687);
nand U12529 (N_12529,N_7944,N_7194);
xor U12530 (N_12530,N_7857,N_6058);
nor U12531 (N_12531,N_5664,N_9715);
nand U12532 (N_12532,N_7433,N_7197);
xor U12533 (N_12533,N_8010,N_5624);
or U12534 (N_12534,N_5887,N_8838);
and U12535 (N_12535,N_7971,N_6561);
xor U12536 (N_12536,N_6792,N_7306);
xor U12537 (N_12537,N_9262,N_8247);
nand U12538 (N_12538,N_6023,N_6481);
xor U12539 (N_12539,N_6079,N_6388);
nor U12540 (N_12540,N_5440,N_8645);
and U12541 (N_12541,N_9522,N_8527);
nand U12542 (N_12542,N_9920,N_6468);
nand U12543 (N_12543,N_7276,N_5063);
or U12544 (N_12544,N_8020,N_6344);
or U12545 (N_12545,N_6641,N_8868);
xnor U12546 (N_12546,N_9651,N_5735);
and U12547 (N_12547,N_6513,N_8035);
xor U12548 (N_12548,N_7595,N_7471);
nand U12549 (N_12549,N_5056,N_9804);
or U12550 (N_12550,N_7062,N_5982);
nand U12551 (N_12551,N_6562,N_6202);
or U12552 (N_12552,N_7883,N_9372);
nor U12553 (N_12553,N_5005,N_7294);
nor U12554 (N_12554,N_6900,N_7267);
nand U12555 (N_12555,N_9425,N_5608);
nor U12556 (N_12556,N_7077,N_9288);
or U12557 (N_12557,N_8577,N_5378);
nand U12558 (N_12558,N_7878,N_8313);
and U12559 (N_12559,N_5412,N_8360);
and U12560 (N_12560,N_8323,N_9549);
xor U12561 (N_12561,N_5193,N_6641);
or U12562 (N_12562,N_5282,N_6694);
and U12563 (N_12563,N_7023,N_6343);
nor U12564 (N_12564,N_9710,N_7956);
and U12565 (N_12565,N_8980,N_9271);
or U12566 (N_12566,N_8942,N_5753);
or U12567 (N_12567,N_6028,N_8346);
or U12568 (N_12568,N_8327,N_7965);
and U12569 (N_12569,N_8913,N_8925);
and U12570 (N_12570,N_9820,N_9372);
or U12571 (N_12571,N_7586,N_7722);
nor U12572 (N_12572,N_9936,N_9692);
and U12573 (N_12573,N_8105,N_6100);
and U12574 (N_12574,N_9604,N_6902);
or U12575 (N_12575,N_5733,N_6459);
nand U12576 (N_12576,N_6690,N_5798);
or U12577 (N_12577,N_8658,N_8453);
nand U12578 (N_12578,N_5470,N_8483);
xor U12579 (N_12579,N_6642,N_6427);
and U12580 (N_12580,N_5657,N_9171);
xor U12581 (N_12581,N_5895,N_9941);
nor U12582 (N_12582,N_9046,N_8361);
and U12583 (N_12583,N_8280,N_6369);
or U12584 (N_12584,N_7316,N_6215);
nor U12585 (N_12585,N_7462,N_8578);
nor U12586 (N_12586,N_6131,N_7060);
nand U12587 (N_12587,N_7209,N_9068);
and U12588 (N_12588,N_6322,N_5950);
or U12589 (N_12589,N_5994,N_5313);
xor U12590 (N_12590,N_8942,N_7658);
nand U12591 (N_12591,N_7007,N_6590);
xnor U12592 (N_12592,N_6212,N_5333);
xor U12593 (N_12593,N_7348,N_9628);
and U12594 (N_12594,N_8592,N_6172);
nand U12595 (N_12595,N_9560,N_8700);
xor U12596 (N_12596,N_5680,N_8123);
xnor U12597 (N_12597,N_9389,N_5932);
and U12598 (N_12598,N_8265,N_5849);
or U12599 (N_12599,N_7737,N_9873);
xnor U12600 (N_12600,N_6044,N_6716);
nor U12601 (N_12601,N_6823,N_8727);
and U12602 (N_12602,N_5265,N_7056);
or U12603 (N_12603,N_9543,N_8166);
nor U12604 (N_12604,N_6489,N_7862);
xnor U12605 (N_12605,N_5846,N_5009);
and U12606 (N_12606,N_6845,N_8331);
nand U12607 (N_12607,N_7108,N_6927);
xor U12608 (N_12608,N_5462,N_5188);
nand U12609 (N_12609,N_5327,N_9079);
and U12610 (N_12610,N_5166,N_8287);
nor U12611 (N_12611,N_5802,N_6788);
and U12612 (N_12612,N_8169,N_8697);
or U12613 (N_12613,N_6245,N_7698);
nand U12614 (N_12614,N_8364,N_9184);
nor U12615 (N_12615,N_8990,N_5635);
nor U12616 (N_12616,N_5545,N_6812);
nor U12617 (N_12617,N_8285,N_8709);
or U12618 (N_12618,N_5742,N_9098);
nor U12619 (N_12619,N_8100,N_7502);
nand U12620 (N_12620,N_7327,N_7394);
or U12621 (N_12621,N_9100,N_6499);
or U12622 (N_12622,N_8721,N_7084);
xor U12623 (N_12623,N_9036,N_9092);
and U12624 (N_12624,N_8581,N_7731);
or U12625 (N_12625,N_8499,N_8063);
or U12626 (N_12626,N_8790,N_9983);
nand U12627 (N_12627,N_9070,N_7283);
nor U12628 (N_12628,N_9242,N_7812);
nor U12629 (N_12629,N_8703,N_9160);
nand U12630 (N_12630,N_7462,N_7707);
or U12631 (N_12631,N_6441,N_7624);
nand U12632 (N_12632,N_6739,N_9753);
xor U12633 (N_12633,N_7715,N_5294);
or U12634 (N_12634,N_8897,N_8746);
or U12635 (N_12635,N_6034,N_8408);
and U12636 (N_12636,N_6296,N_5934);
and U12637 (N_12637,N_8464,N_8374);
nand U12638 (N_12638,N_5825,N_6404);
xnor U12639 (N_12639,N_9044,N_8771);
nor U12640 (N_12640,N_9720,N_7892);
and U12641 (N_12641,N_6025,N_6226);
nor U12642 (N_12642,N_8274,N_8090);
and U12643 (N_12643,N_7838,N_7431);
nand U12644 (N_12644,N_8802,N_6549);
xor U12645 (N_12645,N_9177,N_5871);
xor U12646 (N_12646,N_8984,N_8465);
and U12647 (N_12647,N_5712,N_9047);
nor U12648 (N_12648,N_6944,N_6582);
and U12649 (N_12649,N_7094,N_6952);
xor U12650 (N_12650,N_6998,N_5626);
xor U12651 (N_12651,N_5279,N_6207);
or U12652 (N_12652,N_6986,N_8827);
nand U12653 (N_12653,N_6037,N_9408);
xor U12654 (N_12654,N_6297,N_9320);
nand U12655 (N_12655,N_9360,N_7771);
and U12656 (N_12656,N_9305,N_8075);
nor U12657 (N_12657,N_8832,N_8336);
nand U12658 (N_12658,N_6390,N_9982);
or U12659 (N_12659,N_9621,N_9966);
or U12660 (N_12660,N_6320,N_6690);
nor U12661 (N_12661,N_6483,N_6196);
nor U12662 (N_12662,N_7139,N_7762);
nor U12663 (N_12663,N_6962,N_9702);
nor U12664 (N_12664,N_5392,N_5093);
and U12665 (N_12665,N_6398,N_9202);
nand U12666 (N_12666,N_8902,N_6961);
nand U12667 (N_12667,N_6916,N_8487);
xnor U12668 (N_12668,N_6493,N_5816);
and U12669 (N_12669,N_9597,N_5160);
nor U12670 (N_12670,N_8460,N_8597);
nand U12671 (N_12671,N_7056,N_9780);
and U12672 (N_12672,N_5640,N_6706);
or U12673 (N_12673,N_5581,N_8268);
or U12674 (N_12674,N_6661,N_9952);
nand U12675 (N_12675,N_6578,N_6326);
or U12676 (N_12676,N_9867,N_7503);
or U12677 (N_12677,N_9255,N_6384);
or U12678 (N_12678,N_9879,N_9356);
and U12679 (N_12679,N_8306,N_7756);
and U12680 (N_12680,N_6083,N_8912);
and U12681 (N_12681,N_5109,N_7392);
or U12682 (N_12682,N_8068,N_6699);
nand U12683 (N_12683,N_7322,N_9775);
nand U12684 (N_12684,N_8851,N_8051);
and U12685 (N_12685,N_6858,N_5792);
or U12686 (N_12686,N_9688,N_8815);
nand U12687 (N_12687,N_7087,N_7074);
nor U12688 (N_12688,N_5096,N_8191);
nand U12689 (N_12689,N_5672,N_7390);
xor U12690 (N_12690,N_7927,N_9614);
xor U12691 (N_12691,N_6503,N_8569);
nand U12692 (N_12692,N_8472,N_9576);
nand U12693 (N_12693,N_8903,N_8492);
xnor U12694 (N_12694,N_6031,N_7923);
nor U12695 (N_12695,N_8997,N_6603);
and U12696 (N_12696,N_9484,N_9997);
nor U12697 (N_12697,N_9481,N_8592);
and U12698 (N_12698,N_8198,N_7033);
and U12699 (N_12699,N_6574,N_7765);
xor U12700 (N_12700,N_6189,N_6358);
nand U12701 (N_12701,N_7200,N_6459);
nor U12702 (N_12702,N_5780,N_5249);
nand U12703 (N_12703,N_7702,N_9225);
xnor U12704 (N_12704,N_5332,N_8600);
and U12705 (N_12705,N_9261,N_8211);
nor U12706 (N_12706,N_5540,N_9759);
nand U12707 (N_12707,N_5086,N_8293);
and U12708 (N_12708,N_9220,N_7489);
and U12709 (N_12709,N_9744,N_5913);
xor U12710 (N_12710,N_5180,N_9080);
and U12711 (N_12711,N_7756,N_6056);
nor U12712 (N_12712,N_9051,N_5800);
and U12713 (N_12713,N_9015,N_5051);
xnor U12714 (N_12714,N_8556,N_9101);
xor U12715 (N_12715,N_5670,N_9504);
nand U12716 (N_12716,N_7385,N_8874);
and U12717 (N_12717,N_5845,N_6987);
and U12718 (N_12718,N_8657,N_6954);
xor U12719 (N_12719,N_6148,N_9816);
and U12720 (N_12720,N_5721,N_9630);
or U12721 (N_12721,N_5637,N_6184);
xnor U12722 (N_12722,N_8437,N_5812);
nand U12723 (N_12723,N_7701,N_7493);
nand U12724 (N_12724,N_6494,N_8409);
xnor U12725 (N_12725,N_9705,N_5396);
nand U12726 (N_12726,N_5258,N_5387);
and U12727 (N_12727,N_5468,N_9176);
and U12728 (N_12728,N_7757,N_6795);
xnor U12729 (N_12729,N_9737,N_8028);
and U12730 (N_12730,N_6465,N_8972);
and U12731 (N_12731,N_7733,N_6849);
nand U12732 (N_12732,N_9641,N_9823);
nand U12733 (N_12733,N_9045,N_8310);
nor U12734 (N_12734,N_9261,N_8102);
nor U12735 (N_12735,N_6787,N_9619);
nor U12736 (N_12736,N_5965,N_8733);
xor U12737 (N_12737,N_7953,N_6289);
nor U12738 (N_12738,N_7605,N_5692);
or U12739 (N_12739,N_9500,N_7103);
nand U12740 (N_12740,N_8911,N_6318);
nor U12741 (N_12741,N_8521,N_8499);
nand U12742 (N_12742,N_6954,N_5918);
and U12743 (N_12743,N_7524,N_7353);
nand U12744 (N_12744,N_9969,N_5816);
or U12745 (N_12745,N_8263,N_7032);
xnor U12746 (N_12746,N_6036,N_7334);
and U12747 (N_12747,N_9798,N_8411);
nand U12748 (N_12748,N_9917,N_6658);
xor U12749 (N_12749,N_9048,N_8285);
or U12750 (N_12750,N_5489,N_9019);
nand U12751 (N_12751,N_6008,N_5137);
xnor U12752 (N_12752,N_8898,N_9137);
xor U12753 (N_12753,N_5579,N_6493);
or U12754 (N_12754,N_7379,N_5135);
nor U12755 (N_12755,N_7547,N_9932);
nand U12756 (N_12756,N_9267,N_7571);
or U12757 (N_12757,N_6355,N_6810);
nand U12758 (N_12758,N_6851,N_6546);
xor U12759 (N_12759,N_9095,N_9172);
xnor U12760 (N_12760,N_9158,N_7061);
nor U12761 (N_12761,N_5149,N_5586);
or U12762 (N_12762,N_9626,N_9835);
nand U12763 (N_12763,N_9015,N_9363);
nand U12764 (N_12764,N_8502,N_8908);
nor U12765 (N_12765,N_6632,N_5697);
nand U12766 (N_12766,N_5324,N_7375);
nand U12767 (N_12767,N_9383,N_8704);
and U12768 (N_12768,N_5619,N_5890);
or U12769 (N_12769,N_6819,N_9777);
and U12770 (N_12770,N_9191,N_6521);
and U12771 (N_12771,N_7830,N_6840);
nor U12772 (N_12772,N_5647,N_6415);
xnor U12773 (N_12773,N_9445,N_6411);
and U12774 (N_12774,N_6128,N_6318);
or U12775 (N_12775,N_7153,N_8187);
nor U12776 (N_12776,N_5990,N_6118);
nor U12777 (N_12777,N_5027,N_8148);
and U12778 (N_12778,N_6411,N_5500);
and U12779 (N_12779,N_5148,N_6911);
or U12780 (N_12780,N_6908,N_9526);
nor U12781 (N_12781,N_6309,N_7578);
xnor U12782 (N_12782,N_7870,N_5967);
nor U12783 (N_12783,N_7749,N_6217);
xnor U12784 (N_12784,N_8441,N_9906);
nor U12785 (N_12785,N_8529,N_7836);
nor U12786 (N_12786,N_6120,N_7197);
and U12787 (N_12787,N_7902,N_7684);
and U12788 (N_12788,N_7620,N_7485);
xnor U12789 (N_12789,N_7285,N_8392);
xnor U12790 (N_12790,N_7430,N_5099);
nand U12791 (N_12791,N_8854,N_8104);
and U12792 (N_12792,N_6939,N_7313);
and U12793 (N_12793,N_6484,N_8874);
and U12794 (N_12794,N_8334,N_5447);
nand U12795 (N_12795,N_5614,N_8703);
nor U12796 (N_12796,N_8146,N_7255);
nor U12797 (N_12797,N_8140,N_7101);
and U12798 (N_12798,N_6440,N_5333);
and U12799 (N_12799,N_7371,N_9585);
nand U12800 (N_12800,N_7036,N_6103);
and U12801 (N_12801,N_5216,N_7330);
nand U12802 (N_12802,N_9574,N_8178);
xnor U12803 (N_12803,N_5459,N_9866);
nand U12804 (N_12804,N_8843,N_7374);
xnor U12805 (N_12805,N_5002,N_6690);
or U12806 (N_12806,N_6509,N_5842);
nand U12807 (N_12807,N_8216,N_5319);
nor U12808 (N_12808,N_7998,N_6806);
nor U12809 (N_12809,N_6241,N_9990);
xnor U12810 (N_12810,N_8870,N_5209);
nor U12811 (N_12811,N_9783,N_8195);
and U12812 (N_12812,N_7412,N_9873);
and U12813 (N_12813,N_9090,N_7008);
nand U12814 (N_12814,N_7631,N_7206);
xnor U12815 (N_12815,N_5274,N_5971);
nor U12816 (N_12816,N_5846,N_5489);
nor U12817 (N_12817,N_8574,N_8165);
or U12818 (N_12818,N_6172,N_6607);
or U12819 (N_12819,N_7014,N_9513);
xnor U12820 (N_12820,N_5440,N_9388);
xnor U12821 (N_12821,N_7225,N_5406);
xor U12822 (N_12822,N_7595,N_7482);
or U12823 (N_12823,N_6389,N_7678);
and U12824 (N_12824,N_5437,N_8651);
nand U12825 (N_12825,N_9094,N_8794);
nor U12826 (N_12826,N_8579,N_9180);
and U12827 (N_12827,N_6529,N_8914);
or U12828 (N_12828,N_6605,N_5158);
or U12829 (N_12829,N_9349,N_7884);
nor U12830 (N_12830,N_8258,N_9505);
nor U12831 (N_12831,N_8106,N_6841);
nand U12832 (N_12832,N_8338,N_7499);
nor U12833 (N_12833,N_6421,N_5240);
and U12834 (N_12834,N_5864,N_6869);
nor U12835 (N_12835,N_6467,N_5644);
or U12836 (N_12836,N_5988,N_6935);
nor U12837 (N_12837,N_6344,N_9324);
and U12838 (N_12838,N_9151,N_7519);
nand U12839 (N_12839,N_6818,N_6458);
and U12840 (N_12840,N_9795,N_7141);
and U12841 (N_12841,N_6570,N_9739);
and U12842 (N_12842,N_9769,N_7093);
and U12843 (N_12843,N_6063,N_9916);
nand U12844 (N_12844,N_8530,N_7202);
nor U12845 (N_12845,N_9673,N_5040);
and U12846 (N_12846,N_9341,N_9037);
xnor U12847 (N_12847,N_7002,N_6462);
or U12848 (N_12848,N_5096,N_6413);
nor U12849 (N_12849,N_7399,N_7680);
nand U12850 (N_12850,N_9021,N_8891);
xnor U12851 (N_12851,N_5434,N_9242);
nand U12852 (N_12852,N_7252,N_8596);
nor U12853 (N_12853,N_5358,N_7384);
nor U12854 (N_12854,N_9050,N_9765);
nor U12855 (N_12855,N_8428,N_6168);
xor U12856 (N_12856,N_8270,N_9461);
nand U12857 (N_12857,N_5126,N_5617);
xor U12858 (N_12858,N_9325,N_8989);
nor U12859 (N_12859,N_5344,N_8362);
or U12860 (N_12860,N_7387,N_9525);
nand U12861 (N_12861,N_6329,N_5977);
xor U12862 (N_12862,N_7826,N_7599);
and U12863 (N_12863,N_7122,N_8607);
or U12864 (N_12864,N_6891,N_8859);
or U12865 (N_12865,N_9813,N_6961);
nor U12866 (N_12866,N_9451,N_9704);
or U12867 (N_12867,N_5817,N_9018);
xnor U12868 (N_12868,N_5066,N_5033);
and U12869 (N_12869,N_7475,N_5770);
nand U12870 (N_12870,N_5478,N_8981);
nor U12871 (N_12871,N_5875,N_7995);
or U12872 (N_12872,N_8622,N_7110);
or U12873 (N_12873,N_7553,N_7460);
and U12874 (N_12874,N_5921,N_8530);
or U12875 (N_12875,N_6746,N_6533);
xor U12876 (N_12876,N_9143,N_5332);
and U12877 (N_12877,N_7747,N_8881);
nor U12878 (N_12878,N_5395,N_7450);
or U12879 (N_12879,N_9964,N_6652);
nand U12880 (N_12880,N_7549,N_6285);
nor U12881 (N_12881,N_9333,N_5879);
and U12882 (N_12882,N_9662,N_7830);
and U12883 (N_12883,N_8779,N_6651);
nand U12884 (N_12884,N_6117,N_9183);
nor U12885 (N_12885,N_9114,N_7218);
nand U12886 (N_12886,N_6027,N_6407);
and U12887 (N_12887,N_6968,N_6938);
xnor U12888 (N_12888,N_6576,N_7178);
nor U12889 (N_12889,N_9261,N_9973);
nor U12890 (N_12890,N_5583,N_8162);
nand U12891 (N_12891,N_5038,N_5313);
nand U12892 (N_12892,N_7335,N_7891);
or U12893 (N_12893,N_6558,N_5879);
nand U12894 (N_12894,N_7451,N_9638);
or U12895 (N_12895,N_5799,N_9342);
or U12896 (N_12896,N_5894,N_5149);
or U12897 (N_12897,N_8711,N_7416);
nor U12898 (N_12898,N_9356,N_9402);
and U12899 (N_12899,N_5343,N_9990);
nand U12900 (N_12900,N_7851,N_7464);
and U12901 (N_12901,N_6077,N_7354);
nor U12902 (N_12902,N_9740,N_5281);
xor U12903 (N_12903,N_8395,N_5494);
xor U12904 (N_12904,N_6395,N_8083);
and U12905 (N_12905,N_9469,N_9581);
or U12906 (N_12906,N_7601,N_6380);
and U12907 (N_12907,N_6058,N_8963);
nand U12908 (N_12908,N_5560,N_9912);
xnor U12909 (N_12909,N_9623,N_9859);
and U12910 (N_12910,N_5040,N_8179);
xnor U12911 (N_12911,N_5379,N_6827);
nor U12912 (N_12912,N_8400,N_9628);
xnor U12913 (N_12913,N_7740,N_7411);
xor U12914 (N_12914,N_5810,N_7713);
or U12915 (N_12915,N_9974,N_6638);
or U12916 (N_12916,N_7141,N_9546);
nor U12917 (N_12917,N_9786,N_8742);
or U12918 (N_12918,N_5633,N_6044);
or U12919 (N_12919,N_9961,N_7945);
or U12920 (N_12920,N_6854,N_9083);
and U12921 (N_12921,N_6835,N_5111);
or U12922 (N_12922,N_9236,N_7427);
nand U12923 (N_12923,N_6887,N_9738);
and U12924 (N_12924,N_6291,N_8375);
or U12925 (N_12925,N_9996,N_8642);
xor U12926 (N_12926,N_6395,N_6002);
and U12927 (N_12927,N_8250,N_7001);
xnor U12928 (N_12928,N_5363,N_7806);
or U12929 (N_12929,N_8797,N_7722);
xor U12930 (N_12930,N_7886,N_7302);
and U12931 (N_12931,N_8674,N_9299);
and U12932 (N_12932,N_7617,N_9163);
and U12933 (N_12933,N_9272,N_6100);
nand U12934 (N_12934,N_5157,N_5306);
or U12935 (N_12935,N_6602,N_8447);
and U12936 (N_12936,N_5241,N_9112);
or U12937 (N_12937,N_7042,N_6498);
or U12938 (N_12938,N_7818,N_9547);
or U12939 (N_12939,N_7514,N_8445);
or U12940 (N_12940,N_5919,N_6346);
or U12941 (N_12941,N_6209,N_5287);
nor U12942 (N_12942,N_8663,N_5381);
or U12943 (N_12943,N_7905,N_5566);
xnor U12944 (N_12944,N_9514,N_6671);
or U12945 (N_12945,N_6478,N_7826);
or U12946 (N_12946,N_5341,N_7672);
or U12947 (N_12947,N_7612,N_8766);
or U12948 (N_12948,N_6647,N_9708);
or U12949 (N_12949,N_8371,N_6897);
nor U12950 (N_12950,N_9098,N_7824);
and U12951 (N_12951,N_6784,N_7119);
and U12952 (N_12952,N_6952,N_9506);
and U12953 (N_12953,N_8975,N_6593);
and U12954 (N_12954,N_7267,N_6747);
nor U12955 (N_12955,N_7354,N_7169);
nor U12956 (N_12956,N_7341,N_5661);
and U12957 (N_12957,N_9811,N_5381);
xor U12958 (N_12958,N_5380,N_9065);
xor U12959 (N_12959,N_9460,N_8904);
nor U12960 (N_12960,N_8882,N_9656);
and U12961 (N_12961,N_5270,N_5981);
nand U12962 (N_12962,N_5570,N_5785);
nor U12963 (N_12963,N_8039,N_7217);
nor U12964 (N_12964,N_8332,N_7993);
nand U12965 (N_12965,N_8143,N_7988);
nor U12966 (N_12966,N_6635,N_9602);
nand U12967 (N_12967,N_8237,N_6359);
xnor U12968 (N_12968,N_9304,N_9588);
nand U12969 (N_12969,N_6758,N_7413);
nor U12970 (N_12970,N_7681,N_5098);
nand U12971 (N_12971,N_7739,N_6515);
nor U12972 (N_12972,N_5842,N_9254);
nor U12973 (N_12973,N_6237,N_7845);
or U12974 (N_12974,N_7655,N_6668);
nor U12975 (N_12975,N_7901,N_9890);
or U12976 (N_12976,N_7353,N_7553);
or U12977 (N_12977,N_9018,N_8856);
nor U12978 (N_12978,N_5037,N_5497);
nand U12979 (N_12979,N_5416,N_6840);
nor U12980 (N_12980,N_6484,N_6600);
and U12981 (N_12981,N_6785,N_9377);
and U12982 (N_12982,N_6144,N_9527);
nand U12983 (N_12983,N_9832,N_8154);
nor U12984 (N_12984,N_6778,N_9011);
xnor U12985 (N_12985,N_8995,N_8191);
xnor U12986 (N_12986,N_6107,N_9865);
and U12987 (N_12987,N_6010,N_9362);
xor U12988 (N_12988,N_6918,N_7073);
and U12989 (N_12989,N_8643,N_9420);
and U12990 (N_12990,N_5473,N_6021);
or U12991 (N_12991,N_8108,N_6621);
xor U12992 (N_12992,N_5722,N_9477);
xnor U12993 (N_12993,N_9479,N_6921);
or U12994 (N_12994,N_5676,N_9596);
xnor U12995 (N_12995,N_6656,N_5120);
or U12996 (N_12996,N_8154,N_8138);
or U12997 (N_12997,N_8116,N_5138);
nor U12998 (N_12998,N_7931,N_9115);
nor U12999 (N_12999,N_6530,N_6607);
nand U13000 (N_13000,N_7805,N_5852);
nand U13001 (N_13001,N_8959,N_8967);
xor U13002 (N_13002,N_5294,N_6904);
nor U13003 (N_13003,N_7205,N_7680);
nor U13004 (N_13004,N_5675,N_5768);
xor U13005 (N_13005,N_6724,N_8728);
nor U13006 (N_13006,N_9995,N_7678);
and U13007 (N_13007,N_5092,N_8405);
and U13008 (N_13008,N_7533,N_6380);
xor U13009 (N_13009,N_5077,N_6927);
and U13010 (N_13010,N_9544,N_5269);
nor U13011 (N_13011,N_6853,N_9887);
xnor U13012 (N_13012,N_7748,N_6129);
xor U13013 (N_13013,N_7922,N_6747);
xnor U13014 (N_13014,N_8963,N_9753);
nor U13015 (N_13015,N_7654,N_7025);
nor U13016 (N_13016,N_9035,N_8724);
nand U13017 (N_13017,N_5723,N_8013);
nor U13018 (N_13018,N_6824,N_9033);
or U13019 (N_13019,N_5589,N_9266);
and U13020 (N_13020,N_7294,N_9131);
xor U13021 (N_13021,N_9089,N_6842);
or U13022 (N_13022,N_5007,N_9397);
nor U13023 (N_13023,N_9149,N_7105);
and U13024 (N_13024,N_5021,N_6150);
or U13025 (N_13025,N_7588,N_6876);
nand U13026 (N_13026,N_7088,N_5397);
xnor U13027 (N_13027,N_6169,N_7405);
nor U13028 (N_13028,N_5540,N_8704);
and U13029 (N_13029,N_9523,N_5616);
nand U13030 (N_13030,N_7561,N_5020);
nand U13031 (N_13031,N_9002,N_9522);
nor U13032 (N_13032,N_8493,N_6417);
xnor U13033 (N_13033,N_5519,N_6617);
or U13034 (N_13034,N_7888,N_9090);
and U13035 (N_13035,N_8988,N_7763);
or U13036 (N_13036,N_5652,N_5074);
nand U13037 (N_13037,N_7448,N_6772);
and U13038 (N_13038,N_6536,N_7989);
and U13039 (N_13039,N_5950,N_5227);
nand U13040 (N_13040,N_9583,N_6858);
xnor U13041 (N_13041,N_7014,N_9041);
or U13042 (N_13042,N_8147,N_8004);
nand U13043 (N_13043,N_7550,N_9697);
nor U13044 (N_13044,N_9033,N_9191);
or U13045 (N_13045,N_9348,N_5629);
nand U13046 (N_13046,N_8695,N_7146);
nor U13047 (N_13047,N_6083,N_7763);
nand U13048 (N_13048,N_5722,N_6882);
and U13049 (N_13049,N_5835,N_6050);
nand U13050 (N_13050,N_6774,N_8275);
nand U13051 (N_13051,N_5987,N_9745);
nand U13052 (N_13052,N_7792,N_9775);
nor U13053 (N_13053,N_7594,N_6090);
nor U13054 (N_13054,N_6488,N_8601);
and U13055 (N_13055,N_9107,N_8905);
nand U13056 (N_13056,N_6538,N_5639);
and U13057 (N_13057,N_5752,N_7413);
xor U13058 (N_13058,N_8351,N_8326);
nor U13059 (N_13059,N_6839,N_9192);
or U13060 (N_13060,N_8791,N_6209);
xnor U13061 (N_13061,N_8739,N_8618);
and U13062 (N_13062,N_7763,N_9430);
nor U13063 (N_13063,N_7724,N_6010);
xnor U13064 (N_13064,N_9966,N_6308);
and U13065 (N_13065,N_5903,N_6469);
nand U13066 (N_13066,N_5968,N_8042);
nand U13067 (N_13067,N_7101,N_9929);
and U13068 (N_13068,N_5546,N_9418);
or U13069 (N_13069,N_5945,N_5151);
or U13070 (N_13070,N_6077,N_8382);
and U13071 (N_13071,N_9264,N_9602);
nand U13072 (N_13072,N_6756,N_7515);
nand U13073 (N_13073,N_5911,N_5094);
xnor U13074 (N_13074,N_5030,N_6134);
or U13075 (N_13075,N_8966,N_6154);
and U13076 (N_13076,N_9995,N_9378);
and U13077 (N_13077,N_5595,N_9579);
and U13078 (N_13078,N_8687,N_7561);
and U13079 (N_13079,N_8766,N_5653);
nand U13080 (N_13080,N_5112,N_9625);
nand U13081 (N_13081,N_7939,N_6763);
xor U13082 (N_13082,N_5203,N_9199);
or U13083 (N_13083,N_7929,N_9092);
nand U13084 (N_13084,N_6439,N_9404);
or U13085 (N_13085,N_9104,N_9577);
or U13086 (N_13086,N_6379,N_7034);
nor U13087 (N_13087,N_5746,N_5747);
xnor U13088 (N_13088,N_5888,N_6283);
nand U13089 (N_13089,N_9919,N_5121);
and U13090 (N_13090,N_6264,N_5759);
nor U13091 (N_13091,N_9614,N_8729);
and U13092 (N_13092,N_6184,N_6490);
and U13093 (N_13093,N_7983,N_6037);
and U13094 (N_13094,N_5575,N_7139);
nand U13095 (N_13095,N_7613,N_6876);
nor U13096 (N_13096,N_7585,N_6497);
nor U13097 (N_13097,N_9958,N_5136);
nor U13098 (N_13098,N_6227,N_9368);
and U13099 (N_13099,N_7665,N_9697);
nand U13100 (N_13100,N_6154,N_9726);
nand U13101 (N_13101,N_6390,N_6859);
nand U13102 (N_13102,N_8593,N_9441);
xnor U13103 (N_13103,N_8471,N_6642);
and U13104 (N_13104,N_7016,N_6876);
or U13105 (N_13105,N_6943,N_7584);
nor U13106 (N_13106,N_8874,N_6578);
nand U13107 (N_13107,N_7073,N_8247);
and U13108 (N_13108,N_6298,N_9021);
nand U13109 (N_13109,N_9382,N_5367);
nor U13110 (N_13110,N_8170,N_6087);
nor U13111 (N_13111,N_9254,N_6424);
xor U13112 (N_13112,N_6455,N_7752);
xor U13113 (N_13113,N_9999,N_7310);
or U13114 (N_13114,N_7622,N_7101);
nor U13115 (N_13115,N_7187,N_7103);
nor U13116 (N_13116,N_6977,N_9195);
and U13117 (N_13117,N_5882,N_7043);
xor U13118 (N_13118,N_9687,N_5963);
nand U13119 (N_13119,N_7164,N_5371);
nand U13120 (N_13120,N_9226,N_5113);
xor U13121 (N_13121,N_7371,N_8143);
and U13122 (N_13122,N_5788,N_5207);
nand U13123 (N_13123,N_6240,N_7830);
xor U13124 (N_13124,N_6424,N_7372);
xnor U13125 (N_13125,N_5881,N_5289);
or U13126 (N_13126,N_9420,N_7176);
nor U13127 (N_13127,N_7471,N_6129);
and U13128 (N_13128,N_9850,N_9132);
xnor U13129 (N_13129,N_5872,N_6785);
xor U13130 (N_13130,N_8450,N_7036);
or U13131 (N_13131,N_6958,N_8010);
nor U13132 (N_13132,N_8600,N_8446);
or U13133 (N_13133,N_7706,N_9246);
nor U13134 (N_13134,N_9360,N_6549);
xor U13135 (N_13135,N_6864,N_9895);
or U13136 (N_13136,N_9021,N_7663);
and U13137 (N_13137,N_8612,N_8754);
and U13138 (N_13138,N_6746,N_9225);
nand U13139 (N_13139,N_9151,N_8787);
or U13140 (N_13140,N_6632,N_8675);
or U13141 (N_13141,N_5793,N_6491);
and U13142 (N_13142,N_5100,N_9122);
and U13143 (N_13143,N_7411,N_5363);
and U13144 (N_13144,N_7481,N_5528);
xor U13145 (N_13145,N_9960,N_5741);
or U13146 (N_13146,N_6179,N_8991);
and U13147 (N_13147,N_7970,N_5776);
nor U13148 (N_13148,N_5433,N_9877);
nor U13149 (N_13149,N_9420,N_8389);
and U13150 (N_13150,N_9523,N_7739);
xor U13151 (N_13151,N_7845,N_5132);
nand U13152 (N_13152,N_5955,N_7508);
xnor U13153 (N_13153,N_7912,N_8978);
or U13154 (N_13154,N_5337,N_5435);
nand U13155 (N_13155,N_8789,N_6693);
and U13156 (N_13156,N_6197,N_5130);
or U13157 (N_13157,N_8982,N_7242);
nor U13158 (N_13158,N_6743,N_6318);
and U13159 (N_13159,N_9772,N_9347);
or U13160 (N_13160,N_5872,N_8235);
or U13161 (N_13161,N_5957,N_8956);
or U13162 (N_13162,N_7038,N_8241);
nor U13163 (N_13163,N_6382,N_5493);
nand U13164 (N_13164,N_7128,N_7635);
xor U13165 (N_13165,N_8102,N_8804);
or U13166 (N_13166,N_5269,N_7408);
or U13167 (N_13167,N_5291,N_6211);
nand U13168 (N_13168,N_9751,N_6288);
nor U13169 (N_13169,N_8347,N_7161);
nand U13170 (N_13170,N_5481,N_5340);
xnor U13171 (N_13171,N_7969,N_5465);
or U13172 (N_13172,N_7077,N_6117);
and U13173 (N_13173,N_6827,N_5662);
xnor U13174 (N_13174,N_7339,N_8185);
nand U13175 (N_13175,N_8863,N_9447);
and U13176 (N_13176,N_5768,N_8243);
nor U13177 (N_13177,N_6267,N_7273);
xnor U13178 (N_13178,N_9183,N_7374);
nand U13179 (N_13179,N_6744,N_7412);
nor U13180 (N_13180,N_7939,N_5462);
nor U13181 (N_13181,N_6880,N_8130);
nor U13182 (N_13182,N_7645,N_9122);
nand U13183 (N_13183,N_5396,N_9310);
nor U13184 (N_13184,N_5826,N_9641);
and U13185 (N_13185,N_5490,N_9202);
nor U13186 (N_13186,N_7233,N_8278);
and U13187 (N_13187,N_7194,N_8177);
and U13188 (N_13188,N_7421,N_9451);
and U13189 (N_13189,N_9590,N_5146);
xnor U13190 (N_13190,N_8204,N_8417);
or U13191 (N_13191,N_9261,N_5517);
nand U13192 (N_13192,N_7469,N_5208);
nand U13193 (N_13193,N_7903,N_8679);
or U13194 (N_13194,N_7505,N_5049);
xnor U13195 (N_13195,N_6540,N_6609);
or U13196 (N_13196,N_9937,N_5124);
and U13197 (N_13197,N_5300,N_8609);
and U13198 (N_13198,N_9070,N_9926);
xor U13199 (N_13199,N_7999,N_6219);
nor U13200 (N_13200,N_8981,N_5684);
or U13201 (N_13201,N_8886,N_9472);
or U13202 (N_13202,N_7381,N_6572);
or U13203 (N_13203,N_7192,N_5292);
xor U13204 (N_13204,N_7713,N_5984);
xor U13205 (N_13205,N_6276,N_9487);
or U13206 (N_13206,N_7186,N_8340);
and U13207 (N_13207,N_9284,N_7909);
nor U13208 (N_13208,N_6136,N_7039);
or U13209 (N_13209,N_5937,N_8457);
nand U13210 (N_13210,N_6788,N_7739);
and U13211 (N_13211,N_5401,N_6008);
and U13212 (N_13212,N_5779,N_6804);
or U13213 (N_13213,N_9766,N_8745);
or U13214 (N_13214,N_6041,N_9116);
or U13215 (N_13215,N_8186,N_9053);
or U13216 (N_13216,N_9246,N_5312);
and U13217 (N_13217,N_9357,N_7664);
nand U13218 (N_13218,N_5353,N_6868);
nor U13219 (N_13219,N_8282,N_8434);
or U13220 (N_13220,N_6232,N_6255);
and U13221 (N_13221,N_7835,N_5864);
nor U13222 (N_13222,N_5783,N_6666);
xnor U13223 (N_13223,N_6339,N_6149);
and U13224 (N_13224,N_6317,N_9451);
xnor U13225 (N_13225,N_7746,N_7538);
or U13226 (N_13226,N_8455,N_6051);
nor U13227 (N_13227,N_5814,N_7732);
nand U13228 (N_13228,N_5591,N_6884);
nand U13229 (N_13229,N_6479,N_8112);
xnor U13230 (N_13230,N_5697,N_9153);
and U13231 (N_13231,N_7112,N_6517);
or U13232 (N_13232,N_7369,N_9186);
nand U13233 (N_13233,N_5226,N_5830);
xor U13234 (N_13234,N_6513,N_7770);
nand U13235 (N_13235,N_9431,N_8653);
nor U13236 (N_13236,N_5018,N_8080);
and U13237 (N_13237,N_8050,N_9182);
xor U13238 (N_13238,N_7330,N_8973);
nor U13239 (N_13239,N_5156,N_5555);
or U13240 (N_13240,N_8219,N_9095);
nand U13241 (N_13241,N_8140,N_8166);
xor U13242 (N_13242,N_7598,N_8118);
or U13243 (N_13243,N_5746,N_8801);
nor U13244 (N_13244,N_5643,N_9544);
or U13245 (N_13245,N_8722,N_6464);
nand U13246 (N_13246,N_7264,N_7116);
and U13247 (N_13247,N_6047,N_8372);
xnor U13248 (N_13248,N_9192,N_9295);
or U13249 (N_13249,N_5915,N_6211);
nand U13250 (N_13250,N_6597,N_6781);
nor U13251 (N_13251,N_8797,N_6286);
xor U13252 (N_13252,N_9379,N_6603);
xnor U13253 (N_13253,N_7165,N_5320);
or U13254 (N_13254,N_8819,N_8752);
nor U13255 (N_13255,N_7684,N_5603);
nand U13256 (N_13256,N_7277,N_5432);
nand U13257 (N_13257,N_9311,N_6302);
and U13258 (N_13258,N_7221,N_5332);
xnor U13259 (N_13259,N_5055,N_7251);
nand U13260 (N_13260,N_9693,N_9408);
and U13261 (N_13261,N_6512,N_7928);
nand U13262 (N_13262,N_8944,N_7203);
nor U13263 (N_13263,N_6093,N_6444);
xnor U13264 (N_13264,N_8624,N_9365);
and U13265 (N_13265,N_6577,N_8275);
xnor U13266 (N_13266,N_5776,N_7814);
and U13267 (N_13267,N_7285,N_6571);
or U13268 (N_13268,N_9782,N_6376);
and U13269 (N_13269,N_9903,N_8916);
nand U13270 (N_13270,N_9184,N_5352);
xor U13271 (N_13271,N_9268,N_6240);
nor U13272 (N_13272,N_7078,N_5830);
or U13273 (N_13273,N_7228,N_5418);
nor U13274 (N_13274,N_5549,N_5285);
and U13275 (N_13275,N_5452,N_5990);
nand U13276 (N_13276,N_9922,N_6967);
or U13277 (N_13277,N_5980,N_6006);
nand U13278 (N_13278,N_8283,N_7087);
and U13279 (N_13279,N_8016,N_7478);
or U13280 (N_13280,N_7262,N_5342);
or U13281 (N_13281,N_9350,N_8395);
or U13282 (N_13282,N_6751,N_6046);
nand U13283 (N_13283,N_8076,N_7399);
nand U13284 (N_13284,N_9453,N_7510);
and U13285 (N_13285,N_7092,N_5643);
nand U13286 (N_13286,N_6921,N_5973);
nand U13287 (N_13287,N_8448,N_9321);
nand U13288 (N_13288,N_7141,N_7380);
or U13289 (N_13289,N_7572,N_7348);
nand U13290 (N_13290,N_6251,N_7307);
nand U13291 (N_13291,N_6895,N_7066);
nor U13292 (N_13292,N_7377,N_5546);
nor U13293 (N_13293,N_8710,N_8415);
and U13294 (N_13294,N_6735,N_8071);
xor U13295 (N_13295,N_5840,N_6278);
nor U13296 (N_13296,N_5397,N_7455);
nand U13297 (N_13297,N_8490,N_9887);
nand U13298 (N_13298,N_9959,N_9789);
and U13299 (N_13299,N_8747,N_5738);
xnor U13300 (N_13300,N_9427,N_9853);
nor U13301 (N_13301,N_8435,N_5088);
xor U13302 (N_13302,N_6911,N_9806);
and U13303 (N_13303,N_8125,N_8407);
xnor U13304 (N_13304,N_6949,N_9452);
or U13305 (N_13305,N_5496,N_7810);
xor U13306 (N_13306,N_8937,N_9582);
or U13307 (N_13307,N_8834,N_7316);
and U13308 (N_13308,N_5773,N_5668);
and U13309 (N_13309,N_7684,N_7596);
or U13310 (N_13310,N_8249,N_5811);
and U13311 (N_13311,N_8475,N_8612);
xnor U13312 (N_13312,N_8516,N_6642);
nand U13313 (N_13313,N_6038,N_8289);
nor U13314 (N_13314,N_5858,N_5584);
or U13315 (N_13315,N_9370,N_8658);
nor U13316 (N_13316,N_6223,N_5535);
nor U13317 (N_13317,N_6322,N_5348);
or U13318 (N_13318,N_8214,N_6150);
nor U13319 (N_13319,N_5688,N_8348);
or U13320 (N_13320,N_6558,N_8428);
xnor U13321 (N_13321,N_7360,N_6161);
nand U13322 (N_13322,N_6979,N_8993);
and U13323 (N_13323,N_9180,N_8901);
xnor U13324 (N_13324,N_7668,N_7190);
and U13325 (N_13325,N_6653,N_9463);
and U13326 (N_13326,N_6318,N_9464);
xnor U13327 (N_13327,N_5953,N_9288);
nor U13328 (N_13328,N_9221,N_9920);
xnor U13329 (N_13329,N_6146,N_5447);
nor U13330 (N_13330,N_5413,N_5270);
xnor U13331 (N_13331,N_9501,N_6404);
xor U13332 (N_13332,N_8244,N_7390);
xnor U13333 (N_13333,N_8749,N_6890);
nand U13334 (N_13334,N_9038,N_8536);
xnor U13335 (N_13335,N_9357,N_6471);
or U13336 (N_13336,N_9473,N_7838);
xnor U13337 (N_13337,N_6564,N_9291);
or U13338 (N_13338,N_9337,N_5573);
xnor U13339 (N_13339,N_6924,N_8272);
nor U13340 (N_13340,N_7476,N_6245);
nand U13341 (N_13341,N_8812,N_9215);
or U13342 (N_13342,N_6615,N_6928);
or U13343 (N_13343,N_7459,N_5165);
and U13344 (N_13344,N_8904,N_8913);
nor U13345 (N_13345,N_6742,N_8912);
nand U13346 (N_13346,N_7938,N_9514);
or U13347 (N_13347,N_5749,N_5730);
nor U13348 (N_13348,N_7079,N_5319);
nor U13349 (N_13349,N_6632,N_6007);
and U13350 (N_13350,N_9210,N_7179);
or U13351 (N_13351,N_7627,N_9475);
xnor U13352 (N_13352,N_8902,N_9886);
nor U13353 (N_13353,N_9008,N_7440);
nor U13354 (N_13354,N_5951,N_9421);
nand U13355 (N_13355,N_6802,N_9793);
nor U13356 (N_13356,N_9930,N_7028);
nor U13357 (N_13357,N_5011,N_7319);
nand U13358 (N_13358,N_7427,N_7108);
nand U13359 (N_13359,N_7200,N_8874);
xnor U13360 (N_13360,N_6676,N_5643);
nor U13361 (N_13361,N_8915,N_8213);
nand U13362 (N_13362,N_5866,N_7680);
nor U13363 (N_13363,N_5682,N_5598);
or U13364 (N_13364,N_5353,N_9870);
and U13365 (N_13365,N_9513,N_9276);
nor U13366 (N_13366,N_6955,N_9942);
nand U13367 (N_13367,N_8048,N_6288);
and U13368 (N_13368,N_8954,N_5675);
or U13369 (N_13369,N_5124,N_9182);
and U13370 (N_13370,N_6819,N_8061);
and U13371 (N_13371,N_9095,N_6376);
xnor U13372 (N_13372,N_6945,N_7520);
and U13373 (N_13373,N_8510,N_7658);
nor U13374 (N_13374,N_8732,N_6801);
nor U13375 (N_13375,N_9389,N_8626);
xnor U13376 (N_13376,N_7853,N_7489);
nor U13377 (N_13377,N_8576,N_5692);
and U13378 (N_13378,N_6315,N_5164);
and U13379 (N_13379,N_7203,N_6387);
and U13380 (N_13380,N_9199,N_8531);
nand U13381 (N_13381,N_5203,N_5501);
and U13382 (N_13382,N_6655,N_8347);
nand U13383 (N_13383,N_6803,N_9940);
and U13384 (N_13384,N_8553,N_7394);
or U13385 (N_13385,N_5136,N_5365);
and U13386 (N_13386,N_8217,N_6998);
nand U13387 (N_13387,N_9267,N_5681);
and U13388 (N_13388,N_6997,N_9967);
nand U13389 (N_13389,N_5756,N_6922);
xnor U13390 (N_13390,N_8774,N_5188);
and U13391 (N_13391,N_5641,N_6879);
nand U13392 (N_13392,N_6268,N_6878);
nand U13393 (N_13393,N_8864,N_9486);
xnor U13394 (N_13394,N_5415,N_6292);
xnor U13395 (N_13395,N_5771,N_5333);
nand U13396 (N_13396,N_8041,N_7481);
and U13397 (N_13397,N_6522,N_5750);
xor U13398 (N_13398,N_7270,N_9962);
nor U13399 (N_13399,N_8789,N_7439);
or U13400 (N_13400,N_6163,N_9143);
nand U13401 (N_13401,N_5997,N_5075);
xnor U13402 (N_13402,N_8853,N_7044);
or U13403 (N_13403,N_6697,N_8759);
or U13404 (N_13404,N_9626,N_9870);
nor U13405 (N_13405,N_9379,N_5949);
nand U13406 (N_13406,N_8885,N_6225);
nand U13407 (N_13407,N_8964,N_9010);
and U13408 (N_13408,N_9784,N_8501);
nor U13409 (N_13409,N_8122,N_7217);
or U13410 (N_13410,N_7404,N_7856);
and U13411 (N_13411,N_9557,N_5501);
nor U13412 (N_13412,N_8344,N_5723);
nand U13413 (N_13413,N_6570,N_6353);
or U13414 (N_13414,N_9959,N_5999);
and U13415 (N_13415,N_8240,N_6035);
xnor U13416 (N_13416,N_5922,N_6853);
nor U13417 (N_13417,N_6191,N_6637);
and U13418 (N_13418,N_8505,N_8341);
or U13419 (N_13419,N_6459,N_8279);
nand U13420 (N_13420,N_8114,N_7736);
nor U13421 (N_13421,N_5016,N_6419);
xnor U13422 (N_13422,N_9561,N_6444);
or U13423 (N_13423,N_7737,N_8834);
xnor U13424 (N_13424,N_9897,N_9289);
or U13425 (N_13425,N_8502,N_5850);
xor U13426 (N_13426,N_7140,N_7083);
and U13427 (N_13427,N_9624,N_5056);
nand U13428 (N_13428,N_5405,N_9381);
nand U13429 (N_13429,N_5994,N_9967);
nor U13430 (N_13430,N_7546,N_7886);
and U13431 (N_13431,N_5042,N_5258);
xnor U13432 (N_13432,N_8881,N_7469);
or U13433 (N_13433,N_5172,N_9940);
or U13434 (N_13434,N_5626,N_7513);
xnor U13435 (N_13435,N_7399,N_6395);
nand U13436 (N_13436,N_7274,N_9310);
and U13437 (N_13437,N_8257,N_5303);
or U13438 (N_13438,N_7262,N_7435);
nand U13439 (N_13439,N_7468,N_8108);
and U13440 (N_13440,N_9863,N_9430);
xnor U13441 (N_13441,N_9393,N_7787);
and U13442 (N_13442,N_9724,N_7394);
nand U13443 (N_13443,N_6549,N_5416);
nor U13444 (N_13444,N_5946,N_8508);
and U13445 (N_13445,N_6338,N_6974);
nor U13446 (N_13446,N_6584,N_6929);
or U13447 (N_13447,N_8150,N_7038);
xor U13448 (N_13448,N_8049,N_5234);
or U13449 (N_13449,N_8656,N_9839);
nor U13450 (N_13450,N_8933,N_8310);
nor U13451 (N_13451,N_7440,N_7024);
or U13452 (N_13452,N_6583,N_8305);
or U13453 (N_13453,N_5788,N_9967);
or U13454 (N_13454,N_9356,N_5959);
xor U13455 (N_13455,N_8568,N_9855);
xnor U13456 (N_13456,N_7033,N_5480);
xor U13457 (N_13457,N_8616,N_7769);
or U13458 (N_13458,N_5029,N_5545);
and U13459 (N_13459,N_9568,N_6967);
and U13460 (N_13460,N_8742,N_5398);
and U13461 (N_13461,N_8790,N_6147);
nor U13462 (N_13462,N_5424,N_5343);
or U13463 (N_13463,N_8549,N_5830);
and U13464 (N_13464,N_5960,N_9449);
and U13465 (N_13465,N_8991,N_9419);
and U13466 (N_13466,N_7091,N_8524);
nand U13467 (N_13467,N_5711,N_7210);
xnor U13468 (N_13468,N_8902,N_9266);
or U13469 (N_13469,N_8815,N_7914);
nor U13470 (N_13470,N_7647,N_7957);
and U13471 (N_13471,N_7901,N_8285);
nand U13472 (N_13472,N_9397,N_6719);
nand U13473 (N_13473,N_9037,N_6872);
and U13474 (N_13474,N_6980,N_8872);
nand U13475 (N_13475,N_5093,N_6441);
nor U13476 (N_13476,N_9075,N_5108);
xnor U13477 (N_13477,N_7584,N_8817);
and U13478 (N_13478,N_6127,N_5731);
xor U13479 (N_13479,N_9544,N_9969);
nand U13480 (N_13480,N_9756,N_6482);
and U13481 (N_13481,N_5589,N_6132);
nor U13482 (N_13482,N_6701,N_8548);
or U13483 (N_13483,N_7081,N_5391);
nor U13484 (N_13484,N_9747,N_5510);
xnor U13485 (N_13485,N_5575,N_9436);
nand U13486 (N_13486,N_6153,N_9236);
xor U13487 (N_13487,N_5490,N_6328);
xor U13488 (N_13488,N_9639,N_8252);
or U13489 (N_13489,N_5947,N_5633);
nand U13490 (N_13490,N_8423,N_8039);
and U13491 (N_13491,N_9931,N_5191);
and U13492 (N_13492,N_7488,N_9826);
and U13493 (N_13493,N_8933,N_8664);
nor U13494 (N_13494,N_7535,N_7582);
nand U13495 (N_13495,N_7839,N_8709);
and U13496 (N_13496,N_8924,N_5585);
and U13497 (N_13497,N_7374,N_6269);
or U13498 (N_13498,N_9723,N_8324);
nor U13499 (N_13499,N_6244,N_7085);
nor U13500 (N_13500,N_5030,N_7154);
and U13501 (N_13501,N_5679,N_6918);
and U13502 (N_13502,N_5646,N_7784);
and U13503 (N_13503,N_8552,N_7357);
nor U13504 (N_13504,N_8964,N_9135);
and U13505 (N_13505,N_9344,N_7179);
nor U13506 (N_13506,N_6661,N_7388);
xnor U13507 (N_13507,N_7328,N_8943);
or U13508 (N_13508,N_5578,N_7975);
or U13509 (N_13509,N_5929,N_8744);
or U13510 (N_13510,N_7484,N_9849);
nand U13511 (N_13511,N_9157,N_5848);
or U13512 (N_13512,N_6283,N_8675);
and U13513 (N_13513,N_9424,N_7695);
nor U13514 (N_13514,N_8442,N_9320);
and U13515 (N_13515,N_7088,N_8585);
nor U13516 (N_13516,N_8325,N_8724);
and U13517 (N_13517,N_8190,N_5501);
xnor U13518 (N_13518,N_5997,N_6091);
and U13519 (N_13519,N_8700,N_7101);
nand U13520 (N_13520,N_5976,N_6734);
xnor U13521 (N_13521,N_8576,N_5540);
xor U13522 (N_13522,N_5306,N_9793);
nand U13523 (N_13523,N_8061,N_5213);
nor U13524 (N_13524,N_6523,N_9983);
xor U13525 (N_13525,N_7015,N_8313);
or U13526 (N_13526,N_5434,N_5816);
or U13527 (N_13527,N_6990,N_7153);
xnor U13528 (N_13528,N_7024,N_6262);
and U13529 (N_13529,N_7618,N_8877);
and U13530 (N_13530,N_9033,N_8970);
nor U13531 (N_13531,N_5595,N_7358);
nand U13532 (N_13532,N_5560,N_6739);
or U13533 (N_13533,N_5307,N_7784);
xor U13534 (N_13534,N_7975,N_7016);
nor U13535 (N_13535,N_8308,N_9650);
xor U13536 (N_13536,N_6008,N_8623);
xnor U13537 (N_13537,N_9236,N_6246);
xnor U13538 (N_13538,N_6848,N_7212);
or U13539 (N_13539,N_9201,N_5776);
xor U13540 (N_13540,N_8860,N_5951);
and U13541 (N_13541,N_9055,N_5809);
xnor U13542 (N_13542,N_8315,N_6185);
nor U13543 (N_13543,N_7561,N_5203);
nand U13544 (N_13544,N_5203,N_5508);
xnor U13545 (N_13545,N_7005,N_5414);
nor U13546 (N_13546,N_5238,N_9567);
nor U13547 (N_13547,N_6157,N_9505);
xor U13548 (N_13548,N_8532,N_5051);
and U13549 (N_13549,N_5798,N_7990);
nand U13550 (N_13550,N_8830,N_8558);
xnor U13551 (N_13551,N_8385,N_6146);
and U13552 (N_13552,N_9993,N_5671);
nand U13553 (N_13553,N_5847,N_6608);
nand U13554 (N_13554,N_5869,N_5738);
and U13555 (N_13555,N_8824,N_9694);
nor U13556 (N_13556,N_9971,N_7680);
nor U13557 (N_13557,N_9149,N_9867);
or U13558 (N_13558,N_8708,N_7941);
nor U13559 (N_13559,N_6097,N_9343);
nand U13560 (N_13560,N_9446,N_6282);
nand U13561 (N_13561,N_7195,N_7276);
nor U13562 (N_13562,N_9536,N_5202);
nand U13563 (N_13563,N_6313,N_8377);
nand U13564 (N_13564,N_5481,N_9612);
or U13565 (N_13565,N_7564,N_7109);
xor U13566 (N_13566,N_5830,N_7248);
or U13567 (N_13567,N_5342,N_5014);
nand U13568 (N_13568,N_8863,N_6455);
nand U13569 (N_13569,N_7933,N_5459);
nand U13570 (N_13570,N_5034,N_8774);
nor U13571 (N_13571,N_5435,N_9390);
xnor U13572 (N_13572,N_7688,N_8733);
or U13573 (N_13573,N_6097,N_6424);
nor U13574 (N_13574,N_9883,N_8195);
or U13575 (N_13575,N_6721,N_5630);
xnor U13576 (N_13576,N_8631,N_8061);
xnor U13577 (N_13577,N_6422,N_5831);
nand U13578 (N_13578,N_9690,N_7933);
nor U13579 (N_13579,N_9741,N_7863);
xnor U13580 (N_13580,N_8113,N_9912);
nand U13581 (N_13581,N_8132,N_8334);
nor U13582 (N_13582,N_5043,N_6478);
or U13583 (N_13583,N_7871,N_5607);
nand U13584 (N_13584,N_6600,N_9457);
or U13585 (N_13585,N_7557,N_5509);
xnor U13586 (N_13586,N_5051,N_7106);
nor U13587 (N_13587,N_5756,N_5441);
xnor U13588 (N_13588,N_5319,N_7259);
or U13589 (N_13589,N_7995,N_7275);
and U13590 (N_13590,N_8817,N_6985);
nand U13591 (N_13591,N_7145,N_6589);
and U13592 (N_13592,N_7877,N_9125);
or U13593 (N_13593,N_8762,N_6646);
nor U13594 (N_13594,N_5302,N_6343);
and U13595 (N_13595,N_8069,N_6042);
xnor U13596 (N_13596,N_5327,N_5717);
nor U13597 (N_13597,N_8209,N_5606);
xor U13598 (N_13598,N_6924,N_8403);
or U13599 (N_13599,N_7131,N_5752);
or U13600 (N_13600,N_7803,N_9549);
xnor U13601 (N_13601,N_7507,N_5877);
xor U13602 (N_13602,N_5768,N_7671);
nand U13603 (N_13603,N_9008,N_7664);
nand U13604 (N_13604,N_7053,N_8795);
or U13605 (N_13605,N_6459,N_6385);
or U13606 (N_13606,N_5527,N_5433);
nand U13607 (N_13607,N_8964,N_8378);
xnor U13608 (N_13608,N_7835,N_6245);
xor U13609 (N_13609,N_5748,N_7310);
and U13610 (N_13610,N_7458,N_8585);
xnor U13611 (N_13611,N_5795,N_7512);
nor U13612 (N_13612,N_5930,N_9537);
nand U13613 (N_13613,N_9930,N_8761);
xor U13614 (N_13614,N_9817,N_8719);
xor U13615 (N_13615,N_9965,N_9850);
nand U13616 (N_13616,N_9198,N_8572);
and U13617 (N_13617,N_9223,N_8446);
nor U13618 (N_13618,N_5865,N_6438);
nor U13619 (N_13619,N_9188,N_8657);
nor U13620 (N_13620,N_5960,N_7021);
and U13621 (N_13621,N_7001,N_7110);
xnor U13622 (N_13622,N_6046,N_9694);
xor U13623 (N_13623,N_6977,N_9771);
xnor U13624 (N_13624,N_9996,N_7829);
nand U13625 (N_13625,N_9984,N_8334);
nand U13626 (N_13626,N_9214,N_9432);
xnor U13627 (N_13627,N_6800,N_7609);
nor U13628 (N_13628,N_6262,N_8207);
nand U13629 (N_13629,N_7097,N_5017);
and U13630 (N_13630,N_9627,N_7367);
or U13631 (N_13631,N_9148,N_8408);
nand U13632 (N_13632,N_5095,N_5148);
and U13633 (N_13633,N_8475,N_6709);
xnor U13634 (N_13634,N_8089,N_8470);
nor U13635 (N_13635,N_5943,N_5873);
nor U13636 (N_13636,N_9756,N_5798);
nor U13637 (N_13637,N_9192,N_6513);
and U13638 (N_13638,N_7768,N_7430);
and U13639 (N_13639,N_8306,N_6685);
or U13640 (N_13640,N_9588,N_8723);
nand U13641 (N_13641,N_6405,N_6663);
nand U13642 (N_13642,N_7055,N_6147);
xor U13643 (N_13643,N_5285,N_5199);
nand U13644 (N_13644,N_5536,N_6251);
nor U13645 (N_13645,N_5023,N_5723);
or U13646 (N_13646,N_5055,N_8922);
or U13647 (N_13647,N_9669,N_8657);
nor U13648 (N_13648,N_6468,N_9098);
xnor U13649 (N_13649,N_5595,N_8059);
nand U13650 (N_13650,N_8539,N_5272);
and U13651 (N_13651,N_9391,N_8765);
nor U13652 (N_13652,N_7238,N_5093);
xor U13653 (N_13653,N_7292,N_8295);
nand U13654 (N_13654,N_7176,N_9247);
xnor U13655 (N_13655,N_6426,N_9258);
xnor U13656 (N_13656,N_6251,N_8442);
xor U13657 (N_13657,N_9523,N_6232);
xor U13658 (N_13658,N_6616,N_9616);
xor U13659 (N_13659,N_9245,N_5148);
nand U13660 (N_13660,N_7123,N_8106);
nor U13661 (N_13661,N_8026,N_7521);
nand U13662 (N_13662,N_7218,N_7922);
xnor U13663 (N_13663,N_6431,N_5355);
nor U13664 (N_13664,N_6385,N_5596);
or U13665 (N_13665,N_6736,N_8438);
nor U13666 (N_13666,N_5488,N_7455);
nor U13667 (N_13667,N_5398,N_7713);
and U13668 (N_13668,N_6817,N_9979);
and U13669 (N_13669,N_7458,N_8060);
xor U13670 (N_13670,N_8447,N_6365);
or U13671 (N_13671,N_8272,N_9207);
or U13672 (N_13672,N_5890,N_6470);
xnor U13673 (N_13673,N_6982,N_8071);
nand U13674 (N_13674,N_7110,N_6891);
nand U13675 (N_13675,N_5198,N_8558);
and U13676 (N_13676,N_8682,N_6898);
or U13677 (N_13677,N_9301,N_8622);
and U13678 (N_13678,N_7547,N_8259);
xnor U13679 (N_13679,N_7780,N_6148);
and U13680 (N_13680,N_7626,N_6926);
xnor U13681 (N_13681,N_7999,N_5165);
nor U13682 (N_13682,N_6243,N_9061);
or U13683 (N_13683,N_5516,N_5598);
and U13684 (N_13684,N_8990,N_7011);
and U13685 (N_13685,N_5602,N_8870);
nand U13686 (N_13686,N_8239,N_8254);
and U13687 (N_13687,N_5349,N_6517);
and U13688 (N_13688,N_5518,N_5752);
xor U13689 (N_13689,N_9664,N_7490);
nor U13690 (N_13690,N_5208,N_8807);
and U13691 (N_13691,N_9544,N_7884);
nand U13692 (N_13692,N_5003,N_9753);
xnor U13693 (N_13693,N_9231,N_9283);
or U13694 (N_13694,N_6958,N_7983);
xor U13695 (N_13695,N_5338,N_6854);
xor U13696 (N_13696,N_8240,N_8767);
and U13697 (N_13697,N_6115,N_7462);
nand U13698 (N_13698,N_7927,N_6265);
nand U13699 (N_13699,N_5557,N_6422);
nand U13700 (N_13700,N_6171,N_5127);
nand U13701 (N_13701,N_7731,N_8330);
and U13702 (N_13702,N_9750,N_5839);
nand U13703 (N_13703,N_9783,N_8066);
nor U13704 (N_13704,N_8066,N_8380);
nor U13705 (N_13705,N_5533,N_9460);
nand U13706 (N_13706,N_6662,N_6934);
xor U13707 (N_13707,N_6250,N_8781);
and U13708 (N_13708,N_7466,N_8495);
xor U13709 (N_13709,N_6004,N_6922);
nand U13710 (N_13710,N_7472,N_9316);
nand U13711 (N_13711,N_5963,N_6408);
or U13712 (N_13712,N_7017,N_7131);
and U13713 (N_13713,N_7064,N_8233);
xor U13714 (N_13714,N_8630,N_8262);
and U13715 (N_13715,N_7265,N_7930);
nor U13716 (N_13716,N_9998,N_7383);
nor U13717 (N_13717,N_7643,N_9947);
nand U13718 (N_13718,N_7278,N_5219);
xor U13719 (N_13719,N_7225,N_6237);
and U13720 (N_13720,N_5626,N_7285);
nand U13721 (N_13721,N_5436,N_5520);
and U13722 (N_13722,N_5532,N_9285);
nor U13723 (N_13723,N_5621,N_8558);
or U13724 (N_13724,N_7409,N_6795);
nand U13725 (N_13725,N_9908,N_8390);
xnor U13726 (N_13726,N_5379,N_7564);
xor U13727 (N_13727,N_8922,N_7535);
nand U13728 (N_13728,N_9641,N_7451);
xnor U13729 (N_13729,N_6114,N_8164);
and U13730 (N_13730,N_5443,N_5369);
nand U13731 (N_13731,N_8431,N_6311);
nand U13732 (N_13732,N_6920,N_5362);
and U13733 (N_13733,N_8924,N_5237);
or U13734 (N_13734,N_6245,N_7810);
nand U13735 (N_13735,N_6654,N_9957);
nand U13736 (N_13736,N_9256,N_8080);
and U13737 (N_13737,N_9969,N_8031);
or U13738 (N_13738,N_5520,N_9346);
nor U13739 (N_13739,N_9756,N_9603);
and U13740 (N_13740,N_8994,N_6319);
nand U13741 (N_13741,N_7458,N_9848);
nor U13742 (N_13742,N_7909,N_9526);
nor U13743 (N_13743,N_9473,N_5004);
nand U13744 (N_13744,N_6719,N_8816);
and U13745 (N_13745,N_9832,N_6736);
nor U13746 (N_13746,N_8980,N_6931);
and U13747 (N_13747,N_9242,N_9913);
or U13748 (N_13748,N_9501,N_8299);
xor U13749 (N_13749,N_9521,N_9110);
nor U13750 (N_13750,N_6977,N_8679);
or U13751 (N_13751,N_7710,N_8209);
xor U13752 (N_13752,N_5118,N_6456);
or U13753 (N_13753,N_9567,N_8197);
and U13754 (N_13754,N_9921,N_5350);
nand U13755 (N_13755,N_5241,N_6082);
nor U13756 (N_13756,N_9161,N_8255);
nor U13757 (N_13757,N_9144,N_6658);
or U13758 (N_13758,N_5597,N_8300);
nor U13759 (N_13759,N_8568,N_6669);
nand U13760 (N_13760,N_6036,N_8058);
or U13761 (N_13761,N_9560,N_6008);
and U13762 (N_13762,N_5027,N_9544);
nand U13763 (N_13763,N_8855,N_6710);
or U13764 (N_13764,N_6101,N_6486);
nor U13765 (N_13765,N_6269,N_5026);
nand U13766 (N_13766,N_6130,N_9787);
or U13767 (N_13767,N_8449,N_5969);
and U13768 (N_13768,N_7274,N_9364);
nor U13769 (N_13769,N_9807,N_6093);
or U13770 (N_13770,N_7812,N_6250);
or U13771 (N_13771,N_9762,N_5904);
nand U13772 (N_13772,N_6075,N_9848);
nor U13773 (N_13773,N_6001,N_9419);
nand U13774 (N_13774,N_6465,N_5171);
nand U13775 (N_13775,N_5318,N_8892);
xnor U13776 (N_13776,N_9936,N_5900);
xnor U13777 (N_13777,N_6848,N_6907);
nor U13778 (N_13778,N_6846,N_7145);
or U13779 (N_13779,N_7872,N_8977);
xnor U13780 (N_13780,N_8154,N_8140);
xor U13781 (N_13781,N_5767,N_8974);
or U13782 (N_13782,N_6776,N_8698);
nor U13783 (N_13783,N_9213,N_8951);
nor U13784 (N_13784,N_5470,N_6159);
or U13785 (N_13785,N_9613,N_5355);
nand U13786 (N_13786,N_9448,N_9916);
or U13787 (N_13787,N_9913,N_8574);
and U13788 (N_13788,N_6297,N_5121);
or U13789 (N_13789,N_6652,N_9710);
nor U13790 (N_13790,N_8811,N_7734);
and U13791 (N_13791,N_9648,N_5314);
nor U13792 (N_13792,N_7111,N_9229);
xnor U13793 (N_13793,N_5771,N_8384);
and U13794 (N_13794,N_5220,N_7420);
nor U13795 (N_13795,N_6619,N_9894);
and U13796 (N_13796,N_9082,N_5093);
nor U13797 (N_13797,N_6181,N_8093);
nor U13798 (N_13798,N_5655,N_5393);
nand U13799 (N_13799,N_6163,N_9240);
xnor U13800 (N_13800,N_9637,N_7967);
and U13801 (N_13801,N_7282,N_6789);
nand U13802 (N_13802,N_6931,N_5309);
nor U13803 (N_13803,N_9680,N_5834);
xnor U13804 (N_13804,N_6174,N_7063);
and U13805 (N_13805,N_6639,N_8445);
xnor U13806 (N_13806,N_5921,N_6280);
or U13807 (N_13807,N_5661,N_5163);
and U13808 (N_13808,N_7809,N_8882);
xnor U13809 (N_13809,N_6711,N_5763);
nand U13810 (N_13810,N_5367,N_5889);
xor U13811 (N_13811,N_6516,N_7566);
or U13812 (N_13812,N_7006,N_7917);
or U13813 (N_13813,N_7708,N_6542);
and U13814 (N_13814,N_5732,N_9425);
nor U13815 (N_13815,N_8228,N_5629);
or U13816 (N_13816,N_6430,N_7571);
xnor U13817 (N_13817,N_8951,N_5883);
xnor U13818 (N_13818,N_5310,N_8461);
nor U13819 (N_13819,N_5246,N_7725);
and U13820 (N_13820,N_6111,N_7727);
or U13821 (N_13821,N_7319,N_6678);
nor U13822 (N_13822,N_8036,N_5084);
and U13823 (N_13823,N_9085,N_6766);
nand U13824 (N_13824,N_5633,N_7860);
and U13825 (N_13825,N_5099,N_5954);
xor U13826 (N_13826,N_7378,N_9381);
nor U13827 (N_13827,N_8982,N_7883);
xnor U13828 (N_13828,N_8003,N_9382);
nand U13829 (N_13829,N_9771,N_7657);
and U13830 (N_13830,N_9083,N_7273);
nand U13831 (N_13831,N_5901,N_7078);
nand U13832 (N_13832,N_5243,N_7192);
and U13833 (N_13833,N_5868,N_7048);
xnor U13834 (N_13834,N_6715,N_8564);
and U13835 (N_13835,N_8502,N_5490);
and U13836 (N_13836,N_7601,N_9577);
xnor U13837 (N_13837,N_7569,N_7377);
nor U13838 (N_13838,N_7397,N_9234);
or U13839 (N_13839,N_9748,N_9019);
xor U13840 (N_13840,N_8076,N_9771);
nor U13841 (N_13841,N_6116,N_9078);
nor U13842 (N_13842,N_9962,N_7973);
nand U13843 (N_13843,N_9345,N_8270);
and U13844 (N_13844,N_5888,N_6367);
and U13845 (N_13845,N_8410,N_7565);
and U13846 (N_13846,N_6954,N_6737);
xor U13847 (N_13847,N_9850,N_9552);
nor U13848 (N_13848,N_5678,N_6940);
or U13849 (N_13849,N_9176,N_8288);
and U13850 (N_13850,N_8583,N_8712);
nand U13851 (N_13851,N_5432,N_9919);
nand U13852 (N_13852,N_9797,N_5526);
nand U13853 (N_13853,N_9985,N_6675);
or U13854 (N_13854,N_9764,N_9592);
nand U13855 (N_13855,N_5824,N_6814);
and U13856 (N_13856,N_6265,N_8236);
nand U13857 (N_13857,N_8837,N_9309);
xnor U13858 (N_13858,N_6101,N_6795);
and U13859 (N_13859,N_6801,N_5622);
xor U13860 (N_13860,N_6225,N_9435);
xnor U13861 (N_13861,N_6708,N_8975);
nand U13862 (N_13862,N_9314,N_9350);
nand U13863 (N_13863,N_5759,N_5537);
nor U13864 (N_13864,N_5410,N_9514);
nand U13865 (N_13865,N_9816,N_7755);
nor U13866 (N_13866,N_6369,N_5594);
or U13867 (N_13867,N_6895,N_5467);
or U13868 (N_13868,N_6385,N_8085);
xor U13869 (N_13869,N_5449,N_9006);
nor U13870 (N_13870,N_5655,N_9417);
or U13871 (N_13871,N_9428,N_8105);
and U13872 (N_13872,N_9953,N_9830);
and U13873 (N_13873,N_8259,N_5565);
xor U13874 (N_13874,N_9320,N_5912);
nand U13875 (N_13875,N_9680,N_8481);
and U13876 (N_13876,N_7205,N_8724);
nor U13877 (N_13877,N_5745,N_5064);
nor U13878 (N_13878,N_9710,N_5451);
nor U13879 (N_13879,N_8066,N_7749);
and U13880 (N_13880,N_8716,N_6080);
nand U13881 (N_13881,N_6470,N_5711);
or U13882 (N_13882,N_9017,N_7471);
nor U13883 (N_13883,N_7217,N_5721);
nand U13884 (N_13884,N_6814,N_8749);
nand U13885 (N_13885,N_7011,N_7481);
and U13886 (N_13886,N_6811,N_8433);
xnor U13887 (N_13887,N_6873,N_5582);
or U13888 (N_13888,N_8072,N_7773);
or U13889 (N_13889,N_9280,N_8480);
and U13890 (N_13890,N_9144,N_9997);
xor U13891 (N_13891,N_5582,N_5741);
and U13892 (N_13892,N_5075,N_6239);
and U13893 (N_13893,N_5120,N_8966);
xor U13894 (N_13894,N_6793,N_7987);
nor U13895 (N_13895,N_9016,N_9550);
nor U13896 (N_13896,N_9587,N_9910);
nand U13897 (N_13897,N_8492,N_6941);
and U13898 (N_13898,N_8721,N_8864);
nand U13899 (N_13899,N_7596,N_5069);
nand U13900 (N_13900,N_5941,N_7463);
xor U13901 (N_13901,N_6063,N_9973);
xor U13902 (N_13902,N_7684,N_9121);
and U13903 (N_13903,N_7304,N_8102);
nand U13904 (N_13904,N_5227,N_6339);
nand U13905 (N_13905,N_9769,N_8053);
nor U13906 (N_13906,N_5365,N_5315);
xnor U13907 (N_13907,N_7734,N_9142);
xor U13908 (N_13908,N_6040,N_5643);
xor U13909 (N_13909,N_6199,N_8660);
nor U13910 (N_13910,N_7572,N_6327);
nor U13911 (N_13911,N_6548,N_6528);
xnor U13912 (N_13912,N_5838,N_6592);
or U13913 (N_13913,N_8609,N_5005);
xnor U13914 (N_13914,N_9227,N_6263);
xnor U13915 (N_13915,N_7348,N_9944);
and U13916 (N_13916,N_9909,N_9329);
nor U13917 (N_13917,N_9834,N_6346);
nor U13918 (N_13918,N_7191,N_6264);
nor U13919 (N_13919,N_9248,N_7857);
xor U13920 (N_13920,N_7420,N_8677);
nor U13921 (N_13921,N_5123,N_6344);
xor U13922 (N_13922,N_6718,N_5082);
nand U13923 (N_13923,N_7402,N_6570);
nor U13924 (N_13924,N_9062,N_9313);
and U13925 (N_13925,N_9705,N_7807);
or U13926 (N_13926,N_8655,N_6239);
nand U13927 (N_13927,N_5808,N_5755);
and U13928 (N_13928,N_9582,N_9954);
nor U13929 (N_13929,N_8114,N_9512);
xnor U13930 (N_13930,N_7721,N_8166);
or U13931 (N_13931,N_6578,N_6434);
or U13932 (N_13932,N_9379,N_8487);
xor U13933 (N_13933,N_8388,N_7679);
or U13934 (N_13934,N_7687,N_8678);
nand U13935 (N_13935,N_8134,N_5748);
nand U13936 (N_13936,N_5780,N_7776);
or U13937 (N_13937,N_5932,N_5851);
and U13938 (N_13938,N_7072,N_7046);
xor U13939 (N_13939,N_7974,N_7528);
nand U13940 (N_13940,N_5745,N_8111);
nor U13941 (N_13941,N_5861,N_9787);
nand U13942 (N_13942,N_7652,N_5056);
nand U13943 (N_13943,N_8063,N_5699);
nand U13944 (N_13944,N_8194,N_8808);
nor U13945 (N_13945,N_9354,N_7005);
nor U13946 (N_13946,N_6027,N_5605);
nand U13947 (N_13947,N_6217,N_9332);
or U13948 (N_13948,N_8092,N_7137);
nor U13949 (N_13949,N_7065,N_6328);
nor U13950 (N_13950,N_9673,N_6380);
xor U13951 (N_13951,N_5492,N_5514);
nor U13952 (N_13952,N_7283,N_6521);
or U13953 (N_13953,N_9040,N_6884);
xor U13954 (N_13954,N_6882,N_6945);
xor U13955 (N_13955,N_8211,N_9622);
nor U13956 (N_13956,N_9483,N_5380);
and U13957 (N_13957,N_7174,N_6282);
nand U13958 (N_13958,N_6776,N_5756);
or U13959 (N_13959,N_5361,N_6520);
and U13960 (N_13960,N_9355,N_6606);
or U13961 (N_13961,N_7980,N_6172);
and U13962 (N_13962,N_6938,N_8440);
or U13963 (N_13963,N_8393,N_9943);
and U13964 (N_13964,N_7372,N_6756);
nand U13965 (N_13965,N_9754,N_9531);
nor U13966 (N_13966,N_5969,N_7413);
and U13967 (N_13967,N_5061,N_5016);
nor U13968 (N_13968,N_9924,N_9381);
or U13969 (N_13969,N_8835,N_7786);
or U13970 (N_13970,N_6156,N_6391);
xnor U13971 (N_13971,N_5067,N_9529);
nor U13972 (N_13972,N_5562,N_5693);
xor U13973 (N_13973,N_6381,N_5948);
xor U13974 (N_13974,N_5786,N_7550);
or U13975 (N_13975,N_6450,N_6736);
nand U13976 (N_13976,N_8770,N_9101);
and U13977 (N_13977,N_7414,N_7982);
or U13978 (N_13978,N_6083,N_8136);
or U13979 (N_13979,N_8334,N_7204);
xor U13980 (N_13980,N_8645,N_6822);
and U13981 (N_13981,N_7225,N_8397);
nand U13982 (N_13982,N_6980,N_9085);
nand U13983 (N_13983,N_8336,N_6310);
nor U13984 (N_13984,N_9214,N_9973);
or U13985 (N_13985,N_6104,N_6511);
nand U13986 (N_13986,N_5118,N_7101);
nand U13987 (N_13987,N_6881,N_5537);
nor U13988 (N_13988,N_9571,N_5576);
or U13989 (N_13989,N_5766,N_9092);
and U13990 (N_13990,N_9001,N_8630);
nand U13991 (N_13991,N_9624,N_8141);
nand U13992 (N_13992,N_5922,N_7506);
and U13993 (N_13993,N_5591,N_8996);
xor U13994 (N_13994,N_7146,N_7916);
nor U13995 (N_13995,N_8966,N_6148);
and U13996 (N_13996,N_8142,N_9382);
or U13997 (N_13997,N_7072,N_8935);
nor U13998 (N_13998,N_5318,N_8837);
or U13999 (N_13999,N_5379,N_6266);
nand U14000 (N_14000,N_8272,N_5460);
or U14001 (N_14001,N_8479,N_7451);
nand U14002 (N_14002,N_7359,N_8741);
nor U14003 (N_14003,N_8761,N_6439);
nand U14004 (N_14004,N_9105,N_7440);
nor U14005 (N_14005,N_6178,N_8460);
xor U14006 (N_14006,N_8014,N_5048);
or U14007 (N_14007,N_7040,N_8009);
nand U14008 (N_14008,N_6256,N_5867);
or U14009 (N_14009,N_5291,N_6009);
nor U14010 (N_14010,N_7460,N_8217);
nand U14011 (N_14011,N_5560,N_8361);
xnor U14012 (N_14012,N_8105,N_6803);
xnor U14013 (N_14013,N_7940,N_8494);
nor U14014 (N_14014,N_5085,N_9190);
and U14015 (N_14015,N_9970,N_9074);
and U14016 (N_14016,N_5223,N_7985);
xor U14017 (N_14017,N_5565,N_8645);
nor U14018 (N_14018,N_6277,N_6951);
and U14019 (N_14019,N_5968,N_6467);
and U14020 (N_14020,N_7164,N_9297);
or U14021 (N_14021,N_5680,N_8055);
nor U14022 (N_14022,N_6762,N_7662);
xor U14023 (N_14023,N_7204,N_6547);
and U14024 (N_14024,N_9172,N_5027);
xor U14025 (N_14025,N_5362,N_7492);
xor U14026 (N_14026,N_6562,N_6345);
and U14027 (N_14027,N_5072,N_7713);
or U14028 (N_14028,N_5108,N_8623);
nor U14029 (N_14029,N_5571,N_9964);
or U14030 (N_14030,N_8069,N_8395);
and U14031 (N_14031,N_8821,N_9663);
nor U14032 (N_14032,N_8112,N_7096);
nor U14033 (N_14033,N_6736,N_8139);
nor U14034 (N_14034,N_5716,N_5931);
nor U14035 (N_14035,N_6979,N_5366);
nor U14036 (N_14036,N_5174,N_8140);
nand U14037 (N_14037,N_8851,N_5192);
nand U14038 (N_14038,N_8567,N_8348);
and U14039 (N_14039,N_7946,N_6577);
and U14040 (N_14040,N_9898,N_8576);
and U14041 (N_14041,N_8610,N_9382);
or U14042 (N_14042,N_6412,N_6405);
and U14043 (N_14043,N_5499,N_7219);
nand U14044 (N_14044,N_8259,N_9252);
nor U14045 (N_14045,N_5816,N_5122);
xnor U14046 (N_14046,N_7638,N_5478);
nand U14047 (N_14047,N_6818,N_7283);
nor U14048 (N_14048,N_8498,N_9787);
nand U14049 (N_14049,N_9322,N_5931);
and U14050 (N_14050,N_6210,N_7745);
and U14051 (N_14051,N_7009,N_7907);
nor U14052 (N_14052,N_6936,N_6046);
xor U14053 (N_14053,N_7700,N_5877);
nand U14054 (N_14054,N_6917,N_9179);
xnor U14055 (N_14055,N_6818,N_7070);
nand U14056 (N_14056,N_6214,N_7683);
nor U14057 (N_14057,N_8280,N_5750);
nand U14058 (N_14058,N_6839,N_9465);
nand U14059 (N_14059,N_9533,N_7407);
or U14060 (N_14060,N_5090,N_9406);
nor U14061 (N_14061,N_5282,N_5631);
and U14062 (N_14062,N_8863,N_7191);
nand U14063 (N_14063,N_6938,N_7919);
and U14064 (N_14064,N_9469,N_5396);
and U14065 (N_14065,N_8960,N_7231);
xnor U14066 (N_14066,N_9766,N_9777);
xnor U14067 (N_14067,N_5309,N_9575);
or U14068 (N_14068,N_8098,N_7711);
nand U14069 (N_14069,N_5633,N_8086);
nand U14070 (N_14070,N_6375,N_9206);
nand U14071 (N_14071,N_8079,N_5746);
xnor U14072 (N_14072,N_6470,N_6594);
nand U14073 (N_14073,N_5711,N_5684);
xnor U14074 (N_14074,N_7666,N_8887);
nor U14075 (N_14075,N_9138,N_7342);
and U14076 (N_14076,N_8930,N_5676);
nand U14077 (N_14077,N_7823,N_5338);
and U14078 (N_14078,N_9029,N_7540);
nand U14079 (N_14079,N_8694,N_5639);
nand U14080 (N_14080,N_9194,N_7613);
and U14081 (N_14081,N_5556,N_5432);
and U14082 (N_14082,N_5873,N_7100);
or U14083 (N_14083,N_6885,N_9409);
and U14084 (N_14084,N_5007,N_5141);
or U14085 (N_14085,N_9832,N_8967);
nor U14086 (N_14086,N_5985,N_5563);
or U14087 (N_14087,N_8496,N_5939);
or U14088 (N_14088,N_5354,N_6809);
or U14089 (N_14089,N_6930,N_5415);
nor U14090 (N_14090,N_5209,N_9923);
nor U14091 (N_14091,N_5856,N_8635);
nand U14092 (N_14092,N_9531,N_9232);
xor U14093 (N_14093,N_9075,N_6221);
nand U14094 (N_14094,N_6932,N_5585);
or U14095 (N_14095,N_8523,N_6954);
and U14096 (N_14096,N_8451,N_5855);
nor U14097 (N_14097,N_9325,N_9259);
or U14098 (N_14098,N_8755,N_9089);
xor U14099 (N_14099,N_6404,N_5736);
or U14100 (N_14100,N_6168,N_5627);
nand U14101 (N_14101,N_5255,N_6704);
or U14102 (N_14102,N_6488,N_9650);
or U14103 (N_14103,N_8814,N_6567);
xor U14104 (N_14104,N_6616,N_8183);
nor U14105 (N_14105,N_8090,N_5429);
and U14106 (N_14106,N_5313,N_8866);
xor U14107 (N_14107,N_6349,N_9188);
nor U14108 (N_14108,N_7607,N_5529);
or U14109 (N_14109,N_6993,N_6474);
nand U14110 (N_14110,N_5715,N_7695);
xnor U14111 (N_14111,N_8913,N_9753);
xnor U14112 (N_14112,N_6930,N_5942);
nor U14113 (N_14113,N_8572,N_9446);
xor U14114 (N_14114,N_8038,N_9292);
nand U14115 (N_14115,N_9307,N_5474);
nor U14116 (N_14116,N_7423,N_5364);
and U14117 (N_14117,N_6749,N_7539);
xor U14118 (N_14118,N_7290,N_6544);
nor U14119 (N_14119,N_6953,N_5172);
or U14120 (N_14120,N_7787,N_7114);
nand U14121 (N_14121,N_6315,N_7459);
nor U14122 (N_14122,N_5571,N_6518);
and U14123 (N_14123,N_9343,N_8693);
nor U14124 (N_14124,N_5340,N_5866);
and U14125 (N_14125,N_8574,N_8225);
xor U14126 (N_14126,N_9868,N_9903);
and U14127 (N_14127,N_8104,N_5634);
xnor U14128 (N_14128,N_6288,N_7681);
and U14129 (N_14129,N_6937,N_8288);
nor U14130 (N_14130,N_6938,N_9634);
nor U14131 (N_14131,N_6024,N_6235);
nand U14132 (N_14132,N_8521,N_7944);
nand U14133 (N_14133,N_5028,N_8579);
nand U14134 (N_14134,N_9838,N_6387);
and U14135 (N_14135,N_7449,N_6256);
nor U14136 (N_14136,N_8431,N_9048);
nand U14137 (N_14137,N_8087,N_7291);
and U14138 (N_14138,N_7128,N_5501);
nor U14139 (N_14139,N_8428,N_7430);
xnor U14140 (N_14140,N_6158,N_7341);
xor U14141 (N_14141,N_7039,N_5780);
or U14142 (N_14142,N_8600,N_8896);
nor U14143 (N_14143,N_9702,N_6702);
xor U14144 (N_14144,N_9565,N_6861);
xnor U14145 (N_14145,N_8041,N_5052);
and U14146 (N_14146,N_5602,N_8381);
nand U14147 (N_14147,N_5649,N_8038);
nor U14148 (N_14148,N_8372,N_7624);
or U14149 (N_14149,N_8932,N_9896);
and U14150 (N_14150,N_8961,N_5012);
and U14151 (N_14151,N_6148,N_5436);
nor U14152 (N_14152,N_9852,N_6043);
nor U14153 (N_14153,N_8445,N_9396);
or U14154 (N_14154,N_7938,N_5004);
nand U14155 (N_14155,N_5384,N_5859);
xnor U14156 (N_14156,N_9360,N_9036);
and U14157 (N_14157,N_6843,N_7168);
xor U14158 (N_14158,N_7527,N_7218);
xnor U14159 (N_14159,N_8784,N_8251);
or U14160 (N_14160,N_9917,N_9218);
or U14161 (N_14161,N_5203,N_5826);
xnor U14162 (N_14162,N_7921,N_8508);
or U14163 (N_14163,N_8634,N_7652);
nand U14164 (N_14164,N_8959,N_9126);
xor U14165 (N_14165,N_9118,N_8999);
nor U14166 (N_14166,N_6929,N_7414);
nand U14167 (N_14167,N_5727,N_8130);
xnor U14168 (N_14168,N_6310,N_5840);
nand U14169 (N_14169,N_6703,N_9254);
nor U14170 (N_14170,N_5024,N_5650);
or U14171 (N_14171,N_6595,N_6893);
and U14172 (N_14172,N_5549,N_5621);
and U14173 (N_14173,N_5877,N_8362);
xor U14174 (N_14174,N_7929,N_7525);
nor U14175 (N_14175,N_5708,N_7879);
xor U14176 (N_14176,N_7531,N_7462);
or U14177 (N_14177,N_8580,N_9577);
nand U14178 (N_14178,N_5335,N_5205);
or U14179 (N_14179,N_6812,N_8092);
nand U14180 (N_14180,N_5579,N_6188);
or U14181 (N_14181,N_7640,N_6583);
or U14182 (N_14182,N_8053,N_7073);
or U14183 (N_14183,N_8666,N_7228);
nand U14184 (N_14184,N_7666,N_7655);
and U14185 (N_14185,N_9355,N_7293);
nand U14186 (N_14186,N_6984,N_7100);
nor U14187 (N_14187,N_6839,N_6701);
or U14188 (N_14188,N_7426,N_9226);
xor U14189 (N_14189,N_5901,N_9114);
or U14190 (N_14190,N_6684,N_5007);
or U14191 (N_14191,N_8429,N_6714);
or U14192 (N_14192,N_6542,N_6208);
and U14193 (N_14193,N_5221,N_6069);
nand U14194 (N_14194,N_6257,N_8291);
nand U14195 (N_14195,N_8818,N_7226);
or U14196 (N_14196,N_9594,N_6826);
nand U14197 (N_14197,N_5656,N_8338);
or U14198 (N_14198,N_8827,N_9354);
and U14199 (N_14199,N_9778,N_7213);
nand U14200 (N_14200,N_9715,N_6920);
xor U14201 (N_14201,N_6907,N_5112);
or U14202 (N_14202,N_7625,N_8473);
and U14203 (N_14203,N_9006,N_7133);
nand U14204 (N_14204,N_8785,N_6226);
nand U14205 (N_14205,N_6406,N_8464);
nor U14206 (N_14206,N_5785,N_8561);
or U14207 (N_14207,N_7568,N_9518);
nor U14208 (N_14208,N_6312,N_9516);
nor U14209 (N_14209,N_6114,N_7237);
or U14210 (N_14210,N_7611,N_9023);
xnor U14211 (N_14211,N_6882,N_9840);
or U14212 (N_14212,N_5437,N_7266);
or U14213 (N_14213,N_5539,N_8074);
xor U14214 (N_14214,N_8123,N_8804);
and U14215 (N_14215,N_6727,N_6444);
xor U14216 (N_14216,N_9957,N_7929);
xor U14217 (N_14217,N_7721,N_5224);
nor U14218 (N_14218,N_9776,N_6414);
nor U14219 (N_14219,N_9662,N_9702);
xnor U14220 (N_14220,N_8152,N_7492);
nand U14221 (N_14221,N_6814,N_7313);
nor U14222 (N_14222,N_8396,N_5596);
nor U14223 (N_14223,N_5159,N_5728);
nor U14224 (N_14224,N_8358,N_9499);
and U14225 (N_14225,N_6597,N_6584);
nand U14226 (N_14226,N_6182,N_9888);
nand U14227 (N_14227,N_6229,N_6274);
and U14228 (N_14228,N_9556,N_8978);
nor U14229 (N_14229,N_5574,N_5103);
nand U14230 (N_14230,N_8506,N_7073);
nand U14231 (N_14231,N_9282,N_6117);
nand U14232 (N_14232,N_6162,N_9700);
nand U14233 (N_14233,N_8942,N_8163);
nor U14234 (N_14234,N_5925,N_6436);
and U14235 (N_14235,N_5939,N_5053);
and U14236 (N_14236,N_6037,N_9896);
xnor U14237 (N_14237,N_8950,N_5200);
and U14238 (N_14238,N_9217,N_5593);
nand U14239 (N_14239,N_6552,N_5926);
or U14240 (N_14240,N_7390,N_8840);
xor U14241 (N_14241,N_7857,N_9432);
nor U14242 (N_14242,N_6383,N_5532);
nor U14243 (N_14243,N_6004,N_6628);
or U14244 (N_14244,N_8807,N_6649);
xor U14245 (N_14245,N_5107,N_9774);
or U14246 (N_14246,N_6609,N_9371);
xor U14247 (N_14247,N_5969,N_7317);
nor U14248 (N_14248,N_5448,N_5073);
or U14249 (N_14249,N_7542,N_7158);
and U14250 (N_14250,N_9886,N_8464);
nand U14251 (N_14251,N_5977,N_5903);
xnor U14252 (N_14252,N_5389,N_8428);
nand U14253 (N_14253,N_5793,N_7618);
nand U14254 (N_14254,N_8316,N_6973);
nor U14255 (N_14255,N_7042,N_9730);
or U14256 (N_14256,N_6134,N_6877);
nor U14257 (N_14257,N_5984,N_9192);
xnor U14258 (N_14258,N_9533,N_5720);
xor U14259 (N_14259,N_9921,N_9481);
and U14260 (N_14260,N_9258,N_9919);
and U14261 (N_14261,N_9982,N_6268);
or U14262 (N_14262,N_8595,N_9358);
or U14263 (N_14263,N_9441,N_6370);
or U14264 (N_14264,N_6988,N_5999);
and U14265 (N_14265,N_9793,N_7020);
or U14266 (N_14266,N_6363,N_6543);
and U14267 (N_14267,N_9450,N_6074);
or U14268 (N_14268,N_5162,N_5935);
nor U14269 (N_14269,N_7340,N_5346);
or U14270 (N_14270,N_9439,N_8324);
nand U14271 (N_14271,N_5029,N_9471);
xor U14272 (N_14272,N_9012,N_9061);
nor U14273 (N_14273,N_7586,N_9669);
or U14274 (N_14274,N_6862,N_6020);
and U14275 (N_14275,N_5971,N_7710);
or U14276 (N_14276,N_8110,N_8419);
nor U14277 (N_14277,N_8780,N_6231);
nand U14278 (N_14278,N_7000,N_9428);
and U14279 (N_14279,N_6129,N_7610);
nand U14280 (N_14280,N_5089,N_7457);
or U14281 (N_14281,N_6864,N_6147);
xor U14282 (N_14282,N_5678,N_5026);
nand U14283 (N_14283,N_7526,N_5652);
or U14284 (N_14284,N_7010,N_7447);
xnor U14285 (N_14285,N_9368,N_5614);
or U14286 (N_14286,N_8831,N_8481);
and U14287 (N_14287,N_8025,N_7353);
nor U14288 (N_14288,N_9682,N_5107);
xor U14289 (N_14289,N_8281,N_8403);
nand U14290 (N_14290,N_6091,N_8310);
xor U14291 (N_14291,N_6513,N_5706);
xor U14292 (N_14292,N_6958,N_6285);
xor U14293 (N_14293,N_6789,N_6808);
xor U14294 (N_14294,N_5271,N_9775);
and U14295 (N_14295,N_7642,N_8098);
xnor U14296 (N_14296,N_6019,N_6612);
nor U14297 (N_14297,N_5295,N_5766);
nor U14298 (N_14298,N_5992,N_9407);
nand U14299 (N_14299,N_8947,N_6381);
nand U14300 (N_14300,N_7585,N_6465);
xnor U14301 (N_14301,N_6905,N_8227);
nand U14302 (N_14302,N_5112,N_6425);
or U14303 (N_14303,N_6008,N_6426);
nand U14304 (N_14304,N_8147,N_5504);
and U14305 (N_14305,N_7257,N_9222);
and U14306 (N_14306,N_7477,N_8073);
xnor U14307 (N_14307,N_6171,N_6509);
or U14308 (N_14308,N_6080,N_7591);
or U14309 (N_14309,N_7808,N_5052);
or U14310 (N_14310,N_5050,N_5793);
nand U14311 (N_14311,N_8909,N_5642);
and U14312 (N_14312,N_8843,N_9196);
and U14313 (N_14313,N_8562,N_9684);
and U14314 (N_14314,N_6873,N_7662);
xor U14315 (N_14315,N_7170,N_8927);
or U14316 (N_14316,N_5926,N_7197);
xnor U14317 (N_14317,N_5888,N_9982);
xnor U14318 (N_14318,N_8732,N_6781);
xor U14319 (N_14319,N_8798,N_6983);
and U14320 (N_14320,N_9246,N_8395);
xnor U14321 (N_14321,N_7021,N_9545);
nor U14322 (N_14322,N_6562,N_9953);
or U14323 (N_14323,N_5253,N_6828);
xnor U14324 (N_14324,N_7388,N_6128);
or U14325 (N_14325,N_8835,N_9655);
and U14326 (N_14326,N_6113,N_9962);
nand U14327 (N_14327,N_9150,N_9602);
and U14328 (N_14328,N_6205,N_8567);
or U14329 (N_14329,N_5132,N_9296);
nor U14330 (N_14330,N_9927,N_5643);
nor U14331 (N_14331,N_7578,N_7543);
nand U14332 (N_14332,N_7551,N_8197);
nor U14333 (N_14333,N_9780,N_7756);
xor U14334 (N_14334,N_9505,N_5110);
nor U14335 (N_14335,N_7669,N_9331);
nand U14336 (N_14336,N_9147,N_8752);
and U14337 (N_14337,N_6217,N_6956);
or U14338 (N_14338,N_5893,N_7469);
or U14339 (N_14339,N_6387,N_8670);
nand U14340 (N_14340,N_8332,N_7765);
nor U14341 (N_14341,N_8723,N_6290);
and U14342 (N_14342,N_8746,N_5031);
and U14343 (N_14343,N_8394,N_9992);
xor U14344 (N_14344,N_5219,N_9587);
nand U14345 (N_14345,N_8034,N_7192);
nor U14346 (N_14346,N_5648,N_7010);
nand U14347 (N_14347,N_6494,N_8082);
nand U14348 (N_14348,N_7770,N_7703);
nor U14349 (N_14349,N_5449,N_8016);
nand U14350 (N_14350,N_5518,N_5252);
nor U14351 (N_14351,N_6506,N_5330);
xnor U14352 (N_14352,N_9547,N_7763);
nand U14353 (N_14353,N_5738,N_8311);
and U14354 (N_14354,N_6549,N_5151);
nand U14355 (N_14355,N_6480,N_8795);
nand U14356 (N_14356,N_5932,N_8863);
nor U14357 (N_14357,N_7205,N_8992);
nand U14358 (N_14358,N_6546,N_7086);
or U14359 (N_14359,N_5602,N_6573);
nand U14360 (N_14360,N_8074,N_7760);
nand U14361 (N_14361,N_7747,N_5945);
xor U14362 (N_14362,N_5604,N_7779);
nor U14363 (N_14363,N_8512,N_9746);
nor U14364 (N_14364,N_7563,N_6030);
or U14365 (N_14365,N_7991,N_9041);
and U14366 (N_14366,N_7471,N_7525);
xor U14367 (N_14367,N_6746,N_7873);
and U14368 (N_14368,N_6875,N_8627);
nor U14369 (N_14369,N_7673,N_9781);
and U14370 (N_14370,N_6672,N_8383);
nand U14371 (N_14371,N_5417,N_9973);
nand U14372 (N_14372,N_7358,N_9214);
xnor U14373 (N_14373,N_6429,N_9988);
or U14374 (N_14374,N_7486,N_7679);
nor U14375 (N_14375,N_8576,N_7235);
xnor U14376 (N_14376,N_8284,N_5160);
nor U14377 (N_14377,N_5114,N_5955);
xnor U14378 (N_14378,N_8332,N_9305);
xor U14379 (N_14379,N_8644,N_7936);
or U14380 (N_14380,N_7093,N_9194);
xor U14381 (N_14381,N_6257,N_7146);
or U14382 (N_14382,N_8921,N_5335);
nor U14383 (N_14383,N_6675,N_8420);
nand U14384 (N_14384,N_7081,N_6071);
nand U14385 (N_14385,N_6113,N_6377);
nor U14386 (N_14386,N_7324,N_8749);
nor U14387 (N_14387,N_6625,N_9498);
and U14388 (N_14388,N_6460,N_9499);
xor U14389 (N_14389,N_5491,N_9201);
nand U14390 (N_14390,N_5460,N_5769);
and U14391 (N_14391,N_5441,N_9155);
or U14392 (N_14392,N_7028,N_5076);
nor U14393 (N_14393,N_7182,N_6102);
or U14394 (N_14394,N_5214,N_6416);
or U14395 (N_14395,N_9214,N_6577);
xor U14396 (N_14396,N_7747,N_9522);
or U14397 (N_14397,N_8964,N_7879);
xor U14398 (N_14398,N_9428,N_6050);
or U14399 (N_14399,N_7304,N_8114);
and U14400 (N_14400,N_5670,N_6418);
nand U14401 (N_14401,N_9688,N_8525);
xnor U14402 (N_14402,N_8427,N_5739);
nand U14403 (N_14403,N_9243,N_8346);
xnor U14404 (N_14404,N_7763,N_8572);
xnor U14405 (N_14405,N_9674,N_5215);
nor U14406 (N_14406,N_7718,N_5736);
nand U14407 (N_14407,N_6625,N_5831);
or U14408 (N_14408,N_7336,N_5985);
nand U14409 (N_14409,N_5598,N_9297);
and U14410 (N_14410,N_6817,N_7254);
or U14411 (N_14411,N_8970,N_8004);
or U14412 (N_14412,N_7445,N_9657);
xor U14413 (N_14413,N_5406,N_5233);
xnor U14414 (N_14414,N_9775,N_8103);
or U14415 (N_14415,N_5805,N_6072);
or U14416 (N_14416,N_6309,N_7888);
nand U14417 (N_14417,N_6553,N_5696);
xor U14418 (N_14418,N_6647,N_9471);
nand U14419 (N_14419,N_8460,N_8142);
nor U14420 (N_14420,N_5389,N_9004);
or U14421 (N_14421,N_7570,N_6946);
and U14422 (N_14422,N_7389,N_8696);
nand U14423 (N_14423,N_7572,N_6748);
and U14424 (N_14424,N_9337,N_7503);
nand U14425 (N_14425,N_9675,N_7006);
nand U14426 (N_14426,N_6004,N_6008);
nor U14427 (N_14427,N_7035,N_6519);
or U14428 (N_14428,N_6333,N_6630);
or U14429 (N_14429,N_6262,N_9263);
and U14430 (N_14430,N_5762,N_9101);
and U14431 (N_14431,N_8132,N_6397);
nand U14432 (N_14432,N_9907,N_6319);
and U14433 (N_14433,N_9750,N_7913);
nand U14434 (N_14434,N_8892,N_5687);
or U14435 (N_14435,N_9452,N_5737);
or U14436 (N_14436,N_6930,N_6870);
xnor U14437 (N_14437,N_8887,N_8610);
xor U14438 (N_14438,N_7787,N_5752);
and U14439 (N_14439,N_5191,N_6461);
nand U14440 (N_14440,N_5478,N_6661);
and U14441 (N_14441,N_5320,N_6654);
nor U14442 (N_14442,N_6771,N_8795);
or U14443 (N_14443,N_8524,N_7370);
nor U14444 (N_14444,N_5422,N_9143);
nor U14445 (N_14445,N_5401,N_8570);
nand U14446 (N_14446,N_7958,N_7279);
nand U14447 (N_14447,N_9182,N_9996);
xnor U14448 (N_14448,N_6234,N_9212);
or U14449 (N_14449,N_7469,N_6633);
and U14450 (N_14450,N_9566,N_7236);
xnor U14451 (N_14451,N_8669,N_7562);
nand U14452 (N_14452,N_5694,N_8709);
nand U14453 (N_14453,N_9233,N_7376);
or U14454 (N_14454,N_8130,N_9471);
nand U14455 (N_14455,N_7422,N_7300);
nand U14456 (N_14456,N_6465,N_9386);
or U14457 (N_14457,N_7155,N_6912);
xor U14458 (N_14458,N_5895,N_5475);
nand U14459 (N_14459,N_5472,N_6478);
nor U14460 (N_14460,N_5333,N_5441);
nor U14461 (N_14461,N_8972,N_5667);
nand U14462 (N_14462,N_7595,N_5429);
or U14463 (N_14463,N_8495,N_7574);
and U14464 (N_14464,N_9702,N_7399);
xor U14465 (N_14465,N_6787,N_8927);
and U14466 (N_14466,N_7487,N_9383);
nor U14467 (N_14467,N_7721,N_8552);
or U14468 (N_14468,N_6141,N_7098);
or U14469 (N_14469,N_7536,N_5722);
nand U14470 (N_14470,N_7552,N_8922);
nand U14471 (N_14471,N_9348,N_8622);
or U14472 (N_14472,N_8603,N_8939);
nor U14473 (N_14473,N_5762,N_9472);
nor U14474 (N_14474,N_7480,N_7973);
and U14475 (N_14475,N_7475,N_6282);
nand U14476 (N_14476,N_5722,N_6046);
and U14477 (N_14477,N_5766,N_5482);
xnor U14478 (N_14478,N_5152,N_6698);
and U14479 (N_14479,N_7778,N_7863);
nor U14480 (N_14480,N_7469,N_5682);
nand U14481 (N_14481,N_6895,N_6496);
or U14482 (N_14482,N_5498,N_5011);
xor U14483 (N_14483,N_6957,N_6461);
xor U14484 (N_14484,N_9058,N_6120);
xor U14485 (N_14485,N_7656,N_5693);
or U14486 (N_14486,N_6629,N_7535);
xnor U14487 (N_14487,N_5655,N_8239);
xnor U14488 (N_14488,N_9872,N_5592);
nand U14489 (N_14489,N_9847,N_6932);
nor U14490 (N_14490,N_6234,N_6746);
nand U14491 (N_14491,N_6704,N_8000);
and U14492 (N_14492,N_6827,N_7450);
and U14493 (N_14493,N_7895,N_5930);
and U14494 (N_14494,N_8531,N_9895);
nor U14495 (N_14495,N_8867,N_6928);
or U14496 (N_14496,N_9269,N_8968);
nor U14497 (N_14497,N_9007,N_5070);
nor U14498 (N_14498,N_8202,N_9843);
and U14499 (N_14499,N_9787,N_7454);
nor U14500 (N_14500,N_5820,N_9904);
nand U14501 (N_14501,N_7819,N_8214);
and U14502 (N_14502,N_6989,N_7556);
and U14503 (N_14503,N_9711,N_6439);
xnor U14504 (N_14504,N_9353,N_5319);
xor U14505 (N_14505,N_6632,N_8840);
or U14506 (N_14506,N_8439,N_8659);
nand U14507 (N_14507,N_5345,N_5399);
nand U14508 (N_14508,N_7196,N_9466);
and U14509 (N_14509,N_5384,N_6473);
nand U14510 (N_14510,N_5602,N_9531);
nand U14511 (N_14511,N_9723,N_7792);
nor U14512 (N_14512,N_6190,N_7990);
nor U14513 (N_14513,N_9265,N_9917);
xor U14514 (N_14514,N_7941,N_7985);
xor U14515 (N_14515,N_6093,N_9780);
nor U14516 (N_14516,N_5579,N_8946);
nand U14517 (N_14517,N_9282,N_8245);
and U14518 (N_14518,N_9595,N_6579);
xor U14519 (N_14519,N_7377,N_7522);
nor U14520 (N_14520,N_7977,N_9923);
nor U14521 (N_14521,N_5985,N_6535);
nor U14522 (N_14522,N_6206,N_8137);
xor U14523 (N_14523,N_7575,N_6003);
and U14524 (N_14524,N_7293,N_7936);
nand U14525 (N_14525,N_7246,N_9194);
nand U14526 (N_14526,N_8964,N_9693);
nand U14527 (N_14527,N_7290,N_6334);
nor U14528 (N_14528,N_7545,N_6162);
or U14529 (N_14529,N_8724,N_7113);
or U14530 (N_14530,N_6699,N_6294);
and U14531 (N_14531,N_8490,N_8567);
or U14532 (N_14532,N_8737,N_8530);
or U14533 (N_14533,N_7471,N_6820);
nand U14534 (N_14534,N_6564,N_8387);
nor U14535 (N_14535,N_5693,N_8146);
nor U14536 (N_14536,N_9786,N_6347);
and U14537 (N_14537,N_9995,N_6908);
nand U14538 (N_14538,N_6066,N_8648);
or U14539 (N_14539,N_8262,N_6430);
or U14540 (N_14540,N_8159,N_5346);
nor U14541 (N_14541,N_6796,N_6015);
or U14542 (N_14542,N_6411,N_5922);
nor U14543 (N_14543,N_8981,N_8697);
and U14544 (N_14544,N_7330,N_9662);
xnor U14545 (N_14545,N_9310,N_9171);
nand U14546 (N_14546,N_8893,N_9504);
or U14547 (N_14547,N_5257,N_5870);
nand U14548 (N_14548,N_7568,N_8919);
or U14549 (N_14549,N_9046,N_8529);
nand U14550 (N_14550,N_7485,N_6129);
nor U14551 (N_14551,N_9597,N_6063);
xor U14552 (N_14552,N_6289,N_8327);
nand U14553 (N_14553,N_8352,N_8560);
or U14554 (N_14554,N_9022,N_5401);
or U14555 (N_14555,N_5973,N_7808);
or U14556 (N_14556,N_9474,N_9985);
nor U14557 (N_14557,N_5037,N_8030);
nor U14558 (N_14558,N_7622,N_7363);
nand U14559 (N_14559,N_8301,N_7899);
nand U14560 (N_14560,N_9317,N_7190);
and U14561 (N_14561,N_8025,N_9268);
or U14562 (N_14562,N_6998,N_6322);
nor U14563 (N_14563,N_7506,N_7381);
nor U14564 (N_14564,N_9625,N_6849);
nor U14565 (N_14565,N_6301,N_6355);
nand U14566 (N_14566,N_5354,N_7855);
or U14567 (N_14567,N_5184,N_5566);
xnor U14568 (N_14568,N_6110,N_6469);
xor U14569 (N_14569,N_8510,N_6239);
and U14570 (N_14570,N_5960,N_9319);
nor U14571 (N_14571,N_9326,N_9819);
nand U14572 (N_14572,N_5511,N_8858);
or U14573 (N_14573,N_7210,N_7487);
nand U14574 (N_14574,N_7613,N_5127);
and U14575 (N_14575,N_6343,N_9962);
nor U14576 (N_14576,N_8094,N_6253);
nor U14577 (N_14577,N_9273,N_9702);
nor U14578 (N_14578,N_5804,N_8828);
or U14579 (N_14579,N_9900,N_6606);
and U14580 (N_14580,N_8846,N_8401);
and U14581 (N_14581,N_9414,N_9346);
xnor U14582 (N_14582,N_5596,N_8490);
nor U14583 (N_14583,N_5503,N_6577);
or U14584 (N_14584,N_6343,N_6744);
xnor U14585 (N_14585,N_6819,N_7186);
xnor U14586 (N_14586,N_9628,N_6962);
or U14587 (N_14587,N_7193,N_9936);
nor U14588 (N_14588,N_7368,N_8312);
and U14589 (N_14589,N_8945,N_7060);
xor U14590 (N_14590,N_5563,N_5118);
or U14591 (N_14591,N_8110,N_5839);
or U14592 (N_14592,N_8434,N_5776);
or U14593 (N_14593,N_6341,N_7060);
nand U14594 (N_14594,N_5491,N_6876);
and U14595 (N_14595,N_9750,N_5788);
nor U14596 (N_14596,N_9741,N_5587);
nand U14597 (N_14597,N_8257,N_5247);
or U14598 (N_14598,N_5508,N_9337);
nor U14599 (N_14599,N_8222,N_7843);
nor U14600 (N_14600,N_9642,N_9955);
xnor U14601 (N_14601,N_7392,N_9073);
nand U14602 (N_14602,N_8202,N_5553);
or U14603 (N_14603,N_5759,N_6179);
nand U14604 (N_14604,N_5286,N_9097);
and U14605 (N_14605,N_7021,N_5409);
nor U14606 (N_14606,N_9814,N_6994);
or U14607 (N_14607,N_8573,N_7428);
nor U14608 (N_14608,N_9336,N_9427);
nand U14609 (N_14609,N_6926,N_7393);
nor U14610 (N_14610,N_7737,N_5206);
xnor U14611 (N_14611,N_5028,N_6625);
and U14612 (N_14612,N_6765,N_5598);
xnor U14613 (N_14613,N_9250,N_9172);
nand U14614 (N_14614,N_8221,N_5153);
xor U14615 (N_14615,N_7281,N_9955);
and U14616 (N_14616,N_9136,N_6985);
nor U14617 (N_14617,N_9842,N_8038);
or U14618 (N_14618,N_6973,N_8110);
or U14619 (N_14619,N_6505,N_7794);
nor U14620 (N_14620,N_9359,N_9248);
nand U14621 (N_14621,N_9393,N_9280);
xnor U14622 (N_14622,N_5095,N_7676);
xnor U14623 (N_14623,N_9013,N_6424);
and U14624 (N_14624,N_5799,N_9148);
nand U14625 (N_14625,N_8515,N_9324);
xor U14626 (N_14626,N_8290,N_5840);
nand U14627 (N_14627,N_8473,N_7692);
or U14628 (N_14628,N_6954,N_5817);
or U14629 (N_14629,N_5632,N_8603);
or U14630 (N_14630,N_8906,N_9518);
nor U14631 (N_14631,N_7169,N_5488);
nand U14632 (N_14632,N_6239,N_7427);
nor U14633 (N_14633,N_6428,N_8932);
xor U14634 (N_14634,N_9818,N_5352);
nand U14635 (N_14635,N_7075,N_5723);
nor U14636 (N_14636,N_8447,N_9662);
or U14637 (N_14637,N_7148,N_7012);
or U14638 (N_14638,N_8809,N_8092);
or U14639 (N_14639,N_9162,N_9038);
or U14640 (N_14640,N_5331,N_9897);
nand U14641 (N_14641,N_7746,N_8417);
nand U14642 (N_14642,N_9139,N_8300);
nor U14643 (N_14643,N_6707,N_7367);
nor U14644 (N_14644,N_9959,N_7457);
nand U14645 (N_14645,N_5022,N_6936);
or U14646 (N_14646,N_9135,N_6121);
xor U14647 (N_14647,N_9025,N_9004);
or U14648 (N_14648,N_8914,N_8327);
nand U14649 (N_14649,N_5063,N_9071);
nor U14650 (N_14650,N_7381,N_6140);
nor U14651 (N_14651,N_6813,N_9726);
nor U14652 (N_14652,N_5580,N_5114);
xor U14653 (N_14653,N_6018,N_8507);
nand U14654 (N_14654,N_5704,N_9580);
nand U14655 (N_14655,N_9591,N_7957);
nor U14656 (N_14656,N_8475,N_9264);
or U14657 (N_14657,N_8503,N_6866);
and U14658 (N_14658,N_7984,N_9802);
and U14659 (N_14659,N_5170,N_9612);
nor U14660 (N_14660,N_8491,N_5408);
xnor U14661 (N_14661,N_8827,N_5925);
or U14662 (N_14662,N_7490,N_5221);
xor U14663 (N_14663,N_6696,N_5357);
nor U14664 (N_14664,N_8707,N_9974);
nor U14665 (N_14665,N_5226,N_8740);
xor U14666 (N_14666,N_7572,N_7776);
and U14667 (N_14667,N_7678,N_5767);
or U14668 (N_14668,N_6881,N_9523);
and U14669 (N_14669,N_7001,N_8381);
nand U14670 (N_14670,N_8639,N_6398);
or U14671 (N_14671,N_7181,N_6048);
or U14672 (N_14672,N_9108,N_9868);
xor U14673 (N_14673,N_5339,N_7409);
and U14674 (N_14674,N_5084,N_5209);
and U14675 (N_14675,N_8698,N_7943);
nand U14676 (N_14676,N_9257,N_9378);
or U14677 (N_14677,N_5670,N_8013);
xor U14678 (N_14678,N_6580,N_5664);
xor U14679 (N_14679,N_6556,N_9796);
nor U14680 (N_14680,N_5673,N_9734);
xnor U14681 (N_14681,N_7029,N_7608);
or U14682 (N_14682,N_9316,N_6486);
or U14683 (N_14683,N_9139,N_9633);
nand U14684 (N_14684,N_9377,N_6896);
nor U14685 (N_14685,N_5041,N_7295);
and U14686 (N_14686,N_8882,N_5867);
and U14687 (N_14687,N_9932,N_6234);
or U14688 (N_14688,N_6722,N_5015);
nand U14689 (N_14689,N_7546,N_7442);
or U14690 (N_14690,N_7520,N_9197);
or U14691 (N_14691,N_5218,N_9368);
nor U14692 (N_14692,N_9436,N_6107);
xnor U14693 (N_14693,N_6865,N_7466);
or U14694 (N_14694,N_9179,N_5799);
nand U14695 (N_14695,N_5127,N_6743);
nor U14696 (N_14696,N_9627,N_9109);
nor U14697 (N_14697,N_8203,N_8873);
nand U14698 (N_14698,N_7346,N_9624);
xnor U14699 (N_14699,N_5840,N_9186);
nand U14700 (N_14700,N_8466,N_9698);
xor U14701 (N_14701,N_9646,N_9820);
nor U14702 (N_14702,N_8672,N_7449);
and U14703 (N_14703,N_7472,N_7936);
and U14704 (N_14704,N_9924,N_9632);
or U14705 (N_14705,N_9948,N_6781);
xor U14706 (N_14706,N_9847,N_5754);
nand U14707 (N_14707,N_9265,N_6302);
nand U14708 (N_14708,N_8016,N_8304);
or U14709 (N_14709,N_8928,N_8556);
nor U14710 (N_14710,N_5047,N_8198);
xnor U14711 (N_14711,N_6528,N_7716);
nor U14712 (N_14712,N_6096,N_6594);
xnor U14713 (N_14713,N_7571,N_5776);
or U14714 (N_14714,N_8994,N_7483);
nand U14715 (N_14715,N_6307,N_7843);
and U14716 (N_14716,N_9023,N_7344);
and U14717 (N_14717,N_5949,N_7664);
xnor U14718 (N_14718,N_9108,N_8547);
nand U14719 (N_14719,N_7937,N_6314);
and U14720 (N_14720,N_5394,N_6438);
nand U14721 (N_14721,N_7972,N_9881);
nand U14722 (N_14722,N_5015,N_5475);
nor U14723 (N_14723,N_7402,N_5563);
nand U14724 (N_14724,N_9561,N_6123);
or U14725 (N_14725,N_8444,N_5328);
xnor U14726 (N_14726,N_8136,N_7823);
and U14727 (N_14727,N_5626,N_8290);
or U14728 (N_14728,N_9287,N_5928);
and U14729 (N_14729,N_9590,N_9492);
nor U14730 (N_14730,N_8769,N_6525);
nor U14731 (N_14731,N_8495,N_8456);
and U14732 (N_14732,N_5163,N_8964);
or U14733 (N_14733,N_5065,N_5898);
or U14734 (N_14734,N_7412,N_7575);
nand U14735 (N_14735,N_5958,N_8715);
nor U14736 (N_14736,N_7555,N_7327);
and U14737 (N_14737,N_5432,N_5628);
and U14738 (N_14738,N_6584,N_6144);
or U14739 (N_14739,N_5319,N_9940);
nor U14740 (N_14740,N_5092,N_5273);
and U14741 (N_14741,N_8125,N_8685);
and U14742 (N_14742,N_9795,N_6565);
nor U14743 (N_14743,N_6999,N_6680);
nand U14744 (N_14744,N_8994,N_8453);
nor U14745 (N_14745,N_7655,N_8615);
nor U14746 (N_14746,N_9028,N_5846);
nand U14747 (N_14747,N_7122,N_7064);
and U14748 (N_14748,N_7936,N_5935);
or U14749 (N_14749,N_8239,N_9726);
or U14750 (N_14750,N_7603,N_7579);
and U14751 (N_14751,N_7642,N_7111);
nand U14752 (N_14752,N_8504,N_7289);
and U14753 (N_14753,N_8207,N_6238);
xnor U14754 (N_14754,N_7079,N_6970);
and U14755 (N_14755,N_7120,N_9254);
and U14756 (N_14756,N_7330,N_8685);
or U14757 (N_14757,N_7077,N_5831);
or U14758 (N_14758,N_8580,N_5544);
xor U14759 (N_14759,N_8746,N_8736);
or U14760 (N_14760,N_6073,N_6266);
nor U14761 (N_14761,N_8203,N_6442);
nor U14762 (N_14762,N_8893,N_8854);
nor U14763 (N_14763,N_7671,N_8677);
or U14764 (N_14764,N_6435,N_8289);
nand U14765 (N_14765,N_6876,N_9615);
xnor U14766 (N_14766,N_6035,N_7253);
or U14767 (N_14767,N_6977,N_7009);
and U14768 (N_14768,N_6761,N_5469);
or U14769 (N_14769,N_9953,N_8269);
and U14770 (N_14770,N_9037,N_9557);
and U14771 (N_14771,N_8019,N_9699);
xnor U14772 (N_14772,N_7621,N_8449);
or U14773 (N_14773,N_7171,N_9785);
and U14774 (N_14774,N_6215,N_6528);
xnor U14775 (N_14775,N_5090,N_8829);
xnor U14776 (N_14776,N_9639,N_6944);
and U14777 (N_14777,N_9160,N_5001);
nand U14778 (N_14778,N_6164,N_7699);
or U14779 (N_14779,N_5346,N_5943);
nand U14780 (N_14780,N_8595,N_9864);
xnor U14781 (N_14781,N_8189,N_5503);
and U14782 (N_14782,N_7302,N_6269);
and U14783 (N_14783,N_9974,N_8197);
nand U14784 (N_14784,N_8881,N_8770);
xnor U14785 (N_14785,N_6233,N_9533);
or U14786 (N_14786,N_9585,N_5626);
or U14787 (N_14787,N_9282,N_9570);
and U14788 (N_14788,N_6590,N_8686);
nand U14789 (N_14789,N_8433,N_9202);
nor U14790 (N_14790,N_9836,N_9309);
nand U14791 (N_14791,N_8056,N_6424);
nor U14792 (N_14792,N_8190,N_9387);
nor U14793 (N_14793,N_9762,N_5061);
or U14794 (N_14794,N_9121,N_7759);
or U14795 (N_14795,N_6067,N_7781);
or U14796 (N_14796,N_9019,N_6937);
nand U14797 (N_14797,N_9965,N_5555);
xor U14798 (N_14798,N_9537,N_9674);
nor U14799 (N_14799,N_7117,N_5828);
nor U14800 (N_14800,N_9098,N_9124);
nor U14801 (N_14801,N_8298,N_9823);
xnor U14802 (N_14802,N_8168,N_5983);
nand U14803 (N_14803,N_7464,N_8157);
nand U14804 (N_14804,N_8868,N_5807);
nor U14805 (N_14805,N_9269,N_9772);
nor U14806 (N_14806,N_8564,N_8983);
or U14807 (N_14807,N_5689,N_7950);
nand U14808 (N_14808,N_6606,N_7782);
nand U14809 (N_14809,N_9042,N_5126);
nor U14810 (N_14810,N_9055,N_5606);
nor U14811 (N_14811,N_7910,N_7576);
nand U14812 (N_14812,N_5309,N_7368);
nand U14813 (N_14813,N_5614,N_5229);
and U14814 (N_14814,N_7078,N_7782);
nor U14815 (N_14815,N_5178,N_6046);
and U14816 (N_14816,N_8275,N_9579);
nand U14817 (N_14817,N_6603,N_6395);
or U14818 (N_14818,N_5064,N_9717);
or U14819 (N_14819,N_8565,N_6468);
nor U14820 (N_14820,N_6269,N_9939);
xnor U14821 (N_14821,N_6081,N_6943);
nand U14822 (N_14822,N_8137,N_6770);
xnor U14823 (N_14823,N_6256,N_6408);
nor U14824 (N_14824,N_6029,N_6679);
xor U14825 (N_14825,N_9887,N_8170);
nor U14826 (N_14826,N_7984,N_8486);
nand U14827 (N_14827,N_6193,N_8172);
and U14828 (N_14828,N_5874,N_9889);
nor U14829 (N_14829,N_8550,N_7908);
and U14830 (N_14830,N_8209,N_6702);
or U14831 (N_14831,N_6811,N_9560);
or U14832 (N_14832,N_8961,N_7422);
nand U14833 (N_14833,N_7369,N_5709);
xor U14834 (N_14834,N_5875,N_6990);
nand U14835 (N_14835,N_8961,N_8679);
nor U14836 (N_14836,N_5442,N_7857);
nor U14837 (N_14837,N_7038,N_6583);
and U14838 (N_14838,N_6146,N_8262);
nor U14839 (N_14839,N_5742,N_8241);
and U14840 (N_14840,N_9500,N_8417);
and U14841 (N_14841,N_9776,N_8049);
and U14842 (N_14842,N_9542,N_6663);
nand U14843 (N_14843,N_9045,N_7242);
xnor U14844 (N_14844,N_9177,N_7678);
or U14845 (N_14845,N_5954,N_7035);
xor U14846 (N_14846,N_9013,N_7591);
xor U14847 (N_14847,N_5938,N_5353);
nor U14848 (N_14848,N_8010,N_7731);
xor U14849 (N_14849,N_6147,N_9894);
and U14850 (N_14850,N_9092,N_9598);
nand U14851 (N_14851,N_8599,N_8707);
and U14852 (N_14852,N_9222,N_7199);
nand U14853 (N_14853,N_7483,N_7407);
or U14854 (N_14854,N_6867,N_5151);
or U14855 (N_14855,N_9701,N_7425);
nand U14856 (N_14856,N_9693,N_6931);
nor U14857 (N_14857,N_7972,N_9363);
or U14858 (N_14858,N_8459,N_5603);
xor U14859 (N_14859,N_7349,N_9101);
or U14860 (N_14860,N_5890,N_7553);
or U14861 (N_14861,N_5986,N_7935);
nand U14862 (N_14862,N_7917,N_6019);
nand U14863 (N_14863,N_7305,N_7129);
nand U14864 (N_14864,N_6458,N_7425);
nor U14865 (N_14865,N_6659,N_9293);
nor U14866 (N_14866,N_9266,N_5209);
xnor U14867 (N_14867,N_9689,N_7762);
xor U14868 (N_14868,N_7509,N_7206);
and U14869 (N_14869,N_6340,N_5342);
nand U14870 (N_14870,N_6254,N_5843);
nor U14871 (N_14871,N_9115,N_9895);
and U14872 (N_14872,N_8144,N_7216);
and U14873 (N_14873,N_9718,N_9594);
xor U14874 (N_14874,N_7424,N_8148);
and U14875 (N_14875,N_6708,N_7812);
nor U14876 (N_14876,N_5021,N_8183);
xor U14877 (N_14877,N_6549,N_6399);
nand U14878 (N_14878,N_7157,N_9563);
nand U14879 (N_14879,N_8754,N_7168);
or U14880 (N_14880,N_8636,N_5574);
or U14881 (N_14881,N_9341,N_6386);
nor U14882 (N_14882,N_8288,N_9577);
nand U14883 (N_14883,N_5508,N_8165);
nor U14884 (N_14884,N_9333,N_6543);
nand U14885 (N_14885,N_8447,N_8692);
nor U14886 (N_14886,N_8865,N_5779);
nor U14887 (N_14887,N_7542,N_5238);
xor U14888 (N_14888,N_7365,N_8623);
and U14889 (N_14889,N_6109,N_8680);
nor U14890 (N_14890,N_9607,N_5931);
xnor U14891 (N_14891,N_7486,N_9496);
nor U14892 (N_14892,N_5489,N_9225);
nor U14893 (N_14893,N_6700,N_8880);
and U14894 (N_14894,N_6727,N_8686);
nor U14895 (N_14895,N_7939,N_5376);
or U14896 (N_14896,N_9319,N_9700);
xor U14897 (N_14897,N_5907,N_9584);
nor U14898 (N_14898,N_6999,N_7660);
nor U14899 (N_14899,N_8950,N_7712);
or U14900 (N_14900,N_9242,N_8222);
nor U14901 (N_14901,N_7212,N_8435);
nor U14902 (N_14902,N_9641,N_8369);
xnor U14903 (N_14903,N_7353,N_8083);
nor U14904 (N_14904,N_9562,N_6270);
and U14905 (N_14905,N_7690,N_9361);
and U14906 (N_14906,N_5129,N_6217);
nand U14907 (N_14907,N_5583,N_5995);
nand U14908 (N_14908,N_8731,N_7727);
xor U14909 (N_14909,N_7640,N_9685);
or U14910 (N_14910,N_7292,N_6829);
or U14911 (N_14911,N_7887,N_7299);
nor U14912 (N_14912,N_5392,N_6575);
and U14913 (N_14913,N_7463,N_7150);
nor U14914 (N_14914,N_6279,N_7716);
xor U14915 (N_14915,N_8036,N_5516);
nand U14916 (N_14916,N_9668,N_6164);
and U14917 (N_14917,N_6279,N_8577);
or U14918 (N_14918,N_5522,N_8488);
nand U14919 (N_14919,N_7431,N_6601);
nor U14920 (N_14920,N_8193,N_9155);
xor U14921 (N_14921,N_9924,N_7672);
and U14922 (N_14922,N_5231,N_9850);
xnor U14923 (N_14923,N_7683,N_9814);
xnor U14924 (N_14924,N_6961,N_5841);
or U14925 (N_14925,N_5349,N_6784);
or U14926 (N_14926,N_8170,N_7391);
nor U14927 (N_14927,N_9736,N_7250);
nand U14928 (N_14928,N_7502,N_6535);
nand U14929 (N_14929,N_9108,N_5824);
and U14930 (N_14930,N_5115,N_9560);
and U14931 (N_14931,N_7101,N_5411);
nand U14932 (N_14932,N_7684,N_8522);
nand U14933 (N_14933,N_6181,N_5823);
nor U14934 (N_14934,N_5106,N_8288);
nor U14935 (N_14935,N_8409,N_7284);
or U14936 (N_14936,N_8030,N_6978);
nor U14937 (N_14937,N_7134,N_7692);
nand U14938 (N_14938,N_8705,N_6835);
or U14939 (N_14939,N_6688,N_6390);
or U14940 (N_14940,N_9129,N_8230);
or U14941 (N_14941,N_5931,N_7065);
or U14942 (N_14942,N_7203,N_7493);
nand U14943 (N_14943,N_6832,N_8792);
nor U14944 (N_14944,N_6502,N_9691);
nand U14945 (N_14945,N_6359,N_6753);
nor U14946 (N_14946,N_7971,N_9600);
or U14947 (N_14947,N_7834,N_8906);
or U14948 (N_14948,N_9526,N_8819);
and U14949 (N_14949,N_5314,N_5418);
xor U14950 (N_14950,N_8155,N_7108);
nand U14951 (N_14951,N_9750,N_9085);
nor U14952 (N_14952,N_6770,N_6476);
nand U14953 (N_14953,N_7428,N_5585);
xor U14954 (N_14954,N_7712,N_8067);
nor U14955 (N_14955,N_9845,N_5248);
nand U14956 (N_14956,N_8115,N_7676);
nand U14957 (N_14957,N_7001,N_5191);
or U14958 (N_14958,N_8195,N_9218);
and U14959 (N_14959,N_7492,N_8868);
and U14960 (N_14960,N_8642,N_6510);
and U14961 (N_14961,N_7565,N_8359);
nand U14962 (N_14962,N_6984,N_6718);
or U14963 (N_14963,N_8165,N_5883);
nand U14964 (N_14964,N_5519,N_6576);
and U14965 (N_14965,N_5024,N_6940);
nand U14966 (N_14966,N_5659,N_7482);
xnor U14967 (N_14967,N_7885,N_8612);
or U14968 (N_14968,N_7179,N_7627);
or U14969 (N_14969,N_7902,N_8814);
or U14970 (N_14970,N_5840,N_6336);
xnor U14971 (N_14971,N_7402,N_8947);
or U14972 (N_14972,N_5955,N_8960);
or U14973 (N_14973,N_6211,N_8210);
nand U14974 (N_14974,N_9638,N_5274);
and U14975 (N_14975,N_6732,N_6099);
nand U14976 (N_14976,N_7614,N_8879);
and U14977 (N_14977,N_9293,N_7347);
nor U14978 (N_14978,N_5477,N_6785);
nand U14979 (N_14979,N_9566,N_5377);
or U14980 (N_14980,N_8820,N_8691);
xnor U14981 (N_14981,N_8951,N_8073);
nand U14982 (N_14982,N_8278,N_9946);
and U14983 (N_14983,N_5155,N_5782);
nand U14984 (N_14984,N_5613,N_6225);
and U14985 (N_14985,N_8411,N_7392);
xor U14986 (N_14986,N_8115,N_9370);
xor U14987 (N_14987,N_5473,N_6763);
nor U14988 (N_14988,N_8311,N_6181);
xor U14989 (N_14989,N_5677,N_8298);
or U14990 (N_14990,N_6287,N_7116);
xnor U14991 (N_14991,N_6487,N_5249);
nor U14992 (N_14992,N_7736,N_9821);
or U14993 (N_14993,N_8037,N_5834);
xnor U14994 (N_14994,N_8955,N_9219);
and U14995 (N_14995,N_9671,N_8247);
nand U14996 (N_14996,N_6342,N_7737);
and U14997 (N_14997,N_8662,N_5284);
and U14998 (N_14998,N_7665,N_9345);
xnor U14999 (N_14999,N_7791,N_5280);
xnor U15000 (N_15000,N_14793,N_13808);
nand U15001 (N_15001,N_13962,N_12817);
nor U15002 (N_15002,N_14145,N_14702);
xnor U15003 (N_15003,N_10654,N_14634);
or U15004 (N_15004,N_12568,N_11830);
nand U15005 (N_15005,N_13426,N_10082);
nor U15006 (N_15006,N_14823,N_12443);
nor U15007 (N_15007,N_13671,N_10104);
xor U15008 (N_15008,N_10608,N_11540);
nand U15009 (N_15009,N_14657,N_13550);
xnor U15010 (N_15010,N_11730,N_13476);
nor U15011 (N_15011,N_14952,N_10070);
or U15012 (N_15012,N_10190,N_13509);
nor U15013 (N_15013,N_11538,N_13387);
or U15014 (N_15014,N_10626,N_13713);
nor U15015 (N_15015,N_10307,N_11990);
nand U15016 (N_15016,N_10250,N_10246);
and U15017 (N_15017,N_11073,N_14306);
xor U15018 (N_15018,N_13002,N_14625);
and U15019 (N_15019,N_12695,N_13371);
xnor U15020 (N_15020,N_14051,N_11769);
nand U15021 (N_15021,N_11052,N_13822);
xor U15022 (N_15022,N_14640,N_12221);
and U15023 (N_15023,N_12234,N_10803);
nand U15024 (N_15024,N_12828,N_10516);
or U15025 (N_15025,N_13538,N_12654);
xnor U15026 (N_15026,N_14860,N_11718);
nor U15027 (N_15027,N_13493,N_13996);
nor U15028 (N_15028,N_10646,N_12414);
or U15029 (N_15029,N_12025,N_11989);
nor U15030 (N_15030,N_10549,N_13866);
and U15031 (N_15031,N_13777,N_14023);
nand U15032 (N_15032,N_14915,N_12115);
xor U15033 (N_15033,N_13574,N_10942);
nor U15034 (N_15034,N_12750,N_14307);
nor U15035 (N_15035,N_11648,N_10097);
and U15036 (N_15036,N_12330,N_12906);
nand U15037 (N_15037,N_10592,N_12882);
nand U15038 (N_15038,N_13174,N_10181);
nor U15039 (N_15039,N_12953,N_10829);
nand U15040 (N_15040,N_10796,N_11758);
and U15041 (N_15041,N_14311,N_11124);
xor U15042 (N_15042,N_10333,N_10691);
or U15043 (N_15043,N_12966,N_10088);
nor U15044 (N_15044,N_13389,N_13961);
xor U15045 (N_15045,N_10438,N_14862);
nand U15046 (N_15046,N_14650,N_14365);
nand U15047 (N_15047,N_13297,N_11654);
or U15048 (N_15048,N_10739,N_14120);
and U15049 (N_15049,N_14973,N_11234);
or U15050 (N_15050,N_14598,N_12451);
xnor U15051 (N_15051,N_13906,N_12758);
or U15052 (N_15052,N_13074,N_14845);
xor U15053 (N_15053,N_11995,N_14799);
or U15054 (N_15054,N_12297,N_10192);
nor U15055 (N_15055,N_10450,N_11745);
nor U15056 (N_15056,N_10282,N_13212);
nor U15057 (N_15057,N_13510,N_11802);
or U15058 (N_15058,N_11222,N_14909);
or U15059 (N_15059,N_11529,N_10969);
xor U15060 (N_15060,N_12202,N_14758);
and U15061 (N_15061,N_12674,N_12170);
xor U15062 (N_15062,N_11587,N_14322);
and U15063 (N_15063,N_14810,N_14515);
and U15064 (N_15064,N_13825,N_11897);
xor U15065 (N_15065,N_12641,N_12062);
and U15066 (N_15066,N_10934,N_10576);
or U15067 (N_15067,N_14813,N_10189);
or U15068 (N_15068,N_13065,N_10021);
and U15069 (N_15069,N_11108,N_14500);
or U15070 (N_15070,N_12023,N_13467);
nand U15071 (N_15071,N_13666,N_14644);
nand U15072 (N_15072,N_13726,N_10947);
and U15073 (N_15073,N_11095,N_11454);
or U15074 (N_15074,N_14054,N_14140);
or U15075 (N_15075,N_12970,N_12343);
nand U15076 (N_15076,N_12305,N_14774);
or U15077 (N_15077,N_12603,N_11221);
xor U15078 (N_15078,N_14544,N_11186);
nand U15079 (N_15079,N_12217,N_14609);
nand U15080 (N_15080,N_12254,N_13632);
xor U15081 (N_15081,N_14525,N_14804);
nor U15082 (N_15082,N_13531,N_12005);
nor U15083 (N_15083,N_11231,N_12892);
nor U15084 (N_15084,N_14847,N_10052);
or U15085 (N_15085,N_14729,N_10918);
and U15086 (N_15086,N_10083,N_12047);
and U15087 (N_15087,N_13228,N_11739);
and U15088 (N_15088,N_14377,N_12309);
xor U15089 (N_15089,N_13670,N_14773);
xnor U15090 (N_15090,N_14997,N_11023);
or U15091 (N_15091,N_13357,N_12308);
xnor U15092 (N_15092,N_11592,N_12404);
and U15093 (N_15093,N_14250,N_12904);
nand U15094 (N_15094,N_10092,N_12168);
nand U15095 (N_15095,N_14911,N_10962);
and U15096 (N_15096,N_14331,N_10213);
xor U15097 (N_15097,N_13169,N_14627);
nand U15098 (N_15098,N_11494,N_10504);
or U15099 (N_15099,N_10440,N_13977);
and U15100 (N_15100,N_11384,N_11584);
or U15101 (N_15101,N_14652,N_11316);
and U15102 (N_15102,N_11539,N_14205);
and U15103 (N_15103,N_14792,N_11203);
or U15104 (N_15104,N_10783,N_11344);
or U15105 (N_15105,N_12755,N_11062);
xnor U15106 (N_15106,N_13117,N_13934);
nand U15107 (N_15107,N_12689,N_10114);
and U15108 (N_15108,N_11328,N_12619);
or U15109 (N_15109,N_10804,N_11649);
and U15110 (N_15110,N_10764,N_14849);
xnor U15111 (N_15111,N_11544,N_13741);
xor U15112 (N_15112,N_14111,N_11345);
or U15113 (N_15113,N_13751,N_13583);
xor U15114 (N_15114,N_10583,N_13573);
nand U15115 (N_15115,N_11775,N_10343);
or U15116 (N_15116,N_10749,N_13784);
and U15117 (N_15117,N_12307,N_14299);
and U15118 (N_15118,N_10567,N_10472);
xor U15119 (N_15119,N_12652,N_12719);
and U15120 (N_15120,N_11304,N_13756);
xor U15121 (N_15121,N_12395,N_13193);
and U15122 (N_15122,N_13162,N_10732);
nand U15123 (N_15123,N_13805,N_10179);
nor U15124 (N_15124,N_12699,N_13941);
or U15125 (N_15125,N_10142,N_13149);
nor U15126 (N_15126,N_13986,N_11597);
nor U15127 (N_15127,N_10538,N_13708);
or U15128 (N_15128,N_11247,N_14421);
and U15129 (N_15129,N_14876,N_13515);
nor U15130 (N_15130,N_13705,N_10356);
or U15131 (N_15131,N_13436,N_12713);
or U15132 (N_15132,N_13855,N_14242);
nor U15133 (N_15133,N_14541,N_10768);
nand U15134 (N_15134,N_12140,N_10134);
nor U15135 (N_15135,N_10988,N_14057);
or U15136 (N_15136,N_10030,N_12160);
nor U15137 (N_15137,N_12176,N_12809);
xnor U15138 (N_15138,N_11303,N_13305);
nand U15139 (N_15139,N_14933,N_12955);
xor U15140 (N_15140,N_11914,N_10841);
xor U15141 (N_15141,N_14654,N_12665);
nor U15142 (N_15142,N_11781,N_13852);
xnor U15143 (N_15143,N_12725,N_12219);
and U15144 (N_15144,N_13195,N_10191);
or U15145 (N_15145,N_13706,N_12857);
or U15146 (N_15146,N_13703,N_13564);
or U15147 (N_15147,N_11562,N_10766);
nor U15148 (N_15148,N_14536,N_10446);
xor U15149 (N_15149,N_12071,N_14375);
and U15150 (N_15150,N_11050,N_13469);
or U15151 (N_15151,N_13891,N_12651);
nor U15152 (N_15152,N_10387,N_14759);
nand U15153 (N_15153,N_13124,N_13685);
nand U15154 (N_15154,N_11958,N_12960);
nand U15155 (N_15155,N_13710,N_14519);
xnor U15156 (N_15156,N_11090,N_10582);
nor U15157 (N_15157,N_12123,N_11284);
and U15158 (N_15158,N_14919,N_11139);
nor U15159 (N_15159,N_14717,N_12776);
nand U15160 (N_15160,N_12905,N_14342);
and U15161 (N_15161,N_10500,N_14868);
nor U15162 (N_15162,N_11188,N_13998);
and U15163 (N_15163,N_11148,N_11717);
nand U15164 (N_15164,N_10844,N_10615);
xnor U15165 (N_15165,N_11294,N_13353);
nand U15166 (N_15166,N_11438,N_12535);
nor U15167 (N_15167,N_10017,N_14070);
and U15168 (N_15168,N_13965,N_11513);
xnor U15169 (N_15169,N_12945,N_13115);
nor U15170 (N_15170,N_12749,N_14583);
xnor U15171 (N_15171,N_10166,N_11978);
nor U15172 (N_15172,N_12473,N_10106);
nand U15173 (N_15173,N_12702,N_13092);
xnor U15174 (N_15174,N_14581,N_14679);
nor U15175 (N_15175,N_12060,N_12035);
or U15176 (N_15176,N_10895,N_13270);
and U15177 (N_15177,N_14763,N_10743);
xnor U15178 (N_15178,N_11078,N_10912);
nor U15179 (N_15179,N_13407,N_12597);
and U15180 (N_15180,N_13660,N_14402);
and U15181 (N_15181,N_11939,N_12396);
or U15182 (N_15182,N_11907,N_12764);
or U15183 (N_15183,N_11827,N_13975);
or U15184 (N_15184,N_12293,N_14485);
xnor U15185 (N_15185,N_14942,N_12072);
and U15186 (N_15186,N_12363,N_14084);
xnor U15187 (N_15187,N_14188,N_10596);
xnor U15188 (N_15188,N_14434,N_11474);
nand U15189 (N_15189,N_14113,N_11690);
xor U15190 (N_15190,N_13448,N_11038);
xor U15191 (N_15191,N_12190,N_11554);
xnor U15192 (N_15192,N_11032,N_13361);
or U15193 (N_15193,N_12406,N_10720);
xnor U15194 (N_15194,N_14556,N_11674);
nand U15195 (N_15195,N_14943,N_13529);
nor U15196 (N_15196,N_14596,N_14280);
nand U15197 (N_15197,N_10065,N_10311);
or U15198 (N_15198,N_10394,N_12034);
nand U15199 (N_15199,N_11468,N_14286);
xor U15200 (N_15200,N_11744,N_11751);
nand U15201 (N_15201,N_14570,N_12681);
and U15202 (N_15202,N_13138,N_13443);
nor U15203 (N_15203,N_12258,N_10421);
nor U15204 (N_15204,N_13046,N_11133);
and U15205 (N_15205,N_13060,N_11624);
nor U15206 (N_15206,N_14341,N_12638);
nor U15207 (N_15207,N_12173,N_13902);
nand U15208 (N_15208,N_13017,N_10231);
nand U15209 (N_15209,N_10744,N_13834);
or U15210 (N_15210,N_10442,N_12562);
xor U15211 (N_15211,N_10610,N_10825);
and U15212 (N_15212,N_11224,N_10284);
xnor U15213 (N_15213,N_11464,N_13245);
nor U15214 (N_15214,N_10584,N_14410);
xor U15215 (N_15215,N_11973,N_14474);
nand U15216 (N_15216,N_14103,N_13932);
or U15217 (N_15217,N_12716,N_14175);
nor U15218 (N_15218,N_12565,N_12679);
or U15219 (N_15219,N_14545,N_10229);
nand U15220 (N_15220,N_14337,N_13480);
or U15221 (N_15221,N_12383,N_10581);
or U15222 (N_15222,N_12605,N_14394);
xnor U15223 (N_15223,N_10882,N_14529);
nor U15224 (N_15224,N_11576,N_13328);
xnor U15225 (N_15225,N_13376,N_12497);
or U15226 (N_15226,N_11706,N_10754);
nor U15227 (N_15227,N_11503,N_11080);
or U15228 (N_15228,N_13455,N_12030);
nor U15229 (N_15229,N_13616,N_11312);
and U15230 (N_15230,N_12420,N_10884);
xnor U15231 (N_15231,N_11952,N_13942);
nand U15232 (N_15232,N_10420,N_11593);
or U15233 (N_15233,N_11496,N_13661);
nor U15234 (N_15234,N_14202,N_10270);
nor U15235 (N_15235,N_13796,N_12762);
xnor U15236 (N_15236,N_14802,N_13129);
nor U15237 (N_15237,N_14964,N_12526);
nor U15238 (N_15238,N_10028,N_12121);
xor U15239 (N_15239,N_10120,N_13182);
xor U15240 (N_15240,N_11024,N_13680);
and U15241 (N_15241,N_13653,N_11832);
nand U15242 (N_15242,N_12840,N_13696);
nand U15243 (N_15243,N_13076,N_12126);
and U15244 (N_15244,N_14451,N_13641);
xor U15245 (N_15245,N_12718,N_10636);
or U15246 (N_15246,N_11877,N_12663);
xnor U15247 (N_15247,N_13240,N_10780);
nand U15248 (N_15248,N_10366,N_12317);
or U15249 (N_15249,N_10422,N_13552);
nor U15250 (N_15250,N_13134,N_11182);
nor U15251 (N_15251,N_13350,N_11013);
nand U15252 (N_15252,N_13207,N_13080);
nor U15253 (N_15253,N_14159,N_14446);
and U15254 (N_15254,N_12038,N_13056);
and U15255 (N_15255,N_10319,N_12261);
nor U15256 (N_15256,N_14607,N_10041);
nor U15257 (N_15257,N_14201,N_10367);
xor U15258 (N_15258,N_11015,N_12073);
nor U15259 (N_15259,N_12238,N_13179);
nand U15260 (N_15260,N_10999,N_13893);
nor U15261 (N_15261,N_12639,N_14630);
nand U15262 (N_15262,N_10268,N_14495);
and U15263 (N_15263,N_11109,N_10223);
or U15264 (N_15264,N_10908,N_13012);
nand U15265 (N_15265,N_13917,N_13927);
nor U15266 (N_15266,N_11026,N_11789);
and U15267 (N_15267,N_12417,N_11381);
and U15268 (N_15268,N_13023,N_12130);
nor U15269 (N_15269,N_13412,N_14803);
nor U15270 (N_15270,N_12901,N_11376);
and U15271 (N_15271,N_11356,N_11266);
and U15272 (N_15272,N_12606,N_13268);
nand U15273 (N_15273,N_10435,N_13444);
or U15274 (N_15274,N_14819,N_10337);
nand U15275 (N_15275,N_11515,N_12582);
and U15276 (N_15276,N_11166,N_14769);
or U15277 (N_15277,N_10023,N_10630);
nand U15278 (N_15278,N_12649,N_11664);
nor U15279 (N_15279,N_14701,N_10119);
xor U15280 (N_15280,N_13229,N_11364);
nand U15281 (N_15281,N_11811,N_13449);
and U15282 (N_15282,N_10465,N_10045);
and U15283 (N_15283,N_10534,N_10972);
or U15284 (N_15284,N_12339,N_12978);
nand U15285 (N_15285,N_13931,N_11840);
or U15286 (N_15286,N_11588,N_10130);
nor U15287 (N_15287,N_10699,N_10124);
nand U15288 (N_15288,N_12647,N_13020);
nand U15289 (N_15289,N_10009,N_10980);
xnor U15290 (N_15290,N_11887,N_13924);
or U15291 (N_15291,N_10839,N_11969);
xor U15292 (N_15292,N_12493,N_11324);
xnor U15293 (N_15293,N_11608,N_14852);
nand U15294 (N_15294,N_10715,N_13140);
xnor U15295 (N_15295,N_13596,N_12561);
nand U15296 (N_15296,N_14971,N_12943);
nand U15297 (N_15297,N_11457,N_10556);
nand U15298 (N_15298,N_10171,N_14703);
or U15299 (N_15299,N_13522,N_13085);
xor U15300 (N_15300,N_13404,N_14014);
xnor U15301 (N_15301,N_11964,N_12502);
nor U15302 (N_15302,N_14994,N_10943);
nand U15303 (N_15303,N_14653,N_13209);
and U15304 (N_15304,N_11020,N_13275);
or U15305 (N_15305,N_14199,N_13463);
or U15306 (N_15306,N_10087,N_11350);
nand U15307 (N_15307,N_11697,N_12657);
nor U15308 (N_15308,N_14624,N_12494);
nand U15309 (N_15309,N_10545,N_14472);
and U15310 (N_15310,N_13241,N_14207);
and U15311 (N_15311,N_11253,N_13997);
nand U15312 (N_15312,N_10671,N_14872);
nor U15313 (N_15313,N_11453,N_12885);
xor U15314 (N_15314,N_11705,N_13086);
or U15315 (N_15315,N_13004,N_12010);
xor U15316 (N_15316,N_10536,N_10154);
nor U15317 (N_15317,N_12212,N_13516);
and U15318 (N_15318,N_13694,N_13049);
or U15319 (N_15319,N_10898,N_11152);
xnor U15320 (N_15320,N_12893,N_14887);
or U15321 (N_15321,N_10386,N_10704);
and U15322 (N_15322,N_14327,N_12350);
xnor U15323 (N_15323,N_12430,N_10676);
nor U15324 (N_15324,N_11534,N_10930);
and U15325 (N_15325,N_11000,N_13249);
and U15326 (N_15326,N_12867,N_14212);
and U15327 (N_15327,N_10115,N_10248);
nand U15328 (N_15328,N_10016,N_13576);
or U15329 (N_15329,N_10903,N_13611);
nor U15330 (N_15330,N_14597,N_14222);
and U15331 (N_15331,N_11202,N_11027);
nand U15332 (N_15332,N_11146,N_13344);
nor U15333 (N_15333,N_10721,N_14439);
and U15334 (N_15334,N_13257,N_13373);
xnor U15335 (N_15335,N_13592,N_13078);
nand U15336 (N_15336,N_11699,N_14420);
xnor U15337 (N_15337,N_10860,N_13453);
nor U15338 (N_15338,N_12042,N_12491);
and U15339 (N_15339,N_10728,N_14240);
nor U15340 (N_15340,N_13155,N_12045);
xor U15341 (N_15341,N_13544,N_10327);
xnor U15342 (N_15342,N_10354,N_14494);
and U15343 (N_15343,N_14007,N_12723);
and U15344 (N_15344,N_11719,N_12564);
or U15345 (N_15345,N_14459,N_10352);
and U15346 (N_15346,N_13987,N_11693);
nor U15347 (N_15347,N_14906,N_10886);
nand U15348 (N_15348,N_14429,N_13075);
nor U15349 (N_15349,N_12822,N_13900);
and U15350 (N_15350,N_12250,N_11683);
nand U15351 (N_15351,N_12896,N_14505);
and U15352 (N_15352,N_10819,N_11472);
or U15353 (N_15353,N_11710,N_11550);
and U15354 (N_15354,N_14809,N_14149);
xor U15355 (N_15355,N_14038,N_12472);
nand U15356 (N_15356,N_10278,N_13466);
xnor U15357 (N_15357,N_10089,N_12359);
and U15358 (N_15358,N_13401,N_11486);
nor U15359 (N_15359,N_10836,N_10123);
xnor U15360 (N_15360,N_13461,N_11113);
and U15361 (N_15361,N_10194,N_13141);
nand U15362 (N_15362,N_14540,N_12696);
or U15363 (N_15363,N_12440,N_11640);
nor U15364 (N_15364,N_13517,N_10346);
and U15365 (N_15365,N_12986,N_13069);
and U15366 (N_15366,N_10981,N_13771);
xnor U15367 (N_15367,N_11422,N_12411);
or U15368 (N_15368,N_13470,N_14508);
or U15369 (N_15369,N_10176,N_14699);
and U15370 (N_15370,N_10531,N_13041);
xnor U15371 (N_15371,N_13722,N_14696);
nor U15372 (N_15372,N_14521,N_10987);
nand U15373 (N_15373,N_13501,N_11319);
or U15374 (N_15374,N_10588,N_12599);
nor U15375 (N_15375,N_13752,N_11196);
nor U15376 (N_15376,N_14243,N_14733);
xnor U15377 (N_15377,N_14245,N_11059);
and U15378 (N_15378,N_13603,N_11728);
and U15379 (N_15379,N_12643,N_13951);
nor U15380 (N_15380,N_14339,N_12024);
or U15381 (N_15381,N_12530,N_12629);
nor U15382 (N_15382,N_11003,N_11365);
or U15383 (N_15383,N_13945,N_14176);
nor U15384 (N_15384,N_11371,N_13848);
nand U15385 (N_15385,N_11835,N_14718);
nor U15386 (N_15386,N_13619,N_14692);
nor U15387 (N_15387,N_14066,N_13799);
nor U15388 (N_15388,N_13079,N_10936);
nand U15389 (N_15389,N_12028,N_13173);
and U15390 (N_15390,N_13359,N_10568);
or U15391 (N_15391,N_13486,N_10497);
nor U15392 (N_15392,N_12251,N_10416);
nand U15393 (N_15393,N_12578,N_13905);
or U15394 (N_15394,N_14514,N_11843);
or U15395 (N_15395,N_14266,N_13219);
and U15396 (N_15396,N_14655,N_13928);
and U15397 (N_15397,N_10694,N_10058);
nor U15398 (N_15398,N_10081,N_12720);
or U15399 (N_15399,N_13397,N_13309);
and U15400 (N_15400,N_10632,N_13783);
and U15401 (N_15401,N_12656,N_10785);
xnor U15402 (N_15402,N_14620,N_14928);
and U15403 (N_15403,N_12490,N_14835);
nand U15404 (N_15404,N_13302,N_12065);
nand U15405 (N_15405,N_13456,N_12925);
xnor U15406 (N_15406,N_10855,N_14927);
nor U15407 (N_15407,N_13205,N_12968);
nor U15408 (N_15408,N_12400,N_11339);
and U15409 (N_15409,N_13283,N_14021);
nand U15410 (N_15410,N_14381,N_10380);
nor U15411 (N_15411,N_14831,N_13781);
and U15412 (N_15412,N_13579,N_14641);
or U15413 (N_15413,N_12505,N_11732);
or U15414 (N_15414,N_14164,N_11042);
nand U15415 (N_15415,N_14391,N_10910);
xnor U15416 (N_15416,N_11582,N_13658);
and U15417 (N_15417,N_10653,N_14189);
or U15418 (N_15418,N_14848,N_14916);
nand U15419 (N_15419,N_11612,N_12391);
xor U15420 (N_15420,N_14601,N_12516);
or U15421 (N_15421,N_13643,N_12120);
nor U15422 (N_15422,N_13686,N_13250);
or U15423 (N_15423,N_12185,N_13790);
or U15424 (N_15424,N_13018,N_10672);
xor U15425 (N_15425,N_11197,N_11533);
nor U15426 (N_15426,N_10220,N_14400);
xnor U15427 (N_15427,N_12742,N_10564);
nand U15428 (N_15428,N_10160,N_14468);
nand U15429 (N_15429,N_11101,N_10414);
or U15430 (N_15430,N_14816,N_14470);
nand U15431 (N_15431,N_14343,N_14840);
nor U15432 (N_15432,N_13154,N_14059);
or U15433 (N_15433,N_12832,N_14213);
or U15434 (N_15434,N_13868,N_10614);
and U15435 (N_15435,N_10431,N_11401);
and U15436 (N_15436,N_11954,N_10187);
and U15437 (N_15437,N_14036,N_11317);
or U15438 (N_15438,N_12640,N_10024);
nor U15439 (N_15439,N_14844,N_13743);
xor U15440 (N_15440,N_14304,N_12813);
nor U15441 (N_15441,N_14636,N_10528);
nand U15442 (N_15442,N_10227,N_13044);
xor U15443 (N_15443,N_11797,N_12004);
or U15444 (N_15444,N_10827,N_12177);
and U15445 (N_15445,N_11111,N_14052);
nor U15446 (N_15446,N_14384,N_11543);
xnor U15447 (N_15447,N_13340,N_13881);
and U15448 (N_15448,N_13070,N_12553);
xor U15449 (N_15449,N_11030,N_11721);
or U15450 (N_15450,N_11006,N_14531);
or U15451 (N_15451,N_14035,N_11418);
nor U15452 (N_15452,N_14364,N_11063);
or U15453 (N_15453,N_14839,N_12402);
or U15454 (N_15454,N_10896,N_12866);
and U15455 (N_15455,N_14160,N_11210);
or U15456 (N_15456,N_13859,N_11707);
xnor U15457 (N_15457,N_12392,N_12093);
nor U15458 (N_15458,N_12436,N_11971);
or U15459 (N_15459,N_14842,N_10403);
xnor U15460 (N_15460,N_13352,N_13896);
nor U15461 (N_15461,N_14762,N_14885);
and U15462 (N_15462,N_13667,N_10383);
nor U15463 (N_15463,N_11738,N_11581);
nand U15464 (N_15464,N_12596,N_11741);
or U15465 (N_15465,N_10503,N_14288);
or U15466 (N_15466,N_13939,N_12087);
nand U15467 (N_15467,N_11591,N_11277);
xor U15468 (N_15468,N_14542,N_11564);
or U15469 (N_15469,N_14912,N_10008);
nor U15470 (N_15470,N_14133,N_11734);
xnor U15471 (N_15471,N_10480,N_11089);
xor U15472 (N_15472,N_13161,N_14656);
xnor U15473 (N_15473,N_12407,N_14206);
and U15474 (N_15474,N_11848,N_14918);
or U15475 (N_15475,N_12364,N_12495);
nand U15476 (N_15476,N_12801,N_13102);
xnor U15477 (N_15477,N_11268,N_10973);
nor U15478 (N_15478,N_12541,N_14574);
and U15479 (N_15479,N_10648,N_11439);
or U15480 (N_15480,N_13640,N_14333);
xor U15481 (N_15481,N_12448,N_12791);
nand U15482 (N_15482,N_10817,N_10360);
and U15483 (N_15483,N_14877,N_14223);
xor U15484 (N_15484,N_14440,N_11763);
and U15485 (N_15485,N_14075,N_12031);
nand U15486 (N_15486,N_14349,N_12029);
nand U15487 (N_15487,N_13160,N_14516);
xnor U15488 (N_15488,N_13291,N_10113);
xnor U15489 (N_15489,N_11526,N_10575);
nor U15490 (N_15490,N_14368,N_13024);
or U15491 (N_15491,N_10237,N_13804);
nor U15492 (N_15492,N_13903,N_13739);
and U15493 (N_15493,N_10883,N_10161);
xnor U15494 (N_15494,N_10390,N_13499);
xnor U15495 (N_15495,N_13880,N_11735);
nor U15496 (N_15496,N_10655,N_13370);
xor U15497 (N_15497,N_14547,N_13142);
or U15498 (N_15498,N_12159,N_10997);
and U15499 (N_15499,N_14504,N_10384);
xor U15500 (N_15500,N_14261,N_12733);
and U15501 (N_15501,N_12819,N_13465);
or U15502 (N_15502,N_10927,N_10055);
nor U15503 (N_15503,N_14881,N_14215);
or U15504 (N_15504,N_14354,N_10490);
or U15505 (N_15505,N_12456,N_11168);
xor U15506 (N_15506,N_10527,N_11369);
and U15507 (N_15507,N_11869,N_11191);
nor U15508 (N_15508,N_12683,N_10953);
and U15509 (N_15509,N_14191,N_12325);
or U15510 (N_15510,N_10741,N_13675);
or U15511 (N_15511,N_11747,N_10598);
or U15512 (N_15512,N_10759,N_10322);
xnor U15513 (N_15513,N_13622,N_10251);
nand U15514 (N_15514,N_14851,N_13243);
nand U15515 (N_15515,N_13541,N_12903);
nor U15516 (N_15516,N_14479,N_12486);
xor U15517 (N_15517,N_10795,N_12790);
nor U15518 (N_15518,N_10595,N_11002);
nand U15519 (N_15519,N_11514,N_13187);
xor U15520 (N_15520,N_10714,N_11670);
xnor U15521 (N_15521,N_13491,N_12838);
nor U15522 (N_15522,N_11267,N_10977);
and U15523 (N_15523,N_10210,N_13633);
xor U15524 (N_15524,N_12974,N_13873);
or U15525 (N_15525,N_11308,N_12015);
or U15526 (N_15526,N_11983,N_10924);
and U15527 (N_15527,N_12447,N_12598);
and U15528 (N_15528,N_14501,N_11643);
xnor U15529 (N_15529,N_12610,N_14005);
and U15530 (N_15530,N_14962,N_14659);
nor U15531 (N_15531,N_13264,N_12153);
xnor U15532 (N_15532,N_10578,N_14555);
nand U15533 (N_15533,N_14317,N_10286);
and U15534 (N_15534,N_11207,N_14246);
or U15535 (N_15535,N_11571,N_11780);
nor U15536 (N_15536,N_12253,N_13801);
xor U15537 (N_15537,N_13894,N_11658);
nand U15538 (N_15538,N_12275,N_10443);
nor U15539 (N_15539,N_11449,N_11784);
nor U15540 (N_15540,N_14678,N_12055);
or U15541 (N_15541,N_10523,N_12315);
nor U15542 (N_15542,N_12579,N_14277);
xnor U15543 (N_15543,N_12961,N_10498);
nor U15544 (N_15544,N_11313,N_11777);
nor U15545 (N_15545,N_11236,N_12511);
and U15546 (N_15546,N_11143,N_12128);
and U15547 (N_15547,N_12637,N_10985);
nand U15548 (N_15548,N_14548,N_14720);
xor U15549 (N_15549,N_14253,N_14507);
xnor U15550 (N_15550,N_13729,N_12848);
nor U15551 (N_15551,N_12233,N_13192);
or U15552 (N_15552,N_10389,N_11047);
xor U15553 (N_15553,N_14783,N_10513);
xor U15554 (N_15554,N_10922,N_13323);
or U15555 (N_15555,N_12239,N_11676);
and U15556 (N_15556,N_12950,N_12247);
nand U15557 (N_15557,N_11519,N_13534);
and U15558 (N_15558,N_13035,N_10643);
nand U15559 (N_15559,N_13021,N_11105);
nor U15560 (N_15560,N_10048,N_14670);
or U15561 (N_15561,N_10169,N_14565);
nand U15562 (N_15562,N_12255,N_10002);
and U15563 (N_15563,N_11037,N_13045);
nor U15564 (N_15564,N_13248,N_11946);
xnor U15565 (N_15565,N_10628,N_13256);
or U15566 (N_15566,N_10426,N_13213);
or U15567 (N_15567,N_11878,N_12487);
or U15568 (N_15568,N_11774,N_12134);
xor U15569 (N_15569,N_14389,N_10960);
and U15570 (N_15570,N_14183,N_11348);
xnor U15571 (N_15571,N_13523,N_10811);
and U15572 (N_15572,N_10226,N_11659);
nor U15573 (N_15573,N_13791,N_12573);
nor U15574 (N_15574,N_14826,N_11785);
nand U15575 (N_15575,N_11845,N_12670);
and U15576 (N_15576,N_11242,N_13774);
nand U15577 (N_15577,N_13612,N_12139);
nor U15578 (N_15578,N_12739,N_11322);
nand U15579 (N_15579,N_11257,N_12455);
nand U15580 (N_15580,N_12546,N_13969);
nor U15581 (N_15581,N_10958,N_11028);
and U15582 (N_15582,N_10148,N_12936);
xor U15583 (N_15583,N_12666,N_10396);
and U15584 (N_15584,N_14947,N_14344);
and U15585 (N_15585,N_14580,N_14572);
nor U15586 (N_15586,N_14715,N_12252);
or U15587 (N_15587,N_13665,N_12285);
nand U15588 (N_15588,N_11181,N_10428);
xnor U15589 (N_15589,N_13923,N_12119);
nor U15590 (N_15590,N_11373,N_12424);
nand U15591 (N_15591,N_10823,N_14267);
or U15592 (N_15592,N_10230,N_13645);
nand U15593 (N_15593,N_13769,N_14579);
or U15594 (N_15594,N_14273,N_11645);
nand U15595 (N_15595,N_11888,N_11289);
xnor U15596 (N_15596,N_14101,N_11894);
and U15597 (N_15597,N_11749,N_11298);
and U15598 (N_15598,N_12192,N_12795);
xnor U15599 (N_15599,N_10395,N_12284);
and U15600 (N_15600,N_10335,N_14006);
xor U15601 (N_15601,N_13818,N_13064);
xnor U15602 (N_15602,N_12356,N_10075);
nand U15603 (N_15603,N_14027,N_14939);
xnor U15604 (N_15604,N_14085,N_14611);
and U15605 (N_15605,N_11123,N_13322);
nor U15606 (N_15606,N_12027,N_12104);
or U15607 (N_15607,N_13477,N_10849);
or U15608 (N_15608,N_13527,N_12467);
nor U15609 (N_15609,N_12224,N_10143);
xnor U15610 (N_15610,N_12680,N_12513);
nand U15611 (N_15611,N_13431,N_10571);
nor U15612 (N_15612,N_13806,N_10970);
nor U15613 (N_15613,N_13335,N_10462);
xor U15614 (N_15614,N_13582,N_13382);
and U15615 (N_15615,N_12149,N_14883);
xnor U15616 (N_15616,N_14995,N_11504);
nor U15617 (N_15617,N_10479,N_13101);
nand U15618 (N_15618,N_12097,N_14138);
nand U15619 (N_15619,N_10990,N_14012);
and U15620 (N_15620,N_12235,N_12418);
nor U15621 (N_15621,N_10051,N_13704);
and U15622 (N_15622,N_14454,N_14041);
nand U15623 (N_15623,N_14413,N_12653);
xor U15624 (N_15624,N_10520,N_14496);
nand U15625 (N_15625,N_14447,N_11499);
xnor U15626 (N_15626,N_14211,N_12063);
nand U15627 (N_15627,N_12590,N_12854);
or U15628 (N_15628,N_11071,N_14922);
or U15629 (N_15629,N_13068,N_12600);
or U15630 (N_15630,N_14999,N_13838);
or U15631 (N_15631,N_10535,N_12310);
nor U15632 (N_15632,N_11917,N_10637);
nor U15633 (N_15633,N_13410,N_11931);
or U15634 (N_15634,N_13367,N_14464);
xnor U15635 (N_15635,N_14741,N_10126);
xnor U15636 (N_15636,N_11068,N_13865);
xor U15637 (N_15637,N_10093,N_11723);
or U15638 (N_15638,N_14262,N_12947);
xnor U15639 (N_15639,N_14099,N_13964);
nor U15640 (N_15640,N_10062,N_10467);
or U15641 (N_15641,N_13750,N_11067);
and U15642 (N_15642,N_14030,N_11500);
xor U15643 (N_15643,N_14270,N_13111);
nand U15644 (N_15644,N_10837,N_14298);
and U15645 (N_15645,N_14642,N_13853);
and U15646 (N_15646,N_13211,N_13265);
xor U15647 (N_15647,N_12940,N_11691);
and U15648 (N_15648,N_10848,N_13849);
xnor U15649 (N_15649,N_11161,N_11295);
xor U15650 (N_15650,N_12633,N_13439);
nor U15651 (N_15651,N_13196,N_13957);
and U15652 (N_15652,N_13290,N_12738);
nor U15653 (N_15653,N_10499,N_14600);
nor U15654 (N_15654,N_11684,N_14661);
xor U15655 (N_15655,N_11941,N_13472);
or U15656 (N_15656,N_13617,N_10357);
nor U15657 (N_15657,N_12081,N_10579);
xnor U15658 (N_15658,N_10540,N_11226);
nor U15659 (N_15659,N_13759,N_10207);
nor U15660 (N_15660,N_12797,N_10666);
or U15661 (N_15661,N_14988,N_12724);
nor U15662 (N_15662,N_12244,N_11270);
or U15663 (N_15663,N_10103,N_10488);
or U15664 (N_15664,N_14503,N_13776);
and U15665 (N_15665,N_11563,N_13537);
or U15666 (N_15666,N_14673,N_12057);
nand U15667 (N_15667,N_11467,N_14781);
and U15668 (N_15668,N_14081,N_12355);
or U15669 (N_15669,N_12923,N_14244);
nand U15670 (N_15670,N_14276,N_14083);
or U15671 (N_15671,N_13446,N_14594);
nor U15672 (N_15672,N_12939,N_12941);
and U15673 (N_15673,N_12981,N_14871);
nor U15674 (N_15674,N_14958,N_10966);
and U15675 (N_15675,N_12731,N_10701);
or U15676 (N_15676,N_11021,N_12942);
nand U15677 (N_15677,N_11875,N_11427);
nor U15678 (N_15678,N_11934,N_13447);
nor U15679 (N_15679,N_13526,N_11104);
and U15680 (N_15680,N_10863,N_14903);
or U15681 (N_15681,N_13007,N_11114);
xor U15682 (N_15682,N_14838,N_14197);
nand U15683 (N_15683,N_11491,N_11014);
and U15684 (N_15684,N_14608,N_10801);
or U15685 (N_15685,N_14551,N_10786);
nand U15686 (N_15686,N_12114,N_12468);
xor U15687 (N_15687,N_12482,N_12995);
xnor U15688 (N_15688,N_10170,N_12559);
nor U15689 (N_15689,N_14074,N_10436);
and U15690 (N_15690,N_14040,N_11916);
or U15691 (N_15691,N_11107,N_12910);
or U15692 (N_15692,N_14170,N_14272);
or U15693 (N_15693,N_14675,N_12527);
nand U15694 (N_15694,N_12156,N_10457);
or U15695 (N_15695,N_12937,N_14613);
and U15696 (N_15696,N_12617,N_14707);
xor U15697 (N_15697,N_13755,N_13882);
or U15698 (N_15698,N_10225,N_11791);
nor U15699 (N_15699,N_12220,N_11299);
nand U15700 (N_15700,N_11414,N_11859);
or U15701 (N_15701,N_12550,N_11471);
or U15702 (N_15702,N_11429,N_10639);
nor U15703 (N_15703,N_10351,N_14260);
or U15704 (N_15704,N_12708,N_13887);
nor U15705 (N_15705,N_11380,N_14914);
nand U15706 (N_15706,N_13940,N_11240);
or U15707 (N_15707,N_14704,N_10348);
or U15708 (N_15708,N_12660,N_12998);
and U15709 (N_15709,N_14398,N_11871);
nand U15710 (N_15710,N_10392,N_10570);
nor U15711 (N_15711,N_12753,N_12329);
or U15712 (N_15712,N_11219,N_11823);
and U15713 (N_15713,N_13317,N_10209);
nor U15714 (N_15714,N_13681,N_12198);
xnor U15715 (N_15715,N_10832,N_12125);
xnor U15716 (N_15716,N_13067,N_11668);
or U15717 (N_15717,N_11927,N_13724);
nand U15718 (N_15718,N_12821,N_14614);
xor U15719 (N_15719,N_12118,N_13539);
xnor U15720 (N_15720,N_11211,N_14166);
and U15721 (N_15721,N_12888,N_12810);
and U15722 (N_15722,N_13649,N_14355);
nor U15723 (N_15723,N_12658,N_12403);
and U15724 (N_15724,N_12834,N_11378);
nand U15725 (N_15725,N_13450,N_10781);
nand U15726 (N_15726,N_14229,N_13296);
and U15727 (N_15727,N_11583,N_12839);
and U15728 (N_15728,N_14359,N_11686);
xnor U15729 (N_15729,N_14694,N_14332);
and U15730 (N_15730,N_11810,N_11974);
xnor U15731 (N_15731,N_11755,N_11327);
and U15732 (N_15732,N_14978,N_11433);
xnor U15733 (N_15733,N_12286,N_14935);
nand U15734 (N_15734,N_10167,N_12187);
nor U15735 (N_15735,N_14682,N_11106);
xnor U15736 (N_15736,N_13112,N_13642);
xnor U15737 (N_15737,N_11613,N_11981);
nand U15738 (N_15738,N_13133,N_13895);
or U15739 (N_15739,N_12826,N_10580);
nand U15740 (N_15740,N_11665,N_12222);
or U15741 (N_15741,N_10259,N_13307);
xnor U15742 (N_15742,N_11980,N_14861);
xnor U15743 (N_15743,N_12225,N_10921);
nand U15744 (N_15744,N_12706,N_10405);
xnor U15745 (N_15745,N_10808,N_12921);
or U15746 (N_15746,N_10870,N_11960);
and U15747 (N_15747,N_13232,N_12655);
nand U15748 (N_15748,N_14239,N_13123);
xor U15749 (N_15749,N_11982,N_13294);
and U15750 (N_15750,N_10301,N_12897);
nand U15751 (N_15751,N_12879,N_10555);
nor U15752 (N_15752,N_12180,N_14386);
and U15753 (N_15753,N_13829,N_12962);
xnor U15754 (N_15754,N_12122,N_14345);
and U15755 (N_15755,N_13870,N_11031);
nor U15756 (N_15756,N_13587,N_11056);
xor U15757 (N_15757,N_13507,N_14795);
nor U15758 (N_15758,N_11199,N_13948);
and U15759 (N_15759,N_10751,N_12829);
or U15760 (N_15760,N_13273,N_10271);
and U15761 (N_15761,N_11001,N_12398);
and U15762 (N_15762,N_10310,N_13110);
or U15763 (N_15763,N_10234,N_14963);
and U15764 (N_15764,N_13548,N_13876);
xor U15765 (N_15765,N_12191,N_11395);
or U15766 (N_15766,N_13107,N_10149);
xor U15767 (N_15767,N_14821,N_10878);
nand U15768 (N_15768,N_14200,N_13202);
nor U15769 (N_15769,N_11855,N_13732);
nor U15770 (N_15770,N_12053,N_10014);
xor U15771 (N_15771,N_11359,N_12510);
or U15772 (N_15772,N_11883,N_13749);
or U15773 (N_15773,N_12849,N_13148);
nand U15774 (N_15774,N_14970,N_13234);
or U15775 (N_15775,N_10777,N_12963);
nand U15776 (N_15776,N_13221,N_10834);
nor U15777 (N_15777,N_13131,N_14455);
nand U15778 (N_15778,N_10697,N_11216);
xnor U15779 (N_15779,N_11205,N_12358);
nor U15780 (N_15780,N_10791,N_12200);
xnor U15781 (N_15781,N_11631,N_12784);
or U15782 (N_15782,N_12860,N_14180);
and U15783 (N_15783,N_14811,N_10214);
nor U15784 (N_15784,N_14818,N_14957);
nand U15785 (N_15785,N_11672,N_12169);
and U15786 (N_15786,N_11300,N_14649);
xor U15787 (N_15787,N_13904,N_12620);
xnor U15788 (N_15788,N_10178,N_12685);
xor U15789 (N_15789,N_12335,N_10034);
nand U15790 (N_15790,N_13116,N_10318);
nand U15791 (N_15791,N_13098,N_12429);
nor U15792 (N_15792,N_11407,N_10155);
nor U15793 (N_15793,N_13745,N_12372);
xnor U15794 (N_15794,N_10612,N_14728);
and U15795 (N_15795,N_11374,N_14352);
nor U15796 (N_15796,N_10453,N_11607);
and U15797 (N_15797,N_11963,N_10258);
and U15798 (N_15798,N_14136,N_10965);
and U15799 (N_15799,N_14363,N_11425);
and U15800 (N_15800,N_13530,N_11644);
or U15801 (N_15801,N_11687,N_12847);
xor U15802 (N_15802,N_12442,N_13835);
nor U15803 (N_15803,N_12618,N_11968);
nor U15804 (N_15804,N_14034,N_10368);
nand U15805 (N_15805,N_13988,N_11807);
xnor U15806 (N_15806,N_13707,N_12091);
nand U15807 (N_15807,N_13333,N_11521);
nand U15808 (N_15808,N_10879,N_13789);
and U15809 (N_15809,N_10525,N_10303);
and U15810 (N_15810,N_10941,N_13490);
nand U15811 (N_15811,N_12313,N_12979);
or U15812 (N_15812,N_10515,N_11479);
nor U15813 (N_15813,N_10144,N_14487);
nor U15814 (N_15814,N_13139,N_13003);
or U15815 (N_15815,N_11892,N_11209);
nand U15816 (N_15816,N_14533,N_13254);
nor U15817 (N_15817,N_11604,N_14892);
nor U15818 (N_15818,N_10889,N_13863);
nand U15819 (N_15819,N_12956,N_12743);
and U15820 (N_15820,N_10874,N_14234);
nand U15821 (N_15821,N_11122,N_11904);
or U15822 (N_15822,N_10355,N_10577);
and U15823 (N_15823,N_11517,N_14740);
and U15824 (N_15824,N_11084,N_10730);
xor U15825 (N_15825,N_10238,N_10399);
nand U15826 (N_15826,N_14366,N_14562);
and U15827 (N_15827,N_12808,N_14241);
nand U15828 (N_15828,N_12705,N_13166);
nand U15829 (N_15829,N_11153,N_10328);
and U15830 (N_15830,N_12825,N_11595);
nor U15831 (N_15831,N_11018,N_14290);
and U15832 (N_15832,N_13992,N_14302);
and U15833 (N_15833,N_10853,N_13701);
nand U15834 (N_15834,N_14237,N_13734);
nor U15835 (N_15835,N_13419,N_12917);
and U15836 (N_15836,N_12711,N_12803);
and U15837 (N_15837,N_14902,N_13584);
or U15838 (N_15838,N_12668,N_12585);
and U15839 (N_15839,N_13949,N_13601);
nand U15840 (N_15840,N_10091,N_13702);
nand U15841 (N_15841,N_14238,N_14452);
or U15842 (N_15842,N_13424,N_10264);
or U15843 (N_15843,N_13857,N_11141);
xnor U15844 (N_15844,N_13657,N_13494);
and U15845 (N_15845,N_11935,N_13795);
nor U15846 (N_15846,N_14382,N_13989);
nor U15847 (N_15847,N_12560,N_11772);
and U15848 (N_15848,N_10893,N_10789);
xnor U15849 (N_15849,N_14443,N_11278);
nand U15850 (N_15850,N_10145,N_12017);
xnor U15851 (N_15851,N_13960,N_14941);
nand U15852 (N_15852,N_12969,N_10090);
or U15853 (N_15853,N_12999,N_13772);
or U15854 (N_15854,N_13377,N_11323);
nor U15855 (N_15855,N_14346,N_11998);
nand U15856 (N_15856,N_10689,N_14329);
nand U15857 (N_15857,N_12032,N_14721);
or U15858 (N_15858,N_11757,N_14629);
nand U15859 (N_15859,N_12360,N_12506);
nand U15860 (N_15860,N_14991,N_13735);
nor U15861 (N_15861,N_13454,N_11545);
nor U15862 (N_15862,N_11502,N_11394);
or U15863 (N_15863,N_13766,N_13929);
and U15864 (N_15864,N_14463,N_13363);
nand U15865 (N_15865,N_13782,N_11786);
and U15866 (N_15866,N_12043,N_10748);
nand U15867 (N_15867,N_11787,N_14415);
or U15868 (N_15868,N_12836,N_14967);
or U15869 (N_15869,N_14271,N_13324);
xor U15870 (N_15870,N_10459,N_10334);
nor U15871 (N_15871,N_12769,N_10606);
nor U15872 (N_15872,N_13099,N_11703);
xor U15873 (N_15873,N_12786,N_14499);
or U15874 (N_15874,N_14488,N_11709);
and U15875 (N_15875,N_14779,N_11600);
xor U15876 (N_15876,N_14039,N_14747);
nor U15877 (N_15877,N_13298,N_11933);
and U15878 (N_15878,N_11377,N_10901);
and U15879 (N_15879,N_12982,N_13867);
nand U15880 (N_15880,N_14748,N_14297);
xnor U15881 (N_15881,N_14460,N_11689);
xnor U15882 (N_15882,N_11985,N_12326);
or U15883 (N_15883,N_12760,N_14905);
nand U15884 (N_15884,N_14895,N_14134);
and U15885 (N_15885,N_10673,N_14418);
and U15886 (N_15886,N_11972,N_12781);
nand U15887 (N_15887,N_13301,N_12549);
nand U15888 (N_15888,N_13108,N_11296);
and U15889 (N_15889,N_13770,N_13360);
xnor U15890 (N_15890,N_12394,N_12571);
nand U15891 (N_15891,N_13618,N_10652);
and U15892 (N_15892,N_11505,N_14760);
nand U15893 (N_15893,N_14667,N_11396);
nor U15894 (N_15894,N_10332,N_13425);
nor U15895 (N_15895,N_10059,N_14824);
or U15896 (N_15896,N_11814,N_10138);
nor U15897 (N_15897,N_13554,N_13955);
or U15898 (N_15898,N_11572,N_12474);
or U15899 (N_15899,N_13215,N_12672);
nor U15900 (N_15900,N_11265,N_10557);
nand U15901 (N_15901,N_12806,N_10350);
or U15902 (N_15902,N_13005,N_11552);
or U15903 (N_15903,N_13011,N_12375);
and U15904 (N_15904,N_12020,N_14936);
and U15905 (N_15905,N_10758,N_10718);
or U15906 (N_15906,N_13647,N_11854);
xnor U15907 (N_15907,N_12223,N_14019);
xor U15908 (N_15908,N_10412,N_11928);
nand U15909 (N_15909,N_10007,N_13521);
nand U15910 (N_15910,N_13451,N_10954);
xor U15911 (N_15911,N_11923,N_11198);
or U15912 (N_15912,N_11389,N_11158);
nand U15913 (N_15913,N_10799,N_10905);
xor U15914 (N_15914,N_13973,N_11444);
or U15915 (N_15915,N_12835,N_10644);
xor U15916 (N_15916,N_12129,N_10022);
nand U15917 (N_15917,N_12092,N_11498);
or U15918 (N_15918,N_13604,N_14147);
or U15919 (N_15919,N_14462,N_14475);
nor U15920 (N_15920,N_10012,N_12166);
and U15921 (N_15921,N_11556,N_11652);
nand U15922 (N_15922,N_11366,N_12197);
nand U15923 (N_15923,N_12461,N_12682);
or U15924 (N_15924,N_14513,N_11510);
nand U15925 (N_15925,N_13271,N_14122);
and U15926 (N_15926,N_14635,N_10232);
nor U15927 (N_15927,N_11793,N_12475);
or U15928 (N_15928,N_13922,N_13709);
or U15929 (N_15929,N_14278,N_10573);
nand U15930 (N_15930,N_12213,N_11655);
xor U15931 (N_15931,N_10313,N_12916);
nand U15932 (N_15932,N_12993,N_11057);
xnor U15933 (N_15933,N_12994,N_12018);
nand U15934 (N_15934,N_11950,N_14198);
nand U15935 (N_15935,N_13747,N_14537);
nand U15936 (N_15936,N_10788,N_12435);
or U15937 (N_15937,N_12712,N_14808);
nor U15938 (N_15938,N_10439,N_11367);
xor U15939 (N_15939,N_10454,N_10274);
xor U15940 (N_15940,N_13883,N_10267);
or U15941 (N_15941,N_14664,N_14750);
nor U15942 (N_15942,N_11049,N_12873);
or U15943 (N_15943,N_11145,N_11404);
xnor U15944 (N_15944,N_14406,N_10650);
xnor U15945 (N_15945,N_12622,N_12277);
and U15946 (N_15946,N_12145,N_10430);
and U15947 (N_15947,N_14404,N_14193);
nand U15948 (N_15948,N_14734,N_12387);
and U15949 (N_15949,N_13656,N_14930);
and U15950 (N_15950,N_13077,N_11117);
nand U15951 (N_15951,N_10815,N_11630);
nand U15952 (N_15952,N_10558,N_13568);
or U15953 (N_15953,N_12673,N_14893);
xnor U15954 (N_15954,N_14569,N_13803);
and U15955 (N_15955,N_14282,N_10590);
nand U15956 (N_15956,N_10208,N_13811);
or U15957 (N_15957,N_12301,N_12958);
nand U15958 (N_15958,N_11956,N_14056);
nand U15959 (N_15959,N_10110,N_12524);
nand U15960 (N_15960,N_14372,N_11269);
xnor U15961 (N_15961,N_13779,N_11096);
nor U15962 (N_15962,N_13406,N_13038);
nand U15963 (N_15963,N_14526,N_13416);
nor U15964 (N_15964,N_10887,N_13203);
or U15965 (N_15965,N_11440,N_13817);
xnor U15966 (N_15966,N_13577,N_11497);
xor U15967 (N_15967,N_10358,N_12338);
and U15968 (N_15968,N_10517,N_12952);
nor U15969 (N_15969,N_11590,N_12498);
nor U15970 (N_15970,N_11666,N_14003);
nor U15971 (N_15971,N_12688,N_11841);
xor U15972 (N_15972,N_13815,N_11121);
and U15973 (N_15973,N_14938,N_12378);
xor U15974 (N_15974,N_11729,N_12437);
xor U15975 (N_15975,N_13897,N_14367);
nand U15976 (N_15976,N_13420,N_12677);
or U15977 (N_15977,N_11007,N_10064);
or U15978 (N_15978,N_14621,N_10477);
and U15979 (N_15979,N_14428,N_14772);
or U15980 (N_15980,N_14154,N_11437);
nand U15981 (N_15981,N_10397,N_10444);
nand U15982 (N_15982,N_12844,N_14669);
or U15983 (N_15983,N_13126,N_10066);
nand U15984 (N_15984,N_10369,N_14115);
and U15985 (N_15985,N_10658,N_12876);
xor U15986 (N_15986,N_10681,N_13334);
xnor U15987 (N_15987,N_11737,N_14771);
and U15988 (N_15988,N_14119,N_14998);
nor U15989 (N_15989,N_11488,N_12008);
nor U15990 (N_15990,N_10814,N_14204);
nor U15991 (N_15991,N_13963,N_12920);
xor U15992 (N_15992,N_12184,N_10629);
or U15993 (N_15993,N_11837,N_13433);
and U15994 (N_15994,N_14492,N_10661);
or U15995 (N_15995,N_11388,N_12282);
or U15996 (N_15996,N_10553,N_10607);
and U15997 (N_15997,N_13723,N_12697);
or U15998 (N_15998,N_13034,N_11081);
nor U15999 (N_15999,N_13725,N_10413);
and U16000 (N_16000,N_13282,N_12036);
nand U16001 (N_16001,N_12266,N_13990);
nor U16002 (N_16002,N_13194,N_13886);
nand U16003 (N_16003,N_13114,N_13717);
xor U16004 (N_16004,N_11134,N_10593);
nor U16005 (N_16005,N_12268,N_11701);
and U16006 (N_16006,N_13238,N_10432);
or U16007 (N_16007,N_10861,N_13320);
or U16008 (N_16008,N_10810,N_10215);
nor U16009 (N_16009,N_10929,N_11940);
or U16010 (N_16010,N_13417,N_11766);
xor U16011 (N_16011,N_10687,N_11911);
and U16012 (N_16012,N_13106,N_12175);
or U16013 (N_16013,N_11137,N_14401);
and U16014 (N_16014,N_14532,N_10339);
nor U16015 (N_16015,N_13230,N_10624);
nor U16016 (N_16016,N_10299,N_12693);
nand U16017 (N_16017,N_12471,N_14185);
nor U16018 (N_16018,N_11074,N_14279);
nor U16019 (N_16019,N_10585,N_12070);
nor U16020 (N_16020,N_11896,N_13936);
xnor U16021 (N_16021,N_13850,N_10199);
nor U16022 (N_16022,N_13514,N_12730);
or U16023 (N_16023,N_10173,N_11764);
and U16024 (N_16024,N_12083,N_12218);
and U16025 (N_16025,N_11601,N_12748);
nor U16026 (N_16026,N_12281,N_14643);
nor U16027 (N_16027,N_11893,N_12410);
and U16028 (N_16028,N_11863,N_10057);
xnor U16029 (N_16029,N_13974,N_14605);
xor U16030 (N_16030,N_14127,N_11286);
xor U16031 (N_16031,N_13627,N_12137);
and U16032 (N_16032,N_11403,N_11419);
xor U16033 (N_16033,N_14742,N_13809);
or U16034 (N_16034,N_13146,N_13982);
and U16035 (N_16035,N_14046,N_11463);
or U16036 (N_16036,N_11370,N_11206);
xnor U16037 (N_16037,N_10487,N_10733);
nand U16038 (N_16038,N_14589,N_14869);
or U16039 (N_16039,N_14444,N_10805);
and U16040 (N_16040,N_10127,N_10105);
nor U16041 (N_16041,N_12103,N_12907);
xnor U16042 (N_16042,N_12698,N_13580);
or U16043 (N_16043,N_11673,N_12751);
and U16044 (N_16044,N_13242,N_10378);
nor U16045 (N_16045,N_13913,N_11577);
or U16046 (N_16046,N_13346,N_10964);
and U16047 (N_16047,N_11682,N_10850);
nor U16048 (N_16048,N_11252,N_11694);
nor U16049 (N_16049,N_11575,N_10314);
nor U16050 (N_16050,N_11287,N_13025);
nand U16051 (N_16051,N_14000,N_11873);
or U16052 (N_16052,N_10094,N_12548);
nand U16053 (N_16053,N_14461,N_14419);
or U16054 (N_16054,N_14142,N_10631);
and U16055 (N_16055,N_10100,N_14591);
nor U16056 (N_16056,N_13427,N_10137);
nor U16057 (N_16057,N_11828,N_11945);
nor U16058 (N_16058,N_12778,N_11477);
and U16059 (N_16059,N_14274,N_14181);
nor U16060 (N_16060,N_13058,N_11653);
xor U16061 (N_16061,N_14296,N_13862);
and U16062 (N_16062,N_14314,N_14681);
and U16063 (N_16063,N_10724,N_11633);
xor U16064 (N_16064,N_14713,N_13137);
xnor U16065 (N_16065,N_13600,N_14062);
or U16066 (N_16066,N_13676,N_14498);
nand U16067 (N_16067,N_10086,N_10080);
or U16068 (N_16068,N_13888,N_14859);
nand U16069 (N_16069,N_14959,N_12412);
or U16070 (N_16070,N_12540,N_14714);
nand U16071 (N_16071,N_11886,N_13047);
and U16072 (N_16072,N_13628,N_13188);
and U16073 (N_16073,N_10939,N_10364);
nor U16074 (N_16074,N_12990,N_10277);
and U16075 (N_16075,N_11947,N_12384);
nand U16076 (N_16076,N_11159,N_14135);
xnor U16077 (N_16077,N_10756,N_11884);
and U16078 (N_16078,N_14458,N_10995);
nand U16079 (N_16079,N_12291,N_10175);
nor U16080 (N_16080,N_13489,N_11248);
xnor U16081 (N_16081,N_14226,N_13754);
or U16082 (N_16082,N_10408,N_13858);
nand U16083 (N_16083,N_13843,N_12470);
or U16084 (N_16084,N_10717,N_11929);
nor U16085 (N_16085,N_12050,N_10821);
or U16086 (N_16086,N_14387,N_14901);
and U16087 (N_16087,N_11862,N_10027);
and U16088 (N_16088,N_12804,N_11054);
and U16089 (N_16089,N_12944,N_12800);
or U16090 (N_16090,N_10324,N_11410);
or U16091 (N_16091,N_12662,N_13700);
nand U16092 (N_16092,N_13687,N_11616);
xnor U16093 (N_16093,N_11868,N_12311);
nand U16094 (N_16094,N_12457,N_13252);
xnor U16095 (N_16095,N_14053,N_13201);
and U16096 (N_16096,N_12607,N_12388);
nand U16097 (N_16097,N_14866,N_11493);
and U16098 (N_16098,N_14814,N_14776);
or U16099 (N_16099,N_12229,N_13418);
nor U16100 (N_16100,N_13946,N_10933);
nand U16101 (N_16101,N_11157,N_13094);
or U16102 (N_16102,N_10544,N_13438);
and U16103 (N_16103,N_13009,N_11275);
nand U16104 (N_16104,N_14528,N_11861);
nand U16105 (N_16105,N_10146,N_12631);
nor U16106 (N_16106,N_10862,N_11858);
and U16107 (N_16107,N_11305,N_11334);
nand U16108 (N_16108,N_12985,N_11343);
or U16109 (N_16109,N_13689,N_13908);
and U16110 (N_16110,N_11906,N_12595);
xnor U16111 (N_16111,N_12064,N_13746);
or U16112 (N_16112,N_14638,N_12312);
nand U16113 (N_16113,N_12262,N_10634);
or U16114 (N_16114,N_12740,N_10018);
or U16115 (N_16115,N_11903,N_12519);
or U16116 (N_16116,N_14543,N_13561);
nor U16117 (N_16117,N_12704,N_12279);
nand U16118 (N_16118,N_10550,N_13163);
nor U16119 (N_16119,N_14423,N_13269);
xor U16120 (N_16120,N_14469,N_13947);
nand U16121 (N_16121,N_11565,N_10812);
and U16122 (N_16122,N_12669,N_11255);
nand U16123 (N_16123,N_10678,N_14002);
and U16124 (N_16124,N_12248,N_13218);
xnor U16125 (N_16125,N_13971,N_12612);
nor U16126 (N_16126,N_12734,N_14782);
or U16127 (N_16127,N_14225,N_11155);
or U16128 (N_16128,N_10505,N_12132);
and U16129 (N_16129,N_11385,N_13342);
nor U16130 (N_16130,N_12376,N_12863);
nor U16131 (N_16131,N_11857,N_11302);
nor U16132 (N_16132,N_10272,N_10959);
nor U16133 (N_16133,N_12300,N_10293);
and U16134 (N_16134,N_10136,N_13072);
nand U16135 (N_16135,N_14326,N_11230);
and U16136 (N_16136,N_12260,N_14825);
or U16137 (N_16137,N_13555,N_14380);
xnor U16138 (N_16138,N_13528,N_13716);
nand U16139 (N_16139,N_14028,N_11011);
and U16140 (N_16140,N_11596,N_11227);
nor U16141 (N_16141,N_13624,N_12241);
xor U16142 (N_16142,N_11621,N_10740);
nor U16143 (N_16143,N_12875,N_11816);
and U16144 (N_16144,N_10833,N_14209);
or U16145 (N_16145,N_11495,N_14812);
and U16146 (N_16146,N_11120,N_10121);
xnor U16147 (N_16147,N_13306,N_12263);
xnor U16148 (N_16148,N_11860,N_12090);
and U16149 (N_16149,N_13362,N_13022);
nand U16150 (N_16150,N_10682,N_13432);
nor U16151 (N_16151,N_13381,N_14552);
nand U16152 (N_16152,N_11898,N_10095);
nand U16153 (N_16153,N_11016,N_12022);
and U16154 (N_16154,N_12116,N_11900);
nor U16155 (N_16155,N_12922,N_13677);
nand U16156 (N_16156,N_12370,N_11301);
nand U16157 (N_16157,N_11657,N_11966);
nor U16158 (N_16158,N_11112,N_11239);
xor U16159 (N_16159,N_13524,N_13400);
nor U16160 (N_16160,N_14550,N_10955);
xor U16161 (N_16161,N_11970,N_10036);
or U16162 (N_16162,N_13214,N_11986);
or U16163 (N_16163,N_12586,N_10635);
xor U16164 (N_16164,N_13308,N_11813);
nor U16165 (N_16165,N_11118,N_10537);
nand U16166 (N_16166,N_12193,N_10347);
and U16167 (N_16167,N_12352,N_13030);
or U16168 (N_16168,N_12380,N_11060);
and U16169 (N_16169,N_14623,N_14044);
and U16170 (N_16170,N_14078,N_11470);
nand U16171 (N_16171,N_10502,N_10419);
and U16172 (N_16172,N_14786,N_11826);
nor U16173 (N_16173,N_11636,N_13314);
or U16174 (N_16174,N_13391,N_13312);
or U16175 (N_16175,N_14465,N_11361);
or U16176 (N_16176,N_14320,N_10068);
xor U16177 (N_16177,N_12431,N_10522);
nand U16178 (N_16178,N_14658,N_14685);
nor U16179 (N_16179,N_14370,N_12908);
and U16180 (N_16180,N_12353,N_11333);
and U16181 (N_16181,N_12886,N_12722);
or U16182 (N_16182,N_12445,N_14409);
nand U16183 (N_16183,N_11921,N_11442);
nand U16184 (N_16184,N_11092,N_14990);
xor U16185 (N_16185,N_14008,N_10492);
and U16186 (N_16186,N_13090,N_13386);
nand U16187 (N_16187,N_12636,N_11853);
xor U16188 (N_16188,N_12016,N_14383);
nor U16189 (N_16189,N_11204,N_12351);
and U16190 (N_16190,N_12537,N_10159);
nand U16191 (N_16191,N_10605,N_11770);
xnor U16192 (N_16192,N_11353,N_11185);
nand U16193 (N_16193,N_10713,N_10851);
or U16194 (N_16194,N_14144,N_11005);
xnor U16195 (N_16195,N_10029,N_11850);
nand U16196 (N_16196,N_11795,N_13122);
or U16197 (N_16197,N_14336,N_10101);
nor U16198 (N_16198,N_10112,N_14073);
nor U16199 (N_16199,N_10393,N_12989);
xor U16200 (N_16200,N_13277,N_10521);
nor U16201 (N_16201,N_11879,N_14948);
or U16202 (N_16202,N_13688,N_13199);
xor U16203 (N_16203,N_13457,N_14637);
and U16204 (N_16204,N_14921,N_14833);
nor U16205 (N_16205,N_13492,N_13198);
or U16206 (N_16206,N_14227,N_11326);
nand U16207 (N_16207,N_10204,N_13156);
xor U16208 (N_16208,N_12520,N_10304);
nand U16209 (N_16209,N_13008,N_14378);
and U16210 (N_16210,N_10532,N_13119);
nor U16211 (N_16211,N_10913,N_10072);
and U16212 (N_16212,N_12460,N_12278);
nand U16213 (N_16213,N_14013,N_11809);
and U16214 (N_16214,N_12296,N_10526);
or U16215 (N_16215,N_11594,N_10359);
nand U16216 (N_16216,N_13031,N_12077);
nor U16217 (N_16217,N_12432,N_12577);
xor U16218 (N_16218,N_12466,N_13938);
or U16219 (N_16219,N_14985,N_12189);
xor U16220 (N_16220,N_11083,N_14944);
xnor U16221 (N_16221,N_13384,N_10493);
nand U16222 (N_16222,N_11357,N_13820);
or U16223 (N_16223,N_12066,N_14663);
or U16224 (N_16224,N_11822,N_13655);
nand U16225 (N_16225,N_13220,N_13281);
xnor U16226 (N_16226,N_11017,N_13285);
xnor U16227 (N_16227,N_12855,N_11132);
nand U16228 (N_16228,N_14908,N_14604);
or U16229 (N_16229,N_12525,N_14486);
and U16230 (N_16230,N_11663,N_13585);
nor U16231 (N_16231,N_14374,N_13937);
xor U16232 (N_16232,N_14328,N_11271);
nor U16233 (N_16233,N_12141,N_12650);
nor U16234 (N_16234,N_10362,N_10686);
or U16235 (N_16235,N_14616,N_13593);
or U16236 (N_16236,N_12003,N_12959);
nor U16237 (N_16237,N_13468,N_13411);
nor U16238 (N_16238,N_14735,N_14559);
nand U16239 (N_16239,N_11390,N_12438);
nand U16240 (N_16240,N_12452,N_12464);
and U16241 (N_16241,N_10415,N_11012);
xor U16242 (N_16242,N_10205,N_14224);
nand U16243 (N_16243,N_14676,N_11154);
nand U16244 (N_16244,N_12727,N_10945);
xnor U16245 (N_16245,N_10433,N_11237);
and U16246 (N_16246,N_11872,N_13823);
or U16247 (N_16247,N_11805,N_13097);
xnor U16248 (N_16248,N_11671,N_12089);
nand U16249 (N_16249,N_13757,N_12927);
nand U16250 (N_16250,N_10099,N_10289);
nor U16251 (N_16251,N_10153,N_14867);
nand U16252 (N_16252,N_13177,N_14977);
nand U16253 (N_16253,N_13217,N_10349);
or U16254 (N_16254,N_11720,N_10700);
nor U16255 (N_16255,N_10937,N_13565);
nand U16256 (N_16256,N_12133,N_11901);
xor U16257 (N_16257,N_12798,N_12754);
or U16258 (N_16258,N_11431,N_10651);
nand U16259 (N_16259,N_11035,N_11506);
nand U16260 (N_16260,N_13679,N_10784);
or U16261 (N_16261,N_10660,N_10049);
nand U16262 (N_16262,N_12557,N_12154);
nor U16263 (N_16263,N_12374,N_12208);
nand U16264 (N_16264,N_13013,N_11451);
and U16265 (N_16265,N_14390,N_10491);
nor U16266 (N_16266,N_11909,N_12214);
nor U16267 (N_16267,N_13132,N_11936);
nand U16268 (N_16268,N_12977,N_12856);
and U16269 (N_16269,N_12872,N_13311);
nand U16270 (N_16270,N_13120,N_11446);
nand U16271 (N_16271,N_11053,N_10038);
and U16272 (N_16272,N_12246,N_11408);
and U16273 (N_16273,N_11480,N_11999);
xnor U16274 (N_16274,N_10325,N_12869);
or U16275 (N_16275,N_11010,N_13286);
nor U16276 (N_16276,N_11489,N_12794);
and U16277 (N_16277,N_13488,N_11036);
xnor U16278 (N_16278,N_11615,N_12346);
nand U16279 (N_16279,N_12816,N_12625);
and U16280 (N_16280,N_12465,N_14764);
nor U16281 (N_16281,N_11347,N_10616);
xor U16282 (N_16282,N_10530,N_13184);
and U16283 (N_16283,N_12264,N_12299);
nor U16284 (N_16284,N_11069,N_14285);
xor U16285 (N_16285,N_12399,N_12367);
nand U16286 (N_16286,N_11836,N_14534);
nand U16287 (N_16287,N_13263,N_14602);
xnor U16288 (N_16288,N_14258,N_14106);
nand U16289 (N_16289,N_10109,N_13520);
nand U16290 (N_16290,N_12207,N_12938);
nand U16291 (N_16291,N_10601,N_13639);
nor U16292 (N_16292,N_14894,N_13837);
or U16293 (N_16293,N_12230,N_11602);
xor U16294 (N_16294,N_14807,N_13944);
or U16295 (N_16295,N_14626,N_11635);
and U16296 (N_16296,N_13396,N_10247);
nand U16297 (N_16297,N_11208,N_11393);
nand U16298 (N_16298,N_12581,N_14293);
or U16299 (N_16299,N_11178,N_11201);
nor U16300 (N_16300,N_13016,N_13602);
nor U16301 (N_16301,N_10757,N_13919);
xor U16302 (N_16302,N_13226,N_11724);
or U16303 (N_16303,N_11179,N_10344);
or U16304 (N_16304,N_14303,N_14080);
nand U16305 (N_16305,N_14335,N_11175);
xnor U16306 (N_16306,N_14784,N_14397);
or U16307 (N_16307,N_13235,N_13445);
nor U16308 (N_16308,N_10469,N_12267);
nand U16309 (N_16309,N_11272,N_10869);
xnor U16310 (N_16310,N_10460,N_11606);
nand U16311 (N_16311,N_11818,N_12932);
nor U16312 (N_16312,N_12040,N_13566);
and U16313 (N_16313,N_13208,N_11585);
nand U16314 (N_16314,N_13800,N_14817);
nand U16315 (N_16315,N_12324,N_14955);
xor U16316 (N_16316,N_11405,N_12485);
nor U16317 (N_16317,N_10391,N_11870);
and U16318 (N_16318,N_10554,N_11151);
or U16319 (N_16319,N_11397,N_14442);
nor U16320 (N_16320,N_11548,N_10261);
xnor U16321 (N_16321,N_10778,N_11743);
and U16322 (N_16322,N_12543,N_14399);
or U16323 (N_16323,N_11783,N_14248);
xnor U16324 (N_16324,N_11679,N_12614);
or U16325 (N_16325,N_11569,N_13040);
xor U16326 (N_16326,N_14929,N_12333);
and U16327 (N_16327,N_14619,N_12009);
nor U16328 (N_16328,N_14780,N_12257);
or U16329 (N_16329,N_12086,N_12744);
nor U16330 (N_16330,N_10760,N_10484);
and U16331 (N_16331,N_12349,N_11915);
xor U16332 (N_16332,N_12707,N_10374);
nor U16333 (N_16333,N_10447,N_11949);
nand U16334 (N_16334,N_11573,N_11192);
and U16335 (N_16335,N_12095,N_13378);
or U16336 (N_16336,N_13001,N_10552);
nand U16337 (N_16337,N_13478,N_10674);
nand U16338 (N_16338,N_12684,N_10407);
nand U16339 (N_16339,N_13910,N_10543);
or U16340 (N_16340,N_10186,N_12775);
xor U16341 (N_16341,N_14476,N_14064);
nor U16342 (N_16342,N_13597,N_11077);
nor U16343 (N_16343,N_11487,N_10917);
or U16344 (N_16344,N_13121,N_12014);
nand U16345 (N_16345,N_11620,N_14984);
nand U16346 (N_16346,N_12428,N_14511);
and U16347 (N_16347,N_12788,N_14048);
and U16348 (N_16348,N_10627,N_10476);
xnor U16349 (N_16349,N_13875,N_10507);
nor U16350 (N_16350,N_11279,N_14247);
xnor U16351 (N_16351,N_14433,N_12729);
nand U16352 (N_16352,N_11773,N_10931);
xor U16353 (N_16353,N_13553,N_11310);
xnor U16354 (N_16354,N_12334,N_14256);
or U16355 (N_16355,N_11609,N_12563);
or U16356 (N_16356,N_13036,N_14069);
and U16357 (N_16357,N_12046,N_14882);
nor U16358 (N_16358,N_11867,N_12594);
xnor U16359 (N_16359,N_14156,N_12914);
and U16360 (N_16360,N_12895,N_11511);
xor U16361 (N_16361,N_10563,N_11819);
or U16362 (N_16362,N_12080,N_13171);
or U16363 (N_16363,N_11524,N_10010);
nand U16364 (N_16364,N_10609,N_10269);
or U16365 (N_16365,N_12601,N_12228);
nor U16366 (N_16366,N_10956,N_14680);
or U16367 (N_16367,N_14109,N_11662);
xnor U16368 (N_16368,N_13827,N_11354);
nor U16369 (N_16369,N_11215,N_10275);
xor U16370 (N_16370,N_12774,N_14178);
or U16371 (N_16371,N_13280,N_14121);
or U16372 (N_16372,N_12409,N_10998);
nor U16373 (N_16373,N_14898,N_13050);
nor U16374 (N_16374,N_12554,N_13954);
and U16375 (N_16375,N_10217,N_14618);
nor U16376 (N_16376,N_14566,N_12736);
or U16377 (N_16377,N_14438,N_10020);
and U16378 (N_16378,N_10693,N_10425);
nand U16379 (N_16379,N_13246,N_13816);
nand U16380 (N_16380,N_14445,N_10379);
xnor U16381 (N_16381,N_11551,N_14698);
nand U16382 (N_16382,N_14295,N_11342);
xnor U16383 (N_16383,N_11360,N_10257);
and U16384 (N_16384,N_14071,N_10769);
or U16385 (N_16385,N_10288,N_11195);
nor U16386 (N_16386,N_12183,N_13856);
or U16387 (N_16387,N_14549,N_12690);
nor U16388 (N_16388,N_14450,N_12864);
or U16389 (N_16389,N_12646,N_12996);
and U16390 (N_16390,N_14489,N_11957);
and U16391 (N_16391,N_12303,N_14584);
nor U16392 (N_16392,N_14890,N_10031);
nand U16393 (N_16393,N_13172,N_11736);
nor U16394 (N_16394,N_12678,N_10411);
nor U16395 (N_16395,N_10429,N_13536);
nor U16396 (N_16396,N_13355,N_14427);
xnor U16397 (N_16397,N_12802,N_11475);
or U16398 (N_16398,N_14001,N_14077);
nor U16399 (N_16399,N_10198,N_10542);
nor U16400 (N_16400,N_12209,N_14931);
xor U16401 (N_16401,N_10734,N_14108);
nand U16402 (N_16402,N_14203,N_10147);
and U16403 (N_16403,N_14674,N_13216);
and U16404 (N_16404,N_10892,N_11019);
and U16405 (N_16405,N_13609,N_12287);
nor U16406 (N_16406,N_11441,N_10845);
or U16407 (N_16407,N_11274,N_14289);
and U16408 (N_16408,N_10388,N_11225);
nand U16409 (N_16409,N_12413,N_14216);
nor U16410 (N_16410,N_11518,N_14093);
nor U16411 (N_16411,N_11283,N_13062);
and U16412 (N_16412,N_11258,N_11716);
nor U16413 (N_16413,N_13279,N_12703);
nor U16414 (N_16414,N_13318,N_11599);
nand U16415 (N_16415,N_11790,N_11119);
nor U16416 (N_16416,N_13093,N_13976);
or U16417 (N_16417,N_13459,N_10424);
nand U16418 (N_16418,N_10365,N_14049);
xor U16419 (N_16419,N_13762,N_13292);
xor U16420 (N_16420,N_13662,N_11905);
xnor U16421 (N_16421,N_14677,N_13691);
nand U16422 (N_16422,N_10486,N_10249);
nand U16423 (N_16423,N_11778,N_10312);
xor U16424 (N_16424,N_11254,N_13814);
xor U16425 (N_16425,N_10129,N_12575);
nor U16426 (N_16426,N_10623,N_12094);
nand U16427 (N_16427,N_13303,N_12167);
nand U16428 (N_16428,N_11306,N_10725);
and U16429 (N_16429,N_13299,N_14982);
xnor U16430 (N_16430,N_11767,N_14960);
or U16431 (N_16431,N_10662,N_14969);
or U16432 (N_16432,N_14092,N_13109);
nor U16433 (N_16433,N_12158,N_13727);
or U16434 (N_16434,N_13505,N_11091);
and U16435 (N_16435,N_10622,N_13026);
nor U16436 (N_16436,N_14416,N_13869);
or U16437 (N_16437,N_11889,N_12919);
xor U16438 (N_16438,N_12949,N_12013);
nor U16439 (N_16439,N_10771,N_12862);
and U16440 (N_16440,N_10409,N_11692);
or U16441 (N_16441,N_14666,N_12870);
and U16442 (N_16442,N_10708,N_10468);
xnor U16443 (N_16443,N_12157,N_14865);
and U16444 (N_16444,N_14208,N_11099);
nand U16445 (N_16445,N_13399,N_13742);
nand U16446 (N_16446,N_13502,N_13223);
and U16447 (N_16447,N_10992,N_14689);
nand U16448 (N_16448,N_14292,N_11910);
and U16449 (N_16449,N_13958,N_13654);
nand U16450 (N_16450,N_11532,N_11432);
and U16451 (N_16451,N_11097,N_14425);
nor U16452 (N_16452,N_13626,N_10736);
or U16453 (N_16453,N_12991,N_12499);
nor U16454 (N_16454,N_10994,N_12098);
xor U16455 (N_16455,N_13181,N_12934);
and U16456 (N_16456,N_13967,N_14300);
xnor U16457 (N_16457,N_14857,N_14411);
nand U16458 (N_16458,N_11130,N_11782);
nand U16459 (N_16459,N_14192,N_11460);
and U16460 (N_16460,N_11415,N_13423);
xor U16461 (N_16461,N_11944,N_10047);
and U16462 (N_16462,N_13775,N_14751);
and U16463 (N_16463,N_11194,N_14360);
nand U16464 (N_16464,N_13630,N_14255);
or U16465 (N_16465,N_12100,N_13591);
and U16466 (N_16466,N_13063,N_13547);
and U16467 (N_16467,N_11245,N_14319);
nor U16468 (N_16468,N_13785,N_10056);
xor U16469 (N_16469,N_12898,N_14843);
and U16470 (N_16470,N_10974,N_14321);
and U16471 (N_16471,N_12845,N_12700);
nand U16472 (N_16472,N_13170,N_10984);
nand U16473 (N_16473,N_14060,N_11851);
nor U16474 (N_16474,N_13084,N_12347);
and U16475 (N_16475,N_13952,N_10185);
nor U16476 (N_16476,N_10787,N_12196);
nor U16477 (N_16477,N_11235,N_10611);
and U16478 (N_16478,N_11363,N_12362);
xor U16479 (N_16479,N_11598,N_14585);
xnor U16480 (N_16480,N_13943,N_14403);
nand U16481 (N_16481,N_11561,N_11536);
nand U16482 (N_16482,N_11402,N_11398);
or U16483 (N_16483,N_13331,N_10539);
or U16484 (N_16484,N_10385,N_12761);
and U16485 (N_16485,N_11406,N_13892);
and U16486 (N_16486,N_12147,N_14350);
nor U16487 (N_16487,N_11566,N_13402);
and U16488 (N_16488,N_13798,N_14129);
and U16489 (N_16489,N_10719,N_14794);
and U16490 (N_16490,N_14090,N_11065);
and U16491 (N_16491,N_14777,N_11627);
nor U16492 (N_16492,N_14055,N_14975);
nand U16493 (N_16493,N_11808,N_11742);
nor U16494 (N_16494,N_12076,N_14564);
or U16495 (N_16495,N_14190,N_11066);
and U16496 (N_16496,N_10216,N_14151);
xnor U16497 (N_16497,N_10512,N_11880);
or U16498 (N_16498,N_13508,N_11834);
or U16499 (N_16499,N_13153,N_14086);
nand U16500 (N_16500,N_14582,N_14063);
or U16501 (N_16501,N_12529,N_10600);
nand U16502 (N_16502,N_11048,N_13165);
xor U16503 (N_16503,N_11399,N_10309);
or U16504 (N_16504,N_14863,N_11332);
nor U16505 (N_16505,N_14832,N_10280);
nand U16506 (N_16506,N_14184,N_13673);
or U16507 (N_16507,N_10716,N_12964);
or U16508 (N_16508,N_14665,N_14828);
nor U16509 (N_16509,N_10737,N_10782);
and U16510 (N_16510,N_11746,N_14745);
nor U16511 (N_16511,N_14230,N_14805);
nand U16512 (N_16512,N_13365,N_11512);
and U16513 (N_16513,N_13764,N_13846);
nand U16514 (N_16514,N_13325,N_10377);
or U16515 (N_16515,N_12274,N_10370);
nand U16516 (N_16516,N_11864,N_11815);
or U16517 (N_16517,N_13437,N_14884);
nand U16518 (N_16518,N_14308,N_14362);
or U16519 (N_16519,N_14599,N_13698);
or U16520 (N_16520,N_14730,N_10696);
nand U16521 (N_16521,N_12827,N_13398);
and U16522 (N_16522,N_13570,N_13664);
xor U16523 (N_16523,N_12891,N_12161);
xor U16524 (N_16524,N_11714,N_13262);
and U16525 (N_16525,N_13605,N_11461);
nor U16526 (N_16526,N_11919,N_14088);
and U16527 (N_16527,N_13304,N_11831);
nor U16528 (N_16528,N_14338,N_13810);
nor U16529 (N_16529,N_13118,N_11428);
nand U16530 (N_16530,N_12002,N_10822);
or U16531 (N_16531,N_12101,N_10872);
nand U16532 (N_16532,N_14095,N_11509);
nand U16533 (N_16533,N_14926,N_12186);
or U16534 (N_16534,N_11951,N_13663);
xor U16535 (N_16535,N_12608,N_10122);
and U16536 (N_16536,N_14388,N_14126);
nand U16537 (N_16537,N_12450,N_13719);
and U16538 (N_16538,N_11450,N_13266);
xnor U16539 (N_16539,N_13503,N_14889);
nor U16540 (N_16540,N_11150,N_14218);
nor U16541 (N_16541,N_14174,N_13589);
or U16542 (N_16542,N_10382,N_13926);
and U16543 (N_16543,N_10180,N_10755);
and U16544 (N_16544,N_14141,N_11330);
and U16545 (N_16545,N_12405,N_11127);
xnor U16546 (N_16546,N_12314,N_12512);
xor U16547 (N_16547,N_13968,N_13329);
nor U16548 (N_16548,N_12899,N_11865);
xor U16549 (N_16549,N_10983,N_14194);
nand U16550 (N_16550,N_10919,N_12883);
and U16551 (N_16551,N_12240,N_12644);
xnor U16552 (N_16552,N_12481,N_13844);
and U16553 (N_16553,N_12569,N_13332);
xor U16554 (N_16554,N_12165,N_11200);
nand U16555 (N_16555,N_14477,N_14167);
or U16556 (N_16556,N_13010,N_11656);
xnor U16557 (N_16557,N_13422,N_12051);
or U16558 (N_16558,N_12745,N_10711);
xor U16559 (N_16559,N_10794,N_14631);
nand U16560 (N_16560,N_12611,N_13546);
and U16561 (N_16561,N_13278,N_12687);
nand U16562 (N_16562,N_12815,N_11256);
nor U16563 (N_16563,N_10904,N_14340);
nor U16564 (N_16564,N_14880,N_13644);
xnor U16565 (N_16565,N_13442,N_11541);
and U16566 (N_16566,N_10296,N_14829);
nand U16567 (N_16567,N_10797,N_13551);
nand U16568 (N_16568,N_14100,N_10763);
nand U16569 (N_16569,N_12108,N_14856);
xnor U16570 (N_16570,N_11812,N_11926);
and U16571 (N_16571,N_11228,N_12304);
nor U16572 (N_16572,N_11291,N_12195);
or U16573 (N_16573,N_13247,N_12476);
nand U16574 (N_16574,N_12954,N_14232);
xor U16575 (N_16575,N_12983,N_14557);
nor U16576 (N_16576,N_12000,N_11309);
or U16577 (N_16577,N_11372,N_12105);
or U16578 (N_16578,N_13327,N_13440);
or U16579 (N_16579,N_12837,N_14996);
xor U16580 (N_16580,N_10820,N_11733);
xor U16581 (N_16581,N_14954,N_14152);
xnor U16582 (N_16582,N_13222,N_11961);
nor U16583 (N_16583,N_13128,N_13014);
or U16584 (N_16584,N_11610,N_10619);
or U16585 (N_16585,N_11726,N_10330);
nor U16586 (N_16586,N_13571,N_11147);
or U16587 (N_16587,N_14004,N_10139);
nor U16588 (N_16588,N_14453,N_10989);
and U16589 (N_16589,N_14471,N_14765);
nand U16590 (N_16590,N_10371,N_11391);
xnor U16591 (N_16591,N_14738,N_11988);
and U16592 (N_16592,N_14091,N_12242);
xnor U16593 (N_16593,N_13594,N_11046);
nand U16594 (N_16594,N_10752,N_14323);
and U16595 (N_16595,N_10044,N_13981);
xnor U16596 (N_16596,N_14139,N_13168);
and U16597 (N_16597,N_10824,N_11469);
and U16598 (N_16598,N_14945,N_12933);
and U16599 (N_16599,N_13695,N_12812);
and U16600 (N_16600,N_13164,N_14493);
nor U16601 (N_16601,N_12971,N_12188);
nor U16602 (N_16602,N_14571,N_12782);
or U16603 (N_16603,N_12508,N_11932);
nor U16604 (N_16604,N_11800,N_10300);
and U16605 (N_16605,N_11866,N_14357);
xnor U16606 (N_16606,N_11125,N_13871);
nor U16607 (N_16607,N_11531,N_12373);
nor U16608 (N_16608,N_10547,N_13267);
nand U16609 (N_16609,N_14263,N_13562);
xnor U16610 (N_16610,N_12545,N_10342);
xnor U16611 (N_16611,N_12289,N_14506);
or U16612 (N_16612,N_13186,N_10079);
xnor U16613 (N_16613,N_10252,N_13066);
nand U16614 (N_16614,N_14150,N_14923);
nand U16615 (N_16615,N_14098,N_13054);
nand U16616 (N_16616,N_11997,N_12366);
xnor U16617 (N_16617,N_12272,N_13159);
or U16618 (N_16618,N_14568,N_10649);
and U16619 (N_16619,N_10935,N_12270);
nor U16620 (N_16620,N_14305,N_10078);
nor U16621 (N_16621,N_13567,N_14130);
nand U16622 (N_16622,N_13634,N_14015);
nor U16623 (N_16623,N_13915,N_13690);
nand U16624 (N_16624,N_12276,N_12951);
and U16625 (N_16625,N_13830,N_14968);
xor U16626 (N_16626,N_11987,N_14875);
nor U16627 (N_16627,N_14217,N_10858);
and U16628 (N_16628,N_10541,N_10118);
and U16629 (N_16629,N_13569,N_11251);
xor U16630 (N_16630,N_14686,N_13819);
and U16631 (N_16631,N_12422,N_10729);
or U16632 (N_16632,N_13464,N_11695);
xor U16633 (N_16633,N_10372,N_10239);
or U16634 (N_16634,N_11520,N_12113);
nand U16635 (N_16635,N_12336,N_14466);
nor U16636 (N_16636,N_14925,N_12459);
xor U16637 (N_16637,N_13558,N_11748);
nor U16638 (N_16638,N_12379,N_14117);
nor U16639 (N_16639,N_12841,N_13388);
xor U16640 (N_16640,N_13403,N_13358);
and U16641 (N_16641,N_11528,N_13408);
and U16642 (N_16642,N_13575,N_12935);
or U16643 (N_16643,N_13383,N_12331);
xnor U16644 (N_16644,N_10473,N_10566);
and U16645 (N_16645,N_13578,N_10004);
and U16646 (N_16646,N_10599,N_13053);
nand U16647 (N_16647,N_14778,N_11492);
and U16648 (N_16648,N_10587,N_13606);
or U16649 (N_16649,N_12580,N_13636);
nand U16650 (N_16650,N_10745,N_11341);
and U16651 (N_16651,N_11034,N_11135);
xor U16652 (N_16652,N_11530,N_10859);
nor U16653 (N_16653,N_11311,N_14265);
xor U16654 (N_16654,N_13143,N_10690);
and U16655 (N_16655,N_11847,N_10952);
nand U16656 (N_16656,N_11796,N_13736);
or U16657 (N_16657,N_13351,N_11174);
nand U16658 (N_16658,N_11358,N_10157);
xor U16659 (N_16659,N_12871,N_13864);
xnor U16660 (N_16660,N_10489,N_14684);
and U16661 (N_16661,N_12136,N_12226);
xor U16662 (N_16662,N_14116,N_14578);
xor U16663 (N_16663,N_14789,N_12587);
nand U16664 (N_16664,N_13284,N_10926);
xnor U16665 (N_16665,N_14236,N_12667);
xnor U16666 (N_16666,N_11260,N_10211);
nor U16667 (N_16667,N_14025,N_12348);
nand U16668 (N_16668,N_10427,N_12054);
or U16669 (N_16669,N_14318,N_12591);
and U16670 (N_16670,N_14102,N_11722);
nand U16671 (N_16671,N_12259,N_13833);
or U16672 (N_16672,N_12890,N_14913);
nand U16673 (N_16673,N_13651,N_14131);
nand U16674 (N_16674,N_11603,N_10957);
xnor U16675 (N_16675,N_13542,N_11632);
or U16676 (N_16676,N_10302,N_11614);
nor U16677 (N_16677,N_14989,N_11485);
and U16678 (N_16678,N_12820,N_11704);
xnor U16679 (N_16679,N_10253,N_11967);
nor U16680 (N_16680,N_13794,N_14757);
and U16681 (N_16681,N_14112,N_14491);
or U16682 (N_16682,N_11218,N_12496);
and U16683 (N_16683,N_13088,N_11250);
nor U16684 (N_16684,N_10518,N_14554);
nor U16685 (N_16685,N_13513,N_11619);
xnor U16686 (N_16686,N_12642,N_13983);
xnor U16687 (N_16687,N_12433,N_13874);
nor U16688 (N_16688,N_12069,N_10317);
or U16689 (N_16689,N_10162,N_13714);
nand U16690 (N_16690,N_14214,N_10283);
xnor U16691 (N_16691,N_12830,N_10495);
xnor U16692 (N_16692,N_12902,N_11522);
or U16693 (N_16693,N_11622,N_12256);
nor U16694 (N_16694,N_11156,N_13559);
nor U16695 (N_16695,N_11542,N_11126);
nor U16696 (N_16696,N_14693,N_13623);
nand U16697 (N_16697,N_14746,N_11553);
nor U16698 (N_16698,N_11660,N_11129);
and U16699 (N_16699,N_14706,N_12661);
nor U16700 (N_16700,N_10726,N_11140);
or U16701 (N_16701,N_10633,N_14900);
and U16702 (N_16702,N_14768,N_11617);
or U16703 (N_16703,N_14484,N_13167);
nor U16704 (N_16704,N_10406,N_13103);
xnor U16705 (N_16705,N_14712,N_11618);
or U16706 (N_16706,N_14724,N_12041);
or U16707 (N_16707,N_14510,N_13227);
and U16708 (N_16708,N_12865,N_14736);
or U16709 (N_16709,N_10695,N_12536);
or U16710 (N_16710,N_14878,N_14512);
nand U16711 (N_16711,N_13473,N_10659);
or U16712 (N_16712,N_12551,N_10040);
nand U16713 (N_16713,N_13720,N_14668);
nand U16714 (N_16714,N_13861,N_10015);
nor U16715 (N_16715,N_14257,N_12150);
or U16716 (N_16716,N_11993,N_10875);
nor U16717 (N_16717,N_10172,N_11578);
xor U16718 (N_16718,N_13608,N_12645);
or U16719 (N_16719,N_11516,N_13260);
or U16720 (N_16720,N_14509,N_11527);
and U16721 (N_16721,N_12393,N_12868);
nand U16722 (N_16722,N_12106,N_12833);
nor U16723 (N_16723,N_12709,N_10620);
nor U16724 (N_16724,N_12850,N_14716);
nor U16725 (N_16725,N_10069,N_10865);
xor U16726 (N_16726,N_10046,N_13845);
or U16727 (N_16727,N_12852,N_10551);
nor U16728 (N_16728,N_11925,N_12288);
and U16729 (N_16729,N_14373,N_11072);
xnor U16730 (N_16730,N_12385,N_11794);
nor U16731 (N_16731,N_14065,N_13375);
or U16732 (N_16732,N_13813,N_11315);
and U16733 (N_16733,N_12859,N_12676);
or U16734 (N_16734,N_12924,N_10738);
nor U16735 (N_16735,N_11908,N_13413);
and U16736 (N_16736,N_10165,N_14358);
and U16737 (N_16737,N_10254,N_11821);
or U16738 (N_16738,N_11994,N_10891);
nand U16739 (N_16739,N_10474,N_11325);
nor U16740 (N_16740,N_14153,N_10001);
nor U16741 (N_16741,N_11264,N_13504);
xnor U16742 (N_16742,N_10331,N_11064);
nor U16743 (N_16743,N_12521,N_14497);
or U16744 (N_16744,N_13295,N_13953);
xor U16745 (N_16745,N_11678,N_12026);
and U16746 (N_16746,N_13043,N_11362);
or U16747 (N_16747,N_10920,N_14143);
xor U16748 (N_16748,N_11881,N_11753);
xor U16749 (N_16749,N_10445,N_10265);
xnor U16750 (N_16750,N_10533,N_10285);
nor U16751 (N_16751,N_14744,N_13831);
xor U16752 (N_16752,N_14436,N_12691);
nor U16753 (N_16753,N_13599,N_12732);
nand U16754 (N_16754,N_11183,N_13276);
or U16755 (N_16755,N_11639,N_13083);
nand U16756 (N_16756,N_10641,N_14687);
or U16757 (N_16757,N_14523,N_12957);
nand U16758 (N_16758,N_12107,N_14934);
nand U16759 (N_16759,N_12878,N_11434);
nor U16760 (N_16760,N_13347,N_12164);
or U16761 (N_16761,N_10212,N_11623);
and U16762 (N_16762,N_14118,N_13409);
nor U16763 (N_16763,N_12542,N_10647);
nand U16764 (N_16764,N_14691,N_12480);
or U16765 (N_16765,N_12626,N_13607);
nor U16766 (N_16766,N_13828,N_12881);
and U16767 (N_16767,N_11420,N_14467);
nor U16768 (N_16768,N_13460,N_13994);
xor U16769 (N_16769,N_13659,N_12425);
or U16770 (N_16770,N_10376,N_11383);
xnor U16771 (N_16771,N_14891,N_12162);
or U16772 (N_16772,N_13394,N_13474);
nor U16773 (N_16773,N_12785,N_11165);
nor U16774 (N_16774,N_11246,N_12538);
or U16775 (N_16775,N_12215,N_13191);
nor U16776 (N_16776,N_10975,N_11164);
and U16777 (N_16777,N_11285,N_11138);
nor U16778 (N_16778,N_11314,N_13081);
and U16779 (N_16779,N_11937,N_14456);
or U16780 (N_16780,N_10746,N_11088);
nand U16781 (N_16781,N_12909,N_11243);
nor U16782 (N_16782,N_14897,N_10675);
or U16783 (N_16783,N_13787,N_14301);
nand U16784 (N_16784,N_14836,N_11400);
nand U16785 (N_16785,N_11756,N_12602);
nand U16786 (N_16786,N_10772,N_10410);
xor U16787 (N_16787,N_10826,N_12911);
xor U16788 (N_16788,N_10982,N_12079);
and U16789 (N_16789,N_14430,N_10885);
xnor U16790 (N_16790,N_10158,N_10976);
nor U16791 (N_16791,N_11750,N_12369);
nand U16792 (N_16792,N_10228,N_10852);
nor U16793 (N_16793,N_12477,N_11144);
or U16794 (N_16794,N_12931,N_14009);
and U16795 (N_16795,N_13316,N_14520);
and U16796 (N_16796,N_12386,N_11839);
or U16797 (N_16797,N_10618,N_12444);
nand U16798 (N_16798,N_12874,N_11501);
and U16799 (N_16799,N_13430,N_12163);
nor U16800 (N_16800,N_11163,N_10894);
nor U16801 (N_16801,N_13157,N_12039);
and U16802 (N_16802,N_10569,N_10003);
and U16803 (N_16803,N_10098,N_12397);
nor U16804 (N_16804,N_13935,N_13158);
nor U16805 (N_16805,N_13956,N_13581);
nor U16806 (N_16806,N_12805,N_14437);
nand U16807 (N_16807,N_12068,N_10128);
nor U16808 (N_16808,N_13368,N_13091);
nor U16809 (N_16809,N_14651,N_11259);
and U16810 (N_16810,N_12458,N_12522);
nand U16811 (N_16811,N_12227,N_14235);
xnor U16812 (N_16812,N_10560,N_11638);
or U16813 (N_16813,N_10096,N_10747);
or U16814 (N_16814,N_10642,N_11189);
xor U16815 (N_16815,N_11149,N_10316);
nand U16816 (N_16816,N_14567,N_13693);
and U16817 (N_16817,N_11992,N_10206);
or U16818 (N_16818,N_12576,N_10773);
nor U16819 (N_16819,N_10471,N_10731);
or U16820 (N_16820,N_10574,N_10842);
xnor U16821 (N_16821,N_12421,N_12427);
nand U16822 (N_16822,N_14950,N_12523);
or U16823 (N_16823,N_11490,N_12984);
nor U16824 (N_16824,N_10338,N_14182);
nor U16825 (N_16825,N_14983,N_10494);
or U16826 (N_16826,N_10501,N_12752);
nand U16827 (N_16827,N_11094,N_10866);
nor U16828 (N_16828,N_10071,N_13793);
nor U16829 (N_16829,N_13339,N_12056);
or U16830 (N_16830,N_10978,N_10519);
nand U16831 (N_16831,N_14940,N_10950);
and U16832 (N_16832,N_14592,N_10968);
nor U16833 (N_16833,N_14457,N_10831);
nor U16834 (N_16834,N_14026,N_10856);
and U16835 (N_16835,N_14577,N_14031);
or U16836 (N_16836,N_10195,N_13684);
nand U16837 (N_16837,N_12199,N_13674);
and U16838 (N_16838,N_14797,N_11008);
nand U16839 (N_16839,N_11798,N_14033);
nand U16840 (N_16840,N_12948,N_11212);
xor U16841 (N_16841,N_14379,N_10873);
or U16842 (N_16842,N_11176,N_14886);
nor U16843 (N_16843,N_11680,N_11899);
and U16844 (N_16844,N_10793,N_10073);
nand U16845 (N_16845,N_11669,N_13051);
nor U16846 (N_16846,N_13731,N_10877);
and U16847 (N_16847,N_13730,N_13136);
xnor U16848 (N_16848,N_11233,N_12019);
nand U16849 (N_16849,N_10470,N_10679);
nand U16850 (N_16850,N_13635,N_14538);
xor U16851 (N_16851,N_10591,N_10323);
xor U16852 (N_16852,N_12624,N_10135);
nor U16853 (N_16853,N_10164,N_11426);
xnor U16854 (N_16854,N_13435,N_11776);
nand U16855 (N_16855,N_11942,N_10168);
xor U16856 (N_16856,N_13999,N_14756);
or U16857 (N_16857,N_14846,N_12117);
nor U16858 (N_16858,N_10779,N_14157);
xnor U16859 (N_16859,N_12544,N_14082);
xor U16860 (N_16860,N_12534,N_11386);
nor U16861 (N_16861,N_14622,N_14356);
nor U16862 (N_16862,N_12127,N_10657);
nor U16863 (N_16863,N_10838,N_14309);
nand U16864 (N_16864,N_12204,N_12928);
nor U16865 (N_16865,N_14732,N_12306);
nor U16866 (N_16866,N_10373,N_13721);
or U16867 (N_16867,N_14546,N_14173);
nand U16868 (N_16868,N_12814,N_10025);
nand U16869 (N_16869,N_11351,N_10125);
and U16870 (N_16870,N_10294,N_10565);
and U16871 (N_16871,N_12976,N_11912);
xor U16872 (N_16872,N_13500,N_12715);
and U16873 (N_16873,N_10235,N_10260);
xnor U16874 (N_16874,N_10037,N_11244);
nand U16875 (N_16875,N_14853,N_11413);
nand U16876 (N_16876,N_11288,N_12818);
nor U16877 (N_16877,N_12500,N_13185);
nor U16878 (N_16878,N_11079,N_11681);
nor U16879 (N_16879,N_13518,N_13511);
xnor U16880 (N_16880,N_12492,N_13836);
xor U16881 (N_16881,N_11051,N_13224);
xnor U16882 (N_16882,N_12747,N_10971);
nor U16883 (N_16883,N_11193,N_11190);
or U16884 (N_16884,N_12930,N_12001);
nor U16885 (N_16885,N_11473,N_11725);
and U16886 (N_16886,N_13807,N_10846);
nor U16887 (N_16887,N_12887,N_13535);
nand U16888 (N_16888,N_13073,N_14775);
nand U16889 (N_16889,N_14146,N_11329);
xor U16890 (N_16890,N_14986,N_14961);
and U16891 (N_16891,N_10867,N_13909);
nand U16892 (N_16892,N_10400,N_10291);
or U16893 (N_16893,N_13914,N_13921);
or U16894 (N_16894,N_10326,N_13525);
xor U16895 (N_16895,N_10617,N_11452);
nand U16896 (N_16896,N_10245,N_11752);
nand U16897 (N_16897,N_10864,N_10670);
xor U16898 (N_16898,N_10753,N_13369);
nor U16899 (N_16899,N_14089,N_12777);
or U16900 (N_16900,N_10262,N_11445);
or U16901 (N_16901,N_14045,N_14042);
nand U16902 (N_16902,N_11557,N_14268);
xnor U16903 (N_16903,N_12737,N_11549);
nor U16904 (N_16904,N_10508,N_10765);
nor U16905 (N_16905,N_13348,N_11628);
nor U16906 (N_16906,N_12831,N_12290);
or U16907 (N_16907,N_13200,N_11412);
xnor U16908 (N_16908,N_13251,N_14395);
xor U16909 (N_16909,N_14251,N_11115);
and U16910 (N_16910,N_13907,N_12630);
nor U16911 (N_16911,N_10506,N_11647);
and U16912 (N_16912,N_14749,N_14294);
nand U16913 (N_16913,N_12265,N_11842);
nor U16914 (N_16914,N_11698,N_11238);
nor U16915 (N_16915,N_14169,N_12509);
nor U16916 (N_16916,N_14593,N_14315);
nand U16917 (N_16917,N_10899,N_13151);
nand U16918 (N_16918,N_11677,N_11184);
xnor U16919 (N_16919,N_12566,N_14610);
or U16920 (N_16920,N_14316,N_13028);
or U16921 (N_16921,N_12007,N_14123);
nor U16922 (N_16922,N_10336,N_14210);
and U16923 (N_16923,N_10967,N_11754);
nand U16924 (N_16924,N_11996,N_12980);
and U16925 (N_16925,N_13851,N_13767);
and U16926 (N_16926,N_10986,N_13458);
and U16927 (N_16927,N_13812,N_12138);
or U16928 (N_16928,N_13595,N_12011);
or U16929 (N_16929,N_13374,N_10857);
and U16930 (N_16930,N_10703,N_14016);
or U16931 (N_16931,N_11646,N_13995);
nand U16932 (N_16932,N_14558,N_10140);
or U16933 (N_16933,N_14539,N_13481);
xnor U16934 (N_16934,N_12390,N_11340);
and U16935 (N_16935,N_14723,N_10572);
nand U16936 (N_16936,N_14264,N_13586);
or U16937 (N_16937,N_14854,N_14107);
nand U16938 (N_16938,N_13089,N_14615);
and U16939 (N_16939,N_14132,N_14177);
or U16940 (N_16940,N_14697,N_14392);
nand U16941 (N_16941,N_10854,N_12792);
and U16942 (N_16942,N_11483,N_11160);
nor U16943 (N_16943,N_14527,N_14424);
xnor U16944 (N_16944,N_13669,N_11307);
or U16945 (N_16945,N_12894,N_14219);
nor U16946 (N_16946,N_10880,N_14137);
nand U16947 (N_16947,N_14815,N_14020);
nor U16948 (N_16948,N_12269,N_14727);
xor U16949 (N_16949,N_11761,N_10451);
nor U16950 (N_16950,N_10932,N_14287);
and U16951 (N_16951,N_12292,N_13625);
nor U16952 (N_16952,N_14324,N_14483);
or U16953 (N_16953,N_12124,N_10224);
xor U16954 (N_16954,N_14396,N_11765);
xor U16955 (N_16955,N_12152,N_13672);
nand U16956 (N_16956,N_11580,N_13984);
xnor U16957 (N_16957,N_10117,N_14076);
nand U16958 (N_16958,N_12061,N_12142);
or U16959 (N_16959,N_11320,N_11110);
nor U16960 (N_16960,N_10683,N_14791);
and U16961 (N_16961,N_12988,N_12131);
and U16962 (N_16962,N_11874,N_10684);
or U16963 (N_16963,N_13753,N_10478);
nand U16964 (N_16964,N_14647,N_10233);
xor U16965 (N_16965,N_12111,N_12143);
nor U16966 (N_16966,N_10292,N_10131);
nand U16967 (N_16967,N_14104,N_13244);
nor U16968 (N_16968,N_10363,N_12851);
nand U16969 (N_16969,N_14632,N_12302);
nand U16970 (N_16970,N_10455,N_12453);
xnor U16971 (N_16971,N_10638,N_12434);
nand U16972 (N_16972,N_12462,N_12972);
and U16973 (N_16973,N_11959,N_10792);
nor U16974 (N_16974,N_13792,N_14017);
xor U16975 (N_16975,N_12357,N_13763);
and U16976 (N_16976,N_11022,N_12692);
xnor U16977 (N_16977,N_10669,N_10510);
xor U16978 (N_16978,N_12178,N_14612);
nor U16979 (N_16979,N_14310,N_11586);
or U16980 (N_16980,N_13183,N_12099);
nand U16981 (N_16981,N_11885,N_12489);
and U16982 (N_16982,N_10761,N_14022);
or U16983 (N_16983,N_13631,N_10218);
and U16984 (N_16984,N_11131,N_12913);
xor U16985 (N_16985,N_11667,N_14628);
or U16986 (N_16986,N_10039,N_12245);
nand U16987 (N_16987,N_12717,N_11448);
nand U16988 (N_16988,N_11537,N_13832);
and U16989 (N_16989,N_13415,N_10665);
xnor U16990 (N_16990,N_11170,N_12710);
nand U16991 (N_16991,N_14369,N_10461);
nor U16992 (N_16992,N_12236,N_13854);
and U16993 (N_16993,N_14162,N_10184);
nor U16994 (N_16994,N_12918,N_10255);
nand U16995 (N_16995,N_10868,N_12048);
or U16996 (N_16996,N_10514,N_13071);
xor U16997 (N_16997,N_11276,N_13233);
nand U16998 (N_16998,N_10890,N_12478);
nor U16999 (N_16999,N_13797,N_12088);
and U17000 (N_17000,N_14096,N_11792);
nor U17001 (N_17001,N_10305,N_14490);
nand U17002 (N_17002,N_12469,N_10361);
and U17003 (N_17003,N_12846,N_14753);
or U17004 (N_17004,N_12583,N_12365);
or U17005 (N_17005,N_13042,N_14987);
or U17006 (N_17006,N_12635,N_11525);
and U17007 (N_17007,N_12074,N_13506);
or U17008 (N_17008,N_10236,N_14325);
nor U17009 (N_17009,N_13321,N_14937);
xor U17010 (N_17010,N_12377,N_13549);
or U17011 (N_17011,N_11768,N_10242);
nand U17012 (N_17012,N_10809,N_10843);
and U17013 (N_17013,N_14432,N_13337);
or U17014 (N_17014,N_13841,N_14448);
nand U17015 (N_17015,N_14414,N_13175);
nor U17016 (N_17016,N_10107,N_12416);
and U17017 (N_17017,N_11172,N_12858);
nor U17018 (N_17018,N_10434,N_12627);
xnor U17019 (N_17019,N_11423,N_12155);
nand U17020 (N_17020,N_13057,N_11075);
xor U17021 (N_17021,N_11058,N_14535);
or U17022 (N_17022,N_13512,N_11625);
xnor U17023 (N_17023,N_14165,N_12179);
nor U17024 (N_17024,N_11727,N_13778);
or U17025 (N_17025,N_11833,N_13293);
nor U17026 (N_17026,N_14907,N_12361);
nor U17027 (N_17027,N_10452,N_12823);
nor U17028 (N_17028,N_13152,N_14032);
nand U17029 (N_17029,N_12694,N_11965);
and U17030 (N_17030,N_12616,N_10688);
xor U17031 (N_17031,N_12929,N_12613);
or U17032 (N_17032,N_12514,N_10951);
nor U17033 (N_17033,N_11055,N_14561);
xor U17034 (N_17034,N_13434,N_13482);
nand U17035 (N_17035,N_12006,N_11349);
and U17036 (N_17036,N_14426,N_10201);
nor U17037 (N_17037,N_10266,N_11465);
or U17038 (N_17038,N_12381,N_13839);
and U17039 (N_17039,N_12555,N_10948);
and U17040 (N_17040,N_12210,N_13027);
nor U17041 (N_17041,N_11611,N_14259);
and U17042 (N_17042,N_13879,N_13485);
nand U17043 (N_17043,N_12946,N_10613);
nand U17044 (N_17044,N_10524,N_13842);
or U17045 (N_17045,N_10871,N_12746);
xor U17046 (N_17046,N_13471,N_14700);
and U17047 (N_17047,N_12319,N_12112);
xor U17048 (N_17048,N_12965,N_10496);
or U17049 (N_17049,N_12824,N_11817);
and U17050 (N_17050,N_10418,N_11220);
xor U17051 (N_17051,N_14097,N_14334);
or U17052 (N_17052,N_10698,N_13692);
or U17053 (N_17053,N_11040,N_14079);
or U17054 (N_17054,N_11508,N_13475);
and U17055 (N_17055,N_10353,N_13560);
nor U17056 (N_17056,N_13354,N_13288);
nand U17057 (N_17057,N_14161,N_12389);
and U17058 (N_17058,N_14896,N_14376);
and U17059 (N_17059,N_14220,N_13135);
and U17060 (N_17060,N_13646,N_12686);
nor U17061 (N_17061,N_14951,N_12997);
xor U17062 (N_17062,N_11223,N_13744);
or U17063 (N_17063,N_14037,N_10482);
xor U17064 (N_17064,N_13479,N_11335);
and U17065 (N_17065,N_12967,N_13916);
and U17066 (N_17066,N_14976,N_13190);
nor U17067 (N_17067,N_10043,N_14575);
xnor U17068 (N_17068,N_10925,N_14473);
and U17069 (N_17069,N_10961,N_13540);
and U17070 (N_17070,N_10907,N_13557);
or U17071 (N_17071,N_11788,N_11045);
and U17072 (N_17072,N_13718,N_12766);
xnor U17073 (N_17073,N_11702,N_14482);
or U17074 (N_17074,N_13697,N_12328);
nand U17075 (N_17075,N_11642,N_14662);
xor U17076 (N_17076,N_10256,N_14932);
xnor U17077 (N_17077,N_11844,N_13519);
nor U17078 (N_17078,N_12861,N_11100);
and U17079 (N_17079,N_11352,N_12572);
xor U17080 (N_17080,N_11626,N_12756);
nand U17081 (N_17081,N_14148,N_13847);
or U17082 (N_17082,N_11570,N_11004);
and U17083 (N_17083,N_12322,N_10000);
nand U17084 (N_17084,N_11943,N_10663);
and U17085 (N_17085,N_11629,N_13610);
and U17086 (N_17086,N_13979,N_13970);
nand U17087 (N_17087,N_10108,N_11804);
xor U17088 (N_17088,N_11297,N_13872);
and U17089 (N_17089,N_11846,N_13556);
and U17090 (N_17090,N_11688,N_10723);
nand U17091 (N_17091,N_13338,N_13738);
and U17092 (N_17092,N_14683,N_12621);
or U17093 (N_17093,N_12194,N_11824);
xnor U17094 (N_17094,N_13733,N_13255);
or U17095 (N_17095,N_11338,N_11799);
xor U17096 (N_17096,N_13087,N_13802);
xnor U17097 (N_17097,N_14560,N_13343);
nor U17098 (N_17098,N_11466,N_13613);
xor U17099 (N_17099,N_12973,N_14435);
or U17100 (N_17100,N_13015,N_14761);
or U17101 (N_17101,N_13598,N_13372);
xor U17102 (N_17102,N_11558,N_10116);
or U17103 (N_17103,N_14796,N_12789);
nand U17104 (N_17104,N_10914,N_13563);
or U17105 (N_17105,N_13033,N_13760);
xnor U17106 (N_17106,N_14441,N_13225);
nand U17107 (N_17107,N_14330,N_14785);
xnor U17108 (N_17108,N_10458,N_13925);
nor U17109 (N_17109,N_13773,N_12446);
or U17110 (N_17110,N_11567,N_11991);
nor U17111 (N_17111,N_14050,N_14870);
xor U17112 (N_17112,N_13204,N_11455);
nand U17113 (N_17113,N_12203,N_13144);
nand U17114 (N_17114,N_14291,N_14072);
nor U17115 (N_17115,N_14755,N_10742);
xor U17116 (N_17116,N_14094,N_11984);
nor U17117 (N_17117,N_10589,N_14672);
xor U17118 (N_17118,N_10750,N_13210);
and U17119 (N_17119,N_12415,N_10668);
xnor U17120 (N_17120,N_12574,N_10702);
nor U17121 (N_17121,N_10341,N_14168);
or U17122 (N_17122,N_13006,N_11922);
xnor U17123 (N_17123,N_11574,N_14646);
xor U17124 (N_17124,N_10946,N_13715);
and U17125 (N_17125,N_14820,N_14313);
and U17126 (N_17126,N_10464,N_12558);
nand U17127 (N_17127,N_11478,N_10881);
xnor U17128 (N_17128,N_11806,N_11416);
and U17129 (N_17129,N_12294,N_12201);
nand U17130 (N_17130,N_14822,N_13543);
nand U17131 (N_17131,N_13349,N_10840);
nand U17132 (N_17132,N_11484,N_13319);
and U17133 (N_17133,N_11180,N_13096);
or U17134 (N_17134,N_13261,N_11375);
xnor U17135 (N_17135,N_12243,N_10902);
nor U17136 (N_17136,N_12058,N_12518);
nor U17137 (N_17137,N_14249,N_12479);
nand U17138 (N_17138,N_10182,N_13300);
xnor U17139 (N_17139,N_11167,N_13933);
and U17140 (N_17140,N_14801,N_13037);
and U17141 (N_17141,N_12368,N_14660);
xnor U17142 (N_17142,N_10297,N_11430);
nor U17143 (N_17143,N_11876,N_10196);
nand U17144 (N_17144,N_11102,N_14588);
nand U17145 (N_17145,N_10900,N_12078);
or U17146 (N_17146,N_14478,N_12426);
xnor U17147 (N_17147,N_12634,N_11009);
and U17148 (N_17148,N_12232,N_10888);
or U17149 (N_17149,N_14873,N_12082);
nand U17150 (N_17150,N_12408,N_11387);
nor U17151 (N_17151,N_14522,N_11700);
or U17152 (N_17152,N_14695,N_14966);
or U17153 (N_17153,N_13648,N_12454);
xor U17154 (N_17154,N_10102,N_13972);
xnor U17155 (N_17155,N_11232,N_14743);
or U17156 (N_17156,N_10042,N_12547);
xor U17157 (N_17157,N_12151,N_12779);
nand U17158 (N_17158,N_11249,N_10475);
xor U17159 (N_17159,N_11459,N_12488);
nand U17160 (N_17160,N_13130,N_13061);
nand U17161 (N_17161,N_14888,N_13189);
nand U17162 (N_17162,N_13840,N_10050);
nor U17163 (N_17163,N_11838,N_12912);
nor U17164 (N_17164,N_12771,N_11852);
or U17165 (N_17165,N_10279,N_11443);
and U17166 (N_17166,N_12033,N_14431);
xnor U17167 (N_17167,N_10013,N_11803);
nand U17168 (N_17168,N_11476,N_11955);
nor U17169 (N_17169,N_12021,N_12623);
and U17170 (N_17170,N_11128,N_10993);
nor U17171 (N_17171,N_13315,N_11579);
nand U17172 (N_17172,N_13452,N_12337);
and U17173 (N_17173,N_10561,N_10273);
nand U17174 (N_17174,N_10806,N_14171);
or U17175 (N_17175,N_11685,N_12975);
nand U17176 (N_17176,N_14128,N_11482);
nor U17177 (N_17177,N_10340,N_11033);
nand U17178 (N_17178,N_13650,N_14087);
or U17179 (N_17179,N_14371,N_13532);
and U17180 (N_17180,N_12504,N_10219);
or U17181 (N_17181,N_12515,N_10150);
nand U17182 (N_17182,N_10329,N_14920);
nor U17183 (N_17183,N_13180,N_14879);
nor U17184 (N_17184,N_12517,N_13912);
nor U17185 (N_17185,N_10712,N_11650);
and U17186 (N_17186,N_11962,N_12726);
nand U17187 (N_17187,N_10979,N_13231);
nor U17188 (N_17188,N_11217,N_13993);
nand U17189 (N_17189,N_13786,N_14058);
nor U17190 (N_17190,N_14481,N_13901);
or U17191 (N_17191,N_12273,N_14124);
or U17192 (N_17192,N_10456,N_14449);
nor U17193 (N_17193,N_14899,N_12172);
nor U17194 (N_17194,N_14231,N_10807);
xnor U17195 (N_17195,N_14573,N_13272);
or U17196 (N_17196,N_14770,N_11409);
nand U17197 (N_17197,N_14754,N_14233);
nor U17198 (N_17198,N_10911,N_12182);
nor U17199 (N_17199,N_10727,N_12463);
and U17200 (N_17200,N_13366,N_13758);
xnor U17201 (N_17201,N_10485,N_12584);
or U17202 (N_17202,N_10800,N_11589);
nand U17203 (N_17203,N_13237,N_10005);
and U17204 (N_17204,N_10221,N_11116);
or U17205 (N_17205,N_12441,N_12171);
or U17206 (N_17206,N_12567,N_13699);
nor U17207 (N_17207,N_14221,N_12109);
and U17208 (N_17208,N_13728,N_11953);
nor U17209 (N_17209,N_11417,N_13885);
nand U17210 (N_17210,N_12768,N_13032);
xor U17211 (N_17211,N_12721,N_14949);
nand U17212 (N_17212,N_14633,N_12880);
and U17213 (N_17213,N_10054,N_12059);
and U17214 (N_17214,N_11162,N_12589);
nor U17215 (N_17215,N_11546,N_10133);
and U17216 (N_17216,N_11041,N_11708);
xor U17217 (N_17217,N_14530,N_12811);
or U17218 (N_17218,N_10938,N_13712);
or U17219 (N_17219,N_11098,N_14827);
and U17220 (N_17220,N_10562,N_14752);
and U17221 (N_17221,N_12075,N_10828);
nand U17222 (N_17222,N_12110,N_11273);
or U17223 (N_17223,N_13985,N_13405);
nor U17224 (N_17224,N_13629,N_12609);
nand U17225 (N_17225,N_10509,N_10011);
xnor U17226 (N_17226,N_10345,N_11979);
xnor U17227 (N_17227,N_14502,N_11712);
or U17228 (N_17228,N_14690,N_12728);
or U17229 (N_17229,N_14830,N_12843);
xor U17230 (N_17230,N_13392,N_14563);
nor U17231 (N_17231,N_12484,N_10298);
or U17232 (N_17232,N_14767,N_10906);
xnor U17233 (N_17233,N_14874,N_13127);
or U17234 (N_17234,N_12342,N_10705);
or U17235 (N_17235,N_12757,N_12340);
nand U17236 (N_17236,N_10200,N_13824);
xnor U17237 (N_17237,N_13039,N_13991);
nor U17238 (N_17238,N_12783,N_14974);
or U17239 (N_17239,N_14953,N_12884);
and U17240 (N_17240,N_14606,N_13441);
nor U17241 (N_17241,N_11605,N_11829);
nand U17242 (N_17242,N_11424,N_10586);
and U17243 (N_17243,N_11280,N_11711);
xnor U17244 (N_17244,N_10026,N_14972);
nand U17245 (N_17245,N_13059,N_12615);
or U17246 (N_17246,N_10423,N_11187);
or U17247 (N_17247,N_13821,N_10991);
nand U17248 (N_17248,N_14834,N_10141);
and U17249 (N_17249,N_10188,N_12531);
nand U17250 (N_17250,N_13379,N_11321);
xnor U17251 (N_17251,N_12148,N_13918);
or U17252 (N_17252,N_13682,N_11229);
and U17253 (N_17253,N_12439,N_14155);
nand U17254 (N_17254,N_14858,N_11382);
xor U17255 (N_17255,N_12767,N_11029);
nand U17256 (N_17256,N_14125,N_10276);
and U17257 (N_17257,N_12807,N_13638);
nand U17258 (N_17258,N_13889,N_10163);
xor U17259 (N_17259,N_10321,N_14553);
or U17260 (N_17260,N_14412,N_13259);
nand U17261 (N_17261,N_10243,N_11895);
nand U17262 (N_17262,N_10909,N_10594);
nor U17263 (N_17263,N_11675,N_13326);
nor U17264 (N_17264,N_12283,N_14283);
and U17265 (N_17265,N_12085,N_10061);
and U17266 (N_17266,N_10222,N_12211);
nor U17267 (N_17267,N_12770,N_11891);
or U17268 (N_17268,N_10692,N_14348);
or U17269 (N_17269,N_11336,N_12354);
and U17270 (N_17270,N_10404,N_10437);
and U17271 (N_17271,N_10722,N_10483);
nor U17272 (N_17272,N_12341,N_13274);
or U17273 (N_17273,N_10603,N_11637);
xnor U17274 (N_17274,N_13289,N_13668);
nor U17275 (N_17275,N_11262,N_13930);
nor U17276 (N_17276,N_10006,N_10441);
nor U17277 (N_17277,N_12528,N_14806);
xor U17278 (N_17278,N_13428,N_14351);
and U17279 (N_17279,N_14163,N_13019);
xnor U17280 (N_17280,N_12759,N_11355);
or U17281 (N_17281,N_10417,N_12320);
xnor U17282 (N_17282,N_10835,N_11435);
nor U17283 (N_17283,N_13253,N_14068);
and U17284 (N_17284,N_11025,N_12701);
nand U17285 (N_17285,N_13380,N_14639);
and U17286 (N_17286,N_12332,N_11555);
xor U17287 (N_17287,N_11421,N_12915);
xnor U17288 (N_17288,N_11086,N_12174);
xnor U17289 (N_17289,N_13878,N_14725);
nand U17290 (N_17290,N_11261,N_14587);
nand U17291 (N_17291,N_10315,N_12503);
xnor U17292 (N_17292,N_14993,N_14671);
xnor U17293 (N_17293,N_10996,N_11890);
xnor U17294 (N_17294,N_10035,N_14645);
nand U17295 (N_17295,N_14705,N_11070);
or U17296 (N_17296,N_10053,N_10625);
and U17297 (N_17297,N_13082,N_14281);
and U17298 (N_17298,N_12877,N_10511);
nand U17299 (N_17299,N_13100,N_13150);
nand U17300 (N_17300,N_11103,N_11290);
and U17301 (N_17301,N_10940,N_10916);
nor U17302 (N_17302,N_11214,N_12604);
and U17303 (N_17303,N_12216,N_10295);
nor U17304 (N_17304,N_13105,N_14417);
xnor U17305 (N_17305,N_14910,N_13055);
nor U17306 (N_17306,N_10084,N_13052);
xnor U17307 (N_17307,N_12763,N_13258);
and U17308 (N_17308,N_14067,N_14347);
or U17309 (N_17309,N_13737,N_14924);
xnor U17310 (N_17310,N_13588,N_10735);
and U17311 (N_17311,N_14228,N_14850);
xnor U17312 (N_17312,N_12102,N_10802);
nor U17313 (N_17313,N_14586,N_13178);
nor U17314 (N_17314,N_10602,N_12344);
and U17315 (N_17315,N_11462,N_11801);
or U17316 (N_17316,N_13429,N_14196);
nand U17317 (N_17317,N_13950,N_11292);
or U17318 (N_17318,N_12793,N_13385);
nand U17319 (N_17319,N_13768,N_14061);
xor U17320 (N_17320,N_12889,N_11379);
and U17321 (N_17321,N_14904,N_13029);
xor U17322 (N_17322,N_14719,N_10816);
or U17323 (N_17323,N_12632,N_10320);
or U17324 (N_17324,N_11507,N_14422);
and U17325 (N_17325,N_10770,N_14590);
xnor U17326 (N_17326,N_13621,N_10529);
or U17327 (N_17327,N_13313,N_11535);
nor U17328 (N_17328,N_10019,N_12084);
nand U17329 (N_17329,N_10402,N_10398);
and U17330 (N_17330,N_11771,N_11142);
nand U17331 (N_17331,N_12037,N_11976);
and U17332 (N_17332,N_11458,N_13498);
or U17333 (N_17333,N_14864,N_13393);
or U17334 (N_17334,N_10063,N_12787);
nor U17335 (N_17335,N_14946,N_12206);
nor U17336 (N_17336,N_11093,N_10546);
xnor U17337 (N_17337,N_12556,N_13740);
nor U17338 (N_17338,N_10847,N_11975);
nand U17339 (N_17339,N_14790,N_13572);
and U17340 (N_17340,N_12853,N_13890);
or U17341 (N_17341,N_10706,N_11696);
or U17342 (N_17342,N_13487,N_10762);
xnor U17343 (N_17343,N_12507,N_12327);
nor U17344 (N_17344,N_11762,N_13959);
nor U17345 (N_17345,N_11641,N_11346);
xor U17346 (N_17346,N_12231,N_14731);
or U17347 (N_17347,N_10928,N_11820);
xor U17348 (N_17348,N_11173,N_10375);
or U17349 (N_17349,N_12671,N_11136);
and U17350 (N_17350,N_12532,N_12714);
nand U17351 (N_17351,N_10240,N_13966);
xor U17352 (N_17352,N_11213,N_11337);
or U17353 (N_17353,N_10381,N_11568);
and U17354 (N_17354,N_14788,N_10174);
and U17355 (N_17355,N_12987,N_10156);
or U17356 (N_17356,N_11715,N_12780);
or U17357 (N_17357,N_12135,N_13206);
and U17358 (N_17358,N_14172,N_14710);
nand U17359 (N_17359,N_11920,N_13197);
nand U17360 (N_17360,N_13095,N_12900);
nor U17361 (N_17361,N_11085,N_12419);
and U17362 (N_17362,N_14800,N_12664);
or U17363 (N_17363,N_14158,N_10664);
nor U17364 (N_17364,N_14517,N_14841);
or U17365 (N_17365,N_13483,N_12146);
nand U17366 (N_17366,N_12593,N_12628);
nor U17367 (N_17367,N_11740,N_10798);
or U17368 (N_17368,N_10183,N_13497);
and U17369 (N_17369,N_10060,N_10774);
nor U17370 (N_17370,N_13748,N_12796);
xor U17371 (N_17371,N_10830,N_13330);
and U17372 (N_17372,N_10466,N_10597);
or U17373 (N_17373,N_12588,N_14711);
nor U17374 (N_17374,N_14353,N_14739);
nor U17375 (N_17375,N_14708,N_14603);
xnor U17376 (N_17376,N_13336,N_10710);
xor U17377 (N_17377,N_12012,N_11560);
nand U17378 (N_17378,N_12401,N_13898);
nor U17379 (N_17379,N_14284,N_14787);
and U17380 (N_17380,N_13176,N_12144);
nor U17381 (N_17381,N_14361,N_10449);
and U17382 (N_17382,N_13533,N_10281);
nor U17383 (N_17383,N_13125,N_10897);
or U17384 (N_17384,N_14524,N_14179);
or U17385 (N_17385,N_11948,N_11779);
nand U17386 (N_17386,N_10085,N_12926);
nor U17387 (N_17387,N_10202,N_14408);
xnor U17388 (N_17388,N_14766,N_11436);
xnor U17389 (N_17389,N_10604,N_12205);
or U17390 (N_17390,N_12249,N_14855);
and U17391 (N_17391,N_10244,N_11411);
xor U17392 (N_17392,N_13765,N_14043);
or U17393 (N_17393,N_10203,N_14595);
nor U17394 (N_17394,N_13000,N_14648);
and U17395 (N_17395,N_12049,N_10151);
and U17396 (N_17396,N_10709,N_13978);
nand U17397 (N_17397,N_10033,N_10667);
and U17398 (N_17398,N_12044,N_10111);
xor U17399 (N_17399,N_14254,N_11447);
nor U17400 (N_17400,N_10963,N_12237);
nor U17401 (N_17401,N_11523,N_11087);
nand U17402 (N_17402,N_12842,N_10032);
xor U17403 (N_17403,N_11293,N_13414);
nor U17404 (N_17404,N_14105,N_14726);
or U17405 (N_17405,N_10767,N_14688);
or U17406 (N_17406,N_10813,N_14393);
nor U17407 (N_17407,N_10448,N_13614);
nor U17408 (N_17408,N_10076,N_12570);
xnor U17409 (N_17409,N_14010,N_10656);
nand U17410 (N_17410,N_10645,N_14186);
nor U17411 (N_17411,N_14405,N_11759);
nor U17412 (N_17412,N_11731,N_13495);
or U17413 (N_17413,N_14110,N_14981);
and U17414 (N_17414,N_10463,N_13678);
and U17415 (N_17415,N_12271,N_11651);
nand U17416 (N_17416,N_12295,N_13788);
or U17417 (N_17417,N_12318,N_11849);
nor U17418 (N_17418,N_11713,N_14965);
and U17419 (N_17419,N_14385,N_14992);
and U17420 (N_17420,N_10193,N_11938);
and U17421 (N_17421,N_11177,N_14980);
nor U17422 (N_17422,N_12539,N_12323);
nand U17423 (N_17423,N_11392,N_14917);
and U17424 (N_17424,N_12345,N_14187);
xor U17425 (N_17425,N_12316,N_14979);
nand U17426 (N_17426,N_13310,N_12772);
xor U17427 (N_17427,N_14114,N_11318);
nor U17428 (N_17428,N_13884,N_13395);
nor U17429 (N_17429,N_14737,N_12321);
nand U17430 (N_17430,N_11902,N_11368);
nand U17431 (N_17431,N_12483,N_11924);
xor U17432 (N_17432,N_12659,N_11171);
nor U17433 (N_17433,N_11856,N_10818);
nand U17434 (N_17434,N_13356,N_12592);
or U17435 (N_17435,N_10287,N_11661);
or U17436 (N_17436,N_11282,N_13364);
xor U17437 (N_17437,N_11825,N_14576);
or U17438 (N_17438,N_11043,N_11076);
and U17439 (N_17439,N_10680,N_10685);
xor U17440 (N_17440,N_12648,N_10177);
nand U17441 (N_17441,N_11281,N_10401);
nand U17442 (N_17442,N_10621,N_13637);
or U17443 (N_17443,N_10775,N_11082);
nor U17444 (N_17444,N_10915,N_13877);
or U17445 (N_17445,N_14518,N_11331);
or U17446 (N_17446,N_11456,N_12371);
nor U17447 (N_17447,N_12501,N_13761);
nor U17448 (N_17448,N_10077,N_13484);
nand U17449 (N_17449,N_12992,N_10548);
nand U17450 (N_17450,N_11977,N_12096);
xor U17451 (N_17451,N_10640,N_13652);
xor U17452 (N_17452,N_12735,N_10306);
xor U17453 (N_17453,N_13239,N_11044);
xor U17454 (N_17454,N_10707,N_11882);
and U17455 (N_17455,N_13287,N_10132);
and U17456 (N_17456,N_13920,N_12280);
nor U17457 (N_17457,N_10776,N_13390);
nand U17458 (N_17458,N_13341,N_13147);
xor U17459 (N_17459,N_10197,N_10923);
nor U17460 (N_17460,N_13113,N_14275);
nor U17461 (N_17461,N_12382,N_11481);
nand U17462 (N_17462,N_12773,N_13711);
and U17463 (N_17463,N_14024,N_13462);
nor U17464 (N_17464,N_11760,N_13620);
or U17465 (N_17465,N_12449,N_11169);
or U17466 (N_17466,N_12675,N_13236);
nor U17467 (N_17467,N_10790,N_14617);
or U17468 (N_17468,N_11241,N_12052);
or U17469 (N_17469,N_10481,N_14480);
or U17470 (N_17470,N_13496,N_14722);
nand U17471 (N_17471,N_13421,N_10074);
xnor U17472 (N_17472,N_14709,N_11930);
or U17473 (N_17473,N_12552,N_10067);
and U17474 (N_17474,N_13683,N_14956);
nor U17475 (N_17475,N_10559,N_13545);
nand U17476 (N_17476,N_11918,N_12067);
and U17477 (N_17477,N_12533,N_14312);
or U17478 (N_17478,N_10263,N_10677);
nand U17479 (N_17479,N_14047,N_10949);
xnor U17480 (N_17480,N_10876,N_14798);
xnor U17481 (N_17481,N_10152,N_13345);
or U17482 (N_17482,N_12181,N_12741);
nor U17483 (N_17483,N_13980,N_11039);
xnor U17484 (N_17484,N_14195,N_10308);
xnor U17485 (N_17485,N_13860,N_11061);
and U17486 (N_17486,N_14252,N_11263);
or U17487 (N_17487,N_14407,N_11547);
and U17488 (N_17488,N_11559,N_14018);
xnor U17489 (N_17489,N_10241,N_10944);
nor U17490 (N_17490,N_13048,N_14011);
xor U17491 (N_17491,N_12765,N_12423);
or U17492 (N_17492,N_12799,N_13826);
or U17493 (N_17493,N_14029,N_13590);
xor U17494 (N_17494,N_14837,N_13899);
nor U17495 (N_17495,N_13780,N_13911);
xor U17496 (N_17496,N_12298,N_11634);
nor U17497 (N_17497,N_14269,N_11913);
or U17498 (N_17498,N_13615,N_10290);
or U17499 (N_17499,N_13104,N_13145);
nand U17500 (N_17500,N_12500,N_14596);
nor U17501 (N_17501,N_11932,N_14532);
nor U17502 (N_17502,N_12409,N_12702);
nand U17503 (N_17503,N_12428,N_13129);
xnor U17504 (N_17504,N_10694,N_12784);
nor U17505 (N_17505,N_13477,N_14821);
xor U17506 (N_17506,N_12262,N_13899);
and U17507 (N_17507,N_12606,N_11682);
or U17508 (N_17508,N_12771,N_11910);
nand U17509 (N_17509,N_11444,N_14431);
xnor U17510 (N_17510,N_14765,N_13020);
and U17511 (N_17511,N_14635,N_13085);
and U17512 (N_17512,N_13253,N_12490);
and U17513 (N_17513,N_11166,N_14240);
or U17514 (N_17514,N_12471,N_14572);
nand U17515 (N_17515,N_12401,N_11902);
and U17516 (N_17516,N_10008,N_11743);
xnor U17517 (N_17517,N_11282,N_10867);
nand U17518 (N_17518,N_13138,N_10776);
or U17519 (N_17519,N_12128,N_13629);
xor U17520 (N_17520,N_14779,N_12219);
nor U17521 (N_17521,N_13155,N_13361);
xnor U17522 (N_17522,N_12152,N_14389);
xor U17523 (N_17523,N_11620,N_11094);
or U17524 (N_17524,N_11109,N_14722);
xnor U17525 (N_17525,N_11207,N_10406);
or U17526 (N_17526,N_14659,N_10942);
nor U17527 (N_17527,N_12393,N_10341);
and U17528 (N_17528,N_12909,N_12950);
or U17529 (N_17529,N_11248,N_10037);
and U17530 (N_17530,N_12417,N_12480);
nand U17531 (N_17531,N_11190,N_10534);
xor U17532 (N_17532,N_12017,N_11283);
nor U17533 (N_17533,N_10466,N_10512);
xor U17534 (N_17534,N_14551,N_13231);
nand U17535 (N_17535,N_14737,N_13229);
nand U17536 (N_17536,N_14697,N_10378);
or U17537 (N_17537,N_14719,N_12161);
xnor U17538 (N_17538,N_14762,N_12146);
and U17539 (N_17539,N_13841,N_14275);
xnor U17540 (N_17540,N_14533,N_14417);
nand U17541 (N_17541,N_13861,N_10293);
nor U17542 (N_17542,N_14672,N_13119);
and U17543 (N_17543,N_14762,N_14704);
xnor U17544 (N_17544,N_11850,N_14907);
nand U17545 (N_17545,N_12606,N_11573);
and U17546 (N_17546,N_13757,N_13242);
xor U17547 (N_17547,N_13540,N_12942);
nand U17548 (N_17548,N_12630,N_13880);
nand U17549 (N_17549,N_10472,N_12331);
nand U17550 (N_17550,N_12977,N_12616);
and U17551 (N_17551,N_11166,N_10466);
nand U17552 (N_17552,N_14529,N_11469);
nor U17553 (N_17553,N_10108,N_14327);
nor U17554 (N_17554,N_13799,N_11265);
xor U17555 (N_17555,N_11460,N_11253);
and U17556 (N_17556,N_13658,N_11683);
nand U17557 (N_17557,N_11759,N_14167);
xor U17558 (N_17558,N_13762,N_11340);
and U17559 (N_17559,N_11164,N_14607);
nor U17560 (N_17560,N_10619,N_13494);
and U17561 (N_17561,N_10352,N_14917);
nand U17562 (N_17562,N_10345,N_10997);
and U17563 (N_17563,N_12645,N_13276);
and U17564 (N_17564,N_11957,N_13979);
nand U17565 (N_17565,N_11388,N_14930);
or U17566 (N_17566,N_13102,N_12459);
or U17567 (N_17567,N_10460,N_12894);
xnor U17568 (N_17568,N_11325,N_14440);
and U17569 (N_17569,N_10768,N_13096);
nor U17570 (N_17570,N_14263,N_13652);
nor U17571 (N_17571,N_14147,N_13672);
and U17572 (N_17572,N_10468,N_13589);
xnor U17573 (N_17573,N_12263,N_14820);
and U17574 (N_17574,N_10240,N_10166);
and U17575 (N_17575,N_13375,N_12372);
nand U17576 (N_17576,N_10623,N_14187);
nand U17577 (N_17577,N_11056,N_12392);
and U17578 (N_17578,N_11258,N_10374);
nor U17579 (N_17579,N_10082,N_14428);
or U17580 (N_17580,N_10655,N_11175);
nor U17581 (N_17581,N_12686,N_12803);
and U17582 (N_17582,N_10310,N_10512);
xnor U17583 (N_17583,N_11334,N_10583);
and U17584 (N_17584,N_10581,N_13440);
and U17585 (N_17585,N_13286,N_10100);
or U17586 (N_17586,N_13148,N_11316);
nor U17587 (N_17587,N_13405,N_13690);
and U17588 (N_17588,N_12826,N_13917);
xor U17589 (N_17589,N_12543,N_13011);
or U17590 (N_17590,N_11758,N_11008);
and U17591 (N_17591,N_11982,N_10587);
and U17592 (N_17592,N_10350,N_11953);
or U17593 (N_17593,N_13714,N_10249);
nand U17594 (N_17594,N_12138,N_13804);
nand U17595 (N_17595,N_10623,N_11464);
xor U17596 (N_17596,N_12363,N_14466);
or U17597 (N_17597,N_11781,N_11179);
or U17598 (N_17598,N_13329,N_10229);
and U17599 (N_17599,N_13714,N_12096);
nand U17600 (N_17600,N_11422,N_10376);
nor U17601 (N_17601,N_14846,N_11406);
xnor U17602 (N_17602,N_13532,N_11769);
or U17603 (N_17603,N_11817,N_10670);
and U17604 (N_17604,N_13940,N_10819);
or U17605 (N_17605,N_14802,N_12489);
or U17606 (N_17606,N_13942,N_10417);
nand U17607 (N_17607,N_10982,N_11554);
xor U17608 (N_17608,N_12694,N_12871);
and U17609 (N_17609,N_12699,N_10654);
xnor U17610 (N_17610,N_12539,N_12406);
nand U17611 (N_17611,N_13273,N_14957);
nand U17612 (N_17612,N_11088,N_12919);
and U17613 (N_17613,N_12967,N_11678);
or U17614 (N_17614,N_13416,N_10671);
nor U17615 (N_17615,N_13447,N_11899);
or U17616 (N_17616,N_10538,N_12768);
xnor U17617 (N_17617,N_12243,N_14132);
nand U17618 (N_17618,N_12743,N_11633);
and U17619 (N_17619,N_14093,N_10342);
or U17620 (N_17620,N_13909,N_13916);
nor U17621 (N_17621,N_14918,N_10433);
nor U17622 (N_17622,N_11663,N_13832);
or U17623 (N_17623,N_10678,N_10953);
or U17624 (N_17624,N_13511,N_11342);
or U17625 (N_17625,N_11972,N_10438);
xnor U17626 (N_17626,N_12614,N_10428);
nor U17627 (N_17627,N_12766,N_10952);
nand U17628 (N_17628,N_12731,N_10823);
or U17629 (N_17629,N_10893,N_13946);
nor U17630 (N_17630,N_13254,N_14272);
and U17631 (N_17631,N_13750,N_14951);
or U17632 (N_17632,N_10980,N_10397);
xor U17633 (N_17633,N_14649,N_13622);
nor U17634 (N_17634,N_13983,N_10778);
xor U17635 (N_17635,N_14871,N_10828);
and U17636 (N_17636,N_10249,N_11650);
xor U17637 (N_17637,N_10929,N_13743);
or U17638 (N_17638,N_13896,N_14191);
nor U17639 (N_17639,N_12672,N_10952);
and U17640 (N_17640,N_11737,N_13197);
nand U17641 (N_17641,N_10603,N_10279);
or U17642 (N_17642,N_10737,N_13292);
nand U17643 (N_17643,N_10261,N_10022);
nor U17644 (N_17644,N_10894,N_14393);
xor U17645 (N_17645,N_14467,N_14607);
and U17646 (N_17646,N_14703,N_10876);
nor U17647 (N_17647,N_13471,N_14372);
xnor U17648 (N_17648,N_12612,N_12253);
nor U17649 (N_17649,N_11567,N_10307);
nand U17650 (N_17650,N_14092,N_13781);
nand U17651 (N_17651,N_14676,N_11999);
and U17652 (N_17652,N_12959,N_10079);
or U17653 (N_17653,N_14260,N_12137);
nor U17654 (N_17654,N_14020,N_12287);
and U17655 (N_17655,N_10261,N_14400);
nand U17656 (N_17656,N_10581,N_14789);
and U17657 (N_17657,N_10282,N_12514);
and U17658 (N_17658,N_11133,N_10245);
and U17659 (N_17659,N_14890,N_13484);
nor U17660 (N_17660,N_13973,N_11450);
or U17661 (N_17661,N_11448,N_14880);
or U17662 (N_17662,N_13372,N_14451);
xor U17663 (N_17663,N_11370,N_12243);
nand U17664 (N_17664,N_13294,N_10140);
and U17665 (N_17665,N_12370,N_13000);
nand U17666 (N_17666,N_11628,N_11151);
and U17667 (N_17667,N_12410,N_11228);
xnor U17668 (N_17668,N_10692,N_10125);
xnor U17669 (N_17669,N_13203,N_12759);
nor U17670 (N_17670,N_10387,N_13529);
and U17671 (N_17671,N_14044,N_10243);
or U17672 (N_17672,N_11097,N_14836);
or U17673 (N_17673,N_11168,N_13410);
or U17674 (N_17674,N_13593,N_14414);
or U17675 (N_17675,N_12028,N_14791);
and U17676 (N_17676,N_13902,N_14910);
and U17677 (N_17677,N_13672,N_13224);
nor U17678 (N_17678,N_12025,N_12962);
or U17679 (N_17679,N_14116,N_10272);
nand U17680 (N_17680,N_13875,N_11994);
nor U17681 (N_17681,N_14876,N_13584);
and U17682 (N_17682,N_11926,N_12669);
nor U17683 (N_17683,N_12687,N_11785);
xor U17684 (N_17684,N_12733,N_13238);
and U17685 (N_17685,N_10388,N_10514);
and U17686 (N_17686,N_13006,N_12648);
nor U17687 (N_17687,N_12095,N_12382);
and U17688 (N_17688,N_10558,N_10567);
nor U17689 (N_17689,N_13490,N_10304);
nand U17690 (N_17690,N_10788,N_10006);
nand U17691 (N_17691,N_12386,N_14103);
or U17692 (N_17692,N_11984,N_12110);
xnor U17693 (N_17693,N_11137,N_14837);
nand U17694 (N_17694,N_10823,N_10778);
nand U17695 (N_17695,N_14526,N_14570);
nor U17696 (N_17696,N_12332,N_11881);
xor U17697 (N_17697,N_12744,N_13392);
nand U17698 (N_17698,N_12699,N_12806);
or U17699 (N_17699,N_10570,N_14787);
and U17700 (N_17700,N_10509,N_10515);
nor U17701 (N_17701,N_12700,N_12285);
nor U17702 (N_17702,N_12427,N_11740);
nor U17703 (N_17703,N_14366,N_12888);
nand U17704 (N_17704,N_14168,N_14057);
and U17705 (N_17705,N_10822,N_12607);
or U17706 (N_17706,N_14786,N_10291);
xnor U17707 (N_17707,N_12727,N_13107);
and U17708 (N_17708,N_14190,N_14563);
or U17709 (N_17709,N_11363,N_10152);
or U17710 (N_17710,N_13653,N_10804);
xnor U17711 (N_17711,N_10776,N_10401);
or U17712 (N_17712,N_14015,N_10097);
nor U17713 (N_17713,N_10557,N_13563);
and U17714 (N_17714,N_11159,N_14483);
nor U17715 (N_17715,N_11220,N_10313);
nand U17716 (N_17716,N_11811,N_14894);
xor U17717 (N_17717,N_11143,N_13360);
and U17718 (N_17718,N_11933,N_13597);
nor U17719 (N_17719,N_10775,N_10967);
or U17720 (N_17720,N_12430,N_10582);
nor U17721 (N_17721,N_13470,N_13581);
nor U17722 (N_17722,N_11787,N_12567);
or U17723 (N_17723,N_11973,N_12524);
nor U17724 (N_17724,N_11062,N_12534);
xnor U17725 (N_17725,N_13119,N_10619);
nor U17726 (N_17726,N_12134,N_13944);
or U17727 (N_17727,N_10749,N_14121);
nand U17728 (N_17728,N_13381,N_13512);
xnor U17729 (N_17729,N_13811,N_14251);
nand U17730 (N_17730,N_10736,N_13137);
nor U17731 (N_17731,N_11210,N_12191);
nor U17732 (N_17732,N_11279,N_14615);
and U17733 (N_17733,N_10114,N_11199);
and U17734 (N_17734,N_11385,N_12990);
nand U17735 (N_17735,N_12069,N_13508);
or U17736 (N_17736,N_10542,N_14462);
xnor U17737 (N_17737,N_14012,N_10382);
nand U17738 (N_17738,N_13152,N_10624);
xor U17739 (N_17739,N_10565,N_10163);
xor U17740 (N_17740,N_12153,N_14918);
nand U17741 (N_17741,N_11247,N_12967);
xor U17742 (N_17742,N_11094,N_13527);
and U17743 (N_17743,N_11954,N_11115);
or U17744 (N_17744,N_13737,N_14179);
and U17745 (N_17745,N_11922,N_13729);
or U17746 (N_17746,N_14753,N_11334);
xnor U17747 (N_17747,N_13854,N_14050);
nor U17748 (N_17748,N_12869,N_11532);
nor U17749 (N_17749,N_14776,N_13478);
nor U17750 (N_17750,N_14832,N_14864);
xor U17751 (N_17751,N_13793,N_14887);
or U17752 (N_17752,N_11535,N_11341);
nor U17753 (N_17753,N_12820,N_10731);
xnor U17754 (N_17754,N_13858,N_10325);
or U17755 (N_17755,N_11529,N_13631);
or U17756 (N_17756,N_13581,N_11265);
xnor U17757 (N_17757,N_14576,N_12269);
xor U17758 (N_17758,N_11911,N_13151);
xor U17759 (N_17759,N_12807,N_12052);
nor U17760 (N_17760,N_14405,N_13909);
xor U17761 (N_17761,N_10954,N_12683);
nor U17762 (N_17762,N_13855,N_12394);
nor U17763 (N_17763,N_10236,N_11825);
and U17764 (N_17764,N_13096,N_14225);
nand U17765 (N_17765,N_10101,N_14885);
nand U17766 (N_17766,N_11926,N_14980);
nand U17767 (N_17767,N_13485,N_11131);
and U17768 (N_17768,N_14773,N_14879);
xor U17769 (N_17769,N_10413,N_14639);
or U17770 (N_17770,N_14688,N_10117);
nand U17771 (N_17771,N_11282,N_10853);
nand U17772 (N_17772,N_10662,N_12625);
or U17773 (N_17773,N_14405,N_11649);
nor U17774 (N_17774,N_12367,N_12389);
nand U17775 (N_17775,N_13111,N_13725);
nor U17776 (N_17776,N_12152,N_12581);
or U17777 (N_17777,N_11455,N_11944);
nand U17778 (N_17778,N_11113,N_14747);
xor U17779 (N_17779,N_12588,N_14476);
or U17780 (N_17780,N_10123,N_11494);
nand U17781 (N_17781,N_13130,N_14188);
xor U17782 (N_17782,N_12508,N_14555);
and U17783 (N_17783,N_12417,N_11633);
xor U17784 (N_17784,N_12899,N_11569);
nor U17785 (N_17785,N_14864,N_13267);
and U17786 (N_17786,N_11523,N_14124);
xor U17787 (N_17787,N_10512,N_13742);
or U17788 (N_17788,N_12200,N_10032);
nor U17789 (N_17789,N_13318,N_11062);
nand U17790 (N_17790,N_10401,N_13877);
nor U17791 (N_17791,N_10334,N_12845);
nand U17792 (N_17792,N_12369,N_14551);
nand U17793 (N_17793,N_13561,N_11595);
nor U17794 (N_17794,N_14719,N_12299);
nor U17795 (N_17795,N_12500,N_12300);
and U17796 (N_17796,N_14089,N_11779);
and U17797 (N_17797,N_10430,N_10744);
or U17798 (N_17798,N_12569,N_14105);
nor U17799 (N_17799,N_13453,N_13345);
nand U17800 (N_17800,N_13709,N_10551);
or U17801 (N_17801,N_10517,N_10295);
xnor U17802 (N_17802,N_13740,N_14423);
or U17803 (N_17803,N_13813,N_13283);
xnor U17804 (N_17804,N_13796,N_10797);
or U17805 (N_17805,N_11332,N_11393);
nand U17806 (N_17806,N_12804,N_10544);
and U17807 (N_17807,N_11927,N_12817);
xor U17808 (N_17808,N_13844,N_10527);
and U17809 (N_17809,N_14529,N_14553);
xnor U17810 (N_17810,N_12483,N_14176);
or U17811 (N_17811,N_13732,N_11611);
or U17812 (N_17812,N_14503,N_13275);
nand U17813 (N_17813,N_12742,N_11369);
and U17814 (N_17814,N_10400,N_11816);
or U17815 (N_17815,N_13181,N_11832);
xnor U17816 (N_17816,N_10340,N_13632);
nand U17817 (N_17817,N_11997,N_12104);
nor U17818 (N_17818,N_13737,N_12175);
nor U17819 (N_17819,N_12514,N_11519);
or U17820 (N_17820,N_13882,N_13221);
nor U17821 (N_17821,N_10037,N_12174);
and U17822 (N_17822,N_11406,N_14984);
and U17823 (N_17823,N_13675,N_13364);
nor U17824 (N_17824,N_14528,N_13571);
and U17825 (N_17825,N_10563,N_13515);
and U17826 (N_17826,N_14758,N_11221);
nor U17827 (N_17827,N_11172,N_13225);
nor U17828 (N_17828,N_12221,N_13545);
and U17829 (N_17829,N_13994,N_13333);
nor U17830 (N_17830,N_12669,N_13225);
nand U17831 (N_17831,N_14960,N_11144);
and U17832 (N_17832,N_14707,N_12771);
xnor U17833 (N_17833,N_11495,N_12346);
nand U17834 (N_17834,N_10583,N_14612);
and U17835 (N_17835,N_12336,N_12265);
nor U17836 (N_17836,N_11218,N_13640);
nand U17837 (N_17837,N_14904,N_13492);
and U17838 (N_17838,N_13221,N_14554);
and U17839 (N_17839,N_11500,N_11464);
nor U17840 (N_17840,N_10106,N_10385);
nor U17841 (N_17841,N_12905,N_13926);
or U17842 (N_17842,N_14294,N_11560);
and U17843 (N_17843,N_12979,N_14472);
nor U17844 (N_17844,N_11675,N_11780);
or U17845 (N_17845,N_14591,N_10998);
nand U17846 (N_17846,N_12997,N_11566);
and U17847 (N_17847,N_13251,N_13409);
xor U17848 (N_17848,N_12070,N_12870);
or U17849 (N_17849,N_10578,N_11034);
nand U17850 (N_17850,N_14272,N_12944);
or U17851 (N_17851,N_10986,N_11815);
nand U17852 (N_17852,N_12266,N_11324);
xnor U17853 (N_17853,N_14836,N_12325);
nand U17854 (N_17854,N_14243,N_14819);
nor U17855 (N_17855,N_10251,N_12614);
nand U17856 (N_17856,N_11593,N_10043);
xnor U17857 (N_17857,N_11018,N_14184);
and U17858 (N_17858,N_13046,N_12897);
or U17859 (N_17859,N_13597,N_13172);
nor U17860 (N_17860,N_10416,N_13138);
or U17861 (N_17861,N_13407,N_12088);
and U17862 (N_17862,N_14832,N_12061);
nor U17863 (N_17863,N_10616,N_12208);
nand U17864 (N_17864,N_14256,N_10218);
xnor U17865 (N_17865,N_14233,N_14987);
nor U17866 (N_17866,N_12405,N_12823);
xor U17867 (N_17867,N_14861,N_14056);
xnor U17868 (N_17868,N_10149,N_11884);
and U17869 (N_17869,N_14773,N_10517);
xnor U17870 (N_17870,N_14908,N_14350);
or U17871 (N_17871,N_12173,N_11039);
nand U17872 (N_17872,N_11382,N_12433);
or U17873 (N_17873,N_13630,N_10303);
xor U17874 (N_17874,N_13674,N_12181);
nor U17875 (N_17875,N_12858,N_14776);
and U17876 (N_17876,N_10082,N_12919);
or U17877 (N_17877,N_14348,N_13143);
nand U17878 (N_17878,N_12777,N_14091);
or U17879 (N_17879,N_14704,N_14485);
nand U17880 (N_17880,N_13655,N_12589);
nand U17881 (N_17881,N_10984,N_12997);
nand U17882 (N_17882,N_14665,N_11452);
or U17883 (N_17883,N_10952,N_13241);
xnor U17884 (N_17884,N_10665,N_11176);
nand U17885 (N_17885,N_13147,N_11092);
xor U17886 (N_17886,N_10233,N_13112);
nor U17887 (N_17887,N_10579,N_10618);
or U17888 (N_17888,N_12712,N_13152);
or U17889 (N_17889,N_10783,N_10507);
nand U17890 (N_17890,N_12741,N_10626);
xor U17891 (N_17891,N_11266,N_10941);
and U17892 (N_17892,N_13891,N_14962);
or U17893 (N_17893,N_10676,N_13825);
nand U17894 (N_17894,N_11041,N_14699);
nor U17895 (N_17895,N_11260,N_13103);
xnor U17896 (N_17896,N_14716,N_13579);
and U17897 (N_17897,N_14057,N_14055);
and U17898 (N_17898,N_11032,N_13871);
xor U17899 (N_17899,N_13599,N_10471);
or U17900 (N_17900,N_12350,N_13110);
nor U17901 (N_17901,N_14218,N_11907);
and U17902 (N_17902,N_10605,N_14626);
nor U17903 (N_17903,N_10640,N_11552);
nor U17904 (N_17904,N_12800,N_10077);
and U17905 (N_17905,N_10640,N_10401);
or U17906 (N_17906,N_14066,N_10930);
nand U17907 (N_17907,N_11328,N_14318);
nor U17908 (N_17908,N_13326,N_11545);
nor U17909 (N_17909,N_11303,N_13149);
nand U17910 (N_17910,N_10208,N_10343);
xor U17911 (N_17911,N_11857,N_10169);
xnor U17912 (N_17912,N_10914,N_14490);
nand U17913 (N_17913,N_13977,N_11485);
and U17914 (N_17914,N_14291,N_12893);
nor U17915 (N_17915,N_14174,N_11138);
xor U17916 (N_17916,N_13287,N_14687);
and U17917 (N_17917,N_10109,N_14558);
nor U17918 (N_17918,N_13073,N_10691);
xor U17919 (N_17919,N_14600,N_10750);
nand U17920 (N_17920,N_10344,N_12525);
nor U17921 (N_17921,N_10609,N_10172);
nand U17922 (N_17922,N_13233,N_12327);
or U17923 (N_17923,N_10883,N_13179);
nor U17924 (N_17924,N_10586,N_13337);
nor U17925 (N_17925,N_11927,N_13513);
nand U17926 (N_17926,N_12222,N_14940);
xnor U17927 (N_17927,N_10953,N_11739);
nor U17928 (N_17928,N_12920,N_11421);
or U17929 (N_17929,N_10113,N_14622);
and U17930 (N_17930,N_10816,N_12118);
or U17931 (N_17931,N_11254,N_10167);
and U17932 (N_17932,N_14432,N_10480);
and U17933 (N_17933,N_14915,N_14431);
and U17934 (N_17934,N_12394,N_12943);
nand U17935 (N_17935,N_14418,N_12184);
nand U17936 (N_17936,N_10452,N_12219);
and U17937 (N_17937,N_11015,N_12585);
nor U17938 (N_17938,N_11298,N_12448);
nor U17939 (N_17939,N_14555,N_10420);
nand U17940 (N_17940,N_13405,N_10482);
nand U17941 (N_17941,N_14092,N_10480);
or U17942 (N_17942,N_12514,N_12730);
xor U17943 (N_17943,N_13724,N_14279);
and U17944 (N_17944,N_10459,N_11102);
nand U17945 (N_17945,N_14078,N_14063);
or U17946 (N_17946,N_14620,N_13840);
xnor U17947 (N_17947,N_10148,N_11763);
or U17948 (N_17948,N_11337,N_12313);
nand U17949 (N_17949,N_14633,N_11061);
nor U17950 (N_17950,N_12773,N_11180);
or U17951 (N_17951,N_14545,N_14693);
or U17952 (N_17952,N_13280,N_12261);
nor U17953 (N_17953,N_13469,N_10110);
and U17954 (N_17954,N_10625,N_11466);
nand U17955 (N_17955,N_13928,N_13693);
nand U17956 (N_17956,N_10706,N_13567);
nor U17957 (N_17957,N_12502,N_11710);
and U17958 (N_17958,N_14024,N_11263);
or U17959 (N_17959,N_11859,N_14054);
nor U17960 (N_17960,N_12637,N_14376);
xnor U17961 (N_17961,N_10556,N_10335);
nor U17962 (N_17962,N_13430,N_11653);
xnor U17963 (N_17963,N_11304,N_13086);
and U17964 (N_17964,N_11583,N_13262);
xor U17965 (N_17965,N_12617,N_11252);
nor U17966 (N_17966,N_10770,N_10994);
nor U17967 (N_17967,N_10644,N_10399);
or U17968 (N_17968,N_14397,N_11849);
nand U17969 (N_17969,N_12860,N_10863);
xor U17970 (N_17970,N_10038,N_11417);
nand U17971 (N_17971,N_11370,N_10936);
or U17972 (N_17972,N_13984,N_14480);
xnor U17973 (N_17973,N_12255,N_12003);
and U17974 (N_17974,N_13152,N_13565);
xor U17975 (N_17975,N_10383,N_11357);
and U17976 (N_17976,N_11642,N_11052);
xor U17977 (N_17977,N_10198,N_10493);
nor U17978 (N_17978,N_13152,N_11683);
xnor U17979 (N_17979,N_12994,N_13073);
or U17980 (N_17980,N_12268,N_14153);
and U17981 (N_17981,N_14061,N_14072);
nand U17982 (N_17982,N_10764,N_10502);
nand U17983 (N_17983,N_10658,N_14824);
or U17984 (N_17984,N_11381,N_14729);
and U17985 (N_17985,N_13932,N_10188);
or U17986 (N_17986,N_11396,N_11333);
and U17987 (N_17987,N_14667,N_10045);
nand U17988 (N_17988,N_12375,N_12437);
xor U17989 (N_17989,N_13006,N_12058);
or U17990 (N_17990,N_11423,N_14190);
nand U17991 (N_17991,N_11443,N_12561);
and U17992 (N_17992,N_10013,N_14949);
xor U17993 (N_17993,N_12454,N_14372);
and U17994 (N_17994,N_11564,N_12237);
xnor U17995 (N_17995,N_14442,N_12138);
or U17996 (N_17996,N_13467,N_12382);
and U17997 (N_17997,N_10906,N_13283);
nand U17998 (N_17998,N_13526,N_11815);
and U17999 (N_17999,N_12365,N_13426);
xnor U18000 (N_18000,N_11958,N_10861);
or U18001 (N_18001,N_12228,N_13297);
and U18002 (N_18002,N_13846,N_10402);
nand U18003 (N_18003,N_13570,N_12839);
xnor U18004 (N_18004,N_13132,N_13407);
and U18005 (N_18005,N_14033,N_14182);
and U18006 (N_18006,N_14477,N_13742);
nor U18007 (N_18007,N_10964,N_14417);
nor U18008 (N_18008,N_12797,N_13381);
nand U18009 (N_18009,N_13826,N_12934);
xor U18010 (N_18010,N_11507,N_11738);
nor U18011 (N_18011,N_11001,N_13086);
nor U18012 (N_18012,N_12285,N_11298);
xor U18013 (N_18013,N_14761,N_14018);
nor U18014 (N_18014,N_11957,N_11474);
nand U18015 (N_18015,N_12714,N_14172);
or U18016 (N_18016,N_11652,N_14004);
nor U18017 (N_18017,N_13828,N_10337);
and U18018 (N_18018,N_14523,N_13665);
and U18019 (N_18019,N_13207,N_13217);
and U18020 (N_18020,N_11270,N_14785);
nor U18021 (N_18021,N_12917,N_11904);
and U18022 (N_18022,N_11611,N_13545);
nor U18023 (N_18023,N_11038,N_11597);
or U18024 (N_18024,N_12432,N_11839);
nor U18025 (N_18025,N_14572,N_14798);
nand U18026 (N_18026,N_10445,N_11240);
nand U18027 (N_18027,N_13393,N_12899);
nor U18028 (N_18028,N_11312,N_13748);
nor U18029 (N_18029,N_12477,N_13251);
nor U18030 (N_18030,N_14418,N_10345);
nand U18031 (N_18031,N_13092,N_12872);
nand U18032 (N_18032,N_14165,N_13555);
nand U18033 (N_18033,N_11891,N_14559);
nand U18034 (N_18034,N_12608,N_11925);
nor U18035 (N_18035,N_12971,N_12281);
and U18036 (N_18036,N_11208,N_11270);
and U18037 (N_18037,N_11624,N_12411);
and U18038 (N_18038,N_10878,N_14143);
nor U18039 (N_18039,N_12755,N_12776);
nor U18040 (N_18040,N_10744,N_12181);
nand U18041 (N_18041,N_14862,N_10528);
xor U18042 (N_18042,N_11932,N_14696);
xor U18043 (N_18043,N_14694,N_13104);
and U18044 (N_18044,N_10493,N_14544);
xnor U18045 (N_18045,N_13035,N_14590);
nor U18046 (N_18046,N_11929,N_14051);
and U18047 (N_18047,N_10220,N_14443);
or U18048 (N_18048,N_14817,N_10173);
and U18049 (N_18049,N_12702,N_12795);
or U18050 (N_18050,N_11026,N_13529);
nand U18051 (N_18051,N_12519,N_10345);
or U18052 (N_18052,N_13082,N_13387);
or U18053 (N_18053,N_13974,N_12745);
xor U18054 (N_18054,N_10283,N_11511);
nor U18055 (N_18055,N_10881,N_13310);
nor U18056 (N_18056,N_13423,N_10264);
xor U18057 (N_18057,N_11133,N_10711);
nor U18058 (N_18058,N_11613,N_14868);
or U18059 (N_18059,N_13235,N_10334);
or U18060 (N_18060,N_10516,N_12444);
nand U18061 (N_18061,N_14497,N_13790);
or U18062 (N_18062,N_11997,N_10306);
nand U18063 (N_18063,N_13203,N_11528);
nand U18064 (N_18064,N_11614,N_13734);
nand U18065 (N_18065,N_13197,N_12926);
nand U18066 (N_18066,N_12190,N_13000);
or U18067 (N_18067,N_10363,N_14610);
nand U18068 (N_18068,N_14323,N_12872);
xnor U18069 (N_18069,N_14777,N_11438);
or U18070 (N_18070,N_14593,N_12687);
nor U18071 (N_18071,N_13154,N_12272);
and U18072 (N_18072,N_11487,N_12979);
nor U18073 (N_18073,N_14015,N_10417);
xnor U18074 (N_18074,N_13479,N_12631);
xor U18075 (N_18075,N_13303,N_13704);
nor U18076 (N_18076,N_10902,N_12355);
nand U18077 (N_18077,N_11053,N_13915);
xor U18078 (N_18078,N_14217,N_12246);
and U18079 (N_18079,N_10316,N_13468);
xor U18080 (N_18080,N_10840,N_14604);
xor U18081 (N_18081,N_10054,N_13893);
nor U18082 (N_18082,N_12777,N_11056);
xnor U18083 (N_18083,N_14275,N_12939);
xnor U18084 (N_18084,N_11105,N_14549);
xor U18085 (N_18085,N_13450,N_13722);
nor U18086 (N_18086,N_11302,N_11538);
nor U18087 (N_18087,N_14944,N_12063);
xor U18088 (N_18088,N_12044,N_13255);
nor U18089 (N_18089,N_11527,N_14990);
and U18090 (N_18090,N_14895,N_10178);
and U18091 (N_18091,N_11740,N_10258);
or U18092 (N_18092,N_11932,N_10508);
nor U18093 (N_18093,N_13400,N_12981);
nor U18094 (N_18094,N_10305,N_10636);
nor U18095 (N_18095,N_11100,N_14303);
nor U18096 (N_18096,N_11227,N_12233);
and U18097 (N_18097,N_12101,N_13765);
xor U18098 (N_18098,N_12637,N_13114);
or U18099 (N_18099,N_13782,N_12635);
and U18100 (N_18100,N_10371,N_12493);
nand U18101 (N_18101,N_12420,N_14299);
and U18102 (N_18102,N_13516,N_13015);
or U18103 (N_18103,N_12694,N_10270);
and U18104 (N_18104,N_12899,N_14476);
nor U18105 (N_18105,N_11580,N_14991);
nand U18106 (N_18106,N_13370,N_14929);
and U18107 (N_18107,N_11141,N_11307);
nand U18108 (N_18108,N_11084,N_14382);
nor U18109 (N_18109,N_12792,N_13863);
or U18110 (N_18110,N_12341,N_11010);
or U18111 (N_18111,N_10706,N_14556);
or U18112 (N_18112,N_14354,N_10392);
or U18113 (N_18113,N_13102,N_10749);
nor U18114 (N_18114,N_11536,N_11383);
xnor U18115 (N_18115,N_12170,N_13801);
nand U18116 (N_18116,N_10303,N_14690);
or U18117 (N_18117,N_11823,N_14662);
nand U18118 (N_18118,N_10771,N_10252);
xnor U18119 (N_18119,N_11673,N_13736);
nor U18120 (N_18120,N_11459,N_12134);
nand U18121 (N_18121,N_13446,N_13460);
or U18122 (N_18122,N_10679,N_12965);
xnor U18123 (N_18123,N_11273,N_13878);
nor U18124 (N_18124,N_12217,N_13797);
xnor U18125 (N_18125,N_11713,N_12798);
nor U18126 (N_18126,N_14780,N_12274);
xnor U18127 (N_18127,N_13706,N_11861);
or U18128 (N_18128,N_10378,N_13984);
or U18129 (N_18129,N_10434,N_10995);
or U18130 (N_18130,N_13139,N_12295);
xnor U18131 (N_18131,N_14855,N_10586);
xor U18132 (N_18132,N_10992,N_13923);
nor U18133 (N_18133,N_14516,N_12487);
nand U18134 (N_18134,N_10579,N_10627);
or U18135 (N_18135,N_10984,N_10846);
xnor U18136 (N_18136,N_14520,N_13552);
nand U18137 (N_18137,N_10230,N_14630);
and U18138 (N_18138,N_11093,N_12718);
and U18139 (N_18139,N_10148,N_11296);
nand U18140 (N_18140,N_11755,N_11735);
nor U18141 (N_18141,N_10038,N_12422);
xnor U18142 (N_18142,N_12341,N_10742);
or U18143 (N_18143,N_12603,N_11818);
nand U18144 (N_18144,N_14940,N_10553);
nor U18145 (N_18145,N_10950,N_12382);
nor U18146 (N_18146,N_10409,N_10994);
xor U18147 (N_18147,N_12186,N_14240);
and U18148 (N_18148,N_13552,N_10444);
or U18149 (N_18149,N_12891,N_11424);
or U18150 (N_18150,N_10180,N_13572);
nor U18151 (N_18151,N_13007,N_14087);
nand U18152 (N_18152,N_14796,N_10362);
or U18153 (N_18153,N_11693,N_14091);
xor U18154 (N_18154,N_14493,N_14260);
or U18155 (N_18155,N_11399,N_12622);
nor U18156 (N_18156,N_10959,N_12749);
nand U18157 (N_18157,N_12732,N_12514);
xor U18158 (N_18158,N_12483,N_14640);
nor U18159 (N_18159,N_12876,N_13298);
or U18160 (N_18160,N_13327,N_10822);
nand U18161 (N_18161,N_10680,N_10839);
xnor U18162 (N_18162,N_12697,N_10424);
nor U18163 (N_18163,N_13630,N_12296);
nand U18164 (N_18164,N_13108,N_11120);
or U18165 (N_18165,N_11854,N_13526);
nor U18166 (N_18166,N_11697,N_14426);
or U18167 (N_18167,N_12924,N_10392);
and U18168 (N_18168,N_13856,N_12806);
nand U18169 (N_18169,N_14528,N_14069);
nor U18170 (N_18170,N_12823,N_14640);
or U18171 (N_18171,N_10624,N_10651);
nand U18172 (N_18172,N_13685,N_12366);
or U18173 (N_18173,N_12270,N_12730);
or U18174 (N_18174,N_14841,N_11837);
nand U18175 (N_18175,N_10028,N_10462);
or U18176 (N_18176,N_10978,N_14451);
nor U18177 (N_18177,N_10253,N_13524);
or U18178 (N_18178,N_13715,N_12365);
nor U18179 (N_18179,N_13824,N_11600);
and U18180 (N_18180,N_12172,N_12949);
and U18181 (N_18181,N_13005,N_11463);
xnor U18182 (N_18182,N_10361,N_13917);
xnor U18183 (N_18183,N_14337,N_10778);
xnor U18184 (N_18184,N_12235,N_13653);
nand U18185 (N_18185,N_10692,N_10391);
nand U18186 (N_18186,N_13345,N_13334);
and U18187 (N_18187,N_13992,N_14929);
and U18188 (N_18188,N_10904,N_13733);
nor U18189 (N_18189,N_10074,N_13262);
and U18190 (N_18190,N_11890,N_12971);
and U18191 (N_18191,N_13378,N_13797);
or U18192 (N_18192,N_11791,N_10272);
nor U18193 (N_18193,N_12092,N_11399);
xnor U18194 (N_18194,N_12836,N_11115);
or U18195 (N_18195,N_12740,N_10648);
or U18196 (N_18196,N_13584,N_14475);
and U18197 (N_18197,N_11160,N_11119);
xnor U18198 (N_18198,N_11886,N_12214);
xnor U18199 (N_18199,N_14997,N_12311);
nor U18200 (N_18200,N_10659,N_13946);
and U18201 (N_18201,N_14568,N_13599);
nand U18202 (N_18202,N_12097,N_13329);
and U18203 (N_18203,N_14076,N_12785);
xor U18204 (N_18204,N_13199,N_13111);
xnor U18205 (N_18205,N_13029,N_11328);
and U18206 (N_18206,N_13777,N_12978);
xor U18207 (N_18207,N_12693,N_12014);
and U18208 (N_18208,N_13619,N_11604);
or U18209 (N_18209,N_10839,N_12764);
nor U18210 (N_18210,N_14850,N_14620);
nand U18211 (N_18211,N_12678,N_10893);
nand U18212 (N_18212,N_11095,N_12857);
or U18213 (N_18213,N_12850,N_12437);
nor U18214 (N_18214,N_14039,N_11181);
nand U18215 (N_18215,N_11579,N_10206);
and U18216 (N_18216,N_10683,N_13746);
and U18217 (N_18217,N_13879,N_10765);
and U18218 (N_18218,N_14282,N_11471);
and U18219 (N_18219,N_11276,N_14799);
and U18220 (N_18220,N_11930,N_12540);
nand U18221 (N_18221,N_13436,N_10393);
and U18222 (N_18222,N_14566,N_13093);
or U18223 (N_18223,N_11336,N_12136);
and U18224 (N_18224,N_10496,N_11572);
or U18225 (N_18225,N_12391,N_10333);
or U18226 (N_18226,N_10605,N_11515);
xor U18227 (N_18227,N_14798,N_13521);
and U18228 (N_18228,N_12207,N_10107);
and U18229 (N_18229,N_10993,N_10112);
nor U18230 (N_18230,N_12565,N_14268);
nand U18231 (N_18231,N_11841,N_11338);
xor U18232 (N_18232,N_13895,N_14095);
nor U18233 (N_18233,N_11104,N_14132);
nand U18234 (N_18234,N_13804,N_13333);
xnor U18235 (N_18235,N_10233,N_13043);
or U18236 (N_18236,N_14052,N_12248);
nand U18237 (N_18237,N_11636,N_10611);
and U18238 (N_18238,N_14716,N_12374);
xor U18239 (N_18239,N_13103,N_12410);
and U18240 (N_18240,N_13743,N_13300);
xnor U18241 (N_18241,N_11629,N_14866);
xnor U18242 (N_18242,N_12365,N_10035);
nor U18243 (N_18243,N_12988,N_13023);
xnor U18244 (N_18244,N_13233,N_11691);
or U18245 (N_18245,N_10715,N_11631);
and U18246 (N_18246,N_12838,N_12956);
nand U18247 (N_18247,N_12391,N_14069);
nand U18248 (N_18248,N_10821,N_10466);
nor U18249 (N_18249,N_10544,N_14091);
nor U18250 (N_18250,N_14785,N_11115);
or U18251 (N_18251,N_11720,N_14200);
nor U18252 (N_18252,N_10281,N_12359);
or U18253 (N_18253,N_12367,N_12337);
or U18254 (N_18254,N_13958,N_11542);
nor U18255 (N_18255,N_12958,N_13710);
or U18256 (N_18256,N_11057,N_11178);
nor U18257 (N_18257,N_11510,N_12541);
nor U18258 (N_18258,N_11057,N_12819);
nand U18259 (N_18259,N_12561,N_12178);
and U18260 (N_18260,N_10778,N_10614);
and U18261 (N_18261,N_12906,N_14650);
or U18262 (N_18262,N_12085,N_10316);
xor U18263 (N_18263,N_12631,N_11242);
and U18264 (N_18264,N_13524,N_13731);
nor U18265 (N_18265,N_10536,N_13625);
xor U18266 (N_18266,N_10864,N_14174);
nand U18267 (N_18267,N_14967,N_11353);
nor U18268 (N_18268,N_12454,N_13189);
nor U18269 (N_18269,N_13750,N_10267);
or U18270 (N_18270,N_12424,N_10540);
nand U18271 (N_18271,N_12051,N_10808);
xor U18272 (N_18272,N_12936,N_12263);
nor U18273 (N_18273,N_13588,N_10857);
xor U18274 (N_18274,N_11116,N_12988);
and U18275 (N_18275,N_12177,N_14309);
nand U18276 (N_18276,N_12295,N_12659);
or U18277 (N_18277,N_11086,N_10832);
nor U18278 (N_18278,N_10486,N_11707);
or U18279 (N_18279,N_13365,N_13890);
and U18280 (N_18280,N_12507,N_13839);
and U18281 (N_18281,N_10120,N_10953);
nand U18282 (N_18282,N_11897,N_14804);
nand U18283 (N_18283,N_13552,N_14893);
nand U18284 (N_18284,N_12756,N_10702);
nand U18285 (N_18285,N_12167,N_12271);
nor U18286 (N_18286,N_10352,N_14236);
nor U18287 (N_18287,N_12204,N_11711);
or U18288 (N_18288,N_13761,N_10458);
nand U18289 (N_18289,N_10270,N_13118);
nand U18290 (N_18290,N_10394,N_13700);
xor U18291 (N_18291,N_14871,N_10237);
nor U18292 (N_18292,N_10260,N_14583);
nor U18293 (N_18293,N_10441,N_10123);
or U18294 (N_18294,N_10760,N_14141);
nor U18295 (N_18295,N_12375,N_14604);
xnor U18296 (N_18296,N_12221,N_12285);
nor U18297 (N_18297,N_13254,N_12090);
nand U18298 (N_18298,N_14849,N_11931);
xor U18299 (N_18299,N_14061,N_10018);
xor U18300 (N_18300,N_13583,N_13260);
nand U18301 (N_18301,N_13352,N_10985);
nand U18302 (N_18302,N_14296,N_12421);
xor U18303 (N_18303,N_10127,N_14638);
or U18304 (N_18304,N_14466,N_14819);
or U18305 (N_18305,N_14885,N_13955);
and U18306 (N_18306,N_13123,N_13247);
xor U18307 (N_18307,N_10859,N_13419);
nor U18308 (N_18308,N_14476,N_10801);
or U18309 (N_18309,N_14599,N_10077);
nor U18310 (N_18310,N_13000,N_10752);
and U18311 (N_18311,N_12313,N_14315);
nand U18312 (N_18312,N_14069,N_13873);
nand U18313 (N_18313,N_11488,N_14366);
nand U18314 (N_18314,N_10275,N_12765);
xnor U18315 (N_18315,N_14684,N_11714);
or U18316 (N_18316,N_10530,N_11591);
or U18317 (N_18317,N_11622,N_14285);
xor U18318 (N_18318,N_10766,N_13919);
nor U18319 (N_18319,N_10227,N_13777);
and U18320 (N_18320,N_11324,N_13919);
nor U18321 (N_18321,N_10888,N_11970);
nand U18322 (N_18322,N_10032,N_13942);
and U18323 (N_18323,N_14248,N_11170);
or U18324 (N_18324,N_13519,N_12739);
or U18325 (N_18325,N_10377,N_12936);
nor U18326 (N_18326,N_13125,N_10528);
and U18327 (N_18327,N_14000,N_11291);
nand U18328 (N_18328,N_11348,N_12763);
xor U18329 (N_18329,N_12377,N_10572);
nand U18330 (N_18330,N_11109,N_11448);
nor U18331 (N_18331,N_14164,N_11430);
or U18332 (N_18332,N_11319,N_11978);
or U18333 (N_18333,N_13206,N_13708);
nor U18334 (N_18334,N_14225,N_12141);
nand U18335 (N_18335,N_10811,N_11684);
or U18336 (N_18336,N_11707,N_13730);
and U18337 (N_18337,N_13739,N_13050);
or U18338 (N_18338,N_12816,N_14965);
nand U18339 (N_18339,N_14002,N_14088);
and U18340 (N_18340,N_10975,N_13650);
nand U18341 (N_18341,N_10056,N_13593);
nor U18342 (N_18342,N_14467,N_10968);
nor U18343 (N_18343,N_14840,N_12504);
xnor U18344 (N_18344,N_13705,N_14566);
nor U18345 (N_18345,N_13585,N_10835);
xor U18346 (N_18346,N_14217,N_10095);
nand U18347 (N_18347,N_10027,N_13355);
or U18348 (N_18348,N_12409,N_12266);
and U18349 (N_18349,N_12146,N_14108);
nor U18350 (N_18350,N_11415,N_10769);
xor U18351 (N_18351,N_11775,N_12966);
and U18352 (N_18352,N_14163,N_13046);
nor U18353 (N_18353,N_12000,N_13877);
nand U18354 (N_18354,N_11673,N_11044);
nor U18355 (N_18355,N_13893,N_13443);
and U18356 (N_18356,N_11104,N_10186);
or U18357 (N_18357,N_12756,N_10067);
nor U18358 (N_18358,N_11099,N_11267);
nand U18359 (N_18359,N_14147,N_10144);
nor U18360 (N_18360,N_10995,N_13522);
and U18361 (N_18361,N_10421,N_11084);
or U18362 (N_18362,N_10642,N_12126);
and U18363 (N_18363,N_13849,N_14831);
xnor U18364 (N_18364,N_10726,N_11628);
or U18365 (N_18365,N_14597,N_14990);
xor U18366 (N_18366,N_14333,N_13862);
and U18367 (N_18367,N_12083,N_11238);
xnor U18368 (N_18368,N_11139,N_12280);
and U18369 (N_18369,N_13999,N_13114);
and U18370 (N_18370,N_13740,N_12196);
and U18371 (N_18371,N_11376,N_11100);
and U18372 (N_18372,N_13913,N_11691);
and U18373 (N_18373,N_13640,N_10585);
xor U18374 (N_18374,N_10720,N_14048);
xor U18375 (N_18375,N_12423,N_13653);
or U18376 (N_18376,N_12020,N_10379);
and U18377 (N_18377,N_13577,N_11568);
nor U18378 (N_18378,N_14260,N_13845);
nand U18379 (N_18379,N_11340,N_12827);
and U18380 (N_18380,N_14452,N_11280);
xor U18381 (N_18381,N_12298,N_10815);
nand U18382 (N_18382,N_14274,N_12879);
nand U18383 (N_18383,N_14492,N_10658);
and U18384 (N_18384,N_14993,N_13305);
xnor U18385 (N_18385,N_14110,N_11188);
or U18386 (N_18386,N_12884,N_12898);
nor U18387 (N_18387,N_12718,N_12265);
or U18388 (N_18388,N_12234,N_10074);
or U18389 (N_18389,N_12274,N_10873);
xnor U18390 (N_18390,N_11987,N_13281);
and U18391 (N_18391,N_13606,N_11944);
and U18392 (N_18392,N_12740,N_14036);
nand U18393 (N_18393,N_14531,N_14374);
and U18394 (N_18394,N_10485,N_12701);
xnor U18395 (N_18395,N_10479,N_12335);
nor U18396 (N_18396,N_14451,N_14689);
and U18397 (N_18397,N_12823,N_12929);
nand U18398 (N_18398,N_14668,N_10882);
nand U18399 (N_18399,N_12510,N_13488);
xor U18400 (N_18400,N_13283,N_12965);
nor U18401 (N_18401,N_12621,N_13961);
nor U18402 (N_18402,N_13367,N_14618);
or U18403 (N_18403,N_13044,N_12993);
nand U18404 (N_18404,N_12546,N_14544);
or U18405 (N_18405,N_11651,N_13486);
nor U18406 (N_18406,N_11733,N_12613);
or U18407 (N_18407,N_14672,N_13524);
or U18408 (N_18408,N_12550,N_11967);
and U18409 (N_18409,N_11263,N_13391);
nand U18410 (N_18410,N_10693,N_11396);
or U18411 (N_18411,N_12445,N_11226);
nand U18412 (N_18412,N_11605,N_13394);
nand U18413 (N_18413,N_11005,N_11619);
nor U18414 (N_18414,N_13371,N_11497);
nor U18415 (N_18415,N_10036,N_13735);
or U18416 (N_18416,N_12710,N_13486);
and U18417 (N_18417,N_14663,N_11531);
nand U18418 (N_18418,N_11794,N_13992);
nand U18419 (N_18419,N_12670,N_12198);
nor U18420 (N_18420,N_10936,N_11425);
or U18421 (N_18421,N_14808,N_13725);
xnor U18422 (N_18422,N_13841,N_10498);
xor U18423 (N_18423,N_11183,N_14478);
xnor U18424 (N_18424,N_10807,N_14401);
xor U18425 (N_18425,N_10633,N_14898);
and U18426 (N_18426,N_13790,N_10898);
and U18427 (N_18427,N_11678,N_11197);
xor U18428 (N_18428,N_11739,N_12462);
nand U18429 (N_18429,N_12151,N_11968);
xnor U18430 (N_18430,N_14454,N_11684);
or U18431 (N_18431,N_13910,N_13574);
or U18432 (N_18432,N_14566,N_14019);
or U18433 (N_18433,N_13146,N_11045);
nor U18434 (N_18434,N_11157,N_14550);
xor U18435 (N_18435,N_12457,N_12041);
and U18436 (N_18436,N_10753,N_14376);
nor U18437 (N_18437,N_11586,N_10759);
xor U18438 (N_18438,N_13057,N_13710);
xnor U18439 (N_18439,N_10254,N_11200);
xnor U18440 (N_18440,N_12083,N_10676);
nor U18441 (N_18441,N_11073,N_11221);
nand U18442 (N_18442,N_13195,N_12076);
nand U18443 (N_18443,N_12780,N_13359);
xor U18444 (N_18444,N_14904,N_13789);
and U18445 (N_18445,N_10313,N_14546);
nand U18446 (N_18446,N_10330,N_13367);
and U18447 (N_18447,N_12529,N_12618);
xor U18448 (N_18448,N_14847,N_13119);
xor U18449 (N_18449,N_14712,N_14236);
nor U18450 (N_18450,N_13930,N_10696);
xor U18451 (N_18451,N_10651,N_11923);
nor U18452 (N_18452,N_11010,N_12655);
nand U18453 (N_18453,N_13405,N_10609);
or U18454 (N_18454,N_12809,N_10474);
or U18455 (N_18455,N_11332,N_10364);
and U18456 (N_18456,N_13131,N_13817);
nand U18457 (N_18457,N_10844,N_13476);
xnor U18458 (N_18458,N_11571,N_10062);
nand U18459 (N_18459,N_12744,N_14125);
or U18460 (N_18460,N_12044,N_14347);
and U18461 (N_18461,N_11683,N_12878);
nand U18462 (N_18462,N_10034,N_11509);
xor U18463 (N_18463,N_14016,N_13299);
or U18464 (N_18464,N_13523,N_10316);
nand U18465 (N_18465,N_12260,N_13765);
nor U18466 (N_18466,N_11941,N_14101);
nor U18467 (N_18467,N_10529,N_13151);
or U18468 (N_18468,N_12398,N_10328);
or U18469 (N_18469,N_12813,N_12122);
and U18470 (N_18470,N_12818,N_11552);
xnor U18471 (N_18471,N_13516,N_13993);
and U18472 (N_18472,N_10444,N_10371);
or U18473 (N_18473,N_11637,N_14813);
nor U18474 (N_18474,N_10711,N_10500);
and U18475 (N_18475,N_12730,N_12906);
xnor U18476 (N_18476,N_13665,N_13558);
and U18477 (N_18477,N_13340,N_12764);
xor U18478 (N_18478,N_12643,N_13892);
xnor U18479 (N_18479,N_12218,N_14597);
and U18480 (N_18480,N_10019,N_10043);
xnor U18481 (N_18481,N_13533,N_13075);
xor U18482 (N_18482,N_13987,N_13691);
xor U18483 (N_18483,N_11790,N_13581);
and U18484 (N_18484,N_13550,N_14356);
xor U18485 (N_18485,N_11247,N_10327);
nor U18486 (N_18486,N_10643,N_11170);
nor U18487 (N_18487,N_13186,N_10463);
or U18488 (N_18488,N_13681,N_10747);
and U18489 (N_18489,N_10604,N_14048);
nand U18490 (N_18490,N_12129,N_10113);
and U18491 (N_18491,N_12973,N_11365);
nand U18492 (N_18492,N_10883,N_12379);
or U18493 (N_18493,N_10282,N_14256);
and U18494 (N_18494,N_13091,N_14728);
nor U18495 (N_18495,N_13433,N_11569);
nor U18496 (N_18496,N_12593,N_14428);
xnor U18497 (N_18497,N_14356,N_12477);
and U18498 (N_18498,N_12992,N_11263);
nor U18499 (N_18499,N_13271,N_13546);
nor U18500 (N_18500,N_11827,N_13326);
nand U18501 (N_18501,N_13049,N_10259);
nand U18502 (N_18502,N_13680,N_10706);
nand U18503 (N_18503,N_13552,N_10647);
and U18504 (N_18504,N_11474,N_13530);
nand U18505 (N_18505,N_11885,N_11482);
xnor U18506 (N_18506,N_14734,N_13837);
and U18507 (N_18507,N_11056,N_13436);
and U18508 (N_18508,N_12715,N_12770);
xnor U18509 (N_18509,N_14500,N_10419);
nor U18510 (N_18510,N_12912,N_10944);
nor U18511 (N_18511,N_10502,N_11227);
nand U18512 (N_18512,N_11569,N_12415);
nand U18513 (N_18513,N_14992,N_10515);
xor U18514 (N_18514,N_11011,N_14670);
or U18515 (N_18515,N_14642,N_11086);
or U18516 (N_18516,N_13881,N_11740);
nand U18517 (N_18517,N_14411,N_13882);
xor U18518 (N_18518,N_14829,N_10549);
xnor U18519 (N_18519,N_11115,N_14265);
nor U18520 (N_18520,N_12579,N_11560);
nand U18521 (N_18521,N_11118,N_14350);
nand U18522 (N_18522,N_11299,N_10329);
and U18523 (N_18523,N_10860,N_12485);
nand U18524 (N_18524,N_10556,N_11679);
or U18525 (N_18525,N_14847,N_12420);
or U18526 (N_18526,N_14402,N_11568);
and U18527 (N_18527,N_11105,N_11828);
xor U18528 (N_18528,N_14139,N_14965);
xor U18529 (N_18529,N_13110,N_11305);
nor U18530 (N_18530,N_14359,N_11213);
nor U18531 (N_18531,N_10605,N_11808);
and U18532 (N_18532,N_10618,N_13592);
and U18533 (N_18533,N_14354,N_14785);
or U18534 (N_18534,N_11962,N_11431);
and U18535 (N_18535,N_10754,N_14254);
or U18536 (N_18536,N_14203,N_12683);
or U18537 (N_18537,N_10388,N_11040);
and U18538 (N_18538,N_13034,N_10891);
xnor U18539 (N_18539,N_11500,N_10584);
xnor U18540 (N_18540,N_12988,N_11489);
nand U18541 (N_18541,N_11619,N_12652);
xnor U18542 (N_18542,N_10544,N_13435);
xor U18543 (N_18543,N_11279,N_10742);
and U18544 (N_18544,N_13089,N_10611);
or U18545 (N_18545,N_10689,N_13437);
or U18546 (N_18546,N_13738,N_13611);
nor U18547 (N_18547,N_11418,N_13011);
nand U18548 (N_18548,N_11657,N_13424);
xor U18549 (N_18549,N_12055,N_12184);
and U18550 (N_18550,N_10147,N_14231);
and U18551 (N_18551,N_12226,N_11754);
xnor U18552 (N_18552,N_11805,N_11891);
and U18553 (N_18553,N_13189,N_10318);
nor U18554 (N_18554,N_14660,N_12025);
nor U18555 (N_18555,N_14454,N_11958);
or U18556 (N_18556,N_13505,N_14324);
nor U18557 (N_18557,N_12284,N_14292);
xor U18558 (N_18558,N_14259,N_10319);
nor U18559 (N_18559,N_12732,N_11625);
nand U18560 (N_18560,N_11578,N_14914);
nand U18561 (N_18561,N_13263,N_14289);
or U18562 (N_18562,N_11553,N_14110);
nor U18563 (N_18563,N_14522,N_12783);
xor U18564 (N_18564,N_11462,N_12770);
and U18565 (N_18565,N_12549,N_11413);
and U18566 (N_18566,N_12071,N_13727);
xnor U18567 (N_18567,N_11526,N_10011);
and U18568 (N_18568,N_13032,N_13624);
nand U18569 (N_18569,N_10817,N_14836);
and U18570 (N_18570,N_13264,N_10032);
xor U18571 (N_18571,N_13167,N_13934);
or U18572 (N_18572,N_11549,N_12523);
nand U18573 (N_18573,N_12278,N_10216);
or U18574 (N_18574,N_12130,N_13774);
nand U18575 (N_18575,N_10751,N_11117);
and U18576 (N_18576,N_10034,N_10025);
and U18577 (N_18577,N_12452,N_13771);
nand U18578 (N_18578,N_11906,N_10350);
nand U18579 (N_18579,N_11227,N_12529);
nand U18580 (N_18580,N_10713,N_13221);
nor U18581 (N_18581,N_11482,N_10910);
or U18582 (N_18582,N_11237,N_10964);
xor U18583 (N_18583,N_13270,N_11893);
or U18584 (N_18584,N_12277,N_13419);
or U18585 (N_18585,N_13945,N_11215);
nor U18586 (N_18586,N_11661,N_14987);
and U18587 (N_18587,N_12284,N_10679);
xnor U18588 (N_18588,N_14645,N_11033);
or U18589 (N_18589,N_10586,N_13010);
xnor U18590 (N_18590,N_12909,N_11173);
or U18591 (N_18591,N_13629,N_10520);
nand U18592 (N_18592,N_11943,N_14908);
and U18593 (N_18593,N_10027,N_12455);
or U18594 (N_18594,N_14935,N_13693);
nand U18595 (N_18595,N_14278,N_11014);
xnor U18596 (N_18596,N_10045,N_12349);
or U18597 (N_18597,N_11639,N_10417);
nand U18598 (N_18598,N_14054,N_12879);
xnor U18599 (N_18599,N_10642,N_11569);
or U18600 (N_18600,N_14522,N_12751);
or U18601 (N_18601,N_14743,N_13925);
nor U18602 (N_18602,N_14536,N_13512);
and U18603 (N_18603,N_11991,N_12578);
xnor U18604 (N_18604,N_13674,N_14042);
nor U18605 (N_18605,N_10628,N_11763);
nand U18606 (N_18606,N_10187,N_12989);
xnor U18607 (N_18607,N_10789,N_10425);
and U18608 (N_18608,N_12751,N_10027);
and U18609 (N_18609,N_13152,N_12066);
nand U18610 (N_18610,N_12908,N_12870);
or U18611 (N_18611,N_10836,N_13192);
nor U18612 (N_18612,N_10819,N_13811);
and U18613 (N_18613,N_13750,N_10014);
nor U18614 (N_18614,N_14844,N_12136);
and U18615 (N_18615,N_14822,N_14620);
and U18616 (N_18616,N_14523,N_12851);
nand U18617 (N_18617,N_14323,N_13427);
and U18618 (N_18618,N_12979,N_12944);
and U18619 (N_18619,N_14416,N_12584);
nor U18620 (N_18620,N_14445,N_12975);
xor U18621 (N_18621,N_13947,N_12535);
xnor U18622 (N_18622,N_12870,N_14108);
or U18623 (N_18623,N_13057,N_10401);
nand U18624 (N_18624,N_10469,N_14006);
xor U18625 (N_18625,N_13804,N_10995);
or U18626 (N_18626,N_10301,N_12228);
or U18627 (N_18627,N_14968,N_12446);
xnor U18628 (N_18628,N_14053,N_12895);
xor U18629 (N_18629,N_14587,N_12823);
nor U18630 (N_18630,N_13986,N_12402);
nand U18631 (N_18631,N_13010,N_11725);
nand U18632 (N_18632,N_11541,N_12069);
nor U18633 (N_18633,N_12649,N_14711);
or U18634 (N_18634,N_14254,N_10446);
and U18635 (N_18635,N_14765,N_10176);
nor U18636 (N_18636,N_14850,N_11392);
xor U18637 (N_18637,N_10522,N_10459);
or U18638 (N_18638,N_11254,N_11488);
nand U18639 (N_18639,N_14915,N_11265);
and U18640 (N_18640,N_14534,N_11388);
and U18641 (N_18641,N_11975,N_11578);
nor U18642 (N_18642,N_14929,N_14074);
nand U18643 (N_18643,N_13590,N_13567);
nand U18644 (N_18644,N_10196,N_13244);
and U18645 (N_18645,N_11876,N_13711);
xnor U18646 (N_18646,N_12308,N_12461);
or U18647 (N_18647,N_10151,N_14069);
xnor U18648 (N_18648,N_12816,N_14191);
nand U18649 (N_18649,N_12145,N_13539);
or U18650 (N_18650,N_11235,N_13966);
or U18651 (N_18651,N_11397,N_11520);
nand U18652 (N_18652,N_11728,N_14950);
and U18653 (N_18653,N_14358,N_13472);
nand U18654 (N_18654,N_12089,N_13681);
or U18655 (N_18655,N_14590,N_12895);
or U18656 (N_18656,N_14134,N_14704);
or U18657 (N_18657,N_12662,N_13659);
and U18658 (N_18658,N_12423,N_14611);
and U18659 (N_18659,N_12492,N_12795);
xnor U18660 (N_18660,N_10243,N_12657);
nor U18661 (N_18661,N_11114,N_13173);
nand U18662 (N_18662,N_12688,N_13131);
nor U18663 (N_18663,N_13092,N_14296);
xnor U18664 (N_18664,N_12681,N_13516);
nor U18665 (N_18665,N_10492,N_13389);
nand U18666 (N_18666,N_12794,N_11758);
or U18667 (N_18667,N_10948,N_12119);
xor U18668 (N_18668,N_12934,N_12466);
nand U18669 (N_18669,N_13006,N_14047);
or U18670 (N_18670,N_11150,N_12008);
nand U18671 (N_18671,N_14954,N_13067);
and U18672 (N_18672,N_11097,N_14499);
nand U18673 (N_18673,N_11350,N_13147);
or U18674 (N_18674,N_11179,N_11191);
nor U18675 (N_18675,N_13346,N_12812);
or U18676 (N_18676,N_10165,N_13036);
or U18677 (N_18677,N_10790,N_11509);
xnor U18678 (N_18678,N_14320,N_13468);
nand U18679 (N_18679,N_10978,N_13552);
and U18680 (N_18680,N_10448,N_11150);
xor U18681 (N_18681,N_14770,N_12924);
or U18682 (N_18682,N_14428,N_12980);
xor U18683 (N_18683,N_14289,N_10979);
nand U18684 (N_18684,N_13193,N_12477);
nand U18685 (N_18685,N_10231,N_12801);
nand U18686 (N_18686,N_12448,N_11292);
xnor U18687 (N_18687,N_11184,N_14464);
or U18688 (N_18688,N_13616,N_12485);
nand U18689 (N_18689,N_10427,N_10442);
xor U18690 (N_18690,N_13226,N_14107);
nor U18691 (N_18691,N_14401,N_10154);
or U18692 (N_18692,N_11484,N_13861);
or U18693 (N_18693,N_14008,N_14157);
xnor U18694 (N_18694,N_10168,N_14604);
nor U18695 (N_18695,N_14856,N_10125);
and U18696 (N_18696,N_14798,N_12604);
nand U18697 (N_18697,N_13120,N_11967);
or U18698 (N_18698,N_14930,N_13333);
nand U18699 (N_18699,N_13383,N_12705);
and U18700 (N_18700,N_11404,N_14485);
xor U18701 (N_18701,N_13645,N_11865);
or U18702 (N_18702,N_14638,N_14675);
or U18703 (N_18703,N_12642,N_14488);
nor U18704 (N_18704,N_13636,N_13872);
nor U18705 (N_18705,N_12789,N_14947);
and U18706 (N_18706,N_12806,N_11453);
nand U18707 (N_18707,N_10484,N_10780);
xnor U18708 (N_18708,N_13623,N_13367);
nand U18709 (N_18709,N_10815,N_11705);
xor U18710 (N_18710,N_10348,N_10855);
nor U18711 (N_18711,N_10446,N_14851);
xnor U18712 (N_18712,N_11523,N_13654);
and U18713 (N_18713,N_11622,N_14778);
nand U18714 (N_18714,N_10331,N_14809);
and U18715 (N_18715,N_14557,N_13396);
xnor U18716 (N_18716,N_14655,N_10249);
xor U18717 (N_18717,N_12929,N_10155);
nand U18718 (N_18718,N_14647,N_14244);
nand U18719 (N_18719,N_12881,N_11714);
nor U18720 (N_18720,N_12329,N_14565);
xnor U18721 (N_18721,N_11541,N_13780);
and U18722 (N_18722,N_14134,N_13766);
and U18723 (N_18723,N_10475,N_13831);
xnor U18724 (N_18724,N_13048,N_11540);
or U18725 (N_18725,N_12917,N_12771);
xor U18726 (N_18726,N_10617,N_13269);
and U18727 (N_18727,N_12635,N_14268);
nor U18728 (N_18728,N_13110,N_12053);
nand U18729 (N_18729,N_13744,N_11797);
and U18730 (N_18730,N_12681,N_10713);
nor U18731 (N_18731,N_10517,N_11872);
nand U18732 (N_18732,N_12938,N_14085);
nor U18733 (N_18733,N_11530,N_10292);
nand U18734 (N_18734,N_14926,N_11021);
nor U18735 (N_18735,N_11967,N_11505);
xor U18736 (N_18736,N_12634,N_11488);
xnor U18737 (N_18737,N_12788,N_11433);
nor U18738 (N_18738,N_14995,N_14119);
or U18739 (N_18739,N_11430,N_11824);
xnor U18740 (N_18740,N_13641,N_10425);
nor U18741 (N_18741,N_12021,N_14729);
and U18742 (N_18742,N_10014,N_10475);
or U18743 (N_18743,N_12057,N_11819);
or U18744 (N_18744,N_12515,N_11596);
nand U18745 (N_18745,N_10118,N_13579);
nand U18746 (N_18746,N_11088,N_11269);
nor U18747 (N_18747,N_13949,N_14596);
nand U18748 (N_18748,N_12310,N_11358);
xor U18749 (N_18749,N_14478,N_10268);
nor U18750 (N_18750,N_11999,N_12444);
nor U18751 (N_18751,N_13210,N_11850);
nand U18752 (N_18752,N_12981,N_12370);
xor U18753 (N_18753,N_13045,N_13511);
nor U18754 (N_18754,N_13044,N_12303);
nor U18755 (N_18755,N_10088,N_10900);
nor U18756 (N_18756,N_13408,N_14648);
nor U18757 (N_18757,N_10746,N_12106);
and U18758 (N_18758,N_10490,N_12378);
or U18759 (N_18759,N_12267,N_13204);
xor U18760 (N_18760,N_11451,N_13541);
and U18761 (N_18761,N_12049,N_12108);
xnor U18762 (N_18762,N_10517,N_12966);
and U18763 (N_18763,N_14037,N_12606);
and U18764 (N_18764,N_13503,N_10533);
or U18765 (N_18765,N_11229,N_13481);
and U18766 (N_18766,N_14688,N_10174);
nand U18767 (N_18767,N_10111,N_13067);
nor U18768 (N_18768,N_12495,N_13739);
nor U18769 (N_18769,N_11999,N_12959);
xnor U18770 (N_18770,N_12417,N_14468);
nor U18771 (N_18771,N_11603,N_11791);
nor U18772 (N_18772,N_12329,N_11899);
or U18773 (N_18773,N_11607,N_10189);
or U18774 (N_18774,N_12296,N_10746);
and U18775 (N_18775,N_13447,N_13348);
xor U18776 (N_18776,N_12323,N_12369);
nand U18777 (N_18777,N_11616,N_11955);
and U18778 (N_18778,N_12864,N_10454);
nor U18779 (N_18779,N_12469,N_10777);
nand U18780 (N_18780,N_13872,N_13216);
and U18781 (N_18781,N_11884,N_11148);
and U18782 (N_18782,N_10998,N_10591);
xor U18783 (N_18783,N_10401,N_14588);
nand U18784 (N_18784,N_11428,N_11647);
nor U18785 (N_18785,N_13632,N_12142);
xnor U18786 (N_18786,N_13098,N_12174);
xnor U18787 (N_18787,N_13250,N_10832);
nand U18788 (N_18788,N_12191,N_10871);
or U18789 (N_18789,N_13302,N_13238);
and U18790 (N_18790,N_14264,N_13989);
xor U18791 (N_18791,N_14106,N_14490);
nand U18792 (N_18792,N_10775,N_10364);
xor U18793 (N_18793,N_12750,N_12228);
or U18794 (N_18794,N_10567,N_10560);
xnor U18795 (N_18795,N_10388,N_13618);
and U18796 (N_18796,N_13717,N_11050);
xnor U18797 (N_18797,N_14279,N_14651);
or U18798 (N_18798,N_10612,N_11920);
or U18799 (N_18799,N_14998,N_13105);
and U18800 (N_18800,N_13632,N_10632);
nand U18801 (N_18801,N_10067,N_13249);
or U18802 (N_18802,N_14702,N_13032);
nor U18803 (N_18803,N_12135,N_12387);
nand U18804 (N_18804,N_10955,N_13338);
nand U18805 (N_18805,N_14700,N_11231);
nand U18806 (N_18806,N_14013,N_11406);
xnor U18807 (N_18807,N_13279,N_11914);
nor U18808 (N_18808,N_13083,N_13298);
nand U18809 (N_18809,N_10052,N_11607);
nand U18810 (N_18810,N_14280,N_12999);
xnor U18811 (N_18811,N_14524,N_14893);
nor U18812 (N_18812,N_11097,N_14073);
xor U18813 (N_18813,N_12659,N_13379);
and U18814 (N_18814,N_11877,N_10846);
nor U18815 (N_18815,N_12675,N_10671);
nor U18816 (N_18816,N_13939,N_12226);
xnor U18817 (N_18817,N_13268,N_10060);
nand U18818 (N_18818,N_13290,N_13422);
or U18819 (N_18819,N_13352,N_12967);
nor U18820 (N_18820,N_12320,N_11503);
or U18821 (N_18821,N_13987,N_14651);
and U18822 (N_18822,N_13647,N_13391);
xor U18823 (N_18823,N_13769,N_10911);
nor U18824 (N_18824,N_13614,N_13189);
or U18825 (N_18825,N_13415,N_10417);
xnor U18826 (N_18826,N_11359,N_12500);
xnor U18827 (N_18827,N_11541,N_14076);
xor U18828 (N_18828,N_11954,N_11288);
nand U18829 (N_18829,N_11717,N_11031);
and U18830 (N_18830,N_14927,N_14268);
nand U18831 (N_18831,N_11329,N_11038);
xor U18832 (N_18832,N_11962,N_13888);
xnor U18833 (N_18833,N_10826,N_13762);
and U18834 (N_18834,N_13995,N_12804);
or U18835 (N_18835,N_11265,N_13956);
xnor U18836 (N_18836,N_13405,N_13443);
and U18837 (N_18837,N_14983,N_10533);
nand U18838 (N_18838,N_13052,N_13855);
and U18839 (N_18839,N_10227,N_11396);
and U18840 (N_18840,N_12611,N_12780);
nand U18841 (N_18841,N_12219,N_14227);
and U18842 (N_18842,N_12113,N_12815);
and U18843 (N_18843,N_14428,N_13306);
nor U18844 (N_18844,N_11922,N_10567);
xnor U18845 (N_18845,N_14491,N_10650);
and U18846 (N_18846,N_14342,N_11486);
xnor U18847 (N_18847,N_12200,N_11242);
nor U18848 (N_18848,N_13592,N_10952);
and U18849 (N_18849,N_11517,N_13732);
or U18850 (N_18850,N_13953,N_12860);
nor U18851 (N_18851,N_10534,N_11981);
nand U18852 (N_18852,N_13910,N_13391);
nor U18853 (N_18853,N_14012,N_13782);
or U18854 (N_18854,N_13470,N_12333);
nand U18855 (N_18855,N_10156,N_11014);
or U18856 (N_18856,N_11086,N_11258);
nand U18857 (N_18857,N_12246,N_10585);
or U18858 (N_18858,N_14382,N_13074);
or U18859 (N_18859,N_12071,N_12974);
xor U18860 (N_18860,N_13889,N_12109);
or U18861 (N_18861,N_14611,N_11951);
or U18862 (N_18862,N_12928,N_10094);
or U18863 (N_18863,N_13181,N_10840);
or U18864 (N_18864,N_11227,N_14382);
or U18865 (N_18865,N_11852,N_13133);
and U18866 (N_18866,N_12856,N_11276);
and U18867 (N_18867,N_12661,N_11061);
nand U18868 (N_18868,N_12352,N_10914);
and U18869 (N_18869,N_12286,N_11912);
nand U18870 (N_18870,N_14510,N_14035);
or U18871 (N_18871,N_11643,N_12215);
nor U18872 (N_18872,N_13331,N_11807);
nand U18873 (N_18873,N_11398,N_14493);
or U18874 (N_18874,N_12753,N_11129);
nand U18875 (N_18875,N_13611,N_14822);
or U18876 (N_18876,N_12466,N_11040);
xor U18877 (N_18877,N_13392,N_10564);
nand U18878 (N_18878,N_14444,N_10010);
nor U18879 (N_18879,N_11496,N_12871);
nand U18880 (N_18880,N_13914,N_13356);
xor U18881 (N_18881,N_14135,N_11113);
nor U18882 (N_18882,N_10046,N_13708);
and U18883 (N_18883,N_12566,N_11025);
and U18884 (N_18884,N_11779,N_14042);
nand U18885 (N_18885,N_13665,N_10678);
and U18886 (N_18886,N_10743,N_12446);
xnor U18887 (N_18887,N_12380,N_12483);
xnor U18888 (N_18888,N_14634,N_14526);
and U18889 (N_18889,N_10459,N_11410);
or U18890 (N_18890,N_11749,N_10362);
and U18891 (N_18891,N_13541,N_13748);
and U18892 (N_18892,N_11903,N_13506);
and U18893 (N_18893,N_13422,N_11530);
nor U18894 (N_18894,N_14589,N_11153);
xnor U18895 (N_18895,N_13395,N_11277);
and U18896 (N_18896,N_13887,N_10526);
xor U18897 (N_18897,N_11626,N_11298);
or U18898 (N_18898,N_12514,N_13261);
or U18899 (N_18899,N_11742,N_11242);
or U18900 (N_18900,N_14954,N_10521);
or U18901 (N_18901,N_10396,N_14872);
or U18902 (N_18902,N_14294,N_10360);
or U18903 (N_18903,N_13019,N_10904);
and U18904 (N_18904,N_12286,N_14778);
xor U18905 (N_18905,N_13847,N_14269);
nand U18906 (N_18906,N_12850,N_13267);
and U18907 (N_18907,N_13051,N_10614);
xor U18908 (N_18908,N_14584,N_10841);
nor U18909 (N_18909,N_12984,N_10694);
and U18910 (N_18910,N_12238,N_11995);
nor U18911 (N_18911,N_10417,N_10037);
or U18912 (N_18912,N_11395,N_12334);
nor U18913 (N_18913,N_11311,N_10694);
nor U18914 (N_18914,N_13307,N_11815);
nand U18915 (N_18915,N_13781,N_11657);
or U18916 (N_18916,N_11749,N_10798);
nand U18917 (N_18917,N_11793,N_12961);
and U18918 (N_18918,N_12178,N_14393);
and U18919 (N_18919,N_10798,N_14800);
or U18920 (N_18920,N_10847,N_13555);
nor U18921 (N_18921,N_14887,N_14043);
xor U18922 (N_18922,N_13200,N_12372);
and U18923 (N_18923,N_10336,N_12399);
xor U18924 (N_18924,N_10631,N_11714);
and U18925 (N_18925,N_10729,N_10393);
nor U18926 (N_18926,N_13026,N_10647);
and U18927 (N_18927,N_10187,N_11154);
nand U18928 (N_18928,N_10142,N_14845);
nor U18929 (N_18929,N_10098,N_10586);
nand U18930 (N_18930,N_13702,N_10912);
xor U18931 (N_18931,N_10316,N_10496);
and U18932 (N_18932,N_14845,N_12584);
nor U18933 (N_18933,N_12720,N_13725);
nor U18934 (N_18934,N_14214,N_13761);
or U18935 (N_18935,N_11012,N_12970);
or U18936 (N_18936,N_10913,N_13598);
and U18937 (N_18937,N_14025,N_12913);
and U18938 (N_18938,N_11029,N_12052);
and U18939 (N_18939,N_14191,N_10702);
nand U18940 (N_18940,N_13833,N_14133);
or U18941 (N_18941,N_14108,N_13250);
xor U18942 (N_18942,N_11842,N_12516);
xor U18943 (N_18943,N_13990,N_11160);
or U18944 (N_18944,N_11909,N_11753);
xnor U18945 (N_18945,N_11937,N_14236);
or U18946 (N_18946,N_12010,N_14649);
xor U18947 (N_18947,N_13388,N_10961);
or U18948 (N_18948,N_10388,N_13746);
xnor U18949 (N_18949,N_12391,N_10928);
nand U18950 (N_18950,N_11760,N_13541);
and U18951 (N_18951,N_11788,N_14008);
xor U18952 (N_18952,N_11229,N_13855);
or U18953 (N_18953,N_10036,N_14133);
and U18954 (N_18954,N_10419,N_14800);
nor U18955 (N_18955,N_12727,N_13458);
or U18956 (N_18956,N_13246,N_12499);
or U18957 (N_18957,N_11476,N_11888);
and U18958 (N_18958,N_14859,N_11988);
and U18959 (N_18959,N_14588,N_11789);
nor U18960 (N_18960,N_14280,N_14103);
xnor U18961 (N_18961,N_13183,N_13458);
nand U18962 (N_18962,N_11070,N_14198);
nand U18963 (N_18963,N_10804,N_13113);
nand U18964 (N_18964,N_12438,N_14272);
and U18965 (N_18965,N_13988,N_11474);
nor U18966 (N_18966,N_11827,N_11589);
nand U18967 (N_18967,N_12076,N_14895);
or U18968 (N_18968,N_13574,N_14890);
xnor U18969 (N_18969,N_14045,N_14469);
or U18970 (N_18970,N_12859,N_12814);
nand U18971 (N_18971,N_13922,N_12524);
nand U18972 (N_18972,N_10586,N_14849);
xnor U18973 (N_18973,N_14630,N_12627);
nand U18974 (N_18974,N_14572,N_13658);
and U18975 (N_18975,N_10582,N_13237);
nand U18976 (N_18976,N_13176,N_11148);
nand U18977 (N_18977,N_14191,N_10654);
nand U18978 (N_18978,N_14068,N_10913);
nand U18979 (N_18979,N_14937,N_14833);
and U18980 (N_18980,N_14711,N_10666);
xnor U18981 (N_18981,N_14021,N_14009);
nor U18982 (N_18982,N_13031,N_10838);
nand U18983 (N_18983,N_13447,N_10604);
nand U18984 (N_18984,N_10836,N_14465);
or U18985 (N_18985,N_11266,N_10993);
xnor U18986 (N_18986,N_10860,N_11980);
xnor U18987 (N_18987,N_11292,N_13738);
xnor U18988 (N_18988,N_13831,N_10352);
nand U18989 (N_18989,N_11108,N_14912);
nand U18990 (N_18990,N_12819,N_14606);
or U18991 (N_18991,N_12167,N_13402);
or U18992 (N_18992,N_12373,N_14049);
and U18993 (N_18993,N_13669,N_10455);
xor U18994 (N_18994,N_10734,N_11843);
nand U18995 (N_18995,N_10283,N_10517);
xnor U18996 (N_18996,N_11634,N_13506);
and U18997 (N_18997,N_11886,N_13406);
or U18998 (N_18998,N_10149,N_11925);
nand U18999 (N_18999,N_14877,N_13962);
or U19000 (N_19000,N_11527,N_11821);
and U19001 (N_19001,N_11251,N_12130);
nor U19002 (N_19002,N_10690,N_13270);
nor U19003 (N_19003,N_13934,N_12409);
and U19004 (N_19004,N_11133,N_12147);
xnor U19005 (N_19005,N_11192,N_11767);
nand U19006 (N_19006,N_14735,N_13631);
or U19007 (N_19007,N_12038,N_11197);
and U19008 (N_19008,N_14536,N_12799);
nor U19009 (N_19009,N_11588,N_11717);
or U19010 (N_19010,N_11789,N_14031);
xnor U19011 (N_19011,N_13027,N_13479);
nor U19012 (N_19012,N_10809,N_12161);
and U19013 (N_19013,N_11646,N_14003);
nor U19014 (N_19014,N_10547,N_12186);
and U19015 (N_19015,N_11991,N_14033);
nor U19016 (N_19016,N_14258,N_14279);
xnor U19017 (N_19017,N_10566,N_13564);
nor U19018 (N_19018,N_12748,N_12255);
and U19019 (N_19019,N_11649,N_12414);
and U19020 (N_19020,N_12962,N_10058);
and U19021 (N_19021,N_12214,N_12425);
or U19022 (N_19022,N_11341,N_10641);
or U19023 (N_19023,N_11090,N_14554);
nand U19024 (N_19024,N_11687,N_11814);
and U19025 (N_19025,N_11433,N_12231);
or U19026 (N_19026,N_13436,N_10458);
and U19027 (N_19027,N_11475,N_13354);
nand U19028 (N_19028,N_12241,N_12219);
and U19029 (N_19029,N_13048,N_14738);
nand U19030 (N_19030,N_14718,N_11964);
nor U19031 (N_19031,N_12429,N_10792);
nor U19032 (N_19032,N_14266,N_10178);
nor U19033 (N_19033,N_12150,N_13844);
xnor U19034 (N_19034,N_14299,N_14381);
nor U19035 (N_19035,N_12655,N_14711);
or U19036 (N_19036,N_13457,N_11031);
nor U19037 (N_19037,N_12009,N_13258);
nor U19038 (N_19038,N_10261,N_13735);
and U19039 (N_19039,N_13569,N_13484);
nand U19040 (N_19040,N_13214,N_13016);
and U19041 (N_19041,N_10214,N_12995);
or U19042 (N_19042,N_14621,N_14385);
nor U19043 (N_19043,N_13563,N_12981);
nand U19044 (N_19044,N_10957,N_11009);
nor U19045 (N_19045,N_11113,N_14423);
xor U19046 (N_19046,N_11988,N_14092);
or U19047 (N_19047,N_14749,N_12472);
nor U19048 (N_19048,N_11891,N_12962);
xor U19049 (N_19049,N_11587,N_10568);
nor U19050 (N_19050,N_14805,N_14881);
or U19051 (N_19051,N_11963,N_11054);
and U19052 (N_19052,N_10423,N_12634);
nor U19053 (N_19053,N_13016,N_10597);
or U19054 (N_19054,N_14708,N_10989);
nand U19055 (N_19055,N_10908,N_13511);
nand U19056 (N_19056,N_14363,N_12129);
or U19057 (N_19057,N_11045,N_13081);
nor U19058 (N_19058,N_14366,N_10251);
xor U19059 (N_19059,N_13109,N_13857);
nor U19060 (N_19060,N_14964,N_10278);
and U19061 (N_19061,N_13113,N_13832);
nor U19062 (N_19062,N_11804,N_12507);
nand U19063 (N_19063,N_12031,N_11961);
xor U19064 (N_19064,N_11341,N_10534);
xnor U19065 (N_19065,N_14405,N_10250);
nor U19066 (N_19066,N_10451,N_12423);
nor U19067 (N_19067,N_13868,N_11547);
nor U19068 (N_19068,N_11150,N_12977);
and U19069 (N_19069,N_14096,N_11145);
and U19070 (N_19070,N_14351,N_13729);
xor U19071 (N_19071,N_14046,N_11096);
xor U19072 (N_19072,N_14173,N_14539);
nor U19073 (N_19073,N_10442,N_10729);
nand U19074 (N_19074,N_10898,N_11996);
xnor U19075 (N_19075,N_14386,N_10857);
nand U19076 (N_19076,N_14322,N_12260);
nor U19077 (N_19077,N_10553,N_12638);
or U19078 (N_19078,N_13185,N_13726);
and U19079 (N_19079,N_13359,N_13143);
or U19080 (N_19080,N_14248,N_12907);
nand U19081 (N_19081,N_11796,N_11996);
nor U19082 (N_19082,N_12503,N_12875);
nand U19083 (N_19083,N_14253,N_14799);
nor U19084 (N_19084,N_11117,N_14482);
nand U19085 (N_19085,N_14337,N_13243);
nor U19086 (N_19086,N_13205,N_11676);
or U19087 (N_19087,N_10124,N_13182);
xor U19088 (N_19088,N_12418,N_10132);
nor U19089 (N_19089,N_13489,N_14945);
nand U19090 (N_19090,N_12923,N_10299);
xnor U19091 (N_19091,N_14793,N_12150);
nor U19092 (N_19092,N_13259,N_11653);
nand U19093 (N_19093,N_11565,N_12347);
xnor U19094 (N_19094,N_14735,N_13783);
nor U19095 (N_19095,N_11717,N_14891);
xnor U19096 (N_19096,N_14491,N_10738);
nor U19097 (N_19097,N_13224,N_13552);
and U19098 (N_19098,N_14851,N_12052);
and U19099 (N_19099,N_14567,N_14443);
xor U19100 (N_19100,N_11380,N_14168);
xor U19101 (N_19101,N_13392,N_11582);
or U19102 (N_19102,N_13289,N_10948);
and U19103 (N_19103,N_13186,N_13187);
or U19104 (N_19104,N_13582,N_11497);
and U19105 (N_19105,N_10496,N_13309);
nor U19106 (N_19106,N_13843,N_14105);
nand U19107 (N_19107,N_13658,N_13510);
xnor U19108 (N_19108,N_12073,N_10244);
xor U19109 (N_19109,N_14438,N_14411);
or U19110 (N_19110,N_14272,N_13910);
or U19111 (N_19111,N_11923,N_10252);
nand U19112 (N_19112,N_10863,N_13647);
or U19113 (N_19113,N_13849,N_14901);
or U19114 (N_19114,N_12974,N_10516);
nor U19115 (N_19115,N_13403,N_13882);
xnor U19116 (N_19116,N_10788,N_14479);
xnor U19117 (N_19117,N_10992,N_14289);
and U19118 (N_19118,N_11515,N_12583);
xor U19119 (N_19119,N_11794,N_10571);
xnor U19120 (N_19120,N_14581,N_12777);
or U19121 (N_19121,N_12126,N_14531);
or U19122 (N_19122,N_13899,N_12130);
nor U19123 (N_19123,N_12298,N_11570);
xnor U19124 (N_19124,N_14140,N_10832);
and U19125 (N_19125,N_10889,N_13554);
nor U19126 (N_19126,N_10005,N_14920);
xnor U19127 (N_19127,N_11101,N_10867);
or U19128 (N_19128,N_13451,N_11212);
nand U19129 (N_19129,N_12715,N_13169);
or U19130 (N_19130,N_12138,N_14809);
or U19131 (N_19131,N_13794,N_13450);
or U19132 (N_19132,N_12107,N_12570);
and U19133 (N_19133,N_13430,N_11454);
xor U19134 (N_19134,N_11399,N_12472);
xor U19135 (N_19135,N_12390,N_14296);
xor U19136 (N_19136,N_11306,N_14252);
xor U19137 (N_19137,N_13395,N_11609);
xnor U19138 (N_19138,N_10973,N_14157);
xor U19139 (N_19139,N_14253,N_12055);
xor U19140 (N_19140,N_11977,N_10772);
xnor U19141 (N_19141,N_13115,N_13219);
nor U19142 (N_19142,N_11294,N_10990);
xor U19143 (N_19143,N_14316,N_10022);
and U19144 (N_19144,N_14603,N_13122);
or U19145 (N_19145,N_11057,N_11635);
xor U19146 (N_19146,N_14437,N_12329);
or U19147 (N_19147,N_13623,N_13373);
or U19148 (N_19148,N_11168,N_13626);
or U19149 (N_19149,N_11093,N_12669);
or U19150 (N_19150,N_10448,N_13462);
nand U19151 (N_19151,N_10400,N_10112);
or U19152 (N_19152,N_10944,N_14033);
nor U19153 (N_19153,N_10003,N_14688);
nor U19154 (N_19154,N_13628,N_11256);
and U19155 (N_19155,N_14920,N_11823);
or U19156 (N_19156,N_11255,N_10642);
nor U19157 (N_19157,N_10674,N_14769);
and U19158 (N_19158,N_13906,N_13339);
or U19159 (N_19159,N_11091,N_11293);
and U19160 (N_19160,N_10493,N_10356);
xor U19161 (N_19161,N_12354,N_11848);
nor U19162 (N_19162,N_12892,N_11609);
xor U19163 (N_19163,N_14021,N_12753);
and U19164 (N_19164,N_11164,N_12377);
and U19165 (N_19165,N_14166,N_12344);
or U19166 (N_19166,N_14959,N_14313);
xnor U19167 (N_19167,N_11147,N_14300);
xnor U19168 (N_19168,N_11582,N_10364);
nand U19169 (N_19169,N_13503,N_12530);
nand U19170 (N_19170,N_14673,N_13382);
or U19171 (N_19171,N_11359,N_10334);
and U19172 (N_19172,N_10064,N_13783);
xor U19173 (N_19173,N_12260,N_14538);
or U19174 (N_19174,N_13854,N_10898);
nand U19175 (N_19175,N_13438,N_11530);
xor U19176 (N_19176,N_11779,N_10811);
nor U19177 (N_19177,N_10292,N_11996);
xnor U19178 (N_19178,N_13510,N_12909);
or U19179 (N_19179,N_11955,N_14375);
nor U19180 (N_19180,N_10658,N_14765);
nor U19181 (N_19181,N_11285,N_14194);
xnor U19182 (N_19182,N_12522,N_13391);
and U19183 (N_19183,N_10507,N_10420);
nor U19184 (N_19184,N_12855,N_13214);
xor U19185 (N_19185,N_13071,N_11103);
xor U19186 (N_19186,N_12035,N_10043);
nor U19187 (N_19187,N_14999,N_12324);
and U19188 (N_19188,N_12034,N_14545);
or U19189 (N_19189,N_14731,N_10604);
nand U19190 (N_19190,N_12865,N_11193);
and U19191 (N_19191,N_10283,N_12267);
or U19192 (N_19192,N_11118,N_13566);
nand U19193 (N_19193,N_13800,N_10899);
or U19194 (N_19194,N_13520,N_14110);
or U19195 (N_19195,N_12004,N_11191);
and U19196 (N_19196,N_13229,N_12962);
xor U19197 (N_19197,N_10839,N_13856);
xnor U19198 (N_19198,N_11484,N_14745);
nand U19199 (N_19199,N_11104,N_11147);
nor U19200 (N_19200,N_13084,N_11521);
nor U19201 (N_19201,N_10813,N_11121);
nand U19202 (N_19202,N_10170,N_12320);
and U19203 (N_19203,N_10370,N_14026);
and U19204 (N_19204,N_10905,N_11410);
and U19205 (N_19205,N_14087,N_13992);
and U19206 (N_19206,N_14861,N_13464);
xor U19207 (N_19207,N_14845,N_14331);
nor U19208 (N_19208,N_11179,N_10389);
xor U19209 (N_19209,N_12404,N_12545);
xor U19210 (N_19210,N_13935,N_10137);
or U19211 (N_19211,N_12841,N_14247);
and U19212 (N_19212,N_10931,N_12426);
or U19213 (N_19213,N_14018,N_12789);
and U19214 (N_19214,N_13894,N_14504);
nor U19215 (N_19215,N_11472,N_12790);
xor U19216 (N_19216,N_13335,N_11358);
and U19217 (N_19217,N_12978,N_13708);
or U19218 (N_19218,N_13874,N_10267);
xor U19219 (N_19219,N_13628,N_10837);
and U19220 (N_19220,N_12196,N_13155);
nand U19221 (N_19221,N_11746,N_13983);
and U19222 (N_19222,N_10963,N_11152);
or U19223 (N_19223,N_14328,N_11381);
xor U19224 (N_19224,N_12208,N_13736);
or U19225 (N_19225,N_14187,N_12897);
nor U19226 (N_19226,N_13570,N_10150);
nor U19227 (N_19227,N_14284,N_11711);
and U19228 (N_19228,N_14413,N_13679);
or U19229 (N_19229,N_10371,N_14520);
or U19230 (N_19230,N_12492,N_12405);
and U19231 (N_19231,N_14051,N_11541);
or U19232 (N_19232,N_10203,N_11049);
nor U19233 (N_19233,N_11671,N_13536);
or U19234 (N_19234,N_14699,N_11896);
and U19235 (N_19235,N_14020,N_14471);
and U19236 (N_19236,N_10120,N_12718);
xnor U19237 (N_19237,N_12651,N_11369);
nand U19238 (N_19238,N_11045,N_12221);
xor U19239 (N_19239,N_14214,N_11505);
nand U19240 (N_19240,N_11994,N_11421);
xnor U19241 (N_19241,N_11391,N_12443);
nand U19242 (N_19242,N_10545,N_11414);
xor U19243 (N_19243,N_12290,N_10536);
nand U19244 (N_19244,N_14229,N_12583);
and U19245 (N_19245,N_14316,N_11243);
xnor U19246 (N_19246,N_11494,N_13331);
and U19247 (N_19247,N_13550,N_13059);
and U19248 (N_19248,N_13613,N_12689);
xor U19249 (N_19249,N_10056,N_13192);
nor U19250 (N_19250,N_10268,N_10175);
or U19251 (N_19251,N_12642,N_14471);
and U19252 (N_19252,N_10043,N_14885);
and U19253 (N_19253,N_11748,N_13004);
xor U19254 (N_19254,N_13171,N_11733);
and U19255 (N_19255,N_11425,N_10852);
nand U19256 (N_19256,N_13887,N_12463);
nand U19257 (N_19257,N_11380,N_12225);
nand U19258 (N_19258,N_12230,N_13952);
or U19259 (N_19259,N_13566,N_11912);
nor U19260 (N_19260,N_10426,N_14347);
or U19261 (N_19261,N_13478,N_13130);
nand U19262 (N_19262,N_13298,N_14931);
and U19263 (N_19263,N_12535,N_13661);
nand U19264 (N_19264,N_12479,N_14754);
nor U19265 (N_19265,N_11731,N_13563);
or U19266 (N_19266,N_10876,N_14997);
and U19267 (N_19267,N_14208,N_11575);
nor U19268 (N_19268,N_13605,N_13227);
or U19269 (N_19269,N_11509,N_12897);
and U19270 (N_19270,N_12026,N_10975);
xor U19271 (N_19271,N_14640,N_13439);
nor U19272 (N_19272,N_10541,N_14578);
nand U19273 (N_19273,N_14333,N_11377);
xor U19274 (N_19274,N_13445,N_11367);
nand U19275 (N_19275,N_10469,N_11944);
and U19276 (N_19276,N_14311,N_12078);
nor U19277 (N_19277,N_13452,N_13546);
xor U19278 (N_19278,N_11380,N_12412);
xnor U19279 (N_19279,N_10718,N_12217);
nand U19280 (N_19280,N_11124,N_12882);
or U19281 (N_19281,N_10970,N_12296);
and U19282 (N_19282,N_12876,N_14842);
nand U19283 (N_19283,N_11611,N_10164);
xor U19284 (N_19284,N_10553,N_12964);
or U19285 (N_19285,N_10946,N_13844);
or U19286 (N_19286,N_11040,N_14450);
and U19287 (N_19287,N_13414,N_11464);
nand U19288 (N_19288,N_11804,N_14153);
nand U19289 (N_19289,N_12507,N_10805);
or U19290 (N_19290,N_11799,N_13890);
nor U19291 (N_19291,N_11137,N_10477);
nand U19292 (N_19292,N_12714,N_10826);
or U19293 (N_19293,N_10548,N_14602);
xor U19294 (N_19294,N_14164,N_12071);
xnor U19295 (N_19295,N_14211,N_13682);
nor U19296 (N_19296,N_13555,N_11605);
xor U19297 (N_19297,N_12827,N_13232);
nand U19298 (N_19298,N_11655,N_10841);
and U19299 (N_19299,N_11033,N_11151);
nor U19300 (N_19300,N_10507,N_10756);
nor U19301 (N_19301,N_11194,N_14911);
xnor U19302 (N_19302,N_11662,N_14318);
or U19303 (N_19303,N_13187,N_12945);
nor U19304 (N_19304,N_11274,N_10005);
nand U19305 (N_19305,N_14373,N_12341);
nor U19306 (N_19306,N_12424,N_12133);
xnor U19307 (N_19307,N_12272,N_14579);
nand U19308 (N_19308,N_13004,N_11386);
nor U19309 (N_19309,N_14331,N_12529);
xor U19310 (N_19310,N_10798,N_10128);
nor U19311 (N_19311,N_14398,N_14074);
or U19312 (N_19312,N_13556,N_12238);
xnor U19313 (N_19313,N_13437,N_12386);
nand U19314 (N_19314,N_11001,N_10106);
xnor U19315 (N_19315,N_11739,N_14836);
xor U19316 (N_19316,N_13139,N_10248);
nor U19317 (N_19317,N_13054,N_14353);
and U19318 (N_19318,N_10072,N_14292);
nor U19319 (N_19319,N_11606,N_13641);
nand U19320 (N_19320,N_10711,N_13840);
and U19321 (N_19321,N_14026,N_12968);
and U19322 (N_19322,N_12746,N_13339);
and U19323 (N_19323,N_10477,N_13893);
or U19324 (N_19324,N_10167,N_13743);
and U19325 (N_19325,N_12820,N_13966);
nor U19326 (N_19326,N_11736,N_14606);
nor U19327 (N_19327,N_11320,N_10834);
nand U19328 (N_19328,N_11367,N_12366);
or U19329 (N_19329,N_12365,N_14091);
nor U19330 (N_19330,N_13978,N_11960);
nor U19331 (N_19331,N_13708,N_11553);
or U19332 (N_19332,N_12767,N_10570);
or U19333 (N_19333,N_13781,N_10867);
and U19334 (N_19334,N_12996,N_13673);
or U19335 (N_19335,N_10438,N_10883);
and U19336 (N_19336,N_10693,N_14901);
nand U19337 (N_19337,N_13649,N_12324);
nand U19338 (N_19338,N_11721,N_11825);
nor U19339 (N_19339,N_11112,N_14971);
or U19340 (N_19340,N_12455,N_11318);
and U19341 (N_19341,N_11097,N_13133);
or U19342 (N_19342,N_11529,N_11078);
nor U19343 (N_19343,N_14667,N_13228);
nand U19344 (N_19344,N_10695,N_14218);
xor U19345 (N_19345,N_12714,N_12826);
and U19346 (N_19346,N_12600,N_13977);
xor U19347 (N_19347,N_14648,N_10405);
or U19348 (N_19348,N_14050,N_11678);
or U19349 (N_19349,N_13218,N_13070);
nor U19350 (N_19350,N_14109,N_12710);
xor U19351 (N_19351,N_13885,N_13212);
nand U19352 (N_19352,N_10400,N_13142);
nand U19353 (N_19353,N_12846,N_11095);
or U19354 (N_19354,N_11657,N_12347);
and U19355 (N_19355,N_12342,N_10955);
nand U19356 (N_19356,N_14913,N_13460);
xnor U19357 (N_19357,N_11073,N_12507);
nor U19358 (N_19358,N_12854,N_14878);
or U19359 (N_19359,N_12214,N_12741);
nor U19360 (N_19360,N_14436,N_11040);
nand U19361 (N_19361,N_10584,N_13098);
nand U19362 (N_19362,N_11028,N_12398);
or U19363 (N_19363,N_11003,N_11058);
nand U19364 (N_19364,N_10614,N_14026);
nand U19365 (N_19365,N_13512,N_11040);
and U19366 (N_19366,N_14118,N_13752);
nand U19367 (N_19367,N_14584,N_12038);
xor U19368 (N_19368,N_12449,N_10222);
nand U19369 (N_19369,N_12309,N_14477);
nand U19370 (N_19370,N_10741,N_11139);
xnor U19371 (N_19371,N_13439,N_10356);
nor U19372 (N_19372,N_11463,N_13740);
and U19373 (N_19373,N_10845,N_10205);
xnor U19374 (N_19374,N_12402,N_11541);
xnor U19375 (N_19375,N_13476,N_14452);
and U19376 (N_19376,N_13318,N_11150);
xnor U19377 (N_19377,N_12066,N_12704);
nand U19378 (N_19378,N_11320,N_14521);
xor U19379 (N_19379,N_10375,N_11008);
or U19380 (N_19380,N_11871,N_12945);
nor U19381 (N_19381,N_12887,N_10539);
and U19382 (N_19382,N_12523,N_13531);
xor U19383 (N_19383,N_11324,N_11627);
and U19384 (N_19384,N_13602,N_11821);
or U19385 (N_19385,N_14466,N_12185);
and U19386 (N_19386,N_10324,N_13532);
nor U19387 (N_19387,N_13730,N_12480);
or U19388 (N_19388,N_12356,N_14794);
nor U19389 (N_19389,N_10890,N_12058);
nand U19390 (N_19390,N_10305,N_11362);
or U19391 (N_19391,N_11282,N_12568);
and U19392 (N_19392,N_10089,N_13166);
xnor U19393 (N_19393,N_12626,N_11278);
and U19394 (N_19394,N_10131,N_13649);
xor U19395 (N_19395,N_12346,N_11305);
nor U19396 (N_19396,N_12235,N_10822);
or U19397 (N_19397,N_10177,N_11738);
or U19398 (N_19398,N_11380,N_11423);
xor U19399 (N_19399,N_14881,N_14233);
and U19400 (N_19400,N_13251,N_14774);
xnor U19401 (N_19401,N_12180,N_14430);
nand U19402 (N_19402,N_12224,N_14889);
and U19403 (N_19403,N_12153,N_11061);
nor U19404 (N_19404,N_14907,N_13526);
nor U19405 (N_19405,N_13921,N_11513);
nand U19406 (N_19406,N_12553,N_11401);
or U19407 (N_19407,N_10221,N_11043);
nand U19408 (N_19408,N_11547,N_13374);
nor U19409 (N_19409,N_12360,N_10756);
or U19410 (N_19410,N_13096,N_13232);
nand U19411 (N_19411,N_12049,N_11769);
and U19412 (N_19412,N_13139,N_11833);
nor U19413 (N_19413,N_14050,N_10592);
nand U19414 (N_19414,N_13274,N_11137);
xnor U19415 (N_19415,N_12643,N_11699);
nand U19416 (N_19416,N_13700,N_14693);
or U19417 (N_19417,N_12213,N_10485);
nand U19418 (N_19418,N_10587,N_11319);
nor U19419 (N_19419,N_10582,N_12817);
nand U19420 (N_19420,N_10355,N_13016);
nor U19421 (N_19421,N_11906,N_13739);
nor U19422 (N_19422,N_11683,N_11287);
xor U19423 (N_19423,N_11729,N_13902);
nand U19424 (N_19424,N_11563,N_13957);
nor U19425 (N_19425,N_13023,N_13786);
xor U19426 (N_19426,N_10050,N_14041);
or U19427 (N_19427,N_13108,N_14905);
xnor U19428 (N_19428,N_14473,N_12713);
nor U19429 (N_19429,N_14354,N_12270);
nor U19430 (N_19430,N_11932,N_12385);
or U19431 (N_19431,N_13488,N_14963);
xor U19432 (N_19432,N_12953,N_14733);
xor U19433 (N_19433,N_14917,N_10591);
xnor U19434 (N_19434,N_12354,N_10727);
xnor U19435 (N_19435,N_11216,N_11335);
nor U19436 (N_19436,N_13045,N_14520);
xnor U19437 (N_19437,N_14111,N_10160);
nor U19438 (N_19438,N_10688,N_12151);
and U19439 (N_19439,N_13868,N_12438);
and U19440 (N_19440,N_12936,N_14513);
nor U19441 (N_19441,N_14409,N_11138);
or U19442 (N_19442,N_14289,N_11675);
nor U19443 (N_19443,N_10070,N_12352);
or U19444 (N_19444,N_14704,N_11417);
and U19445 (N_19445,N_10026,N_13885);
nand U19446 (N_19446,N_11846,N_11563);
xor U19447 (N_19447,N_13110,N_10637);
xnor U19448 (N_19448,N_12319,N_14760);
nand U19449 (N_19449,N_12943,N_14040);
nor U19450 (N_19450,N_13885,N_12778);
or U19451 (N_19451,N_14218,N_13307);
xnor U19452 (N_19452,N_11873,N_14960);
and U19453 (N_19453,N_14483,N_13961);
nand U19454 (N_19454,N_10118,N_12423);
nand U19455 (N_19455,N_10652,N_14056);
and U19456 (N_19456,N_11893,N_14185);
or U19457 (N_19457,N_11193,N_11400);
or U19458 (N_19458,N_10153,N_11234);
xnor U19459 (N_19459,N_10797,N_10453);
nand U19460 (N_19460,N_12714,N_14067);
or U19461 (N_19461,N_14680,N_13167);
xor U19462 (N_19462,N_14065,N_10662);
nand U19463 (N_19463,N_11680,N_10128);
or U19464 (N_19464,N_11135,N_11833);
or U19465 (N_19465,N_10456,N_13942);
and U19466 (N_19466,N_13380,N_13752);
or U19467 (N_19467,N_10892,N_10810);
nand U19468 (N_19468,N_12255,N_12829);
or U19469 (N_19469,N_10617,N_11163);
or U19470 (N_19470,N_13577,N_12646);
or U19471 (N_19471,N_14232,N_10582);
or U19472 (N_19472,N_12511,N_10230);
nand U19473 (N_19473,N_10904,N_12331);
and U19474 (N_19474,N_10364,N_12611);
and U19475 (N_19475,N_13017,N_13790);
nor U19476 (N_19476,N_11872,N_14954);
nand U19477 (N_19477,N_10066,N_13089);
xor U19478 (N_19478,N_14290,N_10696);
xnor U19479 (N_19479,N_12251,N_12236);
nor U19480 (N_19480,N_12440,N_11088);
xor U19481 (N_19481,N_14562,N_10044);
and U19482 (N_19482,N_10905,N_13837);
nand U19483 (N_19483,N_13909,N_11726);
or U19484 (N_19484,N_13841,N_13681);
nor U19485 (N_19485,N_11339,N_12392);
nand U19486 (N_19486,N_14920,N_13383);
nand U19487 (N_19487,N_13248,N_13674);
xnor U19488 (N_19488,N_11364,N_11416);
and U19489 (N_19489,N_10701,N_12006);
xnor U19490 (N_19490,N_14437,N_11920);
xor U19491 (N_19491,N_13365,N_11804);
nand U19492 (N_19492,N_10991,N_11686);
or U19493 (N_19493,N_10934,N_11370);
or U19494 (N_19494,N_12385,N_14840);
or U19495 (N_19495,N_11684,N_10568);
and U19496 (N_19496,N_11530,N_11338);
nand U19497 (N_19497,N_14027,N_12656);
xnor U19498 (N_19498,N_12651,N_10935);
and U19499 (N_19499,N_11636,N_14263);
xnor U19500 (N_19500,N_14131,N_11912);
nand U19501 (N_19501,N_12937,N_13098);
and U19502 (N_19502,N_10118,N_11389);
xor U19503 (N_19503,N_13438,N_10256);
xor U19504 (N_19504,N_12513,N_13321);
xor U19505 (N_19505,N_12139,N_10243);
and U19506 (N_19506,N_12756,N_12680);
and U19507 (N_19507,N_10599,N_10798);
nor U19508 (N_19508,N_10467,N_11447);
xnor U19509 (N_19509,N_12587,N_13878);
and U19510 (N_19510,N_14711,N_13384);
nor U19511 (N_19511,N_14974,N_14427);
nand U19512 (N_19512,N_11705,N_14360);
or U19513 (N_19513,N_14892,N_12801);
nand U19514 (N_19514,N_13998,N_13692);
nor U19515 (N_19515,N_14927,N_14130);
nor U19516 (N_19516,N_14734,N_10168);
xor U19517 (N_19517,N_11994,N_10339);
and U19518 (N_19518,N_14306,N_11592);
or U19519 (N_19519,N_12906,N_13124);
nor U19520 (N_19520,N_14715,N_13411);
nor U19521 (N_19521,N_11119,N_10452);
nand U19522 (N_19522,N_13362,N_13589);
and U19523 (N_19523,N_14469,N_10844);
or U19524 (N_19524,N_12974,N_13259);
xor U19525 (N_19525,N_11154,N_13714);
nand U19526 (N_19526,N_12211,N_14594);
nor U19527 (N_19527,N_10937,N_12092);
or U19528 (N_19528,N_12274,N_14571);
or U19529 (N_19529,N_10567,N_14511);
nand U19530 (N_19530,N_10709,N_12244);
and U19531 (N_19531,N_10712,N_11172);
nor U19532 (N_19532,N_13155,N_13372);
or U19533 (N_19533,N_13768,N_13952);
nand U19534 (N_19534,N_13459,N_11368);
and U19535 (N_19535,N_11806,N_11825);
xnor U19536 (N_19536,N_11351,N_11405);
nor U19537 (N_19537,N_14296,N_10210);
xnor U19538 (N_19538,N_10923,N_14364);
xor U19539 (N_19539,N_13197,N_13521);
or U19540 (N_19540,N_14899,N_10722);
or U19541 (N_19541,N_10189,N_14960);
xnor U19542 (N_19542,N_13950,N_10392);
nor U19543 (N_19543,N_11705,N_11114);
or U19544 (N_19544,N_14051,N_13653);
and U19545 (N_19545,N_14425,N_14932);
or U19546 (N_19546,N_12632,N_10087);
nor U19547 (N_19547,N_11557,N_12376);
or U19548 (N_19548,N_14510,N_11846);
nor U19549 (N_19549,N_13411,N_11427);
and U19550 (N_19550,N_11597,N_12813);
nor U19551 (N_19551,N_14549,N_14411);
xor U19552 (N_19552,N_10547,N_12056);
nand U19553 (N_19553,N_12142,N_12498);
nor U19554 (N_19554,N_13066,N_10480);
and U19555 (N_19555,N_13664,N_10607);
or U19556 (N_19556,N_10755,N_14401);
nor U19557 (N_19557,N_12841,N_10032);
xnor U19558 (N_19558,N_14693,N_13563);
or U19559 (N_19559,N_11046,N_10621);
and U19560 (N_19560,N_10793,N_11644);
or U19561 (N_19561,N_10137,N_14264);
and U19562 (N_19562,N_12753,N_14458);
nand U19563 (N_19563,N_14753,N_14928);
or U19564 (N_19564,N_10019,N_14774);
or U19565 (N_19565,N_10669,N_11648);
nand U19566 (N_19566,N_14337,N_10024);
nor U19567 (N_19567,N_14544,N_11185);
or U19568 (N_19568,N_12710,N_10674);
and U19569 (N_19569,N_10745,N_14502);
nand U19570 (N_19570,N_14696,N_10319);
or U19571 (N_19571,N_14086,N_10499);
or U19572 (N_19572,N_13004,N_10768);
nor U19573 (N_19573,N_14196,N_11863);
or U19574 (N_19574,N_12921,N_10866);
nor U19575 (N_19575,N_10426,N_11302);
and U19576 (N_19576,N_10524,N_12108);
and U19577 (N_19577,N_13806,N_10117);
and U19578 (N_19578,N_11271,N_11382);
or U19579 (N_19579,N_10007,N_14316);
or U19580 (N_19580,N_13095,N_11399);
xnor U19581 (N_19581,N_11222,N_12585);
nor U19582 (N_19582,N_14252,N_12761);
or U19583 (N_19583,N_11890,N_14942);
xnor U19584 (N_19584,N_11686,N_13462);
and U19585 (N_19585,N_14428,N_13392);
nor U19586 (N_19586,N_13568,N_13552);
nor U19587 (N_19587,N_13724,N_14204);
and U19588 (N_19588,N_10635,N_13537);
nor U19589 (N_19589,N_12563,N_13542);
xnor U19590 (N_19590,N_13187,N_14693);
xnor U19591 (N_19591,N_11217,N_13292);
or U19592 (N_19592,N_10437,N_13244);
or U19593 (N_19593,N_11421,N_14775);
xnor U19594 (N_19594,N_11127,N_13511);
and U19595 (N_19595,N_13610,N_14298);
nor U19596 (N_19596,N_10341,N_13063);
nand U19597 (N_19597,N_12762,N_14893);
nand U19598 (N_19598,N_11480,N_13324);
nor U19599 (N_19599,N_11741,N_13530);
nor U19600 (N_19600,N_13170,N_12004);
or U19601 (N_19601,N_12291,N_10355);
nor U19602 (N_19602,N_10055,N_13025);
nor U19603 (N_19603,N_11037,N_12344);
or U19604 (N_19604,N_10570,N_12988);
or U19605 (N_19605,N_11340,N_10221);
nand U19606 (N_19606,N_14325,N_10659);
nor U19607 (N_19607,N_10335,N_13583);
and U19608 (N_19608,N_12846,N_10014);
xor U19609 (N_19609,N_11054,N_12249);
nand U19610 (N_19610,N_13423,N_10947);
and U19611 (N_19611,N_11656,N_14921);
nand U19612 (N_19612,N_10277,N_10128);
nand U19613 (N_19613,N_12678,N_12923);
and U19614 (N_19614,N_12472,N_10365);
or U19615 (N_19615,N_11176,N_13464);
and U19616 (N_19616,N_12202,N_12763);
or U19617 (N_19617,N_11926,N_11630);
or U19618 (N_19618,N_14492,N_10504);
or U19619 (N_19619,N_12430,N_11267);
nor U19620 (N_19620,N_10209,N_13220);
or U19621 (N_19621,N_12544,N_10990);
xor U19622 (N_19622,N_11323,N_11001);
nand U19623 (N_19623,N_14779,N_11333);
or U19624 (N_19624,N_10669,N_10331);
nand U19625 (N_19625,N_10193,N_11723);
xnor U19626 (N_19626,N_12230,N_13978);
and U19627 (N_19627,N_10938,N_11138);
or U19628 (N_19628,N_12960,N_12373);
nor U19629 (N_19629,N_13606,N_12431);
or U19630 (N_19630,N_13871,N_12580);
xnor U19631 (N_19631,N_11099,N_10504);
nor U19632 (N_19632,N_10071,N_13248);
xor U19633 (N_19633,N_10762,N_14106);
xor U19634 (N_19634,N_13102,N_13426);
and U19635 (N_19635,N_12895,N_13091);
and U19636 (N_19636,N_10264,N_10830);
nand U19637 (N_19637,N_13021,N_14924);
nor U19638 (N_19638,N_10880,N_12360);
nand U19639 (N_19639,N_14656,N_10152);
nor U19640 (N_19640,N_11046,N_10753);
nand U19641 (N_19641,N_12461,N_13831);
nor U19642 (N_19642,N_14492,N_10955);
and U19643 (N_19643,N_12071,N_11696);
and U19644 (N_19644,N_13292,N_13519);
and U19645 (N_19645,N_11762,N_14624);
nor U19646 (N_19646,N_10839,N_12170);
and U19647 (N_19647,N_14918,N_10811);
xnor U19648 (N_19648,N_13901,N_11269);
nor U19649 (N_19649,N_14006,N_13785);
or U19650 (N_19650,N_11458,N_10063);
nand U19651 (N_19651,N_12190,N_12846);
nand U19652 (N_19652,N_11297,N_12071);
and U19653 (N_19653,N_12034,N_10778);
nor U19654 (N_19654,N_11990,N_11904);
nand U19655 (N_19655,N_12898,N_13986);
nand U19656 (N_19656,N_13608,N_13232);
xnor U19657 (N_19657,N_13144,N_13009);
xor U19658 (N_19658,N_14666,N_11146);
xnor U19659 (N_19659,N_12661,N_12551);
xnor U19660 (N_19660,N_11873,N_10266);
or U19661 (N_19661,N_10392,N_12857);
and U19662 (N_19662,N_12321,N_14779);
and U19663 (N_19663,N_12021,N_14305);
or U19664 (N_19664,N_13478,N_10632);
nand U19665 (N_19665,N_14121,N_10675);
nand U19666 (N_19666,N_13681,N_12640);
nand U19667 (N_19667,N_13267,N_13138);
nand U19668 (N_19668,N_13062,N_10955);
nand U19669 (N_19669,N_13250,N_10760);
and U19670 (N_19670,N_14815,N_12706);
and U19671 (N_19671,N_11076,N_11697);
and U19672 (N_19672,N_14922,N_14871);
nor U19673 (N_19673,N_10384,N_11493);
nor U19674 (N_19674,N_12246,N_10055);
and U19675 (N_19675,N_10301,N_11909);
xor U19676 (N_19676,N_13302,N_10370);
xor U19677 (N_19677,N_13719,N_13581);
and U19678 (N_19678,N_13604,N_10148);
nor U19679 (N_19679,N_11438,N_13158);
nor U19680 (N_19680,N_11299,N_14891);
nor U19681 (N_19681,N_10898,N_11730);
or U19682 (N_19682,N_13763,N_12483);
xor U19683 (N_19683,N_14451,N_11850);
nor U19684 (N_19684,N_11282,N_14504);
or U19685 (N_19685,N_10821,N_11739);
xor U19686 (N_19686,N_10491,N_10803);
or U19687 (N_19687,N_13550,N_14499);
and U19688 (N_19688,N_14922,N_13036);
nor U19689 (N_19689,N_10830,N_14377);
and U19690 (N_19690,N_10608,N_11692);
and U19691 (N_19691,N_10656,N_14612);
or U19692 (N_19692,N_13981,N_11985);
and U19693 (N_19693,N_11691,N_13554);
xor U19694 (N_19694,N_13829,N_13447);
or U19695 (N_19695,N_13828,N_14293);
xor U19696 (N_19696,N_11129,N_11374);
xor U19697 (N_19697,N_11116,N_14358);
xnor U19698 (N_19698,N_14236,N_10973);
nand U19699 (N_19699,N_12326,N_11224);
or U19700 (N_19700,N_13519,N_13732);
nand U19701 (N_19701,N_11770,N_11360);
nand U19702 (N_19702,N_11174,N_11761);
nor U19703 (N_19703,N_10747,N_12513);
or U19704 (N_19704,N_10849,N_11252);
nand U19705 (N_19705,N_13290,N_11813);
nor U19706 (N_19706,N_11948,N_13252);
xnor U19707 (N_19707,N_14802,N_13471);
xor U19708 (N_19708,N_10758,N_10890);
nor U19709 (N_19709,N_12098,N_13384);
nor U19710 (N_19710,N_10450,N_11103);
or U19711 (N_19711,N_13188,N_10037);
nand U19712 (N_19712,N_14692,N_14281);
nand U19713 (N_19713,N_12671,N_14167);
nor U19714 (N_19714,N_10177,N_12618);
or U19715 (N_19715,N_10056,N_14962);
and U19716 (N_19716,N_13816,N_14509);
or U19717 (N_19717,N_13675,N_10563);
and U19718 (N_19718,N_12359,N_12030);
and U19719 (N_19719,N_14878,N_10792);
and U19720 (N_19720,N_10291,N_11668);
or U19721 (N_19721,N_12980,N_10104);
nor U19722 (N_19722,N_11228,N_11716);
and U19723 (N_19723,N_11534,N_13661);
xor U19724 (N_19724,N_14949,N_13465);
or U19725 (N_19725,N_10154,N_10001);
nand U19726 (N_19726,N_13073,N_13118);
or U19727 (N_19727,N_10113,N_13138);
nor U19728 (N_19728,N_11757,N_14664);
xor U19729 (N_19729,N_11700,N_12709);
xor U19730 (N_19730,N_11931,N_12094);
and U19731 (N_19731,N_14089,N_13255);
and U19732 (N_19732,N_11144,N_10986);
and U19733 (N_19733,N_10813,N_10534);
nand U19734 (N_19734,N_14325,N_10776);
xnor U19735 (N_19735,N_14525,N_10483);
nor U19736 (N_19736,N_14463,N_10988);
nor U19737 (N_19737,N_12460,N_14458);
xnor U19738 (N_19738,N_14444,N_12766);
and U19739 (N_19739,N_11013,N_13128);
nor U19740 (N_19740,N_10568,N_14660);
or U19741 (N_19741,N_12263,N_13789);
nor U19742 (N_19742,N_14621,N_12225);
nor U19743 (N_19743,N_11211,N_13168);
or U19744 (N_19744,N_14642,N_13829);
xor U19745 (N_19745,N_12620,N_13204);
and U19746 (N_19746,N_12142,N_10331);
and U19747 (N_19747,N_13440,N_12283);
nor U19748 (N_19748,N_10422,N_11690);
and U19749 (N_19749,N_11240,N_11085);
or U19750 (N_19750,N_14039,N_14133);
or U19751 (N_19751,N_14347,N_10258);
or U19752 (N_19752,N_10884,N_14035);
or U19753 (N_19753,N_10504,N_12289);
nor U19754 (N_19754,N_13432,N_12153);
nand U19755 (N_19755,N_10550,N_10086);
and U19756 (N_19756,N_14543,N_11842);
nand U19757 (N_19757,N_13032,N_13397);
xnor U19758 (N_19758,N_11317,N_12903);
nor U19759 (N_19759,N_14458,N_12656);
or U19760 (N_19760,N_10562,N_14448);
or U19761 (N_19761,N_11869,N_14928);
xnor U19762 (N_19762,N_14910,N_13451);
and U19763 (N_19763,N_14941,N_12955);
xnor U19764 (N_19764,N_13188,N_14215);
and U19765 (N_19765,N_11890,N_11892);
or U19766 (N_19766,N_11612,N_10152);
nor U19767 (N_19767,N_14955,N_13095);
nor U19768 (N_19768,N_12255,N_10865);
xor U19769 (N_19769,N_11218,N_10375);
nor U19770 (N_19770,N_14851,N_11584);
nor U19771 (N_19771,N_10352,N_13774);
xor U19772 (N_19772,N_10473,N_10469);
xor U19773 (N_19773,N_14418,N_14777);
nor U19774 (N_19774,N_13289,N_14028);
nor U19775 (N_19775,N_13804,N_10160);
or U19776 (N_19776,N_10482,N_13296);
or U19777 (N_19777,N_13589,N_14126);
nand U19778 (N_19778,N_11585,N_12332);
nor U19779 (N_19779,N_10583,N_14607);
and U19780 (N_19780,N_12662,N_10186);
xnor U19781 (N_19781,N_14260,N_13895);
nand U19782 (N_19782,N_10325,N_14312);
nand U19783 (N_19783,N_10497,N_14849);
and U19784 (N_19784,N_10500,N_13051);
nor U19785 (N_19785,N_13451,N_11005);
xor U19786 (N_19786,N_12924,N_12329);
and U19787 (N_19787,N_11735,N_13762);
nor U19788 (N_19788,N_11053,N_13286);
nor U19789 (N_19789,N_11095,N_10793);
nor U19790 (N_19790,N_10861,N_11875);
or U19791 (N_19791,N_13932,N_13285);
or U19792 (N_19792,N_12420,N_14441);
nand U19793 (N_19793,N_11743,N_14703);
nor U19794 (N_19794,N_10456,N_10428);
nand U19795 (N_19795,N_11899,N_10409);
nand U19796 (N_19796,N_12852,N_14542);
or U19797 (N_19797,N_10952,N_13200);
or U19798 (N_19798,N_12347,N_10661);
nand U19799 (N_19799,N_10297,N_10433);
or U19800 (N_19800,N_13067,N_12976);
nand U19801 (N_19801,N_10842,N_10262);
or U19802 (N_19802,N_14892,N_14539);
nand U19803 (N_19803,N_12870,N_13068);
and U19804 (N_19804,N_13903,N_13722);
nor U19805 (N_19805,N_14203,N_13522);
or U19806 (N_19806,N_10404,N_13447);
nand U19807 (N_19807,N_10967,N_14531);
or U19808 (N_19808,N_10086,N_10611);
nand U19809 (N_19809,N_12669,N_13262);
nor U19810 (N_19810,N_13849,N_10823);
nor U19811 (N_19811,N_10380,N_13195);
nor U19812 (N_19812,N_14357,N_14481);
or U19813 (N_19813,N_12699,N_11482);
nor U19814 (N_19814,N_10364,N_14839);
or U19815 (N_19815,N_10726,N_14236);
and U19816 (N_19816,N_13141,N_13337);
nor U19817 (N_19817,N_13593,N_11626);
and U19818 (N_19818,N_12652,N_12064);
and U19819 (N_19819,N_12323,N_11793);
xor U19820 (N_19820,N_14102,N_10499);
and U19821 (N_19821,N_11026,N_13227);
nand U19822 (N_19822,N_10608,N_14164);
nor U19823 (N_19823,N_12494,N_13046);
and U19824 (N_19824,N_14999,N_11813);
xor U19825 (N_19825,N_10748,N_11364);
nor U19826 (N_19826,N_10349,N_13995);
xnor U19827 (N_19827,N_11004,N_14218);
or U19828 (N_19828,N_13581,N_13686);
and U19829 (N_19829,N_13104,N_11766);
and U19830 (N_19830,N_12711,N_10610);
nand U19831 (N_19831,N_14640,N_14502);
xnor U19832 (N_19832,N_13297,N_14092);
nor U19833 (N_19833,N_14168,N_11490);
or U19834 (N_19834,N_14228,N_10455);
or U19835 (N_19835,N_11200,N_14386);
or U19836 (N_19836,N_14053,N_13069);
or U19837 (N_19837,N_10964,N_11481);
and U19838 (N_19838,N_12806,N_11930);
and U19839 (N_19839,N_13899,N_13478);
xor U19840 (N_19840,N_13724,N_10570);
nor U19841 (N_19841,N_14588,N_13798);
xnor U19842 (N_19842,N_10286,N_11942);
or U19843 (N_19843,N_10397,N_10923);
nor U19844 (N_19844,N_14218,N_10114);
and U19845 (N_19845,N_11291,N_11523);
or U19846 (N_19846,N_11065,N_12031);
nor U19847 (N_19847,N_12696,N_14311);
or U19848 (N_19848,N_14506,N_14043);
nor U19849 (N_19849,N_10604,N_10643);
or U19850 (N_19850,N_11097,N_14548);
xor U19851 (N_19851,N_10852,N_10592);
nand U19852 (N_19852,N_14519,N_12018);
and U19853 (N_19853,N_10773,N_12862);
nand U19854 (N_19854,N_13300,N_13734);
and U19855 (N_19855,N_13585,N_13358);
nand U19856 (N_19856,N_12359,N_12634);
nand U19857 (N_19857,N_11927,N_13862);
or U19858 (N_19858,N_14650,N_13133);
xor U19859 (N_19859,N_11670,N_13207);
or U19860 (N_19860,N_11513,N_13640);
and U19861 (N_19861,N_10110,N_11306);
and U19862 (N_19862,N_14000,N_10243);
and U19863 (N_19863,N_13849,N_13181);
or U19864 (N_19864,N_10107,N_11174);
xnor U19865 (N_19865,N_11610,N_11618);
and U19866 (N_19866,N_11483,N_13397);
xor U19867 (N_19867,N_12873,N_12285);
and U19868 (N_19868,N_11098,N_12756);
or U19869 (N_19869,N_11152,N_13831);
or U19870 (N_19870,N_10586,N_14063);
nand U19871 (N_19871,N_14060,N_10998);
nor U19872 (N_19872,N_11289,N_14975);
nand U19873 (N_19873,N_10456,N_12262);
nor U19874 (N_19874,N_10897,N_10644);
xor U19875 (N_19875,N_14321,N_10726);
and U19876 (N_19876,N_11832,N_13763);
or U19877 (N_19877,N_12220,N_13954);
xor U19878 (N_19878,N_12155,N_13578);
xnor U19879 (N_19879,N_10058,N_10348);
and U19880 (N_19880,N_14968,N_13180);
nand U19881 (N_19881,N_11209,N_12020);
or U19882 (N_19882,N_12943,N_12409);
xor U19883 (N_19883,N_10746,N_14117);
and U19884 (N_19884,N_10824,N_12768);
nand U19885 (N_19885,N_14720,N_14837);
nand U19886 (N_19886,N_14111,N_11930);
nor U19887 (N_19887,N_11531,N_11950);
xnor U19888 (N_19888,N_12748,N_13811);
nor U19889 (N_19889,N_13172,N_11514);
xnor U19890 (N_19890,N_11093,N_12651);
and U19891 (N_19891,N_11941,N_13438);
nand U19892 (N_19892,N_14282,N_13448);
nand U19893 (N_19893,N_11666,N_10352);
or U19894 (N_19894,N_10403,N_13477);
and U19895 (N_19895,N_12344,N_13351);
nand U19896 (N_19896,N_13158,N_13131);
and U19897 (N_19897,N_10165,N_12989);
xor U19898 (N_19898,N_13029,N_11358);
nand U19899 (N_19899,N_11703,N_11212);
and U19900 (N_19900,N_14681,N_13826);
xnor U19901 (N_19901,N_11058,N_14927);
and U19902 (N_19902,N_12755,N_14239);
or U19903 (N_19903,N_11263,N_10696);
nor U19904 (N_19904,N_11280,N_12149);
or U19905 (N_19905,N_11473,N_11588);
and U19906 (N_19906,N_13081,N_13819);
nand U19907 (N_19907,N_13301,N_10506);
xor U19908 (N_19908,N_12447,N_11429);
xor U19909 (N_19909,N_12632,N_14543);
and U19910 (N_19910,N_13004,N_10846);
xor U19911 (N_19911,N_13877,N_14335);
xnor U19912 (N_19912,N_11968,N_13999);
or U19913 (N_19913,N_10390,N_13268);
nor U19914 (N_19914,N_10456,N_13650);
and U19915 (N_19915,N_13890,N_12953);
xor U19916 (N_19916,N_14687,N_10941);
and U19917 (N_19917,N_13358,N_13937);
xnor U19918 (N_19918,N_11858,N_13723);
nand U19919 (N_19919,N_14819,N_11749);
xor U19920 (N_19920,N_10478,N_12094);
or U19921 (N_19921,N_11793,N_10985);
and U19922 (N_19922,N_13669,N_11263);
nor U19923 (N_19923,N_13941,N_13912);
and U19924 (N_19924,N_12245,N_14218);
and U19925 (N_19925,N_11447,N_14167);
nor U19926 (N_19926,N_13526,N_13319);
nor U19927 (N_19927,N_14145,N_11962);
nand U19928 (N_19928,N_14145,N_13667);
xnor U19929 (N_19929,N_11199,N_12285);
nand U19930 (N_19930,N_14438,N_11742);
xor U19931 (N_19931,N_10037,N_11311);
nor U19932 (N_19932,N_14932,N_13740);
nor U19933 (N_19933,N_14763,N_12443);
nand U19934 (N_19934,N_10136,N_11645);
or U19935 (N_19935,N_14453,N_14400);
and U19936 (N_19936,N_11901,N_13666);
xor U19937 (N_19937,N_11808,N_12794);
nor U19938 (N_19938,N_10691,N_13858);
and U19939 (N_19939,N_11217,N_10240);
xnor U19940 (N_19940,N_14174,N_13274);
nor U19941 (N_19941,N_11325,N_13525);
xor U19942 (N_19942,N_11290,N_11276);
and U19943 (N_19943,N_13603,N_12389);
and U19944 (N_19944,N_14928,N_13275);
nand U19945 (N_19945,N_11762,N_10659);
or U19946 (N_19946,N_11652,N_12658);
nand U19947 (N_19947,N_12075,N_13342);
nand U19948 (N_19948,N_13755,N_13089);
nand U19949 (N_19949,N_14047,N_11733);
and U19950 (N_19950,N_13375,N_14359);
xor U19951 (N_19951,N_12392,N_10243);
and U19952 (N_19952,N_14315,N_11600);
and U19953 (N_19953,N_13576,N_13276);
nand U19954 (N_19954,N_10813,N_14560);
nand U19955 (N_19955,N_14675,N_12307);
or U19956 (N_19956,N_13760,N_14711);
or U19957 (N_19957,N_10929,N_14381);
or U19958 (N_19958,N_11990,N_10296);
nand U19959 (N_19959,N_12576,N_10927);
nand U19960 (N_19960,N_10293,N_10885);
nor U19961 (N_19961,N_14250,N_10642);
xor U19962 (N_19962,N_10326,N_12183);
xnor U19963 (N_19963,N_13394,N_12938);
or U19964 (N_19964,N_10223,N_13230);
nand U19965 (N_19965,N_11890,N_13003);
nand U19966 (N_19966,N_10718,N_14033);
or U19967 (N_19967,N_12443,N_13587);
and U19968 (N_19968,N_10613,N_14756);
xor U19969 (N_19969,N_13445,N_11033);
or U19970 (N_19970,N_12599,N_10643);
xnor U19971 (N_19971,N_12325,N_14535);
nor U19972 (N_19972,N_12138,N_14136);
nor U19973 (N_19973,N_13323,N_10420);
or U19974 (N_19974,N_14385,N_11150);
or U19975 (N_19975,N_14772,N_12265);
xor U19976 (N_19976,N_13503,N_13398);
and U19977 (N_19977,N_10215,N_12244);
xnor U19978 (N_19978,N_11228,N_11471);
and U19979 (N_19979,N_11394,N_12842);
and U19980 (N_19980,N_13850,N_12101);
and U19981 (N_19981,N_12666,N_13232);
and U19982 (N_19982,N_11870,N_12576);
nand U19983 (N_19983,N_11889,N_14299);
and U19984 (N_19984,N_13288,N_14214);
nand U19985 (N_19985,N_11688,N_13034);
or U19986 (N_19986,N_10977,N_13403);
xnor U19987 (N_19987,N_14117,N_13219);
nor U19988 (N_19988,N_14481,N_13358);
and U19989 (N_19989,N_12152,N_12904);
or U19990 (N_19990,N_14388,N_14043);
and U19991 (N_19991,N_10505,N_13020);
and U19992 (N_19992,N_14601,N_14754);
nor U19993 (N_19993,N_10448,N_12840);
and U19994 (N_19994,N_11413,N_11960);
nand U19995 (N_19995,N_13065,N_10801);
or U19996 (N_19996,N_10460,N_12382);
or U19997 (N_19997,N_14553,N_14023);
nor U19998 (N_19998,N_10930,N_13363);
or U19999 (N_19999,N_10281,N_13123);
and UO_0 (O_0,N_16910,N_19085);
and UO_1 (O_1,N_16423,N_17165);
nor UO_2 (O_2,N_19502,N_16242);
and UO_3 (O_3,N_15805,N_17964);
xor UO_4 (O_4,N_18926,N_16376);
nor UO_5 (O_5,N_15650,N_15905);
and UO_6 (O_6,N_18797,N_19733);
and UO_7 (O_7,N_18612,N_15318);
nor UO_8 (O_8,N_17267,N_15064);
or UO_9 (O_9,N_15604,N_17934);
or UO_10 (O_10,N_18683,N_19542);
xor UO_11 (O_11,N_17240,N_17461);
xor UO_12 (O_12,N_18234,N_15871);
nor UO_13 (O_13,N_15101,N_17684);
or UO_14 (O_14,N_18897,N_17062);
or UO_15 (O_15,N_15019,N_16264);
or UO_16 (O_16,N_19462,N_17086);
nor UO_17 (O_17,N_15723,N_16571);
and UO_18 (O_18,N_19411,N_17121);
nor UO_19 (O_19,N_17638,N_17604);
nand UO_20 (O_20,N_16879,N_16535);
xnor UO_21 (O_21,N_19440,N_19267);
xor UO_22 (O_22,N_16666,N_16846);
xor UO_23 (O_23,N_15610,N_16247);
or UO_24 (O_24,N_18125,N_15726);
xor UO_25 (O_25,N_15363,N_18957);
xor UO_26 (O_26,N_16709,N_19949);
or UO_27 (O_27,N_19753,N_17988);
nand UO_28 (O_28,N_16133,N_18698);
and UO_29 (O_29,N_16634,N_18143);
or UO_30 (O_30,N_19985,N_19190);
or UO_31 (O_31,N_17677,N_17715);
or UO_32 (O_32,N_19548,N_15455);
nor UO_33 (O_33,N_16266,N_15502);
nor UO_34 (O_34,N_18667,N_18755);
and UO_35 (O_35,N_15342,N_19645);
or UO_36 (O_36,N_18166,N_19869);
xor UO_37 (O_37,N_18813,N_15985);
nand UO_38 (O_38,N_16620,N_19025);
nand UO_39 (O_39,N_18986,N_19602);
nand UO_40 (O_40,N_16805,N_19461);
nand UO_41 (O_41,N_19931,N_19076);
nand UO_42 (O_42,N_17469,N_18705);
xnor UO_43 (O_43,N_18261,N_17324);
nand UO_44 (O_44,N_16861,N_16842);
and UO_45 (O_45,N_18331,N_19957);
or UO_46 (O_46,N_18588,N_16436);
nor UO_47 (O_47,N_16733,N_16308);
nor UO_48 (O_48,N_17361,N_19684);
and UO_49 (O_49,N_19594,N_19620);
and UO_50 (O_50,N_19766,N_19323);
or UO_51 (O_51,N_18914,N_15808);
nand UO_52 (O_52,N_19705,N_17236);
or UO_53 (O_53,N_17411,N_19675);
xnor UO_54 (O_54,N_18183,N_15850);
nand UO_55 (O_55,N_18735,N_17234);
nand UO_56 (O_56,N_19337,N_18927);
or UO_57 (O_57,N_17380,N_19146);
nor UO_58 (O_58,N_16375,N_16475);
nand UO_59 (O_59,N_17562,N_17465);
or UO_60 (O_60,N_15111,N_15922);
nand UO_61 (O_61,N_15216,N_17076);
or UO_62 (O_62,N_17342,N_19976);
nor UO_63 (O_63,N_16031,N_19748);
xor UO_64 (O_64,N_18244,N_19689);
or UO_65 (O_65,N_18589,N_17610);
and UO_66 (O_66,N_18966,N_18117);
xor UO_67 (O_67,N_16501,N_19954);
nand UO_68 (O_68,N_17967,N_17237);
nand UO_69 (O_69,N_18992,N_17285);
or UO_70 (O_70,N_18163,N_19149);
nand UO_71 (O_71,N_19824,N_19324);
xnor UO_72 (O_72,N_18587,N_19372);
nand UO_73 (O_73,N_16131,N_17831);
xor UO_74 (O_74,N_19909,N_18446);
nor UO_75 (O_75,N_19830,N_17835);
or UO_76 (O_76,N_17453,N_16896);
or UO_77 (O_77,N_18723,N_18322);
and UO_78 (O_78,N_18795,N_19807);
nor UO_79 (O_79,N_16224,N_17245);
or UO_80 (O_80,N_17116,N_16276);
xnor UO_81 (O_81,N_16100,N_19095);
nor UO_82 (O_82,N_19662,N_19368);
nand UO_83 (O_83,N_19427,N_18655);
nand UO_84 (O_84,N_19537,N_19104);
and UO_85 (O_85,N_19589,N_19086);
nand UO_86 (O_86,N_16459,N_15740);
nand UO_87 (O_87,N_18389,N_19993);
and UO_88 (O_88,N_19357,N_18790);
xnor UO_89 (O_89,N_18057,N_17363);
and UO_90 (O_90,N_17806,N_16366);
nor UO_91 (O_91,N_15947,N_17707);
nand UO_92 (O_92,N_15538,N_18732);
nand UO_93 (O_93,N_18314,N_19642);
nor UO_94 (O_94,N_17326,N_17785);
nor UO_95 (O_95,N_18842,N_17358);
nand UO_96 (O_96,N_16442,N_18879);
nand UO_97 (O_97,N_17972,N_15340);
xor UO_98 (O_98,N_15063,N_17450);
and UO_99 (O_99,N_19338,N_18046);
or UO_100 (O_100,N_19582,N_15500);
xnor UO_101 (O_101,N_15837,N_19451);
or UO_102 (O_102,N_17654,N_17115);
nand UO_103 (O_103,N_19133,N_18930);
nor UO_104 (O_104,N_17049,N_15371);
and UO_105 (O_105,N_17286,N_17878);
nand UO_106 (O_106,N_16560,N_16233);
and UO_107 (O_107,N_17403,N_17860);
nor UO_108 (O_108,N_15184,N_16854);
nor UO_109 (O_109,N_16585,N_16927);
nand UO_110 (O_110,N_15280,N_18558);
or UO_111 (O_111,N_15081,N_15427);
or UO_112 (O_112,N_16255,N_19196);
xnor UO_113 (O_113,N_19541,N_19102);
and UO_114 (O_114,N_18369,N_19288);
nand UO_115 (O_115,N_16121,N_17222);
and UO_116 (O_116,N_18048,N_19607);
and UO_117 (O_117,N_18083,N_15335);
or UO_118 (O_118,N_17656,N_17879);
and UO_119 (O_119,N_17817,N_17529);
or UO_120 (O_120,N_18523,N_16533);
xnor UO_121 (O_121,N_15497,N_19261);
nand UO_122 (O_122,N_18283,N_16104);
nor UO_123 (O_123,N_16532,N_19965);
nand UO_124 (O_124,N_18448,N_18603);
and UO_125 (O_125,N_19371,N_17619);
and UO_126 (O_126,N_15482,N_16174);
or UO_127 (O_127,N_16294,N_16074);
or UO_128 (O_128,N_18037,N_17940);
or UO_129 (O_129,N_19191,N_18292);
xor UO_130 (O_130,N_19867,N_18704);
nand UO_131 (O_131,N_17740,N_15705);
or UO_132 (O_132,N_16341,N_16984);
or UO_133 (O_133,N_17352,N_15444);
and UO_134 (O_134,N_18379,N_15205);
and UO_135 (O_135,N_18002,N_19446);
xor UO_136 (O_136,N_18786,N_19844);
nand UO_137 (O_137,N_16768,N_15972);
or UO_138 (O_138,N_18171,N_16939);
and UO_139 (O_139,N_17392,N_19050);
or UO_140 (O_140,N_16340,N_18654);
or UO_141 (O_141,N_15720,N_19055);
and UO_142 (O_142,N_19916,N_16950);
nor UO_143 (O_143,N_19961,N_19121);
nand UO_144 (O_144,N_19552,N_17241);
xnor UO_145 (O_145,N_19900,N_16850);
or UO_146 (O_146,N_15954,N_17330);
or UO_147 (O_147,N_17601,N_18095);
and UO_148 (O_148,N_16346,N_19235);
or UO_149 (O_149,N_18127,N_15667);
and UO_150 (O_150,N_16913,N_18093);
nand UO_151 (O_151,N_16057,N_18264);
and UO_152 (O_152,N_16093,N_19304);
nor UO_153 (O_153,N_18895,N_17744);
nor UO_154 (O_154,N_15975,N_18186);
nor UO_155 (O_155,N_16623,N_18373);
xor UO_156 (O_156,N_17252,N_15087);
and UO_157 (O_157,N_16193,N_15319);
and UO_158 (O_158,N_16140,N_15440);
nand UO_159 (O_159,N_19504,N_17094);
or UO_160 (O_160,N_19680,N_16961);
and UO_161 (O_161,N_16214,N_18661);
nand UO_162 (O_162,N_17451,N_19886);
or UO_163 (O_163,N_18228,N_17600);
and UO_164 (O_164,N_15199,N_16662);
or UO_165 (O_165,N_17145,N_18069);
xnor UO_166 (O_166,N_16138,N_17910);
nor UO_167 (O_167,N_16428,N_19227);
or UO_168 (O_168,N_15886,N_15161);
xnor UO_169 (O_169,N_18101,N_16277);
xnor UO_170 (O_170,N_15707,N_18642);
nor UO_171 (O_171,N_18567,N_15283);
nand UO_172 (O_172,N_16010,N_19718);
or UO_173 (O_173,N_19518,N_15459);
and UO_174 (O_174,N_17590,N_15771);
and UO_175 (O_175,N_16184,N_19405);
nor UO_176 (O_176,N_19113,N_18853);
xor UO_177 (O_177,N_16336,N_15879);
nand UO_178 (O_178,N_19818,N_18335);
and UO_179 (O_179,N_16988,N_16364);
xnor UO_180 (O_180,N_19801,N_15800);
and UO_181 (O_181,N_16643,N_19852);
and UO_182 (O_182,N_17553,N_16631);
nand UO_183 (O_183,N_19084,N_19699);
and UO_184 (O_184,N_15944,N_16026);
nor UO_185 (O_185,N_19181,N_19460);
or UO_186 (O_186,N_16418,N_15825);
or UO_187 (O_187,N_16251,N_18787);
nor UO_188 (O_188,N_19401,N_15036);
and UO_189 (O_189,N_17107,N_16484);
and UO_190 (O_190,N_16622,N_17555);
and UO_191 (O_191,N_16180,N_17746);
nand UO_192 (O_192,N_15169,N_19800);
or UO_193 (O_193,N_16168,N_19299);
xor UO_194 (O_194,N_16593,N_17368);
xnor UO_195 (O_195,N_17249,N_19981);
nand UO_196 (O_196,N_18226,N_19698);
nand UO_197 (O_197,N_16246,N_15020);
xnor UO_198 (O_198,N_15366,N_15343);
xnor UO_199 (O_199,N_16655,N_17081);
nor UO_200 (O_200,N_15926,N_17536);
nand UO_201 (O_201,N_17385,N_19658);
xor UO_202 (O_202,N_16359,N_17008);
or UO_203 (O_203,N_18504,N_18598);
nor UO_204 (O_204,N_15328,N_15594);
nand UO_205 (O_205,N_18395,N_16853);
or UO_206 (O_206,N_17768,N_16818);
or UO_207 (O_207,N_19041,N_15992);
nor UO_208 (O_208,N_15209,N_15960);
nand UO_209 (O_209,N_18794,N_18266);
nor UO_210 (O_210,N_15661,N_19962);
xnor UO_211 (O_211,N_17560,N_19535);
nor UO_212 (O_212,N_18063,N_16176);
nand UO_213 (O_213,N_18952,N_16367);
nand UO_214 (O_214,N_18616,N_16330);
xnor UO_215 (O_215,N_17609,N_16740);
nor UO_216 (O_216,N_19621,N_17036);
or UO_217 (O_217,N_18991,N_18769);
nand UO_218 (O_218,N_19914,N_17797);
xor UO_219 (O_219,N_16273,N_17023);
and UO_220 (O_220,N_16189,N_15748);
or UO_221 (O_221,N_18542,N_18110);
and UO_222 (O_222,N_17690,N_17843);
nand UO_223 (O_223,N_17979,N_19119);
and UO_224 (O_224,N_15387,N_19361);
or UO_225 (O_225,N_18235,N_16043);
nand UO_226 (O_226,N_16157,N_18575);
and UO_227 (O_227,N_16786,N_18424);
nor UO_228 (O_228,N_19287,N_18672);
or UO_229 (O_229,N_19613,N_16384);
nand UO_230 (O_230,N_18832,N_15969);
xor UO_231 (O_231,N_17623,N_17966);
and UO_232 (O_232,N_19210,N_15406);
xor UO_233 (O_233,N_17615,N_18820);
or UO_234 (O_234,N_17752,N_16765);
nor UO_235 (O_235,N_15362,N_18281);
nor UO_236 (O_236,N_16029,N_16125);
nor UO_237 (O_237,N_19078,N_17111);
xnor UO_238 (O_238,N_15701,N_18195);
or UO_239 (O_239,N_18249,N_15562);
nand UO_240 (O_240,N_17221,N_17870);
and UO_241 (O_241,N_16612,N_19874);
nand UO_242 (O_242,N_15861,N_19285);
nor UO_243 (O_243,N_16117,N_17779);
and UO_244 (O_244,N_16414,N_18595);
or UO_245 (O_245,N_18144,N_17833);
and UO_246 (O_246,N_15256,N_18321);
nor UO_247 (O_247,N_17956,N_18791);
and UO_248 (O_248,N_18131,N_18086);
or UO_249 (O_249,N_17635,N_17194);
nor UO_250 (O_250,N_19184,N_15419);
nor UO_251 (O_251,N_18541,N_18601);
and UO_252 (O_252,N_17331,N_17837);
and UO_253 (O_253,N_15865,N_17945);
xor UO_254 (O_254,N_18524,N_16441);
nor UO_255 (O_255,N_17304,N_19489);
and UO_256 (O_256,N_15460,N_17563);
nor UO_257 (O_257,N_16943,N_17215);
xor UO_258 (O_258,N_18625,N_16099);
or UO_259 (O_259,N_17132,N_19855);
nor UO_260 (O_260,N_19348,N_16672);
nand UO_261 (O_261,N_16290,N_19245);
or UO_262 (O_262,N_16695,N_15620);
and UO_263 (O_263,N_19100,N_17495);
and UO_264 (O_264,N_15799,N_16997);
and UO_265 (O_265,N_18118,N_15269);
and UO_266 (O_266,N_16163,N_16555);
xor UO_267 (O_267,N_17112,N_16975);
nand UO_268 (O_268,N_17416,N_16582);
nand UO_269 (O_269,N_18647,N_15791);
or UO_270 (O_270,N_18818,N_15742);
or UO_271 (O_271,N_15483,N_15421);
xnor UO_272 (O_272,N_19030,N_18089);
nand UO_273 (O_273,N_17181,N_19204);
nor UO_274 (O_274,N_15465,N_19960);
xnor UO_275 (O_275,N_15076,N_18464);
and UO_276 (O_276,N_18351,N_15962);
nand UO_277 (O_277,N_17171,N_19683);
and UO_278 (O_278,N_18332,N_17751);
nor UO_279 (O_279,N_18475,N_18490);
nand UO_280 (O_280,N_17724,N_17268);
nand UO_281 (O_281,N_19665,N_15030);
nand UO_282 (O_282,N_17976,N_18531);
nor UO_283 (O_283,N_18922,N_18682);
and UO_284 (O_284,N_17127,N_18646);
nand UO_285 (O_285,N_17935,N_19688);
nor UO_286 (O_286,N_16385,N_19606);
or UO_287 (O_287,N_19180,N_18695);
and UO_288 (O_288,N_17144,N_16938);
xor UO_289 (O_289,N_18840,N_19561);
and UO_290 (O_290,N_18586,N_16335);
nor UO_291 (O_291,N_18271,N_19595);
or UO_292 (O_292,N_18837,N_18688);
nand UO_293 (O_293,N_17586,N_19177);
or UO_294 (O_294,N_19885,N_17104);
or UO_295 (O_295,N_17454,N_18354);
nor UO_296 (O_296,N_16307,N_15289);
nand UO_297 (O_297,N_15875,N_17986);
xor UO_298 (O_298,N_18297,N_18337);
and UO_299 (O_299,N_18802,N_16198);
or UO_300 (O_300,N_16921,N_15505);
or UO_301 (O_301,N_16956,N_15598);
xnor UO_302 (O_302,N_18707,N_19270);
or UO_303 (O_303,N_17630,N_18554);
nand UO_304 (O_304,N_15566,N_16457);
xor UO_305 (O_305,N_15626,N_15860);
nor UO_306 (O_306,N_16159,N_15047);
and UO_307 (O_307,N_15390,N_15980);
nor UO_308 (O_308,N_17253,N_16937);
nand UO_309 (O_309,N_16507,N_17977);
or UO_310 (O_310,N_16706,N_16628);
nand UO_311 (O_311,N_18296,N_17647);
or UO_312 (O_312,N_17649,N_17761);
or UO_313 (O_313,N_16312,N_18461);
nand UO_314 (O_314,N_17517,N_16406);
and UO_315 (O_315,N_16637,N_16248);
nor UO_316 (O_316,N_18154,N_16386);
or UO_317 (O_317,N_16617,N_15512);
nand UO_318 (O_318,N_18062,N_16035);
nor UO_319 (O_319,N_17841,N_19301);
or UO_320 (O_320,N_18877,N_19298);
xnor UO_321 (O_321,N_15520,N_19482);
or UO_322 (O_322,N_16080,N_15925);
or UO_323 (O_323,N_15264,N_18725);
nor UO_324 (O_324,N_16746,N_16109);
xnor UO_325 (O_325,N_17223,N_18906);
and UO_326 (O_326,N_15422,N_16887);
and UO_327 (O_327,N_18416,N_16470);
nand UO_328 (O_328,N_19546,N_16985);
nor UO_329 (O_329,N_17384,N_15055);
xnor UO_330 (O_330,N_19033,N_19789);
nor UO_331 (O_331,N_16916,N_16542);
xnor UO_332 (O_332,N_16841,N_17942);
and UO_333 (O_333,N_18078,N_15545);
xnor UO_334 (O_334,N_15163,N_18363);
xor UO_335 (O_335,N_16050,N_19765);
nand UO_336 (O_336,N_16068,N_18451);
nor UO_337 (O_337,N_17265,N_19796);
and UO_338 (O_338,N_18483,N_19964);
nor UO_339 (O_339,N_15525,N_15593);
or UO_340 (O_340,N_19467,N_16016);
or UO_341 (O_341,N_16941,N_17731);
or UO_342 (O_342,N_16280,N_16439);
and UO_343 (O_343,N_17711,N_17031);
nor UO_344 (O_344,N_19501,N_18810);
and UO_345 (O_345,N_18339,N_17754);
nand UO_346 (O_346,N_15431,N_17357);
and UO_347 (O_347,N_16333,N_15333);
xnor UO_348 (O_348,N_17418,N_19841);
or UO_349 (O_349,N_19506,N_18724);
nor UO_350 (O_350,N_16696,N_19938);
xor UO_351 (O_351,N_19399,N_17152);
nor UO_352 (O_352,N_18663,N_18900);
nand UO_353 (O_353,N_19329,N_18910);
nor UO_354 (O_354,N_16142,N_17749);
xnor UO_355 (O_355,N_17533,N_19445);
or UO_356 (O_356,N_18834,N_16027);
nor UO_357 (O_357,N_18020,N_19407);
and UO_358 (O_358,N_15190,N_17446);
nor UO_359 (O_359,N_15696,N_19802);
or UO_360 (O_360,N_16134,N_17160);
xnor UO_361 (O_361,N_16419,N_19466);
nand UO_362 (O_362,N_15652,N_17655);
or UO_363 (O_363,N_18773,N_18718);
nor UO_364 (O_364,N_16565,N_18259);
and UO_365 (O_365,N_15416,N_15339);
xor UO_366 (O_366,N_19540,N_16570);
xor UO_367 (O_367,N_16636,N_18066);
and UO_368 (O_368,N_16394,N_17309);
nand UO_369 (O_369,N_16583,N_18948);
nand UO_370 (O_370,N_18613,N_17695);
or UO_371 (O_371,N_18177,N_19478);
and UO_372 (O_372,N_19409,N_16102);
nand UO_373 (O_373,N_19334,N_16285);
nand UO_374 (O_374,N_18227,N_19963);
nor UO_375 (O_375,N_17991,N_18254);
and UO_376 (O_376,N_16949,N_19311);
nor UO_377 (O_377,N_17733,N_19381);
xor UO_378 (O_378,N_19206,N_15494);
xnor UO_379 (O_379,N_19282,N_18324);
or UO_380 (O_380,N_18611,N_18135);
or UO_381 (O_381,N_17428,N_17516);
or UO_382 (O_382,N_17261,N_18286);
and UO_383 (O_383,N_15029,N_19866);
xor UO_384 (O_384,N_16085,N_16855);
nand UO_385 (O_385,N_19107,N_16714);
and UO_386 (O_386,N_18053,N_16795);
nor UO_387 (O_387,N_17925,N_18427);
nor UO_388 (O_388,N_19721,N_19168);
nor UO_389 (O_389,N_16592,N_19643);
or UO_390 (O_390,N_18942,N_19160);
nand UO_391 (O_391,N_16569,N_17931);
and UO_392 (O_392,N_17013,N_15107);
nor UO_393 (O_393,N_15041,N_15716);
nor UO_394 (O_394,N_15766,N_18711);
xnor UO_395 (O_395,N_16712,N_17508);
and UO_396 (O_396,N_16191,N_19375);
nor UO_397 (O_397,N_19322,N_16078);
xnor UO_398 (O_398,N_19070,N_16177);
nand UO_399 (O_399,N_17786,N_18027);
xnor UO_400 (O_400,N_19937,N_19269);
nand UO_401 (O_401,N_17321,N_19890);
nand UO_402 (O_402,N_15734,N_15847);
xnor UO_403 (O_403,N_19488,N_19252);
or UO_404 (O_404,N_17079,N_17566);
and UO_405 (O_405,N_16807,N_16503);
or UO_406 (O_406,N_19116,N_19336);
nand UO_407 (O_407,N_15352,N_18277);
nand UO_408 (O_408,N_15392,N_16584);
nand UO_409 (O_409,N_19707,N_17394);
nand UO_410 (O_410,N_16328,N_19536);
and UO_411 (O_411,N_18931,N_15900);
nor UO_412 (O_412,N_15329,N_18623);
xnor UO_413 (O_413,N_17891,N_17681);
and UO_414 (O_414,N_19719,N_19862);
or UO_415 (O_415,N_19942,N_16674);
nand UO_416 (O_416,N_15842,N_19264);
and UO_417 (O_417,N_15389,N_15220);
and UO_418 (O_418,N_19215,N_15065);
nor UO_419 (O_419,N_15931,N_16865);
nor UO_420 (O_420,N_18674,N_17857);
xor UO_421 (O_421,N_18352,N_17381);
xor UO_422 (O_422,N_19392,N_16630);
or UO_423 (O_423,N_18460,N_16812);
nor UO_424 (O_424,N_18013,N_18176);
and UO_425 (O_425,N_18447,N_18081);
nand UO_426 (O_426,N_16034,N_15874);
xor UO_427 (O_427,N_17796,N_15784);
or UO_428 (O_428,N_19414,N_19522);
or UO_429 (O_429,N_19520,N_18898);
and UO_430 (O_430,N_18382,N_15524);
and UO_431 (O_431,N_17825,N_19850);
nand UO_432 (O_432,N_17633,N_15348);
xor UO_433 (O_433,N_17067,N_17686);
and UO_434 (O_434,N_15388,N_19693);
or UO_435 (O_435,N_19218,N_15298);
nor UO_436 (O_436,N_17073,N_18726);
and UO_437 (O_437,N_17435,N_15834);
or UO_438 (O_438,N_16751,N_15173);
and UO_439 (O_439,N_16421,N_18675);
nor UO_440 (O_440,N_17227,N_19017);
and UO_441 (O_441,N_18391,N_18164);
xor UO_442 (O_442,N_19975,N_16310);
nor UO_443 (O_443,N_15675,N_15051);
nand UO_444 (O_444,N_17608,N_16263);
and UO_445 (O_445,N_17757,N_15178);
or UO_446 (O_446,N_17387,N_17770);
and UO_447 (O_447,N_16095,N_16116);
or UO_448 (O_448,N_16815,N_16410);
nand UO_449 (O_449,N_18604,N_17958);
xor UO_450 (O_450,N_19058,N_17414);
or UO_451 (O_451,N_16045,N_15100);
xor UO_452 (O_452,N_19363,N_19587);
nor UO_453 (O_453,N_15779,N_19545);
nand UO_454 (O_454,N_18882,N_19835);
nor UO_455 (O_455,N_18445,N_19555);
nand UO_456 (O_456,N_15133,N_18233);
xnor UO_457 (O_457,N_15832,N_15284);
xnor UO_458 (O_458,N_16862,N_19290);
nor UO_459 (O_459,N_15773,N_19563);
or UO_460 (O_460,N_17110,N_16828);
or UO_461 (O_461,N_15804,N_19925);
nand UO_462 (O_462,N_19230,N_17612);
and UO_463 (O_463,N_19007,N_18963);
nor UO_464 (O_464,N_19984,N_16929);
nor UO_465 (O_465,N_16574,N_15257);
and UO_466 (O_466,N_18153,N_15844);
nand UO_467 (O_467,N_19767,N_15909);
nor UO_468 (O_468,N_18540,N_16811);
and UO_469 (O_469,N_18894,N_17844);
xnor UO_470 (O_470,N_16651,N_16368);
xnor UO_471 (O_471,N_19758,N_16126);
or UO_472 (O_472,N_18720,N_18771);
nand UO_473 (O_473,N_16388,N_16909);
and UO_474 (O_474,N_17808,N_18302);
and UO_475 (O_475,N_19921,N_18859);
xor UO_476 (O_476,N_15088,N_19697);
nand UO_477 (O_477,N_19247,N_19172);
xor UO_478 (O_478,N_18516,N_17278);
nor UO_479 (O_479,N_17277,N_15203);
nand UO_480 (O_480,N_15619,N_16401);
and UO_481 (O_481,N_15449,N_18715);
xnor UO_482 (O_482,N_18309,N_19366);
xnor UO_483 (O_483,N_17621,N_19876);
nand UO_484 (O_484,N_19878,N_16413);
or UO_485 (O_485,N_18319,N_16567);
or UO_486 (O_486,N_17175,N_15086);
nor UO_487 (O_487,N_16953,N_18643);
nor UO_488 (O_488,N_17420,N_18741);
xor UO_489 (O_489,N_15447,N_18462);
xor UO_490 (O_490,N_16652,N_18861);
or UO_491 (O_491,N_17541,N_15515);
xnor UO_492 (O_492,N_19592,N_17210);
and UO_493 (O_493,N_16741,N_19112);
xor UO_494 (O_494,N_16882,N_15364);
nand UO_495 (O_495,N_19428,N_15462);
xor UO_496 (O_496,N_18417,N_18824);
nor UO_497 (O_497,N_19918,N_17396);
or UO_498 (O_498,N_15827,N_18169);
or UO_499 (O_499,N_16028,N_18518);
and UO_500 (O_500,N_16389,N_18232);
nand UO_501 (O_501,N_16973,N_16001);
xor UO_502 (O_502,N_15144,N_15246);
and UO_503 (O_503,N_19067,N_19532);
nor UO_504 (O_504,N_16370,N_19724);
xnor UO_505 (O_505,N_18156,N_15835);
and UO_506 (O_506,N_17054,N_16185);
and UO_507 (O_507,N_17741,N_19879);
xor UO_508 (O_508,N_17374,N_15979);
or UO_509 (O_509,N_16424,N_15755);
nor UO_510 (O_510,N_15225,N_17123);
or UO_511 (O_511,N_15774,N_18536);
and UO_512 (O_512,N_18560,N_19842);
and UO_513 (O_513,N_19672,N_15300);
nor UO_514 (O_514,N_19819,N_15457);
nor UO_515 (O_515,N_15655,N_18848);
or UO_516 (O_516,N_15783,N_15785);
xor UO_517 (O_517,N_19562,N_17100);
nand UO_518 (O_518,N_18916,N_18023);
and UO_519 (O_519,N_18624,N_15223);
nand UO_520 (O_520,N_15495,N_19933);
nand UO_521 (O_521,N_18493,N_15239);
xnor UO_522 (O_522,N_17226,N_15657);
or UO_523 (O_523,N_15633,N_18355);
or UO_524 (O_524,N_17791,N_16902);
nor UO_525 (O_525,N_17103,N_15775);
nand UO_526 (O_526,N_17472,N_15991);
and UO_527 (O_527,N_19054,N_18669);
nand UO_528 (O_528,N_17128,N_18912);
or UO_529 (O_529,N_16014,N_15547);
xnor UO_530 (O_530,N_17047,N_15400);
or UO_531 (O_531,N_16092,N_18222);
nand UO_532 (O_532,N_16249,N_18781);
nor UO_533 (O_533,N_18320,N_15288);
nor UO_534 (O_534,N_17447,N_15105);
and UO_535 (O_535,N_16797,N_15893);
nor UO_536 (O_536,N_18673,N_15396);
nand UO_537 (O_537,N_17691,N_16201);
or UO_538 (O_538,N_17663,N_16237);
nand UO_539 (O_539,N_17017,N_18392);
nand UO_540 (O_540,N_15439,N_16947);
nand UO_541 (O_541,N_17137,N_18471);
xor UO_542 (O_542,N_19286,N_17706);
nor UO_543 (O_543,N_17642,N_19081);
or UO_544 (O_544,N_18733,N_15595);
nor UO_545 (O_545,N_18179,N_15623);
nor UO_546 (O_546,N_16875,N_17433);
nor UO_547 (O_547,N_18237,N_17509);
nor UO_548 (O_548,N_16239,N_15822);
or UO_549 (O_549,N_18032,N_18344);
nand UO_550 (O_550,N_18433,N_17238);
nand UO_551 (O_551,N_16474,N_17548);
and UO_552 (O_552,N_19028,N_16101);
nand UO_553 (O_553,N_18430,N_15591);
nor UO_554 (O_554,N_17375,N_18617);
and UO_555 (O_555,N_15132,N_15083);
and UO_556 (O_556,N_17888,N_17760);
nand UO_557 (O_557,N_16979,N_16356);
nand UO_558 (O_558,N_17676,N_19155);
and UO_559 (O_559,N_15709,N_19514);
nor UO_560 (O_560,N_17528,N_17355);
or UO_561 (O_561,N_19732,N_19704);
xnor UO_562 (O_562,N_15222,N_17329);
and UO_563 (O_563,N_15202,N_16864);
and UO_564 (O_564,N_18985,N_18317);
and UO_565 (O_565,N_15005,N_16250);
nor UO_566 (O_566,N_18090,N_19720);
xor UO_567 (O_567,N_15942,N_18476);
nor UO_568 (O_568,N_16256,N_16279);
and UO_569 (O_569,N_18678,N_19397);
xnor UO_570 (O_570,N_18058,N_18021);
nor UO_571 (O_571,N_15430,N_17921);
and UO_572 (O_572,N_18744,N_16179);
and UO_573 (O_573,N_16325,N_17102);
or UO_574 (O_574,N_16781,N_18602);
xnor UO_575 (O_575,N_17781,N_16734);
nor UO_576 (O_576,N_19158,N_15790);
and UO_577 (O_577,N_18644,N_19741);
nand UO_578 (O_578,N_17719,N_17954);
xor UO_579 (O_579,N_16155,N_16132);
nor UO_580 (O_580,N_19560,N_17356);
or UO_581 (O_581,N_17183,N_16331);
xor UO_582 (O_582,N_18357,N_17009);
nor UO_583 (O_583,N_18989,N_15079);
nor UO_584 (O_584,N_17320,N_15091);
xnor UO_585 (O_585,N_15853,N_15404);
or UO_586 (O_586,N_19473,N_18147);
and UO_587 (O_587,N_19778,N_16486);
and UO_588 (O_588,N_17313,N_16297);
nand UO_589 (O_589,N_15188,N_15628);
nand UO_590 (O_590,N_18734,N_19123);
or UO_591 (O_591,N_17971,N_19632);
nand UO_592 (O_592,N_19432,N_18494);
nor UO_593 (O_593,N_19509,N_17486);
nor UO_594 (O_594,N_17704,N_15978);
nand UO_595 (O_595,N_18425,N_19894);
and UO_596 (O_596,N_16422,N_18075);
and UO_597 (O_597,N_17895,N_18189);
nor UO_598 (O_598,N_18736,N_18619);
xor UO_599 (O_599,N_16599,N_16378);
nor UO_600 (O_600,N_19659,N_18050);
or UO_601 (O_601,N_15863,N_17788);
nand UO_602 (O_602,N_19803,N_17605);
nor UO_603 (O_603,N_16880,N_15112);
xor UO_604 (O_604,N_18767,N_16520);
xor UO_605 (O_605,N_17502,N_19060);
nand UO_606 (O_606,N_15772,N_15224);
xnor UO_607 (O_607,N_15367,N_19284);
xnor UO_608 (O_608,N_19439,N_16692);
nand UO_609 (O_609,N_16742,N_18641);
and UO_610 (O_610,N_15870,N_17675);
or UO_611 (O_611,N_19453,N_17595);
and UO_612 (O_612,N_18330,N_15561);
and UO_613 (O_613,N_18632,N_17873);
or UO_614 (O_614,N_19496,N_15743);
and UO_615 (O_615,N_15833,N_16369);
xnor UO_616 (O_616,N_18977,N_15458);
and UO_617 (O_617,N_18491,N_19549);
nand UO_618 (O_618,N_18913,N_17410);
nor UO_619 (O_619,N_17907,N_17544);
nor UO_620 (O_620,N_19306,N_19547);
nor UO_621 (O_621,N_15732,N_15058);
or UO_622 (O_622,N_17543,N_18645);
xnor UO_623 (O_623,N_18936,N_19309);
nor UO_624 (O_624,N_18774,N_18811);
xnor UO_625 (O_625,N_17874,N_19339);
nand UO_626 (O_626,N_19584,N_17620);
xnor UO_627 (O_627,N_17498,N_18938);
nand UO_628 (O_628,N_19174,N_16650);
xor UO_629 (O_629,N_15405,N_18770);
xnor UO_630 (O_630,N_18808,N_15078);
or UO_631 (O_631,N_19099,N_17371);
nand UO_632 (O_632,N_17134,N_19888);
nand UO_633 (O_633,N_17060,N_15237);
nor UO_634 (O_634,N_19024,N_16225);
nor UO_635 (O_635,N_17193,N_19701);
nor UO_636 (O_636,N_19932,N_16519);
and UO_637 (O_637,N_15736,N_17148);
xnor UO_638 (O_638,N_16411,N_19000);
xnor UO_639 (O_639,N_18262,N_19822);
nor UO_640 (O_640,N_17559,N_17572);
and UO_641 (O_641,N_15946,N_19036);
nand UO_642 (O_642,N_18231,N_16989);
nand UO_643 (O_643,N_16113,N_19421);
xnor UO_644 (O_644,N_15207,N_19328);
and UO_645 (O_645,N_16430,N_15901);
or UO_646 (O_646,N_19838,N_15303);
or UO_647 (O_647,N_17307,N_16833);
xnor UO_648 (O_648,N_16845,N_15843);
nor UO_649 (O_649,N_16767,N_18854);
xor UO_650 (O_650,N_15508,N_19679);
nor UO_651 (O_651,N_17665,N_16986);
and UO_652 (O_652,N_16923,N_16645);
and UO_653 (O_653,N_15892,N_17598);
and UO_654 (O_654,N_15026,N_18294);
nand UO_655 (O_655,N_15649,N_16365);
or UO_656 (O_656,N_16877,N_17184);
nor UO_657 (O_657,N_15453,N_18001);
or UO_658 (O_658,N_18520,N_17674);
nand UO_659 (O_659,N_16338,N_16453);
or UO_660 (O_660,N_16429,N_19736);
xnor UO_661 (O_661,N_16586,N_17002);
or UO_662 (O_662,N_16087,N_17968);
nand UO_663 (O_663,N_15729,N_17561);
and UO_664 (O_664,N_19182,N_19650);
and UO_665 (O_665,N_15093,N_19412);
xor UO_666 (O_666,N_18485,N_17989);
nand UO_667 (O_667,N_19193,N_18061);
nor UO_668 (O_668,N_19438,N_15008);
or UO_669 (O_669,N_16918,N_18489);
nor UO_670 (O_670,N_19226,N_17993);
or UO_671 (O_671,N_15571,N_15252);
and UO_672 (O_672,N_19739,N_17306);
nor UO_673 (O_673,N_17696,N_15151);
or UO_674 (O_674,N_17263,N_15956);
nand UO_675 (O_675,N_19202,N_15070);
or UO_676 (O_676,N_17807,N_16173);
nor UO_677 (O_677,N_17231,N_19833);
nand UO_678 (O_678,N_15877,N_19212);
nor UO_679 (O_679,N_19811,N_16488);
nor UO_680 (O_680,N_17577,N_16701);
nor UO_681 (O_681,N_17197,N_18280);
nand UO_682 (O_682,N_18003,N_19088);
nand UO_683 (O_683,N_19185,N_16613);
xor UO_684 (O_684,N_17494,N_17007);
nor UO_685 (O_685,N_15891,N_19791);
or UO_686 (O_686,N_18621,N_15197);
or UO_687 (O_687,N_18103,N_15118);
xnor UO_688 (O_688,N_15911,N_15471);
nand UO_689 (O_689,N_16402,N_16888);
nor UO_690 (O_690,N_16464,N_17432);
or UO_691 (O_691,N_16576,N_18634);
nor UO_692 (O_692,N_17671,N_19941);
nor UO_693 (O_693,N_15728,N_19839);
and UO_694 (O_694,N_17985,N_19877);
nand UO_695 (O_695,N_19591,N_19408);
or UO_696 (O_696,N_16258,N_18148);
and UO_697 (O_697,N_18064,N_17892);
or UO_698 (O_698,N_19576,N_17489);
nor UO_699 (O_699,N_15052,N_17168);
nand UO_700 (O_700,N_17748,N_18405);
nand UO_701 (O_701,N_19300,N_17445);
nor UO_702 (O_702,N_16903,N_18009);
and UO_703 (O_703,N_17510,N_19858);
and UO_704 (O_704,N_16883,N_19608);
and UO_705 (O_705,N_17087,N_17201);
nor UO_706 (O_706,N_17325,N_16849);
xor UO_707 (O_707,N_19893,N_16536);
xor UO_708 (O_708,N_17068,N_15386);
nand UO_709 (O_709,N_19234,N_17994);
nand UO_710 (O_710,N_17312,N_15350);
or UO_711 (O_711,N_16377,N_19075);
nand UO_712 (O_712,N_18030,N_18123);
nand UO_713 (O_713,N_18610,N_17003);
or UO_714 (O_714,N_18772,N_18782);
or UO_715 (O_715,N_19051,N_19823);
xnor UO_716 (O_716,N_19687,N_16420);
xnor UO_717 (O_717,N_17712,N_17596);
nor UO_718 (O_718,N_18126,N_15022);
and UO_719 (O_719,N_19690,N_15399);
nor UO_720 (O_720,N_15579,N_16164);
or UO_721 (O_721,N_16483,N_15688);
nand UO_722 (O_722,N_17750,N_16412);
nor UO_723 (O_723,N_18846,N_16788);
xnor UO_724 (O_724,N_18596,N_19061);
nand UO_725 (O_725,N_19875,N_15710);
or UO_726 (O_726,N_17980,N_16200);
and UO_727 (O_727,N_17272,N_15316);
and UO_728 (O_728,N_18128,N_18035);
nand UO_729 (O_729,N_17581,N_16186);
or UO_730 (O_730,N_17289,N_15485);
nor UO_731 (O_731,N_16496,N_18188);
xnor UO_732 (O_732,N_19859,N_19426);
and UO_733 (O_733,N_19967,N_17095);
nand UO_734 (O_734,N_15745,N_19686);
or UO_735 (O_735,N_15856,N_16195);
nor UO_736 (O_736,N_15606,N_18055);
nand UO_737 (O_737,N_18158,N_17531);
xnor UO_738 (O_738,N_17395,N_19612);
nor UO_739 (O_739,N_17296,N_18289);
and UO_740 (O_740,N_17195,N_18085);
xor UO_741 (O_741,N_15238,N_15446);
and UO_742 (O_742,N_18325,N_19769);
nand UO_743 (O_743,N_16676,N_17061);
nor UO_744 (O_744,N_16146,N_17923);
nor UO_745 (O_745,N_16607,N_18775);
xor UO_746 (O_746,N_19785,N_15928);
xor UO_747 (O_747,N_15415,N_17092);
and UO_748 (O_748,N_15308,N_19383);
nor UO_749 (O_749,N_16881,N_18551);
nand UO_750 (O_750,N_17518,N_15687);
and UO_751 (O_751,N_15168,N_17129);
and UO_752 (O_752,N_15636,N_16391);
and UO_753 (O_753,N_15480,N_16573);
or UO_754 (O_754,N_15479,N_19619);
xor UO_755 (O_755,N_16626,N_18829);
and UO_756 (O_756,N_17011,N_15680);
nand UO_757 (O_757,N_15072,N_15027);
nor UO_758 (O_758,N_19125,N_15206);
nor UO_759 (O_759,N_17669,N_19080);
and UO_760 (O_760,N_17897,N_15689);
and UO_761 (O_761,N_16188,N_17349);
xnor UO_762 (O_762,N_18209,N_18282);
nor UO_763 (O_763,N_18974,N_19843);
nand UO_764 (O_764,N_17041,N_19799);
or UO_765 (O_765,N_19332,N_19251);
xnor UO_766 (O_766,N_16079,N_18284);
or UO_767 (O_767,N_18178,N_19458);
and UO_768 (O_768,N_15868,N_15473);
nand UO_769 (O_769,N_19996,N_16287);
or UO_770 (O_770,N_18970,N_19278);
or UO_771 (O_771,N_19709,N_15527);
nor UO_772 (O_772,N_15381,N_19188);
nand UO_773 (O_773,N_18394,N_16575);
or UO_774 (O_774,N_18367,N_17119);
nor UO_775 (O_775,N_16928,N_18559);
or UO_776 (O_776,N_17303,N_16925);
nor UO_777 (O_777,N_17190,N_19905);
or UO_778 (O_778,N_15630,N_15988);
xor UO_779 (O_779,N_18679,N_17383);
nor UO_780 (O_780,N_18323,N_16703);
nor UO_781 (O_781,N_17708,N_17801);
nand UO_782 (O_782,N_15839,N_18071);
or UO_783 (O_783,N_18138,N_19706);
or UO_784 (O_784,N_19810,N_15312);
xor UO_785 (O_785,N_18470,N_18114);
nor UO_786 (O_786,N_16466,N_15254);
nand UO_787 (O_787,N_19779,N_19114);
or UO_788 (O_788,N_16379,N_17153);
xor UO_789 (O_789,N_15477,N_17444);
nand UO_790 (O_790,N_15271,N_15539);
or UO_791 (O_791,N_16914,N_15582);
nor UO_792 (O_792,N_17082,N_17298);
xor UO_793 (O_793,N_17783,N_18935);
or UO_794 (O_794,N_18562,N_15690);
or UO_795 (O_795,N_17800,N_18010);
nand UO_796 (O_796,N_18386,N_19064);
nor UO_797 (O_797,N_18505,N_15442);
or UO_798 (O_798,N_17736,N_17248);
xnor UO_799 (O_799,N_17946,N_17499);
xnor UO_800 (O_800,N_15073,N_16096);
nand UO_801 (O_801,N_19516,N_19795);
or UO_802 (O_802,N_16405,N_19487);
nand UO_803 (O_803,N_17480,N_16284);
and UO_804 (O_804,N_16669,N_17636);
or UO_805 (O_805,N_19143,N_19127);
nand UO_806 (O_806,N_15260,N_19640);
xnor UO_807 (O_807,N_16244,N_16175);
or UO_808 (O_808,N_15621,N_17101);
or UO_809 (O_809,N_16160,N_18640);
or UO_810 (O_810,N_18535,N_19471);
nor UO_811 (O_811,N_15551,N_17846);
and UO_812 (O_812,N_17662,N_17276);
nand UO_813 (O_813,N_17650,N_19376);
or UO_814 (O_814,N_18236,N_19231);
or UO_815 (O_815,N_15085,N_15050);
xnor UO_816 (O_816,N_19244,N_18962);
xnor UO_817 (O_817,N_18513,N_19258);
nor UO_818 (O_818,N_18361,N_16587);
and UO_819 (O_819,N_15934,N_19087);
xnor UO_820 (O_820,N_17188,N_19015);
and UO_821 (O_821,N_16036,N_17066);
xor UO_822 (O_822,N_17063,N_16679);
nor UO_823 (O_823,N_18742,N_15176);
nor UO_824 (O_824,N_19834,N_18702);
or UO_825 (O_825,N_15369,N_15121);
nand UO_826 (O_826,N_16639,N_15614);
or UO_827 (O_827,N_18785,N_18225);
and UO_828 (O_828,N_18615,N_19583);
and UO_829 (O_829,N_18574,N_19250);
or UO_830 (O_830,N_15491,N_15746);
nor UO_831 (O_831,N_15454,N_15888);
nand UO_832 (O_832,N_15607,N_18496);
or UO_833 (O_833,N_18517,N_16445);
or UO_834 (O_834,N_16752,N_18527);
and UO_835 (O_835,N_16900,N_19730);
nand UO_836 (O_836,N_16206,N_17462);
or UO_837 (O_837,N_18511,N_15533);
nor UO_838 (O_838,N_16403,N_19737);
or UO_839 (O_839,N_17220,N_17078);
xnor UO_840 (O_840,N_19870,N_17481);
and UO_841 (O_841,N_18200,N_19840);
and UO_842 (O_842,N_17348,N_18788);
and UO_843 (O_843,N_18018,N_15681);
nor UO_844 (O_844,N_16885,N_17950);
or UO_845 (O_845,N_17767,N_15098);
nand UO_846 (O_846,N_15276,N_17467);
and UO_847 (O_847,N_17056,N_15986);
nand UO_848 (O_848,N_18637,N_17315);
nand UO_849 (O_849,N_19615,N_16697);
xnor UO_850 (O_850,N_18486,N_18187);
xnor UO_851 (O_851,N_16737,N_18146);
xor UO_852 (O_852,N_17851,N_17365);
xor UO_853 (O_853,N_17027,N_18731);
or UO_854 (O_854,N_18946,N_15243);
nor UO_855 (O_855,N_17709,N_16322);
nand UO_856 (O_856,N_15544,N_17822);
xnor UO_857 (O_857,N_18017,N_16606);
xnor UO_858 (O_858,N_15417,N_16726);
xor UO_859 (O_859,N_17440,N_16624);
or UO_860 (O_860,N_15857,N_16139);
xnor UO_861 (O_861,N_17701,N_18529);
xor UO_862 (O_862,N_17269,N_15914);
nand UO_863 (O_863,N_16192,N_16537);
nand UO_864 (O_864,N_16874,N_18329);
nand UO_865 (O_865,N_16813,N_18174);
or UO_866 (O_866,N_17497,N_18334);
or UO_867 (O_867,N_15990,N_17154);
and UO_868 (O_868,N_15060,N_15854);
xor UO_869 (O_869,N_15142,N_16578);
xor UO_870 (O_870,N_17850,N_19098);
and UO_871 (O_871,N_19310,N_17710);
nand UO_872 (O_872,N_19138,N_17077);
and UO_873 (O_873,N_16962,N_16047);
and UO_874 (O_874,N_19105,N_18890);
nand UO_875 (O_875,N_19742,N_15625);
and UO_876 (O_876,N_16824,N_18639);
or UO_877 (O_877,N_17699,N_19902);
or UO_878 (O_878,N_16506,N_19904);
nand UO_879 (O_879,N_19935,N_19579);
xor UO_880 (O_880,N_16736,N_16148);
and UO_881 (O_881,N_15658,N_16397);
nand UO_882 (O_882,N_16572,N_15115);
or UO_883 (O_883,N_18850,N_17626);
and UO_884 (O_884,N_15426,N_19274);
and UO_885 (O_885,N_18500,N_19132);
or UO_886 (O_886,N_17549,N_16694);
and UO_887 (O_887,N_19783,N_19165);
and UO_888 (O_888,N_18313,N_18800);
xnor UO_889 (O_889,N_19853,N_19297);
xnor UO_890 (O_890,N_19343,N_19717);
xor UO_891 (O_891,N_15738,N_17545);
or UO_892 (O_892,N_15816,N_15000);
and UO_893 (O_893,N_17351,N_16303);
nand UO_894 (O_894,N_16042,N_19848);
nor UO_895 (O_895,N_17550,N_18047);
xnor UO_896 (O_896,N_15824,N_15012);
or UO_897 (O_897,N_19969,N_17680);
nand UO_898 (O_898,N_16708,N_18571);
or UO_899 (O_899,N_15718,N_15624);
nand UO_900 (O_900,N_19447,N_18550);
and UO_901 (O_901,N_16931,N_15379);
and UO_902 (O_902,N_16725,N_15492);
xnor UO_903 (O_903,N_18996,N_19347);
or UO_904 (O_904,N_15821,N_16810);
nor UO_905 (O_905,N_18370,N_19437);
or UO_906 (O_906,N_17339,N_18253);
or UO_907 (O_907,N_18396,N_15296);
xnor UO_908 (O_908,N_17141,N_16067);
or UO_909 (O_909,N_17698,N_15177);
xnor UO_910 (O_910,N_19892,N_18303);
or UO_911 (O_911,N_19611,N_15851);
or UO_912 (O_912,N_17959,N_19669);
and UO_913 (O_913,N_19868,N_19479);
nand UO_914 (O_914,N_17855,N_15812);
nor UO_915 (O_915,N_19021,N_15974);
nand UO_916 (O_916,N_18468,N_18076);
nand UO_917 (O_917,N_17960,N_19930);
or UO_918 (O_918,N_19083,N_18659);
and UO_919 (O_919,N_18004,N_19574);
nand UO_920 (O_920,N_16683,N_18487);
and UO_921 (O_921,N_17282,N_16127);
nor UO_922 (O_922,N_19425,N_17540);
nand UO_923 (O_923,N_16693,N_15698);
xor UO_924 (O_924,N_17173,N_16274);
nand UO_925 (O_925,N_15071,N_17573);
or UO_926 (O_926,N_18564,N_18658);
xor UO_927 (O_927,N_19847,N_17802);
nand UO_928 (O_928,N_18932,N_18124);
nor UO_929 (O_929,N_19623,N_15671);
or UO_930 (O_930,N_17804,N_19920);
or UO_931 (O_931,N_15255,N_19530);
or UO_932 (O_932,N_18484,N_16891);
xnor UO_933 (O_933,N_16111,N_15004);
and UO_934 (O_934,N_17794,N_16739);
or UO_935 (O_935,N_18839,N_19846);
nand UO_936 (O_936,N_15164,N_17334);
and UO_937 (O_937,N_19148,N_18687);
nor UO_938 (O_938,N_18552,N_15189);
or UO_939 (O_939,N_17667,N_17599);
and UO_940 (O_940,N_15964,N_15683);
and UO_941 (O_941,N_17199,N_17981);
nor UO_942 (O_942,N_16744,N_17827);
or UO_943 (O_943,N_18753,N_16106);
or UO_944 (O_944,N_15691,N_18219);
nor UO_945 (O_945,N_16500,N_17936);
or UO_946 (O_946,N_18175,N_15382);
nand UO_947 (O_947,N_17146,N_15331);
and UO_948 (O_948,N_17224,N_17242);
or UO_949 (O_949,N_16878,N_18727);
and UO_950 (O_950,N_19952,N_16710);
or UO_951 (O_951,N_18721,N_16245);
and UO_952 (O_952,N_15370,N_15951);
or UO_953 (O_953,N_16832,N_16238);
and UO_954 (O_954,N_18299,N_19221);
and UO_955 (O_955,N_16868,N_17281);
xnor UO_956 (O_956,N_19229,N_19341);
or UO_957 (O_957,N_18691,N_18269);
nor UO_958 (O_958,N_19523,N_18212);
or UO_959 (O_959,N_19131,N_16844);
xnor UO_960 (O_960,N_16505,N_17212);
and UO_961 (O_961,N_17233,N_17730);
or UO_962 (O_962,N_18426,N_19089);
nor UO_963 (O_963,N_17521,N_18409);
or UO_964 (O_964,N_17885,N_18909);
nor UO_965 (O_965,N_17039,N_16771);
xor UO_966 (O_966,N_16048,N_18198);
nor UO_967 (O_967,N_16292,N_15245);
nand UO_968 (O_968,N_15433,N_15410);
and UO_969 (O_969,N_18402,N_19043);
nand UO_970 (O_970,N_16720,N_15730);
or UO_971 (O_971,N_15611,N_17952);
and UO_972 (O_972,N_16664,N_16088);
nor UO_973 (O_973,N_18039,N_16353);
xor UO_974 (O_974,N_18152,N_16763);
nand UO_975 (O_975,N_15513,N_15368);
nand UO_976 (O_976,N_18893,N_18275);
xnor UO_977 (O_977,N_15126,N_19910);
nor UO_978 (O_978,N_19924,N_15314);
and UO_979 (O_979,N_17664,N_17915);
or UO_980 (O_980,N_18353,N_17225);
nor UO_981 (O_981,N_15514,N_19194);
nand UO_982 (O_982,N_17015,N_15936);
and UO_983 (O_983,N_15155,N_17089);
or UO_984 (O_984,N_15391,N_18419);
nor UO_985 (O_985,N_17311,N_18803);
nand UO_986 (O_986,N_18383,N_15357);
nand UO_987 (O_987,N_15638,N_17759);
xor UO_988 (O_988,N_17948,N_18815);
nand UO_989 (O_989,N_18056,N_15703);
nor UO_990 (O_990,N_16382,N_16657);
nor UO_991 (O_991,N_18959,N_15420);
xnor UO_992 (O_992,N_19956,N_19416);
xor UO_993 (O_993,N_17743,N_17828);
nor UO_994 (O_994,N_18184,N_19597);
xor UO_995 (O_995,N_18905,N_17064);
or UO_996 (O_996,N_17125,N_17771);
xor UO_997 (O_997,N_18988,N_18388);
nor UO_998 (O_998,N_16473,N_17914);
nand UO_999 (O_999,N_19677,N_16219);
nor UO_1000 (O_1000,N_15963,N_17042);
xnor UO_1001 (O_1001,N_17020,N_17526);
nor UO_1002 (O_1002,N_17344,N_19825);
or UO_1003 (O_1003,N_17147,N_19167);
nand UO_1004 (O_1004,N_16158,N_19817);
and UO_1005 (O_1005,N_16407,N_19660);
nand UO_1006 (O_1006,N_15217,N_15920);
and UO_1007 (O_1007,N_16857,N_17668);
and UO_1008 (O_1008,N_16872,N_19289);
and UO_1009 (O_1009,N_18929,N_19668);
nand UO_1010 (O_1010,N_17504,N_17496);
nand UO_1011 (O_1011,N_17159,N_19936);
and UO_1012 (O_1012,N_18092,N_19012);
or UO_1013 (O_1013,N_18925,N_19272);
or UO_1014 (O_1014,N_19593,N_19225);
nand UO_1015 (O_1015,N_16063,N_16064);
nor UO_1016 (O_1016,N_16448,N_17546);
nand UO_1017 (O_1017,N_15463,N_19533);
and UO_1018 (O_1018,N_18343,N_19360);
nor UO_1019 (O_1019,N_18421,N_19388);
and UO_1020 (O_1020,N_18276,N_15109);
xor UO_1021 (O_1021,N_15156,N_18501);
nand UO_1022 (O_1022,N_15583,N_17350);
nand UO_1023 (O_1023,N_19176,N_15818);
xnor UO_1024 (O_1024,N_16020,N_18028);
xnor UO_1025 (O_1025,N_17611,N_18965);
nand UO_1026 (O_1026,N_19118,N_19821);
nand UO_1027 (O_1027,N_18581,N_16234);
nor UO_1028 (O_1028,N_15798,N_18310);
or UO_1029 (O_1029,N_18580,N_16450);
nand UO_1030 (O_1030,N_19386,N_18958);
nand UO_1031 (O_1031,N_17883,N_15552);
nor UO_1032 (O_1032,N_16959,N_19346);
and UO_1033 (O_1033,N_19553,N_17722);
nor UO_1034 (O_1034,N_17574,N_18155);
or UO_1035 (O_1035,N_17211,N_18220);
nand UO_1036 (O_1036,N_19749,N_19410);
nand UO_1037 (O_1037,N_16524,N_18211);
or UO_1038 (O_1038,N_17911,N_15456);
or UO_1039 (O_1039,N_17864,N_16323);
xnor UO_1040 (O_1040,N_18761,N_18943);
nand UO_1041 (O_1041,N_19510,N_16907);
or UO_1042 (O_1042,N_16564,N_18975);
nor UO_1043 (O_1043,N_15792,N_19380);
nor UO_1044 (O_1044,N_16416,N_19856);
nand UO_1045 (O_1045,N_17941,N_18107);
nand UO_1046 (O_1046,N_18122,N_16595);
xnor UO_1047 (O_1047,N_17192,N_19771);
nand UO_1048 (O_1048,N_18453,N_17346);
nor UO_1049 (O_1049,N_17789,N_19154);
and UO_1050 (O_1050,N_18561,N_19013);
nor UO_1051 (O_1051,N_16523,N_15193);
nor UO_1052 (O_1052,N_16196,N_16803);
nand UO_1053 (O_1053,N_19647,N_17205);
nor UO_1054 (O_1054,N_16351,N_19213);
and UO_1055 (O_1055,N_16659,N_18662);
xor UO_1056 (O_1056,N_17872,N_19122);
nand UO_1057 (O_1057,N_15397,N_15375);
or UO_1058 (O_1058,N_16301,N_17438);
nand UO_1059 (O_1059,N_15568,N_16625);
and UO_1060 (O_1060,N_15760,N_18413);
or UO_1061 (O_1061,N_18359,N_15913);
or UO_1062 (O_1062,N_17524,N_16546);
and UO_1063 (O_1063,N_17511,N_18706);
or UO_1064 (O_1064,N_18748,N_18982);
nand UO_1065 (O_1065,N_18224,N_18557);
or UO_1066 (O_1066,N_16337,N_15849);
and UO_1067 (O_1067,N_15501,N_16764);
and UO_1068 (O_1068,N_17273,N_17470);
xor UO_1069 (O_1069,N_18134,N_17271);
or UO_1070 (O_1070,N_19074,N_18137);
nand UO_1071 (O_1071,N_17639,N_15862);
nor UO_1072 (O_1072,N_18229,N_15546);
or UO_1073 (O_1073,N_17232,N_18404);
nand UO_1074 (O_1074,N_18680,N_17593);
nand UO_1075 (O_1075,N_15059,N_16785);
nor UO_1076 (O_1076,N_18008,N_15213);
or UO_1077 (O_1077,N_19831,N_19944);
and UO_1078 (O_1078,N_17607,N_16796);
nor UO_1079 (O_1079,N_18902,N_18326);
and UO_1080 (O_1080,N_17406,N_15136);
xor UO_1081 (O_1081,N_18290,N_15735);
or UO_1082 (O_1082,N_15038,N_16922);
xnor UO_1083 (O_1083,N_18579,N_15137);
nand UO_1084 (O_1084,N_16432,N_19404);
nor UO_1085 (O_1085,N_15737,N_17747);
xor UO_1086 (O_1086,N_17984,N_18257);
xor UO_1087 (O_1087,N_17890,N_16400);
nand UO_1088 (O_1088,N_16002,N_19023);
nand UO_1089 (O_1089,N_17254,N_18094);
xor UO_1090 (O_1090,N_16502,N_19784);
and UO_1091 (O_1091,N_15437,N_15102);
xnor UO_1092 (O_1092,N_17987,N_19203);
or UO_1093 (O_1093,N_19394,N_17963);
nand UO_1094 (O_1094,N_15970,N_15787);
nand UO_1095 (O_1095,N_15504,N_17133);
and UO_1096 (O_1096,N_19757,N_19691);
xnor UO_1097 (O_1097,N_16830,N_19774);
or UO_1098 (O_1098,N_17539,N_18950);
and UO_1099 (O_1099,N_18630,N_16999);
nor UO_1100 (O_1100,N_19805,N_16128);
or UO_1101 (O_1101,N_16462,N_15301);
nor UO_1102 (O_1102,N_16153,N_16012);
nand UO_1103 (O_1103,N_18428,N_18838);
and UO_1104 (O_1104,N_16780,N_19657);
and UO_1105 (O_1105,N_16278,N_17955);
nor UO_1106 (O_1106,N_19519,N_15434);
nand UO_1107 (O_1107,N_18278,N_17294);
or UO_1108 (O_1108,N_18293,N_16105);
xnor UO_1109 (O_1109,N_18307,N_16228);
xnor UO_1110 (O_1110,N_19145,N_16769);
xnor UO_1111 (O_1111,N_19164,N_15903);
xor UO_1112 (O_1112,N_19256,N_15326);
or UO_1113 (O_1113,N_15104,N_15971);
and UO_1114 (O_1114,N_18247,N_16444);
xnor UO_1115 (O_1115,N_15143,N_15204);
nor UO_1116 (O_1116,N_17848,N_15248);
nand UO_1117 (O_1117,N_19998,N_17646);
nor UO_1118 (O_1118,N_18801,N_17360);
and UO_1119 (O_1119,N_18696,N_15094);
nor UO_1120 (O_1120,N_16596,N_16963);
xor UO_1121 (O_1121,N_15618,N_18173);
or UO_1122 (O_1122,N_19670,N_18981);
nand UO_1123 (O_1123,N_17430,N_15057);
nor UO_1124 (O_1124,N_16008,N_15996);
nand UO_1125 (O_1125,N_19664,N_16236);
or UO_1126 (O_1126,N_15639,N_15578);
xnor UO_1127 (O_1127,N_15106,N_19763);
nor UO_1128 (O_1128,N_16952,N_16717);
or UO_1129 (O_1129,N_16745,N_16481);
nand UO_1130 (O_1130,N_15803,N_16527);
nor UO_1131 (O_1131,N_17404,N_19836);
nor UO_1132 (O_1132,N_18686,N_15496);
nor UO_1133 (O_1133,N_15749,N_18548);
xor UO_1134 (O_1134,N_16081,N_18435);
and UO_1135 (O_1135,N_15793,N_19790);
and UO_1136 (O_1136,N_18026,N_15466);
or UO_1137 (O_1137,N_15037,N_18568);
and UO_1138 (O_1138,N_18999,N_16633);
nand UO_1139 (O_1139,N_17402,N_15414);
and UO_1140 (O_1140,N_16216,N_15325);
or UO_1141 (O_1141,N_15506,N_15398);
xnor UO_1142 (O_1142,N_17473,N_15966);
and UO_1143 (O_1143,N_19271,N_15899);
or UO_1144 (O_1144,N_18102,N_15317);
or UO_1145 (O_1145,N_17436,N_15981);
xnor UO_1146 (O_1146,N_15383,N_19201);
nor UO_1147 (O_1147,N_15219,N_17769);
and UO_1148 (O_1148,N_16794,N_19813);
xnor UO_1149 (O_1149,N_19884,N_18578);
nand UO_1150 (O_1150,N_19475,N_19863);
nor UO_1151 (O_1151,N_17016,N_16750);
nand UO_1152 (O_1152,N_16347,N_16272);
nand UO_1153 (O_1153,N_17969,N_19880);
xnor UO_1154 (O_1154,N_17927,N_17030);
or UO_1155 (O_1155,N_15487,N_18526);
nor UO_1156 (O_1156,N_17679,N_19344);
nand UO_1157 (O_1157,N_17932,N_19400);
or UO_1158 (O_1158,N_19333,N_15664);
and UO_1159 (O_1159,N_18538,N_16493);
or UO_1160 (O_1160,N_19515,N_15858);
nor UO_1161 (O_1161,N_19951,N_18347);
nor UO_1162 (O_1162,N_19987,N_19147);
and UO_1163 (O_1163,N_19178,N_17142);
xor UO_1164 (O_1164,N_17957,N_16354);
and UO_1165 (O_1165,N_16062,N_15338);
and UO_1166 (O_1166,N_17424,N_17179);
nand UO_1167 (O_1167,N_17475,N_18566);
nor UO_1168 (O_1168,N_16137,N_16122);
or UO_1169 (O_1169,N_19187,N_19911);
or UO_1170 (O_1170,N_19768,N_18749);
and UO_1171 (O_1171,N_16075,N_16601);
or UO_1172 (O_1172,N_16817,N_16309);
xor UO_1173 (O_1173,N_17028,N_19891);
nor UO_1174 (O_1174,N_16793,N_16404);
xor UO_1175 (O_1175,N_18546,N_19556);
xnor UO_1176 (O_1176,N_15349,N_15122);
nand UO_1177 (O_1177,N_15567,N_17018);
nand UO_1178 (O_1178,N_19525,N_15907);
nor UO_1179 (O_1179,N_17943,N_16467);
xor UO_1180 (O_1180,N_18883,N_19974);
or UO_1181 (O_1181,N_16904,N_15311);
nand UO_1182 (O_1182,N_15830,N_16472);
nand UO_1183 (O_1183,N_17459,N_18979);
xnor UO_1184 (O_1184,N_17845,N_18246);
and UO_1185 (O_1185,N_17322,N_15165);
nand UO_1186 (O_1186,N_17214,N_15418);
or UO_1187 (O_1187,N_18285,N_16261);
and UO_1188 (O_1188,N_15806,N_17821);
nor UO_1189 (O_1189,N_18831,N_16946);
and UO_1190 (O_1190,N_18657,N_15565);
and UO_1191 (O_1191,N_16151,N_18288);
xnor UO_1192 (O_1192,N_19170,N_17863);
and UO_1193 (O_1193,N_19559,N_16876);
and UO_1194 (O_1194,N_16054,N_17139);
nand UO_1195 (O_1195,N_17965,N_15183);
nor UO_1196 (O_1196,N_15345,N_19435);
or UO_1197 (O_1197,N_19101,N_18701);
xnor UO_1198 (O_1198,N_15939,N_15542);
or UO_1199 (O_1199,N_18305,N_16315);
and UO_1200 (O_1200,N_15097,N_18036);
and UO_1201 (O_1201,N_18449,N_18054);
nand UO_1202 (O_1202,N_16487,N_15763);
or UO_1203 (O_1203,N_15315,N_18474);
nor UO_1204 (O_1204,N_17568,N_15187);
nand UO_1205 (O_1205,N_15075,N_19223);
nor UO_1206 (O_1206,N_18876,N_19108);
xor UO_1207 (O_1207,N_16066,N_18406);
and UO_1208 (O_1208,N_18250,N_18492);
xnor UO_1209 (O_1209,N_15194,N_18031);
xnor UO_1210 (O_1210,N_19379,N_18287);
nor UO_1211 (O_1211,N_15915,N_17345);
nor UO_1212 (O_1212,N_19266,N_19512);
and UO_1213 (O_1213,N_16461,N_16118);
and UO_1214 (O_1214,N_15175,N_15577);
xor UO_1215 (O_1215,N_18044,N_19494);
and UO_1216 (O_1216,N_17301,N_19678);
and UO_1217 (O_1217,N_19627,N_15432);
or UO_1218 (O_1218,N_19581,N_16077);
or UO_1219 (O_1219,N_15240,N_16729);
nor UO_1220 (O_1220,N_15230,N_15605);
or UO_1221 (O_1221,N_15930,N_17995);
nand UO_1222 (O_1222,N_16051,N_18185);
nand UO_1223 (O_1223,N_17762,N_19806);
xor UO_1224 (O_1224,N_19093,N_18034);
xnor UO_1225 (O_1225,N_19524,N_15517);
and UO_1226 (O_1226,N_16856,N_19947);
nor UO_1227 (O_1227,N_16253,N_16314);
and UO_1228 (O_1228,N_16267,N_18903);
xnor UO_1229 (O_1229,N_15987,N_19599);
xor UO_1230 (O_1230,N_19486,N_17575);
or UO_1231 (O_1231,N_19503,N_19354);
or UO_1232 (O_1232,N_16704,N_15559);
and UO_1233 (O_1233,N_18584,N_16058);
nor UO_1234 (O_1234,N_15778,N_15233);
nor UO_1235 (O_1235,N_17250,N_17207);
nand UO_1236 (O_1236,N_19430,N_16760);
or UO_1237 (O_1237,N_16271,N_19395);
and UO_1238 (O_1238,N_16119,N_17672);
or UO_1239 (O_1239,N_18993,N_15977);
nor UO_1240 (O_1240,N_16531,N_17328);
nor UO_1241 (O_1241,N_17460,N_18328);
and UO_1242 (O_1242,N_18479,N_19006);
nand UO_1243 (O_1243,N_17255,N_15526);
or UO_1244 (O_1244,N_16425,N_17466);
or UO_1245 (O_1245,N_17648,N_19216);
nor UO_1246 (O_1246,N_17569,N_17973);
nand UO_1247 (O_1247,N_16544,N_19715);
or UO_1248 (O_1248,N_16688,N_15353);
and UO_1249 (O_1249,N_18358,N_18390);
nor UO_1250 (O_1250,N_18265,N_17659);
or UO_1251 (O_1251,N_18240,N_15448);
nand UO_1252 (O_1252,N_19422,N_19899);
xor UO_1253 (O_1253,N_15721,N_16753);
nand UO_1254 (O_1254,N_15344,N_18514);
nor UO_1255 (O_1255,N_15534,N_16492);
or UO_1256 (O_1256,N_18508,N_18097);
or UO_1257 (O_1257,N_17852,N_16580);
or UO_1258 (O_1258,N_15139,N_16390);
xnor UO_1259 (O_1259,N_16232,N_19815);
nand UO_1260 (O_1260,N_17723,N_16288);
nand UO_1261 (O_1261,N_15185,N_19505);
nor UO_1262 (O_1262,N_16589,N_15117);
nor UO_1263 (O_1263,N_17505,N_18889);
nand UO_1264 (O_1264,N_15941,N_19586);
nor UO_1265 (O_1265,N_17742,N_15385);
nand UO_1266 (O_1266,N_17834,N_16073);
and UO_1267 (O_1267,N_18964,N_18132);
and UO_1268 (O_1268,N_19211,N_16262);
nor UO_1269 (O_1269,N_15172,N_17666);
xnor UO_1270 (O_1270,N_15033,N_17084);
or UO_1271 (O_1271,N_17949,N_15796);
or UO_1272 (O_1272,N_15108,N_15200);
or UO_1273 (O_1273,N_15813,N_19685);
nand UO_1274 (O_1274,N_18349,N_15519);
or UO_1275 (O_1275,N_19882,N_16656);
nand UO_1276 (O_1276,N_17218,N_19129);
and UO_1277 (O_1277,N_17717,N_16859);
xor UO_1278 (O_1278,N_18650,N_19387);
nor UO_1279 (O_1279,N_16522,N_18756);
nand UO_1280 (O_1280,N_17917,N_19531);
or UO_1281 (O_1281,N_15923,N_16908);
and UO_1282 (O_1282,N_19483,N_19103);
nand UO_1283 (O_1283,N_16009,N_18049);
nor UO_1284 (O_1284,N_18377,N_15080);
nor UO_1285 (O_1285,N_16826,N_15585);
or UO_1286 (O_1286,N_16415,N_15904);
nand UO_1287 (O_1287,N_19600,N_19110);
and UO_1288 (O_1288,N_17046,N_16178);
xnor UO_1289 (O_1289,N_18088,N_17918);
or UO_1290 (O_1290,N_15895,N_16013);
nor UO_1291 (O_1291,N_16352,N_17640);
nand UO_1292 (O_1292,N_17055,N_18631);
or UO_1293 (O_1293,N_16836,N_15261);
nand UO_1294 (O_1294,N_15634,N_15242);
xor UO_1295 (O_1295,N_16534,N_16721);
and UO_1296 (O_1296,N_18865,N_16269);
nor UO_1297 (O_1297,N_18677,N_18019);
and UO_1298 (O_1298,N_16821,N_19331);
and UO_1299 (O_1299,N_19232,N_19047);
xnor UO_1300 (O_1300,N_16082,N_16779);
or UO_1301 (O_1301,N_19016,N_18442);
or UO_1302 (O_1302,N_19319,N_18255);
xnor UO_1303 (O_1303,N_17809,N_19279);
nor UO_1304 (O_1304,N_19927,N_18378);
nor UO_1305 (O_1305,N_15757,N_16556);
and UO_1306 (O_1306,N_19010,N_16342);
nand UO_1307 (O_1307,N_18139,N_15159);
nor UO_1308 (O_1308,N_16747,N_16498);
xor UO_1309 (O_1309,N_19092,N_19162);
xor UO_1310 (O_1310,N_19156,N_15695);
and UO_1311 (O_1311,N_16282,N_19820);
or UO_1312 (O_1312,N_18213,N_19069);
and UO_1313 (O_1313,N_15945,N_17778);
nor UO_1314 (O_1314,N_15581,N_17262);
nand UO_1315 (O_1315,N_19255,N_15855);
nand UO_1316 (O_1316,N_16183,N_18012);
xor UO_1317 (O_1317,N_17702,N_15601);
and UO_1318 (O_1318,N_19303,N_16434);
or UO_1319 (O_1319,N_18745,N_18267);
nand UO_1320 (O_1320,N_16529,N_16642);
nor UO_1321 (O_1321,N_18423,N_15758);
xor UO_1322 (O_1322,N_15445,N_18585);
xor UO_1323 (O_1323,N_18628,N_19782);
and UO_1324 (O_1324,N_17790,N_15692);
nand UO_1325 (O_1325,N_16684,N_16863);
xnor UO_1326 (O_1326,N_19728,N_16969);
or UO_1327 (O_1327,N_17185,N_17764);
and UO_1328 (O_1328,N_17021,N_16766);
nor UO_1329 (O_1329,N_18863,N_16667);
and UO_1330 (O_1330,N_15616,N_17734);
nand UO_1331 (O_1331,N_16504,N_15795);
nor UO_1332 (O_1332,N_19746,N_16086);
nand UO_1333 (O_1333,N_18162,N_17122);
nand UO_1334 (O_1334,N_16668,N_17876);
xor UO_1335 (O_1335,N_17155,N_18896);
and UO_1336 (O_1336,N_15068,N_15668);
nor UO_1337 (O_1337,N_16313,N_19302);
and UO_1338 (O_1338,N_15660,N_18754);
xor UO_1339 (O_1339,N_15642,N_18341);
nand UO_1340 (O_1340,N_16935,N_16743);
nor UO_1341 (O_1341,N_19418,N_19094);
nor UO_1342 (O_1342,N_19972,N_19978);
or UO_1343 (O_1343,N_18274,N_18626);
and UO_1344 (O_1344,N_19955,N_18141);
xor UO_1345 (O_1345,N_19320,N_17186);
xor UO_1346 (O_1346,N_18751,N_19610);
or UO_1347 (O_1347,N_18594,N_17689);
xnor UO_1348 (O_1348,N_17811,N_16289);
xor UO_1349 (O_1349,N_18515,N_16912);
nand UO_1350 (O_1350,N_15146,N_18593);
or UO_1351 (O_1351,N_16658,N_15018);
or UO_1352 (O_1352,N_16431,N_18572);
or UO_1353 (O_1353,N_16663,N_15140);
or UO_1354 (O_1354,N_15599,N_18618);
or UO_1355 (O_1355,N_19571,N_19695);
and UO_1356 (O_1356,N_15236,N_15395);
xnor UO_1357 (O_1357,N_18258,N_16458);
xor UO_1358 (O_1358,N_17182,N_18374);
or UO_1359 (O_1359,N_17434,N_19276);
nand UO_1360 (O_1360,N_15472,N_17335);
or UO_1361 (O_1361,N_18418,N_19169);
and UO_1362 (O_1362,N_18823,N_17130);
nor UO_1363 (O_1363,N_17124,N_18336);
and UO_1364 (O_1364,N_15275,N_19915);
nand UO_1365 (O_1365,N_17069,N_17347);
or UO_1366 (O_1366,N_16616,N_18768);
or UO_1367 (O_1367,N_15918,N_18133);
or UO_1368 (O_1368,N_19059,N_19837);
nand UO_1369 (O_1369,N_15826,N_17442);
xnor UO_1370 (O_1370,N_16690,N_15150);
nor UO_1371 (O_1371,N_16635,N_19217);
and UO_1372 (O_1372,N_15876,N_19452);
nor UO_1373 (O_1373,N_18555,N_15304);
nor UO_1374 (O_1374,N_18565,N_16772);
and UO_1375 (O_1375,N_15166,N_16044);
xor UO_1376 (O_1376,N_17727,N_16053);
xnor UO_1377 (O_1377,N_17051,N_16770);
and UO_1378 (O_1378,N_18070,N_19906);
nor UO_1379 (O_1379,N_16559,N_17576);
or UO_1380 (O_1380,N_15129,N_18065);
xnor UO_1381 (O_1381,N_15747,N_19490);
nand UO_1382 (O_1382,N_19469,N_18660);
and UO_1383 (O_1383,N_15119,N_19751);
and UO_1384 (O_1384,N_19979,N_16296);
and UO_1385 (O_1385,N_15282,N_17579);
nor UO_1386 (O_1386,N_19040,N_18648);
nor UO_1387 (O_1387,N_17838,N_15880);
xor UO_1388 (O_1388,N_18119,N_18304);
nand UO_1389 (O_1389,N_19631,N_17823);
nor UO_1390 (O_1390,N_16226,N_15927);
or UO_1391 (O_1391,N_19048,N_15464);
nand UO_1392 (O_1392,N_19943,N_19588);
or UO_1393 (O_1393,N_15235,N_17006);
nand UO_1394 (O_1394,N_16716,N_19472);
xor UO_1395 (O_1395,N_15921,N_19513);
or UO_1396 (O_1396,N_15884,N_18530);
nand UO_1397 (O_1397,N_19617,N_17370);
and UO_1398 (O_1398,N_19444,N_19362);
nor UO_1399 (O_1399,N_18308,N_17816);
and UO_1400 (O_1400,N_19318,N_17096);
and UO_1401 (O_1401,N_16893,N_16561);
xnor UO_1402 (O_1402,N_15299,N_18533);
nor UO_1403 (O_1403,N_18722,N_16417);
nor UO_1404 (O_1404,N_18084,N_18583);
or UO_1405 (O_1405,N_16843,N_19468);
nor UO_1406 (O_1406,N_16678,N_18685);
and UO_1407 (O_1407,N_15488,N_18636);
nor UO_1408 (O_1408,N_16114,N_18006);
xnor UO_1409 (O_1409,N_19495,N_15120);
and UO_1410 (O_1410,N_19674,N_17862);
xor UO_1411 (O_1411,N_15467,N_16890);
xor UO_1412 (O_1412,N_15007,N_15377);
nor UO_1413 (O_1413,N_16408,N_19171);
xnor UO_1414 (O_1414,N_15789,N_17739);
or UO_1415 (O_1415,N_15478,N_19692);
nor UO_1416 (O_1416,N_15509,N_15887);
nand UO_1417 (O_1417,N_18059,N_18432);
nand UO_1418 (O_1418,N_17482,N_18956);
xor UO_1419 (O_1419,N_16698,N_15522);
nand UO_1420 (O_1420,N_18954,N_19097);
nand UO_1421 (O_1421,N_17391,N_19770);
xor UO_1422 (O_1422,N_17478,N_17455);
or UO_1423 (O_1423,N_16510,N_16037);
or UO_1424 (O_1424,N_15556,N_17483);
or UO_1425 (O_1425,N_16071,N_15503);
or UO_1426 (O_1426,N_16005,N_15171);
nor UO_1427 (O_1427,N_17274,N_18864);
or UO_1428 (O_1428,N_16597,N_16514);
nor UO_1429 (O_1429,N_16171,N_15906);
xnor UO_1430 (O_1430,N_18609,N_19804);
nor UO_1431 (O_1431,N_15077,N_16229);
nand UO_1432 (O_1432,N_15372,N_19305);
nor UO_1433 (O_1433,N_16748,N_17398);
and UO_1434 (O_1434,N_15035,N_18150);
xnor UO_1435 (O_1435,N_19345,N_18480);
nand UO_1436 (O_1436,N_15617,N_15560);
xnor UO_1437 (O_1437,N_17978,N_18263);
or UO_1438 (O_1438,N_17080,N_15937);
nor UO_1439 (O_1439,N_17091,N_16648);
or UO_1440 (O_1440,N_17425,N_15024);
nor UO_1441 (O_1441,N_15531,N_18990);
xor UO_1442 (O_1442,N_16298,N_18251);
nor UO_1443 (O_1443,N_17228,N_16387);
or UO_1444 (O_1444,N_17097,N_17697);
or UO_1445 (O_1445,N_18509,N_17728);
nor UO_1446 (O_1446,N_18521,N_16754);
nor UO_1447 (O_1447,N_16478,N_16320);
nand UO_1448 (O_1448,N_17587,N_18828);
xnor UO_1449 (O_1449,N_18544,N_17106);
nand UO_1450 (O_1450,N_17682,N_17109);
or UO_1451 (O_1451,N_16161,N_17400);
xor UO_1452 (O_1452,N_16355,N_16981);
or UO_1453 (O_1453,N_17501,N_15147);
nor UO_1454 (O_1454,N_15741,N_15231);
xnor UO_1455 (O_1455,N_16089,N_17288);
nor UO_1456 (O_1456,N_15435,N_18796);
and UO_1457 (O_1457,N_15229,N_16252);
nand UO_1458 (O_1458,N_19263,N_15016);
nor UO_1459 (O_1459,N_19968,N_16072);
or UO_1460 (O_1460,N_16711,N_19992);
or UO_1461 (O_1461,N_18159,N_15622);
nand UO_1462 (O_1462,N_17437,N_18532);
or UO_1463 (O_1463,N_15273,N_17260);
nand UO_1464 (O_1464,N_15873,N_18510);
nand UO_1465 (O_1465,N_16240,N_15550);
nor UO_1466 (O_1466,N_18201,N_15359);
and UO_1467 (O_1467,N_18739,N_18011);
or UO_1468 (O_1468,N_15917,N_17390);
and UO_1469 (O_1469,N_17924,N_18372);
nor UO_1470 (O_1470,N_15686,N_18627);
or UO_1471 (O_1471,N_16515,N_15998);
and UO_1472 (O_1472,N_17287,N_17552);
nor UO_1473 (O_1473,N_15540,N_17525);
or UO_1474 (O_1474,N_15541,N_17052);
xor UO_1475 (O_1475,N_16305,N_15609);
nor UO_1476 (O_1476,N_15321,N_18921);
nor UO_1477 (O_1477,N_18190,N_17953);
nand UO_1478 (O_1478,N_18477,N_18106);
nand UO_1479 (O_1479,N_16598,N_17040);
nand UO_1480 (O_1480,N_17251,N_18888);
xor UO_1481 (O_1481,N_17093,N_18368);
or UO_1482 (O_1482,N_15309,N_16735);
nand UO_1483 (O_1483,N_19772,N_19389);
xor UO_1484 (O_1484,N_17174,N_17213);
or UO_1485 (O_1485,N_15848,N_18995);
nor UO_1486 (O_1486,N_16361,N_17401);
nand UO_1487 (O_1487,N_18466,N_16069);
and UO_1488 (O_1488,N_17468,N_18366);
nand UO_1489 (O_1489,N_16451,N_16557);
and UO_1490 (O_1490,N_19253,N_19293);
and UO_1491 (O_1491,N_17849,N_15378);
xor UO_1492 (O_1492,N_16490,N_15090);
xor UO_1493 (O_1493,N_18041,N_17735);
and UO_1494 (O_1494,N_18814,N_18651);
xnor UO_1495 (O_1495,N_18444,N_17189);
or UO_1496 (O_1496,N_19534,N_19382);
xor UO_1497 (O_1497,N_18607,N_19652);
xor UO_1498 (O_1498,N_18684,N_19710);
and UO_1499 (O_1499,N_18096,N_19249);
and UO_1500 (O_1500,N_19152,N_19897);
and UO_1501 (O_1501,N_17805,N_19860);
nand UO_1502 (O_1502,N_18884,N_17726);
and UO_1503 (O_1503,N_17393,N_17532);
xor UO_1504 (O_1504,N_17906,N_17512);
nor UO_1505 (O_1505,N_17867,N_19378);
and UO_1506 (O_1506,N_15997,N_17024);
nor UO_1507 (O_1507,N_19622,N_17629);
nor UO_1508 (O_1508,N_16594,N_17644);
nand UO_1509 (O_1509,N_18747,N_15528);
nand UO_1510 (O_1510,N_16967,N_18437);
nand UO_1511 (O_1511,N_19456,N_16213);
and UO_1512 (O_1512,N_19470,N_19091);
nor UO_1513 (O_1513,N_18710,N_16299);
and UO_1514 (O_1514,N_15995,N_19773);
nor UO_1515 (O_1515,N_16471,N_18528);
nor UO_1516 (O_1516,N_16000,N_18851);
nand UO_1517 (O_1517,N_18867,N_16349);
xor UO_1518 (O_1518,N_17859,N_19259);
and UO_1519 (O_1519,N_16822,N_18230);
xnor UO_1520 (O_1520,N_16362,N_18400);
nand UO_1521 (O_1521,N_15227,N_16426);
and UO_1522 (O_1522,N_16732,N_18522);
xnor UO_1523 (O_1523,N_15802,N_16621);
nand UO_1524 (O_1524,N_17295,N_17652);
nand UO_1525 (O_1525,N_19873,N_17627);
nor UO_1526 (O_1526,N_19764,N_19403);
nand UO_1527 (O_1527,N_16792,N_17164);
nand UO_1528 (O_1528,N_19794,N_19228);
nand UO_1529 (O_1529,N_15281,N_15191);
or UO_1530 (O_1530,N_18983,N_16547);
and UO_1531 (O_1531,N_16995,N_18488);
and UO_1532 (O_1532,N_18817,N_15866);
and UO_1533 (O_1533,N_16317,N_19039);
nand UO_1534 (O_1534,N_15046,N_16319);
and UO_1535 (O_1535,N_18629,N_19026);
nand UO_1536 (O_1536,N_15124,N_15241);
and UO_1537 (O_1537,N_16965,N_16806);
and UO_1538 (O_1538,N_19307,N_19312);
xor UO_1539 (O_1539,N_18806,N_17880);
xnor UO_1540 (O_1540,N_19314,N_16915);
or UO_1541 (O_1541,N_18869,N_18816);
nor UO_1542 (O_1542,N_15089,N_15828);
nand UO_1543 (O_1543,N_19355,N_19797);
xor UO_1544 (O_1544,N_17426,N_18420);
nor UO_1545 (O_1545,N_18000,N_18024);
nor UO_1546 (O_1546,N_17905,N_17072);
or UO_1547 (O_1547,N_17177,N_19554);
nor UO_1548 (O_1548,N_15002,N_17523);
xor UO_1549 (O_1549,N_16673,N_16860);
xnor UO_1550 (O_1550,N_15916,N_18204);
nand UO_1551 (O_1551,N_19653,N_17614);
and UO_1552 (O_1552,N_19828,N_17264);
nor UO_1553 (O_1553,N_16852,N_18719);
nor UO_1554 (O_1554,N_19596,N_17191);
and UO_1555 (O_1555,N_19901,N_15727);
nor UO_1556 (O_1556,N_16932,N_19236);
nand UO_1557 (O_1557,N_18778,N_18792);
nor UO_1558 (O_1558,N_16371,N_15394);
xnor UO_1559 (O_1559,N_15706,N_17585);
nand UO_1560 (O_1560,N_18260,N_18941);
or UO_1561 (O_1561,N_15380,N_19743);
nand UO_1562 (O_1562,N_16202,N_19603);
and UO_1563 (O_1563,N_16948,N_17448);
or UO_1564 (O_1564,N_18708,N_19106);
or UO_1565 (O_1565,N_16112,N_19630);
and UO_1566 (O_1566,N_18151,N_15602);
and UO_1567 (O_1567,N_16774,N_18784);
nor UO_1568 (O_1568,N_15711,N_19725);
xor UO_1569 (O_1569,N_17377,N_18549);
or UO_1570 (O_1570,N_18620,N_16840);
and UO_1571 (O_1571,N_18217,N_19459);
nand UO_1572 (O_1572,N_19729,N_17999);
or UO_1573 (O_1573,N_15685,N_17720);
nand UO_1574 (O_1574,N_15470,N_16761);
nand UO_1575 (O_1575,N_16538,N_16838);
nor UO_1576 (O_1576,N_15323,N_15752);
nand UO_1577 (O_1577,N_16449,N_16443);
or UO_1578 (O_1578,N_16809,N_16998);
nand UO_1579 (O_1579,N_19491,N_15908);
xor UO_1580 (O_1580,N_19814,N_15532);
or UO_1581 (O_1581,N_18871,N_17597);
nand UO_1582 (O_1582,N_16023,N_15481);
and UO_1583 (O_1583,N_18364,N_18346);
xor UO_1584 (O_1584,N_17939,N_15770);
nand UO_1585 (O_1585,N_19406,N_19308);
xnor UO_1586 (O_1586,N_16713,N_19126);
and UO_1587 (O_1587,N_18969,N_15148);
nor UO_1588 (O_1588,N_17787,N_16311);
xor UO_1589 (O_1589,N_15403,N_17685);
xor UO_1590 (O_1590,N_15670,N_15815);
nor UO_1591 (O_1591,N_16990,N_16465);
xnor UO_1592 (O_1592,N_18826,N_16724);
xor UO_1593 (O_1593,N_19224,N_19809);
nand UO_1594 (O_1594,N_17305,N_18534);
xor UO_1595 (O_1595,N_15291,N_19907);
or UO_1596 (O_1596,N_15092,N_17431);
or UO_1597 (O_1597,N_16671,N_17382);
or UO_1598 (O_1598,N_16265,N_16700);
or UO_1599 (O_1599,N_18998,N_17157);
and UO_1600 (O_1600,N_17187,N_18924);
nand UO_1601 (O_1601,N_17565,N_17032);
nor UO_1602 (O_1602,N_17673,N_19694);
nand UO_1603 (O_1603,N_17894,N_16618);
and UO_1604 (O_1604,N_18196,N_15263);
or UO_1605 (O_1605,N_17871,N_15493);
or UO_1606 (O_1606,N_17057,N_19370);
nor UO_1607 (O_1607,N_19197,N_16435);
or UO_1608 (O_1608,N_17243,N_17176);
or UO_1609 (O_1609,N_16540,N_18809);
xnor UO_1610 (O_1610,N_15564,N_18108);
and UO_1611 (O_1611,N_19151,N_18348);
nand UO_1612 (O_1612,N_18408,N_16968);
and UO_1613 (O_1613,N_16218,N_17135);
nor UO_1614 (O_1614,N_17776,N_19057);
nor UO_1615 (O_1615,N_18693,N_19018);
and UO_1616 (O_1616,N_15461,N_19970);
nor UO_1617 (O_1617,N_18738,N_17162);
xor UO_1618 (O_1618,N_18746,N_17314);
and UO_1619 (O_1619,N_17588,N_16518);
or UO_1620 (O_1620,N_15268,N_18590);
nand UO_1621 (O_1621,N_19175,N_19434);
nand UO_1622 (O_1622,N_18847,N_18606);
and UO_1623 (O_1623,N_17343,N_16715);
xor UO_1624 (O_1624,N_17564,N_15590);
and UO_1625 (O_1625,N_15574,N_15306);
or UO_1626 (O_1626,N_18779,N_16649);
nor UO_1627 (O_1627,N_17247,N_17645);
or UO_1628 (O_1628,N_16455,N_18799);
xnor UO_1629 (O_1629,N_17854,N_18653);
nand UO_1630 (O_1630,N_19661,N_15902);
xor UO_1631 (O_1631,N_19419,N_17780);
xor UO_1632 (O_1632,N_15474,N_16460);
nand UO_1633 (O_1633,N_18860,N_18295);
nor UO_1634 (O_1634,N_15631,N_16129);
nor UO_1635 (O_1635,N_16691,N_17113);
and UO_1636 (O_1636,N_15265,N_19082);
nand UO_1637 (O_1637,N_19005,N_16097);
nor UO_1638 (O_1638,N_18949,N_18729);
xnor UO_1639 (O_1639,N_15994,N_15731);
nand UO_1640 (O_1640,N_15056,N_15881);
nand UO_1641 (O_1641,N_15535,N_15025);
and UO_1642 (O_1642,N_15662,N_15044);
nand UO_1643 (O_1643,N_18045,N_19958);
nor UO_1644 (O_1644,N_16837,N_16357);
nor UO_1645 (O_1645,N_16905,N_16957);
nor UO_1646 (O_1646,N_17877,N_17408);
xnor UO_1647 (O_1647,N_19777,N_17813);
xnor UO_1648 (O_1648,N_15468,N_16993);
xor UO_1649 (O_1649,N_16808,N_16512);
or UO_1650 (O_1650,N_17898,N_18191);
nor UO_1651 (O_1651,N_16060,N_18845);
xnor UO_1652 (O_1652,N_16003,N_18597);
nand UO_1653 (O_1653,N_16545,N_19179);
nor UO_1654 (O_1654,N_15116,N_17624);
xnor UO_1655 (O_1655,N_17997,N_19500);
nor UO_1656 (O_1656,N_19349,N_19356);
nor UO_1657 (O_1657,N_18780,N_18129);
nor UO_1658 (O_1658,N_16579,N_16829);
or UO_1659 (O_1659,N_15759,N_15095);
or UO_1660 (O_1660,N_17206,N_15250);
or UO_1661 (O_1661,N_15523,N_16468);
xor UO_1662 (O_1662,N_15249,N_18082);
nand UO_1663 (O_1663,N_17998,N_18737);
and UO_1664 (O_1664,N_17407,N_18161);
nor UO_1665 (O_1665,N_17886,N_16149);
or UO_1666 (O_1666,N_18987,N_18248);
or UO_1667 (O_1667,N_17962,N_16820);
nor UO_1668 (O_1668,N_19714,N_18911);
xor UO_1669 (O_1669,N_15679,N_17158);
xnor UO_1670 (O_1670,N_16600,N_17075);
or UO_1671 (O_1671,N_18503,N_15346);
nand UO_1672 (O_1672,N_16306,N_15647);
nor UO_1673 (O_1673,N_16358,N_16108);
nand UO_1674 (O_1674,N_16762,N_15469);
xnor UO_1675 (O_1675,N_16926,N_16055);
and UO_1676 (O_1676,N_16480,N_19316);
xor UO_1677 (O_1677,N_18371,N_15983);
or UO_1678 (O_1678,N_15486,N_18777);
nand UO_1679 (O_1679,N_19977,N_15267);
nor UO_1680 (O_1680,N_19651,N_18398);
xnor UO_1681 (O_1681,N_15507,N_17556);
nand UO_1682 (O_1682,N_19199,N_19702);
xor UO_1683 (O_1683,N_16454,N_15484);
and UO_1684 (O_1684,N_18940,N_19142);
or UO_1685 (O_1685,N_16345,N_19424);
or UO_1686 (O_1686,N_16399,N_16165);
nor UO_1687 (O_1687,N_18478,N_19022);
xor UO_1688 (O_1688,N_15232,N_17519);
and UO_1689 (O_1689,N_15767,N_16220);
or UO_1690 (O_1690,N_17803,N_16756);
nor UO_1691 (O_1691,N_15425,N_19317);
nand UO_1692 (O_1692,N_15084,N_15712);
and UO_1693 (O_1693,N_19035,N_16007);
or UO_1694 (O_1694,N_15725,N_16758);
nand UO_1695 (O_1695,N_19062,N_17758);
and UO_1696 (O_1696,N_19485,N_16154);
nand UO_1697 (O_1697,N_18016,N_15006);
nor UO_1698 (O_1698,N_17583,N_16452);
or UO_1699 (O_1699,N_18042,N_15894);
and UO_1700 (O_1700,N_18272,N_16799);
nand UO_1701 (O_1701,N_18608,N_17513);
nor UO_1702 (O_1702,N_17908,N_19273);
xnor UO_1703 (O_1703,N_19529,N_15882);
xnor UO_1704 (O_1704,N_19492,N_18243);
and UO_1705 (O_1705,N_19056,N_17429);
or UO_1706 (O_1706,N_17625,N_17151);
xnor UO_1707 (O_1707,N_15640,N_16870);
or UO_1708 (O_1708,N_16871,N_19750);
nor UO_1709 (O_1709,N_17476,N_15355);
nand UO_1710 (O_1710,N_15074,N_18040);
and UO_1711 (O_1711,N_18315,N_18713);
xnor UO_1712 (O_1712,N_16230,N_16316);
nor UO_1713 (O_1713,N_16558,N_18855);
and UO_1714 (O_1714,N_16610,N_15149);
xor UO_1715 (O_1715,N_16899,N_16730);
nand UO_1716 (O_1716,N_15592,N_18279);
xnor UO_1717 (O_1717,N_19034,N_17196);
or UO_1718 (O_1718,N_18919,N_19497);
xnor UO_1719 (O_1719,N_17035,N_17782);
or UO_1720 (O_1720,N_18060,N_18077);
xnor UO_1721 (O_1721,N_18825,N_17887);
and UO_1722 (O_1722,N_17292,N_18592);
xor UO_1723 (O_1723,N_15653,N_19759);
or UO_1724 (O_1724,N_15756,N_18080);
nand UO_1725 (O_1725,N_17938,N_17353);
nand UO_1726 (O_1726,N_19639,N_15429);
nor UO_1727 (O_1727,N_15933,N_19527);
xnor UO_1728 (O_1728,N_17643,N_18113);
nand UO_1729 (O_1729,N_16197,N_15999);
or UO_1730 (O_1730,N_16936,N_15957);
nor UO_1731 (O_1731,N_19903,N_16205);
nor UO_1732 (O_1732,N_19390,N_16143);
nor UO_1733 (O_1733,N_17293,N_16577);
nand UO_1734 (O_1734,N_15408,N_16825);
or UO_1735 (O_1735,N_16090,N_19864);
or UO_1736 (O_1736,N_16591,N_15327);
or UO_1737 (O_1737,N_15536,N_18665);
or UO_1738 (O_1738,N_16727,N_15330);
or UO_1739 (O_1739,N_19003,N_19550);
or UO_1740 (O_1740,N_15829,N_19335);
and UO_1741 (O_1741,N_15940,N_18072);
nand UO_1742 (O_1742,N_16759,N_19385);
nand UO_1743 (O_1743,N_19637,N_16437);
nor UO_1744 (O_1744,N_18410,N_17022);
and UO_1745 (O_1745,N_16398,N_15573);
and UO_1746 (O_1746,N_15114,N_15554);
nand UO_1747 (O_1747,N_15898,N_19431);
nand UO_1748 (O_1748,N_15713,N_16933);
and UO_1749 (O_1749,N_19292,N_17045);
nor UO_1750 (O_1750,N_16162,N_19186);
nand UO_1751 (O_1751,N_16059,N_17203);
or UO_1752 (O_1752,N_18436,N_15651);
xor UO_1753 (O_1753,N_18238,N_19654);
and UO_1754 (O_1754,N_17487,N_19480);
or UO_1755 (O_1755,N_19922,N_16147);
nor UO_1756 (O_1756,N_15811,N_19009);
nand UO_1757 (O_1757,N_19484,N_17688);
nand UO_1758 (O_1758,N_18340,N_18223);
or UO_1759 (O_1759,N_17118,N_15103);
or UO_1760 (O_1760,N_17913,N_16380);
nor UO_1761 (O_1761,N_18120,N_19066);
or UO_1762 (O_1762,N_18412,N_16025);
xnor UO_1763 (O_1763,N_19711,N_19734);
and UO_1764 (O_1764,N_15684,N_17929);
or UO_1765 (O_1765,N_18210,N_16241);
nand UO_1766 (O_1766,N_15958,N_17098);
or UO_1767 (O_1767,N_15048,N_19786);
or UO_1768 (O_1768,N_18577,N_19735);
and UO_1769 (O_1769,N_17114,N_16019);
xnor UO_1770 (O_1770,N_16866,N_17048);
or UO_1771 (O_1771,N_19727,N_19760);
nor UO_1772 (O_1772,N_15158,N_15910);
and UO_1773 (O_1773,N_18765,N_18955);
xnor UO_1774 (O_1774,N_16681,N_16181);
nor UO_1775 (O_1775,N_18365,N_19240);
nor UO_1776 (O_1776,N_19027,N_17422);
nand UO_1777 (O_1777,N_15989,N_19787);
xor UO_1778 (O_1778,N_15195,N_19526);
nand UO_1779 (O_1779,N_15801,N_17889);
nor UO_1780 (O_1780,N_17824,N_16033);
nand UO_1781 (O_1781,N_18868,N_19448);
nand UO_1782 (O_1782,N_17900,N_15499);
nor UO_1783 (O_1783,N_19241,N_19275);
nand UO_1784 (O_1784,N_18694,N_17903);
nand UO_1785 (O_1785,N_19994,N_17868);
xor UO_1786 (O_1786,N_17413,N_16777);
xor UO_1787 (O_1787,N_17235,N_17772);
and UO_1788 (O_1788,N_16141,N_18676);
xnor UO_1789 (O_1789,N_18980,N_19564);
nor UO_1790 (O_1790,N_15053,N_16816);
nor UO_1791 (O_1791,N_18022,N_17919);
or UO_1792 (O_1792,N_19572,N_15293);
or UO_1793 (O_1793,N_17714,N_19788);
nor UO_1794 (O_1794,N_17912,N_16562);
or UO_1795 (O_1795,N_19991,N_19682);
or UO_1796 (O_1796,N_17922,N_17602);
and UO_1797 (O_1797,N_17899,N_18762);
xor UO_1798 (O_1798,N_17947,N_18928);
nor UO_1799 (O_1799,N_19854,N_19265);
and UO_1800 (O_1800,N_15754,N_16098);
and UO_1801 (O_1801,N_15529,N_15218);
or UO_1802 (O_1802,N_19551,N_19002);
or UO_1803 (O_1803,N_17464,N_15753);
and UO_1804 (O_1804,N_19618,N_17840);
and UO_1805 (O_1805,N_15724,N_17651);
nand UO_1806 (O_1806,N_17537,N_19997);
or UO_1807 (O_1807,N_16038,N_19257);
nand UO_1808 (O_1808,N_16790,N_15973);
nor UO_1809 (O_1809,N_17415,N_17323);
and UO_1810 (O_1810,N_17661,N_16647);
nor UO_1811 (O_1811,N_17893,N_16773);
nand UO_1812 (O_1812,N_16210,N_15212);
nor UO_1813 (O_1813,N_17058,N_19073);
nand UO_1814 (O_1814,N_18194,N_19829);
nor UO_1815 (O_1815,N_17982,N_15360);
xnor UO_1816 (O_1816,N_17279,N_15637);
xnor UO_1817 (O_1817,N_18199,N_18181);
or UO_1818 (O_1818,N_16552,N_16749);
nand UO_1819 (O_1819,N_18443,N_15885);
or UO_1820 (O_1820,N_19754,N_17105);
nor UO_1821 (O_1821,N_16360,N_17527);
nor UO_1822 (O_1822,N_16363,N_15287);
xor UO_1823 (O_1823,N_16521,N_15645);
and UO_1824 (O_1824,N_17866,N_15935);
xnor UO_1825 (O_1825,N_15247,N_18766);
and UO_1826 (O_1826,N_19999,N_18311);
or UO_1827 (O_1827,N_19663,N_19569);
and UO_1828 (O_1828,N_18819,N_18923);
xor UO_1829 (O_1829,N_18822,N_16015);
nor UO_1830 (O_1830,N_18764,N_19340);
nor UO_1831 (O_1831,N_18079,N_19696);
and UO_1832 (O_1832,N_19872,N_18205);
nand UO_1833 (O_1833,N_19352,N_18880);
xnor UO_1834 (O_1834,N_19498,N_17718);
or UO_1835 (O_1835,N_15356,N_19747);
nand UO_1836 (O_1836,N_18783,N_16791);
xnor UO_1837 (O_1837,N_16934,N_15401);
or UO_1838 (O_1838,N_16497,N_16227);
nand UO_1839 (O_1839,N_15929,N_16945);
or UO_1840 (O_1840,N_15663,N_17149);
nand UO_1841 (O_1841,N_18907,N_15897);
nand UO_1842 (O_1842,N_18537,N_17359);
nand UO_1843 (O_1843,N_18499,N_18947);
or UO_1844 (O_1844,N_18136,N_16705);
and UO_1845 (O_1845,N_19646,N_15919);
or UO_1846 (O_1846,N_19161,N_15780);
nand UO_1847 (O_1847,N_17818,N_17318);
nor UO_1848 (O_1848,N_16940,N_17637);
nor UO_1849 (O_1849,N_15521,N_18757);
and UO_1850 (O_1850,N_17379,N_15608);
nor UO_1851 (O_1851,N_19464,N_15361);
and UO_1852 (O_1852,N_17933,N_15201);
or UO_1853 (O_1853,N_15180,N_17492);
xnor UO_1854 (O_1854,N_18789,N_16699);
nand UO_1855 (O_1855,N_18116,N_18874);
nand UO_1856 (O_1856,N_17280,N_18401);
xnor UO_1857 (O_1857,N_17026,N_15096);
nand UO_1858 (O_1858,N_15912,N_15351);
nand UO_1859 (O_1859,N_19929,N_15580);
nand UO_1860 (O_1860,N_19001,N_18350);
xnor UO_1861 (O_1861,N_17774,N_19538);
or UO_1862 (O_1862,N_16847,N_18273);
xnor UO_1863 (O_1863,N_19233,N_17554);
nor UO_1864 (O_1864,N_15131,N_19493);
xor UO_1865 (O_1865,N_15451,N_17208);
nand UO_1866 (O_1866,N_17443,N_16911);
nand UO_1867 (O_1867,N_17558,N_15196);
or UO_1868 (O_1868,N_15846,N_19517);
nor UO_1869 (O_1869,N_19117,N_18121);
xor UO_1870 (O_1870,N_18885,N_17875);
or UO_1871 (O_1871,N_16517,N_18699);
and UO_1872 (O_1872,N_17756,N_17439);
or UO_1873 (O_1873,N_19415,N_19948);
or UO_1874 (O_1874,N_16446,N_19277);
and UO_1875 (O_1875,N_16789,N_19568);
xnor UO_1876 (O_1876,N_15336,N_19208);
xnor UO_1877 (O_1877,N_17567,N_18573);
nand UO_1878 (O_1878,N_19090,N_18015);
xnor UO_1879 (O_1879,N_19543,N_15589);
xor UO_1880 (O_1880,N_17120,N_15167);
nor UO_1881 (O_1881,N_19700,N_18951);
and UO_1882 (O_1882,N_15570,N_19008);
or UO_1883 (O_1883,N_19895,N_17618);
and UO_1884 (O_1884,N_19463,N_15297);
xnor UO_1885 (O_1885,N_18525,N_16438);
nor UO_1886 (O_1886,N_15214,N_15152);
and UO_1887 (O_1887,N_16553,N_16775);
xnor UO_1888 (O_1888,N_18547,N_18759);
nand UO_1889 (O_1889,N_15452,N_15334);
and UO_1890 (O_1890,N_19871,N_18671);
nor UO_1891 (O_1891,N_19364,N_17010);
nand UO_1892 (O_1892,N_19465,N_18495);
nor UO_1893 (O_1893,N_16873,N_18202);
and UO_1894 (O_1894,N_18498,N_17219);
xnor UO_1895 (O_1895,N_15769,N_16295);
and UO_1896 (O_1896,N_17683,N_15258);
xor UO_1897 (O_1897,N_16094,N_18130);
nand UO_1898 (O_1898,N_17376,N_15170);
and UO_1899 (O_1899,N_19042,N_17657);
nor UO_1900 (O_1900,N_18856,N_15635);
nand UO_1901 (O_1901,N_15878,N_19940);
and UO_1902 (O_1902,N_18664,N_18545);
and UO_1903 (O_1903,N_15641,N_18142);
xor UO_1904 (O_1904,N_19655,N_19260);
nand UO_1905 (O_1905,N_18908,N_19291);
nand UO_1906 (O_1906,N_16107,N_15768);
or UO_1907 (O_1907,N_17458,N_19063);
nand UO_1908 (O_1908,N_18207,N_19752);
nand UO_1909 (O_1909,N_15270,N_16951);
xnor UO_1910 (O_1910,N_19745,N_15412);
and UO_1911 (O_1911,N_18703,N_18214);
and UO_1912 (O_1912,N_17259,N_16603);
or UO_1913 (O_1913,N_18972,N_17029);
nor UO_1914 (O_1914,N_15337,N_16011);
or UO_1915 (O_1915,N_18807,N_17784);
nand UO_1916 (O_1916,N_17814,N_15009);
nor UO_1917 (O_1917,N_17613,N_17538);
or UO_1918 (O_1918,N_19183,N_16539);
nor UO_1919 (O_1919,N_15924,N_15682);
xor UO_1920 (O_1920,N_17792,N_16110);
xnor UO_1921 (O_1921,N_15042,N_18467);
or UO_1922 (O_1922,N_18635,N_17126);
nor UO_1923 (O_1923,N_16329,N_19635);
xor UO_1924 (O_1924,N_17755,N_15823);
xor UO_1925 (O_1925,N_18730,N_17300);
xor UO_1926 (O_1926,N_18973,N_15234);
xnor UO_1927 (O_1927,N_15436,N_16632);
nand UO_1928 (O_1928,N_16723,N_15845);
nand UO_1929 (O_1929,N_15302,N_15859);
and UO_1930 (O_1930,N_19294,N_17399);
and UO_1931 (O_1931,N_17337,N_19761);
xnor UO_1932 (O_1932,N_17819,N_18870);
and UO_1933 (O_1933,N_15365,N_19396);
nand UO_1934 (O_1934,N_17388,N_18917);
or UO_1935 (O_1935,N_19032,N_15600);
and UO_1936 (O_1936,N_15776,N_15719);
xnor UO_1937 (O_1937,N_15211,N_18758);
and UO_1938 (O_1938,N_16268,N_18728);
and UO_1939 (O_1939,N_15722,N_15001);
or UO_1940 (O_1940,N_19173,N_17136);
or UO_1941 (O_1941,N_15226,N_16776);
xor UO_1942 (O_1942,N_15831,N_16548);
nor UO_1943 (O_1943,N_17341,N_16017);
xor UO_1944 (O_1944,N_19793,N_16291);
or UO_1945 (O_1945,N_15586,N_19402);
nor UO_1946 (O_1946,N_17514,N_15125);
or UO_1947 (O_1947,N_17317,N_15959);
nor UO_1948 (O_1948,N_15045,N_16440);
nand UO_1949 (O_1949,N_17660,N_16477);
and UO_1950 (O_1950,N_17421,N_18569);
nor UO_1951 (O_1951,N_19973,N_16395);
or UO_1952 (O_1952,N_15694,N_17419);
or UO_1953 (O_1953,N_18506,N_16640);
nor UO_1954 (O_1954,N_16987,N_17389);
nand UO_1955 (O_1955,N_16516,N_16479);
or UO_1956 (O_1956,N_15733,N_18038);
nand UO_1957 (O_1957,N_16886,N_16495);
xor UO_1958 (O_1958,N_17427,N_15794);
nand UO_1959 (O_1959,N_18068,N_16032);
nand UO_1960 (O_1960,N_15021,N_16974);
nand UO_1961 (O_1961,N_15017,N_17209);
or UO_1962 (O_1962,N_19038,N_18387);
xnor UO_1963 (O_1963,N_16482,N_15215);
nand UO_1964 (O_1964,N_17858,N_17738);
nor UO_1965 (O_1965,N_16170,N_16629);
nand UO_1966 (O_1966,N_16392,N_19476);
nor UO_1967 (O_1967,N_17520,N_16374);
nor UO_1968 (O_1968,N_19128,N_18649);
or UO_1969 (O_1969,N_16983,N_18901);
nor UO_1970 (O_1970,N_18835,N_15510);
or UO_1971 (O_1971,N_18291,N_18252);
or UO_1972 (O_1972,N_16958,N_16300);
nor UO_1973 (O_1973,N_15699,N_15864);
xor UO_1974 (O_1974,N_15549,N_15597);
nor UO_1975 (O_1975,N_15613,N_16427);
nand UO_1976 (O_1976,N_17658,N_19326);
nand UO_1977 (O_1977,N_18553,N_17484);
xnor UO_1978 (O_1978,N_17904,N_17239);
nor UO_1979 (O_1979,N_17795,N_15402);
and UO_1980 (O_1980,N_17246,N_18878);
nand UO_1981 (O_1981,N_15693,N_17169);
nand UO_1982 (O_1982,N_15838,N_16123);
nor UO_1983 (O_1983,N_16463,N_18376);
nand UO_1984 (O_1984,N_15040,N_17117);
nand UO_1985 (O_1985,N_16944,N_17670);
and UO_1986 (O_1986,N_18841,N_15557);
and UO_1987 (O_1987,N_18298,N_17557);
nor UO_1988 (O_1988,N_19219,N_16166);
nor UO_1989 (O_1989,N_15555,N_18203);
and UO_1990 (O_1990,N_19511,N_19827);
and UO_1991 (O_1991,N_16456,N_16373);
nand UO_1992 (O_1992,N_18872,N_19135);
or UO_1993 (O_1993,N_17920,N_16182);
nand UO_1994 (O_1994,N_17687,N_18104);
nor UO_1995 (O_1995,N_16800,N_18918);
nor UO_1996 (O_1996,N_19141,N_17547);
nand UO_1997 (O_1997,N_16677,N_19268);
or UO_1998 (O_1998,N_18760,N_15797);
xnor UO_1999 (O_1999,N_15023,N_16052);
xor UO_2000 (O_2000,N_18356,N_16318);
or UO_2001 (O_2001,N_19262,N_19242);
nor UO_2002 (O_2002,N_19029,N_15034);
nor UO_2003 (O_2003,N_15950,N_16588);
nor UO_2004 (O_2004,N_17983,N_18454);
xnor UO_2005 (O_2005,N_15354,N_15840);
and UO_2006 (O_2006,N_18380,N_16778);
nand UO_2007 (O_2007,N_16685,N_17634);
nand UO_2008 (O_2008,N_17108,N_19851);
nor UO_2009 (O_2009,N_18920,N_17578);
or UO_2010 (O_2010,N_17284,N_15869);
or UO_2011 (O_2011,N_17043,N_15576);
and UO_2012 (O_2012,N_15932,N_17386);
and UO_2013 (O_2013,N_15295,N_15782);
and UO_2014 (O_2014,N_17362,N_19609);
nand UO_2015 (O_2015,N_17256,N_19881);
nand UO_2016 (O_2016,N_17180,N_18025);
nand UO_2017 (O_2017,N_18469,N_17340);
and UO_2018 (O_2018,N_16135,N_18570);
xor UO_2019 (O_2019,N_15558,N_17488);
nor UO_2020 (O_2020,N_16103,N_19857);
xor UO_2021 (O_2021,N_16207,N_16641);
and UO_2022 (O_2022,N_16884,N_16006);
nor UO_2023 (O_2023,N_18752,N_15145);
and UO_2024 (O_2024,N_17830,N_18638);
nand UO_2025 (O_2025,N_16209,N_19420);
nor UO_2026 (O_2026,N_17616,N_15762);
or UO_2027 (O_2027,N_18743,N_16281);
xor UO_2028 (O_2028,N_17216,N_18605);
nor UO_2029 (O_2029,N_15162,N_15313);
nand UO_2030 (O_2030,N_15569,N_19499);
nand UO_2031 (O_2031,N_17534,N_19457);
nand UO_2032 (O_2032,N_17853,N_15596);
or UO_2033 (O_2033,N_16350,N_17463);
and UO_2034 (O_2034,N_15700,N_15943);
nand UO_2035 (O_2035,N_15572,N_19200);
nor UO_2036 (O_2036,N_16508,N_18697);
nand UO_2037 (O_2037,N_18997,N_19708);
and UO_2038 (O_2038,N_19634,N_16304);
or UO_2039 (O_2039,N_17138,N_19601);
or UO_2040 (O_2040,N_17266,N_15890);
nand UO_2041 (O_2041,N_19731,N_16199);
xor UO_2042 (O_2042,N_19816,N_19139);
or UO_2043 (O_2043,N_18600,N_15358);
and UO_2044 (O_2044,N_18681,N_16257);
and UO_2045 (O_2045,N_16275,N_17570);
nor UO_2046 (O_2046,N_16396,N_18976);
nor UO_2047 (O_2047,N_18689,N_19781);
nor UO_2048 (O_2048,N_18218,N_19166);
nor UO_2049 (O_2049,N_19528,N_19740);
nor UO_2050 (O_2050,N_17004,N_18051);
or UO_2051 (O_2051,N_19077,N_18934);
nand UO_2052 (O_2052,N_18193,N_17902);
xnor UO_2053 (O_2053,N_18750,N_17628);
nor UO_2054 (O_2054,N_16757,N_18519);
nand UO_2055 (O_2055,N_15612,N_15153);
xor UO_2056 (O_2056,N_15678,N_19037);
and UO_2057 (O_2057,N_19565,N_18714);
nor UO_2058 (O_2058,N_19945,N_15553);
nor UO_2059 (O_2059,N_17930,N_17641);
and UO_2060 (O_2060,N_18666,N_17474);
nand UO_2061 (O_2061,N_19887,N_18431);
and UO_2062 (O_2062,N_17832,N_19713);
or UO_2063 (O_2063,N_18381,N_16260);
nor UO_2064 (O_2064,N_19585,N_16324);
nand UO_2065 (O_2065,N_15672,N_16212);
nor UO_2066 (O_2066,N_15516,N_15244);
or UO_2067 (O_2067,N_17019,N_17229);
nand UO_2068 (O_2068,N_17716,N_17926);
and UO_2069 (O_2069,N_18978,N_17198);
or UO_2070 (O_2070,N_18216,N_19744);
nand UO_2071 (O_2071,N_15259,N_18712);
nor UO_2072 (O_2072,N_18414,N_16321);
or UO_2073 (O_2073,N_19020,N_15015);
nor UO_2074 (O_2074,N_15253,N_17928);
or UO_2075 (O_2075,N_19966,N_15761);
nor UO_2076 (O_2076,N_15014,N_19983);
or UO_2077 (O_2077,N_15786,N_19959);
nand UO_2078 (O_2078,N_19570,N_15310);
nor UO_2079 (O_2079,N_19845,N_17631);
nand UO_2080 (O_2080,N_18385,N_15984);
xor UO_2081 (O_2081,N_15031,N_17799);
nor UO_2082 (O_2082,N_15062,N_19111);
or UO_2083 (O_2083,N_16554,N_16892);
and UO_2084 (O_2084,N_16906,N_15160);
nand UO_2085 (O_2085,N_19450,N_16960);
nor UO_2086 (O_2086,N_17244,N_16784);
or UO_2087 (O_2087,N_18497,N_17372);
nand UO_2088 (O_2088,N_16783,N_15423);
xnor UO_2089 (O_2089,N_15584,N_16689);
nand UO_2090 (O_2090,N_16566,N_15428);
nand UO_2091 (O_2091,N_17793,N_17810);
or UO_2092 (O_2092,N_18182,N_18844);
nor UO_2093 (O_2093,N_16894,N_15272);
xor UO_2094 (O_2094,N_16543,N_17170);
nand UO_2095 (O_2095,N_17522,N_17143);
and UO_2096 (O_2096,N_16469,N_17591);
xnor UO_2097 (O_2097,N_16823,N_17589);
and UO_2098 (O_2098,N_17729,N_19648);
xor UO_2099 (O_2099,N_19861,N_17217);
nand UO_2100 (O_2100,N_18167,N_19157);
xor UO_2101 (O_2101,N_19628,N_16528);
xor UO_2102 (O_2102,N_15836,N_16964);
xnor UO_2103 (O_2103,N_16409,N_19832);
nand UO_2104 (O_2104,N_16605,N_18740);
nor UO_2105 (O_2105,N_16525,N_18984);
nand UO_2106 (O_2106,N_18539,N_17299);
xor UO_2107 (O_2107,N_19995,N_19280);
and UO_2108 (O_2108,N_18316,N_17901);
and UO_2109 (O_2109,N_15489,N_19096);
nand UO_2110 (O_2110,N_17452,N_16343);
and UO_2111 (O_2111,N_16302,N_18014);
and UO_2112 (O_2112,N_18160,N_16327);
xor UO_2113 (O_2113,N_15819,N_19384);
nand UO_2114 (O_2114,N_16608,N_19014);
nor UO_2115 (O_2115,N_17617,N_17369);
or UO_2116 (O_2116,N_19883,N_15677);
or UO_2117 (O_2117,N_17364,N_18709);
nand UO_2118 (O_2118,N_19798,N_17584);
or UO_2119 (O_2119,N_18074,N_15715);
nor UO_2120 (O_2120,N_16802,N_19417);
nand UO_2121 (O_2121,N_16867,N_17884);
nand UO_2122 (O_2122,N_17441,N_16755);
nand UO_2123 (O_2123,N_19315,N_17477);
or UO_2124 (O_2124,N_19454,N_17961);
nand UO_2125 (O_2125,N_19507,N_15666);
xor UO_2126 (O_2126,N_17507,N_16994);
and UO_2127 (O_2127,N_17071,N_18384);
and UO_2128 (O_2128,N_17012,N_18944);
nor UO_2129 (O_2129,N_17085,N_16563);
xnor UO_2130 (O_2130,N_19865,N_19896);
nand UO_2131 (O_2131,N_16339,N_16615);
nand UO_2132 (O_2132,N_17449,N_18455);
and UO_2133 (O_2133,N_18149,N_17530);
xnor UO_2134 (O_2134,N_16491,N_17839);
nand UO_2135 (O_2135,N_16982,N_16217);
and UO_2136 (O_2136,N_15644,N_16172);
xnor UO_2137 (O_2137,N_17283,N_15575);
nand UO_2138 (O_2138,N_17721,N_17457);
and UO_2139 (O_2139,N_17692,N_19912);
nor UO_2140 (O_2140,N_19004,N_19443);
nor UO_2141 (O_2141,N_19455,N_16638);
or UO_2142 (O_2142,N_19071,N_19159);
nor UO_2143 (O_2143,N_19946,N_19557);
xor UO_2144 (O_2144,N_19625,N_19423);
or UO_2145 (O_2145,N_19578,N_19313);
nand UO_2146 (O_2146,N_19049,N_15277);
xnor UO_2147 (O_2147,N_17338,N_16970);
or UO_2148 (O_2148,N_19325,N_16018);
nor UO_2149 (O_2149,N_19726,N_15135);
nand UO_2150 (O_2150,N_18434,N_19192);
xnor UO_2151 (O_2151,N_19065,N_15294);
nand UO_2152 (O_2152,N_16383,N_16670);
and UO_2153 (O_2153,N_17000,N_16136);
nand UO_2154 (O_2154,N_17038,N_16550);
or UO_2155 (O_2155,N_18456,N_15032);
xor UO_2156 (O_2156,N_17678,N_19220);
xor UO_2157 (O_2157,N_18512,N_16040);
xnor UO_2158 (O_2158,N_16215,N_17812);
nand UO_2159 (O_2159,N_15676,N_17829);
and UO_2160 (O_2160,N_17319,N_16901);
and UO_2161 (O_2161,N_15751,N_18614);
nand UO_2162 (O_2162,N_17200,N_17308);
or UO_2163 (O_2163,N_18438,N_17163);
and UO_2164 (O_2164,N_18812,N_15003);
and UO_2165 (O_2165,N_16718,N_15952);
or UO_2166 (O_2166,N_19636,N_19971);
or UO_2167 (O_2167,N_15654,N_18717);
nand UO_2168 (O_2168,N_16660,N_16204);
nor UO_2169 (O_2169,N_16259,N_18968);
nor UO_2170 (O_2170,N_18333,N_17332);
xnor UO_2171 (O_2171,N_19120,N_17310);
nor UO_2172 (O_2172,N_16541,N_17270);
nor UO_2173 (O_2173,N_17316,N_15809);
xor UO_2174 (O_2174,N_17053,N_18776);
nor UO_2175 (O_2175,N_16568,N_18858);
nor UO_2176 (O_2176,N_17479,N_18556);
or UO_2177 (O_2177,N_15968,N_19248);
nor UO_2178 (O_2178,N_16646,N_15852);
and UO_2179 (O_2179,N_17580,N_19667);
and UO_2180 (O_2180,N_17367,N_17178);
nand UO_2181 (O_2181,N_15702,N_15717);
or UO_2182 (O_2182,N_18502,N_17693);
xor UO_2183 (O_2183,N_17456,N_15305);
nand UO_2184 (O_2184,N_17204,N_18145);
xnor UO_2185 (O_2185,N_18633,N_16130);
xnor UO_2186 (O_2186,N_19644,N_17290);
and UO_2187 (O_2187,N_19980,N_18300);
nor UO_2188 (O_2188,N_15518,N_19079);
xnor UO_2189 (O_2189,N_19150,N_15708);
xnor UO_2190 (O_2190,N_16476,N_16447);
nor UO_2191 (O_2191,N_15210,N_15656);
nand UO_2192 (O_2192,N_18345,N_16326);
xnor UO_2193 (O_2193,N_18881,N_15186);
xnor UO_2194 (O_2194,N_19134,N_18994);
nand UO_2195 (O_2195,N_15739,N_16293);
or UO_2196 (O_2196,N_15290,N_19238);
nand UO_2197 (O_2197,N_18716,N_19365);
xor UO_2198 (O_2198,N_16061,N_17397);
and UO_2199 (O_2199,N_15764,N_16489);
nand UO_2200 (O_2200,N_15054,N_18622);
nand UO_2201 (O_2201,N_17542,N_18091);
xor UO_2202 (O_2202,N_15341,N_15113);
xnor UO_2203 (O_2203,N_17490,N_16731);
or UO_2204 (O_2204,N_19053,N_18221);
and UO_2205 (O_2205,N_19374,N_19919);
nand UO_2206 (O_2206,N_18843,N_18961);
nand UO_2207 (O_2207,N_19398,N_19889);
and UO_2208 (O_2208,N_18937,N_19351);
nor UO_2209 (O_2209,N_19342,N_18798);
nor UO_2210 (O_2210,N_16270,N_19605);
and UO_2211 (O_2211,N_19449,N_17099);
xnor UO_2212 (O_2212,N_17090,N_19762);
nor UO_2213 (O_2213,N_18465,N_17847);
nand UO_2214 (O_2214,N_19928,N_15659);
nor UO_2215 (O_2215,N_19923,N_16372);
or UO_2216 (O_2216,N_15066,N_18452);
nor UO_2217 (O_2217,N_19109,N_15714);
or UO_2218 (O_2218,N_17653,N_16254);
or UO_2219 (O_2219,N_16942,N_15646);
xor UO_2220 (O_2220,N_15627,N_18830);
and UO_2221 (O_2221,N_19254,N_19986);
xnor UO_2222 (O_2222,N_18459,N_19926);
or UO_2223 (O_2223,N_16609,N_17826);
and UO_2224 (O_2224,N_18422,N_15443);
or UO_2225 (O_2225,N_16827,N_19144);
or UO_2226 (O_2226,N_19626,N_16835);
nand UO_2227 (O_2227,N_19671,N_16614);
xnor UO_2228 (O_2228,N_16203,N_18411);
nand UO_2229 (O_2229,N_19638,N_17603);
nor UO_2230 (O_2230,N_16971,N_16286);
nor UO_2231 (O_2231,N_18429,N_19044);
xor UO_2232 (O_2232,N_15632,N_19580);
xor UO_2233 (O_2233,N_17992,N_19939);
and UO_2234 (O_2234,N_17713,N_16644);
nand UO_2235 (O_2235,N_18318,N_16485);
nor UO_2236 (O_2236,N_18690,N_19046);
nand UO_2237 (O_2237,N_15198,N_16590);
nor UO_2238 (O_2238,N_17737,N_16509);
and UO_2239 (O_2239,N_17327,N_15174);
and UO_2240 (O_2240,N_18891,N_18256);
or UO_2241 (O_2241,N_18591,N_19908);
or UO_2242 (O_2242,N_18439,N_18866);
xnor UO_2243 (O_2243,N_19566,N_16021);
nor UO_2244 (O_2244,N_16920,N_16897);
nor UO_2245 (O_2245,N_19624,N_16804);
and UO_2246 (O_2246,N_15251,N_16848);
and UO_2247 (O_2247,N_16070,N_15061);
nor UO_2248 (O_2248,N_15563,N_15384);
and UO_2249 (O_2249,N_17775,N_19849);
xor UO_2250 (O_2250,N_19321,N_15322);
and UO_2251 (O_2251,N_16022,N_18301);
or UO_2252 (O_2252,N_17594,N_19775);
nand UO_2253 (O_2253,N_15953,N_15982);
or UO_2254 (O_2254,N_17297,N_16661);
or UO_2255 (O_2255,N_18463,N_16194);
nand UO_2256 (O_2256,N_17703,N_18029);
xor UO_2257 (O_2257,N_15407,N_19792);
and UO_2258 (O_2258,N_15320,N_17861);
nor UO_2259 (O_2259,N_19812,N_16814);
nand UO_2260 (O_2260,N_19393,N_15043);
nor UO_2261 (O_2261,N_16955,N_16499);
xnor UO_2262 (O_2262,N_18692,N_16738);
xor UO_2263 (O_2263,N_17882,N_18836);
nand UO_2264 (O_2264,N_18652,N_15286);
nor UO_2265 (O_2265,N_19391,N_16619);
xnor UO_2266 (O_2266,N_15099,N_17582);
nor UO_2267 (O_2267,N_18109,N_18887);
xnor UO_2268 (O_2268,N_16187,N_18507);
xnor UO_2269 (O_2269,N_18157,N_19917);
or UO_2270 (O_2270,N_15128,N_16494);
nor UO_2271 (O_2271,N_15673,N_17820);
or UO_2272 (O_2272,N_19953,N_15069);
and UO_2273 (O_2273,N_18111,N_16169);
xor UO_2274 (O_2274,N_19649,N_17491);
xor UO_2275 (O_2275,N_19656,N_19616);
xnor UO_2276 (O_2276,N_16144,N_17798);
and UO_2277 (O_2277,N_15697,N_16530);
nand UO_2278 (O_2278,N_16049,N_16167);
nand UO_2279 (O_2279,N_17423,N_17258);
and UO_2280 (O_2280,N_18170,N_19198);
and UO_2281 (O_2281,N_15817,N_19676);
xor UO_2282 (O_2282,N_16150,N_15615);
and UO_2283 (O_2283,N_17970,N_15138);
nor UO_2284 (O_2284,N_18473,N_16839);
or UO_2285 (O_2285,N_17944,N_19433);
or UO_2286 (O_2286,N_18668,N_15130);
and UO_2287 (O_2287,N_15010,N_19295);
and UO_2288 (O_2288,N_18821,N_16930);
nor UO_2289 (O_2289,N_19989,N_18915);
nand UO_2290 (O_2290,N_18576,N_19246);
nand UO_2291 (O_2291,N_19988,N_15498);
or UO_2292 (O_2292,N_15948,N_19508);
or UO_2293 (O_2293,N_16653,N_17700);
or UO_2294 (O_2294,N_15141,N_19629);
nor UO_2295 (O_2295,N_16978,N_16604);
nor UO_2296 (O_2296,N_16602,N_15067);
or UO_2297 (O_2297,N_17025,N_16895);
nor UO_2298 (O_2298,N_19755,N_18270);
xnor UO_2299 (O_2299,N_17172,N_16334);
nor UO_2300 (O_2300,N_15221,N_18793);
or UO_2301 (O_2301,N_17777,N_17856);
or UO_2302 (O_2302,N_19045,N_16056);
or UO_2303 (O_2303,N_19237,N_16039);
or UO_2304 (O_2304,N_18208,N_17937);
or UO_2305 (O_2305,N_17161,N_16687);
or UO_2306 (O_2306,N_19604,N_18239);
and UO_2307 (O_2307,N_15278,N_18399);
nor UO_2308 (O_2308,N_19808,N_17909);
nand UO_2309 (O_2309,N_18241,N_19950);
nor UO_2310 (O_2310,N_19031,N_16992);
or UO_2311 (O_2311,N_16627,N_17001);
nand UO_2312 (O_2312,N_18375,N_17156);
xor UO_2313 (O_2313,N_15965,N_17471);
nor UO_2314 (O_2314,N_16393,N_18849);
or UO_2315 (O_2315,N_18862,N_16719);
or UO_2316 (O_2316,N_19429,N_17765);
and UO_2317 (O_2317,N_15332,N_19214);
and UO_2318 (O_2318,N_17412,N_19072);
and UO_2319 (O_2319,N_16190,N_17622);
xnor UO_2320 (O_2320,N_19723,N_17732);
xor UO_2321 (O_2321,N_15228,N_17291);
nand UO_2322 (O_2322,N_18192,N_18482);
nand UO_2323 (O_2323,N_16581,N_17592);
and UO_2324 (O_2324,N_18971,N_16801);
nor UO_2325 (O_2325,N_18700,N_15807);
and UO_2326 (O_2326,N_16235,N_19137);
nand UO_2327 (O_2327,N_18215,N_16798);
nor UO_2328 (O_2328,N_17694,N_19189);
or UO_2329 (O_2329,N_15841,N_19163);
and UO_2330 (O_2330,N_16041,N_15039);
nor UO_2331 (O_2331,N_18007,N_19296);
nor UO_2332 (O_2332,N_17815,N_16065);
xnor UO_2333 (O_2333,N_18360,N_17773);
nand UO_2334 (O_2334,N_16208,N_19633);
and UO_2335 (O_2335,N_15867,N_16675);
nor UO_2336 (O_2336,N_16917,N_17485);
and UO_2337 (O_2337,N_19990,N_19712);
nor UO_2338 (O_2338,N_15955,N_18115);
nor UO_2339 (O_2339,N_15011,N_15648);
xnor UO_2340 (O_2340,N_17202,N_15750);
or UO_2341 (O_2341,N_15441,N_19477);
xnor UO_2342 (O_2342,N_18052,N_16223);
and UO_2343 (O_2343,N_18873,N_19573);
and UO_2344 (O_2344,N_18099,N_18458);
and UO_2345 (O_2345,N_17140,N_17131);
or UO_2346 (O_2346,N_17070,N_18472);
nand UO_2347 (O_2347,N_19575,N_19052);
and UO_2348 (O_2348,N_17378,N_17044);
nor UO_2349 (O_2349,N_19140,N_18197);
or UO_2350 (O_2350,N_15374,N_16966);
or UO_2351 (O_2351,N_17896,N_16782);
and UO_2352 (O_2352,N_15409,N_15476);
or UO_2353 (O_2353,N_15279,N_16513);
xor UO_2354 (O_2354,N_18563,N_15123);
and UO_2355 (O_2355,N_19413,N_15537);
or UO_2356 (O_2356,N_18441,N_16152);
xor UO_2357 (O_2357,N_15669,N_18100);
and UO_2358 (O_2358,N_19350,N_18342);
xor UO_2359 (O_2359,N_15814,N_16665);
and UO_2360 (O_2360,N_15373,N_19283);
and UO_2361 (O_2361,N_15820,N_17050);
xnor UO_2362 (O_2362,N_17500,N_19441);
nand UO_2363 (O_2363,N_15744,N_18206);
or UO_2364 (O_2364,N_17275,N_18312);
xnor UO_2365 (O_2365,N_19222,N_19195);
xor UO_2366 (O_2366,N_16283,N_18481);
nand UO_2367 (O_2367,N_16120,N_19539);
or UO_2368 (O_2368,N_16977,N_15307);
and UO_2369 (O_2369,N_15450,N_17366);
xnor UO_2370 (O_2370,N_15134,N_19703);
nor UO_2371 (O_2371,N_17974,N_17014);
or UO_2372 (O_2372,N_18327,N_18403);
nor UO_2373 (O_2373,N_15643,N_17166);
or UO_2374 (O_2374,N_18180,N_18582);
nor UO_2375 (O_2375,N_15179,N_16124);
or UO_2376 (O_2376,N_18543,N_16115);
nand UO_2377 (O_2377,N_18852,N_18656);
nand UO_2378 (O_2378,N_18875,N_15704);
or UO_2379 (O_2379,N_17503,N_16707);
or UO_2380 (O_2380,N_15588,N_15967);
and UO_2381 (O_2381,N_16004,N_17836);
and UO_2382 (O_2382,N_16787,N_16654);
xor UO_2383 (O_2383,N_15872,N_18899);
and UO_2384 (O_2384,N_18407,N_17842);
or UO_2385 (O_2385,N_17571,N_17869);
or UO_2386 (O_2386,N_18397,N_18306);
nand UO_2387 (O_2387,N_18242,N_16221);
and UO_2388 (O_2388,N_15781,N_18904);
and UO_2389 (O_2389,N_15938,N_18105);
nor UO_2390 (O_2390,N_15883,N_17034);
or UO_2391 (O_2391,N_16889,N_19716);
or UO_2392 (O_2392,N_17037,N_15475);
or UO_2393 (O_2393,N_19776,N_16344);
xnor UO_2394 (O_2394,N_15511,N_17373);
xor UO_2395 (O_2395,N_19567,N_15665);
nor UO_2396 (O_2396,N_19614,N_18827);
nand UO_2397 (O_2397,N_16919,N_19558);
nand UO_2398 (O_2398,N_18245,N_18005);
and UO_2399 (O_2399,N_18415,N_15548);
xor UO_2400 (O_2400,N_17990,N_17745);
and UO_2401 (O_2401,N_16511,N_17766);
xnor UO_2402 (O_2402,N_16243,N_18892);
xnor UO_2403 (O_2403,N_18953,N_16083);
nand UO_2404 (O_2404,N_17725,N_19590);
nor UO_2405 (O_2405,N_18165,N_18599);
nor UO_2406 (O_2406,N_16996,N_17005);
xor UO_2407 (O_2407,N_18362,N_19011);
or UO_2408 (O_2408,N_18857,N_16831);
nor UO_2409 (O_2409,N_19377,N_15266);
nor UO_2410 (O_2410,N_16332,N_18833);
and UO_2411 (O_2411,N_15543,N_18140);
nand UO_2412 (O_2412,N_18393,N_19239);
or UO_2413 (O_2413,N_18805,N_19780);
xnor UO_2414 (O_2414,N_15674,N_15347);
and UO_2415 (O_2415,N_16222,N_19436);
and UO_2416 (O_2416,N_19068,N_17088);
xor UO_2417 (O_2417,N_17336,N_18763);
or UO_2418 (O_2418,N_17865,N_18804);
nor UO_2419 (O_2419,N_19474,N_17951);
xnor UO_2420 (O_2420,N_17506,N_17065);
and UO_2421 (O_2421,N_17975,N_16819);
and UO_2422 (O_2422,N_15028,N_16551);
nor UO_2423 (O_2423,N_17150,N_17996);
nor UO_2424 (O_2424,N_16549,N_15413);
xor UO_2425 (O_2425,N_17551,N_19367);
nand UO_2426 (O_2426,N_16954,N_19898);
nand UO_2427 (O_2427,N_19209,N_15393);
xor UO_2428 (O_2428,N_17405,N_19130);
and UO_2429 (O_2429,N_19666,N_19358);
or UO_2430 (O_2430,N_18043,N_18087);
or UO_2431 (O_2431,N_18440,N_17417);
nand UO_2432 (O_2432,N_19205,N_17167);
xnor UO_2433 (O_2433,N_17230,N_19207);
and UO_2434 (O_2434,N_15629,N_16076);
and UO_2435 (O_2435,N_19826,N_19359);
or UO_2436 (O_2436,N_16976,N_15049);
xor UO_2437 (O_2437,N_19681,N_17409);
nand UO_2438 (O_2438,N_19544,N_16091);
xor UO_2439 (O_2439,N_18450,N_16924);
xor UO_2440 (O_2440,N_17632,N_19124);
nand UO_2441 (O_2441,N_16722,N_16728);
xnor UO_2442 (O_2442,N_15411,N_16611);
and UO_2443 (O_2443,N_17033,N_16024);
xnor UO_2444 (O_2444,N_19598,N_17059);
nor UO_2445 (O_2445,N_17493,N_15181);
xor UO_2446 (O_2446,N_15587,N_17606);
nor UO_2447 (O_2447,N_15530,N_15961);
nand UO_2448 (O_2448,N_19353,N_15208);
xnor UO_2449 (O_2449,N_19673,N_16682);
nor UO_2450 (O_2450,N_16702,N_15424);
xor UO_2451 (O_2451,N_15262,N_17257);
nand UO_2452 (O_2452,N_15889,N_19442);
or UO_2453 (O_2453,N_16046,N_19934);
nand UO_2454 (O_2454,N_19153,N_19913);
or UO_2455 (O_2455,N_15157,N_19577);
or UO_2456 (O_2456,N_15603,N_16526);
nor UO_2457 (O_2457,N_15777,N_15376);
and UO_2458 (O_2458,N_15292,N_18172);
nor UO_2459 (O_2459,N_19982,N_16898);
xnor UO_2460 (O_2460,N_16869,N_19019);
and UO_2461 (O_2461,N_15082,N_18939);
and UO_2462 (O_2462,N_17074,N_19369);
and UO_2463 (O_2463,N_15993,N_18033);
xnor UO_2464 (O_2464,N_15788,N_15127);
nand UO_2465 (O_2465,N_15765,N_15490);
nor UO_2466 (O_2466,N_18073,N_18112);
xor UO_2467 (O_2467,N_19115,N_18945);
nor UO_2468 (O_2468,N_15274,N_16381);
and UO_2469 (O_2469,N_15154,N_19373);
or UO_2470 (O_2470,N_18067,N_18338);
nand UO_2471 (O_2471,N_19327,N_19481);
nand UO_2472 (O_2472,N_16980,N_16030);
xor UO_2473 (O_2473,N_16433,N_18886);
and UO_2474 (O_2474,N_18457,N_15810);
or UO_2475 (O_2475,N_15285,N_15324);
or UO_2476 (O_2476,N_19722,N_17753);
and UO_2477 (O_2477,N_15976,N_16156);
nor UO_2478 (O_2478,N_17535,N_15110);
and UO_2479 (O_2479,N_16211,N_19641);
xor UO_2480 (O_2480,N_15949,N_19738);
xor UO_2481 (O_2481,N_18098,N_16348);
or UO_2482 (O_2482,N_19756,N_16686);
and UO_2483 (O_2483,N_17302,N_17881);
or UO_2484 (O_2484,N_17916,N_19521);
nor UO_2485 (O_2485,N_16084,N_17354);
or UO_2486 (O_2486,N_18268,N_16231);
and UO_2487 (O_2487,N_17083,N_18960);
or UO_2488 (O_2488,N_17763,N_16145);
nor UO_2489 (O_2489,N_16858,N_16851);
and UO_2490 (O_2490,N_19330,N_17705);
xor UO_2491 (O_2491,N_19136,N_18670);
or UO_2492 (O_2492,N_18967,N_18168);
xor UO_2493 (O_2493,N_16680,N_15013);
and UO_2494 (O_2494,N_15182,N_19243);
or UO_2495 (O_2495,N_15192,N_15438);
nor UO_2496 (O_2496,N_16991,N_15896);
or UO_2497 (O_2497,N_19281,N_16972);
or UO_2498 (O_2498,N_18933,N_16834);
and UO_2499 (O_2499,N_17515,N_17333);
endmodule