module basic_500_3000_500_4_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_185,In_90);
or U1 (N_1,In_252,In_35);
and U2 (N_2,In_391,In_430);
nor U3 (N_3,In_52,In_268);
or U4 (N_4,In_463,In_455);
nor U5 (N_5,In_406,In_471);
nor U6 (N_6,In_341,In_53);
and U7 (N_7,In_177,In_417);
or U8 (N_8,In_258,In_457);
nand U9 (N_9,In_374,In_480);
nor U10 (N_10,In_272,In_155);
nand U11 (N_11,In_367,In_1);
nand U12 (N_12,In_395,In_420);
or U13 (N_13,In_104,In_426);
or U14 (N_14,In_489,In_124);
or U15 (N_15,In_78,In_393);
or U16 (N_16,In_446,In_232);
nor U17 (N_17,In_76,In_449);
and U18 (N_18,In_100,In_415);
nor U19 (N_19,In_483,In_357);
nand U20 (N_20,In_348,In_458);
nand U21 (N_21,In_413,In_254);
or U22 (N_22,In_392,In_102);
or U23 (N_23,In_166,In_265);
or U24 (N_24,In_214,In_125);
and U25 (N_25,In_157,In_68);
nor U26 (N_26,In_353,In_248);
or U27 (N_27,In_262,In_26);
and U28 (N_28,In_88,In_231);
and U29 (N_29,In_158,In_448);
nor U30 (N_30,In_399,In_182);
nand U31 (N_31,In_274,In_93);
nor U32 (N_32,In_461,In_114);
and U33 (N_33,In_2,In_39);
and U34 (N_34,In_336,In_333);
and U35 (N_35,In_494,In_354);
or U36 (N_36,In_159,In_178);
or U37 (N_37,In_221,In_195);
nand U38 (N_38,In_59,In_80);
or U39 (N_39,In_452,In_116);
and U40 (N_40,In_440,In_427);
nand U41 (N_41,In_99,In_183);
and U42 (N_42,In_325,In_223);
nand U43 (N_43,In_329,In_139);
and U44 (N_44,In_263,In_222);
and U45 (N_45,In_138,In_256);
or U46 (N_46,In_210,In_388);
and U47 (N_47,In_441,In_450);
nand U48 (N_48,In_60,In_21);
or U49 (N_49,In_174,In_322);
nand U50 (N_50,In_239,In_300);
and U51 (N_51,In_285,In_69);
or U52 (N_52,In_267,In_12);
and U53 (N_53,In_375,In_10);
or U54 (N_54,In_246,In_144);
nand U55 (N_55,In_295,In_205);
nor U56 (N_56,In_196,In_108);
nand U57 (N_57,In_270,In_435);
and U58 (N_58,In_291,In_218);
and U59 (N_59,In_276,In_151);
nand U60 (N_60,In_189,In_423);
nand U61 (N_61,In_128,In_14);
and U62 (N_62,In_48,In_234);
nand U63 (N_63,In_310,In_16);
or U64 (N_64,In_193,In_360);
nor U65 (N_65,In_240,In_314);
xnor U66 (N_66,In_3,In_358);
or U67 (N_67,In_204,In_192);
nand U68 (N_68,In_451,In_209);
and U69 (N_69,In_408,In_136);
or U70 (N_70,In_475,In_424);
nor U71 (N_71,In_190,In_419);
and U72 (N_72,In_350,In_137);
nor U73 (N_73,In_343,In_473);
and U74 (N_74,In_57,In_131);
and U75 (N_75,In_95,In_171);
nor U76 (N_76,In_122,In_394);
nand U77 (N_77,In_51,In_429);
and U78 (N_78,In_308,In_135);
nand U79 (N_79,In_313,In_127);
nor U80 (N_80,In_207,In_241);
and U81 (N_81,In_289,In_479);
and U82 (N_82,In_6,In_330);
and U83 (N_83,In_172,In_198);
nor U84 (N_84,In_225,In_89);
nor U85 (N_85,In_273,In_113);
or U86 (N_86,In_443,In_324);
or U87 (N_87,In_376,In_352);
nand U88 (N_88,In_453,In_37);
or U89 (N_89,In_47,In_497);
nand U90 (N_90,In_369,In_142);
nor U91 (N_91,In_50,In_436);
or U92 (N_92,In_377,In_154);
and U93 (N_93,In_111,In_175);
and U94 (N_94,In_86,In_302);
or U95 (N_95,In_188,In_275);
and U96 (N_96,In_130,In_485);
or U97 (N_97,In_98,In_191);
nor U98 (N_98,In_20,In_402);
and U99 (N_99,In_347,In_292);
and U100 (N_100,In_34,In_216);
and U101 (N_101,In_107,In_414);
nand U102 (N_102,In_370,In_181);
and U103 (N_103,In_379,In_168);
nor U104 (N_104,In_421,In_219);
nand U105 (N_105,In_318,In_250);
nand U106 (N_106,In_487,In_320);
nand U107 (N_107,In_13,In_444);
nor U108 (N_108,In_495,In_62);
or U109 (N_109,In_288,In_340);
nand U110 (N_110,In_18,In_396);
nor U111 (N_111,In_397,In_167);
and U112 (N_112,In_38,In_74);
and U113 (N_113,In_432,In_206);
nor U114 (N_114,In_244,In_77);
nand U115 (N_115,In_398,In_148);
or U116 (N_116,In_41,In_72);
nand U117 (N_117,In_409,In_442);
and U118 (N_118,In_488,In_149);
nor U119 (N_119,In_381,In_255);
nor U120 (N_120,In_83,In_213);
or U121 (N_121,In_23,In_30);
and U122 (N_122,In_499,In_115);
nor U123 (N_123,In_110,In_266);
nor U124 (N_124,In_301,In_140);
nor U125 (N_125,In_54,In_416);
and U126 (N_126,In_469,In_94);
nand U127 (N_127,In_306,In_387);
and U128 (N_128,In_141,In_227);
nor U129 (N_129,In_378,In_97);
and U130 (N_130,In_44,In_283);
nand U131 (N_131,In_328,In_152);
nand U132 (N_132,In_9,In_344);
nand U133 (N_133,In_119,In_85);
or U134 (N_134,In_307,In_403);
and U135 (N_135,In_327,In_384);
xnor U136 (N_136,In_143,In_278);
or U137 (N_137,In_304,In_386);
xnor U138 (N_138,In_411,In_153);
or U139 (N_139,In_331,In_456);
nor U140 (N_140,In_257,In_472);
or U141 (N_141,In_431,In_297);
nand U142 (N_142,In_303,In_363);
nor U143 (N_143,In_162,In_82);
nand U144 (N_144,In_418,In_293);
nand U145 (N_145,In_132,In_264);
nand U146 (N_146,In_238,In_372);
nor U147 (N_147,In_280,In_467);
and U148 (N_148,In_184,In_260);
and U149 (N_149,In_362,In_120);
nand U150 (N_150,In_242,In_459);
and U151 (N_151,In_383,In_56);
and U152 (N_152,In_359,In_121);
nor U153 (N_153,In_282,In_58);
nand U154 (N_154,In_17,In_164);
nor U155 (N_155,In_271,In_133);
nor U156 (N_156,In_63,In_5);
or U157 (N_157,In_412,In_237);
and U158 (N_158,In_481,In_101);
or U159 (N_159,In_323,In_326);
nor U160 (N_160,In_253,In_390);
and U161 (N_161,In_490,In_315);
nor U162 (N_162,In_476,In_351);
nand U163 (N_163,In_230,In_169);
nand U164 (N_164,In_25,In_299);
nand U165 (N_165,In_211,In_215);
nand U166 (N_166,In_433,In_66);
or U167 (N_167,In_228,In_79);
and U168 (N_168,In_150,In_296);
nand U169 (N_169,In_45,In_349);
nor U170 (N_170,In_84,In_368);
and U171 (N_171,In_28,In_22);
and U172 (N_172,In_478,In_311);
nand U173 (N_173,In_201,In_466);
and U174 (N_174,In_482,In_4);
xor U175 (N_175,In_46,In_202);
nor U176 (N_176,In_339,In_212);
nand U177 (N_177,In_106,In_249);
or U178 (N_178,In_346,In_356);
and U179 (N_179,In_437,In_492);
nand U180 (N_180,In_405,In_220);
nor U181 (N_181,In_484,In_187);
xor U182 (N_182,In_226,In_493);
and U183 (N_183,In_284,In_55);
or U184 (N_184,In_224,In_464);
nor U185 (N_185,In_199,In_468);
and U186 (N_186,In_496,In_160);
nor U187 (N_187,In_281,In_8);
and U188 (N_188,In_31,In_312);
nor U189 (N_189,In_438,In_269);
xor U190 (N_190,In_27,In_361);
and U191 (N_191,In_425,In_261);
nand U192 (N_192,In_103,In_439);
nand U193 (N_193,In_19,In_147);
nand U194 (N_194,In_477,In_316);
and U195 (N_195,In_259,In_447);
nor U196 (N_196,In_422,In_165);
nand U197 (N_197,In_337,In_309);
nor U198 (N_198,In_197,In_7);
nand U199 (N_199,In_134,In_400);
and U200 (N_200,In_338,In_65);
or U201 (N_201,In_33,In_126);
and U202 (N_202,In_454,In_366);
or U203 (N_203,In_11,In_364);
or U204 (N_204,In_15,In_389);
and U205 (N_205,In_434,In_112);
nand U206 (N_206,In_173,In_145);
or U207 (N_207,In_498,In_96);
nand U208 (N_208,In_380,In_92);
nor U209 (N_209,In_410,In_355);
or U210 (N_210,In_382,In_236);
nand U211 (N_211,In_176,In_64);
nor U212 (N_212,In_404,In_73);
and U213 (N_213,In_32,In_203);
nand U214 (N_214,In_123,In_321);
nor U215 (N_215,In_445,In_109);
nand U216 (N_216,In_117,In_286);
nor U217 (N_217,In_332,In_105);
nor U218 (N_218,In_407,In_24);
and U219 (N_219,In_70,In_294);
nand U220 (N_220,In_335,In_161);
nor U221 (N_221,In_371,In_129);
or U222 (N_222,In_279,In_319);
nor U223 (N_223,In_87,In_287);
nor U224 (N_224,In_474,In_91);
and U225 (N_225,In_36,In_163);
or U226 (N_226,In_470,In_385);
and U227 (N_227,In_401,In_67);
nor U228 (N_228,In_235,In_40);
nand U229 (N_229,In_217,In_298);
or U230 (N_230,In_81,In_229);
nor U231 (N_231,In_179,In_42);
xnor U232 (N_232,In_342,In_334);
nor U233 (N_233,In_317,In_43);
or U234 (N_234,In_233,In_373);
or U235 (N_235,In_29,In_208);
or U236 (N_236,In_194,In_345);
and U237 (N_237,In_247,In_251);
and U238 (N_238,In_305,In_170);
and U239 (N_239,In_290,In_243);
nand U240 (N_240,In_365,In_491);
or U241 (N_241,In_71,In_75);
and U242 (N_242,In_200,In_156);
nor U243 (N_243,In_460,In_486);
or U244 (N_244,In_146,In_462);
nand U245 (N_245,In_245,In_0);
and U246 (N_246,In_180,In_428);
and U247 (N_247,In_186,In_49);
or U248 (N_248,In_277,In_465);
and U249 (N_249,In_118,In_61);
nand U250 (N_250,In_103,In_400);
and U251 (N_251,In_246,In_117);
nor U252 (N_252,In_474,In_433);
or U253 (N_253,In_403,In_160);
nand U254 (N_254,In_367,In_450);
nand U255 (N_255,In_185,In_165);
nor U256 (N_256,In_404,In_475);
nor U257 (N_257,In_468,In_328);
or U258 (N_258,In_183,In_282);
nor U259 (N_259,In_68,In_292);
and U260 (N_260,In_59,In_145);
nor U261 (N_261,In_85,In_310);
and U262 (N_262,In_282,In_463);
or U263 (N_263,In_12,In_141);
nand U264 (N_264,In_85,In_210);
nor U265 (N_265,In_369,In_51);
nor U266 (N_266,In_210,In_243);
nand U267 (N_267,In_151,In_354);
nor U268 (N_268,In_191,In_283);
and U269 (N_269,In_411,In_118);
nor U270 (N_270,In_326,In_136);
nor U271 (N_271,In_49,In_8);
nor U272 (N_272,In_97,In_495);
and U273 (N_273,In_51,In_177);
or U274 (N_274,In_47,In_278);
or U275 (N_275,In_445,In_467);
nor U276 (N_276,In_370,In_31);
and U277 (N_277,In_186,In_301);
and U278 (N_278,In_260,In_489);
nand U279 (N_279,In_95,In_476);
nand U280 (N_280,In_192,In_125);
xor U281 (N_281,In_80,In_328);
or U282 (N_282,In_10,In_156);
or U283 (N_283,In_137,In_335);
and U284 (N_284,In_329,In_149);
and U285 (N_285,In_212,In_287);
or U286 (N_286,In_491,In_46);
or U287 (N_287,In_60,In_455);
nand U288 (N_288,In_9,In_324);
nor U289 (N_289,In_319,In_195);
nand U290 (N_290,In_15,In_413);
or U291 (N_291,In_408,In_82);
or U292 (N_292,In_433,In_67);
nor U293 (N_293,In_177,In_383);
nand U294 (N_294,In_27,In_456);
nor U295 (N_295,In_163,In_349);
or U296 (N_296,In_308,In_383);
nor U297 (N_297,In_14,In_47);
nand U298 (N_298,In_309,In_212);
or U299 (N_299,In_404,In_307);
nor U300 (N_300,In_324,In_20);
xnor U301 (N_301,In_115,In_188);
nor U302 (N_302,In_83,In_180);
nand U303 (N_303,In_235,In_323);
or U304 (N_304,In_207,In_458);
and U305 (N_305,In_291,In_391);
nand U306 (N_306,In_359,In_250);
and U307 (N_307,In_16,In_417);
and U308 (N_308,In_282,In_309);
or U309 (N_309,In_493,In_138);
nand U310 (N_310,In_475,In_476);
nand U311 (N_311,In_124,In_111);
and U312 (N_312,In_391,In_436);
and U313 (N_313,In_387,In_287);
and U314 (N_314,In_197,In_411);
and U315 (N_315,In_37,In_380);
or U316 (N_316,In_225,In_51);
nand U317 (N_317,In_18,In_322);
nand U318 (N_318,In_346,In_332);
nand U319 (N_319,In_202,In_83);
nor U320 (N_320,In_63,In_256);
nor U321 (N_321,In_266,In_111);
and U322 (N_322,In_90,In_152);
and U323 (N_323,In_452,In_70);
nand U324 (N_324,In_487,In_426);
and U325 (N_325,In_214,In_40);
or U326 (N_326,In_216,In_428);
or U327 (N_327,In_203,In_280);
nand U328 (N_328,In_210,In_151);
and U329 (N_329,In_221,In_249);
and U330 (N_330,In_194,In_251);
or U331 (N_331,In_453,In_255);
nand U332 (N_332,In_180,In_217);
nor U333 (N_333,In_16,In_281);
and U334 (N_334,In_365,In_42);
nor U335 (N_335,In_486,In_138);
nand U336 (N_336,In_59,In_0);
nor U337 (N_337,In_373,In_290);
xor U338 (N_338,In_499,In_498);
nand U339 (N_339,In_14,In_360);
nand U340 (N_340,In_71,In_299);
nand U341 (N_341,In_272,In_429);
and U342 (N_342,In_297,In_94);
or U343 (N_343,In_223,In_224);
or U344 (N_344,In_69,In_422);
or U345 (N_345,In_126,In_270);
nand U346 (N_346,In_314,In_280);
nand U347 (N_347,In_162,In_412);
and U348 (N_348,In_138,In_339);
and U349 (N_349,In_257,In_264);
and U350 (N_350,In_46,In_313);
or U351 (N_351,In_478,In_438);
nand U352 (N_352,In_7,In_286);
nand U353 (N_353,In_280,In_299);
or U354 (N_354,In_426,In_437);
and U355 (N_355,In_326,In_73);
or U356 (N_356,In_137,In_203);
and U357 (N_357,In_67,In_34);
or U358 (N_358,In_96,In_251);
nand U359 (N_359,In_476,In_138);
nor U360 (N_360,In_349,In_30);
and U361 (N_361,In_283,In_99);
and U362 (N_362,In_469,In_335);
and U363 (N_363,In_378,In_405);
and U364 (N_364,In_426,In_202);
nand U365 (N_365,In_328,In_396);
nor U366 (N_366,In_365,In_40);
xor U367 (N_367,In_376,In_154);
and U368 (N_368,In_417,In_342);
nor U369 (N_369,In_494,In_123);
and U370 (N_370,In_56,In_60);
nand U371 (N_371,In_352,In_431);
nor U372 (N_372,In_63,In_230);
nor U373 (N_373,In_287,In_278);
nand U374 (N_374,In_303,In_427);
and U375 (N_375,In_251,In_273);
nor U376 (N_376,In_451,In_91);
nor U377 (N_377,In_453,In_274);
or U378 (N_378,In_181,In_108);
or U379 (N_379,In_88,In_150);
and U380 (N_380,In_369,In_87);
and U381 (N_381,In_423,In_412);
nor U382 (N_382,In_463,In_4);
and U383 (N_383,In_174,In_402);
nor U384 (N_384,In_271,In_235);
and U385 (N_385,In_300,In_270);
nor U386 (N_386,In_490,In_90);
nor U387 (N_387,In_332,In_27);
or U388 (N_388,In_403,In_271);
nor U389 (N_389,In_121,In_217);
nor U390 (N_390,In_231,In_293);
and U391 (N_391,In_65,In_480);
and U392 (N_392,In_362,In_263);
nand U393 (N_393,In_493,In_475);
or U394 (N_394,In_230,In_46);
nand U395 (N_395,In_69,In_50);
and U396 (N_396,In_486,In_80);
nand U397 (N_397,In_401,In_362);
or U398 (N_398,In_106,In_391);
nor U399 (N_399,In_445,In_312);
or U400 (N_400,In_57,In_327);
nor U401 (N_401,In_103,In_47);
nand U402 (N_402,In_116,In_115);
nand U403 (N_403,In_205,In_46);
and U404 (N_404,In_252,In_106);
or U405 (N_405,In_198,In_199);
nor U406 (N_406,In_295,In_208);
or U407 (N_407,In_168,In_351);
or U408 (N_408,In_210,In_308);
nand U409 (N_409,In_352,In_12);
and U410 (N_410,In_58,In_315);
nand U411 (N_411,In_401,In_60);
or U412 (N_412,In_365,In_151);
and U413 (N_413,In_179,In_199);
nand U414 (N_414,In_382,In_447);
nand U415 (N_415,In_245,In_94);
nand U416 (N_416,In_397,In_235);
or U417 (N_417,In_212,In_436);
or U418 (N_418,In_272,In_131);
nor U419 (N_419,In_165,In_39);
or U420 (N_420,In_329,In_154);
nand U421 (N_421,In_407,In_5);
and U422 (N_422,In_15,In_54);
nor U423 (N_423,In_203,In_62);
and U424 (N_424,In_443,In_271);
nand U425 (N_425,In_135,In_434);
or U426 (N_426,In_339,In_113);
nand U427 (N_427,In_326,In_467);
and U428 (N_428,In_229,In_201);
and U429 (N_429,In_307,In_469);
or U430 (N_430,In_314,In_92);
or U431 (N_431,In_240,In_432);
nand U432 (N_432,In_25,In_298);
nand U433 (N_433,In_272,In_7);
and U434 (N_434,In_130,In_225);
or U435 (N_435,In_295,In_491);
nor U436 (N_436,In_408,In_192);
nor U437 (N_437,In_262,In_422);
nand U438 (N_438,In_209,In_351);
nand U439 (N_439,In_410,In_484);
nand U440 (N_440,In_380,In_280);
and U441 (N_441,In_16,In_96);
nand U442 (N_442,In_429,In_309);
and U443 (N_443,In_67,In_193);
nor U444 (N_444,In_324,In_83);
or U445 (N_445,In_431,In_111);
and U446 (N_446,In_101,In_266);
or U447 (N_447,In_313,In_120);
or U448 (N_448,In_40,In_190);
nor U449 (N_449,In_57,In_55);
and U450 (N_450,In_140,In_396);
nand U451 (N_451,In_82,In_357);
and U452 (N_452,In_383,In_494);
nand U453 (N_453,In_129,In_269);
nor U454 (N_454,In_422,In_421);
nor U455 (N_455,In_210,In_429);
or U456 (N_456,In_158,In_186);
nor U457 (N_457,In_44,In_71);
or U458 (N_458,In_379,In_494);
and U459 (N_459,In_455,In_114);
nand U460 (N_460,In_172,In_461);
xnor U461 (N_461,In_435,In_153);
nand U462 (N_462,In_352,In_451);
and U463 (N_463,In_347,In_211);
nor U464 (N_464,In_481,In_447);
and U465 (N_465,In_89,In_280);
nor U466 (N_466,In_34,In_315);
and U467 (N_467,In_322,In_9);
nor U468 (N_468,In_122,In_48);
or U469 (N_469,In_41,In_89);
nand U470 (N_470,In_14,In_236);
and U471 (N_471,In_387,In_188);
or U472 (N_472,In_21,In_377);
nor U473 (N_473,In_146,In_120);
or U474 (N_474,In_185,In_438);
or U475 (N_475,In_140,In_352);
or U476 (N_476,In_26,In_461);
nand U477 (N_477,In_296,In_466);
nand U478 (N_478,In_366,In_92);
and U479 (N_479,In_301,In_344);
nor U480 (N_480,In_443,In_178);
xnor U481 (N_481,In_100,In_199);
nor U482 (N_482,In_433,In_30);
nor U483 (N_483,In_352,In_413);
nor U484 (N_484,In_209,In_281);
nor U485 (N_485,In_453,In_132);
or U486 (N_486,In_241,In_442);
or U487 (N_487,In_65,In_188);
nor U488 (N_488,In_167,In_488);
nand U489 (N_489,In_261,In_449);
or U490 (N_490,In_141,In_86);
or U491 (N_491,In_491,In_253);
nand U492 (N_492,In_330,In_289);
and U493 (N_493,In_356,In_65);
or U494 (N_494,In_365,In_56);
nor U495 (N_495,In_249,In_432);
or U496 (N_496,In_14,In_424);
and U497 (N_497,In_113,In_76);
and U498 (N_498,In_160,In_389);
or U499 (N_499,In_456,In_271);
and U500 (N_500,In_383,In_152);
and U501 (N_501,In_175,In_453);
or U502 (N_502,In_305,In_341);
or U503 (N_503,In_244,In_68);
or U504 (N_504,In_33,In_421);
or U505 (N_505,In_81,In_69);
nor U506 (N_506,In_165,In_15);
xnor U507 (N_507,In_122,In_303);
nand U508 (N_508,In_182,In_257);
nand U509 (N_509,In_164,In_84);
nand U510 (N_510,In_245,In_212);
xor U511 (N_511,In_131,In_303);
nand U512 (N_512,In_247,In_167);
nand U513 (N_513,In_365,In_13);
and U514 (N_514,In_304,In_279);
nor U515 (N_515,In_27,In_433);
and U516 (N_516,In_439,In_60);
and U517 (N_517,In_481,In_290);
or U518 (N_518,In_281,In_487);
and U519 (N_519,In_225,In_223);
nand U520 (N_520,In_289,In_388);
and U521 (N_521,In_168,In_69);
nand U522 (N_522,In_140,In_424);
nand U523 (N_523,In_437,In_67);
or U524 (N_524,In_107,In_326);
nand U525 (N_525,In_134,In_29);
nor U526 (N_526,In_45,In_117);
nor U527 (N_527,In_333,In_206);
nor U528 (N_528,In_331,In_13);
nor U529 (N_529,In_273,In_457);
nand U530 (N_530,In_452,In_90);
nor U531 (N_531,In_188,In_431);
nand U532 (N_532,In_485,In_270);
and U533 (N_533,In_409,In_479);
and U534 (N_534,In_49,In_147);
nand U535 (N_535,In_466,In_351);
nor U536 (N_536,In_468,In_20);
and U537 (N_537,In_242,In_78);
nand U538 (N_538,In_65,In_489);
nand U539 (N_539,In_295,In_23);
nand U540 (N_540,In_202,In_443);
or U541 (N_541,In_412,In_354);
or U542 (N_542,In_30,In_96);
nor U543 (N_543,In_24,In_443);
nand U544 (N_544,In_319,In_187);
or U545 (N_545,In_476,In_493);
and U546 (N_546,In_126,In_443);
or U547 (N_547,In_211,In_386);
or U548 (N_548,In_316,In_30);
nand U549 (N_549,In_414,In_256);
and U550 (N_550,In_214,In_10);
and U551 (N_551,In_90,In_483);
and U552 (N_552,In_220,In_316);
and U553 (N_553,In_134,In_490);
nand U554 (N_554,In_9,In_439);
nor U555 (N_555,In_306,In_280);
and U556 (N_556,In_47,In_53);
and U557 (N_557,In_408,In_150);
nor U558 (N_558,In_177,In_402);
and U559 (N_559,In_444,In_15);
nand U560 (N_560,In_343,In_65);
nor U561 (N_561,In_424,In_152);
or U562 (N_562,In_359,In_15);
or U563 (N_563,In_111,In_242);
nand U564 (N_564,In_432,In_3);
and U565 (N_565,In_277,In_264);
and U566 (N_566,In_150,In_41);
and U567 (N_567,In_13,In_202);
nor U568 (N_568,In_345,In_491);
or U569 (N_569,In_419,In_443);
or U570 (N_570,In_447,In_281);
nand U571 (N_571,In_264,In_173);
nor U572 (N_572,In_80,In_1);
nand U573 (N_573,In_142,In_53);
and U574 (N_574,In_35,In_177);
nor U575 (N_575,In_292,In_275);
nor U576 (N_576,In_12,In_483);
nand U577 (N_577,In_246,In_236);
and U578 (N_578,In_246,In_208);
and U579 (N_579,In_395,In_29);
and U580 (N_580,In_70,In_282);
nor U581 (N_581,In_337,In_486);
or U582 (N_582,In_201,In_237);
and U583 (N_583,In_274,In_125);
nand U584 (N_584,In_433,In_77);
or U585 (N_585,In_102,In_394);
or U586 (N_586,In_387,In_178);
nor U587 (N_587,In_205,In_324);
xor U588 (N_588,In_289,In_253);
and U589 (N_589,In_345,In_113);
nor U590 (N_590,In_484,In_285);
and U591 (N_591,In_455,In_82);
nor U592 (N_592,In_182,In_123);
nand U593 (N_593,In_303,In_423);
nand U594 (N_594,In_6,In_129);
or U595 (N_595,In_378,In_343);
nand U596 (N_596,In_55,In_214);
and U597 (N_597,In_35,In_386);
xnor U598 (N_598,In_19,In_228);
or U599 (N_599,In_434,In_444);
or U600 (N_600,In_5,In_173);
or U601 (N_601,In_431,In_123);
or U602 (N_602,In_68,In_342);
nor U603 (N_603,In_309,In_343);
nor U604 (N_604,In_136,In_73);
and U605 (N_605,In_326,In_109);
and U606 (N_606,In_27,In_366);
nor U607 (N_607,In_0,In_51);
and U608 (N_608,In_3,In_101);
or U609 (N_609,In_396,In_16);
nor U610 (N_610,In_194,In_198);
and U611 (N_611,In_425,In_165);
nand U612 (N_612,In_262,In_367);
nor U613 (N_613,In_434,In_9);
or U614 (N_614,In_323,In_449);
or U615 (N_615,In_158,In_307);
or U616 (N_616,In_263,In_107);
nand U617 (N_617,In_131,In_347);
nand U618 (N_618,In_319,In_424);
or U619 (N_619,In_340,In_462);
or U620 (N_620,In_230,In_196);
and U621 (N_621,In_384,In_406);
nor U622 (N_622,In_109,In_43);
nand U623 (N_623,In_478,In_440);
or U624 (N_624,In_223,In_61);
and U625 (N_625,In_121,In_234);
and U626 (N_626,In_425,In_278);
nand U627 (N_627,In_262,In_6);
nand U628 (N_628,In_216,In_79);
nand U629 (N_629,In_39,In_295);
nand U630 (N_630,In_254,In_300);
and U631 (N_631,In_324,In_17);
or U632 (N_632,In_124,In_125);
or U633 (N_633,In_455,In_312);
or U634 (N_634,In_417,In_401);
and U635 (N_635,In_235,In_81);
nand U636 (N_636,In_385,In_277);
nand U637 (N_637,In_131,In_220);
nand U638 (N_638,In_63,In_299);
nand U639 (N_639,In_219,In_496);
and U640 (N_640,In_159,In_462);
or U641 (N_641,In_387,In_185);
or U642 (N_642,In_11,In_48);
nor U643 (N_643,In_15,In_83);
nor U644 (N_644,In_393,In_75);
and U645 (N_645,In_195,In_99);
nor U646 (N_646,In_431,In_60);
and U647 (N_647,In_374,In_52);
nand U648 (N_648,In_254,In_378);
nor U649 (N_649,In_99,In_7);
or U650 (N_650,In_202,In_193);
xor U651 (N_651,In_488,In_230);
and U652 (N_652,In_228,In_154);
nor U653 (N_653,In_455,In_359);
and U654 (N_654,In_401,In_165);
and U655 (N_655,In_330,In_240);
or U656 (N_656,In_285,In_85);
nor U657 (N_657,In_42,In_314);
nor U658 (N_658,In_386,In_95);
nand U659 (N_659,In_353,In_491);
and U660 (N_660,In_289,In_29);
nand U661 (N_661,In_21,In_459);
nand U662 (N_662,In_352,In_276);
or U663 (N_663,In_187,In_218);
nand U664 (N_664,In_390,In_150);
or U665 (N_665,In_71,In_445);
and U666 (N_666,In_461,In_486);
nand U667 (N_667,In_315,In_218);
xor U668 (N_668,In_9,In_435);
and U669 (N_669,In_385,In_199);
nor U670 (N_670,In_371,In_60);
nand U671 (N_671,In_245,In_399);
nor U672 (N_672,In_402,In_41);
and U673 (N_673,In_479,In_443);
nor U674 (N_674,In_432,In_148);
or U675 (N_675,In_407,In_414);
nand U676 (N_676,In_184,In_218);
nor U677 (N_677,In_161,In_63);
or U678 (N_678,In_438,In_243);
nor U679 (N_679,In_319,In_324);
xnor U680 (N_680,In_77,In_103);
and U681 (N_681,In_66,In_243);
or U682 (N_682,In_485,In_204);
nor U683 (N_683,In_352,In_342);
or U684 (N_684,In_283,In_365);
nand U685 (N_685,In_69,In_90);
nand U686 (N_686,In_380,In_140);
and U687 (N_687,In_229,In_344);
nor U688 (N_688,In_375,In_84);
xnor U689 (N_689,In_359,In_325);
nor U690 (N_690,In_276,In_207);
nand U691 (N_691,In_496,In_47);
nand U692 (N_692,In_119,In_278);
or U693 (N_693,In_456,In_452);
and U694 (N_694,In_381,In_390);
and U695 (N_695,In_31,In_441);
nor U696 (N_696,In_148,In_232);
and U697 (N_697,In_125,In_118);
and U698 (N_698,In_217,In_172);
or U699 (N_699,In_156,In_389);
nand U700 (N_700,In_339,In_380);
and U701 (N_701,In_443,In_432);
nand U702 (N_702,In_373,In_405);
nor U703 (N_703,In_166,In_7);
nand U704 (N_704,In_312,In_382);
nand U705 (N_705,In_298,In_277);
and U706 (N_706,In_195,In_273);
or U707 (N_707,In_227,In_52);
or U708 (N_708,In_162,In_185);
or U709 (N_709,In_456,In_366);
nand U710 (N_710,In_382,In_116);
or U711 (N_711,In_327,In_29);
nor U712 (N_712,In_250,In_255);
nand U713 (N_713,In_168,In_215);
and U714 (N_714,In_492,In_99);
nor U715 (N_715,In_336,In_343);
nand U716 (N_716,In_231,In_381);
and U717 (N_717,In_320,In_448);
and U718 (N_718,In_107,In_491);
nand U719 (N_719,In_431,In_179);
and U720 (N_720,In_418,In_251);
or U721 (N_721,In_189,In_46);
nor U722 (N_722,In_294,In_59);
nor U723 (N_723,In_90,In_77);
or U724 (N_724,In_206,In_179);
nand U725 (N_725,In_178,In_149);
or U726 (N_726,In_204,In_414);
and U727 (N_727,In_120,In_408);
and U728 (N_728,In_135,In_375);
and U729 (N_729,In_188,In_189);
nand U730 (N_730,In_317,In_341);
or U731 (N_731,In_304,In_363);
nor U732 (N_732,In_474,In_73);
and U733 (N_733,In_18,In_46);
nor U734 (N_734,In_10,In_181);
and U735 (N_735,In_179,In_401);
or U736 (N_736,In_405,In_337);
or U737 (N_737,In_398,In_462);
or U738 (N_738,In_89,In_388);
or U739 (N_739,In_135,In_279);
and U740 (N_740,In_290,In_124);
nand U741 (N_741,In_376,In_484);
and U742 (N_742,In_133,In_8);
nand U743 (N_743,In_208,In_285);
and U744 (N_744,In_145,In_460);
nand U745 (N_745,In_485,In_219);
nand U746 (N_746,In_130,In_210);
nand U747 (N_747,In_361,In_247);
and U748 (N_748,In_375,In_53);
nor U749 (N_749,In_423,In_23);
nand U750 (N_750,N_381,N_338);
nor U751 (N_751,N_67,N_721);
nor U752 (N_752,N_488,N_442);
and U753 (N_753,N_164,N_745);
and U754 (N_754,N_58,N_181);
nand U755 (N_755,N_710,N_341);
nand U756 (N_756,N_129,N_42);
nand U757 (N_757,N_423,N_637);
or U758 (N_758,N_39,N_545);
nand U759 (N_759,N_279,N_621);
nor U760 (N_760,N_91,N_403);
nand U761 (N_761,N_747,N_509);
xor U762 (N_762,N_746,N_298);
and U763 (N_763,N_141,N_521);
and U764 (N_764,N_501,N_567);
nand U765 (N_765,N_477,N_420);
and U766 (N_766,N_331,N_395);
nor U767 (N_767,N_378,N_617);
or U768 (N_768,N_573,N_411);
and U769 (N_769,N_296,N_51);
nand U770 (N_770,N_684,N_169);
or U771 (N_771,N_356,N_28);
or U772 (N_772,N_154,N_78);
nand U773 (N_773,N_512,N_301);
or U774 (N_774,N_278,N_363);
nand U775 (N_775,N_344,N_74);
nand U776 (N_776,N_694,N_446);
nand U777 (N_777,N_466,N_360);
nand U778 (N_778,N_185,N_170);
and U779 (N_779,N_236,N_566);
nor U780 (N_780,N_475,N_43);
nand U781 (N_781,N_66,N_514);
and U782 (N_782,N_744,N_415);
or U783 (N_783,N_166,N_398);
or U784 (N_784,N_30,N_93);
and U785 (N_785,N_741,N_577);
nand U786 (N_786,N_46,N_16);
nand U787 (N_787,N_49,N_602);
nor U788 (N_788,N_693,N_604);
nor U789 (N_789,N_661,N_585);
and U790 (N_790,N_406,N_148);
nand U791 (N_791,N_620,N_699);
nand U792 (N_792,N_561,N_48);
and U793 (N_793,N_242,N_323);
or U794 (N_794,N_649,N_161);
nand U795 (N_795,N_535,N_603);
and U796 (N_796,N_229,N_720);
or U797 (N_797,N_714,N_13);
and U798 (N_798,N_272,N_232);
nand U799 (N_799,N_180,N_64);
and U800 (N_800,N_367,N_332);
nand U801 (N_801,N_438,N_238);
nand U802 (N_802,N_739,N_677);
nor U803 (N_803,N_664,N_17);
nand U804 (N_804,N_625,N_105);
nor U805 (N_805,N_76,N_676);
nand U806 (N_806,N_366,N_708);
and U807 (N_807,N_245,N_412);
and U808 (N_808,N_109,N_276);
and U809 (N_809,N_251,N_510);
nor U810 (N_810,N_294,N_327);
nand U811 (N_811,N_309,N_408);
nor U812 (N_812,N_71,N_80);
and U813 (N_813,N_526,N_613);
nor U814 (N_814,N_100,N_706);
and U815 (N_815,N_84,N_659);
or U816 (N_816,N_686,N_350);
or U817 (N_817,N_128,N_143);
or U818 (N_818,N_86,N_319);
xnor U819 (N_819,N_611,N_565);
nor U820 (N_820,N_287,N_160);
nor U821 (N_821,N_337,N_99);
and U822 (N_822,N_440,N_217);
or U823 (N_823,N_583,N_155);
or U824 (N_824,N_473,N_608);
and U825 (N_825,N_144,N_299);
nor U826 (N_826,N_392,N_18);
or U827 (N_827,N_98,N_303);
and U828 (N_828,N_104,N_179);
and U829 (N_829,N_389,N_671);
nand U830 (N_830,N_549,N_594);
nand U831 (N_831,N_616,N_244);
and U832 (N_832,N_725,N_87);
nor U833 (N_833,N_701,N_667);
or U834 (N_834,N_547,N_639);
nand U835 (N_835,N_347,N_83);
nand U836 (N_836,N_644,N_569);
or U837 (N_837,N_384,N_10);
and U838 (N_838,N_727,N_199);
or U839 (N_839,N_588,N_252);
nand U840 (N_840,N_702,N_692);
xor U841 (N_841,N_543,N_376);
and U842 (N_842,N_24,N_559);
nand U843 (N_843,N_716,N_57);
nor U844 (N_844,N_742,N_665);
nor U845 (N_845,N_162,N_351);
nor U846 (N_846,N_421,N_601);
nand U847 (N_847,N_580,N_352);
or U848 (N_848,N_499,N_4);
or U849 (N_849,N_318,N_19);
and U850 (N_850,N_127,N_231);
and U851 (N_851,N_47,N_270);
or U852 (N_852,N_263,N_503);
or U853 (N_853,N_191,N_189);
nor U854 (N_854,N_623,N_619);
nor U855 (N_855,N_622,N_377);
nor U856 (N_856,N_250,N_142);
or U857 (N_857,N_633,N_106);
or U858 (N_858,N_688,N_461);
nand U859 (N_859,N_192,N_146);
nor U860 (N_860,N_414,N_346);
nand U861 (N_861,N_190,N_541);
or U862 (N_862,N_655,N_120);
xnor U863 (N_863,N_295,N_228);
nor U864 (N_864,N_564,N_738);
or U865 (N_865,N_679,N_648);
nand U866 (N_866,N_218,N_612);
nand U867 (N_867,N_70,N_111);
or U868 (N_868,N_273,N_172);
or U869 (N_869,N_426,N_314);
or U870 (N_870,N_399,N_646);
nor U871 (N_871,N_463,N_454);
or U872 (N_872,N_419,N_570);
and U873 (N_873,N_410,N_530);
and U874 (N_874,N_578,N_221);
nand U875 (N_875,N_416,N_262);
nor U876 (N_876,N_394,N_449);
and U877 (N_877,N_207,N_507);
nand U878 (N_878,N_306,N_134);
or U879 (N_879,N_519,N_125);
nand U880 (N_880,N_464,N_371);
or U881 (N_881,N_364,N_115);
nor U882 (N_882,N_266,N_551);
and U883 (N_883,N_248,N_418);
nor U884 (N_884,N_103,N_660);
nand U885 (N_885,N_370,N_215);
nand U886 (N_886,N_534,N_25);
nand U887 (N_887,N_178,N_3);
nand U888 (N_888,N_224,N_348);
and U889 (N_889,N_736,N_313);
or U890 (N_890,N_428,N_536);
and U891 (N_891,N_568,N_27);
nand U892 (N_892,N_41,N_670);
or U893 (N_893,N_196,N_642);
nand U894 (N_894,N_495,N_44);
nor U895 (N_895,N_246,N_730);
or U896 (N_896,N_167,N_579);
and U897 (N_897,N_304,N_157);
or U898 (N_898,N_293,N_422);
and U899 (N_899,N_544,N_197);
or U900 (N_900,N_525,N_413);
nor U901 (N_901,N_233,N_73);
nand U902 (N_902,N_21,N_479);
or U903 (N_903,N_689,N_139);
or U904 (N_904,N_393,N_606);
and U905 (N_905,N_553,N_733);
or U906 (N_906,N_560,N_322);
or U907 (N_907,N_444,N_65);
nand U908 (N_908,N_433,N_333);
nand U909 (N_909,N_54,N_195);
nand U910 (N_910,N_213,N_200);
nor U911 (N_911,N_374,N_69);
nor U912 (N_912,N_335,N_500);
and U913 (N_913,N_532,N_77);
or U914 (N_914,N_386,N_361);
nor U915 (N_915,N_305,N_235);
nand U916 (N_916,N_237,N_220);
and U917 (N_917,N_581,N_518);
and U918 (N_918,N_307,N_290);
nor U919 (N_919,N_362,N_15);
nor U920 (N_920,N_194,N_523);
and U921 (N_921,N_522,N_88);
or U922 (N_922,N_82,N_268);
nand U923 (N_923,N_432,N_498);
or U924 (N_924,N_615,N_445);
nor U925 (N_925,N_204,N_265);
or U926 (N_926,N_187,N_533);
nor U927 (N_927,N_696,N_112);
nor U928 (N_928,N_516,N_554);
or U929 (N_929,N_425,N_385);
or U930 (N_930,N_586,N_599);
or U931 (N_931,N_528,N_183);
nor U932 (N_932,N_126,N_320);
and U933 (N_933,N_494,N_373);
and U934 (N_934,N_123,N_254);
and U935 (N_935,N_90,N_355);
or U936 (N_936,N_651,N_315);
or U937 (N_937,N_223,N_548);
or U938 (N_938,N_455,N_632);
or U939 (N_939,N_529,N_285);
or U940 (N_940,N_614,N_211);
and U941 (N_941,N_711,N_317);
nor U942 (N_942,N_206,N_85);
or U943 (N_943,N_339,N_508);
nor U944 (N_944,N_102,N_124);
nor U945 (N_945,N_743,N_349);
or U946 (N_946,N_1,N_557);
or U947 (N_947,N_45,N_584);
nor U948 (N_948,N_645,N_424);
nand U949 (N_949,N_214,N_81);
or U950 (N_950,N_343,N_683);
nand U951 (N_951,N_205,N_609);
and U952 (N_952,N_354,N_329);
nand U953 (N_953,N_662,N_291);
or U954 (N_954,N_476,N_216);
nand U955 (N_955,N_277,N_666);
nor U956 (N_956,N_404,N_517);
and U957 (N_957,N_717,N_718);
nor U958 (N_958,N_152,N_435);
nand U959 (N_959,N_647,N_174);
or U960 (N_960,N_537,N_249);
or U961 (N_961,N_118,N_36);
or U962 (N_962,N_219,N_452);
nand U963 (N_963,N_168,N_110);
nor U964 (N_964,N_467,N_643);
nor U965 (N_965,N_629,N_504);
and U966 (N_966,N_540,N_492);
and U967 (N_967,N_558,N_685);
or U968 (N_968,N_133,N_429);
nor U969 (N_969,N_62,N_12);
or U970 (N_970,N_490,N_101);
nand U971 (N_971,N_95,N_258);
or U972 (N_972,N_122,N_531);
nor U973 (N_973,N_470,N_552);
nor U974 (N_974,N_247,N_626);
or U975 (N_975,N_32,N_257);
or U976 (N_976,N_462,N_75);
and U977 (N_977,N_259,N_726);
nand U978 (N_978,N_222,N_486);
and U979 (N_979,N_663,N_14);
or U980 (N_980,N_729,N_22);
or U981 (N_981,N_690,N_695);
nor U982 (N_982,N_198,N_704);
nand U983 (N_983,N_555,N_358);
or U984 (N_984,N_527,N_0);
and U985 (N_985,N_437,N_388);
nand U986 (N_986,N_311,N_596);
nand U987 (N_987,N_177,N_68);
or U988 (N_988,N_723,N_737);
or U989 (N_989,N_63,N_482);
nor U990 (N_990,N_147,N_345);
nor U991 (N_991,N_330,N_260);
nand U992 (N_992,N_130,N_610);
nor U993 (N_993,N_480,N_203);
nand U994 (N_994,N_441,N_156);
nand U995 (N_995,N_59,N_748);
or U996 (N_996,N_740,N_340);
and U997 (N_997,N_669,N_640);
nand U998 (N_998,N_713,N_634);
nand U999 (N_999,N_712,N_587);
nand U1000 (N_1000,N_575,N_539);
and U1001 (N_1001,N_297,N_321);
nor U1002 (N_1002,N_208,N_241);
nor U1003 (N_1003,N_735,N_158);
and U1004 (N_1004,N_401,N_145);
nor U1005 (N_1005,N_505,N_201);
or U1006 (N_1006,N_485,N_402);
nand U1007 (N_1007,N_23,N_357);
nand U1008 (N_1008,N_31,N_675);
and U1009 (N_1009,N_137,N_556);
or U1010 (N_1010,N_448,N_468);
nor U1011 (N_1011,N_472,N_89);
xnor U1012 (N_1012,N_114,N_607);
nand U1013 (N_1013,N_496,N_26);
or U1014 (N_1014,N_453,N_728);
and U1015 (N_1015,N_2,N_227);
and U1016 (N_1016,N_572,N_184);
and U1017 (N_1017,N_538,N_286);
nor U1018 (N_1018,N_369,N_107);
nor U1019 (N_1019,N_40,N_635);
nand U1020 (N_1020,N_308,N_636);
or U1021 (N_1021,N_300,N_546);
nor U1022 (N_1022,N_243,N_230);
and U1023 (N_1023,N_368,N_117);
and U1024 (N_1024,N_34,N_576);
or U1025 (N_1025,N_591,N_724);
nor U1026 (N_1026,N_457,N_202);
nor U1027 (N_1027,N_682,N_439);
nor U1028 (N_1028,N_691,N_149);
nor U1029 (N_1029,N_240,N_407);
or U1030 (N_1030,N_653,N_390);
or U1031 (N_1031,N_605,N_571);
nand U1032 (N_1032,N_52,N_574);
nor U1033 (N_1033,N_328,N_597);
or U1034 (N_1034,N_289,N_175);
nand U1035 (N_1035,N_431,N_732);
and U1036 (N_1036,N_281,N_72);
or U1037 (N_1037,N_282,N_481);
nand U1038 (N_1038,N_478,N_734);
nor U1039 (N_1039,N_20,N_234);
and U1040 (N_1040,N_312,N_600);
nand U1041 (N_1041,N_650,N_590);
nor U1042 (N_1042,N_261,N_61);
and U1043 (N_1043,N_680,N_94);
nor U1044 (N_1044,N_292,N_434);
nand U1045 (N_1045,N_255,N_562);
nor U1046 (N_1046,N_336,N_491);
or U1047 (N_1047,N_372,N_136);
or U1048 (N_1048,N_37,N_627);
nand U1049 (N_1049,N_471,N_334);
and U1050 (N_1050,N_707,N_631);
or U1051 (N_1051,N_209,N_427);
nor U1052 (N_1052,N_474,N_542);
nor U1053 (N_1053,N_119,N_9);
nand U1054 (N_1054,N_397,N_722);
or U1055 (N_1055,N_436,N_698);
nor U1056 (N_1056,N_8,N_96);
nor U1057 (N_1057,N_113,N_359);
and U1058 (N_1058,N_524,N_430);
or U1059 (N_1059,N_165,N_749);
nand U1060 (N_1060,N_135,N_458);
nand U1061 (N_1061,N_697,N_138);
nor U1062 (N_1062,N_630,N_497);
or U1063 (N_1063,N_267,N_657);
or U1064 (N_1064,N_275,N_469);
nor U1065 (N_1065,N_11,N_92);
nand U1066 (N_1066,N_375,N_163);
xor U1067 (N_1067,N_400,N_153);
or U1068 (N_1068,N_654,N_715);
nand U1069 (N_1069,N_38,N_405);
and U1070 (N_1070,N_226,N_487);
or U1071 (N_1071,N_658,N_176);
nand U1072 (N_1072,N_50,N_116);
and U1073 (N_1073,N_210,N_450);
nand U1074 (N_1074,N_283,N_159);
nand U1075 (N_1075,N_193,N_456);
nand U1076 (N_1076,N_97,N_628);
and U1077 (N_1077,N_731,N_687);
and U1078 (N_1078,N_33,N_56);
nand U1079 (N_1079,N_188,N_53);
and U1080 (N_1080,N_563,N_365);
and U1081 (N_1081,N_379,N_29);
nor U1082 (N_1082,N_310,N_171);
or U1083 (N_1083,N_391,N_55);
nor U1084 (N_1084,N_342,N_672);
nand U1085 (N_1085,N_60,N_668);
and U1086 (N_1086,N_451,N_705);
nor U1087 (N_1087,N_225,N_150);
nand U1088 (N_1088,N_513,N_380);
nor U1089 (N_1089,N_520,N_182);
or U1090 (N_1090,N_79,N_326);
or U1091 (N_1091,N_447,N_483);
or U1092 (N_1092,N_284,N_593);
nor U1093 (N_1093,N_6,N_324);
nand U1094 (N_1094,N_151,N_186);
nand U1095 (N_1095,N_239,N_387);
or U1096 (N_1096,N_35,N_592);
nand U1097 (N_1097,N_256,N_465);
and U1098 (N_1098,N_459,N_595);
and U1099 (N_1099,N_489,N_253);
nand U1100 (N_1100,N_484,N_383);
nand U1101 (N_1101,N_652,N_173);
nor U1102 (N_1102,N_641,N_638);
and U1103 (N_1103,N_506,N_719);
nor U1104 (N_1104,N_316,N_264);
or U1105 (N_1105,N_409,N_460);
nor U1106 (N_1106,N_678,N_288);
and U1107 (N_1107,N_7,N_624);
or U1108 (N_1108,N_325,N_108);
nand U1109 (N_1109,N_589,N_674);
or U1110 (N_1110,N_550,N_511);
nand U1111 (N_1111,N_212,N_502);
or U1112 (N_1112,N_700,N_493);
nor U1113 (N_1113,N_709,N_673);
or U1114 (N_1114,N_618,N_271);
nand U1115 (N_1115,N_382,N_582);
and U1116 (N_1116,N_417,N_269);
nor U1117 (N_1117,N_443,N_5);
nor U1118 (N_1118,N_703,N_132);
and U1119 (N_1119,N_280,N_396);
or U1120 (N_1120,N_598,N_656);
nand U1121 (N_1121,N_131,N_681);
and U1122 (N_1122,N_515,N_140);
or U1123 (N_1123,N_274,N_121);
nor U1124 (N_1124,N_353,N_302);
nor U1125 (N_1125,N_85,N_678);
and U1126 (N_1126,N_127,N_421);
or U1127 (N_1127,N_106,N_75);
and U1128 (N_1128,N_87,N_272);
nor U1129 (N_1129,N_326,N_503);
and U1130 (N_1130,N_714,N_255);
nand U1131 (N_1131,N_669,N_314);
and U1132 (N_1132,N_311,N_128);
and U1133 (N_1133,N_663,N_364);
and U1134 (N_1134,N_422,N_326);
nand U1135 (N_1135,N_586,N_250);
or U1136 (N_1136,N_747,N_463);
and U1137 (N_1137,N_728,N_362);
nand U1138 (N_1138,N_392,N_123);
and U1139 (N_1139,N_557,N_556);
nor U1140 (N_1140,N_497,N_38);
nand U1141 (N_1141,N_661,N_120);
nor U1142 (N_1142,N_345,N_267);
and U1143 (N_1143,N_623,N_296);
nor U1144 (N_1144,N_109,N_475);
nand U1145 (N_1145,N_85,N_195);
and U1146 (N_1146,N_181,N_27);
nor U1147 (N_1147,N_335,N_601);
and U1148 (N_1148,N_521,N_135);
nor U1149 (N_1149,N_566,N_539);
nand U1150 (N_1150,N_324,N_392);
nand U1151 (N_1151,N_163,N_14);
or U1152 (N_1152,N_625,N_473);
and U1153 (N_1153,N_671,N_72);
nand U1154 (N_1154,N_110,N_614);
nor U1155 (N_1155,N_23,N_707);
nor U1156 (N_1156,N_138,N_416);
or U1157 (N_1157,N_557,N_475);
nor U1158 (N_1158,N_738,N_338);
or U1159 (N_1159,N_396,N_270);
or U1160 (N_1160,N_419,N_257);
nand U1161 (N_1161,N_334,N_484);
nand U1162 (N_1162,N_402,N_164);
or U1163 (N_1163,N_689,N_278);
and U1164 (N_1164,N_66,N_589);
and U1165 (N_1165,N_490,N_343);
or U1166 (N_1166,N_301,N_579);
and U1167 (N_1167,N_210,N_326);
and U1168 (N_1168,N_436,N_627);
nor U1169 (N_1169,N_625,N_368);
and U1170 (N_1170,N_141,N_388);
and U1171 (N_1171,N_36,N_462);
and U1172 (N_1172,N_306,N_637);
nor U1173 (N_1173,N_438,N_587);
and U1174 (N_1174,N_633,N_235);
or U1175 (N_1175,N_175,N_589);
and U1176 (N_1176,N_164,N_684);
nand U1177 (N_1177,N_665,N_62);
or U1178 (N_1178,N_170,N_695);
xor U1179 (N_1179,N_493,N_316);
nand U1180 (N_1180,N_21,N_638);
and U1181 (N_1181,N_521,N_712);
nand U1182 (N_1182,N_5,N_409);
and U1183 (N_1183,N_239,N_133);
nand U1184 (N_1184,N_579,N_281);
and U1185 (N_1185,N_522,N_268);
nand U1186 (N_1186,N_514,N_382);
and U1187 (N_1187,N_688,N_327);
or U1188 (N_1188,N_96,N_40);
nand U1189 (N_1189,N_274,N_75);
nand U1190 (N_1190,N_96,N_259);
nand U1191 (N_1191,N_104,N_463);
or U1192 (N_1192,N_402,N_701);
nor U1193 (N_1193,N_394,N_242);
or U1194 (N_1194,N_257,N_402);
and U1195 (N_1195,N_162,N_482);
or U1196 (N_1196,N_33,N_517);
or U1197 (N_1197,N_323,N_47);
and U1198 (N_1198,N_279,N_748);
nor U1199 (N_1199,N_298,N_678);
nor U1200 (N_1200,N_121,N_616);
nand U1201 (N_1201,N_81,N_353);
and U1202 (N_1202,N_557,N_331);
nand U1203 (N_1203,N_263,N_366);
or U1204 (N_1204,N_656,N_595);
nand U1205 (N_1205,N_46,N_172);
nor U1206 (N_1206,N_665,N_673);
or U1207 (N_1207,N_478,N_369);
nand U1208 (N_1208,N_14,N_347);
nor U1209 (N_1209,N_547,N_291);
and U1210 (N_1210,N_437,N_328);
and U1211 (N_1211,N_552,N_422);
or U1212 (N_1212,N_102,N_680);
or U1213 (N_1213,N_354,N_9);
nand U1214 (N_1214,N_742,N_326);
and U1215 (N_1215,N_638,N_653);
nor U1216 (N_1216,N_505,N_247);
and U1217 (N_1217,N_580,N_712);
and U1218 (N_1218,N_406,N_546);
and U1219 (N_1219,N_397,N_148);
and U1220 (N_1220,N_749,N_89);
and U1221 (N_1221,N_68,N_307);
nor U1222 (N_1222,N_493,N_319);
and U1223 (N_1223,N_224,N_232);
and U1224 (N_1224,N_286,N_478);
or U1225 (N_1225,N_455,N_75);
or U1226 (N_1226,N_473,N_606);
nand U1227 (N_1227,N_422,N_472);
nor U1228 (N_1228,N_214,N_154);
and U1229 (N_1229,N_167,N_522);
and U1230 (N_1230,N_407,N_531);
nor U1231 (N_1231,N_336,N_663);
nand U1232 (N_1232,N_746,N_266);
or U1233 (N_1233,N_391,N_16);
nor U1234 (N_1234,N_643,N_363);
and U1235 (N_1235,N_398,N_535);
or U1236 (N_1236,N_398,N_602);
nand U1237 (N_1237,N_4,N_703);
nor U1238 (N_1238,N_88,N_436);
and U1239 (N_1239,N_136,N_242);
nor U1240 (N_1240,N_325,N_259);
nand U1241 (N_1241,N_381,N_663);
and U1242 (N_1242,N_292,N_480);
nand U1243 (N_1243,N_624,N_223);
nor U1244 (N_1244,N_487,N_595);
or U1245 (N_1245,N_427,N_719);
and U1246 (N_1246,N_408,N_582);
and U1247 (N_1247,N_22,N_372);
xnor U1248 (N_1248,N_42,N_223);
nand U1249 (N_1249,N_638,N_493);
nand U1250 (N_1250,N_656,N_630);
and U1251 (N_1251,N_528,N_465);
nand U1252 (N_1252,N_416,N_727);
nor U1253 (N_1253,N_320,N_164);
nor U1254 (N_1254,N_653,N_240);
and U1255 (N_1255,N_261,N_414);
nor U1256 (N_1256,N_161,N_6);
nor U1257 (N_1257,N_702,N_161);
nor U1258 (N_1258,N_0,N_130);
and U1259 (N_1259,N_745,N_104);
and U1260 (N_1260,N_53,N_118);
nor U1261 (N_1261,N_740,N_524);
or U1262 (N_1262,N_511,N_398);
nand U1263 (N_1263,N_669,N_383);
and U1264 (N_1264,N_587,N_105);
xnor U1265 (N_1265,N_633,N_107);
or U1266 (N_1266,N_195,N_244);
nand U1267 (N_1267,N_500,N_171);
nand U1268 (N_1268,N_613,N_55);
and U1269 (N_1269,N_189,N_292);
or U1270 (N_1270,N_715,N_164);
nor U1271 (N_1271,N_323,N_292);
and U1272 (N_1272,N_545,N_20);
nand U1273 (N_1273,N_609,N_400);
or U1274 (N_1274,N_631,N_677);
or U1275 (N_1275,N_106,N_646);
and U1276 (N_1276,N_173,N_412);
nand U1277 (N_1277,N_212,N_48);
and U1278 (N_1278,N_301,N_296);
nor U1279 (N_1279,N_735,N_747);
and U1280 (N_1280,N_467,N_726);
nand U1281 (N_1281,N_648,N_14);
or U1282 (N_1282,N_748,N_417);
and U1283 (N_1283,N_194,N_531);
or U1284 (N_1284,N_701,N_578);
and U1285 (N_1285,N_615,N_175);
or U1286 (N_1286,N_658,N_305);
nand U1287 (N_1287,N_46,N_235);
nand U1288 (N_1288,N_201,N_152);
and U1289 (N_1289,N_231,N_475);
nand U1290 (N_1290,N_379,N_743);
nor U1291 (N_1291,N_362,N_665);
or U1292 (N_1292,N_271,N_114);
nand U1293 (N_1293,N_356,N_85);
or U1294 (N_1294,N_353,N_290);
or U1295 (N_1295,N_704,N_210);
and U1296 (N_1296,N_616,N_86);
and U1297 (N_1297,N_624,N_528);
nand U1298 (N_1298,N_45,N_728);
nor U1299 (N_1299,N_486,N_308);
and U1300 (N_1300,N_404,N_99);
or U1301 (N_1301,N_283,N_499);
or U1302 (N_1302,N_708,N_482);
nand U1303 (N_1303,N_296,N_633);
nor U1304 (N_1304,N_14,N_12);
nand U1305 (N_1305,N_130,N_719);
nand U1306 (N_1306,N_123,N_131);
nor U1307 (N_1307,N_208,N_511);
nor U1308 (N_1308,N_439,N_394);
nor U1309 (N_1309,N_576,N_37);
and U1310 (N_1310,N_428,N_600);
and U1311 (N_1311,N_423,N_536);
and U1312 (N_1312,N_342,N_69);
and U1313 (N_1313,N_450,N_458);
nand U1314 (N_1314,N_492,N_169);
nor U1315 (N_1315,N_232,N_356);
or U1316 (N_1316,N_3,N_298);
or U1317 (N_1317,N_89,N_722);
nand U1318 (N_1318,N_418,N_364);
or U1319 (N_1319,N_80,N_585);
nand U1320 (N_1320,N_297,N_16);
nand U1321 (N_1321,N_675,N_129);
or U1322 (N_1322,N_474,N_475);
or U1323 (N_1323,N_384,N_321);
or U1324 (N_1324,N_65,N_695);
and U1325 (N_1325,N_185,N_336);
nor U1326 (N_1326,N_258,N_249);
or U1327 (N_1327,N_417,N_163);
nand U1328 (N_1328,N_513,N_720);
or U1329 (N_1329,N_184,N_345);
or U1330 (N_1330,N_469,N_177);
and U1331 (N_1331,N_67,N_260);
and U1332 (N_1332,N_731,N_404);
nor U1333 (N_1333,N_133,N_64);
or U1334 (N_1334,N_270,N_259);
or U1335 (N_1335,N_620,N_369);
and U1336 (N_1336,N_132,N_254);
nand U1337 (N_1337,N_732,N_288);
nand U1338 (N_1338,N_214,N_456);
nor U1339 (N_1339,N_504,N_728);
and U1340 (N_1340,N_104,N_220);
nor U1341 (N_1341,N_245,N_47);
nand U1342 (N_1342,N_172,N_418);
nand U1343 (N_1343,N_706,N_62);
nor U1344 (N_1344,N_54,N_602);
and U1345 (N_1345,N_120,N_42);
nand U1346 (N_1346,N_496,N_591);
and U1347 (N_1347,N_93,N_110);
or U1348 (N_1348,N_451,N_447);
nand U1349 (N_1349,N_337,N_223);
nand U1350 (N_1350,N_232,N_708);
nand U1351 (N_1351,N_398,N_26);
and U1352 (N_1352,N_362,N_199);
nor U1353 (N_1353,N_92,N_177);
nand U1354 (N_1354,N_387,N_324);
and U1355 (N_1355,N_365,N_205);
or U1356 (N_1356,N_46,N_379);
nand U1357 (N_1357,N_321,N_66);
and U1358 (N_1358,N_449,N_42);
and U1359 (N_1359,N_382,N_737);
nor U1360 (N_1360,N_238,N_205);
or U1361 (N_1361,N_135,N_578);
nand U1362 (N_1362,N_405,N_41);
or U1363 (N_1363,N_476,N_361);
or U1364 (N_1364,N_145,N_234);
nor U1365 (N_1365,N_683,N_166);
or U1366 (N_1366,N_409,N_201);
nor U1367 (N_1367,N_443,N_684);
or U1368 (N_1368,N_358,N_541);
nand U1369 (N_1369,N_427,N_577);
nand U1370 (N_1370,N_180,N_502);
nor U1371 (N_1371,N_645,N_254);
nand U1372 (N_1372,N_330,N_545);
and U1373 (N_1373,N_83,N_615);
and U1374 (N_1374,N_23,N_662);
nor U1375 (N_1375,N_497,N_742);
or U1376 (N_1376,N_110,N_352);
nor U1377 (N_1377,N_234,N_469);
xor U1378 (N_1378,N_252,N_410);
nand U1379 (N_1379,N_292,N_645);
nor U1380 (N_1380,N_371,N_46);
or U1381 (N_1381,N_584,N_501);
nand U1382 (N_1382,N_539,N_274);
or U1383 (N_1383,N_354,N_24);
or U1384 (N_1384,N_268,N_144);
or U1385 (N_1385,N_274,N_390);
or U1386 (N_1386,N_264,N_227);
or U1387 (N_1387,N_333,N_206);
nand U1388 (N_1388,N_95,N_105);
nor U1389 (N_1389,N_634,N_164);
or U1390 (N_1390,N_79,N_89);
or U1391 (N_1391,N_417,N_257);
and U1392 (N_1392,N_441,N_706);
or U1393 (N_1393,N_602,N_573);
nand U1394 (N_1394,N_424,N_560);
nand U1395 (N_1395,N_126,N_617);
nand U1396 (N_1396,N_596,N_267);
and U1397 (N_1397,N_231,N_575);
and U1398 (N_1398,N_198,N_113);
nor U1399 (N_1399,N_503,N_346);
nand U1400 (N_1400,N_53,N_216);
nor U1401 (N_1401,N_333,N_190);
nor U1402 (N_1402,N_481,N_429);
or U1403 (N_1403,N_74,N_303);
or U1404 (N_1404,N_502,N_360);
nand U1405 (N_1405,N_334,N_211);
or U1406 (N_1406,N_488,N_203);
nand U1407 (N_1407,N_436,N_556);
or U1408 (N_1408,N_594,N_158);
nor U1409 (N_1409,N_747,N_8);
nand U1410 (N_1410,N_607,N_585);
or U1411 (N_1411,N_308,N_407);
nor U1412 (N_1412,N_322,N_44);
or U1413 (N_1413,N_104,N_389);
nor U1414 (N_1414,N_370,N_636);
or U1415 (N_1415,N_269,N_59);
and U1416 (N_1416,N_712,N_211);
and U1417 (N_1417,N_138,N_384);
and U1418 (N_1418,N_525,N_139);
nand U1419 (N_1419,N_61,N_565);
nand U1420 (N_1420,N_456,N_627);
or U1421 (N_1421,N_721,N_659);
nor U1422 (N_1422,N_686,N_614);
nor U1423 (N_1423,N_426,N_280);
nand U1424 (N_1424,N_346,N_559);
and U1425 (N_1425,N_711,N_6);
and U1426 (N_1426,N_641,N_57);
or U1427 (N_1427,N_250,N_426);
or U1428 (N_1428,N_139,N_494);
and U1429 (N_1429,N_748,N_307);
nand U1430 (N_1430,N_396,N_222);
or U1431 (N_1431,N_426,N_510);
and U1432 (N_1432,N_326,N_49);
and U1433 (N_1433,N_63,N_295);
or U1434 (N_1434,N_156,N_214);
or U1435 (N_1435,N_122,N_418);
nor U1436 (N_1436,N_346,N_621);
nor U1437 (N_1437,N_472,N_209);
nand U1438 (N_1438,N_15,N_492);
xor U1439 (N_1439,N_217,N_335);
nor U1440 (N_1440,N_525,N_87);
and U1441 (N_1441,N_145,N_314);
nand U1442 (N_1442,N_229,N_200);
or U1443 (N_1443,N_529,N_710);
nor U1444 (N_1444,N_157,N_108);
nand U1445 (N_1445,N_467,N_731);
or U1446 (N_1446,N_227,N_710);
nand U1447 (N_1447,N_113,N_76);
nand U1448 (N_1448,N_189,N_285);
nand U1449 (N_1449,N_265,N_361);
and U1450 (N_1450,N_422,N_375);
or U1451 (N_1451,N_74,N_182);
and U1452 (N_1452,N_715,N_146);
or U1453 (N_1453,N_344,N_558);
and U1454 (N_1454,N_174,N_450);
nor U1455 (N_1455,N_205,N_30);
nand U1456 (N_1456,N_466,N_165);
and U1457 (N_1457,N_159,N_81);
nand U1458 (N_1458,N_726,N_312);
nor U1459 (N_1459,N_729,N_370);
nor U1460 (N_1460,N_556,N_368);
and U1461 (N_1461,N_153,N_749);
and U1462 (N_1462,N_31,N_339);
nor U1463 (N_1463,N_317,N_721);
or U1464 (N_1464,N_684,N_230);
or U1465 (N_1465,N_733,N_574);
nor U1466 (N_1466,N_42,N_417);
nor U1467 (N_1467,N_106,N_331);
nor U1468 (N_1468,N_424,N_392);
nor U1469 (N_1469,N_400,N_492);
or U1470 (N_1470,N_682,N_437);
nor U1471 (N_1471,N_579,N_363);
nand U1472 (N_1472,N_287,N_272);
or U1473 (N_1473,N_732,N_624);
or U1474 (N_1474,N_548,N_46);
nand U1475 (N_1475,N_98,N_740);
or U1476 (N_1476,N_370,N_442);
or U1477 (N_1477,N_538,N_604);
and U1478 (N_1478,N_108,N_10);
and U1479 (N_1479,N_202,N_630);
and U1480 (N_1480,N_563,N_231);
nor U1481 (N_1481,N_722,N_671);
or U1482 (N_1482,N_389,N_349);
or U1483 (N_1483,N_538,N_420);
nor U1484 (N_1484,N_490,N_390);
nor U1485 (N_1485,N_309,N_279);
and U1486 (N_1486,N_656,N_224);
nand U1487 (N_1487,N_8,N_399);
or U1488 (N_1488,N_211,N_656);
nor U1489 (N_1489,N_202,N_391);
nor U1490 (N_1490,N_128,N_449);
nand U1491 (N_1491,N_635,N_211);
and U1492 (N_1492,N_76,N_422);
and U1493 (N_1493,N_41,N_606);
or U1494 (N_1494,N_461,N_746);
or U1495 (N_1495,N_714,N_549);
xnor U1496 (N_1496,N_356,N_486);
nor U1497 (N_1497,N_739,N_115);
and U1498 (N_1498,N_594,N_36);
and U1499 (N_1499,N_627,N_540);
and U1500 (N_1500,N_1479,N_1152);
nor U1501 (N_1501,N_1274,N_1044);
or U1502 (N_1502,N_1473,N_1302);
and U1503 (N_1503,N_908,N_1363);
or U1504 (N_1504,N_1288,N_1066);
nand U1505 (N_1505,N_1039,N_1403);
or U1506 (N_1506,N_1191,N_925);
nand U1507 (N_1507,N_1432,N_796);
or U1508 (N_1508,N_1014,N_1279);
or U1509 (N_1509,N_1172,N_1205);
or U1510 (N_1510,N_791,N_1483);
nand U1511 (N_1511,N_786,N_1093);
nor U1512 (N_1512,N_1412,N_1034);
nor U1513 (N_1513,N_1420,N_1223);
and U1514 (N_1514,N_1416,N_808);
nand U1515 (N_1515,N_901,N_1224);
or U1516 (N_1516,N_833,N_1115);
or U1517 (N_1517,N_1125,N_966);
or U1518 (N_1518,N_1043,N_848);
nor U1519 (N_1519,N_1258,N_964);
or U1520 (N_1520,N_1084,N_787);
and U1521 (N_1521,N_1293,N_1148);
nor U1522 (N_1522,N_1235,N_1489);
nand U1523 (N_1523,N_1445,N_778);
or U1524 (N_1524,N_1475,N_991);
and U1525 (N_1525,N_1026,N_984);
nor U1526 (N_1526,N_1009,N_1312);
nand U1527 (N_1527,N_1341,N_868);
xor U1528 (N_1528,N_820,N_893);
and U1529 (N_1529,N_920,N_869);
nand U1530 (N_1530,N_1315,N_1415);
nor U1531 (N_1531,N_1217,N_1421);
nand U1532 (N_1532,N_911,N_999);
nand U1533 (N_1533,N_1131,N_1332);
or U1534 (N_1534,N_907,N_1095);
nand U1535 (N_1535,N_1270,N_937);
or U1536 (N_1536,N_1248,N_855);
nand U1537 (N_1537,N_1498,N_1466);
and U1538 (N_1538,N_1135,N_1261);
and U1539 (N_1539,N_1019,N_1283);
or U1540 (N_1540,N_842,N_1331);
and U1541 (N_1541,N_1460,N_1068);
nand U1542 (N_1542,N_934,N_1249);
or U1543 (N_1543,N_1370,N_1220);
nand U1544 (N_1544,N_1423,N_1229);
and U1545 (N_1545,N_1247,N_1256);
nand U1546 (N_1546,N_1444,N_1375);
nand U1547 (N_1547,N_864,N_1311);
nor U1548 (N_1548,N_952,N_1454);
xor U1549 (N_1549,N_1083,N_1150);
or U1550 (N_1550,N_1289,N_903);
or U1551 (N_1551,N_969,N_1273);
xor U1552 (N_1552,N_1435,N_1484);
or U1553 (N_1553,N_1253,N_1409);
or U1554 (N_1554,N_943,N_1330);
and U1555 (N_1555,N_1251,N_823);
nor U1556 (N_1556,N_851,N_1378);
or U1557 (N_1557,N_846,N_1380);
or U1558 (N_1558,N_1338,N_1237);
or U1559 (N_1559,N_1101,N_1397);
nor U1560 (N_1560,N_826,N_850);
nand U1561 (N_1561,N_900,N_895);
and U1562 (N_1562,N_1335,N_827);
or U1563 (N_1563,N_870,N_1309);
and U1564 (N_1564,N_1180,N_1181);
nor U1565 (N_1565,N_1336,N_996);
nand U1566 (N_1566,N_780,N_1314);
nor U1567 (N_1567,N_1342,N_1079);
and U1568 (N_1568,N_871,N_917);
nand U1569 (N_1569,N_845,N_1398);
or U1570 (N_1570,N_1465,N_1052);
and U1571 (N_1571,N_1376,N_1243);
nand U1572 (N_1572,N_1428,N_1063);
or U1573 (N_1573,N_1121,N_1255);
and U1574 (N_1574,N_1456,N_844);
nand U1575 (N_1575,N_879,N_1136);
nand U1576 (N_1576,N_959,N_976);
nor U1577 (N_1577,N_849,N_1451);
nor U1578 (N_1578,N_771,N_1036);
nor U1579 (N_1579,N_1410,N_837);
and U1580 (N_1580,N_1174,N_1097);
nand U1581 (N_1581,N_1455,N_789);
nor U1582 (N_1582,N_927,N_817);
nand U1583 (N_1583,N_1140,N_1004);
or U1584 (N_1584,N_1272,N_804);
nand U1585 (N_1585,N_1276,N_1384);
or U1586 (N_1586,N_1468,N_1219);
or U1587 (N_1587,N_861,N_1216);
nand U1588 (N_1588,N_1055,N_1287);
nand U1589 (N_1589,N_857,N_1134);
nor U1590 (N_1590,N_1469,N_1441);
or U1591 (N_1591,N_885,N_1113);
nand U1592 (N_1592,N_798,N_1285);
nand U1593 (N_1593,N_1234,N_1230);
or U1594 (N_1594,N_1240,N_1112);
and U1595 (N_1595,N_918,N_1476);
and U1596 (N_1596,N_1381,N_1141);
and U1597 (N_1597,N_1377,N_1120);
and U1598 (N_1598,N_1269,N_1470);
and U1599 (N_1599,N_1182,N_1367);
nand U1600 (N_1600,N_1306,N_809);
and U1601 (N_1601,N_829,N_1027);
nor U1602 (N_1602,N_1158,N_1076);
nand U1603 (N_1603,N_1316,N_1396);
or U1604 (N_1604,N_1071,N_1427);
nand U1605 (N_1605,N_781,N_949);
nor U1606 (N_1606,N_1277,N_986);
nor U1607 (N_1607,N_1179,N_881);
and U1608 (N_1608,N_1389,N_1005);
or U1609 (N_1609,N_1482,N_1457);
or U1610 (N_1610,N_1442,N_1207);
nor U1611 (N_1611,N_783,N_1352);
and U1612 (N_1612,N_1006,N_1242);
or U1613 (N_1613,N_1284,N_754);
nor U1614 (N_1614,N_1447,N_928);
nand U1615 (N_1615,N_805,N_1139);
and U1616 (N_1616,N_1320,N_1364);
or U1617 (N_1617,N_1245,N_944);
and U1618 (N_1618,N_1183,N_866);
nand U1619 (N_1619,N_1018,N_875);
nor U1620 (N_1620,N_1210,N_1154);
nand U1621 (N_1621,N_899,N_779);
nand U1622 (N_1622,N_1106,N_1357);
or U1623 (N_1623,N_1228,N_1450);
nand U1624 (N_1624,N_750,N_1178);
nand U1625 (N_1625,N_1355,N_1478);
nand U1626 (N_1626,N_854,N_1221);
or U1627 (N_1627,N_792,N_760);
and U1628 (N_1628,N_790,N_1117);
nor U1629 (N_1629,N_1308,N_1128);
nand U1630 (N_1630,N_1414,N_946);
or U1631 (N_1631,N_990,N_883);
nand U1632 (N_1632,N_1058,N_1385);
nand U1633 (N_1633,N_1265,N_876);
nor U1634 (N_1634,N_1078,N_1486);
and U1635 (N_1635,N_1252,N_1091);
nand U1636 (N_1636,N_1098,N_1193);
nand U1637 (N_1637,N_1209,N_1433);
or U1638 (N_1638,N_810,N_1037);
and U1639 (N_1639,N_960,N_1267);
nand U1640 (N_1640,N_1021,N_1383);
or U1641 (N_1641,N_761,N_982);
or U1642 (N_1642,N_770,N_1250);
and U1643 (N_1643,N_1356,N_816);
and U1644 (N_1644,N_1057,N_886);
nand U1645 (N_1645,N_948,N_897);
or U1646 (N_1646,N_777,N_1132);
and U1647 (N_1647,N_1477,N_1496);
and U1648 (N_1648,N_965,N_1218);
nor U1649 (N_1649,N_811,N_894);
nor U1650 (N_1650,N_1048,N_1417);
nand U1651 (N_1651,N_1424,N_772);
nor U1652 (N_1652,N_985,N_1399);
or U1653 (N_1653,N_1013,N_1390);
nor U1654 (N_1654,N_1151,N_1226);
nor U1655 (N_1655,N_882,N_1499);
and U1656 (N_1656,N_1303,N_1175);
nand U1657 (N_1657,N_922,N_1146);
nand U1658 (N_1658,N_812,N_955);
nor U1659 (N_1659,N_1463,N_891);
nor U1660 (N_1660,N_1149,N_793);
nor U1661 (N_1661,N_1163,N_1452);
or U1662 (N_1662,N_1368,N_1379);
and U1663 (N_1663,N_1394,N_1366);
nor U1664 (N_1664,N_1294,N_1046);
or U1665 (N_1665,N_929,N_1434);
nand U1666 (N_1666,N_1426,N_1266);
nand U1667 (N_1667,N_1203,N_1405);
and U1668 (N_1668,N_1080,N_767);
and U1669 (N_1669,N_887,N_788);
and U1670 (N_1670,N_1090,N_1089);
nor U1671 (N_1671,N_878,N_1431);
nor U1672 (N_1672,N_755,N_981);
and U1673 (N_1673,N_974,N_1187);
or U1674 (N_1674,N_1346,N_1343);
or U1675 (N_1675,N_998,N_1129);
and U1676 (N_1676,N_968,N_1438);
nand U1677 (N_1677,N_766,N_1291);
nand U1678 (N_1678,N_1264,N_1028);
nor U1679 (N_1679,N_1096,N_1192);
and U1680 (N_1680,N_1429,N_1166);
nor U1681 (N_1681,N_794,N_1196);
or U1682 (N_1682,N_945,N_1305);
and U1683 (N_1683,N_1177,N_836);
and U1684 (N_1684,N_958,N_1236);
or U1685 (N_1685,N_1081,N_1025);
or U1686 (N_1686,N_935,N_1448);
nor U1687 (N_1687,N_1280,N_1064);
and U1688 (N_1688,N_824,N_801);
nand U1689 (N_1689,N_1413,N_890);
nor U1690 (N_1690,N_1073,N_822);
nor U1691 (N_1691,N_880,N_1404);
nand U1692 (N_1692,N_1238,N_1035);
and U1693 (N_1693,N_1092,N_1329);
nand U1694 (N_1694,N_1231,N_1391);
nand U1695 (N_1695,N_859,N_889);
or U1696 (N_1696,N_799,N_1130);
nand U1697 (N_1697,N_1436,N_1194);
or U1698 (N_1698,N_987,N_1087);
nor U1699 (N_1699,N_1310,N_994);
nor U1700 (N_1700,N_802,N_1145);
or U1701 (N_1701,N_1215,N_905);
or U1702 (N_1702,N_997,N_1023);
nor U1703 (N_1703,N_877,N_1045);
nor U1704 (N_1704,N_1459,N_1016);
nand U1705 (N_1705,N_1030,N_1204);
and U1706 (N_1706,N_873,N_1446);
or U1707 (N_1707,N_1085,N_1392);
nor U1708 (N_1708,N_1173,N_1286);
nand U1709 (N_1709,N_1189,N_785);
or U1710 (N_1710,N_1041,N_1492);
nor U1711 (N_1711,N_1020,N_782);
or U1712 (N_1712,N_1107,N_1127);
nor U1713 (N_1713,N_884,N_1327);
or U1714 (N_1714,N_1165,N_1313);
nor U1715 (N_1715,N_1388,N_1359);
nor U1716 (N_1716,N_1168,N_1222);
or U1717 (N_1717,N_1188,N_902);
nand U1718 (N_1718,N_757,N_1349);
nor U1719 (N_1719,N_1015,N_1102);
and U1720 (N_1720,N_914,N_1105);
nor U1721 (N_1721,N_1202,N_1493);
or U1722 (N_1722,N_1317,N_1062);
or U1723 (N_1723,N_776,N_839);
nor U1724 (N_1724,N_940,N_874);
and U1725 (N_1725,N_983,N_1094);
nor U1726 (N_1726,N_828,N_1297);
and U1727 (N_1727,N_1032,N_1323);
nand U1728 (N_1728,N_971,N_1491);
and U1729 (N_1729,N_904,N_1049);
and U1730 (N_1730,N_759,N_1206);
and U1731 (N_1731,N_1347,N_1012);
and U1732 (N_1732,N_1325,N_1418);
nor U1733 (N_1733,N_1000,N_814);
or U1734 (N_1734,N_1440,N_1156);
and U1735 (N_1735,N_838,N_1268);
and U1736 (N_1736,N_919,N_773);
nand U1737 (N_1737,N_758,N_1225);
nor U1738 (N_1738,N_1407,N_862);
nand U1739 (N_1739,N_1011,N_1116);
nand U1740 (N_1740,N_1462,N_1402);
nor U1741 (N_1741,N_1254,N_813);
or U1742 (N_1742,N_1257,N_1109);
nand U1743 (N_1743,N_1246,N_1373);
nand U1744 (N_1744,N_1002,N_1033);
or U1745 (N_1745,N_1232,N_1001);
and U1746 (N_1746,N_1147,N_1494);
nor U1747 (N_1747,N_977,N_975);
and U1748 (N_1748,N_1208,N_909);
and U1749 (N_1749,N_1365,N_1481);
or U1750 (N_1750,N_1153,N_1155);
nand U1751 (N_1751,N_1449,N_1487);
or U1752 (N_1752,N_1299,N_1467);
and U1753 (N_1753,N_1401,N_1184);
nand U1754 (N_1754,N_910,N_1263);
nor U1755 (N_1755,N_1176,N_1022);
nor U1756 (N_1756,N_1122,N_751);
xor U1757 (N_1757,N_1233,N_1161);
and U1758 (N_1758,N_806,N_1271);
nand U1759 (N_1759,N_936,N_1198);
nor U1760 (N_1760,N_1133,N_860);
nor U1761 (N_1761,N_892,N_1053);
and U1762 (N_1762,N_1111,N_1051);
and U1763 (N_1763,N_1292,N_834);
and U1764 (N_1764,N_953,N_858);
nor U1765 (N_1765,N_970,N_1162);
or U1766 (N_1766,N_1353,N_1077);
and U1767 (N_1767,N_763,N_830);
nor U1768 (N_1768,N_888,N_795);
or U1769 (N_1769,N_1382,N_1164);
nor U1770 (N_1770,N_1422,N_1298);
nor U1771 (N_1771,N_1393,N_843);
or U1772 (N_1772,N_1458,N_1065);
or U1773 (N_1773,N_1328,N_924);
nand U1774 (N_1774,N_1339,N_926);
nand U1775 (N_1775,N_784,N_1318);
nand U1776 (N_1776,N_921,N_1495);
or U1777 (N_1777,N_815,N_835);
nand U1778 (N_1778,N_1110,N_797);
nor U1779 (N_1779,N_1060,N_1301);
and U1780 (N_1780,N_1047,N_947);
nor U1781 (N_1781,N_1103,N_1369);
nand U1782 (N_1782,N_1474,N_1324);
or U1783 (N_1783,N_807,N_1361);
and U1784 (N_1784,N_972,N_1029);
or U1785 (N_1785,N_847,N_933);
and U1786 (N_1786,N_831,N_1197);
or U1787 (N_1787,N_1119,N_775);
and U1788 (N_1788,N_1437,N_1278);
or U1789 (N_1789,N_1137,N_1259);
or U1790 (N_1790,N_1061,N_1472);
or U1791 (N_1791,N_1300,N_1262);
nor U1792 (N_1792,N_1425,N_989);
or U1793 (N_1793,N_1372,N_1443);
nand U1794 (N_1794,N_1010,N_1059);
or U1795 (N_1795,N_1453,N_913);
xor U1796 (N_1796,N_1354,N_1430);
and U1797 (N_1797,N_1340,N_1056);
or U1798 (N_1798,N_988,N_1386);
nand U1799 (N_1799,N_1211,N_1319);
and U1800 (N_1800,N_1143,N_1345);
and U1801 (N_1801,N_1321,N_951);
nand U1802 (N_1802,N_1074,N_1326);
nand U1803 (N_1803,N_1082,N_954);
nor U1804 (N_1804,N_1088,N_993);
nand U1805 (N_1805,N_1160,N_1159);
nand U1806 (N_1806,N_1104,N_1069);
nand U1807 (N_1807,N_1304,N_1124);
nand U1808 (N_1808,N_1050,N_992);
nor U1809 (N_1809,N_1408,N_896);
or U1810 (N_1810,N_1400,N_1171);
nand U1811 (N_1811,N_1490,N_1471);
and U1812 (N_1812,N_1387,N_768);
nor U1813 (N_1813,N_1200,N_856);
or U1814 (N_1814,N_1007,N_1295);
or U1815 (N_1815,N_1334,N_1275);
or U1816 (N_1816,N_1118,N_832);
nand U1817 (N_1817,N_1488,N_939);
or U1818 (N_1818,N_1480,N_1042);
nand U1819 (N_1819,N_973,N_1350);
or U1820 (N_1820,N_941,N_1070);
and U1821 (N_1821,N_753,N_825);
nor U1822 (N_1822,N_906,N_1439);
and U1823 (N_1823,N_803,N_1126);
and U1824 (N_1824,N_1170,N_1260);
or U1825 (N_1825,N_1167,N_1008);
and U1826 (N_1826,N_923,N_1395);
and U1827 (N_1827,N_1114,N_963);
nor U1828 (N_1828,N_1123,N_932);
nor U1829 (N_1829,N_1144,N_1362);
or U1830 (N_1830,N_1360,N_1072);
and U1831 (N_1831,N_1281,N_1024);
nand U1832 (N_1832,N_1344,N_916);
or U1833 (N_1833,N_1358,N_762);
and U1834 (N_1834,N_1017,N_1054);
and U1835 (N_1835,N_1214,N_765);
nor U1836 (N_1836,N_821,N_1333);
nor U1837 (N_1837,N_1213,N_769);
nand U1838 (N_1838,N_1239,N_756);
nand U1839 (N_1839,N_1086,N_995);
and U1840 (N_1840,N_1142,N_1282);
and U1841 (N_1841,N_950,N_1322);
or U1842 (N_1842,N_818,N_867);
and U1843 (N_1843,N_1201,N_840);
nor U1844 (N_1844,N_931,N_764);
or U1845 (N_1845,N_1199,N_956);
nand U1846 (N_1846,N_1406,N_1212);
or U1847 (N_1847,N_1067,N_1337);
and U1848 (N_1848,N_819,N_1157);
nor U1849 (N_1849,N_942,N_752);
nand U1850 (N_1850,N_865,N_1371);
nand U1851 (N_1851,N_980,N_1040);
or U1852 (N_1852,N_978,N_1108);
or U1853 (N_1853,N_1244,N_1003);
or U1854 (N_1854,N_1138,N_1419);
nor U1855 (N_1855,N_1351,N_1099);
and U1856 (N_1856,N_872,N_1100);
or U1857 (N_1857,N_962,N_1227);
or U1858 (N_1858,N_800,N_1497);
or U1859 (N_1859,N_912,N_961);
and U1860 (N_1860,N_930,N_957);
nor U1861 (N_1861,N_1241,N_1464);
nor U1862 (N_1862,N_841,N_1290);
or U1863 (N_1863,N_915,N_979);
or U1864 (N_1864,N_967,N_1075);
or U1865 (N_1865,N_863,N_774);
or U1866 (N_1866,N_1195,N_1485);
nor U1867 (N_1867,N_1169,N_1031);
and U1868 (N_1868,N_1411,N_1296);
or U1869 (N_1869,N_938,N_1348);
or U1870 (N_1870,N_898,N_852);
and U1871 (N_1871,N_1374,N_1461);
or U1872 (N_1872,N_1185,N_1307);
nor U1873 (N_1873,N_1186,N_1190);
and U1874 (N_1874,N_853,N_1038);
nand U1875 (N_1875,N_1388,N_953);
or U1876 (N_1876,N_1016,N_758);
or U1877 (N_1877,N_989,N_930);
and U1878 (N_1878,N_1072,N_808);
or U1879 (N_1879,N_1360,N_1052);
nand U1880 (N_1880,N_1290,N_1114);
nor U1881 (N_1881,N_865,N_970);
nor U1882 (N_1882,N_1293,N_1152);
nor U1883 (N_1883,N_1097,N_998);
nand U1884 (N_1884,N_1065,N_936);
nor U1885 (N_1885,N_806,N_1426);
and U1886 (N_1886,N_1284,N_1110);
and U1887 (N_1887,N_855,N_1313);
or U1888 (N_1888,N_865,N_1104);
or U1889 (N_1889,N_775,N_1180);
or U1890 (N_1890,N_1041,N_840);
nand U1891 (N_1891,N_797,N_845);
nor U1892 (N_1892,N_1096,N_1010);
and U1893 (N_1893,N_876,N_1473);
and U1894 (N_1894,N_1102,N_795);
nand U1895 (N_1895,N_1301,N_1454);
nor U1896 (N_1896,N_1183,N_1348);
or U1897 (N_1897,N_1447,N_912);
and U1898 (N_1898,N_1176,N_1330);
nor U1899 (N_1899,N_1077,N_1258);
nand U1900 (N_1900,N_1226,N_1350);
nand U1901 (N_1901,N_1415,N_1225);
nand U1902 (N_1902,N_1460,N_928);
nor U1903 (N_1903,N_872,N_1016);
and U1904 (N_1904,N_1459,N_809);
nand U1905 (N_1905,N_816,N_1242);
and U1906 (N_1906,N_1245,N_754);
nor U1907 (N_1907,N_1216,N_1070);
and U1908 (N_1908,N_889,N_831);
or U1909 (N_1909,N_1147,N_889);
nor U1910 (N_1910,N_1002,N_820);
nand U1911 (N_1911,N_798,N_871);
nor U1912 (N_1912,N_1015,N_1237);
nor U1913 (N_1913,N_1260,N_979);
nand U1914 (N_1914,N_1254,N_1111);
nand U1915 (N_1915,N_1242,N_1157);
nor U1916 (N_1916,N_990,N_853);
nor U1917 (N_1917,N_1441,N_1072);
nand U1918 (N_1918,N_1380,N_1050);
nand U1919 (N_1919,N_914,N_890);
or U1920 (N_1920,N_1174,N_843);
nor U1921 (N_1921,N_1337,N_1342);
and U1922 (N_1922,N_857,N_1184);
nand U1923 (N_1923,N_1219,N_905);
nor U1924 (N_1924,N_1353,N_935);
or U1925 (N_1925,N_1177,N_1433);
nand U1926 (N_1926,N_843,N_809);
or U1927 (N_1927,N_978,N_1171);
and U1928 (N_1928,N_1286,N_1255);
or U1929 (N_1929,N_1418,N_1028);
nor U1930 (N_1930,N_1283,N_1366);
nand U1931 (N_1931,N_1269,N_1299);
and U1932 (N_1932,N_1272,N_1321);
nor U1933 (N_1933,N_768,N_1100);
or U1934 (N_1934,N_829,N_951);
or U1935 (N_1935,N_1111,N_806);
nor U1936 (N_1936,N_761,N_1055);
or U1937 (N_1937,N_1198,N_1074);
and U1938 (N_1938,N_1346,N_828);
or U1939 (N_1939,N_1404,N_1225);
or U1940 (N_1940,N_1106,N_1156);
and U1941 (N_1941,N_1182,N_910);
nand U1942 (N_1942,N_990,N_1119);
nor U1943 (N_1943,N_1483,N_1130);
and U1944 (N_1944,N_1439,N_1054);
nor U1945 (N_1945,N_1307,N_1119);
and U1946 (N_1946,N_1410,N_792);
and U1947 (N_1947,N_996,N_1329);
nand U1948 (N_1948,N_1117,N_800);
nand U1949 (N_1949,N_1127,N_1497);
and U1950 (N_1950,N_1236,N_1016);
or U1951 (N_1951,N_1493,N_982);
nand U1952 (N_1952,N_1021,N_1443);
and U1953 (N_1953,N_1335,N_1248);
nand U1954 (N_1954,N_800,N_1241);
and U1955 (N_1955,N_1211,N_950);
and U1956 (N_1956,N_921,N_1177);
nand U1957 (N_1957,N_1247,N_862);
nand U1958 (N_1958,N_1268,N_1235);
nand U1959 (N_1959,N_1491,N_1492);
and U1960 (N_1960,N_775,N_1204);
nor U1961 (N_1961,N_1103,N_978);
nor U1962 (N_1962,N_958,N_1312);
or U1963 (N_1963,N_1184,N_1196);
nand U1964 (N_1964,N_1483,N_1306);
or U1965 (N_1965,N_1314,N_775);
nand U1966 (N_1966,N_1431,N_1225);
and U1967 (N_1967,N_1259,N_1155);
nor U1968 (N_1968,N_767,N_1089);
and U1969 (N_1969,N_922,N_1496);
and U1970 (N_1970,N_1424,N_1328);
nand U1971 (N_1971,N_996,N_1230);
nor U1972 (N_1972,N_1107,N_1317);
and U1973 (N_1973,N_785,N_979);
nor U1974 (N_1974,N_1392,N_1208);
or U1975 (N_1975,N_1412,N_785);
or U1976 (N_1976,N_958,N_1168);
and U1977 (N_1977,N_810,N_1498);
nor U1978 (N_1978,N_812,N_1060);
or U1979 (N_1979,N_756,N_1236);
nand U1980 (N_1980,N_1142,N_815);
and U1981 (N_1981,N_1162,N_1361);
nor U1982 (N_1982,N_1187,N_1006);
nor U1983 (N_1983,N_1465,N_1449);
nor U1984 (N_1984,N_1294,N_767);
or U1985 (N_1985,N_1076,N_1365);
nand U1986 (N_1986,N_1373,N_910);
nand U1987 (N_1987,N_1182,N_1236);
nand U1988 (N_1988,N_923,N_920);
and U1989 (N_1989,N_991,N_1396);
or U1990 (N_1990,N_1335,N_1119);
nor U1991 (N_1991,N_1217,N_1321);
nand U1992 (N_1992,N_1274,N_1022);
or U1993 (N_1993,N_1191,N_1240);
nor U1994 (N_1994,N_1098,N_1427);
nand U1995 (N_1995,N_911,N_976);
nand U1996 (N_1996,N_1173,N_1395);
nand U1997 (N_1997,N_801,N_1111);
or U1998 (N_1998,N_1015,N_898);
or U1999 (N_1999,N_1219,N_1318);
and U2000 (N_2000,N_1450,N_813);
nor U2001 (N_2001,N_1294,N_1000);
and U2002 (N_2002,N_1080,N_795);
nand U2003 (N_2003,N_783,N_1300);
or U2004 (N_2004,N_1090,N_947);
nand U2005 (N_2005,N_1223,N_794);
nor U2006 (N_2006,N_853,N_1204);
nor U2007 (N_2007,N_1305,N_1084);
and U2008 (N_2008,N_938,N_1497);
nand U2009 (N_2009,N_1137,N_786);
and U2010 (N_2010,N_1473,N_1428);
and U2011 (N_2011,N_849,N_1405);
and U2012 (N_2012,N_887,N_1056);
and U2013 (N_2013,N_1020,N_1111);
and U2014 (N_2014,N_1488,N_1088);
nor U2015 (N_2015,N_1158,N_784);
nor U2016 (N_2016,N_1041,N_1209);
and U2017 (N_2017,N_1283,N_1168);
and U2018 (N_2018,N_1458,N_1055);
and U2019 (N_2019,N_1139,N_1411);
xnor U2020 (N_2020,N_850,N_1054);
nand U2021 (N_2021,N_1161,N_1277);
or U2022 (N_2022,N_903,N_1339);
nor U2023 (N_2023,N_1485,N_1232);
nor U2024 (N_2024,N_1073,N_800);
and U2025 (N_2025,N_940,N_1334);
or U2026 (N_2026,N_1352,N_1400);
nor U2027 (N_2027,N_1458,N_831);
nand U2028 (N_2028,N_1411,N_1077);
nand U2029 (N_2029,N_1116,N_948);
or U2030 (N_2030,N_1049,N_1479);
and U2031 (N_2031,N_819,N_832);
nand U2032 (N_2032,N_806,N_771);
nor U2033 (N_2033,N_785,N_1019);
or U2034 (N_2034,N_1247,N_1117);
and U2035 (N_2035,N_958,N_1058);
nand U2036 (N_2036,N_821,N_1495);
or U2037 (N_2037,N_1318,N_1326);
and U2038 (N_2038,N_921,N_1116);
nor U2039 (N_2039,N_1087,N_903);
or U2040 (N_2040,N_1374,N_1211);
nor U2041 (N_2041,N_1025,N_1200);
nor U2042 (N_2042,N_952,N_1356);
or U2043 (N_2043,N_1169,N_1445);
nor U2044 (N_2044,N_839,N_750);
nand U2045 (N_2045,N_1267,N_1099);
or U2046 (N_2046,N_1077,N_924);
and U2047 (N_2047,N_826,N_765);
and U2048 (N_2048,N_1458,N_1279);
nand U2049 (N_2049,N_1275,N_825);
nor U2050 (N_2050,N_1303,N_1387);
nand U2051 (N_2051,N_1125,N_1439);
or U2052 (N_2052,N_1134,N_1414);
nand U2053 (N_2053,N_1403,N_854);
nand U2054 (N_2054,N_1276,N_1053);
nand U2055 (N_2055,N_1468,N_1067);
nor U2056 (N_2056,N_997,N_1129);
and U2057 (N_2057,N_1172,N_807);
nand U2058 (N_2058,N_1471,N_976);
or U2059 (N_2059,N_1228,N_787);
and U2060 (N_2060,N_1185,N_974);
nor U2061 (N_2061,N_928,N_894);
nor U2062 (N_2062,N_1068,N_1266);
nand U2063 (N_2063,N_795,N_1029);
and U2064 (N_2064,N_997,N_1337);
nand U2065 (N_2065,N_862,N_880);
and U2066 (N_2066,N_1159,N_1177);
or U2067 (N_2067,N_1466,N_967);
and U2068 (N_2068,N_1231,N_786);
nand U2069 (N_2069,N_1335,N_1055);
and U2070 (N_2070,N_1391,N_1076);
nor U2071 (N_2071,N_829,N_874);
nor U2072 (N_2072,N_878,N_896);
or U2073 (N_2073,N_1324,N_1073);
and U2074 (N_2074,N_1241,N_930);
or U2075 (N_2075,N_1310,N_1238);
nor U2076 (N_2076,N_949,N_1129);
nor U2077 (N_2077,N_1188,N_927);
nor U2078 (N_2078,N_1430,N_834);
or U2079 (N_2079,N_1052,N_904);
or U2080 (N_2080,N_991,N_901);
and U2081 (N_2081,N_862,N_1473);
nand U2082 (N_2082,N_882,N_831);
or U2083 (N_2083,N_877,N_1185);
nand U2084 (N_2084,N_1308,N_1018);
or U2085 (N_2085,N_1410,N_1278);
and U2086 (N_2086,N_764,N_1479);
nor U2087 (N_2087,N_933,N_953);
nor U2088 (N_2088,N_998,N_1482);
nand U2089 (N_2089,N_1363,N_1027);
nor U2090 (N_2090,N_988,N_1326);
and U2091 (N_2091,N_1192,N_832);
nand U2092 (N_2092,N_1258,N_1031);
nand U2093 (N_2093,N_1362,N_895);
and U2094 (N_2094,N_1187,N_772);
nand U2095 (N_2095,N_1362,N_1230);
nand U2096 (N_2096,N_1241,N_1176);
nor U2097 (N_2097,N_923,N_811);
nand U2098 (N_2098,N_1048,N_992);
nor U2099 (N_2099,N_873,N_1395);
or U2100 (N_2100,N_1280,N_884);
or U2101 (N_2101,N_1372,N_808);
nor U2102 (N_2102,N_1180,N_1010);
nor U2103 (N_2103,N_847,N_1019);
nor U2104 (N_2104,N_909,N_1361);
and U2105 (N_2105,N_1298,N_1477);
nor U2106 (N_2106,N_1201,N_1425);
or U2107 (N_2107,N_1397,N_1306);
and U2108 (N_2108,N_1343,N_797);
and U2109 (N_2109,N_938,N_1251);
nand U2110 (N_2110,N_980,N_954);
nand U2111 (N_2111,N_1096,N_1348);
nor U2112 (N_2112,N_1451,N_1023);
and U2113 (N_2113,N_1329,N_1284);
nand U2114 (N_2114,N_945,N_1324);
nand U2115 (N_2115,N_1351,N_1004);
nand U2116 (N_2116,N_1031,N_894);
nand U2117 (N_2117,N_1029,N_1427);
or U2118 (N_2118,N_1324,N_1298);
nand U2119 (N_2119,N_1032,N_1132);
or U2120 (N_2120,N_888,N_1178);
and U2121 (N_2121,N_1016,N_1008);
nand U2122 (N_2122,N_829,N_1351);
or U2123 (N_2123,N_1035,N_1458);
and U2124 (N_2124,N_914,N_1497);
nand U2125 (N_2125,N_1103,N_917);
or U2126 (N_2126,N_1242,N_1021);
and U2127 (N_2127,N_953,N_983);
nor U2128 (N_2128,N_1477,N_798);
nor U2129 (N_2129,N_894,N_799);
or U2130 (N_2130,N_1277,N_1010);
nand U2131 (N_2131,N_783,N_1382);
or U2132 (N_2132,N_1170,N_1335);
or U2133 (N_2133,N_1409,N_1178);
or U2134 (N_2134,N_1331,N_986);
or U2135 (N_2135,N_1285,N_1149);
or U2136 (N_2136,N_956,N_1176);
nand U2137 (N_2137,N_877,N_1059);
nand U2138 (N_2138,N_1234,N_1326);
nor U2139 (N_2139,N_1446,N_1327);
nand U2140 (N_2140,N_1017,N_1297);
nand U2141 (N_2141,N_879,N_1340);
nand U2142 (N_2142,N_1233,N_1073);
nand U2143 (N_2143,N_1385,N_1042);
or U2144 (N_2144,N_1062,N_1261);
and U2145 (N_2145,N_1383,N_987);
nand U2146 (N_2146,N_1485,N_826);
and U2147 (N_2147,N_1167,N_1493);
nand U2148 (N_2148,N_1433,N_1455);
or U2149 (N_2149,N_1461,N_919);
xnor U2150 (N_2150,N_1306,N_898);
nand U2151 (N_2151,N_1380,N_1353);
nand U2152 (N_2152,N_1270,N_1311);
nor U2153 (N_2153,N_1175,N_1449);
or U2154 (N_2154,N_837,N_916);
or U2155 (N_2155,N_1436,N_1308);
and U2156 (N_2156,N_1339,N_1324);
nand U2157 (N_2157,N_831,N_1161);
nand U2158 (N_2158,N_1401,N_947);
nor U2159 (N_2159,N_1095,N_1360);
or U2160 (N_2160,N_912,N_920);
nor U2161 (N_2161,N_1306,N_1320);
nand U2162 (N_2162,N_1371,N_892);
nand U2163 (N_2163,N_1113,N_1216);
nand U2164 (N_2164,N_1187,N_1438);
nand U2165 (N_2165,N_853,N_1147);
nand U2166 (N_2166,N_1282,N_1182);
and U2167 (N_2167,N_909,N_954);
nand U2168 (N_2168,N_1031,N_964);
nor U2169 (N_2169,N_1298,N_1465);
and U2170 (N_2170,N_1066,N_1347);
and U2171 (N_2171,N_1387,N_985);
or U2172 (N_2172,N_1227,N_1285);
or U2173 (N_2173,N_1299,N_902);
or U2174 (N_2174,N_776,N_1343);
nor U2175 (N_2175,N_1379,N_1208);
or U2176 (N_2176,N_1150,N_1006);
and U2177 (N_2177,N_768,N_1203);
or U2178 (N_2178,N_1245,N_1431);
and U2179 (N_2179,N_1327,N_1461);
and U2180 (N_2180,N_773,N_1440);
nand U2181 (N_2181,N_1094,N_943);
or U2182 (N_2182,N_1362,N_1285);
or U2183 (N_2183,N_1214,N_1487);
nor U2184 (N_2184,N_1180,N_1464);
or U2185 (N_2185,N_789,N_1067);
xor U2186 (N_2186,N_803,N_779);
and U2187 (N_2187,N_1008,N_1087);
nor U2188 (N_2188,N_1465,N_899);
nand U2189 (N_2189,N_1491,N_1117);
and U2190 (N_2190,N_1397,N_1003);
and U2191 (N_2191,N_1360,N_1338);
and U2192 (N_2192,N_835,N_752);
or U2193 (N_2193,N_1385,N_1429);
and U2194 (N_2194,N_758,N_785);
nand U2195 (N_2195,N_796,N_1344);
nor U2196 (N_2196,N_1419,N_967);
nor U2197 (N_2197,N_867,N_1280);
and U2198 (N_2198,N_1105,N_1200);
nand U2199 (N_2199,N_958,N_813);
nor U2200 (N_2200,N_1484,N_875);
and U2201 (N_2201,N_1356,N_959);
and U2202 (N_2202,N_1047,N_1192);
or U2203 (N_2203,N_843,N_937);
nor U2204 (N_2204,N_776,N_1499);
nand U2205 (N_2205,N_945,N_827);
or U2206 (N_2206,N_1020,N_1086);
and U2207 (N_2207,N_1417,N_767);
and U2208 (N_2208,N_1027,N_775);
or U2209 (N_2209,N_827,N_1047);
or U2210 (N_2210,N_1481,N_778);
or U2211 (N_2211,N_972,N_1441);
and U2212 (N_2212,N_1012,N_866);
and U2213 (N_2213,N_1152,N_799);
nand U2214 (N_2214,N_791,N_1205);
and U2215 (N_2215,N_825,N_1093);
nor U2216 (N_2216,N_1433,N_1340);
nand U2217 (N_2217,N_1350,N_1348);
nor U2218 (N_2218,N_949,N_1283);
or U2219 (N_2219,N_1232,N_962);
or U2220 (N_2220,N_1219,N_1231);
and U2221 (N_2221,N_1497,N_1356);
nor U2222 (N_2222,N_1269,N_1289);
and U2223 (N_2223,N_1111,N_778);
and U2224 (N_2224,N_1078,N_1438);
xor U2225 (N_2225,N_1015,N_1070);
and U2226 (N_2226,N_1430,N_926);
and U2227 (N_2227,N_1121,N_1438);
nand U2228 (N_2228,N_943,N_1400);
nor U2229 (N_2229,N_1222,N_1127);
or U2230 (N_2230,N_1187,N_1193);
and U2231 (N_2231,N_900,N_809);
or U2232 (N_2232,N_1048,N_882);
or U2233 (N_2233,N_1208,N_964);
nand U2234 (N_2234,N_1043,N_924);
and U2235 (N_2235,N_1216,N_830);
and U2236 (N_2236,N_1053,N_751);
nor U2237 (N_2237,N_1377,N_1422);
and U2238 (N_2238,N_1343,N_1409);
nand U2239 (N_2239,N_1020,N_877);
and U2240 (N_2240,N_1483,N_1360);
and U2241 (N_2241,N_1212,N_1416);
nor U2242 (N_2242,N_987,N_1487);
or U2243 (N_2243,N_889,N_953);
nor U2244 (N_2244,N_1225,N_944);
nor U2245 (N_2245,N_856,N_1211);
nand U2246 (N_2246,N_1397,N_1443);
and U2247 (N_2247,N_784,N_1057);
nor U2248 (N_2248,N_1360,N_1327);
nand U2249 (N_2249,N_1166,N_881);
nor U2250 (N_2250,N_2220,N_2155);
or U2251 (N_2251,N_2199,N_2017);
nand U2252 (N_2252,N_1975,N_1803);
or U2253 (N_2253,N_1525,N_2119);
or U2254 (N_2254,N_1606,N_1514);
or U2255 (N_2255,N_2018,N_1519);
and U2256 (N_2256,N_1729,N_2133);
nor U2257 (N_2257,N_2198,N_1875);
or U2258 (N_2258,N_1566,N_2048);
or U2259 (N_2259,N_2177,N_2137);
or U2260 (N_2260,N_1882,N_1716);
nor U2261 (N_2261,N_1911,N_1705);
nor U2262 (N_2262,N_1877,N_1786);
and U2263 (N_2263,N_2229,N_2062);
and U2264 (N_2264,N_1662,N_2011);
or U2265 (N_2265,N_1778,N_1634);
and U2266 (N_2266,N_2158,N_1874);
nand U2267 (N_2267,N_1502,N_1790);
or U2268 (N_2268,N_2125,N_1869);
nor U2269 (N_2269,N_2073,N_1799);
and U2270 (N_2270,N_1657,N_1533);
or U2271 (N_2271,N_2047,N_1629);
or U2272 (N_2272,N_1542,N_1596);
nor U2273 (N_2273,N_2077,N_1810);
and U2274 (N_2274,N_2214,N_2203);
or U2275 (N_2275,N_1859,N_1547);
and U2276 (N_2276,N_1850,N_1912);
nor U2277 (N_2277,N_2036,N_1749);
nor U2278 (N_2278,N_1954,N_1726);
nand U2279 (N_2279,N_2098,N_1936);
nor U2280 (N_2280,N_1956,N_2081);
nor U2281 (N_2281,N_1658,N_2103);
nand U2282 (N_2282,N_1938,N_2218);
nor U2283 (N_2283,N_2102,N_2222);
nand U2284 (N_2284,N_1955,N_1913);
nand U2285 (N_2285,N_2149,N_2106);
and U2286 (N_2286,N_1709,N_1905);
nor U2287 (N_2287,N_1844,N_2070);
and U2288 (N_2288,N_1500,N_2023);
or U2289 (N_2289,N_1993,N_2019);
nor U2290 (N_2290,N_1899,N_1550);
nor U2291 (N_2291,N_1903,N_1967);
and U2292 (N_2292,N_2215,N_2246);
nand U2293 (N_2293,N_1765,N_1871);
nor U2294 (N_2294,N_1628,N_2108);
nand U2295 (N_2295,N_1605,N_1694);
and U2296 (N_2296,N_1898,N_1923);
nand U2297 (N_2297,N_1641,N_2110);
and U2298 (N_2298,N_1666,N_1580);
nor U2299 (N_2299,N_1696,N_1679);
nor U2300 (N_2300,N_2207,N_2052);
and U2301 (N_2301,N_1536,N_1977);
or U2302 (N_2302,N_1782,N_1623);
and U2303 (N_2303,N_2156,N_1663);
nor U2304 (N_2304,N_1949,N_2117);
nor U2305 (N_2305,N_1681,N_1867);
nor U2306 (N_2306,N_2049,N_2020);
nand U2307 (N_2307,N_1981,N_1573);
or U2308 (N_2308,N_1991,N_1767);
nor U2309 (N_2309,N_1702,N_1831);
and U2310 (N_2310,N_2151,N_2208);
and U2311 (N_2311,N_2058,N_1785);
nor U2312 (N_2312,N_2170,N_1581);
nor U2313 (N_2313,N_2094,N_1748);
nand U2314 (N_2314,N_2244,N_2140);
and U2315 (N_2315,N_1801,N_1939);
nor U2316 (N_2316,N_2076,N_1650);
or U2317 (N_2317,N_1644,N_2172);
nor U2318 (N_2318,N_1540,N_2135);
or U2319 (N_2319,N_1910,N_1558);
nand U2320 (N_2320,N_1529,N_1538);
nand U2321 (N_2321,N_1675,N_1703);
nor U2322 (N_2322,N_2056,N_1612);
and U2323 (N_2323,N_2233,N_2061);
and U2324 (N_2324,N_2004,N_2153);
or U2325 (N_2325,N_1753,N_1659);
or U2326 (N_2326,N_2211,N_2118);
nand U2327 (N_2327,N_1548,N_1597);
and U2328 (N_2328,N_2189,N_1793);
and U2329 (N_2329,N_2029,N_1892);
or U2330 (N_2330,N_2114,N_1611);
or U2331 (N_2331,N_1562,N_1523);
or U2332 (N_2332,N_1928,N_2184);
nor U2333 (N_2333,N_1860,N_1673);
nor U2334 (N_2334,N_1760,N_1727);
and U2335 (N_2335,N_1671,N_2055);
nand U2336 (N_2336,N_1979,N_1797);
and U2337 (N_2337,N_1994,N_2237);
and U2338 (N_2338,N_1823,N_1862);
and U2339 (N_2339,N_1541,N_1660);
nand U2340 (N_2340,N_2115,N_1582);
nand U2341 (N_2341,N_1858,N_1544);
nor U2342 (N_2342,N_1532,N_2213);
nor U2343 (N_2343,N_1642,N_1791);
and U2344 (N_2344,N_2178,N_2206);
and U2345 (N_2345,N_1743,N_1526);
nor U2346 (N_2346,N_1798,N_1942);
or U2347 (N_2347,N_2221,N_1588);
nand U2348 (N_2348,N_1863,N_2174);
nor U2349 (N_2349,N_1812,N_1830);
or U2350 (N_2350,N_1866,N_2075);
nand U2351 (N_2351,N_1944,N_1530);
and U2352 (N_2352,N_1563,N_1808);
nor U2353 (N_2353,N_1895,N_1510);
nor U2354 (N_2354,N_1806,N_1740);
or U2355 (N_2355,N_1843,N_1890);
nor U2356 (N_2356,N_2138,N_2120);
and U2357 (N_2357,N_1908,N_1920);
and U2358 (N_2358,N_1616,N_1651);
xor U2359 (N_2359,N_1554,N_1966);
or U2360 (N_2360,N_1755,N_1725);
or U2361 (N_2361,N_2116,N_1820);
or U2362 (N_2362,N_2054,N_2212);
nor U2363 (N_2363,N_2042,N_1712);
nor U2364 (N_2364,N_1531,N_2249);
and U2365 (N_2365,N_1665,N_1624);
nand U2366 (N_2366,N_2154,N_2030);
or U2367 (N_2367,N_2109,N_1518);
or U2368 (N_2368,N_1774,N_2145);
nand U2369 (N_2369,N_1876,N_1517);
nor U2370 (N_2370,N_2035,N_1501);
nand U2371 (N_2371,N_1985,N_2129);
nand U2372 (N_2372,N_1664,N_1815);
nor U2373 (N_2373,N_1809,N_2150);
nor U2374 (N_2374,N_2111,N_2248);
nand U2375 (N_2375,N_1560,N_1731);
and U2376 (N_2376,N_2083,N_1756);
nor U2377 (N_2377,N_2165,N_2227);
and U2378 (N_2378,N_1515,N_2009);
and U2379 (N_2379,N_1549,N_1940);
nand U2380 (N_2380,N_1686,N_1733);
nor U2381 (N_2381,N_1829,N_1764);
and U2382 (N_2382,N_2014,N_1846);
nor U2383 (N_2383,N_1613,N_1845);
nand U2384 (N_2384,N_2186,N_1959);
and U2385 (N_2385,N_1980,N_1574);
nor U2386 (N_2386,N_2136,N_1948);
nand U2387 (N_2387,N_2033,N_1724);
nor U2388 (N_2388,N_1856,N_2226);
nand U2389 (N_2389,N_2219,N_2112);
nand U2390 (N_2390,N_1901,N_1636);
and U2391 (N_2391,N_1508,N_2239);
xor U2392 (N_2392,N_1992,N_2013);
nand U2393 (N_2393,N_1674,N_1932);
and U2394 (N_2394,N_1924,N_2079);
or U2395 (N_2395,N_1919,N_2192);
nand U2396 (N_2396,N_1640,N_1744);
or U2397 (N_2397,N_1824,N_2113);
and U2398 (N_2398,N_1976,N_1635);
nor U2399 (N_2399,N_1618,N_1896);
nand U2400 (N_2400,N_1656,N_1819);
and U2401 (N_2401,N_1590,N_2182);
nand U2402 (N_2402,N_1568,N_1507);
nand U2403 (N_2403,N_1787,N_1762);
nor U2404 (N_2404,N_2101,N_2123);
nand U2405 (N_2405,N_1600,N_1773);
nor U2406 (N_2406,N_2078,N_1759);
nor U2407 (N_2407,N_1880,N_1946);
nor U2408 (N_2408,N_2068,N_1916);
nor U2409 (N_2409,N_1962,N_1884);
nor U2410 (N_2410,N_1789,N_1556);
or U2411 (N_2411,N_1893,N_1964);
nand U2412 (N_2412,N_2008,N_2241);
and U2413 (N_2413,N_1935,N_1589);
or U2414 (N_2414,N_2216,N_2224);
and U2415 (N_2415,N_1800,N_1870);
and U2416 (N_2416,N_2180,N_1713);
or U2417 (N_2417,N_1909,N_1961);
or U2418 (N_2418,N_1897,N_1689);
and U2419 (N_2419,N_1633,N_1972);
or U2420 (N_2420,N_1851,N_2143);
and U2421 (N_2421,N_2085,N_1617);
or U2422 (N_2422,N_2183,N_1776);
or U2423 (N_2423,N_1775,N_2147);
or U2424 (N_2424,N_1503,N_1676);
or U2425 (N_2425,N_2168,N_1816);
nand U2426 (N_2426,N_1717,N_2016);
and U2427 (N_2427,N_1741,N_2060);
nor U2428 (N_2428,N_2043,N_1678);
nor U2429 (N_2429,N_2092,N_1934);
and U2430 (N_2430,N_2086,N_1957);
nand U2431 (N_2431,N_2089,N_1834);
and U2432 (N_2432,N_1645,N_1963);
nand U2433 (N_2433,N_2041,N_1578);
and U2434 (N_2434,N_2232,N_1608);
or U2435 (N_2435,N_2242,N_1587);
or U2436 (N_2436,N_1952,N_2240);
or U2437 (N_2437,N_1811,N_1814);
nand U2438 (N_2438,N_1854,N_1839);
nand U2439 (N_2439,N_1792,N_1766);
and U2440 (N_2440,N_1833,N_1732);
or U2441 (N_2441,N_2141,N_2022);
nor U2442 (N_2442,N_1742,N_2231);
nand U2443 (N_2443,N_2209,N_1512);
or U2444 (N_2444,N_2134,N_2051);
or U2445 (N_2445,N_1585,N_2082);
nand U2446 (N_2446,N_2139,N_2093);
nand U2447 (N_2447,N_1861,N_1615);
nand U2448 (N_2448,N_1997,N_2234);
and U2449 (N_2449,N_2142,N_2028);
nor U2450 (N_2450,N_2039,N_1917);
nand U2451 (N_2451,N_1627,N_1551);
or U2452 (N_2452,N_2107,N_1677);
or U2453 (N_2453,N_2245,N_1847);
or U2454 (N_2454,N_1545,N_1887);
nand U2455 (N_2455,N_2095,N_2163);
or U2456 (N_2456,N_1734,N_2084);
nor U2457 (N_2457,N_1745,N_1722);
or U2458 (N_2458,N_1736,N_1647);
nand U2459 (N_2459,N_1534,N_1960);
and U2460 (N_2460,N_1886,N_2122);
and U2461 (N_2461,N_2188,N_1706);
nand U2462 (N_2462,N_1777,N_1557);
and U2463 (N_2463,N_1524,N_1594);
nor U2464 (N_2464,N_1865,N_2201);
or U2465 (N_2465,N_1655,N_1828);
and U2466 (N_2466,N_1788,N_1630);
and U2467 (N_2467,N_2179,N_2066);
or U2468 (N_2468,N_2169,N_1715);
or U2469 (N_2469,N_1619,N_1520);
and U2470 (N_2470,N_1718,N_1561);
nor U2471 (N_2471,N_1857,N_1990);
and U2472 (N_2472,N_1539,N_1593);
or U2473 (N_2473,N_2152,N_2126);
or U2474 (N_2474,N_1591,N_1826);
nand U2475 (N_2475,N_1670,N_1953);
nand U2476 (N_2476,N_1951,N_1842);
or U2477 (N_2477,N_1757,N_2175);
and U2478 (N_2478,N_1937,N_1763);
and U2479 (N_2479,N_1970,N_1586);
nand U2480 (N_2480,N_1973,N_1986);
and U2481 (N_2481,N_2087,N_2166);
nor U2482 (N_2482,N_2131,N_1690);
or U2483 (N_2483,N_1754,N_1751);
or U2484 (N_2484,N_2065,N_1931);
or U2485 (N_2485,N_2196,N_1632);
and U2486 (N_2486,N_1930,N_2132);
and U2487 (N_2487,N_1521,N_1684);
or U2488 (N_2488,N_1849,N_2148);
nor U2489 (N_2489,N_1900,N_1595);
nor U2490 (N_2490,N_1750,N_1577);
nor U2491 (N_2491,N_1770,N_1933);
and U2492 (N_2492,N_1758,N_2181);
nor U2493 (N_2493,N_1667,N_1989);
or U2494 (N_2494,N_1771,N_2225);
and U2495 (N_2495,N_2072,N_1701);
and U2496 (N_2496,N_1835,N_1700);
and U2497 (N_2497,N_2197,N_1516);
nand U2498 (N_2498,N_2185,N_1528);
and U2499 (N_2499,N_1987,N_1555);
or U2500 (N_2500,N_1796,N_2090);
nor U2501 (N_2501,N_2002,N_1950);
nand U2502 (N_2502,N_1626,N_1738);
nand U2503 (N_2503,N_2194,N_1723);
nand U2504 (N_2504,N_1735,N_1926);
nor U2505 (N_2505,N_1614,N_2127);
and U2506 (N_2506,N_2130,N_1693);
and U2507 (N_2507,N_1984,N_1739);
and U2508 (N_2508,N_2236,N_2097);
nor U2509 (N_2509,N_1855,N_1968);
nand U2510 (N_2510,N_2202,N_2003);
and U2511 (N_2511,N_1902,N_1553);
and U2512 (N_2512,N_1878,N_2025);
nand U2513 (N_2513,N_1680,N_1625);
or U2514 (N_2514,N_1599,N_1969);
nor U2515 (N_2515,N_1906,N_1978);
and U2516 (N_2516,N_2205,N_1915);
nor U2517 (N_2517,N_2059,N_2157);
and U2518 (N_2518,N_1546,N_1889);
or U2519 (N_2519,N_1837,N_1719);
or U2520 (N_2520,N_2100,N_2223);
and U2521 (N_2521,N_1925,N_1509);
nor U2522 (N_2522,N_1579,N_2010);
nand U2523 (N_2523,N_2124,N_1584);
nand U2524 (N_2524,N_1638,N_2204);
nor U2525 (N_2525,N_1710,N_2096);
nand U2526 (N_2526,N_1646,N_1802);
or U2527 (N_2527,N_2173,N_1768);
nand U2528 (N_2528,N_2024,N_1728);
xor U2529 (N_2529,N_1698,N_1622);
or U2530 (N_2530,N_1922,N_1999);
nand U2531 (N_2531,N_2005,N_1688);
or U2532 (N_2532,N_1691,N_1730);
and U2533 (N_2533,N_1505,N_1711);
nand U2534 (N_2534,N_2167,N_2037);
and U2535 (N_2535,N_1848,N_1840);
nor U2536 (N_2536,N_1564,N_1822);
nand U2537 (N_2537,N_2187,N_1945);
and U2538 (N_2538,N_1669,N_1552);
nor U2539 (N_2539,N_1695,N_2164);
nor U2540 (N_2540,N_1779,N_1592);
and U2541 (N_2541,N_1853,N_1795);
nor U2542 (N_2542,N_1604,N_1832);
and U2543 (N_2543,N_1817,N_1649);
nor U2544 (N_2544,N_1769,N_1995);
and U2545 (N_2545,N_1927,N_2064);
or U2546 (N_2546,N_1575,N_2045);
and U2547 (N_2547,N_1535,N_1572);
nand U2548 (N_2548,N_2021,N_2247);
and U2549 (N_2549,N_2050,N_1752);
or U2550 (N_2550,N_1781,N_1894);
or U2551 (N_2551,N_1836,N_2088);
or U2552 (N_2552,N_1958,N_2031);
nor U2553 (N_2553,N_1610,N_1643);
or U2554 (N_2554,N_2128,N_1827);
and U2555 (N_2555,N_1914,N_1513);
or U2556 (N_2556,N_2006,N_1983);
and U2557 (N_2557,N_1965,N_1537);
nand U2558 (N_2558,N_1747,N_2007);
and U2559 (N_2559,N_2146,N_1872);
nor U2560 (N_2560,N_1941,N_2191);
nor U2561 (N_2561,N_2038,N_1996);
or U2562 (N_2562,N_2063,N_1648);
nand U2563 (N_2563,N_1818,N_1697);
nand U2564 (N_2564,N_2026,N_1883);
and U2565 (N_2565,N_1907,N_2159);
nor U2566 (N_2566,N_2210,N_1571);
nand U2567 (N_2567,N_2238,N_1881);
and U2568 (N_2568,N_1685,N_1720);
and U2569 (N_2569,N_1704,N_1971);
or U2570 (N_2570,N_1888,N_1825);
nand U2571 (N_2571,N_2190,N_2200);
nor U2572 (N_2572,N_1891,N_1783);
nand U2573 (N_2573,N_1672,N_1821);
nor U2574 (N_2574,N_2080,N_1885);
nand U2575 (N_2575,N_2171,N_1602);
and U2576 (N_2576,N_1974,N_1929);
nor U2577 (N_2577,N_1576,N_2053);
or U2578 (N_2578,N_1721,N_1522);
nand U2579 (N_2579,N_1570,N_2046);
nand U2580 (N_2580,N_1807,N_1794);
or U2581 (N_2581,N_1527,N_2032);
and U2582 (N_2582,N_2012,N_2044);
nor U2583 (N_2583,N_2121,N_1661);
nor U2584 (N_2584,N_1772,N_2176);
or U2585 (N_2585,N_1921,N_1598);
or U2586 (N_2586,N_1683,N_1652);
nor U2587 (N_2587,N_1601,N_2217);
nor U2588 (N_2588,N_1620,N_1841);
or U2589 (N_2589,N_2230,N_2160);
nand U2590 (N_2590,N_1988,N_1699);
nand U2591 (N_2591,N_1805,N_1879);
or U2592 (N_2592,N_1631,N_1682);
or U2593 (N_2593,N_1904,N_1852);
nor U2594 (N_2594,N_2067,N_2162);
nor U2595 (N_2595,N_2235,N_1603);
nand U2596 (N_2596,N_1746,N_1868);
nor U2597 (N_2597,N_1559,N_2193);
nor U2598 (N_2598,N_1607,N_1998);
nor U2599 (N_2599,N_1804,N_1943);
nor U2600 (N_2600,N_1692,N_2091);
and U2601 (N_2601,N_1707,N_2069);
or U2602 (N_2602,N_1637,N_1947);
nor U2603 (N_2603,N_2034,N_1780);
and U2604 (N_2604,N_1654,N_2243);
nor U2605 (N_2605,N_1504,N_2105);
or U2606 (N_2606,N_1621,N_1569);
nor U2607 (N_2607,N_2074,N_1708);
and U2608 (N_2608,N_1565,N_1873);
and U2609 (N_2609,N_1506,N_2104);
nor U2610 (N_2610,N_1543,N_1864);
nor U2611 (N_2611,N_2195,N_1609);
nand U2612 (N_2612,N_2071,N_1761);
and U2613 (N_2613,N_1567,N_2015);
nor U2614 (N_2614,N_1737,N_1784);
or U2615 (N_2615,N_1714,N_1982);
and U2616 (N_2616,N_2228,N_2001);
nor U2617 (N_2617,N_1511,N_1838);
and U2618 (N_2618,N_2099,N_1668);
or U2619 (N_2619,N_1813,N_2040);
nor U2620 (N_2620,N_1653,N_2057);
and U2621 (N_2621,N_2144,N_1687);
nand U2622 (N_2622,N_1918,N_1583);
nand U2623 (N_2623,N_2161,N_2027);
and U2624 (N_2624,N_1639,N_2000);
nor U2625 (N_2625,N_1741,N_1545);
nor U2626 (N_2626,N_2245,N_1783);
xor U2627 (N_2627,N_1938,N_1523);
and U2628 (N_2628,N_1775,N_1513);
or U2629 (N_2629,N_1902,N_1612);
nand U2630 (N_2630,N_2059,N_1555);
or U2631 (N_2631,N_1721,N_1914);
or U2632 (N_2632,N_1663,N_1867);
or U2633 (N_2633,N_2098,N_2065);
or U2634 (N_2634,N_1718,N_1984);
and U2635 (N_2635,N_2242,N_1831);
nand U2636 (N_2636,N_2078,N_1752);
or U2637 (N_2637,N_2230,N_2087);
and U2638 (N_2638,N_1889,N_2019);
and U2639 (N_2639,N_2053,N_1868);
nor U2640 (N_2640,N_1547,N_2006);
nor U2641 (N_2641,N_2238,N_2005);
and U2642 (N_2642,N_1848,N_1622);
or U2643 (N_2643,N_2071,N_1663);
nor U2644 (N_2644,N_1630,N_1989);
nand U2645 (N_2645,N_2225,N_1954);
nor U2646 (N_2646,N_1846,N_1692);
or U2647 (N_2647,N_1839,N_1594);
and U2648 (N_2648,N_2188,N_2051);
or U2649 (N_2649,N_1619,N_2249);
or U2650 (N_2650,N_1817,N_2086);
or U2651 (N_2651,N_2041,N_1886);
nor U2652 (N_2652,N_2133,N_1830);
nand U2653 (N_2653,N_1990,N_1731);
nor U2654 (N_2654,N_2165,N_1893);
or U2655 (N_2655,N_1740,N_1590);
and U2656 (N_2656,N_1919,N_1727);
nor U2657 (N_2657,N_2170,N_1520);
or U2658 (N_2658,N_1757,N_2238);
nor U2659 (N_2659,N_2134,N_1755);
nor U2660 (N_2660,N_2062,N_2191);
nand U2661 (N_2661,N_2054,N_2214);
or U2662 (N_2662,N_1639,N_1885);
and U2663 (N_2663,N_1946,N_1553);
nor U2664 (N_2664,N_2179,N_1823);
nor U2665 (N_2665,N_1737,N_2069);
nor U2666 (N_2666,N_1759,N_1800);
nand U2667 (N_2667,N_1943,N_1874);
nor U2668 (N_2668,N_1569,N_2110);
or U2669 (N_2669,N_2115,N_2177);
nor U2670 (N_2670,N_1594,N_2174);
nor U2671 (N_2671,N_1665,N_1591);
nor U2672 (N_2672,N_1728,N_1564);
nand U2673 (N_2673,N_2023,N_1671);
nand U2674 (N_2674,N_1758,N_2201);
and U2675 (N_2675,N_2115,N_1984);
nor U2676 (N_2676,N_1885,N_2152);
nand U2677 (N_2677,N_1872,N_1652);
and U2678 (N_2678,N_1511,N_1737);
nor U2679 (N_2679,N_2078,N_1787);
nor U2680 (N_2680,N_1684,N_1879);
nand U2681 (N_2681,N_2033,N_1515);
or U2682 (N_2682,N_1810,N_1624);
and U2683 (N_2683,N_1932,N_1606);
or U2684 (N_2684,N_1725,N_1906);
nand U2685 (N_2685,N_1833,N_1835);
nor U2686 (N_2686,N_1652,N_2022);
and U2687 (N_2687,N_1849,N_1608);
nor U2688 (N_2688,N_1701,N_1786);
or U2689 (N_2689,N_1917,N_1904);
and U2690 (N_2690,N_1747,N_1507);
and U2691 (N_2691,N_1796,N_2215);
nor U2692 (N_2692,N_2232,N_1506);
or U2693 (N_2693,N_1616,N_1953);
or U2694 (N_2694,N_2008,N_1794);
xnor U2695 (N_2695,N_1856,N_1724);
nor U2696 (N_2696,N_2052,N_2103);
and U2697 (N_2697,N_2219,N_1683);
nand U2698 (N_2698,N_1509,N_1968);
nor U2699 (N_2699,N_2196,N_1707);
or U2700 (N_2700,N_1618,N_1981);
nand U2701 (N_2701,N_1700,N_1608);
or U2702 (N_2702,N_1899,N_1715);
or U2703 (N_2703,N_1601,N_2041);
nor U2704 (N_2704,N_2083,N_1997);
or U2705 (N_2705,N_2068,N_2069);
nand U2706 (N_2706,N_1765,N_1745);
and U2707 (N_2707,N_1732,N_1671);
or U2708 (N_2708,N_2171,N_1733);
xnor U2709 (N_2709,N_1910,N_2234);
nand U2710 (N_2710,N_2204,N_1817);
and U2711 (N_2711,N_2176,N_1564);
nand U2712 (N_2712,N_2023,N_1845);
nand U2713 (N_2713,N_2238,N_2022);
nand U2714 (N_2714,N_2118,N_2205);
nand U2715 (N_2715,N_1974,N_2049);
or U2716 (N_2716,N_2151,N_1729);
nand U2717 (N_2717,N_1620,N_1639);
or U2718 (N_2718,N_2221,N_2063);
nand U2719 (N_2719,N_1872,N_1667);
nand U2720 (N_2720,N_1808,N_2191);
nor U2721 (N_2721,N_1986,N_2073);
nor U2722 (N_2722,N_1519,N_1631);
and U2723 (N_2723,N_2189,N_2026);
nand U2724 (N_2724,N_1505,N_2041);
nor U2725 (N_2725,N_2205,N_2048);
xnor U2726 (N_2726,N_1898,N_2005);
nand U2727 (N_2727,N_2119,N_2008);
nor U2728 (N_2728,N_1944,N_2210);
or U2729 (N_2729,N_1547,N_2193);
and U2730 (N_2730,N_1927,N_2182);
and U2731 (N_2731,N_1541,N_1622);
nor U2732 (N_2732,N_1861,N_1945);
nor U2733 (N_2733,N_1878,N_1601);
and U2734 (N_2734,N_1699,N_2218);
or U2735 (N_2735,N_2148,N_2205);
and U2736 (N_2736,N_1848,N_1880);
nand U2737 (N_2737,N_1825,N_2166);
and U2738 (N_2738,N_1665,N_1630);
or U2739 (N_2739,N_2005,N_1565);
and U2740 (N_2740,N_1781,N_1821);
nand U2741 (N_2741,N_2187,N_1926);
or U2742 (N_2742,N_1633,N_1834);
and U2743 (N_2743,N_1834,N_1505);
and U2744 (N_2744,N_1819,N_1767);
nand U2745 (N_2745,N_1524,N_2005);
or U2746 (N_2746,N_1718,N_1589);
and U2747 (N_2747,N_1967,N_1720);
xnor U2748 (N_2748,N_2209,N_1968);
nand U2749 (N_2749,N_1862,N_1839);
and U2750 (N_2750,N_1570,N_1978);
or U2751 (N_2751,N_2221,N_1728);
nor U2752 (N_2752,N_2081,N_1900);
nand U2753 (N_2753,N_2065,N_2082);
or U2754 (N_2754,N_2076,N_1735);
and U2755 (N_2755,N_1890,N_2185);
nor U2756 (N_2756,N_1556,N_1552);
nand U2757 (N_2757,N_1629,N_2115);
xnor U2758 (N_2758,N_1593,N_2225);
nor U2759 (N_2759,N_1982,N_1534);
nand U2760 (N_2760,N_2071,N_2204);
and U2761 (N_2761,N_1921,N_1544);
nor U2762 (N_2762,N_1680,N_1556);
nor U2763 (N_2763,N_1936,N_2075);
nor U2764 (N_2764,N_1830,N_1829);
or U2765 (N_2765,N_1801,N_1985);
and U2766 (N_2766,N_2203,N_2042);
or U2767 (N_2767,N_1997,N_1567);
nand U2768 (N_2768,N_1701,N_1822);
nor U2769 (N_2769,N_1672,N_2219);
and U2770 (N_2770,N_1814,N_1604);
nor U2771 (N_2771,N_1758,N_1820);
and U2772 (N_2772,N_2098,N_1855);
or U2773 (N_2773,N_1934,N_1785);
nor U2774 (N_2774,N_1768,N_1593);
nand U2775 (N_2775,N_1820,N_1992);
nand U2776 (N_2776,N_2219,N_2020);
nor U2777 (N_2777,N_2081,N_2143);
or U2778 (N_2778,N_1757,N_1611);
nor U2779 (N_2779,N_2036,N_1555);
nor U2780 (N_2780,N_1821,N_2064);
and U2781 (N_2781,N_1609,N_2085);
and U2782 (N_2782,N_1840,N_1852);
nor U2783 (N_2783,N_2133,N_2036);
nor U2784 (N_2784,N_2140,N_1526);
and U2785 (N_2785,N_1814,N_2007);
or U2786 (N_2786,N_2018,N_1591);
or U2787 (N_2787,N_2014,N_1999);
and U2788 (N_2788,N_1856,N_1819);
nor U2789 (N_2789,N_1971,N_1553);
or U2790 (N_2790,N_1859,N_1752);
nor U2791 (N_2791,N_2100,N_1783);
or U2792 (N_2792,N_2080,N_1662);
nor U2793 (N_2793,N_1881,N_2145);
nor U2794 (N_2794,N_1916,N_1934);
nor U2795 (N_2795,N_1566,N_2112);
or U2796 (N_2796,N_2040,N_1592);
nand U2797 (N_2797,N_1824,N_1765);
nor U2798 (N_2798,N_2038,N_1582);
nand U2799 (N_2799,N_1824,N_1790);
nor U2800 (N_2800,N_1630,N_1578);
and U2801 (N_2801,N_1783,N_1975);
or U2802 (N_2802,N_1989,N_1775);
nand U2803 (N_2803,N_1729,N_1855);
or U2804 (N_2804,N_2028,N_2016);
nor U2805 (N_2805,N_1804,N_1651);
nand U2806 (N_2806,N_1647,N_2042);
or U2807 (N_2807,N_2190,N_2204);
xnor U2808 (N_2808,N_2184,N_1528);
or U2809 (N_2809,N_2091,N_1607);
nand U2810 (N_2810,N_2237,N_1684);
and U2811 (N_2811,N_1588,N_1609);
nor U2812 (N_2812,N_1517,N_2080);
nor U2813 (N_2813,N_1506,N_1562);
nand U2814 (N_2814,N_2145,N_2018);
nand U2815 (N_2815,N_2144,N_1734);
or U2816 (N_2816,N_2242,N_1970);
or U2817 (N_2817,N_2247,N_2100);
or U2818 (N_2818,N_1613,N_1863);
or U2819 (N_2819,N_1971,N_1630);
nor U2820 (N_2820,N_2104,N_2143);
nor U2821 (N_2821,N_1706,N_1710);
and U2822 (N_2822,N_1659,N_1661);
or U2823 (N_2823,N_2192,N_2183);
and U2824 (N_2824,N_1968,N_1687);
nor U2825 (N_2825,N_1517,N_1553);
nand U2826 (N_2826,N_1653,N_2096);
or U2827 (N_2827,N_2223,N_1525);
or U2828 (N_2828,N_2158,N_1890);
nand U2829 (N_2829,N_1927,N_2206);
and U2830 (N_2830,N_1769,N_2185);
or U2831 (N_2831,N_1941,N_1703);
nand U2832 (N_2832,N_2103,N_1887);
nor U2833 (N_2833,N_1872,N_1818);
nand U2834 (N_2834,N_2232,N_2062);
nor U2835 (N_2835,N_1851,N_2037);
and U2836 (N_2836,N_1575,N_1721);
nor U2837 (N_2837,N_2229,N_2022);
nand U2838 (N_2838,N_2148,N_2030);
or U2839 (N_2839,N_1800,N_1812);
or U2840 (N_2840,N_1728,N_1729);
and U2841 (N_2841,N_2143,N_2066);
nand U2842 (N_2842,N_1601,N_1734);
or U2843 (N_2843,N_1686,N_1580);
nor U2844 (N_2844,N_2230,N_2034);
nor U2845 (N_2845,N_2078,N_1744);
nor U2846 (N_2846,N_1805,N_1668);
nand U2847 (N_2847,N_1526,N_2247);
nor U2848 (N_2848,N_2186,N_1582);
nand U2849 (N_2849,N_2159,N_2077);
nand U2850 (N_2850,N_2081,N_2127);
or U2851 (N_2851,N_1645,N_2238);
nand U2852 (N_2852,N_1957,N_1927);
and U2853 (N_2853,N_1668,N_1664);
or U2854 (N_2854,N_2213,N_2072);
xnor U2855 (N_2855,N_2171,N_1696);
or U2856 (N_2856,N_2039,N_1594);
nand U2857 (N_2857,N_1658,N_2127);
and U2858 (N_2858,N_1943,N_2005);
or U2859 (N_2859,N_2104,N_2198);
and U2860 (N_2860,N_2113,N_1886);
nor U2861 (N_2861,N_1611,N_1667);
or U2862 (N_2862,N_1962,N_1754);
and U2863 (N_2863,N_1529,N_1602);
and U2864 (N_2864,N_1788,N_2213);
nand U2865 (N_2865,N_2019,N_2113);
nand U2866 (N_2866,N_1695,N_2188);
nand U2867 (N_2867,N_1564,N_2030);
nand U2868 (N_2868,N_1958,N_2096);
or U2869 (N_2869,N_1786,N_1929);
or U2870 (N_2870,N_1984,N_2011);
and U2871 (N_2871,N_1553,N_2067);
or U2872 (N_2872,N_1993,N_1601);
or U2873 (N_2873,N_1525,N_2233);
nor U2874 (N_2874,N_1617,N_2244);
or U2875 (N_2875,N_1997,N_1597);
nand U2876 (N_2876,N_1663,N_1894);
and U2877 (N_2877,N_1842,N_1699);
nand U2878 (N_2878,N_1880,N_1794);
and U2879 (N_2879,N_1960,N_1540);
nand U2880 (N_2880,N_1800,N_2102);
nor U2881 (N_2881,N_2205,N_1531);
and U2882 (N_2882,N_2159,N_2072);
xnor U2883 (N_2883,N_1841,N_1615);
or U2884 (N_2884,N_1562,N_1667);
nand U2885 (N_2885,N_1652,N_1866);
or U2886 (N_2886,N_1885,N_1553);
nor U2887 (N_2887,N_1706,N_1830);
nor U2888 (N_2888,N_1765,N_1761);
nor U2889 (N_2889,N_1766,N_2180);
nand U2890 (N_2890,N_1550,N_2138);
nor U2891 (N_2891,N_1548,N_1643);
nand U2892 (N_2892,N_1556,N_1832);
and U2893 (N_2893,N_2028,N_2214);
or U2894 (N_2894,N_2087,N_1667);
nand U2895 (N_2895,N_1544,N_2192);
nor U2896 (N_2896,N_1829,N_1856);
and U2897 (N_2897,N_1732,N_1831);
nor U2898 (N_2898,N_1665,N_1997);
nor U2899 (N_2899,N_1621,N_2183);
nand U2900 (N_2900,N_1880,N_1958);
nand U2901 (N_2901,N_2231,N_1688);
and U2902 (N_2902,N_1835,N_2212);
and U2903 (N_2903,N_1704,N_1650);
nor U2904 (N_2904,N_2078,N_1738);
nor U2905 (N_2905,N_2054,N_1674);
nand U2906 (N_2906,N_1614,N_1976);
nor U2907 (N_2907,N_2013,N_1845);
and U2908 (N_2908,N_1562,N_1995);
nand U2909 (N_2909,N_1626,N_2212);
and U2910 (N_2910,N_1509,N_1823);
or U2911 (N_2911,N_2017,N_1531);
nor U2912 (N_2912,N_2098,N_1526);
nand U2913 (N_2913,N_1830,N_1576);
and U2914 (N_2914,N_2116,N_2229);
or U2915 (N_2915,N_1535,N_2069);
nand U2916 (N_2916,N_2154,N_1970);
and U2917 (N_2917,N_1923,N_1549);
nand U2918 (N_2918,N_1899,N_1978);
nor U2919 (N_2919,N_1515,N_2025);
nor U2920 (N_2920,N_1959,N_1567);
nand U2921 (N_2921,N_1769,N_1964);
and U2922 (N_2922,N_2226,N_1772);
nand U2923 (N_2923,N_1935,N_1654);
xnor U2924 (N_2924,N_1565,N_1599);
and U2925 (N_2925,N_1802,N_1997);
and U2926 (N_2926,N_1752,N_1932);
nor U2927 (N_2927,N_1505,N_2161);
or U2928 (N_2928,N_1559,N_1764);
or U2929 (N_2929,N_1651,N_1855);
and U2930 (N_2930,N_2249,N_1969);
nor U2931 (N_2931,N_1620,N_1669);
nor U2932 (N_2932,N_2130,N_1709);
or U2933 (N_2933,N_2239,N_1845);
xnor U2934 (N_2934,N_1548,N_1554);
or U2935 (N_2935,N_2095,N_1885);
nand U2936 (N_2936,N_2035,N_1750);
and U2937 (N_2937,N_1537,N_2196);
xnor U2938 (N_2938,N_1754,N_1988);
and U2939 (N_2939,N_2191,N_1856);
nor U2940 (N_2940,N_1706,N_1978);
and U2941 (N_2941,N_2160,N_1656);
nand U2942 (N_2942,N_1986,N_1897);
nand U2943 (N_2943,N_1807,N_1626);
and U2944 (N_2944,N_1808,N_1972);
nor U2945 (N_2945,N_1747,N_1720);
nor U2946 (N_2946,N_1927,N_1936);
nand U2947 (N_2947,N_1948,N_1608);
or U2948 (N_2948,N_2209,N_1680);
nor U2949 (N_2949,N_1891,N_1882);
or U2950 (N_2950,N_1792,N_2078);
nand U2951 (N_2951,N_1856,N_1853);
nand U2952 (N_2952,N_1944,N_1611);
nand U2953 (N_2953,N_1585,N_2208);
nor U2954 (N_2954,N_2087,N_1617);
or U2955 (N_2955,N_1579,N_2052);
or U2956 (N_2956,N_1659,N_1653);
or U2957 (N_2957,N_1848,N_1511);
and U2958 (N_2958,N_2032,N_1703);
nand U2959 (N_2959,N_2035,N_1529);
nand U2960 (N_2960,N_1522,N_1871);
and U2961 (N_2961,N_1727,N_2091);
and U2962 (N_2962,N_1644,N_1976);
and U2963 (N_2963,N_2065,N_2157);
nor U2964 (N_2964,N_2227,N_1689);
and U2965 (N_2965,N_1779,N_1589);
nand U2966 (N_2966,N_1922,N_2046);
nand U2967 (N_2967,N_1576,N_2229);
nand U2968 (N_2968,N_2134,N_2101);
and U2969 (N_2969,N_2134,N_1883);
or U2970 (N_2970,N_1677,N_1842);
nand U2971 (N_2971,N_1531,N_1604);
and U2972 (N_2972,N_1839,N_1544);
nor U2973 (N_2973,N_1736,N_2171);
or U2974 (N_2974,N_1537,N_1735);
or U2975 (N_2975,N_2165,N_2072);
nor U2976 (N_2976,N_1943,N_1830);
and U2977 (N_2977,N_2021,N_2127);
nand U2978 (N_2978,N_1544,N_1944);
nand U2979 (N_2979,N_1917,N_1909);
nand U2980 (N_2980,N_1721,N_2216);
xor U2981 (N_2981,N_1919,N_2196);
or U2982 (N_2982,N_2211,N_1860);
and U2983 (N_2983,N_1550,N_2057);
or U2984 (N_2984,N_1919,N_2044);
or U2985 (N_2985,N_1916,N_1660);
nor U2986 (N_2986,N_1781,N_2068);
nor U2987 (N_2987,N_2089,N_2049);
nand U2988 (N_2988,N_1738,N_1907);
nand U2989 (N_2989,N_2168,N_1720);
nor U2990 (N_2990,N_1748,N_1863);
and U2991 (N_2991,N_1829,N_1793);
nor U2992 (N_2992,N_2096,N_1808);
or U2993 (N_2993,N_1948,N_1849);
or U2994 (N_2994,N_1518,N_1559);
and U2995 (N_2995,N_1795,N_1759);
and U2996 (N_2996,N_2021,N_2047);
or U2997 (N_2997,N_1999,N_1691);
or U2998 (N_2998,N_1890,N_1993);
and U2999 (N_2999,N_1789,N_1678);
or UO_0 (O_0,N_2700,N_2479);
or UO_1 (O_1,N_2749,N_2649);
nand UO_2 (O_2,N_2958,N_2707);
nand UO_3 (O_3,N_2269,N_2303);
or UO_4 (O_4,N_2973,N_2406);
and UO_5 (O_5,N_2447,N_2753);
nand UO_6 (O_6,N_2694,N_2645);
and UO_7 (O_7,N_2853,N_2439);
nand UO_8 (O_8,N_2897,N_2785);
nor UO_9 (O_9,N_2601,N_2567);
and UO_10 (O_10,N_2484,N_2318);
or UO_11 (O_11,N_2326,N_2533);
or UO_12 (O_12,N_2278,N_2481);
and UO_13 (O_13,N_2951,N_2452);
nand UO_14 (O_14,N_2741,N_2959);
nand UO_15 (O_15,N_2540,N_2669);
and UO_16 (O_16,N_2451,N_2290);
and UO_17 (O_17,N_2857,N_2494);
and UO_18 (O_18,N_2713,N_2619);
or UO_19 (O_19,N_2801,N_2756);
nand UO_20 (O_20,N_2935,N_2653);
or UO_21 (O_21,N_2416,N_2841);
nand UO_22 (O_22,N_2666,N_2508);
or UO_23 (O_23,N_2586,N_2317);
and UO_24 (O_24,N_2525,N_2693);
or UO_25 (O_25,N_2992,N_2727);
or UO_26 (O_26,N_2743,N_2957);
nand UO_27 (O_27,N_2850,N_2314);
nor UO_28 (O_28,N_2954,N_2724);
nand UO_29 (O_29,N_2379,N_2275);
and UO_30 (O_30,N_2974,N_2482);
nand UO_31 (O_31,N_2944,N_2916);
nor UO_32 (O_32,N_2469,N_2385);
or UO_33 (O_33,N_2260,N_2579);
nand UO_34 (O_34,N_2972,N_2800);
and UO_35 (O_35,N_2560,N_2852);
or UO_36 (O_36,N_2747,N_2321);
nor UO_37 (O_37,N_2739,N_2389);
and UO_38 (O_38,N_2914,N_2903);
nor UO_39 (O_39,N_2824,N_2812);
and UO_40 (O_40,N_2612,N_2918);
and UO_41 (O_41,N_2263,N_2796);
nor UO_42 (O_42,N_2574,N_2359);
nand UO_43 (O_43,N_2765,N_2689);
or UO_44 (O_44,N_2524,N_2632);
nor UO_45 (O_45,N_2660,N_2426);
and UO_46 (O_46,N_2499,N_2648);
or UO_47 (O_47,N_2840,N_2438);
or UO_48 (O_48,N_2488,N_2310);
nand UO_49 (O_49,N_2827,N_2474);
or UO_50 (O_50,N_2589,N_2883);
and UO_51 (O_51,N_2692,N_2895);
or UO_52 (O_52,N_2329,N_2699);
or UO_53 (O_53,N_2826,N_2558);
nor UO_54 (O_54,N_2950,N_2599);
nor UO_55 (O_55,N_2718,N_2774);
nand UO_56 (O_56,N_2886,N_2289);
nor UO_57 (O_57,N_2614,N_2473);
and UO_58 (O_58,N_2776,N_2596);
nor UO_59 (O_59,N_2503,N_2717);
or UO_60 (O_60,N_2360,N_2584);
or UO_61 (O_61,N_2752,N_2984);
or UO_62 (O_62,N_2334,N_2864);
nor UO_63 (O_63,N_2870,N_2745);
nand UO_64 (O_64,N_2372,N_2608);
nor UO_65 (O_65,N_2414,N_2851);
and UO_66 (O_66,N_2298,N_2548);
and UO_67 (O_67,N_2302,N_2641);
or UO_68 (O_68,N_2513,N_2910);
nand UO_69 (O_69,N_2415,N_2575);
or UO_70 (O_70,N_2705,N_2828);
or UO_71 (O_71,N_2330,N_2375);
and UO_72 (O_72,N_2576,N_2328);
and UO_73 (O_73,N_2993,N_2642);
and UO_74 (O_74,N_2907,N_2799);
nand UO_75 (O_75,N_2673,N_2428);
or UO_76 (O_76,N_2809,N_2740);
nor UO_77 (O_77,N_2647,N_2267);
and UO_78 (O_78,N_2622,N_2408);
nand UO_79 (O_79,N_2404,N_2867);
or UO_80 (O_80,N_2505,N_2448);
or UO_81 (O_81,N_2498,N_2256);
or UO_82 (O_82,N_2273,N_2860);
or UO_83 (O_83,N_2885,N_2412);
or UO_84 (O_84,N_2443,N_2582);
nand UO_85 (O_85,N_2313,N_2701);
nor UO_86 (O_86,N_2901,N_2822);
nor UO_87 (O_87,N_2555,N_2947);
or UO_88 (O_88,N_2478,N_2985);
and UO_89 (O_89,N_2435,N_2549);
and UO_90 (O_90,N_2353,N_2581);
nand UO_91 (O_91,N_2607,N_2899);
nor UO_92 (O_92,N_2345,N_2716);
nand UO_93 (O_93,N_2490,N_2735);
or UO_94 (O_94,N_2783,N_2585);
nor UO_95 (O_95,N_2833,N_2733);
nand UO_96 (O_96,N_2532,N_2876);
xnor UO_97 (O_97,N_2880,N_2388);
nor UO_98 (O_98,N_2356,N_2909);
and UO_99 (O_99,N_2652,N_2489);
nand UO_100 (O_100,N_2967,N_2583);
xor UO_101 (O_101,N_2775,N_2434);
or UO_102 (O_102,N_2915,N_2491);
and UO_103 (O_103,N_2790,N_2299);
nor UO_104 (O_104,N_2687,N_2920);
nor UO_105 (O_105,N_2670,N_2422);
and UO_106 (O_106,N_2455,N_2877);
nor UO_107 (O_107,N_2963,N_2633);
or UO_108 (O_108,N_2336,N_2846);
nor UO_109 (O_109,N_2611,N_2424);
nand UO_110 (O_110,N_2654,N_2308);
and UO_111 (O_111,N_2600,N_2587);
and UO_112 (O_112,N_2358,N_2629);
and UO_113 (O_113,N_2795,N_2520);
or UO_114 (O_114,N_2997,N_2657);
nand UO_115 (O_115,N_2460,N_2571);
nor UO_116 (O_116,N_2517,N_2709);
and UO_117 (O_117,N_2684,N_2397);
nand UO_118 (O_118,N_2613,N_2798);
or UO_119 (O_119,N_2364,N_2971);
nor UO_120 (O_120,N_2616,N_2808);
and UO_121 (O_121,N_2347,N_2676);
nand UO_122 (O_122,N_2392,N_2495);
xor UO_123 (O_123,N_2387,N_2946);
or UO_124 (O_124,N_2931,N_2965);
or UO_125 (O_125,N_2938,N_2624);
and UO_126 (O_126,N_2319,N_2887);
nand UO_127 (O_127,N_2834,N_2282);
or UO_128 (O_128,N_2483,N_2922);
and UO_129 (O_129,N_2295,N_2723);
and UO_130 (O_130,N_2939,N_2773);
nand UO_131 (O_131,N_2602,N_2593);
nand UO_132 (O_132,N_2941,N_2953);
and UO_133 (O_133,N_2988,N_2272);
or UO_134 (O_134,N_2541,N_2871);
and UO_135 (O_135,N_2284,N_2725);
nor UO_136 (O_136,N_2445,N_2450);
or UO_137 (O_137,N_2458,N_2528);
or UO_138 (O_138,N_2442,N_2697);
or UO_139 (O_139,N_2721,N_2526);
and UO_140 (O_140,N_2849,N_2879);
nand UO_141 (O_141,N_2861,N_2547);
and UO_142 (O_142,N_2444,N_2337);
nand UO_143 (O_143,N_2307,N_2814);
nor UO_144 (O_144,N_2875,N_2744);
nand UO_145 (O_145,N_2534,N_2341);
nand UO_146 (O_146,N_2522,N_2480);
nor UO_147 (O_147,N_2573,N_2924);
nor UO_148 (O_148,N_2906,N_2832);
or UO_149 (O_149,N_2651,N_2810);
or UO_150 (O_150,N_2952,N_2748);
and UO_151 (O_151,N_2989,N_2288);
nor UO_152 (O_152,N_2370,N_2769);
nand UO_153 (O_153,N_2511,N_2787);
nand UO_154 (O_154,N_2889,N_2943);
nand UO_155 (O_155,N_2802,N_2276);
nor UO_156 (O_156,N_2896,N_2264);
xor UO_157 (O_157,N_2759,N_2902);
nor UO_158 (O_158,N_2923,N_2312);
and UO_159 (O_159,N_2606,N_2913);
nand UO_160 (O_160,N_2979,N_2767);
and UO_161 (O_161,N_2929,N_2698);
nor UO_162 (O_162,N_2766,N_2493);
nand UO_163 (O_163,N_2515,N_2683);
and UO_164 (O_164,N_2892,N_2323);
nand UO_165 (O_165,N_2615,N_2964);
nor UO_166 (O_166,N_2893,N_2461);
nor UO_167 (O_167,N_2771,N_2381);
or UO_168 (O_168,N_2786,N_2430);
or UO_169 (O_169,N_2501,N_2253);
and UO_170 (O_170,N_2262,N_2566);
nand UO_171 (O_171,N_2572,N_2655);
or UO_172 (O_172,N_2791,N_2859);
or UO_173 (O_173,N_2757,N_2368);
or UO_174 (O_174,N_2704,N_2933);
and UO_175 (O_175,N_2722,N_2559);
and UO_176 (O_176,N_2268,N_2564);
nor UO_177 (O_177,N_2873,N_2836);
nor UO_178 (O_178,N_2325,N_2848);
nor UO_179 (O_179,N_2680,N_2663);
nor UO_180 (O_180,N_2618,N_2750);
and UO_181 (O_181,N_2970,N_2590);
xor UO_182 (O_182,N_2627,N_2409);
nand UO_183 (O_183,N_2485,N_2994);
nor UO_184 (O_184,N_2369,N_2664);
nor UO_185 (O_185,N_2755,N_2921);
and UO_186 (O_186,N_2736,N_2293);
nand UO_187 (O_187,N_2592,N_2306);
and UO_188 (O_188,N_2554,N_2839);
or UO_189 (O_189,N_2603,N_2468);
nand UO_190 (O_190,N_2527,N_2354);
nor UO_191 (O_191,N_2980,N_2975);
nand UO_192 (O_192,N_2565,N_2637);
nand UO_193 (O_193,N_2830,N_2838);
or UO_194 (O_194,N_2620,N_2391);
nand UO_195 (O_195,N_2597,N_2644);
or UO_196 (O_196,N_2456,N_2780);
nor UO_197 (O_197,N_2936,N_2677);
nand UO_198 (O_198,N_2390,N_2667);
and UO_199 (O_199,N_2784,N_2546);
nor UO_200 (O_200,N_2542,N_2333);
or UO_201 (O_201,N_2636,N_2423);
nand UO_202 (O_202,N_2398,N_2316);
nand UO_203 (O_203,N_2371,N_2731);
nand UO_204 (O_204,N_2315,N_2617);
or UO_205 (O_205,N_2431,N_2908);
nor UO_206 (O_206,N_2441,N_2804);
nand UO_207 (O_207,N_2343,N_2728);
and UO_208 (O_208,N_2761,N_2516);
or UO_209 (O_209,N_2311,N_2781);
nand UO_210 (O_210,N_2588,N_2477);
nor UO_211 (O_211,N_2506,N_2578);
and UO_212 (O_212,N_2662,N_2470);
and UO_213 (O_213,N_2598,N_2778);
nor UO_214 (O_214,N_2320,N_2768);
and UO_215 (O_215,N_2543,N_2961);
nor UO_216 (O_216,N_2720,N_2928);
and UO_217 (O_217,N_2674,N_2521);
nor UO_218 (O_218,N_2868,N_2695);
nand UO_219 (O_219,N_2854,N_2348);
and UO_220 (O_220,N_2638,N_2996);
or UO_221 (O_221,N_2726,N_2969);
nand UO_222 (O_222,N_2365,N_2917);
nand UO_223 (O_223,N_2466,N_2668);
nor UO_224 (O_224,N_2259,N_2550);
or UO_225 (O_225,N_2252,N_2563);
and UO_226 (O_226,N_2402,N_2255);
nand UO_227 (O_227,N_2497,N_2811);
or UO_228 (O_228,N_2682,N_2454);
nor UO_229 (O_229,N_2835,N_2817);
and UO_230 (O_230,N_2562,N_2639);
nand UO_231 (O_231,N_2383,N_2283);
nand UO_232 (O_232,N_2300,N_2856);
nand UO_233 (O_233,N_2948,N_2539);
or UO_234 (O_234,N_2715,N_2509);
nand UO_235 (O_235,N_2912,N_2421);
or UO_236 (O_236,N_2955,N_2779);
xor UO_237 (O_237,N_2987,N_2453);
nand UO_238 (O_238,N_2257,N_2681);
or UO_239 (O_239,N_2399,N_2393);
nor UO_240 (O_240,N_2286,N_2536);
xor UO_241 (O_241,N_2281,N_2413);
nor UO_242 (O_242,N_2926,N_2420);
and UO_243 (O_243,N_2377,N_2537);
nor UO_244 (O_244,N_2386,N_2486);
or UO_245 (O_245,N_2410,N_2754);
and UO_246 (O_246,N_2591,N_2340);
nor UO_247 (O_247,N_2782,N_2471);
and UO_248 (O_248,N_2900,N_2380);
xor UO_249 (O_249,N_2976,N_2706);
or UO_250 (O_250,N_2292,N_2339);
or UO_251 (O_251,N_2729,N_2254);
or UO_252 (O_252,N_2990,N_2977);
nor UO_253 (O_253,N_2464,N_2847);
nand UO_254 (O_254,N_2679,N_2888);
or UO_255 (O_255,N_2898,N_2855);
or UO_256 (O_256,N_2465,N_2427);
nor UO_257 (O_257,N_2457,N_2332);
nand UO_258 (O_258,N_2530,N_2512);
and UO_259 (O_259,N_2376,N_2280);
nand UO_260 (O_260,N_2324,N_2894);
and UO_261 (O_261,N_2825,N_2710);
or UO_262 (O_262,N_2758,N_2351);
and UO_263 (O_263,N_2635,N_2594);
nand UO_264 (O_264,N_2361,N_2751);
or UO_265 (O_265,N_2535,N_2763);
nor UO_266 (O_266,N_2772,N_2998);
nand UO_267 (O_267,N_2671,N_2472);
nor UO_268 (O_268,N_2475,N_2940);
or UO_269 (O_269,N_2529,N_2437);
or UO_270 (O_270,N_2696,N_2266);
and UO_271 (O_271,N_2401,N_2986);
nor UO_272 (O_272,N_2665,N_2874);
and UO_273 (O_273,N_2819,N_2265);
nor UO_274 (O_274,N_2349,N_2250);
or UO_275 (O_275,N_2869,N_2925);
nor UO_276 (O_276,N_2793,N_2561);
nand UO_277 (O_277,N_2881,N_2346);
nand UO_278 (O_278,N_2945,N_2609);
or UO_279 (O_279,N_2890,N_2932);
and UO_280 (O_280,N_2764,N_2712);
nand UO_281 (O_281,N_2545,N_2432);
nor UO_282 (O_282,N_2467,N_2842);
and UO_283 (O_283,N_2605,N_2419);
nor UO_284 (O_284,N_2625,N_2338);
and UO_285 (O_285,N_2691,N_2553);
or UO_286 (O_286,N_2982,N_2807);
nor UO_287 (O_287,N_2551,N_2569);
nand UO_288 (O_288,N_2686,N_2803);
and UO_289 (O_289,N_2962,N_2646);
nand UO_290 (O_290,N_2631,N_2685);
or UO_291 (O_291,N_2400,N_2891);
or UO_292 (O_292,N_2407,N_2492);
nand UO_293 (O_293,N_2919,N_2394);
and UO_294 (O_294,N_2770,N_2730);
or UO_295 (O_295,N_2734,N_2823);
and UO_296 (O_296,N_2628,N_2309);
and UO_297 (O_297,N_2703,N_2688);
nand UO_298 (O_298,N_2623,N_2661);
nor UO_299 (O_299,N_2634,N_2258);
nand UO_300 (O_300,N_2746,N_2577);
and UO_301 (O_301,N_2942,N_2797);
and UO_302 (O_302,N_2580,N_2595);
and UO_303 (O_303,N_2251,N_2440);
nor UO_304 (O_304,N_2538,N_2382);
nand UO_305 (O_305,N_2418,N_2331);
and UO_306 (O_306,N_2552,N_2866);
or UO_307 (O_307,N_2350,N_2378);
nand UO_308 (O_308,N_2708,N_2983);
or UO_309 (O_309,N_2297,N_2738);
or UO_310 (O_310,N_2742,N_2487);
and UO_311 (O_311,N_2417,N_2504);
nor UO_312 (O_312,N_2357,N_2831);
nor UO_313 (O_313,N_2995,N_2355);
nand UO_314 (O_314,N_2658,N_2514);
or UO_315 (O_315,N_2403,N_2927);
nor UO_316 (O_316,N_2507,N_2304);
nand UO_317 (O_317,N_2261,N_2271);
nand UO_318 (O_318,N_2436,N_2904);
nand UO_319 (O_319,N_2395,N_2806);
nand UO_320 (O_320,N_2610,N_2433);
and UO_321 (O_321,N_2789,N_2523);
nor UO_322 (O_322,N_2342,N_2865);
nor UO_323 (O_323,N_2843,N_2352);
nand UO_324 (O_324,N_2690,N_2991);
or UO_325 (O_325,N_2296,N_2446);
or UO_326 (O_326,N_2604,N_2405);
and UO_327 (O_327,N_2820,N_2570);
or UO_328 (O_328,N_2285,N_2496);
nor UO_329 (O_329,N_2640,N_2837);
nor UO_330 (O_330,N_2568,N_2463);
and UO_331 (O_331,N_2711,N_2279);
nand UO_332 (O_332,N_2862,N_2678);
or UO_333 (O_333,N_2905,N_2981);
nand UO_334 (O_334,N_2396,N_2999);
nand UO_335 (O_335,N_2737,N_2556);
or UO_336 (O_336,N_2557,N_2816);
and UO_337 (O_337,N_2384,N_2762);
nor UO_338 (O_338,N_2518,N_2858);
nor UO_339 (O_339,N_2813,N_2829);
and UO_340 (O_340,N_2960,N_2777);
nand UO_341 (O_341,N_2815,N_2818);
nand UO_342 (O_342,N_2425,N_2643);
nand UO_343 (O_343,N_2274,N_2656);
and UO_344 (O_344,N_2844,N_2429);
nor UO_345 (O_345,N_2344,N_2626);
and UO_346 (O_346,N_2878,N_2366);
and UO_347 (O_347,N_2794,N_2760);
or UO_348 (O_348,N_2937,N_2291);
nor UO_349 (O_349,N_2821,N_2294);
and UO_350 (O_350,N_2510,N_2863);
nor UO_351 (O_351,N_2675,N_2335);
or UO_352 (O_352,N_2732,N_2531);
nand UO_353 (O_353,N_2373,N_2476);
and UO_354 (O_354,N_2374,N_2956);
and UO_355 (O_355,N_2502,N_2277);
and UO_356 (O_356,N_2792,N_2805);
and UO_357 (O_357,N_2287,N_2702);
nand UO_358 (O_358,N_2449,N_2362);
and UO_359 (O_359,N_2363,N_2519);
or UO_360 (O_360,N_2462,N_2411);
nor UO_361 (O_361,N_2305,N_2968);
nand UO_362 (O_362,N_2788,N_2500);
and UO_363 (O_363,N_2934,N_2301);
and UO_364 (O_364,N_2322,N_2930);
and UO_365 (O_365,N_2621,N_2884);
or UO_366 (O_366,N_2949,N_2659);
or UO_367 (O_367,N_2630,N_2845);
or UO_368 (O_368,N_2882,N_2714);
nand UO_369 (O_369,N_2911,N_2544);
and UO_370 (O_370,N_2270,N_2459);
nor UO_371 (O_371,N_2966,N_2367);
nor UO_372 (O_372,N_2978,N_2327);
or UO_373 (O_373,N_2719,N_2650);
and UO_374 (O_374,N_2672,N_2872);
nor UO_375 (O_375,N_2791,N_2823);
nor UO_376 (O_376,N_2516,N_2558);
or UO_377 (O_377,N_2590,N_2353);
nor UO_378 (O_378,N_2815,N_2355);
and UO_379 (O_379,N_2950,N_2313);
or UO_380 (O_380,N_2667,N_2696);
nand UO_381 (O_381,N_2726,N_2670);
or UO_382 (O_382,N_2404,N_2428);
nor UO_383 (O_383,N_2801,N_2865);
nor UO_384 (O_384,N_2560,N_2899);
nor UO_385 (O_385,N_2915,N_2593);
or UO_386 (O_386,N_2965,N_2729);
nor UO_387 (O_387,N_2702,N_2780);
nand UO_388 (O_388,N_2990,N_2935);
nand UO_389 (O_389,N_2484,N_2310);
nand UO_390 (O_390,N_2376,N_2969);
nor UO_391 (O_391,N_2631,N_2355);
or UO_392 (O_392,N_2869,N_2831);
nor UO_393 (O_393,N_2506,N_2555);
or UO_394 (O_394,N_2465,N_2668);
and UO_395 (O_395,N_2691,N_2479);
or UO_396 (O_396,N_2383,N_2633);
nand UO_397 (O_397,N_2481,N_2378);
nand UO_398 (O_398,N_2949,N_2962);
and UO_399 (O_399,N_2733,N_2291);
nor UO_400 (O_400,N_2620,N_2992);
and UO_401 (O_401,N_2453,N_2661);
xor UO_402 (O_402,N_2396,N_2748);
and UO_403 (O_403,N_2971,N_2757);
or UO_404 (O_404,N_2523,N_2844);
nor UO_405 (O_405,N_2360,N_2440);
and UO_406 (O_406,N_2774,N_2386);
nor UO_407 (O_407,N_2273,N_2782);
nor UO_408 (O_408,N_2636,N_2503);
or UO_409 (O_409,N_2310,N_2556);
nand UO_410 (O_410,N_2377,N_2876);
or UO_411 (O_411,N_2255,N_2986);
or UO_412 (O_412,N_2960,N_2672);
nor UO_413 (O_413,N_2804,N_2847);
or UO_414 (O_414,N_2405,N_2465);
nor UO_415 (O_415,N_2263,N_2407);
and UO_416 (O_416,N_2894,N_2593);
nand UO_417 (O_417,N_2817,N_2433);
xor UO_418 (O_418,N_2597,N_2602);
and UO_419 (O_419,N_2763,N_2718);
or UO_420 (O_420,N_2789,N_2673);
nor UO_421 (O_421,N_2953,N_2291);
nor UO_422 (O_422,N_2517,N_2652);
and UO_423 (O_423,N_2800,N_2688);
and UO_424 (O_424,N_2372,N_2557);
and UO_425 (O_425,N_2902,N_2494);
and UO_426 (O_426,N_2505,N_2780);
or UO_427 (O_427,N_2683,N_2548);
or UO_428 (O_428,N_2741,N_2946);
nor UO_429 (O_429,N_2767,N_2327);
or UO_430 (O_430,N_2298,N_2413);
nor UO_431 (O_431,N_2312,N_2776);
nand UO_432 (O_432,N_2797,N_2491);
nor UO_433 (O_433,N_2703,N_2584);
and UO_434 (O_434,N_2761,N_2616);
or UO_435 (O_435,N_2899,N_2911);
nand UO_436 (O_436,N_2364,N_2962);
or UO_437 (O_437,N_2601,N_2257);
and UO_438 (O_438,N_2903,N_2799);
and UO_439 (O_439,N_2568,N_2923);
nand UO_440 (O_440,N_2698,N_2335);
nand UO_441 (O_441,N_2474,N_2891);
and UO_442 (O_442,N_2856,N_2927);
nor UO_443 (O_443,N_2441,N_2956);
or UO_444 (O_444,N_2576,N_2654);
nand UO_445 (O_445,N_2528,N_2265);
or UO_446 (O_446,N_2999,N_2267);
nor UO_447 (O_447,N_2518,N_2348);
nand UO_448 (O_448,N_2702,N_2418);
xnor UO_449 (O_449,N_2913,N_2806);
and UO_450 (O_450,N_2667,N_2694);
and UO_451 (O_451,N_2626,N_2447);
and UO_452 (O_452,N_2383,N_2426);
nand UO_453 (O_453,N_2786,N_2931);
or UO_454 (O_454,N_2544,N_2822);
and UO_455 (O_455,N_2646,N_2935);
and UO_456 (O_456,N_2939,N_2407);
nand UO_457 (O_457,N_2786,N_2809);
nor UO_458 (O_458,N_2869,N_2658);
or UO_459 (O_459,N_2261,N_2481);
or UO_460 (O_460,N_2323,N_2835);
xnor UO_461 (O_461,N_2495,N_2825);
nand UO_462 (O_462,N_2777,N_2570);
or UO_463 (O_463,N_2287,N_2902);
nor UO_464 (O_464,N_2881,N_2825);
and UO_465 (O_465,N_2883,N_2696);
and UO_466 (O_466,N_2250,N_2542);
nor UO_467 (O_467,N_2987,N_2790);
nor UO_468 (O_468,N_2816,N_2573);
xor UO_469 (O_469,N_2416,N_2515);
and UO_470 (O_470,N_2892,N_2296);
nor UO_471 (O_471,N_2302,N_2445);
nand UO_472 (O_472,N_2700,N_2282);
or UO_473 (O_473,N_2984,N_2282);
nand UO_474 (O_474,N_2445,N_2818);
nand UO_475 (O_475,N_2277,N_2752);
or UO_476 (O_476,N_2819,N_2982);
nor UO_477 (O_477,N_2948,N_2404);
nand UO_478 (O_478,N_2760,N_2277);
nand UO_479 (O_479,N_2268,N_2960);
or UO_480 (O_480,N_2374,N_2748);
nor UO_481 (O_481,N_2343,N_2896);
or UO_482 (O_482,N_2892,N_2602);
nand UO_483 (O_483,N_2911,N_2348);
nand UO_484 (O_484,N_2387,N_2608);
and UO_485 (O_485,N_2604,N_2456);
or UO_486 (O_486,N_2903,N_2269);
and UO_487 (O_487,N_2857,N_2661);
nor UO_488 (O_488,N_2507,N_2264);
nand UO_489 (O_489,N_2760,N_2616);
or UO_490 (O_490,N_2352,N_2689);
nand UO_491 (O_491,N_2975,N_2283);
and UO_492 (O_492,N_2704,N_2302);
nor UO_493 (O_493,N_2728,N_2313);
nand UO_494 (O_494,N_2970,N_2871);
and UO_495 (O_495,N_2974,N_2681);
or UO_496 (O_496,N_2507,N_2793);
or UO_497 (O_497,N_2655,N_2825);
nor UO_498 (O_498,N_2833,N_2769);
and UO_499 (O_499,N_2305,N_2639);
endmodule