module basic_1500_15000_2000_60_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_886,In_26);
nand U1 (N_1,In_1385,In_1114);
nand U2 (N_2,In_1454,In_994);
and U3 (N_3,In_983,In_1029);
or U4 (N_4,In_960,In_464);
or U5 (N_5,In_372,In_1121);
nand U6 (N_6,In_229,In_9);
xor U7 (N_7,In_1178,In_173);
xnor U8 (N_8,In_681,In_1224);
nor U9 (N_9,In_882,In_210);
nor U10 (N_10,In_22,In_530);
nand U11 (N_11,In_680,In_567);
or U12 (N_12,In_1186,In_759);
nor U13 (N_13,In_1147,In_28);
nand U14 (N_14,In_1490,In_866);
or U15 (N_15,In_1372,In_70);
nand U16 (N_16,In_1395,In_671);
nand U17 (N_17,In_1314,In_1246);
xnor U18 (N_18,In_170,In_1280);
or U19 (N_19,In_870,In_390);
nand U20 (N_20,In_590,In_1024);
nor U21 (N_21,In_1034,In_1358);
xor U22 (N_22,In_830,In_1321);
nor U23 (N_23,In_1455,In_1084);
xor U24 (N_24,In_1146,In_754);
nor U25 (N_25,In_1202,In_1182);
nand U26 (N_26,In_1165,In_48);
nor U27 (N_27,In_956,In_1258);
xnor U28 (N_28,In_60,In_1039);
and U29 (N_29,In_1279,In_612);
and U30 (N_30,In_11,In_1016);
nand U31 (N_31,In_230,In_340);
nand U32 (N_32,In_44,In_1278);
nor U33 (N_33,In_88,In_371);
xor U34 (N_34,In_441,In_1036);
nand U35 (N_35,In_707,In_226);
xor U36 (N_36,In_138,In_1382);
nand U37 (N_37,In_72,In_1307);
and U38 (N_38,In_423,In_302);
nand U39 (N_39,In_768,In_402);
nand U40 (N_40,In_770,In_1320);
xnor U41 (N_41,In_510,In_1298);
and U42 (N_42,In_110,In_359);
xor U43 (N_43,In_223,In_731);
nand U44 (N_44,In_512,In_858);
nor U45 (N_45,In_431,In_1379);
nor U46 (N_46,In_664,In_318);
or U47 (N_47,In_1331,In_1119);
nor U48 (N_48,In_96,In_381);
or U49 (N_49,In_500,In_42);
and U50 (N_50,In_191,In_967);
xnor U51 (N_51,In_1482,In_255);
xor U52 (N_52,In_1388,In_1152);
xnor U53 (N_53,In_1135,In_535);
nor U54 (N_54,In_533,In_135);
and U55 (N_55,In_880,In_102);
or U56 (N_56,In_74,In_373);
nor U57 (N_57,In_166,In_41);
or U58 (N_58,In_594,In_1444);
xnor U59 (N_59,In_1412,In_288);
xnor U60 (N_60,In_274,In_905);
nor U61 (N_61,In_1479,In_985);
and U62 (N_62,In_1498,In_5);
nor U63 (N_63,In_774,In_591);
and U64 (N_64,In_851,In_128);
nand U65 (N_65,In_696,In_649);
or U66 (N_66,In_1425,In_669);
nand U67 (N_67,In_1212,In_3);
nand U68 (N_68,In_730,In_311);
and U69 (N_69,In_1335,In_1373);
nor U70 (N_70,In_137,In_293);
and U71 (N_71,In_1023,In_1148);
or U72 (N_72,In_146,In_1248);
or U73 (N_73,In_876,In_1160);
nand U74 (N_74,In_1435,In_805);
nand U75 (N_75,In_623,In_1122);
or U76 (N_76,In_183,In_699);
and U77 (N_77,In_1304,In_838);
nand U78 (N_78,In_747,In_843);
xor U79 (N_79,In_704,In_679);
nor U80 (N_80,In_111,In_122);
nand U81 (N_81,In_321,In_1090);
or U82 (N_82,In_94,In_1459);
xor U83 (N_83,In_239,In_1215);
xor U84 (N_84,In_27,In_234);
xnor U85 (N_85,In_853,In_712);
xnor U86 (N_86,In_1472,In_250);
xor U87 (N_87,In_1339,In_143);
xnor U88 (N_88,In_240,In_236);
and U89 (N_89,In_605,In_1274);
and U90 (N_90,In_1190,In_1452);
xnor U91 (N_91,In_844,In_124);
xnor U92 (N_92,In_663,In_1230);
or U93 (N_93,In_65,In_557);
or U94 (N_94,In_201,In_587);
nor U95 (N_95,In_1447,In_618);
nor U96 (N_96,In_1004,In_30);
and U97 (N_97,In_4,In_803);
or U98 (N_98,In_962,In_452);
nor U99 (N_99,In_499,In_1077);
and U100 (N_100,In_198,In_1170);
and U101 (N_101,In_442,In_936);
nand U102 (N_102,In_192,In_763);
nor U103 (N_103,In_1465,In_369);
xnor U104 (N_104,In_511,In_1464);
nand U105 (N_105,In_523,In_1351);
nor U106 (N_106,In_912,In_46);
nor U107 (N_107,In_1326,In_583);
and U108 (N_108,In_534,In_775);
or U109 (N_109,In_1345,In_465);
and U110 (N_110,In_569,In_168);
or U111 (N_111,In_1021,In_907);
xor U112 (N_112,In_329,In_453);
nand U113 (N_113,In_315,In_644);
or U114 (N_114,In_175,In_1386);
nor U115 (N_115,In_490,In_113);
or U116 (N_116,In_194,In_826);
or U117 (N_117,In_847,In_331);
nor U118 (N_118,In_517,In_1242);
and U119 (N_119,In_1073,In_1245);
xnor U120 (N_120,In_212,In_1002);
xnor U121 (N_121,In_751,In_131);
and U122 (N_122,In_909,In_502);
nor U123 (N_123,In_335,In_1141);
or U124 (N_124,In_613,In_1275);
nor U125 (N_125,In_1474,In_935);
nor U126 (N_126,In_134,In_1154);
and U127 (N_127,In_932,In_29);
and U128 (N_128,In_1456,In_1268);
nor U129 (N_129,In_368,In_364);
xor U130 (N_130,In_1101,In_1204);
and U131 (N_131,In_1005,In_547);
nor U132 (N_132,In_690,In_1017);
xor U133 (N_133,In_616,In_237);
and U134 (N_134,In_1302,In_185);
or U135 (N_135,In_1033,In_596);
nand U136 (N_136,In_455,In_1362);
nand U137 (N_137,In_456,In_692);
nor U138 (N_138,In_1257,In_1006);
nor U139 (N_139,In_548,In_790);
and U140 (N_140,In_560,In_773);
nor U141 (N_141,In_758,In_1111);
and U142 (N_142,In_689,In_1167);
or U143 (N_143,In_881,In_1255);
nor U144 (N_144,In_1284,In_1266);
nor U145 (N_145,In_225,In_1193);
xor U146 (N_146,In_1468,In_808);
nor U147 (N_147,In_1380,In_492);
or U148 (N_148,In_737,In_1422);
nor U149 (N_149,In_1066,In_559);
xor U150 (N_150,In_1420,In_732);
xor U151 (N_151,In_307,In_1003);
nor U152 (N_152,In_743,In_1007);
and U153 (N_153,In_1329,In_889);
nor U154 (N_154,In_718,In_148);
nand U155 (N_155,In_1070,In_670);
nand U156 (N_156,In_894,In_509);
xor U157 (N_157,In_984,In_1383);
xnor U158 (N_158,In_18,In_314);
nand U159 (N_159,In_1060,In_133);
xor U160 (N_160,In_728,In_450);
and U161 (N_161,In_589,In_606);
nand U162 (N_162,In_1113,In_277);
and U163 (N_163,In_604,In_325);
xnor U164 (N_164,In_541,In_103);
xor U165 (N_165,In_1356,In_546);
nor U166 (N_166,In_387,In_834);
xor U167 (N_167,In_1461,In_127);
and U168 (N_168,In_1423,In_682);
nor U169 (N_169,In_823,In_1236);
nand U170 (N_170,In_572,In_933);
and U171 (N_171,In_922,In_697);
or U172 (N_172,In_1120,In_640);
xor U173 (N_173,In_981,In_955);
nor U174 (N_174,In_801,In_193);
and U175 (N_175,In_419,In_1471);
nor U176 (N_176,In_980,In_388);
nor U177 (N_177,In_405,In_1201);
nor U178 (N_178,In_484,In_1475);
or U179 (N_179,In_645,In_429);
xor U180 (N_180,In_323,In_873);
nand U181 (N_181,In_1262,In_1071);
or U182 (N_182,In_875,In_762);
nand U183 (N_183,In_1384,In_1306);
nand U184 (N_184,In_614,In_351);
nand U185 (N_185,In_37,In_352);
or U186 (N_186,In_1225,In_64);
nand U187 (N_187,In_1166,In_472);
nor U188 (N_188,In_538,In_228);
nor U189 (N_189,In_518,In_156);
xor U190 (N_190,In_1484,In_913);
xnor U191 (N_191,In_347,In_1401);
or U192 (N_192,In_693,In_1183);
nand U193 (N_193,In_1238,In_1042);
nand U194 (N_194,In_1481,In_1237);
xor U195 (N_195,In_992,In_1157);
nor U196 (N_196,In_516,In_1429);
xnor U197 (N_197,In_184,In_169);
and U198 (N_198,In_1011,In_1000);
and U199 (N_199,In_711,In_622);
and U200 (N_200,In_678,In_17);
or U201 (N_201,In_241,In_601);
nand U202 (N_202,In_954,In_446);
nand U203 (N_203,In_920,In_982);
nor U204 (N_204,In_24,In_1228);
and U205 (N_205,In_100,In_675);
nand U206 (N_206,In_440,In_1416);
nor U207 (N_207,In_969,In_1098);
or U208 (N_208,In_1174,In_1199);
nand U209 (N_209,In_190,In_488);
and U210 (N_210,In_1480,In_1436);
or U211 (N_211,In_709,In_887);
or U212 (N_212,In_800,In_741);
nor U213 (N_213,In_1001,In_1316);
nand U214 (N_214,In_764,In_471);
xnor U215 (N_215,In_745,In_1318);
nor U216 (N_216,In_459,In_911);
nor U217 (N_217,In_67,In_217);
and U218 (N_218,In_726,In_1270);
nor U219 (N_219,In_330,In_1359);
xor U220 (N_220,In_656,In_69);
nand U221 (N_221,In_1376,In_333);
or U222 (N_222,In_610,In_1408);
nor U223 (N_223,In_1085,In_344);
nand U224 (N_224,In_1108,In_47);
xnor U225 (N_225,In_566,In_326);
xnor U226 (N_226,In_1308,In_427);
nand U227 (N_227,In_460,In_1281);
nor U228 (N_228,In_80,In_813);
or U229 (N_229,In_370,In_1404);
nor U230 (N_230,In_418,In_410);
and U231 (N_231,In_698,In_821);
nand U232 (N_232,In_97,In_301);
and U233 (N_233,In_468,In_537);
xnor U234 (N_234,In_1325,In_434);
nor U235 (N_235,In_1430,In_729);
nor U236 (N_236,In_574,In_508);
xor U237 (N_237,In_82,In_871);
nor U238 (N_238,In_1293,In_683);
nor U239 (N_239,In_897,In_998);
xnor U240 (N_240,In_38,In_973);
nor U241 (N_241,In_104,In_898);
nand U242 (N_242,In_422,In_755);
xor U243 (N_243,In_467,In_1232);
nand U244 (N_244,In_1463,In_1428);
xor U245 (N_245,In_172,In_345);
and U246 (N_246,In_1453,In_761);
nand U247 (N_247,In_87,In_673);
nor U248 (N_248,In_896,In_890);
nand U249 (N_249,In_585,In_959);
or U250 (N_250,In_145,In_792);
or U251 (N_251,In_568,In_458);
xor U252 (N_252,In_32,In_1297);
nor U253 (N_253,N_97,In_109);
xnor U254 (N_254,N_2,In_353);
xor U255 (N_255,In_1451,In_862);
and U256 (N_256,In_501,In_1322);
and U257 (N_257,In_908,In_86);
or U258 (N_258,In_375,In_186);
xor U259 (N_259,In_494,In_931);
xor U260 (N_260,In_1159,In_174);
or U261 (N_261,N_94,In_810);
or U262 (N_262,In_859,In_924);
nor U263 (N_263,In_106,In_1068);
nand U264 (N_264,N_156,In_1432);
xnor U265 (N_265,N_56,In_925);
or U266 (N_266,In_725,In_970);
and U267 (N_267,In_396,In_1264);
and U268 (N_268,In_1483,In_1427);
or U269 (N_269,In_398,In_1125);
nor U270 (N_270,In_1049,In_1218);
nor U271 (N_271,In_401,In_308);
nand U272 (N_272,In_178,In_1124);
xor U273 (N_273,In_1226,In_233);
nand U274 (N_274,In_654,In_1406);
and U275 (N_275,In_2,In_556);
and U276 (N_276,N_126,In_62);
nor U277 (N_277,In_147,In_634);
and U278 (N_278,In_550,In_1038);
nand U279 (N_279,N_201,In_575);
or U280 (N_280,N_32,In_638);
xor U281 (N_281,In_378,In_1243);
nor U282 (N_282,In_611,In_940);
or U283 (N_283,In_577,In_828);
nand U284 (N_284,In_286,In_365);
nand U285 (N_285,N_21,In_1263);
xor U286 (N_286,In_1219,In_337);
xnor U287 (N_287,In_938,In_245);
or U288 (N_288,In_1151,In_159);
xnor U289 (N_289,In_1348,In_1249);
nand U290 (N_290,N_212,In_626);
and U291 (N_291,N_39,In_1233);
nor U292 (N_292,In_1025,In_632);
xnor U293 (N_293,N_53,In_901);
and U294 (N_294,In_619,In_267);
and U295 (N_295,In_287,In_305);
or U296 (N_296,In_714,In_73);
and U297 (N_297,In_794,In_1450);
nor U298 (N_298,In_785,In_688);
or U299 (N_299,In_1256,In_179);
and U300 (N_300,In_385,In_141);
nor U301 (N_301,In_1391,In_529);
nor U302 (N_302,In_904,In_476);
and U303 (N_303,In_701,N_81);
nor U304 (N_304,In_1493,In_625);
nor U305 (N_305,In_408,N_6);
nand U306 (N_306,In_531,In_310);
nor U307 (N_307,In_657,In_99);
xor U308 (N_308,In_343,In_636);
or U309 (N_309,In_1327,In_1171);
nand U310 (N_310,In_295,N_36);
nand U311 (N_311,In_397,In_1305);
or U312 (N_312,In_421,In_139);
and U313 (N_313,In_85,In_571);
nand U314 (N_314,In_1466,N_38);
nand U315 (N_315,In_439,N_112);
nand U316 (N_316,In_51,In_514);
nand U317 (N_317,N_225,In_1487);
and U318 (N_318,In_676,In_1300);
and U319 (N_319,In_1374,In_266);
and U320 (N_320,N_135,In_1096);
or U321 (N_321,In_760,In_766);
nand U322 (N_322,In_197,In_665);
nor U323 (N_323,In_167,In_341);
xor U324 (N_324,In_395,In_1069);
and U325 (N_325,In_1221,In_1074);
xnor U326 (N_326,In_1413,In_1499);
nand U327 (N_327,In_1240,In_642);
xor U328 (N_328,N_204,In_915);
nand U329 (N_329,In_927,In_171);
nand U330 (N_330,In_1433,In_1330);
nand U331 (N_331,In_842,In_1295);
or U332 (N_332,In_921,In_469);
nand U333 (N_333,In_75,In_1045);
and U334 (N_334,N_84,In_1030);
xor U335 (N_335,In_1092,In_668);
and U336 (N_336,In_1375,In_519);
or U337 (N_337,In_45,In_1417);
and U338 (N_338,N_207,N_198);
nand U339 (N_339,In_154,In_1013);
nor U340 (N_340,N_186,In_1477);
xor U341 (N_341,In_979,N_158);
and U342 (N_342,In_637,N_222);
nand U343 (N_343,In_89,In_542);
nor U344 (N_344,In_482,N_190);
nor U345 (N_345,In_58,In_1273);
xnor U346 (N_346,In_449,In_1291);
or U347 (N_347,In_809,In_362);
nand U348 (N_348,In_653,N_110);
or U349 (N_349,In_463,In_961);
or U350 (N_350,In_1008,In_328);
and U351 (N_351,N_169,N_119);
or U352 (N_352,N_34,In_687);
xor U353 (N_353,In_56,In_116);
and U354 (N_354,N_46,In_462);
nand U355 (N_355,In_1253,N_168);
nor U356 (N_356,In_608,In_448);
nor U357 (N_357,In_1462,In_1100);
or U358 (N_358,In_1040,In_735);
or U359 (N_359,N_147,N_12);
and U360 (N_360,In_1019,In_406);
or U361 (N_361,In_1043,In_425);
xnor U362 (N_362,In_23,In_1115);
nor U363 (N_363,In_1261,In_1217);
and U364 (N_364,N_47,In_1173);
and U365 (N_365,In_1223,In_316);
or U366 (N_366,In_1449,In_1445);
xor U367 (N_367,N_24,N_143);
nor U368 (N_368,In_424,In_1099);
and U369 (N_369,In_659,In_0);
xor U370 (N_370,In_702,N_137);
nand U371 (N_371,In_1180,In_98);
xnor U372 (N_372,N_130,In_350);
or U373 (N_373,In_1347,In_1343);
and U374 (N_374,In_498,N_245);
nor U375 (N_375,In_812,In_885);
and U376 (N_376,In_674,In_919);
nor U377 (N_377,In_746,In_1290);
or U378 (N_378,In_1185,N_209);
nand U379 (N_379,In_923,In_1250);
nand U380 (N_380,N_68,N_159);
or U381 (N_381,In_631,N_98);
nor U382 (N_382,N_19,In_1053);
or U383 (N_383,N_140,In_480);
nand U384 (N_384,In_987,N_44);
nor U385 (N_385,N_174,In_263);
nor U386 (N_386,N_22,In_195);
nand U387 (N_387,In_748,In_666);
nor U388 (N_388,In_515,N_181);
and U389 (N_389,In_1355,In_276);
or U390 (N_390,In_617,In_878);
and U391 (N_391,In_1350,In_1370);
nand U392 (N_392,In_1244,In_835);
xnor U393 (N_393,In_78,In_1198);
and U394 (N_394,In_1047,In_312);
xnor U395 (N_395,N_107,In_322);
nand U396 (N_396,In_164,In_261);
or U397 (N_397,In_68,In_953);
nor U398 (N_398,N_229,In_946);
nor U399 (N_399,In_879,N_45);
nor U400 (N_400,In_214,In_1087);
nand U401 (N_401,In_238,In_750);
nor U402 (N_402,In_443,In_119);
nand U403 (N_403,In_61,In_162);
or U404 (N_404,In_121,In_817);
and U405 (N_405,In_767,N_191);
nor U406 (N_406,In_1442,In_265);
or U407 (N_407,In_1488,N_35);
nand U408 (N_408,In_202,In_1207);
nor U409 (N_409,In_1353,In_997);
and U410 (N_410,N_141,In_120);
xor U411 (N_411,In_1426,N_90);
and U412 (N_412,In_1133,In_1368);
nand U413 (N_413,In_420,In_1138);
xnor U414 (N_414,In_968,In_220);
xnor U415 (N_415,In_151,In_695);
xor U416 (N_416,In_1323,In_1402);
nor U417 (N_417,In_1315,In_1407);
nand U418 (N_418,In_1153,In_1272);
or U419 (N_419,N_184,In_34);
or U420 (N_420,N_134,In_965);
xor U421 (N_421,In_971,In_700);
xor U422 (N_422,N_132,In_734);
or U423 (N_423,In_1360,In_112);
or U424 (N_424,In_526,In_521);
nand U425 (N_425,In_1282,In_1142);
nor U426 (N_426,In_1048,In_327);
or U427 (N_427,In_855,In_1081);
and U428 (N_428,In_224,N_155);
or U429 (N_429,In_1076,In_1392);
or U430 (N_430,In_1075,In_436);
or U431 (N_431,In_902,In_1285);
xor U432 (N_432,N_188,In_1156);
or U433 (N_433,N_120,N_208);
and U434 (N_434,N_62,N_128);
and U435 (N_435,N_226,In_1018);
nand U436 (N_436,In_84,In_244);
and U437 (N_437,N_117,In_457);
nor U438 (N_438,In_272,N_187);
or U439 (N_439,N_11,In_651);
nand U440 (N_440,In_749,In_495);
and U441 (N_441,In_600,In_248);
nand U442 (N_442,In_564,In_403);
nor U443 (N_443,In_713,In_1057);
or U444 (N_444,In_1032,In_807);
nor U445 (N_445,In_273,In_740);
xnor U446 (N_446,N_3,In_991);
or U447 (N_447,In_1126,In_1390);
xnor U448 (N_448,In_1381,In_966);
nor U449 (N_449,In_796,In_757);
and U450 (N_450,In_339,In_1162);
and U451 (N_451,In_716,In_602);
nor U452 (N_452,In_1220,In_95);
and U453 (N_453,N_164,N_9);
and U454 (N_454,In_140,In_182);
nor U455 (N_455,In_1163,In_187);
nand U456 (N_456,In_565,N_172);
xnor U457 (N_457,In_477,In_1118);
or U458 (N_458,In_1104,In_125);
or U459 (N_459,In_504,In_204);
or U460 (N_460,In_551,In_818);
nand U461 (N_461,In_283,In_545);
nor U462 (N_462,In_1334,N_31);
and U463 (N_463,In_856,In_1341);
nor U464 (N_464,In_802,N_234);
or U465 (N_465,In_950,N_221);
or U466 (N_466,In_386,In_435);
and U467 (N_467,N_118,In_799);
nand U468 (N_468,In_281,In_466);
nand U469 (N_469,In_354,In_570);
xor U470 (N_470,N_129,In_1411);
nor U471 (N_471,In_285,In_415);
nor U472 (N_472,N_102,In_1378);
nor U473 (N_473,In_366,N_217);
xor U474 (N_474,In_55,In_708);
nand U475 (N_475,In_358,In_189);
and U476 (N_476,In_1409,In_93);
nand U477 (N_477,In_216,N_86);
nand U478 (N_478,In_742,In_1333);
or U479 (N_479,In_1132,In_863);
nand U480 (N_480,In_1441,In_181);
xor U481 (N_481,In_1400,In_6);
and U482 (N_482,In_493,In_836);
and U483 (N_483,In_771,In_660);
or U484 (N_484,In_822,N_29);
nor U485 (N_485,In_685,In_271);
and U486 (N_486,In_264,In_1206);
nand U487 (N_487,In_363,In_643);
nand U488 (N_488,In_756,In_1399);
nor U489 (N_489,In_357,In_1168);
and U490 (N_490,N_139,In_411);
xnor U491 (N_491,N_104,In_739);
or U492 (N_492,In_1403,N_166);
nand U493 (N_493,In_588,In_157);
xnor U494 (N_494,In_1150,In_989);
nor U495 (N_495,In_1421,In_129);
nor U496 (N_496,In_126,In_655);
and U497 (N_497,In_1061,In_815);
and U498 (N_498,N_218,In_753);
or U499 (N_499,In_1496,In_1110);
nor U500 (N_500,N_310,In_672);
and U501 (N_501,N_228,In_941);
and U502 (N_502,In_845,N_269);
nor U503 (N_503,In_1009,In_21);
or U504 (N_504,In_1095,In_360);
or U505 (N_505,In_661,N_333);
nand U506 (N_506,In_1363,In_1397);
and U507 (N_507,N_291,In_470);
and U508 (N_508,N_216,N_152);
nand U509 (N_509,N_450,N_248);
or U510 (N_510,N_493,N_469);
and U511 (N_511,In_294,N_96);
nor U512 (N_512,N_205,In_487);
and U513 (N_513,In_79,N_111);
nor U514 (N_514,In_389,In_1080);
nand U515 (N_515,N_392,N_393);
or U516 (N_516,In_999,In_1396);
or U517 (N_517,In_83,In_1079);
and U518 (N_518,In_483,In_1062);
xor U519 (N_519,In_417,In_624);
and U520 (N_520,N_394,N_412);
xor U521 (N_521,N_271,N_286);
nor U522 (N_522,N_432,In_877);
nor U523 (N_523,In_12,In_444);
nand U524 (N_524,In_957,N_138);
or U525 (N_525,In_320,In_52);
nand U526 (N_526,In_426,In_719);
and U527 (N_527,In_14,In_278);
nand U528 (N_528,N_335,In_917);
nand U529 (N_529,N_452,N_327);
and U530 (N_530,In_235,In_1);
nand U531 (N_531,N_79,In_1222);
xnor U532 (N_532,In_780,In_1319);
xor U533 (N_533,N_320,In_1414);
nor U534 (N_534,N_364,N_268);
nor U535 (N_535,In_290,N_363);
nor U536 (N_536,In_1424,N_379);
or U537 (N_537,In_163,N_480);
nand U538 (N_538,N_325,N_448);
nor U539 (N_539,N_14,N_421);
and U540 (N_540,In_952,In_1489);
or U541 (N_541,N_264,In_486);
xor U542 (N_542,N_332,In_399);
and U543 (N_543,N_57,In_752);
nor U544 (N_544,In_1234,In_1271);
or U545 (N_545,In_218,N_416);
nor U546 (N_546,In_769,N_437);
and U547 (N_547,In_528,In_841);
nand U548 (N_548,N_293,In_652);
nand U549 (N_549,N_37,In_1044);
nor U550 (N_550,In_1254,In_597);
nor U551 (N_551,In_1063,N_58);
nand U552 (N_552,In_860,In_848);
nor U553 (N_553,In_781,In_576);
nor U554 (N_554,In_1097,N_492);
nor U555 (N_555,In_1265,In_1169);
nand U556 (N_556,In_393,N_179);
nor U557 (N_557,N_125,N_40);
nand U558 (N_558,N_481,N_103);
nand U559 (N_559,N_280,N_429);
xnor U560 (N_560,In_945,N_183);
nand U561 (N_561,N_321,In_520);
or U562 (N_562,In_827,N_91);
nor U563 (N_563,In_231,In_1189);
nor U564 (N_564,N_304,In_804);
nor U565 (N_565,N_459,N_76);
nand U566 (N_566,N_100,In_1094);
nand U567 (N_567,In_667,In_1418);
and U568 (N_568,N_465,In_474);
nor U569 (N_569,In_1393,In_491);
and U570 (N_570,In_1188,In_485);
nand U571 (N_571,N_471,N_454);
and U572 (N_572,In_787,In_1103);
and U573 (N_573,N_52,In_1145);
and U574 (N_574,N_163,N_220);
nor U575 (N_575,In_1469,In_279);
xor U576 (N_576,In_888,In_1184);
xor U577 (N_577,N_256,N_238);
xor U578 (N_578,In_149,In_382);
xnor U579 (N_579,In_130,In_144);
or U580 (N_580,In_1497,N_415);
nor U581 (N_581,N_298,In_1203);
nor U582 (N_582,In_795,In_153);
or U583 (N_583,In_778,In_686);
and U584 (N_584,In_1352,N_235);
and U585 (N_585,N_242,In_40);
or U586 (N_586,N_230,In_479);
xnor U587 (N_587,In_1313,N_177);
nor U588 (N_588,N_337,In_246);
or U589 (N_589,In_1143,N_385);
or U590 (N_590,In_926,N_193);
nand U591 (N_591,In_1294,N_367);
or U592 (N_592,N_476,N_439);
nand U593 (N_593,In_35,In_1210);
or U594 (N_594,N_323,N_306);
or U595 (N_595,In_105,N_60);
nand U596 (N_596,N_380,In_662);
nand U597 (N_597,In_1078,In_1083);
xnor U598 (N_598,N_106,In_414);
xnor U599 (N_599,N_498,N_244);
and U600 (N_600,In_20,In_303);
nor U601 (N_601,In_832,N_252);
and U602 (N_602,In_937,N_356);
nand U603 (N_603,N_478,N_383);
nor U604 (N_604,In_1139,In_868);
xnor U605 (N_605,N_449,N_28);
nand U606 (N_606,N_485,In_221);
and U607 (N_607,In_864,In_1035);
nor U608 (N_608,In_789,In_816);
and U609 (N_609,N_440,N_369);
nor U610 (N_610,In_1288,N_301);
nor U611 (N_611,In_503,N_438);
or U612 (N_612,In_1289,In_1410);
xor U613 (N_613,N_223,In_1247);
nor U614 (N_614,In_391,N_266);
and U615 (N_615,In_188,N_425);
nor U616 (N_616,N_355,N_237);
and U617 (N_617,In_1340,In_438);
nor U618 (N_618,N_59,N_414);
and U619 (N_619,In_25,N_289);
or U620 (N_620,N_341,N_292);
or U621 (N_621,N_463,In_797);
nand U622 (N_622,In_282,N_313);
xnor U623 (N_623,In_497,N_247);
or U624 (N_624,In_506,In_1072);
and U625 (N_625,N_381,N_210);
or U626 (N_626,N_307,N_257);
or U627 (N_627,In_684,In_1181);
and U628 (N_628,In_1357,In_861);
xnor U629 (N_629,N_142,N_386);
xor U630 (N_630,In_553,In_1089);
nor U631 (N_631,N_300,In_66);
and U632 (N_632,In_703,N_487);
nand U633 (N_633,In_304,In_1056);
nand U634 (N_634,In_152,In_782);
nor U635 (N_635,In_691,In_409);
and U636 (N_636,N_5,In_1136);
or U637 (N_637,N_93,In_209);
nand U638 (N_638,In_1052,In_289);
xnor U639 (N_639,N_115,In_1312);
nor U640 (N_640,N_302,In_791);
nor U641 (N_641,In_300,In_160);
nand U642 (N_642,In_208,N_354);
or U643 (N_643,N_352,In_213);
xnor U644 (N_644,N_423,In_615);
xor U645 (N_645,N_262,N_467);
nor U646 (N_646,In_1050,In_1354);
or U647 (N_647,In_1259,N_274);
xor U648 (N_648,In_211,N_288);
or U649 (N_649,N_275,N_258);
nor U650 (N_650,In_91,N_443);
nor U651 (N_651,In_1292,In_819);
nor U652 (N_652,In_1277,In_296);
nand U653 (N_653,N_294,N_430);
xor U654 (N_654,In_247,In_249);
or U655 (N_655,In_738,N_494);
or U656 (N_656,N_399,In_275);
nor U657 (N_657,N_334,In_15);
and U658 (N_658,N_150,In_1387);
and U659 (N_659,In_1491,In_1064);
nor U660 (N_660,N_71,N_77);
and U661 (N_661,N_175,In_219);
nand U662 (N_662,N_417,In_478);
nand U663 (N_663,In_1310,N_233);
and U664 (N_664,N_388,In_196);
and U665 (N_665,In_1349,In_177);
nand U666 (N_666,In_852,In_1229);
nor U667 (N_667,N_284,N_251);
xnor U668 (N_668,In_906,In_806);
nor U669 (N_669,In_203,In_1067);
and U670 (N_670,N_374,In_1046);
or U671 (N_671,N_466,N_296);
or U672 (N_672,In_586,N_146);
nor U673 (N_673,In_1200,In_706);
nor U674 (N_674,N_281,In_39);
nand U675 (N_675,N_124,In_1485);
or U676 (N_676,In_1187,N_263);
or U677 (N_677,N_336,N_371);
xnor U678 (N_678,In_1195,In_944);
or U679 (N_679,N_199,In_1431);
xor U680 (N_680,N_42,N_206);
xnor U681 (N_681,N_203,In_496);
or U682 (N_682,In_394,In_895);
nor U683 (N_683,N_23,In_1155);
xnor U684 (N_684,In_1311,N_458);
or U685 (N_685,N_391,In_8);
and U686 (N_686,N_197,N_189);
nor U687 (N_687,In_977,In_1065);
nand U688 (N_688,In_1051,In_833);
nand U689 (N_689,In_1296,N_8);
and U690 (N_690,N_330,In_658);
nor U691 (N_691,N_488,In_1389);
and U692 (N_692,In_599,In_598);
xnor U693 (N_693,N_87,In_840);
or U694 (N_694,In_727,In_939);
nand U695 (N_695,In_227,N_473);
nand U696 (N_696,N_477,In_1022);
or U697 (N_697,In_580,N_185);
or U698 (N_698,In_527,N_372);
xor U699 (N_699,N_462,In_1058);
xor U700 (N_700,In_1239,In_1054);
nor U701 (N_701,In_475,N_444);
xor U702 (N_702,In_1235,In_1439);
nor U703 (N_703,In_1309,In_200);
and U704 (N_704,In_257,In_951);
and U705 (N_705,In_1107,N_460);
or U706 (N_706,In_621,In_284);
xor U707 (N_707,In_1020,In_558);
nand U708 (N_708,In_507,N_312);
nor U709 (N_709,In_313,In_1283);
xor U710 (N_710,N_420,In_891);
xnor U711 (N_711,In_607,N_495);
and U712 (N_712,N_231,N_67);
xor U713 (N_713,In_473,In_332);
and U714 (N_714,In_581,N_30);
or U715 (N_715,In_650,In_81);
and U716 (N_716,N_105,N_18);
nand U717 (N_717,N_161,In_1377);
nor U718 (N_718,In_380,N_136);
and U719 (N_719,In_1082,In_736);
nand U720 (N_720,In_540,In_633);
or U721 (N_721,N_196,In_628);
or U722 (N_722,N_80,In_1317);
nor U723 (N_723,In_258,In_630);
and U724 (N_724,In_1026,N_99);
and U725 (N_725,In_1332,N_360);
nand U726 (N_726,N_171,In_505);
nor U727 (N_727,In_1369,N_26);
and U728 (N_728,N_27,N_315);
nor U729 (N_729,In_280,In_1192);
or U730 (N_730,In_33,N_116);
xor U731 (N_731,N_389,In_1116);
nor U732 (N_732,N_422,N_376);
xor U733 (N_733,N_162,N_431);
nand U734 (N_734,N_456,N_249);
xnor U735 (N_735,N_121,N_377);
nand U736 (N_736,In_71,In_555);
and U737 (N_737,In_379,N_362);
nor U738 (N_738,In_1196,In_1440);
or U739 (N_739,In_447,N_182);
xor U740 (N_740,N_405,N_240);
nor U741 (N_741,In_1194,In_609);
and U742 (N_742,N_178,In_972);
xor U743 (N_743,In_522,In_635);
and U744 (N_744,In_270,N_384);
or U745 (N_745,In_648,In_543);
and U746 (N_746,In_1361,N_418);
xor U747 (N_747,In_928,In_1337);
nor U748 (N_748,In_1251,N_54);
xor U749 (N_749,N_122,N_309);
and U750 (N_750,N_660,In_59);
nand U751 (N_751,In_1197,N_559);
or U752 (N_752,N_628,N_680);
and U753 (N_753,In_1012,N_202);
xnor U754 (N_754,N_746,N_533);
xnor U755 (N_755,N_544,In_292);
xnor U756 (N_756,N_609,In_336);
or U757 (N_757,N_486,N_677);
xnor U758 (N_758,In_309,N_721);
or U759 (N_759,In_1175,N_255);
nor U760 (N_760,In_582,In_910);
and U761 (N_761,N_7,N_282);
xor U762 (N_762,In_513,N_682);
nor U763 (N_763,N_644,N_49);
or U764 (N_764,In_1128,N_491);
nor U765 (N_765,N_570,N_358);
or U766 (N_766,N_74,In_132);
nor U767 (N_767,In_432,In_854);
and U768 (N_768,In_677,N_556);
nor U769 (N_769,In_342,In_1123);
and U770 (N_770,In_811,In_19);
and U771 (N_771,N_512,In_1241);
or U772 (N_772,N_253,N_641);
or U773 (N_773,N_101,N_704);
or U774 (N_774,N_15,In_1134);
or U775 (N_775,In_903,N_114);
or U776 (N_776,In_356,In_242);
and U777 (N_777,In_1473,In_454);
or U778 (N_778,In_412,In_765);
nor U779 (N_779,N_688,N_717);
or U780 (N_780,N_710,N_382);
xor U781 (N_781,In_772,N_436);
xnor U782 (N_782,N_701,In_205);
nand U783 (N_783,N_545,N_537);
nor U784 (N_784,N_48,In_142);
and U785 (N_785,In_733,In_107);
nand U786 (N_786,N_33,In_1055);
xor U787 (N_787,In_1131,N_689);
xor U788 (N_788,In_481,In_1494);
or U789 (N_789,N_490,N_634);
nor U790 (N_790,N_521,N_340);
nor U791 (N_791,In_562,In_251);
and U792 (N_792,In_428,In_786);
nand U793 (N_793,N_508,N_279);
or U794 (N_794,N_708,N_700);
and U795 (N_795,N_621,In_1287);
xnor U796 (N_796,In_117,In_319);
xnor U797 (N_797,In_1398,N_707);
nand U798 (N_798,N_552,In_995);
nor U799 (N_799,In_199,N_85);
and U800 (N_800,In_215,N_602);
nand U801 (N_801,In_850,In_334);
nor U802 (N_802,In_592,N_243);
and U803 (N_803,In_1010,In_1476);
nor U804 (N_804,N_153,N_543);
or U805 (N_805,N_83,In_993);
nand U806 (N_806,In_705,In_930);
or U807 (N_807,N_157,N_517);
and U808 (N_808,N_633,N_507);
xor U809 (N_809,N_17,In_544);
and U810 (N_810,In_798,N_654);
nor U811 (N_811,N_600,In_978);
and U812 (N_812,In_306,N_611);
or U813 (N_813,N_319,N_541);
and U814 (N_814,N_534,In_324);
nor U815 (N_815,In_404,N_326);
nor U816 (N_816,N_215,N_65);
and U817 (N_817,In_1405,N_561);
and U818 (N_818,N_659,In_114);
xor U819 (N_819,N_740,N_749);
nor U820 (N_820,In_1364,N_442);
and U821 (N_821,In_50,In_900);
nor U822 (N_822,In_1102,In_254);
xor U823 (N_823,N_684,N_290);
nor U824 (N_824,N_276,In_561);
xnor U825 (N_825,N_592,In_916);
and U826 (N_826,N_741,In_629);
xnor U827 (N_827,N_665,N_527);
xnor U828 (N_828,In_1216,N_566);
nand U829 (N_829,N_629,N_70);
xnor U830 (N_830,N_154,N_612);
nand U831 (N_831,In_43,N_50);
and U832 (N_832,N_737,In_869);
and U833 (N_833,N_272,N_350);
nand U834 (N_834,In_865,In_824);
xor U835 (N_835,N_123,In_165);
and U836 (N_836,N_697,N_504);
xor U837 (N_837,N_167,In_260);
xnor U838 (N_838,N_61,N_529);
xnor U839 (N_839,N_658,In_1137);
nand U840 (N_840,N_588,In_1109);
nor U841 (N_841,N_525,In_620);
xor U842 (N_842,N_729,N_635);
nand U843 (N_843,N_551,N_373);
and U844 (N_844,N_192,N_668);
or U845 (N_845,N_648,In_1129);
nand U846 (N_846,N_594,N_331);
xor U847 (N_847,N_361,N_696);
and U848 (N_848,N_509,N_406);
or U849 (N_849,In_1446,N_702);
or U850 (N_850,N_395,N_724);
nand U851 (N_851,N_346,N_497);
nand U852 (N_852,N_580,N_747);
xor U853 (N_853,In_549,N_607);
nor U854 (N_854,In_975,N_636);
nor U855 (N_855,N_348,N_649);
and U856 (N_856,N_314,N_671);
and U857 (N_857,In_1208,N_345);
nand U858 (N_858,N_625,N_550);
xor U859 (N_859,In_1286,N_261);
or U860 (N_860,N_347,N_732);
nor U861 (N_861,In_579,N_328);
and U862 (N_862,In_779,N_603);
nor U863 (N_863,In_392,N_522);
and U864 (N_864,N_410,N_591);
and U865 (N_865,In_262,In_1467);
or U866 (N_866,N_419,In_694);
or U867 (N_867,N_267,In_1227);
and U868 (N_868,N_441,N_246);
nor U869 (N_869,In_348,N_627);
nor U870 (N_870,N_170,N_568);
nor U871 (N_871,In_1438,In_1478);
xor U872 (N_872,N_195,In_1140);
or U873 (N_873,N_631,N_630);
and U874 (N_874,N_598,In_1213);
and U875 (N_875,In_839,N_655);
and U876 (N_876,N_0,In_788);
nand U877 (N_877,N_703,N_500);
nor U878 (N_878,N_428,N_638);
or U879 (N_879,N_397,In_1093);
nor U880 (N_880,N_695,N_359);
nor U881 (N_881,N_672,N_344);
and U882 (N_882,N_584,N_194);
nor U883 (N_883,In_383,N_620);
nand U884 (N_884,N_407,In_430);
or U885 (N_885,In_298,N_542);
nand U886 (N_886,N_515,In_1460);
xor U887 (N_887,N_535,N_505);
xnor U888 (N_888,In_232,In_374);
xnor U889 (N_889,N_652,N_311);
nor U890 (N_890,N_565,N_647);
xor U891 (N_891,N_342,In_892);
nand U892 (N_892,In_77,In_777);
and U893 (N_893,N_694,N_259);
nor U894 (N_894,N_581,In_1434);
xor U895 (N_895,N_706,In_948);
nand U896 (N_896,N_511,N_576);
nor U897 (N_897,N_569,N_368);
or U898 (N_898,N_546,N_663);
or U899 (N_899,In_720,In_376);
nor U900 (N_900,N_151,N_468);
or U901 (N_901,N_610,N_73);
and U902 (N_902,In_647,N_173);
xnor U903 (N_903,In_641,N_593);
nand U904 (N_904,N_254,In_1367);
xnor U905 (N_905,N_563,In_1127);
nor U906 (N_906,N_108,N_720);
or U907 (N_907,In_1458,N_624);
nor U908 (N_908,N_66,N_590);
xor U909 (N_909,In_1419,N_308);
nor U910 (N_910,N_531,N_616);
nand U911 (N_911,N_667,N_530);
nor U912 (N_912,N_613,In_1088);
xor U913 (N_913,N_646,N_455);
xnor U914 (N_914,In_1328,N_396);
nand U915 (N_915,N_748,In_1415);
nor U916 (N_916,N_567,N_69);
and U917 (N_917,N_510,In_976);
xnor U918 (N_918,In_884,N_475);
and U919 (N_919,In_1041,In_13);
xor U920 (N_920,In_101,N_472);
or U921 (N_921,N_232,In_603);
and U922 (N_922,In_593,In_715);
nand U923 (N_923,In_820,N_653);
and U924 (N_924,N_540,N_719);
or U925 (N_925,N_236,N_95);
nand U926 (N_926,In_291,N_622);
xor U927 (N_927,N_499,N_709);
and U928 (N_928,N_632,N_351);
and U929 (N_929,In_578,N_273);
and U930 (N_930,N_131,In_118);
nor U931 (N_931,In_793,In_1172);
xnor U932 (N_932,In_1437,In_1091);
nand U933 (N_933,In_252,In_776);
nand U934 (N_934,N_586,N_303);
or U935 (N_935,In_721,N_736);
nor U936 (N_936,N_560,N_408);
xnor U937 (N_937,N_601,N_725);
or U938 (N_938,N_365,In_1015);
or U939 (N_939,N_413,N_145);
xor U940 (N_940,N_211,N_742);
xnor U941 (N_941,N_16,N_433);
or U942 (N_942,N_657,In_338);
xor U943 (N_943,In_461,N_213);
nor U944 (N_944,In_1176,N_317);
nand U945 (N_945,In_710,In_1231);
nor U946 (N_946,In_437,In_627);
nor U947 (N_947,N_241,N_63);
nor U948 (N_948,N_666,N_723);
and U949 (N_949,N_523,In_346);
nand U950 (N_950,In_180,In_573);
and U951 (N_951,In_445,In_837);
nand U952 (N_952,N_82,N_564);
and U953 (N_953,N_285,N_479);
xor U954 (N_954,In_207,In_413);
nand U955 (N_955,In_536,In_1105);
or U956 (N_956,N_133,N_575);
nand U957 (N_957,N_608,In_54);
xor U958 (N_958,In_1161,N_13);
nor U959 (N_959,N_685,In_1269);
nand U960 (N_960,N_160,N_20);
nor U961 (N_961,N_731,N_733);
xnor U962 (N_962,In_899,In_646);
nor U963 (N_963,In_115,N_639);
and U964 (N_964,N_260,N_577);
nand U965 (N_965,In_433,N_692);
and U966 (N_966,N_127,N_519);
nand U967 (N_967,N_299,N_283);
nand U968 (N_968,N_489,N_43);
nand U969 (N_969,In_1299,In_831);
nand U970 (N_970,In_849,N_378);
nand U971 (N_971,In_36,In_943);
nand U972 (N_972,N_390,N_445);
nor U973 (N_973,In_1324,In_1492);
or U974 (N_974,In_1149,N_113);
and U975 (N_975,N_571,N_589);
and U976 (N_976,N_643,In_867);
and U977 (N_977,N_409,N_619);
nand U978 (N_978,N_650,In_63);
nor U979 (N_979,N_387,In_554);
or U980 (N_980,In_872,N_690);
xor U981 (N_981,In_524,N_558);
nand U982 (N_982,In_722,N_457);
xor U983 (N_983,N_516,N_679);
xnor U984 (N_984,N_180,N_375);
nand U985 (N_985,N_349,In_253);
xnor U986 (N_986,In_206,In_958);
or U987 (N_987,In_563,N_403);
xor U988 (N_988,N_343,In_155);
and U989 (N_989,N_318,N_357);
nor U990 (N_990,N_322,N_675);
and U991 (N_991,N_424,In_161);
nor U992 (N_992,In_949,N_728);
nand U993 (N_993,N_474,N_464);
nand U994 (N_994,N_453,N_712);
xnor U995 (N_995,N_693,N_496);
and U996 (N_996,N_539,N_278);
nand U997 (N_997,N_528,In_1267);
xnor U998 (N_998,N_470,In_974);
or U999 (N_999,N_75,In_1211);
and U1000 (N_1000,N_945,N_866);
nand U1001 (N_1001,In_92,N_758);
nand U1002 (N_1002,N_763,In_1177);
and U1003 (N_1003,N_961,N_975);
nor U1004 (N_1004,In_532,N_783);
nand U1005 (N_1005,N_642,N_949);
nor U1006 (N_1006,N_756,N_868);
and U1007 (N_1007,N_51,N_687);
or U1008 (N_1008,N_734,N_353);
and U1009 (N_1009,N_451,In_1037);
nor U1010 (N_1010,N_711,N_447);
nor U1011 (N_1011,N_876,N_804);
nand U1012 (N_1012,N_810,N_548);
or U1013 (N_1013,N_214,In_451);
nand U1014 (N_1014,N_958,N_903);
and U1015 (N_1015,N_969,N_583);
nand U1016 (N_1016,N_503,In_1158);
nor U1017 (N_1017,N_579,In_724);
or U1018 (N_1018,N_963,N_770);
xnor U1019 (N_1019,N_982,In_136);
nor U1020 (N_1020,N_366,N_811);
or U1021 (N_1021,N_858,N_968);
nand U1022 (N_1022,N_714,N_850);
and U1023 (N_1023,In_361,N_587);
and U1024 (N_1024,N_886,N_404);
nor U1025 (N_1025,N_948,In_1394);
xor U1026 (N_1026,N_939,N_954);
and U1027 (N_1027,N_847,N_801);
and U1028 (N_1028,In_996,N_935);
and U1029 (N_1029,N_879,In_942);
xnor U1030 (N_1030,N_865,N_929);
or U1031 (N_1031,N_596,N_109);
and U1032 (N_1032,In_49,N_165);
and U1033 (N_1033,N_893,N_844);
nand U1034 (N_1034,N_873,N_834);
nand U1035 (N_1035,N_841,N_883);
xor U1036 (N_1036,N_744,N_999);
and U1037 (N_1037,N_64,N_585);
xor U1038 (N_1038,N_518,N_41);
nor U1039 (N_1039,In_918,N_572);
nor U1040 (N_1040,N_200,N_786);
xor U1041 (N_1041,N_787,In_639);
nor U1042 (N_1042,In_539,N_735);
nor U1043 (N_1043,N_798,N_92);
and U1044 (N_1044,N_788,In_990);
or U1045 (N_1045,N_857,In_784);
or U1046 (N_1046,N_926,N_914);
or U1047 (N_1047,In_1365,N_980);
and U1048 (N_1048,N_936,N_824);
or U1049 (N_1049,N_997,N_738);
nand U1050 (N_1050,N_678,N_973);
nor U1051 (N_1051,N_501,In_1344);
or U1052 (N_1052,In_1303,N_524);
nor U1053 (N_1053,In_1191,In_1130);
and U1054 (N_1054,N_400,N_881);
nand U1055 (N_1055,N_899,N_854);
xor U1056 (N_1056,N_894,N_887);
nand U1057 (N_1057,N_916,N_775);
nor U1058 (N_1058,N_901,N_784);
xnor U1059 (N_1059,N_645,N_875);
nor U1060 (N_1060,In_883,In_1117);
and U1061 (N_1061,N_864,N_686);
nor U1062 (N_1062,In_1252,N_771);
nor U1063 (N_1063,N_910,N_983);
nor U1064 (N_1064,N_329,N_88);
nor U1065 (N_1065,N_532,N_991);
xnor U1066 (N_1066,N_888,N_859);
and U1067 (N_1067,N_848,In_1495);
xor U1068 (N_1068,N_913,N_989);
nand U1069 (N_1069,N_843,N_821);
or U1070 (N_1070,N_435,N_411);
nor U1071 (N_1071,N_661,N_891);
nor U1072 (N_1072,N_401,N_861);
nand U1073 (N_1073,N_670,N_752);
or U1074 (N_1074,N_751,N_877);
or U1075 (N_1075,N_870,N_553);
nand U1076 (N_1076,N_753,In_317);
nand U1077 (N_1077,In_349,N_716);
nor U1078 (N_1078,N_933,N_791);
nand U1079 (N_1079,N_898,N_815);
xor U1080 (N_1080,N_909,N_889);
nor U1081 (N_1081,N_768,In_16);
nor U1082 (N_1082,N_994,N_996);
xor U1083 (N_1083,In_525,N_970);
or U1084 (N_1084,N_793,N_872);
and U1085 (N_1085,N_962,N_555);
or U1086 (N_1086,N_767,N_998);
nand U1087 (N_1087,N_265,N_802);
nand U1088 (N_1088,In_964,N_927);
xnor U1089 (N_1089,N_977,In_947);
and U1090 (N_1090,In_150,N_606);
nand U1091 (N_1091,In_893,N_842);
or U1092 (N_1092,N_955,In_1448);
nand U1093 (N_1093,N_176,N_906);
nand U1094 (N_1094,N_895,In_299);
xnor U1095 (N_1095,In_1457,N_10);
xor U1096 (N_1096,N_239,N_754);
and U1097 (N_1097,N_514,N_917);
or U1098 (N_1098,N_513,In_367);
xor U1099 (N_1099,In_723,N_818);
and U1100 (N_1100,N_640,In_57);
nor U1101 (N_1101,In_846,N_807);
nand U1102 (N_1102,N_757,N_800);
nand U1103 (N_1103,In_988,In_268);
nand U1104 (N_1104,N_774,N_855);
xnor U1105 (N_1105,N_837,N_912);
nand U1106 (N_1106,N_617,N_880);
or U1107 (N_1107,In_857,N_871);
nand U1108 (N_1108,N_952,N_907);
and U1109 (N_1109,N_799,N_825);
nor U1110 (N_1110,N_874,N_722);
nor U1111 (N_1111,N_930,N_582);
xnor U1112 (N_1112,N_779,In_416);
and U1113 (N_1113,N_316,In_1260);
or U1114 (N_1114,N_549,N_829);
nand U1115 (N_1115,In_783,In_31);
nor U1116 (N_1116,N_148,N_794);
xor U1117 (N_1117,N_946,N_713);
nand U1118 (N_1118,In_256,In_874);
and U1119 (N_1119,N_772,N_626);
xnor U1120 (N_1120,N_940,N_942);
xor U1121 (N_1121,N_911,In_1179);
or U1122 (N_1122,N_778,N_305);
or U1123 (N_1123,N_944,N_673);
nand U1124 (N_1124,N_538,N_905);
and U1125 (N_1125,N_398,N_773);
xnor U1126 (N_1126,N_446,N_931);
xnor U1127 (N_1127,N_915,In_1205);
nor U1128 (N_1128,N_324,N_536);
and U1129 (N_1129,N_920,N_55);
and U1130 (N_1130,N_974,In_1276);
nor U1131 (N_1131,N_683,N_806);
nor U1132 (N_1132,N_727,N_520);
nor U1133 (N_1133,N_573,In_76);
or U1134 (N_1134,In_222,N_484);
and U1135 (N_1135,N_599,N_789);
nor U1136 (N_1136,N_698,N_923);
nand U1137 (N_1137,N_270,N_781);
and U1138 (N_1138,N_578,N_730);
xnor U1139 (N_1139,N_25,N_803);
nor U1140 (N_1140,N_953,In_297);
xnor U1141 (N_1141,N_277,N_1);
and U1142 (N_1142,In_1336,N_981);
xor U1143 (N_1143,N_597,In_1059);
nor U1144 (N_1144,N_149,N_482);
or U1145 (N_1145,N_743,In_584);
or U1146 (N_1146,N_995,N_805);
nor U1147 (N_1147,N_681,N_820);
xor U1148 (N_1148,N_605,N_937);
or U1149 (N_1149,N_840,In_269);
xnor U1150 (N_1150,In_595,N_892);
or U1151 (N_1151,N_4,In_1027);
nor U1152 (N_1152,N_745,N_144);
nor U1153 (N_1153,N_224,N_823);
xnor U1154 (N_1154,N_813,N_574);
xor U1155 (N_1155,N_988,In_377);
xnor U1156 (N_1156,N_762,N_941);
or U1157 (N_1157,In_552,In_829);
or U1158 (N_1158,N_928,N_623);
and U1159 (N_1159,In_1346,N_934);
and U1160 (N_1160,N_782,N_785);
nand U1161 (N_1161,N_902,N_809);
nor U1162 (N_1162,N_819,N_651);
nand U1163 (N_1163,N_434,N_795);
or U1164 (N_1164,In_1342,N_502);
nand U1165 (N_1165,N_669,In_1028);
and U1166 (N_1166,N_554,N_932);
and U1167 (N_1167,N_780,In_1443);
xor U1168 (N_1168,N_856,N_863);
or U1169 (N_1169,N_766,N_426);
or U1170 (N_1170,N_897,In_489);
xor U1171 (N_1171,N_614,N_900);
nand U1172 (N_1172,N_978,N_792);
xor U1173 (N_1173,N_705,N_89);
or U1174 (N_1174,N_72,N_826);
nand U1175 (N_1175,N_828,N_338);
xnor U1176 (N_1176,N_674,N_78);
and U1177 (N_1177,N_845,N_943);
and U1178 (N_1178,N_830,In_1470);
and U1179 (N_1179,N_919,In_108);
or U1180 (N_1180,In_259,In_1106);
and U1181 (N_1181,N_835,N_676);
nor U1182 (N_1182,N_908,N_812);
nor U1183 (N_1183,N_853,In_1366);
xor U1184 (N_1184,N_699,N_967);
or U1185 (N_1185,N_808,N_816);
and U1186 (N_1186,N_833,In_963);
or U1187 (N_1187,N_849,N_979);
nand U1188 (N_1188,N_852,N_890);
nand U1189 (N_1189,N_862,N_951);
and U1190 (N_1190,N_976,N_761);
xnor U1191 (N_1191,N_960,N_526);
xnor U1192 (N_1192,N_604,N_777);
nor U1193 (N_1193,In_158,N_838);
nor U1194 (N_1194,In_407,N_885);
and U1195 (N_1195,N_832,N_922);
and U1196 (N_1196,N_993,N_769);
or U1197 (N_1197,N_797,N_718);
nand U1198 (N_1198,N_921,N_985);
nand U1199 (N_1199,N_959,In_986);
nand U1200 (N_1200,In_744,N_297);
and U1201 (N_1201,N_776,N_562);
and U1202 (N_1202,N_287,N_992);
nand U1203 (N_1203,N_461,In_1338);
xnor U1204 (N_1204,In_400,N_971);
and U1205 (N_1205,N_966,N_339);
and U1206 (N_1206,N_755,In_243);
and U1207 (N_1207,N_656,In_1014);
or U1208 (N_1208,N_938,N_965);
or U1209 (N_1209,N_814,N_884);
xor U1210 (N_1210,N_370,N_595);
xor U1211 (N_1211,N_765,N_925);
nor U1212 (N_1212,In_90,N_759);
nor U1213 (N_1213,N_904,N_764);
nand U1214 (N_1214,N_924,In_814);
or U1215 (N_1215,N_956,N_990);
nand U1216 (N_1216,N_715,N_427);
or U1217 (N_1217,N_557,In_1301);
nand U1218 (N_1218,In_1214,N_739);
nor U1219 (N_1219,N_790,N_947);
xnor U1220 (N_1220,In_934,N_987);
or U1221 (N_1221,N_851,N_846);
and U1222 (N_1222,N_827,N_860);
nor U1223 (N_1223,N_618,In_1112);
or U1224 (N_1224,N_295,N_972);
and U1225 (N_1225,In_929,In_825);
nand U1226 (N_1226,N_918,N_817);
or U1227 (N_1227,N_878,In_53);
nand U1228 (N_1228,In_1086,In_1486);
nor U1229 (N_1229,N_839,N_402);
nand U1230 (N_1230,N_836,N_483);
nor U1231 (N_1231,N_691,N_822);
or U1232 (N_1232,In_717,In_355);
xnor U1233 (N_1233,N_506,In_1031);
nand U1234 (N_1234,In_1371,N_950);
and U1235 (N_1235,In_176,In_7);
nor U1236 (N_1236,N_984,N_219);
and U1237 (N_1237,N_726,In_10);
xor U1238 (N_1238,N_986,In_123);
or U1239 (N_1239,N_957,N_547);
nand U1240 (N_1240,In_384,N_250);
or U1241 (N_1241,N_896,In_1144);
nor U1242 (N_1242,N_637,N_664);
or U1243 (N_1243,N_869,N_760);
xor U1244 (N_1244,In_1209,N_662);
nand U1245 (N_1245,N_964,In_914);
xor U1246 (N_1246,N_831,N_227);
nand U1247 (N_1247,N_796,In_1164);
nand U1248 (N_1248,N_615,N_867);
nand U1249 (N_1249,N_750,N_882);
xnor U1250 (N_1250,N_1114,N_1127);
or U1251 (N_1251,N_1027,N_1034);
xnor U1252 (N_1252,N_1020,N_1026);
xnor U1253 (N_1253,N_1003,N_1172);
nor U1254 (N_1254,N_1204,N_1092);
xnor U1255 (N_1255,N_1017,N_1080);
nor U1256 (N_1256,N_1016,N_1103);
nor U1257 (N_1257,N_1078,N_1203);
nor U1258 (N_1258,N_1219,N_1234);
nand U1259 (N_1259,N_1097,N_1148);
and U1260 (N_1260,N_1106,N_1056);
xnor U1261 (N_1261,N_1049,N_1185);
xnor U1262 (N_1262,N_1140,N_1066);
xnor U1263 (N_1263,N_1210,N_1079);
xnor U1264 (N_1264,N_1058,N_1096);
xor U1265 (N_1265,N_1012,N_1116);
and U1266 (N_1266,N_1032,N_1180);
xnor U1267 (N_1267,N_1142,N_1134);
xor U1268 (N_1268,N_1044,N_1088);
nor U1269 (N_1269,N_1111,N_1248);
or U1270 (N_1270,N_1177,N_1006);
and U1271 (N_1271,N_1075,N_1192);
or U1272 (N_1272,N_1153,N_1060);
nor U1273 (N_1273,N_1184,N_1035);
and U1274 (N_1274,N_1039,N_1231);
xnor U1275 (N_1275,N_1178,N_1091);
or U1276 (N_1276,N_1194,N_1214);
and U1277 (N_1277,N_1155,N_1045);
or U1278 (N_1278,N_1233,N_1014);
or U1279 (N_1279,N_1159,N_1182);
or U1280 (N_1280,N_1181,N_1024);
nor U1281 (N_1281,N_1196,N_1239);
xor U1282 (N_1282,N_1071,N_1110);
nand U1283 (N_1283,N_1098,N_1128);
and U1284 (N_1284,N_1171,N_1113);
and U1285 (N_1285,N_1226,N_1124);
nand U1286 (N_1286,N_1095,N_1161);
or U1287 (N_1287,N_1123,N_1150);
nor U1288 (N_1288,N_1051,N_1023);
xnor U1289 (N_1289,N_1208,N_1074);
nor U1290 (N_1290,N_1048,N_1218);
and U1291 (N_1291,N_1236,N_1120);
nor U1292 (N_1292,N_1223,N_1033);
and U1293 (N_1293,N_1072,N_1089);
nand U1294 (N_1294,N_1037,N_1149);
or U1295 (N_1295,N_1126,N_1130);
xnor U1296 (N_1296,N_1129,N_1015);
xor U1297 (N_1297,N_1087,N_1093);
or U1298 (N_1298,N_1073,N_1001);
nor U1299 (N_1299,N_1013,N_1019);
xor U1300 (N_1300,N_1036,N_1238);
and U1301 (N_1301,N_1246,N_1167);
or U1302 (N_1302,N_1175,N_1002);
or U1303 (N_1303,N_1068,N_1112);
or U1304 (N_1304,N_1216,N_1188);
nand U1305 (N_1305,N_1232,N_1055);
or U1306 (N_1306,N_1086,N_1152);
nand U1307 (N_1307,N_1160,N_1147);
nor U1308 (N_1308,N_1105,N_1243);
and U1309 (N_1309,N_1011,N_1115);
or U1310 (N_1310,N_1122,N_1157);
xnor U1311 (N_1311,N_1146,N_1198);
xnor U1312 (N_1312,N_1010,N_1108);
or U1313 (N_1313,N_1240,N_1067);
xor U1314 (N_1314,N_1061,N_1237);
nand U1315 (N_1315,N_1212,N_1162);
and U1316 (N_1316,N_1195,N_1005);
or U1317 (N_1317,N_1050,N_1144);
or U1318 (N_1318,N_1085,N_1121);
nand U1319 (N_1319,N_1117,N_1007);
or U1320 (N_1320,N_1028,N_1099);
and U1321 (N_1321,N_1158,N_1165);
or U1322 (N_1322,N_1077,N_1000);
xor U1323 (N_1323,N_1009,N_1118);
or U1324 (N_1324,N_1168,N_1052);
nand U1325 (N_1325,N_1164,N_1100);
or U1326 (N_1326,N_1220,N_1174);
or U1327 (N_1327,N_1043,N_1163);
xnor U1328 (N_1328,N_1202,N_1135);
or U1329 (N_1329,N_1054,N_1018);
nand U1330 (N_1330,N_1047,N_1156);
nand U1331 (N_1331,N_1200,N_1053);
xor U1332 (N_1332,N_1057,N_1038);
nand U1333 (N_1333,N_1247,N_1063);
nor U1334 (N_1334,N_1119,N_1143);
or U1335 (N_1335,N_1042,N_1021);
and U1336 (N_1336,N_1094,N_1211);
and U1337 (N_1337,N_1109,N_1221);
and U1338 (N_1338,N_1083,N_1084);
and U1339 (N_1339,N_1030,N_1076);
nand U1340 (N_1340,N_1101,N_1145);
and U1341 (N_1341,N_1125,N_1081);
or U1342 (N_1342,N_1065,N_1070);
or U1343 (N_1343,N_1173,N_1169);
nand U1344 (N_1344,N_1245,N_1069);
and U1345 (N_1345,N_1138,N_1205);
or U1346 (N_1346,N_1229,N_1059);
or U1347 (N_1347,N_1131,N_1206);
and U1348 (N_1348,N_1242,N_1197);
nor U1349 (N_1349,N_1022,N_1107);
and U1350 (N_1350,N_1199,N_1190);
nor U1351 (N_1351,N_1241,N_1191);
xor U1352 (N_1352,N_1249,N_1228);
or U1353 (N_1353,N_1217,N_1179);
nor U1354 (N_1354,N_1176,N_1064);
nor U1355 (N_1355,N_1230,N_1170);
or U1356 (N_1356,N_1166,N_1004);
nand U1357 (N_1357,N_1029,N_1193);
xor U1358 (N_1358,N_1235,N_1224);
and U1359 (N_1359,N_1141,N_1222);
nand U1360 (N_1360,N_1186,N_1046);
or U1361 (N_1361,N_1207,N_1213);
and U1362 (N_1362,N_1041,N_1102);
nand U1363 (N_1363,N_1183,N_1201);
or U1364 (N_1364,N_1104,N_1154);
nor U1365 (N_1365,N_1031,N_1209);
nand U1366 (N_1366,N_1137,N_1139);
or U1367 (N_1367,N_1244,N_1008);
or U1368 (N_1368,N_1215,N_1090);
and U1369 (N_1369,N_1133,N_1132);
nand U1370 (N_1370,N_1187,N_1062);
or U1371 (N_1371,N_1040,N_1227);
or U1372 (N_1372,N_1225,N_1189);
xor U1373 (N_1373,N_1025,N_1151);
or U1374 (N_1374,N_1136,N_1082);
and U1375 (N_1375,N_1199,N_1104);
nor U1376 (N_1376,N_1032,N_1220);
or U1377 (N_1377,N_1042,N_1074);
or U1378 (N_1378,N_1076,N_1174);
xor U1379 (N_1379,N_1047,N_1171);
xor U1380 (N_1380,N_1078,N_1147);
xor U1381 (N_1381,N_1035,N_1057);
or U1382 (N_1382,N_1078,N_1169);
and U1383 (N_1383,N_1182,N_1143);
nand U1384 (N_1384,N_1186,N_1021);
xnor U1385 (N_1385,N_1161,N_1149);
and U1386 (N_1386,N_1243,N_1171);
nand U1387 (N_1387,N_1024,N_1012);
nand U1388 (N_1388,N_1205,N_1189);
and U1389 (N_1389,N_1174,N_1113);
nand U1390 (N_1390,N_1002,N_1113);
or U1391 (N_1391,N_1143,N_1023);
or U1392 (N_1392,N_1196,N_1034);
nand U1393 (N_1393,N_1241,N_1215);
xnor U1394 (N_1394,N_1149,N_1114);
nor U1395 (N_1395,N_1070,N_1043);
and U1396 (N_1396,N_1179,N_1066);
and U1397 (N_1397,N_1145,N_1218);
nand U1398 (N_1398,N_1150,N_1082);
or U1399 (N_1399,N_1100,N_1231);
xnor U1400 (N_1400,N_1034,N_1016);
xor U1401 (N_1401,N_1145,N_1219);
or U1402 (N_1402,N_1076,N_1190);
nor U1403 (N_1403,N_1221,N_1211);
nand U1404 (N_1404,N_1062,N_1206);
and U1405 (N_1405,N_1168,N_1003);
and U1406 (N_1406,N_1135,N_1139);
or U1407 (N_1407,N_1191,N_1155);
nor U1408 (N_1408,N_1093,N_1106);
nor U1409 (N_1409,N_1173,N_1045);
and U1410 (N_1410,N_1110,N_1243);
nor U1411 (N_1411,N_1011,N_1128);
xnor U1412 (N_1412,N_1059,N_1206);
xnor U1413 (N_1413,N_1003,N_1061);
nor U1414 (N_1414,N_1164,N_1066);
xnor U1415 (N_1415,N_1075,N_1016);
or U1416 (N_1416,N_1136,N_1099);
nand U1417 (N_1417,N_1069,N_1088);
nand U1418 (N_1418,N_1238,N_1035);
nor U1419 (N_1419,N_1048,N_1032);
or U1420 (N_1420,N_1165,N_1164);
xor U1421 (N_1421,N_1080,N_1024);
nand U1422 (N_1422,N_1071,N_1076);
nor U1423 (N_1423,N_1216,N_1012);
or U1424 (N_1424,N_1068,N_1054);
or U1425 (N_1425,N_1038,N_1005);
xor U1426 (N_1426,N_1249,N_1031);
xor U1427 (N_1427,N_1140,N_1131);
or U1428 (N_1428,N_1071,N_1227);
nand U1429 (N_1429,N_1107,N_1049);
nand U1430 (N_1430,N_1172,N_1182);
nor U1431 (N_1431,N_1112,N_1034);
nor U1432 (N_1432,N_1179,N_1060);
nand U1433 (N_1433,N_1198,N_1057);
or U1434 (N_1434,N_1191,N_1224);
xnor U1435 (N_1435,N_1246,N_1109);
or U1436 (N_1436,N_1205,N_1022);
or U1437 (N_1437,N_1071,N_1121);
or U1438 (N_1438,N_1102,N_1094);
nor U1439 (N_1439,N_1114,N_1187);
or U1440 (N_1440,N_1090,N_1013);
and U1441 (N_1441,N_1064,N_1182);
nor U1442 (N_1442,N_1225,N_1055);
nand U1443 (N_1443,N_1172,N_1079);
nand U1444 (N_1444,N_1115,N_1162);
and U1445 (N_1445,N_1175,N_1132);
nor U1446 (N_1446,N_1033,N_1061);
or U1447 (N_1447,N_1179,N_1127);
xor U1448 (N_1448,N_1049,N_1003);
nor U1449 (N_1449,N_1018,N_1215);
nand U1450 (N_1450,N_1112,N_1031);
nor U1451 (N_1451,N_1185,N_1146);
nand U1452 (N_1452,N_1045,N_1057);
or U1453 (N_1453,N_1109,N_1227);
xor U1454 (N_1454,N_1192,N_1045);
nor U1455 (N_1455,N_1015,N_1085);
xnor U1456 (N_1456,N_1027,N_1081);
nor U1457 (N_1457,N_1023,N_1131);
nand U1458 (N_1458,N_1098,N_1177);
nor U1459 (N_1459,N_1141,N_1126);
or U1460 (N_1460,N_1022,N_1087);
nand U1461 (N_1461,N_1161,N_1236);
or U1462 (N_1462,N_1180,N_1196);
and U1463 (N_1463,N_1138,N_1064);
or U1464 (N_1464,N_1141,N_1022);
nor U1465 (N_1465,N_1181,N_1072);
xor U1466 (N_1466,N_1173,N_1149);
and U1467 (N_1467,N_1208,N_1112);
and U1468 (N_1468,N_1053,N_1249);
nand U1469 (N_1469,N_1236,N_1204);
nand U1470 (N_1470,N_1061,N_1133);
and U1471 (N_1471,N_1213,N_1077);
nor U1472 (N_1472,N_1150,N_1247);
or U1473 (N_1473,N_1099,N_1049);
or U1474 (N_1474,N_1120,N_1179);
nand U1475 (N_1475,N_1243,N_1195);
or U1476 (N_1476,N_1050,N_1248);
nor U1477 (N_1477,N_1087,N_1116);
xnor U1478 (N_1478,N_1181,N_1210);
or U1479 (N_1479,N_1069,N_1057);
nor U1480 (N_1480,N_1162,N_1074);
xnor U1481 (N_1481,N_1180,N_1014);
and U1482 (N_1482,N_1024,N_1172);
nand U1483 (N_1483,N_1028,N_1089);
or U1484 (N_1484,N_1219,N_1030);
or U1485 (N_1485,N_1000,N_1067);
xnor U1486 (N_1486,N_1103,N_1193);
and U1487 (N_1487,N_1194,N_1080);
or U1488 (N_1488,N_1109,N_1116);
xor U1489 (N_1489,N_1229,N_1205);
and U1490 (N_1490,N_1079,N_1231);
nor U1491 (N_1491,N_1089,N_1003);
and U1492 (N_1492,N_1011,N_1161);
nor U1493 (N_1493,N_1113,N_1234);
and U1494 (N_1494,N_1186,N_1089);
nand U1495 (N_1495,N_1137,N_1052);
xnor U1496 (N_1496,N_1224,N_1039);
nor U1497 (N_1497,N_1173,N_1063);
xnor U1498 (N_1498,N_1046,N_1086);
xor U1499 (N_1499,N_1079,N_1156);
and U1500 (N_1500,N_1496,N_1422);
nor U1501 (N_1501,N_1292,N_1392);
and U1502 (N_1502,N_1449,N_1367);
or U1503 (N_1503,N_1409,N_1260);
nand U1504 (N_1504,N_1405,N_1407);
nand U1505 (N_1505,N_1492,N_1278);
and U1506 (N_1506,N_1438,N_1316);
nor U1507 (N_1507,N_1310,N_1468);
xor U1508 (N_1508,N_1293,N_1432);
nor U1509 (N_1509,N_1300,N_1259);
nor U1510 (N_1510,N_1271,N_1254);
nand U1511 (N_1511,N_1329,N_1305);
nand U1512 (N_1512,N_1301,N_1404);
xor U1513 (N_1513,N_1471,N_1368);
xor U1514 (N_1514,N_1441,N_1378);
nor U1515 (N_1515,N_1261,N_1325);
xnor U1516 (N_1516,N_1448,N_1323);
xor U1517 (N_1517,N_1466,N_1375);
and U1518 (N_1518,N_1332,N_1415);
xor U1519 (N_1519,N_1430,N_1287);
or U1520 (N_1520,N_1490,N_1402);
nor U1521 (N_1521,N_1348,N_1451);
xnor U1522 (N_1522,N_1483,N_1336);
or U1523 (N_1523,N_1250,N_1251);
and U1524 (N_1524,N_1442,N_1253);
xor U1525 (N_1525,N_1341,N_1495);
or U1526 (N_1526,N_1372,N_1414);
or U1527 (N_1527,N_1377,N_1309);
nand U1528 (N_1528,N_1469,N_1347);
and U1529 (N_1529,N_1380,N_1423);
and U1530 (N_1530,N_1411,N_1317);
and U1531 (N_1531,N_1308,N_1333);
xnor U1532 (N_1532,N_1464,N_1339);
xor U1533 (N_1533,N_1327,N_1397);
nor U1534 (N_1534,N_1354,N_1462);
nand U1535 (N_1535,N_1427,N_1344);
nand U1536 (N_1536,N_1296,N_1470);
and U1537 (N_1537,N_1472,N_1491);
nor U1538 (N_1538,N_1330,N_1489);
xnor U1539 (N_1539,N_1290,N_1302);
or U1540 (N_1540,N_1376,N_1312);
nor U1541 (N_1541,N_1303,N_1281);
xor U1542 (N_1542,N_1418,N_1360);
nor U1543 (N_1543,N_1479,N_1369);
or U1544 (N_1544,N_1364,N_1444);
or U1545 (N_1545,N_1357,N_1399);
nor U1546 (N_1546,N_1428,N_1382);
or U1547 (N_1547,N_1389,N_1443);
and U1548 (N_1548,N_1497,N_1484);
nand U1549 (N_1549,N_1450,N_1306);
nand U1550 (N_1550,N_1390,N_1349);
and U1551 (N_1551,N_1431,N_1416);
nand U1552 (N_1552,N_1454,N_1280);
and U1553 (N_1553,N_1365,N_1421);
or U1554 (N_1554,N_1467,N_1353);
or U1555 (N_1555,N_1340,N_1412);
or U1556 (N_1556,N_1352,N_1342);
nand U1557 (N_1557,N_1391,N_1337);
nand U1558 (N_1558,N_1363,N_1410);
and U1559 (N_1559,N_1335,N_1298);
or U1560 (N_1560,N_1493,N_1475);
and U1561 (N_1561,N_1326,N_1328);
and U1562 (N_1562,N_1463,N_1277);
or U1563 (N_1563,N_1371,N_1446);
xnor U1564 (N_1564,N_1366,N_1485);
nand U1565 (N_1565,N_1417,N_1388);
or U1566 (N_1566,N_1264,N_1374);
and U1567 (N_1567,N_1276,N_1262);
and U1568 (N_1568,N_1439,N_1482);
or U1569 (N_1569,N_1370,N_1481);
nand U1570 (N_1570,N_1447,N_1361);
nand U1571 (N_1571,N_1252,N_1313);
xnor U1572 (N_1572,N_1355,N_1486);
and U1573 (N_1573,N_1295,N_1265);
nor U1574 (N_1574,N_1478,N_1358);
nand U1575 (N_1575,N_1291,N_1393);
or U1576 (N_1576,N_1473,N_1315);
nand U1577 (N_1577,N_1429,N_1425);
xor U1578 (N_1578,N_1297,N_1346);
nand U1579 (N_1579,N_1311,N_1474);
nor U1580 (N_1580,N_1272,N_1273);
and U1581 (N_1581,N_1275,N_1322);
nand U1582 (N_1582,N_1387,N_1266);
nor U1583 (N_1583,N_1263,N_1288);
xor U1584 (N_1584,N_1269,N_1437);
or U1585 (N_1585,N_1362,N_1359);
and U1586 (N_1586,N_1279,N_1384);
or U1587 (N_1587,N_1381,N_1258);
and U1588 (N_1588,N_1461,N_1268);
or U1589 (N_1589,N_1319,N_1396);
nor U1590 (N_1590,N_1408,N_1480);
nor U1591 (N_1591,N_1379,N_1320);
nor U1592 (N_1592,N_1285,N_1350);
nand U1593 (N_1593,N_1334,N_1274);
nand U1594 (N_1594,N_1465,N_1385);
or U1595 (N_1595,N_1499,N_1459);
and U1596 (N_1596,N_1304,N_1406);
and U1597 (N_1597,N_1282,N_1324);
nand U1598 (N_1598,N_1420,N_1488);
nor U1599 (N_1599,N_1283,N_1395);
or U1600 (N_1600,N_1256,N_1476);
xnor U1601 (N_1601,N_1419,N_1458);
nor U1602 (N_1602,N_1403,N_1398);
nor U1603 (N_1603,N_1456,N_1294);
xor U1604 (N_1604,N_1356,N_1257);
or U1605 (N_1605,N_1289,N_1321);
nor U1606 (N_1606,N_1452,N_1351);
or U1607 (N_1607,N_1270,N_1477);
xor U1608 (N_1608,N_1440,N_1426);
or U1609 (N_1609,N_1394,N_1457);
nand U1610 (N_1610,N_1424,N_1445);
or U1611 (N_1611,N_1284,N_1373);
and U1612 (N_1612,N_1338,N_1498);
or U1613 (N_1613,N_1383,N_1331);
or U1614 (N_1614,N_1487,N_1400);
and U1615 (N_1615,N_1435,N_1453);
nor U1616 (N_1616,N_1318,N_1345);
nor U1617 (N_1617,N_1401,N_1255);
and U1618 (N_1618,N_1455,N_1434);
nor U1619 (N_1619,N_1436,N_1386);
or U1620 (N_1620,N_1433,N_1314);
and U1621 (N_1621,N_1286,N_1307);
xnor U1622 (N_1622,N_1460,N_1343);
or U1623 (N_1623,N_1299,N_1413);
and U1624 (N_1624,N_1267,N_1494);
nor U1625 (N_1625,N_1372,N_1315);
or U1626 (N_1626,N_1459,N_1321);
xor U1627 (N_1627,N_1415,N_1420);
nor U1628 (N_1628,N_1318,N_1255);
xor U1629 (N_1629,N_1301,N_1360);
nand U1630 (N_1630,N_1250,N_1366);
or U1631 (N_1631,N_1366,N_1497);
or U1632 (N_1632,N_1252,N_1275);
or U1633 (N_1633,N_1345,N_1264);
nor U1634 (N_1634,N_1322,N_1479);
or U1635 (N_1635,N_1400,N_1371);
and U1636 (N_1636,N_1445,N_1288);
nor U1637 (N_1637,N_1348,N_1452);
nand U1638 (N_1638,N_1467,N_1299);
nor U1639 (N_1639,N_1251,N_1386);
nand U1640 (N_1640,N_1493,N_1426);
xnor U1641 (N_1641,N_1362,N_1253);
nand U1642 (N_1642,N_1417,N_1478);
and U1643 (N_1643,N_1397,N_1282);
and U1644 (N_1644,N_1296,N_1412);
xor U1645 (N_1645,N_1334,N_1359);
and U1646 (N_1646,N_1469,N_1288);
or U1647 (N_1647,N_1299,N_1373);
or U1648 (N_1648,N_1430,N_1252);
or U1649 (N_1649,N_1400,N_1320);
nand U1650 (N_1650,N_1327,N_1370);
nor U1651 (N_1651,N_1358,N_1257);
nand U1652 (N_1652,N_1367,N_1308);
xnor U1653 (N_1653,N_1399,N_1473);
xor U1654 (N_1654,N_1404,N_1442);
and U1655 (N_1655,N_1439,N_1277);
or U1656 (N_1656,N_1257,N_1296);
or U1657 (N_1657,N_1297,N_1415);
nor U1658 (N_1658,N_1276,N_1360);
or U1659 (N_1659,N_1263,N_1459);
nor U1660 (N_1660,N_1490,N_1436);
or U1661 (N_1661,N_1454,N_1255);
xor U1662 (N_1662,N_1283,N_1446);
and U1663 (N_1663,N_1458,N_1349);
nor U1664 (N_1664,N_1411,N_1385);
and U1665 (N_1665,N_1433,N_1305);
or U1666 (N_1666,N_1452,N_1464);
xnor U1667 (N_1667,N_1464,N_1497);
and U1668 (N_1668,N_1384,N_1401);
xnor U1669 (N_1669,N_1499,N_1413);
nor U1670 (N_1670,N_1438,N_1465);
and U1671 (N_1671,N_1459,N_1314);
nand U1672 (N_1672,N_1480,N_1491);
nand U1673 (N_1673,N_1455,N_1287);
xnor U1674 (N_1674,N_1462,N_1314);
xnor U1675 (N_1675,N_1268,N_1280);
nor U1676 (N_1676,N_1413,N_1400);
xor U1677 (N_1677,N_1377,N_1474);
nor U1678 (N_1678,N_1264,N_1406);
nand U1679 (N_1679,N_1487,N_1334);
nand U1680 (N_1680,N_1445,N_1273);
nor U1681 (N_1681,N_1419,N_1341);
and U1682 (N_1682,N_1486,N_1419);
and U1683 (N_1683,N_1488,N_1290);
nand U1684 (N_1684,N_1400,N_1373);
nand U1685 (N_1685,N_1281,N_1300);
xnor U1686 (N_1686,N_1447,N_1491);
or U1687 (N_1687,N_1282,N_1373);
and U1688 (N_1688,N_1496,N_1443);
and U1689 (N_1689,N_1448,N_1316);
and U1690 (N_1690,N_1480,N_1417);
xnor U1691 (N_1691,N_1401,N_1481);
xor U1692 (N_1692,N_1495,N_1374);
and U1693 (N_1693,N_1407,N_1316);
or U1694 (N_1694,N_1332,N_1356);
or U1695 (N_1695,N_1369,N_1432);
nand U1696 (N_1696,N_1257,N_1421);
or U1697 (N_1697,N_1282,N_1496);
nor U1698 (N_1698,N_1298,N_1462);
xor U1699 (N_1699,N_1401,N_1447);
xnor U1700 (N_1700,N_1468,N_1274);
and U1701 (N_1701,N_1465,N_1427);
nand U1702 (N_1702,N_1397,N_1376);
nor U1703 (N_1703,N_1382,N_1402);
and U1704 (N_1704,N_1487,N_1269);
nand U1705 (N_1705,N_1372,N_1361);
and U1706 (N_1706,N_1497,N_1332);
or U1707 (N_1707,N_1252,N_1324);
or U1708 (N_1708,N_1375,N_1331);
or U1709 (N_1709,N_1426,N_1408);
and U1710 (N_1710,N_1369,N_1424);
or U1711 (N_1711,N_1329,N_1448);
xnor U1712 (N_1712,N_1318,N_1498);
and U1713 (N_1713,N_1275,N_1400);
xnor U1714 (N_1714,N_1463,N_1374);
nor U1715 (N_1715,N_1378,N_1274);
or U1716 (N_1716,N_1392,N_1413);
xor U1717 (N_1717,N_1357,N_1425);
xnor U1718 (N_1718,N_1363,N_1372);
nand U1719 (N_1719,N_1297,N_1441);
nand U1720 (N_1720,N_1282,N_1346);
and U1721 (N_1721,N_1270,N_1277);
or U1722 (N_1722,N_1278,N_1285);
nor U1723 (N_1723,N_1424,N_1356);
xnor U1724 (N_1724,N_1366,N_1276);
nor U1725 (N_1725,N_1259,N_1401);
nor U1726 (N_1726,N_1480,N_1306);
nand U1727 (N_1727,N_1430,N_1320);
and U1728 (N_1728,N_1470,N_1361);
and U1729 (N_1729,N_1454,N_1330);
nand U1730 (N_1730,N_1360,N_1272);
and U1731 (N_1731,N_1300,N_1250);
or U1732 (N_1732,N_1360,N_1459);
nor U1733 (N_1733,N_1418,N_1453);
and U1734 (N_1734,N_1396,N_1412);
or U1735 (N_1735,N_1419,N_1353);
or U1736 (N_1736,N_1323,N_1310);
nor U1737 (N_1737,N_1460,N_1332);
or U1738 (N_1738,N_1383,N_1252);
or U1739 (N_1739,N_1309,N_1473);
and U1740 (N_1740,N_1357,N_1314);
xnor U1741 (N_1741,N_1352,N_1479);
or U1742 (N_1742,N_1265,N_1478);
xor U1743 (N_1743,N_1383,N_1419);
nor U1744 (N_1744,N_1406,N_1320);
nor U1745 (N_1745,N_1365,N_1307);
xor U1746 (N_1746,N_1385,N_1350);
xor U1747 (N_1747,N_1264,N_1491);
xnor U1748 (N_1748,N_1391,N_1250);
xor U1749 (N_1749,N_1367,N_1335);
or U1750 (N_1750,N_1563,N_1595);
and U1751 (N_1751,N_1600,N_1502);
nand U1752 (N_1752,N_1527,N_1501);
and U1753 (N_1753,N_1657,N_1588);
xor U1754 (N_1754,N_1567,N_1673);
or U1755 (N_1755,N_1503,N_1571);
and U1756 (N_1756,N_1544,N_1558);
and U1757 (N_1757,N_1662,N_1630);
nor U1758 (N_1758,N_1608,N_1510);
or U1759 (N_1759,N_1664,N_1661);
nor U1760 (N_1760,N_1597,N_1640);
xor U1761 (N_1761,N_1678,N_1607);
nor U1762 (N_1762,N_1705,N_1632);
xor U1763 (N_1763,N_1702,N_1591);
nand U1764 (N_1764,N_1746,N_1715);
nand U1765 (N_1765,N_1530,N_1541);
nor U1766 (N_1766,N_1519,N_1634);
nor U1767 (N_1767,N_1564,N_1668);
nor U1768 (N_1768,N_1689,N_1653);
nand U1769 (N_1769,N_1742,N_1701);
or U1770 (N_1770,N_1672,N_1547);
or U1771 (N_1771,N_1726,N_1655);
nand U1772 (N_1772,N_1658,N_1552);
nand U1773 (N_1773,N_1526,N_1575);
and U1774 (N_1774,N_1584,N_1743);
and U1775 (N_1775,N_1718,N_1551);
or U1776 (N_1776,N_1725,N_1507);
and U1777 (N_1777,N_1561,N_1533);
nor U1778 (N_1778,N_1635,N_1627);
xnor U1779 (N_1779,N_1611,N_1679);
and U1780 (N_1780,N_1631,N_1538);
nand U1781 (N_1781,N_1617,N_1589);
and U1782 (N_1782,N_1566,N_1546);
and U1783 (N_1783,N_1537,N_1572);
nand U1784 (N_1784,N_1529,N_1694);
xnor U1785 (N_1785,N_1670,N_1555);
and U1786 (N_1786,N_1578,N_1711);
nor U1787 (N_1787,N_1626,N_1587);
or U1788 (N_1788,N_1666,N_1615);
xnor U1789 (N_1789,N_1594,N_1706);
nand U1790 (N_1790,N_1623,N_1605);
nand U1791 (N_1791,N_1622,N_1698);
nor U1792 (N_1792,N_1565,N_1690);
and U1793 (N_1793,N_1643,N_1739);
or U1794 (N_1794,N_1727,N_1514);
xnor U1795 (N_1795,N_1610,N_1504);
nor U1796 (N_1796,N_1740,N_1534);
nor U1797 (N_1797,N_1676,N_1722);
nand U1798 (N_1798,N_1683,N_1719);
or U1799 (N_1799,N_1599,N_1557);
nand U1800 (N_1800,N_1545,N_1521);
nor U1801 (N_1801,N_1738,N_1515);
xor U1802 (N_1802,N_1590,N_1654);
and U1803 (N_1803,N_1650,N_1637);
xor U1804 (N_1804,N_1665,N_1684);
xnor U1805 (N_1805,N_1542,N_1708);
xor U1806 (N_1806,N_1570,N_1604);
or U1807 (N_1807,N_1586,N_1735);
nor U1808 (N_1808,N_1724,N_1736);
nor U1809 (N_1809,N_1596,N_1512);
or U1810 (N_1810,N_1749,N_1598);
nand U1811 (N_1811,N_1516,N_1629);
nand U1812 (N_1812,N_1697,N_1687);
nor U1813 (N_1813,N_1688,N_1734);
nand U1814 (N_1814,N_1549,N_1531);
nand U1815 (N_1815,N_1638,N_1651);
xor U1816 (N_1816,N_1569,N_1577);
or U1817 (N_1817,N_1576,N_1535);
and U1818 (N_1818,N_1500,N_1737);
or U1819 (N_1819,N_1613,N_1709);
and U1820 (N_1820,N_1671,N_1693);
and U1821 (N_1821,N_1513,N_1508);
xor U1822 (N_1822,N_1729,N_1660);
nor U1823 (N_1823,N_1717,N_1550);
xnor U1824 (N_1824,N_1744,N_1603);
and U1825 (N_1825,N_1641,N_1568);
or U1826 (N_1826,N_1731,N_1525);
and U1827 (N_1827,N_1573,N_1720);
xor U1828 (N_1828,N_1614,N_1520);
nor U1829 (N_1829,N_1579,N_1644);
nor U1830 (N_1830,N_1663,N_1556);
or U1831 (N_1831,N_1609,N_1618);
nand U1832 (N_1832,N_1728,N_1522);
xor U1833 (N_1833,N_1612,N_1625);
xnor U1834 (N_1834,N_1713,N_1677);
or U1835 (N_1835,N_1621,N_1633);
and U1836 (N_1836,N_1692,N_1730);
nand U1837 (N_1837,N_1646,N_1707);
nor U1838 (N_1838,N_1548,N_1710);
nand U1839 (N_1839,N_1656,N_1592);
and U1840 (N_1840,N_1647,N_1582);
and U1841 (N_1841,N_1649,N_1606);
or U1842 (N_1842,N_1562,N_1703);
xnor U1843 (N_1843,N_1511,N_1523);
and U1844 (N_1844,N_1695,N_1636);
or U1845 (N_1845,N_1583,N_1506);
nor U1846 (N_1846,N_1685,N_1691);
and U1847 (N_1847,N_1574,N_1518);
nand U1848 (N_1848,N_1528,N_1741);
xnor U1849 (N_1849,N_1642,N_1721);
xnor U1850 (N_1850,N_1645,N_1532);
nand U1851 (N_1851,N_1659,N_1560);
nand U1852 (N_1852,N_1601,N_1745);
or U1853 (N_1853,N_1524,N_1675);
or U1854 (N_1854,N_1581,N_1593);
xor U1855 (N_1855,N_1559,N_1536);
or U1856 (N_1856,N_1682,N_1716);
or U1857 (N_1857,N_1509,N_1553);
and U1858 (N_1858,N_1733,N_1748);
nor U1859 (N_1859,N_1540,N_1699);
and U1860 (N_1860,N_1616,N_1674);
xor U1861 (N_1861,N_1619,N_1667);
nand U1862 (N_1862,N_1624,N_1686);
nand U1863 (N_1863,N_1648,N_1585);
nand U1864 (N_1864,N_1554,N_1747);
nor U1865 (N_1865,N_1723,N_1669);
nand U1866 (N_1866,N_1696,N_1620);
and U1867 (N_1867,N_1602,N_1732);
or U1868 (N_1868,N_1639,N_1543);
nand U1869 (N_1869,N_1681,N_1539);
and U1870 (N_1870,N_1628,N_1505);
nor U1871 (N_1871,N_1652,N_1712);
nor U1872 (N_1872,N_1680,N_1517);
nand U1873 (N_1873,N_1580,N_1700);
xnor U1874 (N_1874,N_1704,N_1714);
nand U1875 (N_1875,N_1536,N_1598);
and U1876 (N_1876,N_1726,N_1542);
and U1877 (N_1877,N_1518,N_1517);
or U1878 (N_1878,N_1712,N_1563);
nor U1879 (N_1879,N_1550,N_1586);
and U1880 (N_1880,N_1508,N_1572);
nor U1881 (N_1881,N_1573,N_1664);
xnor U1882 (N_1882,N_1569,N_1609);
nor U1883 (N_1883,N_1595,N_1543);
or U1884 (N_1884,N_1607,N_1504);
nand U1885 (N_1885,N_1650,N_1529);
nor U1886 (N_1886,N_1640,N_1711);
or U1887 (N_1887,N_1564,N_1619);
or U1888 (N_1888,N_1719,N_1745);
or U1889 (N_1889,N_1710,N_1735);
xor U1890 (N_1890,N_1518,N_1546);
xnor U1891 (N_1891,N_1564,N_1685);
or U1892 (N_1892,N_1621,N_1658);
nand U1893 (N_1893,N_1672,N_1646);
or U1894 (N_1894,N_1533,N_1601);
nor U1895 (N_1895,N_1679,N_1609);
or U1896 (N_1896,N_1668,N_1696);
nand U1897 (N_1897,N_1735,N_1597);
and U1898 (N_1898,N_1693,N_1719);
xnor U1899 (N_1899,N_1507,N_1552);
nor U1900 (N_1900,N_1665,N_1610);
and U1901 (N_1901,N_1720,N_1652);
nor U1902 (N_1902,N_1649,N_1733);
or U1903 (N_1903,N_1678,N_1652);
and U1904 (N_1904,N_1649,N_1651);
nor U1905 (N_1905,N_1633,N_1651);
nand U1906 (N_1906,N_1581,N_1594);
or U1907 (N_1907,N_1731,N_1542);
xor U1908 (N_1908,N_1717,N_1674);
xnor U1909 (N_1909,N_1738,N_1593);
nor U1910 (N_1910,N_1665,N_1676);
xor U1911 (N_1911,N_1605,N_1606);
nor U1912 (N_1912,N_1744,N_1532);
or U1913 (N_1913,N_1686,N_1666);
or U1914 (N_1914,N_1549,N_1728);
and U1915 (N_1915,N_1572,N_1575);
or U1916 (N_1916,N_1637,N_1684);
and U1917 (N_1917,N_1746,N_1736);
nand U1918 (N_1918,N_1700,N_1667);
xnor U1919 (N_1919,N_1597,N_1630);
nor U1920 (N_1920,N_1661,N_1625);
nor U1921 (N_1921,N_1592,N_1700);
and U1922 (N_1922,N_1705,N_1550);
nand U1923 (N_1923,N_1731,N_1514);
and U1924 (N_1924,N_1591,N_1589);
xnor U1925 (N_1925,N_1699,N_1643);
nor U1926 (N_1926,N_1544,N_1741);
nor U1927 (N_1927,N_1613,N_1746);
or U1928 (N_1928,N_1549,N_1569);
and U1929 (N_1929,N_1512,N_1682);
nor U1930 (N_1930,N_1712,N_1650);
or U1931 (N_1931,N_1665,N_1615);
xnor U1932 (N_1932,N_1650,N_1681);
and U1933 (N_1933,N_1552,N_1506);
nand U1934 (N_1934,N_1559,N_1708);
nor U1935 (N_1935,N_1568,N_1617);
and U1936 (N_1936,N_1606,N_1661);
nand U1937 (N_1937,N_1732,N_1577);
or U1938 (N_1938,N_1741,N_1641);
and U1939 (N_1939,N_1617,N_1550);
nand U1940 (N_1940,N_1749,N_1713);
and U1941 (N_1941,N_1673,N_1689);
nor U1942 (N_1942,N_1548,N_1615);
nand U1943 (N_1943,N_1569,N_1554);
or U1944 (N_1944,N_1721,N_1682);
or U1945 (N_1945,N_1664,N_1718);
nor U1946 (N_1946,N_1655,N_1537);
nor U1947 (N_1947,N_1610,N_1664);
and U1948 (N_1948,N_1547,N_1723);
or U1949 (N_1949,N_1558,N_1699);
nand U1950 (N_1950,N_1517,N_1614);
nor U1951 (N_1951,N_1658,N_1721);
or U1952 (N_1952,N_1736,N_1737);
or U1953 (N_1953,N_1706,N_1747);
nor U1954 (N_1954,N_1642,N_1595);
and U1955 (N_1955,N_1653,N_1607);
nand U1956 (N_1956,N_1587,N_1685);
and U1957 (N_1957,N_1651,N_1558);
nand U1958 (N_1958,N_1665,N_1711);
nand U1959 (N_1959,N_1563,N_1524);
and U1960 (N_1960,N_1717,N_1608);
nor U1961 (N_1961,N_1613,N_1619);
xor U1962 (N_1962,N_1692,N_1557);
nand U1963 (N_1963,N_1534,N_1664);
or U1964 (N_1964,N_1583,N_1629);
nor U1965 (N_1965,N_1555,N_1710);
xor U1966 (N_1966,N_1732,N_1686);
or U1967 (N_1967,N_1607,N_1627);
and U1968 (N_1968,N_1503,N_1715);
nand U1969 (N_1969,N_1711,N_1504);
xor U1970 (N_1970,N_1604,N_1745);
xor U1971 (N_1971,N_1719,N_1705);
nand U1972 (N_1972,N_1524,N_1599);
xor U1973 (N_1973,N_1601,N_1678);
xnor U1974 (N_1974,N_1512,N_1675);
xnor U1975 (N_1975,N_1714,N_1508);
xnor U1976 (N_1976,N_1718,N_1513);
and U1977 (N_1977,N_1723,N_1607);
nand U1978 (N_1978,N_1743,N_1587);
and U1979 (N_1979,N_1555,N_1546);
nand U1980 (N_1980,N_1588,N_1651);
nor U1981 (N_1981,N_1748,N_1685);
nand U1982 (N_1982,N_1738,N_1532);
nand U1983 (N_1983,N_1600,N_1689);
or U1984 (N_1984,N_1678,N_1563);
and U1985 (N_1985,N_1502,N_1709);
nor U1986 (N_1986,N_1555,N_1595);
nand U1987 (N_1987,N_1653,N_1584);
xnor U1988 (N_1988,N_1748,N_1665);
or U1989 (N_1989,N_1637,N_1577);
nor U1990 (N_1990,N_1745,N_1671);
and U1991 (N_1991,N_1605,N_1593);
or U1992 (N_1992,N_1617,N_1512);
xnor U1993 (N_1993,N_1573,N_1533);
nor U1994 (N_1994,N_1567,N_1556);
xor U1995 (N_1995,N_1629,N_1568);
and U1996 (N_1996,N_1572,N_1591);
nand U1997 (N_1997,N_1552,N_1615);
xor U1998 (N_1998,N_1674,N_1518);
nor U1999 (N_1999,N_1687,N_1525);
or U2000 (N_2000,N_1784,N_1750);
xnor U2001 (N_2001,N_1964,N_1904);
nor U2002 (N_2002,N_1871,N_1893);
or U2003 (N_2003,N_1843,N_1921);
or U2004 (N_2004,N_1866,N_1958);
nor U2005 (N_2005,N_1848,N_1889);
xor U2006 (N_2006,N_1795,N_1790);
xnor U2007 (N_2007,N_1973,N_1791);
and U2008 (N_2008,N_1918,N_1880);
nor U2009 (N_2009,N_1854,N_1929);
nor U2010 (N_2010,N_1870,N_1839);
or U2011 (N_2011,N_1951,N_1978);
nor U2012 (N_2012,N_1912,N_1980);
nand U2013 (N_2013,N_1828,N_1997);
xor U2014 (N_2014,N_1922,N_1859);
and U2015 (N_2015,N_1915,N_1829);
nand U2016 (N_2016,N_1924,N_1770);
nor U2017 (N_2017,N_1761,N_1927);
xor U2018 (N_2018,N_1949,N_1936);
and U2019 (N_2019,N_1930,N_1847);
nor U2020 (N_2020,N_1882,N_1776);
or U2021 (N_2021,N_1967,N_1999);
nand U2022 (N_2022,N_1935,N_1852);
and U2023 (N_2023,N_1794,N_1873);
xor U2024 (N_2024,N_1890,N_1768);
or U2025 (N_2025,N_1966,N_1939);
and U2026 (N_2026,N_1832,N_1931);
xnor U2027 (N_2027,N_1867,N_1875);
nor U2028 (N_2028,N_1817,N_1987);
nor U2029 (N_2029,N_1996,N_1914);
or U2030 (N_2030,N_1830,N_1865);
nand U2031 (N_2031,N_1797,N_1986);
nand U2032 (N_2032,N_1900,N_1759);
or U2033 (N_2033,N_1942,N_1968);
or U2034 (N_2034,N_1983,N_1869);
xnor U2035 (N_2035,N_1975,N_1754);
nand U2036 (N_2036,N_1793,N_1998);
or U2037 (N_2037,N_1823,N_1884);
nor U2038 (N_2038,N_1895,N_1952);
and U2039 (N_2039,N_1800,N_1773);
nand U2040 (N_2040,N_1970,N_1940);
and U2041 (N_2041,N_1891,N_1826);
and U2042 (N_2042,N_1801,N_1860);
xnor U2043 (N_2043,N_1899,N_1818);
and U2044 (N_2044,N_1907,N_1979);
nor U2045 (N_2045,N_1863,N_1888);
xnor U2046 (N_2046,N_1756,N_1934);
nand U2047 (N_2047,N_1835,N_1827);
and U2048 (N_2048,N_1954,N_1864);
or U2049 (N_2049,N_1775,N_1868);
and U2050 (N_2050,N_1969,N_1782);
xnor U2051 (N_2051,N_1906,N_1877);
nor U2052 (N_2052,N_1883,N_1887);
or U2053 (N_2053,N_1971,N_1896);
nor U2054 (N_2054,N_1956,N_1909);
or U2055 (N_2055,N_1816,N_1941);
xor U2056 (N_2056,N_1955,N_1851);
and U2057 (N_2057,N_1789,N_1894);
nand U2058 (N_2058,N_1799,N_1985);
or U2059 (N_2059,N_1858,N_1804);
nand U2060 (N_2060,N_1758,N_1903);
nor U2061 (N_2061,N_1994,N_1802);
nor U2062 (N_2062,N_1774,N_1963);
and U2063 (N_2063,N_1783,N_1910);
or U2064 (N_2064,N_1885,N_1777);
or U2065 (N_2065,N_1812,N_1984);
xor U2066 (N_2066,N_1982,N_1861);
nor U2067 (N_2067,N_1913,N_1992);
nand U2068 (N_2068,N_1932,N_1806);
nor U2069 (N_2069,N_1988,N_1905);
nor U2070 (N_2070,N_1995,N_1840);
and U2071 (N_2071,N_1957,N_1944);
or U2072 (N_2072,N_1943,N_1815);
nor U2073 (N_2073,N_1993,N_1961);
xnor U2074 (N_2074,N_1881,N_1925);
or U2075 (N_2075,N_1965,N_1809);
and U2076 (N_2076,N_1796,N_1845);
xor U2077 (N_2077,N_1926,N_1763);
or U2078 (N_2078,N_1902,N_1853);
nand U2079 (N_2079,N_1779,N_1751);
or U2080 (N_2080,N_1976,N_1923);
nor U2081 (N_2081,N_1803,N_1886);
nor U2082 (N_2082,N_1950,N_1916);
xor U2083 (N_2083,N_1762,N_1959);
and U2084 (N_2084,N_1945,N_1781);
nand U2085 (N_2085,N_1821,N_1990);
nor U2086 (N_2086,N_1849,N_1813);
nand U2087 (N_2087,N_1836,N_1947);
nand U2088 (N_2088,N_1911,N_1933);
or U2089 (N_2089,N_1752,N_1937);
xor U2090 (N_2090,N_1938,N_1814);
nand U2091 (N_2091,N_1760,N_1785);
or U2092 (N_2092,N_1972,N_1879);
xnor U2093 (N_2093,N_1946,N_1807);
or U2094 (N_2094,N_1850,N_1876);
and U2095 (N_2095,N_1920,N_1772);
and U2096 (N_2096,N_1798,N_1808);
or U2097 (N_2097,N_1897,N_1767);
nand U2098 (N_2098,N_1991,N_1838);
nor U2099 (N_2099,N_1824,N_1833);
or U2100 (N_2100,N_1822,N_1974);
nor U2101 (N_2101,N_1844,N_1753);
and U2102 (N_2102,N_1928,N_1787);
or U2103 (N_2103,N_1841,N_1917);
xnor U2104 (N_2104,N_1898,N_1856);
and U2105 (N_2105,N_1989,N_1901);
and U2106 (N_2106,N_1820,N_1811);
or U2107 (N_2107,N_1780,N_1953);
nor U2108 (N_2108,N_1962,N_1834);
nor U2109 (N_2109,N_1786,N_1825);
and U2110 (N_2110,N_1764,N_1792);
and U2111 (N_2111,N_1757,N_1842);
xor U2112 (N_2112,N_1788,N_1855);
and U2113 (N_2113,N_1892,N_1981);
and U2114 (N_2114,N_1862,N_1948);
nor U2115 (N_2115,N_1874,N_1857);
xor U2116 (N_2116,N_1805,N_1810);
and U2117 (N_2117,N_1755,N_1765);
nand U2118 (N_2118,N_1872,N_1960);
nor U2119 (N_2119,N_1837,N_1766);
and U2120 (N_2120,N_1846,N_1908);
xnor U2121 (N_2121,N_1977,N_1769);
or U2122 (N_2122,N_1771,N_1919);
or U2123 (N_2123,N_1878,N_1819);
nor U2124 (N_2124,N_1778,N_1831);
nor U2125 (N_2125,N_1846,N_1877);
nor U2126 (N_2126,N_1876,N_1750);
or U2127 (N_2127,N_1799,N_1950);
nand U2128 (N_2128,N_1939,N_1762);
nor U2129 (N_2129,N_1924,N_1793);
xnor U2130 (N_2130,N_1843,N_1988);
nor U2131 (N_2131,N_1909,N_1973);
xor U2132 (N_2132,N_1990,N_1755);
or U2133 (N_2133,N_1863,N_1987);
or U2134 (N_2134,N_1758,N_1847);
nor U2135 (N_2135,N_1890,N_1756);
nor U2136 (N_2136,N_1988,N_1955);
nand U2137 (N_2137,N_1938,N_1830);
nand U2138 (N_2138,N_1826,N_1801);
and U2139 (N_2139,N_1978,N_1861);
xor U2140 (N_2140,N_1998,N_1767);
nor U2141 (N_2141,N_1967,N_1934);
and U2142 (N_2142,N_1824,N_1933);
nand U2143 (N_2143,N_1815,N_1912);
nand U2144 (N_2144,N_1976,N_1789);
and U2145 (N_2145,N_1817,N_1882);
and U2146 (N_2146,N_1769,N_1950);
xnor U2147 (N_2147,N_1772,N_1875);
or U2148 (N_2148,N_1904,N_1858);
and U2149 (N_2149,N_1850,N_1832);
nor U2150 (N_2150,N_1950,N_1961);
nor U2151 (N_2151,N_1847,N_1863);
nor U2152 (N_2152,N_1892,N_1832);
and U2153 (N_2153,N_1836,N_1872);
xor U2154 (N_2154,N_1813,N_1843);
xor U2155 (N_2155,N_1891,N_1773);
and U2156 (N_2156,N_1783,N_1924);
nand U2157 (N_2157,N_1854,N_1849);
and U2158 (N_2158,N_1999,N_1785);
nor U2159 (N_2159,N_1900,N_1950);
nor U2160 (N_2160,N_1815,N_1829);
or U2161 (N_2161,N_1960,N_1826);
xor U2162 (N_2162,N_1883,N_1829);
and U2163 (N_2163,N_1868,N_1808);
nand U2164 (N_2164,N_1971,N_1784);
and U2165 (N_2165,N_1804,N_1920);
nand U2166 (N_2166,N_1872,N_1829);
nor U2167 (N_2167,N_1782,N_1785);
nand U2168 (N_2168,N_1941,N_1993);
or U2169 (N_2169,N_1872,N_1976);
nor U2170 (N_2170,N_1797,N_1998);
nor U2171 (N_2171,N_1760,N_1832);
and U2172 (N_2172,N_1922,N_1798);
nand U2173 (N_2173,N_1986,N_1821);
or U2174 (N_2174,N_1996,N_1800);
nand U2175 (N_2175,N_1859,N_1836);
and U2176 (N_2176,N_1895,N_1959);
and U2177 (N_2177,N_1851,N_1946);
xnor U2178 (N_2178,N_1760,N_1960);
xnor U2179 (N_2179,N_1882,N_1985);
nand U2180 (N_2180,N_1788,N_1818);
or U2181 (N_2181,N_1926,N_1777);
xor U2182 (N_2182,N_1946,N_1855);
xor U2183 (N_2183,N_1958,N_1783);
and U2184 (N_2184,N_1903,N_1787);
nand U2185 (N_2185,N_1916,N_1778);
nor U2186 (N_2186,N_1974,N_1758);
nand U2187 (N_2187,N_1861,N_1785);
and U2188 (N_2188,N_1877,N_1844);
nand U2189 (N_2189,N_1780,N_1894);
xnor U2190 (N_2190,N_1936,N_1871);
xor U2191 (N_2191,N_1991,N_1966);
nor U2192 (N_2192,N_1818,N_1781);
or U2193 (N_2193,N_1864,N_1938);
or U2194 (N_2194,N_1979,N_1824);
nand U2195 (N_2195,N_1865,N_1767);
nand U2196 (N_2196,N_1914,N_1795);
or U2197 (N_2197,N_1919,N_1940);
nand U2198 (N_2198,N_1977,N_1996);
and U2199 (N_2199,N_1822,N_1808);
and U2200 (N_2200,N_1842,N_1750);
or U2201 (N_2201,N_1913,N_1803);
or U2202 (N_2202,N_1989,N_1914);
nor U2203 (N_2203,N_1927,N_1912);
nand U2204 (N_2204,N_1812,N_1947);
xnor U2205 (N_2205,N_1871,N_1921);
nor U2206 (N_2206,N_1923,N_1770);
nor U2207 (N_2207,N_1833,N_1911);
xnor U2208 (N_2208,N_1974,N_1959);
nand U2209 (N_2209,N_1776,N_1894);
xnor U2210 (N_2210,N_1894,N_1846);
nand U2211 (N_2211,N_1866,N_1949);
and U2212 (N_2212,N_1760,N_1780);
nand U2213 (N_2213,N_1796,N_1784);
nor U2214 (N_2214,N_1760,N_1951);
xor U2215 (N_2215,N_1813,N_1828);
xor U2216 (N_2216,N_1950,N_1782);
nand U2217 (N_2217,N_1914,N_1988);
xnor U2218 (N_2218,N_1769,N_1900);
xnor U2219 (N_2219,N_1765,N_1760);
xnor U2220 (N_2220,N_1815,N_1941);
nor U2221 (N_2221,N_1968,N_1913);
and U2222 (N_2222,N_1855,N_1822);
and U2223 (N_2223,N_1802,N_1803);
nand U2224 (N_2224,N_1825,N_1779);
and U2225 (N_2225,N_1766,N_1936);
nand U2226 (N_2226,N_1973,N_1937);
xnor U2227 (N_2227,N_1894,N_1964);
xor U2228 (N_2228,N_1828,N_1800);
nor U2229 (N_2229,N_1846,N_1760);
or U2230 (N_2230,N_1830,N_1965);
nor U2231 (N_2231,N_1763,N_1853);
xor U2232 (N_2232,N_1998,N_1984);
xnor U2233 (N_2233,N_1793,N_1931);
nand U2234 (N_2234,N_1793,N_1995);
nand U2235 (N_2235,N_1899,N_1845);
and U2236 (N_2236,N_1828,N_1771);
and U2237 (N_2237,N_1876,N_1910);
xnor U2238 (N_2238,N_1916,N_1906);
and U2239 (N_2239,N_1793,N_1847);
xnor U2240 (N_2240,N_1891,N_1874);
and U2241 (N_2241,N_1981,N_1794);
nor U2242 (N_2242,N_1808,N_1953);
nor U2243 (N_2243,N_1887,N_1967);
or U2244 (N_2244,N_1938,N_1769);
and U2245 (N_2245,N_1789,N_1750);
nor U2246 (N_2246,N_1920,N_1880);
xor U2247 (N_2247,N_1822,N_1873);
xor U2248 (N_2248,N_1864,N_1984);
xor U2249 (N_2249,N_1754,N_1821);
nand U2250 (N_2250,N_2084,N_2117);
nor U2251 (N_2251,N_2234,N_2114);
xor U2252 (N_2252,N_2238,N_2175);
and U2253 (N_2253,N_2135,N_2094);
or U2254 (N_2254,N_2224,N_2227);
and U2255 (N_2255,N_2170,N_2027);
and U2256 (N_2256,N_2022,N_2233);
and U2257 (N_2257,N_2156,N_2196);
xor U2258 (N_2258,N_2107,N_2204);
xor U2259 (N_2259,N_2006,N_2192);
or U2260 (N_2260,N_2120,N_2216);
xnor U2261 (N_2261,N_2182,N_2174);
nand U2262 (N_2262,N_2051,N_2037);
nand U2263 (N_2263,N_2069,N_2024);
nand U2264 (N_2264,N_2147,N_2173);
xnor U2265 (N_2265,N_2241,N_2000);
or U2266 (N_2266,N_2104,N_2005);
nor U2267 (N_2267,N_2124,N_2091);
nand U2268 (N_2268,N_2245,N_2096);
xnor U2269 (N_2269,N_2103,N_2026);
nor U2270 (N_2270,N_2058,N_2187);
nand U2271 (N_2271,N_2034,N_2001);
and U2272 (N_2272,N_2041,N_2194);
and U2273 (N_2273,N_2039,N_2171);
xor U2274 (N_2274,N_2219,N_2060);
or U2275 (N_2275,N_2186,N_2073);
nor U2276 (N_2276,N_2113,N_2032);
xnor U2277 (N_2277,N_2072,N_2118);
nor U2278 (N_2278,N_2137,N_2098);
or U2279 (N_2279,N_2248,N_2221);
nor U2280 (N_2280,N_2062,N_2089);
and U2281 (N_2281,N_2035,N_2150);
and U2282 (N_2282,N_2016,N_2126);
and U2283 (N_2283,N_2085,N_2212);
nand U2284 (N_2284,N_2217,N_2002);
nand U2285 (N_2285,N_2246,N_2095);
nand U2286 (N_2286,N_2047,N_2213);
and U2287 (N_2287,N_2045,N_2151);
nor U2288 (N_2288,N_2179,N_2097);
and U2289 (N_2289,N_2018,N_2209);
nand U2290 (N_2290,N_2180,N_2009);
and U2291 (N_2291,N_2081,N_2012);
xor U2292 (N_2292,N_2166,N_2243);
xnor U2293 (N_2293,N_2228,N_2049);
nand U2294 (N_2294,N_2230,N_2055);
and U2295 (N_2295,N_2004,N_2019);
nand U2296 (N_2296,N_2141,N_2070);
xnor U2297 (N_2297,N_2057,N_2202);
nor U2298 (N_2298,N_2122,N_2043);
nand U2299 (N_2299,N_2169,N_2152);
xnor U2300 (N_2300,N_2007,N_2010);
nand U2301 (N_2301,N_2242,N_2168);
nor U2302 (N_2302,N_2082,N_2108);
and U2303 (N_2303,N_2249,N_2237);
nand U2304 (N_2304,N_2240,N_2208);
nor U2305 (N_2305,N_2033,N_2076);
nor U2306 (N_2306,N_2079,N_2064);
nand U2307 (N_2307,N_2074,N_2223);
nand U2308 (N_2308,N_2183,N_2106);
and U2309 (N_2309,N_2176,N_2052);
and U2310 (N_2310,N_2139,N_2188);
xnor U2311 (N_2311,N_2046,N_2142);
nor U2312 (N_2312,N_2115,N_2203);
and U2313 (N_2313,N_2112,N_2236);
and U2314 (N_2314,N_2189,N_2028);
nand U2315 (N_2315,N_2083,N_2056);
nor U2316 (N_2316,N_2080,N_2164);
nand U2317 (N_2317,N_2077,N_2144);
and U2318 (N_2318,N_2021,N_2065);
nor U2319 (N_2319,N_2100,N_2201);
nor U2320 (N_2320,N_2232,N_2239);
nand U2321 (N_2321,N_2149,N_2143);
xor U2322 (N_2322,N_2119,N_2133);
nor U2323 (N_2323,N_2071,N_2014);
nand U2324 (N_2324,N_2140,N_2178);
or U2325 (N_2325,N_2042,N_2154);
xor U2326 (N_2326,N_2099,N_2138);
xor U2327 (N_2327,N_2134,N_2226);
or U2328 (N_2328,N_2193,N_2127);
or U2329 (N_2329,N_2092,N_2078);
and U2330 (N_2330,N_2125,N_2054);
or U2331 (N_2331,N_2067,N_2088);
xor U2332 (N_2332,N_2132,N_2093);
xor U2333 (N_2333,N_2148,N_2235);
xor U2334 (N_2334,N_2244,N_2008);
nand U2335 (N_2335,N_2031,N_2185);
or U2336 (N_2336,N_2247,N_2162);
nor U2337 (N_2337,N_2158,N_2214);
nor U2338 (N_2338,N_2190,N_2038);
nor U2339 (N_2339,N_2116,N_2066);
and U2340 (N_2340,N_2068,N_2205);
nor U2341 (N_2341,N_2159,N_2050);
and U2342 (N_2342,N_2109,N_2121);
nand U2343 (N_2343,N_2030,N_2101);
nand U2344 (N_2344,N_2195,N_2200);
or U2345 (N_2345,N_2130,N_2197);
or U2346 (N_2346,N_2044,N_2211);
nor U2347 (N_2347,N_2131,N_2025);
and U2348 (N_2348,N_2123,N_2199);
and U2349 (N_2349,N_2040,N_2129);
and U2350 (N_2350,N_2036,N_2160);
nand U2351 (N_2351,N_2155,N_2015);
nand U2352 (N_2352,N_2048,N_2017);
nand U2353 (N_2353,N_2087,N_2153);
or U2354 (N_2354,N_2231,N_2215);
or U2355 (N_2355,N_2157,N_2229);
xor U2356 (N_2356,N_2172,N_2029);
nand U2357 (N_2357,N_2003,N_2063);
nor U2358 (N_2358,N_2013,N_2090);
nand U2359 (N_2359,N_2206,N_2163);
nor U2360 (N_2360,N_2184,N_2161);
nor U2361 (N_2361,N_2220,N_2105);
nand U2362 (N_2362,N_2177,N_2110);
or U2363 (N_2363,N_2165,N_2020);
nor U2364 (N_2364,N_2167,N_2075);
and U2365 (N_2365,N_2111,N_2128);
xor U2366 (N_2366,N_2061,N_2023);
nor U2367 (N_2367,N_2011,N_2136);
and U2368 (N_2368,N_2181,N_2146);
or U2369 (N_2369,N_2145,N_2207);
nand U2370 (N_2370,N_2053,N_2218);
nand U2371 (N_2371,N_2210,N_2225);
nor U2372 (N_2372,N_2102,N_2222);
or U2373 (N_2373,N_2198,N_2059);
nor U2374 (N_2374,N_2191,N_2086);
nor U2375 (N_2375,N_2153,N_2147);
or U2376 (N_2376,N_2100,N_2037);
xor U2377 (N_2377,N_2094,N_2230);
xor U2378 (N_2378,N_2064,N_2076);
nand U2379 (N_2379,N_2076,N_2056);
nor U2380 (N_2380,N_2202,N_2135);
or U2381 (N_2381,N_2189,N_2151);
or U2382 (N_2382,N_2177,N_2180);
nand U2383 (N_2383,N_2084,N_2161);
and U2384 (N_2384,N_2162,N_2063);
xor U2385 (N_2385,N_2123,N_2183);
nand U2386 (N_2386,N_2163,N_2164);
xnor U2387 (N_2387,N_2046,N_2028);
or U2388 (N_2388,N_2102,N_2121);
nor U2389 (N_2389,N_2007,N_2062);
and U2390 (N_2390,N_2001,N_2020);
nand U2391 (N_2391,N_2144,N_2026);
or U2392 (N_2392,N_2147,N_2012);
and U2393 (N_2393,N_2023,N_2091);
or U2394 (N_2394,N_2194,N_2188);
and U2395 (N_2395,N_2142,N_2198);
and U2396 (N_2396,N_2068,N_2145);
nand U2397 (N_2397,N_2226,N_2247);
nor U2398 (N_2398,N_2020,N_2231);
nand U2399 (N_2399,N_2054,N_2018);
and U2400 (N_2400,N_2220,N_2043);
or U2401 (N_2401,N_2040,N_2089);
nand U2402 (N_2402,N_2206,N_2099);
xnor U2403 (N_2403,N_2078,N_2104);
nand U2404 (N_2404,N_2103,N_2161);
and U2405 (N_2405,N_2106,N_2057);
nor U2406 (N_2406,N_2071,N_2232);
xnor U2407 (N_2407,N_2198,N_2053);
xor U2408 (N_2408,N_2117,N_2205);
or U2409 (N_2409,N_2028,N_2097);
nor U2410 (N_2410,N_2000,N_2081);
nor U2411 (N_2411,N_2225,N_2104);
nand U2412 (N_2412,N_2067,N_2134);
and U2413 (N_2413,N_2244,N_2225);
and U2414 (N_2414,N_2132,N_2024);
nor U2415 (N_2415,N_2007,N_2168);
nor U2416 (N_2416,N_2121,N_2207);
and U2417 (N_2417,N_2044,N_2112);
nand U2418 (N_2418,N_2107,N_2103);
and U2419 (N_2419,N_2040,N_2206);
or U2420 (N_2420,N_2245,N_2076);
or U2421 (N_2421,N_2082,N_2245);
xor U2422 (N_2422,N_2012,N_2215);
or U2423 (N_2423,N_2043,N_2157);
or U2424 (N_2424,N_2225,N_2075);
nand U2425 (N_2425,N_2106,N_2238);
nor U2426 (N_2426,N_2117,N_2063);
xor U2427 (N_2427,N_2249,N_2154);
xor U2428 (N_2428,N_2026,N_2151);
or U2429 (N_2429,N_2051,N_2191);
nor U2430 (N_2430,N_2068,N_2085);
nor U2431 (N_2431,N_2131,N_2141);
or U2432 (N_2432,N_2005,N_2226);
xnor U2433 (N_2433,N_2232,N_2025);
nand U2434 (N_2434,N_2000,N_2217);
and U2435 (N_2435,N_2066,N_2133);
nor U2436 (N_2436,N_2243,N_2057);
nand U2437 (N_2437,N_2162,N_2031);
xnor U2438 (N_2438,N_2091,N_2108);
xnor U2439 (N_2439,N_2099,N_2059);
or U2440 (N_2440,N_2173,N_2209);
nor U2441 (N_2441,N_2159,N_2249);
nor U2442 (N_2442,N_2001,N_2067);
nor U2443 (N_2443,N_2053,N_2247);
or U2444 (N_2444,N_2000,N_2162);
xor U2445 (N_2445,N_2055,N_2148);
nor U2446 (N_2446,N_2236,N_2230);
or U2447 (N_2447,N_2055,N_2147);
nand U2448 (N_2448,N_2111,N_2074);
or U2449 (N_2449,N_2004,N_2150);
xnor U2450 (N_2450,N_2043,N_2076);
and U2451 (N_2451,N_2084,N_2143);
and U2452 (N_2452,N_2019,N_2248);
nand U2453 (N_2453,N_2241,N_2113);
nand U2454 (N_2454,N_2113,N_2046);
and U2455 (N_2455,N_2203,N_2003);
nand U2456 (N_2456,N_2057,N_2181);
nor U2457 (N_2457,N_2249,N_2087);
or U2458 (N_2458,N_2129,N_2079);
and U2459 (N_2459,N_2207,N_2054);
and U2460 (N_2460,N_2057,N_2132);
xor U2461 (N_2461,N_2120,N_2155);
nor U2462 (N_2462,N_2196,N_2008);
nor U2463 (N_2463,N_2046,N_2165);
and U2464 (N_2464,N_2029,N_2068);
and U2465 (N_2465,N_2191,N_2205);
nand U2466 (N_2466,N_2073,N_2109);
nand U2467 (N_2467,N_2162,N_2066);
xnor U2468 (N_2468,N_2213,N_2085);
and U2469 (N_2469,N_2248,N_2044);
or U2470 (N_2470,N_2101,N_2060);
or U2471 (N_2471,N_2025,N_2155);
nor U2472 (N_2472,N_2092,N_2207);
xnor U2473 (N_2473,N_2191,N_2021);
or U2474 (N_2474,N_2025,N_2240);
or U2475 (N_2475,N_2221,N_2166);
xor U2476 (N_2476,N_2211,N_2238);
or U2477 (N_2477,N_2055,N_2042);
nand U2478 (N_2478,N_2046,N_2009);
xor U2479 (N_2479,N_2021,N_2235);
xnor U2480 (N_2480,N_2146,N_2125);
and U2481 (N_2481,N_2162,N_2130);
nand U2482 (N_2482,N_2186,N_2041);
or U2483 (N_2483,N_2068,N_2105);
xor U2484 (N_2484,N_2038,N_2238);
xor U2485 (N_2485,N_2157,N_2155);
and U2486 (N_2486,N_2231,N_2219);
or U2487 (N_2487,N_2205,N_2115);
or U2488 (N_2488,N_2208,N_2143);
nand U2489 (N_2489,N_2228,N_2042);
or U2490 (N_2490,N_2095,N_2202);
nor U2491 (N_2491,N_2049,N_2245);
nand U2492 (N_2492,N_2110,N_2174);
nor U2493 (N_2493,N_2027,N_2204);
or U2494 (N_2494,N_2046,N_2104);
and U2495 (N_2495,N_2104,N_2073);
and U2496 (N_2496,N_2039,N_2137);
and U2497 (N_2497,N_2106,N_2070);
nor U2498 (N_2498,N_2176,N_2182);
and U2499 (N_2499,N_2167,N_2160);
and U2500 (N_2500,N_2428,N_2251);
and U2501 (N_2501,N_2332,N_2317);
xnor U2502 (N_2502,N_2406,N_2469);
nand U2503 (N_2503,N_2350,N_2436);
nor U2504 (N_2504,N_2384,N_2293);
and U2505 (N_2505,N_2298,N_2262);
nor U2506 (N_2506,N_2253,N_2392);
nor U2507 (N_2507,N_2473,N_2365);
or U2508 (N_2508,N_2349,N_2418);
xor U2509 (N_2509,N_2379,N_2300);
nor U2510 (N_2510,N_2296,N_2328);
and U2511 (N_2511,N_2258,N_2311);
xnor U2512 (N_2512,N_2427,N_2401);
nor U2513 (N_2513,N_2285,N_2445);
xor U2514 (N_2514,N_2476,N_2489);
nor U2515 (N_2515,N_2268,N_2290);
nor U2516 (N_2516,N_2439,N_2481);
xnor U2517 (N_2517,N_2419,N_2351);
xnor U2518 (N_2518,N_2386,N_2466);
or U2519 (N_2519,N_2259,N_2441);
and U2520 (N_2520,N_2307,N_2291);
nand U2521 (N_2521,N_2448,N_2432);
or U2522 (N_2522,N_2424,N_2279);
xor U2523 (N_2523,N_2348,N_2316);
nor U2524 (N_2524,N_2366,N_2375);
nand U2525 (N_2525,N_2437,N_2413);
and U2526 (N_2526,N_2312,N_2475);
or U2527 (N_2527,N_2255,N_2455);
or U2528 (N_2528,N_2494,N_2313);
and U2529 (N_2529,N_2373,N_2376);
and U2530 (N_2530,N_2431,N_2256);
and U2531 (N_2531,N_2433,N_2359);
or U2532 (N_2532,N_2381,N_2411);
and U2533 (N_2533,N_2407,N_2389);
or U2534 (N_2534,N_2490,N_2440);
or U2535 (N_2535,N_2370,N_2397);
nor U2536 (N_2536,N_2341,N_2326);
and U2537 (N_2537,N_2415,N_2474);
and U2538 (N_2538,N_2499,N_2402);
nor U2539 (N_2539,N_2382,N_2412);
nand U2540 (N_2540,N_2324,N_2367);
or U2541 (N_2541,N_2453,N_2346);
nand U2542 (N_2542,N_2467,N_2353);
nand U2543 (N_2543,N_2263,N_2340);
xor U2544 (N_2544,N_2327,N_2352);
and U2545 (N_2545,N_2383,N_2292);
and U2546 (N_2546,N_2387,N_2369);
and U2547 (N_2547,N_2484,N_2260);
nor U2548 (N_2548,N_2414,N_2470);
xor U2549 (N_2549,N_2452,N_2498);
or U2550 (N_2550,N_2496,N_2257);
xnor U2551 (N_2551,N_2493,N_2450);
nand U2552 (N_2552,N_2342,N_2462);
xnor U2553 (N_2553,N_2355,N_2425);
or U2554 (N_2554,N_2449,N_2480);
nor U2555 (N_2555,N_2338,N_2495);
or U2556 (N_2556,N_2457,N_2388);
or U2557 (N_2557,N_2354,N_2302);
nor U2558 (N_2558,N_2423,N_2314);
nand U2559 (N_2559,N_2271,N_2408);
and U2560 (N_2560,N_2363,N_2405);
nor U2561 (N_2561,N_2309,N_2461);
nor U2562 (N_2562,N_2451,N_2336);
nand U2563 (N_2563,N_2435,N_2273);
or U2564 (N_2564,N_2357,N_2479);
xnor U2565 (N_2565,N_2409,N_2360);
nor U2566 (N_2566,N_2318,N_2377);
xnor U2567 (N_2567,N_2277,N_2390);
or U2568 (N_2568,N_2400,N_2454);
and U2569 (N_2569,N_2492,N_2456);
nor U2570 (N_2570,N_2358,N_2497);
nor U2571 (N_2571,N_2361,N_2443);
and U2572 (N_2572,N_2344,N_2446);
nor U2573 (N_2573,N_2275,N_2422);
or U2574 (N_2574,N_2305,N_2398);
nand U2575 (N_2575,N_2345,N_2485);
xor U2576 (N_2576,N_2394,N_2334);
and U2577 (N_2577,N_2280,N_2252);
or U2578 (N_2578,N_2491,N_2308);
xnor U2579 (N_2579,N_2274,N_2465);
nor U2580 (N_2580,N_2306,N_2267);
nor U2581 (N_2581,N_2368,N_2269);
xnor U2582 (N_2582,N_2320,N_2458);
xnor U2583 (N_2583,N_2289,N_2270);
nand U2584 (N_2584,N_2347,N_2438);
nor U2585 (N_2585,N_2371,N_2385);
and U2586 (N_2586,N_2281,N_2444);
and U2587 (N_2587,N_2404,N_2323);
xnor U2588 (N_2588,N_2471,N_2319);
or U2589 (N_2589,N_2378,N_2321);
nand U2590 (N_2590,N_2362,N_2297);
and U2591 (N_2591,N_2287,N_2460);
nor U2592 (N_2592,N_2464,N_2356);
nor U2593 (N_2593,N_2488,N_2459);
and U2594 (N_2594,N_2303,N_2393);
nand U2595 (N_2595,N_2261,N_2380);
or U2596 (N_2596,N_2483,N_2468);
xor U2597 (N_2597,N_2487,N_2421);
and U2598 (N_2598,N_2482,N_2330);
nand U2599 (N_2599,N_2343,N_2429);
and U2600 (N_2600,N_2410,N_2286);
nand U2601 (N_2601,N_2301,N_2403);
and U2602 (N_2602,N_2272,N_2265);
nand U2603 (N_2603,N_2283,N_2374);
xor U2604 (N_2604,N_2282,N_2477);
xnor U2605 (N_2605,N_2364,N_2331);
nand U2606 (N_2606,N_2417,N_2276);
xor U2607 (N_2607,N_2420,N_2254);
nor U2608 (N_2608,N_2337,N_2399);
xor U2609 (N_2609,N_2416,N_2434);
and U2610 (N_2610,N_2333,N_2310);
nand U2611 (N_2611,N_2284,N_2335);
xor U2612 (N_2612,N_2322,N_2426);
nand U2613 (N_2613,N_2486,N_2250);
or U2614 (N_2614,N_2391,N_2442);
nor U2615 (N_2615,N_2372,N_2304);
nor U2616 (N_2616,N_2299,N_2430);
or U2617 (N_2617,N_2329,N_2472);
nand U2618 (N_2618,N_2266,N_2294);
xor U2619 (N_2619,N_2339,N_2264);
nor U2620 (N_2620,N_2447,N_2315);
nand U2621 (N_2621,N_2463,N_2325);
or U2622 (N_2622,N_2295,N_2478);
nor U2623 (N_2623,N_2395,N_2396);
and U2624 (N_2624,N_2278,N_2288);
nor U2625 (N_2625,N_2328,N_2369);
xor U2626 (N_2626,N_2429,N_2360);
or U2627 (N_2627,N_2421,N_2491);
or U2628 (N_2628,N_2483,N_2277);
and U2629 (N_2629,N_2344,N_2294);
xnor U2630 (N_2630,N_2492,N_2380);
or U2631 (N_2631,N_2302,N_2281);
nor U2632 (N_2632,N_2348,N_2398);
xor U2633 (N_2633,N_2283,N_2253);
and U2634 (N_2634,N_2297,N_2441);
nand U2635 (N_2635,N_2418,N_2392);
nand U2636 (N_2636,N_2298,N_2487);
and U2637 (N_2637,N_2431,N_2358);
and U2638 (N_2638,N_2467,N_2442);
nor U2639 (N_2639,N_2353,N_2487);
or U2640 (N_2640,N_2287,N_2355);
and U2641 (N_2641,N_2407,N_2374);
and U2642 (N_2642,N_2279,N_2438);
or U2643 (N_2643,N_2473,N_2274);
or U2644 (N_2644,N_2296,N_2433);
xnor U2645 (N_2645,N_2351,N_2319);
and U2646 (N_2646,N_2288,N_2310);
and U2647 (N_2647,N_2273,N_2403);
xnor U2648 (N_2648,N_2414,N_2396);
nand U2649 (N_2649,N_2471,N_2420);
and U2650 (N_2650,N_2270,N_2254);
nor U2651 (N_2651,N_2386,N_2279);
or U2652 (N_2652,N_2318,N_2332);
and U2653 (N_2653,N_2494,N_2280);
and U2654 (N_2654,N_2430,N_2482);
xnor U2655 (N_2655,N_2468,N_2317);
xnor U2656 (N_2656,N_2388,N_2255);
and U2657 (N_2657,N_2455,N_2378);
nand U2658 (N_2658,N_2421,N_2470);
nor U2659 (N_2659,N_2397,N_2476);
nor U2660 (N_2660,N_2328,N_2251);
nor U2661 (N_2661,N_2381,N_2354);
or U2662 (N_2662,N_2302,N_2442);
nand U2663 (N_2663,N_2467,N_2415);
xor U2664 (N_2664,N_2269,N_2328);
nand U2665 (N_2665,N_2373,N_2358);
and U2666 (N_2666,N_2411,N_2311);
nor U2667 (N_2667,N_2271,N_2279);
nand U2668 (N_2668,N_2400,N_2322);
nand U2669 (N_2669,N_2265,N_2273);
xor U2670 (N_2670,N_2309,N_2430);
and U2671 (N_2671,N_2415,N_2343);
and U2672 (N_2672,N_2497,N_2281);
nand U2673 (N_2673,N_2497,N_2410);
or U2674 (N_2674,N_2469,N_2375);
xnor U2675 (N_2675,N_2416,N_2260);
xnor U2676 (N_2676,N_2408,N_2419);
nor U2677 (N_2677,N_2398,N_2473);
and U2678 (N_2678,N_2437,N_2261);
and U2679 (N_2679,N_2439,N_2300);
nand U2680 (N_2680,N_2297,N_2471);
nand U2681 (N_2681,N_2377,N_2409);
nor U2682 (N_2682,N_2394,N_2309);
or U2683 (N_2683,N_2461,N_2437);
xnor U2684 (N_2684,N_2347,N_2371);
and U2685 (N_2685,N_2261,N_2375);
nor U2686 (N_2686,N_2371,N_2332);
nor U2687 (N_2687,N_2390,N_2352);
or U2688 (N_2688,N_2311,N_2402);
nor U2689 (N_2689,N_2452,N_2393);
nor U2690 (N_2690,N_2479,N_2451);
or U2691 (N_2691,N_2402,N_2473);
and U2692 (N_2692,N_2432,N_2326);
or U2693 (N_2693,N_2352,N_2318);
and U2694 (N_2694,N_2354,N_2386);
nor U2695 (N_2695,N_2484,N_2307);
or U2696 (N_2696,N_2468,N_2367);
and U2697 (N_2697,N_2336,N_2468);
and U2698 (N_2698,N_2260,N_2438);
and U2699 (N_2699,N_2266,N_2484);
xor U2700 (N_2700,N_2273,N_2368);
xor U2701 (N_2701,N_2266,N_2437);
or U2702 (N_2702,N_2329,N_2366);
nand U2703 (N_2703,N_2465,N_2265);
and U2704 (N_2704,N_2452,N_2302);
xnor U2705 (N_2705,N_2341,N_2312);
nand U2706 (N_2706,N_2461,N_2495);
or U2707 (N_2707,N_2375,N_2487);
and U2708 (N_2708,N_2326,N_2469);
or U2709 (N_2709,N_2316,N_2498);
and U2710 (N_2710,N_2378,N_2255);
nand U2711 (N_2711,N_2309,N_2301);
xor U2712 (N_2712,N_2265,N_2263);
nor U2713 (N_2713,N_2378,N_2344);
nor U2714 (N_2714,N_2427,N_2314);
nor U2715 (N_2715,N_2488,N_2493);
or U2716 (N_2716,N_2497,N_2363);
xor U2717 (N_2717,N_2438,N_2487);
xnor U2718 (N_2718,N_2355,N_2493);
nor U2719 (N_2719,N_2367,N_2369);
and U2720 (N_2720,N_2398,N_2351);
nand U2721 (N_2721,N_2493,N_2462);
and U2722 (N_2722,N_2276,N_2442);
or U2723 (N_2723,N_2269,N_2457);
or U2724 (N_2724,N_2480,N_2488);
or U2725 (N_2725,N_2472,N_2433);
and U2726 (N_2726,N_2251,N_2482);
nand U2727 (N_2727,N_2313,N_2285);
or U2728 (N_2728,N_2377,N_2265);
nor U2729 (N_2729,N_2266,N_2488);
nand U2730 (N_2730,N_2407,N_2250);
or U2731 (N_2731,N_2462,N_2256);
or U2732 (N_2732,N_2362,N_2350);
or U2733 (N_2733,N_2476,N_2404);
nor U2734 (N_2734,N_2422,N_2430);
and U2735 (N_2735,N_2289,N_2377);
xor U2736 (N_2736,N_2491,N_2306);
nor U2737 (N_2737,N_2295,N_2406);
nand U2738 (N_2738,N_2324,N_2303);
nor U2739 (N_2739,N_2260,N_2266);
nand U2740 (N_2740,N_2308,N_2256);
nand U2741 (N_2741,N_2434,N_2353);
nand U2742 (N_2742,N_2388,N_2250);
nand U2743 (N_2743,N_2349,N_2476);
and U2744 (N_2744,N_2282,N_2288);
nand U2745 (N_2745,N_2422,N_2291);
or U2746 (N_2746,N_2396,N_2352);
or U2747 (N_2747,N_2370,N_2480);
nand U2748 (N_2748,N_2308,N_2301);
nor U2749 (N_2749,N_2442,N_2260);
nand U2750 (N_2750,N_2509,N_2648);
nor U2751 (N_2751,N_2722,N_2698);
nand U2752 (N_2752,N_2712,N_2626);
and U2753 (N_2753,N_2514,N_2718);
and U2754 (N_2754,N_2743,N_2518);
nor U2755 (N_2755,N_2611,N_2738);
nor U2756 (N_2756,N_2553,N_2714);
nand U2757 (N_2757,N_2556,N_2634);
and U2758 (N_2758,N_2713,N_2748);
and U2759 (N_2759,N_2547,N_2739);
nand U2760 (N_2760,N_2542,N_2700);
nor U2761 (N_2761,N_2530,N_2597);
or U2762 (N_2762,N_2536,N_2687);
xnor U2763 (N_2763,N_2614,N_2702);
and U2764 (N_2764,N_2528,N_2507);
nand U2765 (N_2765,N_2574,N_2681);
nor U2766 (N_2766,N_2688,N_2603);
and U2767 (N_2767,N_2564,N_2500);
xor U2768 (N_2768,N_2641,N_2502);
nor U2769 (N_2769,N_2607,N_2744);
nand U2770 (N_2770,N_2708,N_2549);
xor U2771 (N_2771,N_2594,N_2562);
nor U2772 (N_2772,N_2673,N_2538);
xnor U2773 (N_2773,N_2736,N_2621);
nand U2774 (N_2774,N_2545,N_2740);
nor U2775 (N_2775,N_2551,N_2719);
and U2776 (N_2776,N_2587,N_2508);
and U2777 (N_2777,N_2720,N_2657);
nand U2778 (N_2778,N_2620,N_2697);
and U2779 (N_2779,N_2576,N_2644);
nand U2780 (N_2780,N_2646,N_2696);
or U2781 (N_2781,N_2554,N_2604);
nand U2782 (N_2782,N_2664,N_2624);
nor U2783 (N_2783,N_2631,N_2636);
xnor U2784 (N_2784,N_2650,N_2680);
or U2785 (N_2785,N_2655,N_2601);
and U2786 (N_2786,N_2663,N_2622);
nor U2787 (N_2787,N_2511,N_2523);
nor U2788 (N_2788,N_2699,N_2555);
nand U2789 (N_2789,N_2570,N_2591);
and U2790 (N_2790,N_2546,N_2513);
and U2791 (N_2791,N_2584,N_2683);
nand U2792 (N_2792,N_2573,N_2617);
or U2793 (N_2793,N_2541,N_2689);
xnor U2794 (N_2794,N_2625,N_2686);
xor U2795 (N_2795,N_2630,N_2726);
or U2796 (N_2796,N_2717,N_2543);
xnor U2797 (N_2797,N_2710,N_2711);
nand U2798 (N_2798,N_2616,N_2745);
xor U2799 (N_2799,N_2608,N_2525);
or U2800 (N_2800,N_2660,N_2749);
and U2801 (N_2801,N_2588,N_2524);
nor U2802 (N_2802,N_2612,N_2674);
nor U2803 (N_2803,N_2552,N_2535);
or U2804 (N_2804,N_2550,N_2519);
nand U2805 (N_2805,N_2737,N_2672);
nand U2806 (N_2806,N_2732,N_2639);
nor U2807 (N_2807,N_2516,N_2501);
and U2808 (N_2808,N_2593,N_2692);
or U2809 (N_2809,N_2503,N_2522);
nor U2810 (N_2810,N_2504,N_2596);
and U2811 (N_2811,N_2721,N_2619);
xnor U2812 (N_2812,N_2532,N_2623);
xor U2813 (N_2813,N_2701,N_2579);
xor U2814 (N_2814,N_2735,N_2685);
or U2815 (N_2815,N_2747,N_2618);
nor U2816 (N_2816,N_2506,N_2684);
and U2817 (N_2817,N_2565,N_2693);
or U2818 (N_2818,N_2557,N_2558);
xnor U2819 (N_2819,N_2581,N_2635);
nor U2820 (N_2820,N_2651,N_2533);
xnor U2821 (N_2821,N_2716,N_2583);
and U2822 (N_2822,N_2540,N_2690);
and U2823 (N_2823,N_2521,N_2649);
xor U2824 (N_2824,N_2569,N_2561);
xor U2825 (N_2825,N_2647,N_2605);
nand U2826 (N_2826,N_2595,N_2633);
nor U2827 (N_2827,N_2531,N_2582);
or U2828 (N_2828,N_2678,N_2715);
nor U2829 (N_2829,N_2534,N_2707);
nor U2830 (N_2830,N_2728,N_2610);
and U2831 (N_2831,N_2592,N_2602);
xnor U2832 (N_2832,N_2643,N_2586);
and U2833 (N_2833,N_2669,N_2599);
nor U2834 (N_2834,N_2529,N_2640);
xnor U2835 (N_2835,N_2632,N_2703);
nor U2836 (N_2836,N_2666,N_2662);
nand U2837 (N_2837,N_2526,N_2559);
or U2838 (N_2838,N_2637,N_2742);
and U2839 (N_2839,N_2567,N_2677);
xor U2840 (N_2840,N_2682,N_2613);
nor U2841 (N_2841,N_2679,N_2590);
and U2842 (N_2842,N_2571,N_2537);
nor U2843 (N_2843,N_2733,N_2512);
or U2844 (N_2844,N_2642,N_2629);
nand U2845 (N_2845,N_2730,N_2695);
nor U2846 (N_2846,N_2645,N_2675);
nand U2847 (N_2847,N_2691,N_2724);
nor U2848 (N_2848,N_2589,N_2568);
nand U2849 (N_2849,N_2560,N_2704);
or U2850 (N_2850,N_2671,N_2723);
and U2851 (N_2851,N_2598,N_2734);
nand U2852 (N_2852,N_2539,N_2609);
xnor U2853 (N_2853,N_2580,N_2676);
xnor U2854 (N_2854,N_2578,N_2665);
nor U2855 (N_2855,N_2577,N_2638);
and U2856 (N_2856,N_2694,N_2548);
nand U2857 (N_2857,N_2709,N_2731);
nor U2858 (N_2858,N_2520,N_2658);
or U2859 (N_2859,N_2515,N_2566);
nand U2860 (N_2860,N_2670,N_2705);
or U2861 (N_2861,N_2667,N_2606);
xnor U2862 (N_2862,N_2563,N_2628);
xnor U2863 (N_2863,N_2654,N_2729);
and U2864 (N_2864,N_2517,N_2706);
nor U2865 (N_2865,N_2668,N_2746);
xor U2866 (N_2866,N_2725,N_2656);
nor U2867 (N_2867,N_2505,N_2527);
xor U2868 (N_2868,N_2575,N_2727);
or U2869 (N_2869,N_2653,N_2572);
nor U2870 (N_2870,N_2585,N_2615);
xnor U2871 (N_2871,N_2544,N_2741);
nand U2872 (N_2872,N_2659,N_2652);
or U2873 (N_2873,N_2661,N_2600);
or U2874 (N_2874,N_2510,N_2627);
or U2875 (N_2875,N_2712,N_2507);
and U2876 (N_2876,N_2527,N_2515);
and U2877 (N_2877,N_2568,N_2517);
xor U2878 (N_2878,N_2673,N_2501);
nand U2879 (N_2879,N_2656,N_2675);
nand U2880 (N_2880,N_2605,N_2664);
or U2881 (N_2881,N_2591,N_2695);
xor U2882 (N_2882,N_2510,N_2647);
and U2883 (N_2883,N_2601,N_2542);
nor U2884 (N_2884,N_2704,N_2561);
nand U2885 (N_2885,N_2539,N_2644);
nand U2886 (N_2886,N_2715,N_2532);
or U2887 (N_2887,N_2549,N_2691);
nand U2888 (N_2888,N_2739,N_2742);
or U2889 (N_2889,N_2513,N_2603);
and U2890 (N_2890,N_2617,N_2654);
or U2891 (N_2891,N_2619,N_2673);
nor U2892 (N_2892,N_2558,N_2538);
xnor U2893 (N_2893,N_2549,N_2713);
nor U2894 (N_2894,N_2538,N_2549);
or U2895 (N_2895,N_2673,N_2541);
or U2896 (N_2896,N_2506,N_2500);
nor U2897 (N_2897,N_2557,N_2565);
and U2898 (N_2898,N_2561,N_2745);
nand U2899 (N_2899,N_2684,N_2525);
xor U2900 (N_2900,N_2552,N_2639);
nor U2901 (N_2901,N_2684,N_2681);
and U2902 (N_2902,N_2500,N_2642);
and U2903 (N_2903,N_2671,N_2615);
or U2904 (N_2904,N_2585,N_2642);
and U2905 (N_2905,N_2646,N_2683);
nor U2906 (N_2906,N_2692,N_2552);
and U2907 (N_2907,N_2557,N_2749);
nor U2908 (N_2908,N_2580,N_2597);
and U2909 (N_2909,N_2511,N_2612);
xnor U2910 (N_2910,N_2526,N_2658);
and U2911 (N_2911,N_2706,N_2680);
nand U2912 (N_2912,N_2543,N_2571);
nor U2913 (N_2913,N_2672,N_2634);
xnor U2914 (N_2914,N_2603,N_2604);
nand U2915 (N_2915,N_2522,N_2620);
xor U2916 (N_2916,N_2699,N_2653);
nor U2917 (N_2917,N_2684,N_2620);
and U2918 (N_2918,N_2748,N_2616);
or U2919 (N_2919,N_2536,N_2722);
nor U2920 (N_2920,N_2596,N_2566);
xor U2921 (N_2921,N_2743,N_2520);
xnor U2922 (N_2922,N_2628,N_2676);
nand U2923 (N_2923,N_2608,N_2516);
and U2924 (N_2924,N_2545,N_2684);
xor U2925 (N_2925,N_2679,N_2719);
or U2926 (N_2926,N_2631,N_2504);
or U2927 (N_2927,N_2638,N_2680);
xnor U2928 (N_2928,N_2515,N_2736);
nor U2929 (N_2929,N_2513,N_2625);
xor U2930 (N_2930,N_2552,N_2553);
or U2931 (N_2931,N_2575,N_2695);
nand U2932 (N_2932,N_2501,N_2665);
xor U2933 (N_2933,N_2651,N_2736);
nor U2934 (N_2934,N_2699,N_2544);
or U2935 (N_2935,N_2711,N_2532);
and U2936 (N_2936,N_2590,N_2544);
or U2937 (N_2937,N_2717,N_2636);
xnor U2938 (N_2938,N_2505,N_2506);
nand U2939 (N_2939,N_2735,N_2583);
and U2940 (N_2940,N_2656,N_2648);
or U2941 (N_2941,N_2526,N_2652);
and U2942 (N_2942,N_2552,N_2580);
nor U2943 (N_2943,N_2660,N_2717);
nand U2944 (N_2944,N_2666,N_2620);
nand U2945 (N_2945,N_2689,N_2558);
nand U2946 (N_2946,N_2664,N_2709);
nand U2947 (N_2947,N_2600,N_2659);
nor U2948 (N_2948,N_2579,N_2690);
or U2949 (N_2949,N_2677,N_2534);
nor U2950 (N_2950,N_2735,N_2726);
and U2951 (N_2951,N_2613,N_2658);
or U2952 (N_2952,N_2526,N_2500);
xor U2953 (N_2953,N_2506,N_2653);
xnor U2954 (N_2954,N_2727,N_2601);
and U2955 (N_2955,N_2548,N_2524);
nand U2956 (N_2956,N_2643,N_2679);
and U2957 (N_2957,N_2595,N_2661);
and U2958 (N_2958,N_2526,N_2655);
or U2959 (N_2959,N_2583,N_2618);
and U2960 (N_2960,N_2587,N_2604);
nor U2961 (N_2961,N_2614,N_2559);
or U2962 (N_2962,N_2665,N_2616);
xor U2963 (N_2963,N_2594,N_2617);
nand U2964 (N_2964,N_2677,N_2511);
or U2965 (N_2965,N_2706,N_2662);
or U2966 (N_2966,N_2530,N_2515);
xor U2967 (N_2967,N_2572,N_2677);
xor U2968 (N_2968,N_2518,N_2726);
xnor U2969 (N_2969,N_2574,N_2514);
or U2970 (N_2970,N_2704,N_2574);
and U2971 (N_2971,N_2609,N_2514);
nand U2972 (N_2972,N_2692,N_2589);
nor U2973 (N_2973,N_2620,N_2701);
nand U2974 (N_2974,N_2737,N_2739);
xnor U2975 (N_2975,N_2705,N_2657);
and U2976 (N_2976,N_2621,N_2644);
or U2977 (N_2977,N_2652,N_2566);
xor U2978 (N_2978,N_2577,N_2541);
xor U2979 (N_2979,N_2660,N_2711);
or U2980 (N_2980,N_2717,N_2572);
nor U2981 (N_2981,N_2704,N_2537);
nand U2982 (N_2982,N_2597,N_2600);
nor U2983 (N_2983,N_2747,N_2652);
and U2984 (N_2984,N_2706,N_2665);
nand U2985 (N_2985,N_2708,N_2600);
nor U2986 (N_2986,N_2590,N_2537);
nor U2987 (N_2987,N_2561,N_2631);
nor U2988 (N_2988,N_2639,N_2597);
nand U2989 (N_2989,N_2734,N_2615);
xor U2990 (N_2990,N_2577,N_2666);
xor U2991 (N_2991,N_2646,N_2703);
and U2992 (N_2992,N_2623,N_2709);
nor U2993 (N_2993,N_2714,N_2501);
nand U2994 (N_2994,N_2648,N_2632);
or U2995 (N_2995,N_2742,N_2504);
or U2996 (N_2996,N_2660,N_2746);
nor U2997 (N_2997,N_2721,N_2644);
or U2998 (N_2998,N_2670,N_2609);
or U2999 (N_2999,N_2661,N_2680);
xor U3000 (N_3000,N_2781,N_2911);
nor U3001 (N_3001,N_2965,N_2786);
or U3002 (N_3002,N_2969,N_2994);
or U3003 (N_3003,N_2909,N_2847);
and U3004 (N_3004,N_2766,N_2944);
nor U3005 (N_3005,N_2820,N_2876);
nand U3006 (N_3006,N_2912,N_2933);
or U3007 (N_3007,N_2760,N_2787);
nor U3008 (N_3008,N_2993,N_2783);
and U3009 (N_3009,N_2849,N_2812);
and U3010 (N_3010,N_2840,N_2916);
xnor U3011 (N_3011,N_2975,N_2929);
and U3012 (N_3012,N_2997,N_2889);
and U3013 (N_3013,N_2770,N_2875);
or U3014 (N_3014,N_2991,N_2850);
or U3015 (N_3015,N_2952,N_2826);
nor U3016 (N_3016,N_2809,N_2830);
xnor U3017 (N_3017,N_2814,N_2871);
nand U3018 (N_3018,N_2962,N_2788);
nor U3019 (N_3019,N_2832,N_2858);
or U3020 (N_3020,N_2884,N_2996);
and U3021 (N_3021,N_2905,N_2921);
xor U3022 (N_3022,N_2880,N_2947);
or U3023 (N_3023,N_2821,N_2968);
nand U3024 (N_3024,N_2899,N_2751);
nand U3025 (N_3025,N_2979,N_2966);
xnor U3026 (N_3026,N_2792,N_2825);
nor U3027 (N_3027,N_2936,N_2948);
and U3028 (N_3028,N_2913,N_2963);
nor U3029 (N_3029,N_2984,N_2903);
or U3030 (N_3030,N_2853,N_2861);
and U3031 (N_3031,N_2855,N_2867);
and U3032 (N_3032,N_2804,N_2805);
or U3033 (N_3033,N_2836,N_2776);
and U3034 (N_3034,N_2828,N_2846);
or U3035 (N_3035,N_2882,N_2822);
or U3036 (N_3036,N_2824,N_2900);
and U3037 (N_3037,N_2810,N_2773);
and U3038 (N_3038,N_2937,N_2961);
or U3039 (N_3039,N_2753,N_2816);
nor U3040 (N_3040,N_2988,N_2920);
xor U3041 (N_3041,N_2977,N_2922);
or U3042 (N_3042,N_2946,N_2790);
nor U3043 (N_3043,N_2960,N_2928);
nand U3044 (N_3044,N_2872,N_2976);
nand U3045 (N_3045,N_2930,N_2887);
xor U3046 (N_3046,N_2935,N_2955);
xnor U3047 (N_3047,N_2754,N_2794);
nor U3048 (N_3048,N_2798,N_2958);
and U3049 (N_3049,N_2949,N_2778);
and U3050 (N_3050,N_2829,N_2756);
or U3051 (N_3051,N_2995,N_2990);
nor U3052 (N_3052,N_2904,N_2980);
nor U3053 (N_3053,N_2981,N_2763);
xor U3054 (N_3054,N_2764,N_2957);
xnor U3055 (N_3055,N_2885,N_2800);
nand U3056 (N_3056,N_2923,N_2869);
and U3057 (N_3057,N_2806,N_2807);
xnor U3058 (N_3058,N_2823,N_2939);
nand U3059 (N_3059,N_2774,N_2973);
or U3060 (N_3060,N_2964,N_2895);
nand U3061 (N_3061,N_2796,N_2779);
or U3062 (N_3062,N_2978,N_2856);
nand U3063 (N_3063,N_2819,N_2950);
nand U3064 (N_3064,N_2896,N_2862);
or U3065 (N_3065,N_2890,N_2924);
nor U3066 (N_3066,N_2883,N_2902);
or U3067 (N_3067,N_2765,N_2908);
and U3068 (N_3068,N_2940,N_2945);
nor U3069 (N_3069,N_2953,N_2992);
and U3070 (N_3070,N_2951,N_2797);
or U3071 (N_3071,N_2793,N_2888);
nand U3072 (N_3072,N_2892,N_2983);
and U3073 (N_3073,N_2854,N_2803);
or U3074 (N_3074,N_2893,N_2851);
nand U3075 (N_3075,N_2915,N_2927);
xor U3076 (N_3076,N_2942,N_2860);
nor U3077 (N_3077,N_2986,N_2813);
and U3078 (N_3078,N_2906,N_2777);
and U3079 (N_3079,N_2866,N_2897);
xnor U3080 (N_3080,N_2757,N_2917);
xor U3081 (N_3081,N_2934,N_2956);
xor U3082 (N_3082,N_2843,N_2811);
nand U3083 (N_3083,N_2891,N_2931);
xor U3084 (N_3084,N_2989,N_2970);
and U3085 (N_3085,N_2827,N_2772);
nand U3086 (N_3086,N_2780,N_2907);
or U3087 (N_3087,N_2879,N_2918);
xor U3088 (N_3088,N_2795,N_2910);
nand U3089 (N_3089,N_2842,N_2998);
nor U3090 (N_3090,N_2971,N_2967);
xor U3091 (N_3091,N_2761,N_2864);
xnor U3092 (N_3092,N_2857,N_2844);
nand U3093 (N_3093,N_2759,N_2785);
xnor U3094 (N_3094,N_2919,N_2752);
or U3095 (N_3095,N_2987,N_2932);
nor U3096 (N_3096,N_2782,N_2767);
or U3097 (N_3097,N_2874,N_2901);
or U3098 (N_3098,N_2926,N_2762);
and U3099 (N_3099,N_2852,N_2954);
xnor U3100 (N_3100,N_2925,N_2818);
xnor U3101 (N_3101,N_2791,N_2834);
xor U3102 (N_3102,N_2817,N_2985);
xnor U3103 (N_3103,N_2877,N_2755);
xnor U3104 (N_3104,N_2999,N_2894);
xor U3105 (N_3105,N_2943,N_2750);
or U3106 (N_3106,N_2848,N_2898);
and U3107 (N_3107,N_2789,N_2775);
nand U3108 (N_3108,N_2873,N_2801);
xor U3109 (N_3109,N_2831,N_2881);
nor U3110 (N_3110,N_2878,N_2802);
xor U3111 (N_3111,N_2808,N_2833);
nor U3112 (N_3112,N_2982,N_2868);
and U3113 (N_3113,N_2941,N_2838);
nor U3114 (N_3114,N_2771,N_2845);
and U3115 (N_3115,N_2758,N_2914);
nand U3116 (N_3116,N_2886,N_2972);
or U3117 (N_3117,N_2870,N_2974);
and U3118 (N_3118,N_2839,N_2863);
xnor U3119 (N_3119,N_2768,N_2938);
or U3120 (N_3120,N_2959,N_2859);
nand U3121 (N_3121,N_2799,N_2769);
or U3122 (N_3122,N_2837,N_2815);
and U3123 (N_3123,N_2835,N_2865);
nor U3124 (N_3124,N_2784,N_2841);
or U3125 (N_3125,N_2836,N_2782);
or U3126 (N_3126,N_2938,N_2827);
xnor U3127 (N_3127,N_2880,N_2823);
or U3128 (N_3128,N_2836,N_2774);
xnor U3129 (N_3129,N_2939,N_2977);
nand U3130 (N_3130,N_2750,N_2899);
and U3131 (N_3131,N_2846,N_2804);
nor U3132 (N_3132,N_2830,N_2763);
xor U3133 (N_3133,N_2851,N_2864);
and U3134 (N_3134,N_2763,N_2888);
nand U3135 (N_3135,N_2779,N_2803);
or U3136 (N_3136,N_2792,N_2766);
nor U3137 (N_3137,N_2946,N_2970);
xnor U3138 (N_3138,N_2903,N_2964);
nand U3139 (N_3139,N_2868,N_2866);
xnor U3140 (N_3140,N_2962,N_2847);
nand U3141 (N_3141,N_2781,N_2811);
and U3142 (N_3142,N_2852,N_2933);
nand U3143 (N_3143,N_2784,N_2834);
nor U3144 (N_3144,N_2971,N_2815);
nand U3145 (N_3145,N_2881,N_2891);
and U3146 (N_3146,N_2873,N_2958);
nand U3147 (N_3147,N_2797,N_2998);
or U3148 (N_3148,N_2807,N_2907);
nand U3149 (N_3149,N_2934,N_2793);
xor U3150 (N_3150,N_2859,N_2946);
or U3151 (N_3151,N_2864,N_2982);
nor U3152 (N_3152,N_2906,N_2874);
or U3153 (N_3153,N_2776,N_2950);
nor U3154 (N_3154,N_2903,N_2919);
nand U3155 (N_3155,N_2946,N_2922);
or U3156 (N_3156,N_2753,N_2924);
nor U3157 (N_3157,N_2792,N_2770);
nor U3158 (N_3158,N_2976,N_2773);
nor U3159 (N_3159,N_2754,N_2930);
xor U3160 (N_3160,N_2851,N_2806);
nor U3161 (N_3161,N_2918,N_2973);
and U3162 (N_3162,N_2820,N_2946);
nand U3163 (N_3163,N_2881,N_2998);
xor U3164 (N_3164,N_2975,N_2864);
nor U3165 (N_3165,N_2844,N_2888);
nand U3166 (N_3166,N_2823,N_2835);
nand U3167 (N_3167,N_2814,N_2843);
nor U3168 (N_3168,N_2763,N_2821);
or U3169 (N_3169,N_2882,N_2978);
or U3170 (N_3170,N_2769,N_2897);
nand U3171 (N_3171,N_2926,N_2830);
nor U3172 (N_3172,N_2967,N_2904);
nand U3173 (N_3173,N_2931,N_2947);
xnor U3174 (N_3174,N_2939,N_2963);
xor U3175 (N_3175,N_2779,N_2973);
xnor U3176 (N_3176,N_2947,N_2797);
nor U3177 (N_3177,N_2788,N_2757);
and U3178 (N_3178,N_2970,N_2773);
xnor U3179 (N_3179,N_2766,N_2890);
or U3180 (N_3180,N_2939,N_2973);
xnor U3181 (N_3181,N_2904,N_2987);
nor U3182 (N_3182,N_2965,N_2796);
or U3183 (N_3183,N_2816,N_2818);
and U3184 (N_3184,N_2862,N_2883);
and U3185 (N_3185,N_2938,N_2783);
nand U3186 (N_3186,N_2773,N_2961);
nor U3187 (N_3187,N_2983,N_2842);
or U3188 (N_3188,N_2828,N_2967);
and U3189 (N_3189,N_2967,N_2935);
and U3190 (N_3190,N_2857,N_2932);
xnor U3191 (N_3191,N_2977,N_2818);
nor U3192 (N_3192,N_2875,N_2882);
and U3193 (N_3193,N_2964,N_2962);
or U3194 (N_3194,N_2809,N_2915);
or U3195 (N_3195,N_2996,N_2819);
xor U3196 (N_3196,N_2794,N_2867);
or U3197 (N_3197,N_2937,N_2782);
or U3198 (N_3198,N_2819,N_2904);
nor U3199 (N_3199,N_2907,N_2997);
and U3200 (N_3200,N_2885,N_2848);
xor U3201 (N_3201,N_2896,N_2981);
nand U3202 (N_3202,N_2906,N_2806);
xnor U3203 (N_3203,N_2946,N_2788);
and U3204 (N_3204,N_2995,N_2786);
and U3205 (N_3205,N_2751,N_2981);
or U3206 (N_3206,N_2772,N_2800);
nor U3207 (N_3207,N_2867,N_2754);
nand U3208 (N_3208,N_2776,N_2932);
or U3209 (N_3209,N_2768,N_2887);
xnor U3210 (N_3210,N_2952,N_2783);
and U3211 (N_3211,N_2915,N_2755);
xnor U3212 (N_3212,N_2824,N_2820);
and U3213 (N_3213,N_2761,N_2805);
nand U3214 (N_3214,N_2776,N_2828);
xnor U3215 (N_3215,N_2843,N_2866);
xnor U3216 (N_3216,N_2849,N_2814);
xor U3217 (N_3217,N_2934,N_2994);
or U3218 (N_3218,N_2752,N_2954);
xnor U3219 (N_3219,N_2904,N_2997);
xor U3220 (N_3220,N_2903,N_2783);
or U3221 (N_3221,N_2983,N_2900);
and U3222 (N_3222,N_2890,N_2840);
or U3223 (N_3223,N_2824,N_2844);
and U3224 (N_3224,N_2900,N_2858);
and U3225 (N_3225,N_2791,N_2900);
xnor U3226 (N_3226,N_2886,N_2754);
and U3227 (N_3227,N_2826,N_2754);
nor U3228 (N_3228,N_2866,N_2924);
and U3229 (N_3229,N_2756,N_2978);
nand U3230 (N_3230,N_2757,N_2991);
nor U3231 (N_3231,N_2821,N_2879);
xor U3232 (N_3232,N_2794,N_2979);
and U3233 (N_3233,N_2847,N_2781);
nand U3234 (N_3234,N_2913,N_2795);
nand U3235 (N_3235,N_2995,N_2941);
and U3236 (N_3236,N_2908,N_2863);
and U3237 (N_3237,N_2807,N_2809);
nand U3238 (N_3238,N_2758,N_2773);
xnor U3239 (N_3239,N_2854,N_2843);
nand U3240 (N_3240,N_2962,N_2979);
nor U3241 (N_3241,N_2922,N_2902);
and U3242 (N_3242,N_2846,N_2956);
and U3243 (N_3243,N_2865,N_2953);
and U3244 (N_3244,N_2805,N_2879);
and U3245 (N_3245,N_2903,N_2891);
or U3246 (N_3246,N_2847,N_2981);
and U3247 (N_3247,N_2974,N_2789);
nand U3248 (N_3248,N_2839,N_2975);
nor U3249 (N_3249,N_2760,N_2827);
xnor U3250 (N_3250,N_3048,N_3244);
xor U3251 (N_3251,N_3186,N_3246);
nand U3252 (N_3252,N_3100,N_3056);
xnor U3253 (N_3253,N_3070,N_3231);
nor U3254 (N_3254,N_3164,N_3233);
or U3255 (N_3255,N_3055,N_3026);
nor U3256 (N_3256,N_3062,N_3166);
nand U3257 (N_3257,N_3082,N_3086);
xnor U3258 (N_3258,N_3022,N_3134);
nor U3259 (N_3259,N_3207,N_3061);
nand U3260 (N_3260,N_3237,N_3119);
and U3261 (N_3261,N_3049,N_3058);
and U3262 (N_3262,N_3219,N_3121);
and U3263 (N_3263,N_3120,N_3093);
nand U3264 (N_3264,N_3118,N_3102);
and U3265 (N_3265,N_3094,N_3226);
nor U3266 (N_3266,N_3156,N_3034);
nand U3267 (N_3267,N_3227,N_3230);
or U3268 (N_3268,N_3232,N_3092);
nor U3269 (N_3269,N_3115,N_3053);
or U3270 (N_3270,N_3003,N_3200);
nor U3271 (N_3271,N_3160,N_3111);
xor U3272 (N_3272,N_3123,N_3054);
nor U3273 (N_3273,N_3190,N_3008);
xor U3274 (N_3274,N_3150,N_3248);
nand U3275 (N_3275,N_3138,N_3019);
or U3276 (N_3276,N_3223,N_3047);
nor U3277 (N_3277,N_3125,N_3103);
or U3278 (N_3278,N_3240,N_3179);
xnor U3279 (N_3279,N_3066,N_3209);
and U3280 (N_3280,N_3069,N_3158);
xnor U3281 (N_3281,N_3162,N_3130);
nor U3282 (N_3282,N_3038,N_3106);
or U3283 (N_3283,N_3076,N_3001);
and U3284 (N_3284,N_3104,N_3098);
or U3285 (N_3285,N_3228,N_3182);
or U3286 (N_3286,N_3028,N_3107);
xor U3287 (N_3287,N_3029,N_3050);
nand U3288 (N_3288,N_3151,N_3091);
and U3289 (N_3289,N_3024,N_3052);
or U3290 (N_3290,N_3243,N_3080);
or U3291 (N_3291,N_3139,N_3206);
and U3292 (N_3292,N_3204,N_3027);
or U3293 (N_3293,N_3195,N_3057);
and U3294 (N_3294,N_3097,N_3157);
nand U3295 (N_3295,N_3033,N_3073);
and U3296 (N_3296,N_3170,N_3000);
nand U3297 (N_3297,N_3149,N_3222);
or U3298 (N_3298,N_3131,N_3212);
nand U3299 (N_3299,N_3011,N_3239);
or U3300 (N_3300,N_3051,N_3099);
or U3301 (N_3301,N_3032,N_3241);
or U3302 (N_3302,N_3064,N_3216);
nor U3303 (N_3303,N_3105,N_3146);
nand U3304 (N_3304,N_3090,N_3013);
nand U3305 (N_3305,N_3109,N_3199);
nand U3306 (N_3306,N_3060,N_3017);
nand U3307 (N_3307,N_3203,N_3014);
or U3308 (N_3308,N_3124,N_3084);
xnor U3309 (N_3309,N_3089,N_3040);
or U3310 (N_3310,N_3213,N_3087);
or U3311 (N_3311,N_3194,N_3191);
or U3312 (N_3312,N_3180,N_3218);
nor U3313 (N_3313,N_3096,N_3137);
nor U3314 (N_3314,N_3249,N_3023);
nor U3315 (N_3315,N_3175,N_3009);
xor U3316 (N_3316,N_3225,N_3046);
or U3317 (N_3317,N_3020,N_3172);
and U3318 (N_3318,N_3152,N_3221);
nand U3319 (N_3319,N_3101,N_3201);
nor U3320 (N_3320,N_3136,N_3002);
and U3321 (N_3321,N_3178,N_3144);
xnor U3322 (N_3322,N_3129,N_3234);
nor U3323 (N_3323,N_3210,N_3042);
or U3324 (N_3324,N_3154,N_3238);
nor U3325 (N_3325,N_3083,N_3181);
or U3326 (N_3326,N_3193,N_3145);
or U3327 (N_3327,N_3037,N_3116);
nor U3328 (N_3328,N_3128,N_3072);
xnor U3329 (N_3329,N_3078,N_3088);
nand U3330 (N_3330,N_3174,N_3079);
and U3331 (N_3331,N_3196,N_3021);
and U3332 (N_3332,N_3059,N_3171);
and U3333 (N_3333,N_3165,N_3177);
nor U3334 (N_3334,N_3016,N_3224);
or U3335 (N_3335,N_3187,N_3067);
or U3336 (N_3336,N_3242,N_3173);
xnor U3337 (N_3337,N_3236,N_3006);
and U3338 (N_3338,N_3198,N_3077);
or U3339 (N_3339,N_3192,N_3012);
xnor U3340 (N_3340,N_3229,N_3122);
or U3341 (N_3341,N_3202,N_3217);
xnor U3342 (N_3342,N_3074,N_3247);
or U3343 (N_3343,N_3007,N_3035);
and U3344 (N_3344,N_3176,N_3235);
and U3345 (N_3345,N_3141,N_3126);
xor U3346 (N_3346,N_3065,N_3183);
nor U3347 (N_3347,N_3025,N_3169);
or U3348 (N_3348,N_3075,N_3041);
or U3349 (N_3349,N_3132,N_3140);
nor U3350 (N_3350,N_3095,N_3043);
nand U3351 (N_3351,N_3147,N_3197);
nand U3352 (N_3352,N_3167,N_3005);
nor U3353 (N_3353,N_3185,N_3112);
and U3354 (N_3354,N_3015,N_3071);
nor U3355 (N_3355,N_3113,N_3081);
nand U3356 (N_3356,N_3110,N_3031);
xor U3357 (N_3357,N_3114,N_3245);
and U3358 (N_3358,N_3161,N_3159);
or U3359 (N_3359,N_3085,N_3214);
and U3360 (N_3360,N_3108,N_3135);
nand U3361 (N_3361,N_3044,N_3215);
nor U3362 (N_3362,N_3063,N_3168);
or U3363 (N_3363,N_3117,N_3045);
and U3364 (N_3364,N_3188,N_3004);
nand U3365 (N_3365,N_3208,N_3039);
xnor U3366 (N_3366,N_3133,N_3184);
nor U3367 (N_3367,N_3036,N_3220);
nand U3368 (N_3368,N_3030,N_3205);
nand U3369 (N_3369,N_3018,N_3127);
or U3370 (N_3370,N_3155,N_3153);
and U3371 (N_3371,N_3163,N_3068);
nor U3372 (N_3372,N_3189,N_3148);
nor U3373 (N_3373,N_3142,N_3211);
nor U3374 (N_3374,N_3143,N_3010);
nand U3375 (N_3375,N_3046,N_3115);
nand U3376 (N_3376,N_3230,N_3123);
nand U3377 (N_3377,N_3058,N_3180);
nand U3378 (N_3378,N_3212,N_3142);
xor U3379 (N_3379,N_3213,N_3024);
xnor U3380 (N_3380,N_3191,N_3246);
xnor U3381 (N_3381,N_3082,N_3187);
xnor U3382 (N_3382,N_3059,N_3204);
or U3383 (N_3383,N_3032,N_3007);
nor U3384 (N_3384,N_3030,N_3045);
nand U3385 (N_3385,N_3182,N_3223);
nand U3386 (N_3386,N_3058,N_3184);
nor U3387 (N_3387,N_3137,N_3229);
nor U3388 (N_3388,N_3134,N_3239);
nor U3389 (N_3389,N_3091,N_3120);
nor U3390 (N_3390,N_3109,N_3007);
nor U3391 (N_3391,N_3060,N_3067);
xnor U3392 (N_3392,N_3208,N_3237);
nor U3393 (N_3393,N_3176,N_3186);
nor U3394 (N_3394,N_3231,N_3225);
or U3395 (N_3395,N_3202,N_3146);
xnor U3396 (N_3396,N_3249,N_3051);
nor U3397 (N_3397,N_3082,N_3129);
nor U3398 (N_3398,N_3097,N_3009);
nand U3399 (N_3399,N_3027,N_3121);
and U3400 (N_3400,N_3085,N_3030);
and U3401 (N_3401,N_3207,N_3175);
xnor U3402 (N_3402,N_3203,N_3155);
xor U3403 (N_3403,N_3000,N_3211);
nor U3404 (N_3404,N_3021,N_3113);
or U3405 (N_3405,N_3171,N_3145);
or U3406 (N_3406,N_3143,N_3217);
nand U3407 (N_3407,N_3077,N_3002);
xnor U3408 (N_3408,N_3244,N_3030);
nand U3409 (N_3409,N_3106,N_3149);
xnor U3410 (N_3410,N_3106,N_3018);
or U3411 (N_3411,N_3210,N_3175);
nand U3412 (N_3412,N_3073,N_3181);
and U3413 (N_3413,N_3201,N_3072);
or U3414 (N_3414,N_3138,N_3219);
or U3415 (N_3415,N_3145,N_3062);
xnor U3416 (N_3416,N_3011,N_3150);
nand U3417 (N_3417,N_3071,N_3124);
and U3418 (N_3418,N_3007,N_3070);
xor U3419 (N_3419,N_3249,N_3116);
xor U3420 (N_3420,N_3069,N_3215);
xor U3421 (N_3421,N_3102,N_3211);
or U3422 (N_3422,N_3072,N_3067);
and U3423 (N_3423,N_3192,N_3205);
xnor U3424 (N_3424,N_3077,N_3214);
nor U3425 (N_3425,N_3244,N_3054);
or U3426 (N_3426,N_3248,N_3008);
xor U3427 (N_3427,N_3248,N_3091);
xnor U3428 (N_3428,N_3179,N_3004);
nand U3429 (N_3429,N_3060,N_3181);
and U3430 (N_3430,N_3194,N_3242);
nor U3431 (N_3431,N_3117,N_3205);
and U3432 (N_3432,N_3166,N_3188);
xnor U3433 (N_3433,N_3102,N_3232);
or U3434 (N_3434,N_3148,N_3116);
nor U3435 (N_3435,N_3242,N_3066);
nor U3436 (N_3436,N_3032,N_3149);
and U3437 (N_3437,N_3213,N_3117);
nor U3438 (N_3438,N_3197,N_3178);
nor U3439 (N_3439,N_3141,N_3186);
or U3440 (N_3440,N_3131,N_3015);
and U3441 (N_3441,N_3146,N_3007);
xor U3442 (N_3442,N_3046,N_3008);
nor U3443 (N_3443,N_3178,N_3024);
and U3444 (N_3444,N_3195,N_3110);
nor U3445 (N_3445,N_3160,N_3123);
nand U3446 (N_3446,N_3030,N_3097);
nor U3447 (N_3447,N_3080,N_3238);
nor U3448 (N_3448,N_3166,N_3042);
xnor U3449 (N_3449,N_3080,N_3206);
xnor U3450 (N_3450,N_3175,N_3008);
xor U3451 (N_3451,N_3099,N_3108);
nand U3452 (N_3452,N_3150,N_3021);
and U3453 (N_3453,N_3224,N_3070);
and U3454 (N_3454,N_3207,N_3115);
and U3455 (N_3455,N_3035,N_3145);
or U3456 (N_3456,N_3002,N_3143);
xnor U3457 (N_3457,N_3247,N_3044);
and U3458 (N_3458,N_3064,N_3248);
nor U3459 (N_3459,N_3106,N_3161);
nand U3460 (N_3460,N_3233,N_3179);
nand U3461 (N_3461,N_3027,N_3248);
xnor U3462 (N_3462,N_3204,N_3057);
xor U3463 (N_3463,N_3111,N_3039);
nor U3464 (N_3464,N_3142,N_3116);
and U3465 (N_3465,N_3096,N_3107);
nor U3466 (N_3466,N_3069,N_3016);
or U3467 (N_3467,N_3117,N_3174);
and U3468 (N_3468,N_3082,N_3016);
or U3469 (N_3469,N_3006,N_3186);
xor U3470 (N_3470,N_3181,N_3190);
nor U3471 (N_3471,N_3184,N_3087);
nand U3472 (N_3472,N_3103,N_3182);
nand U3473 (N_3473,N_3108,N_3247);
or U3474 (N_3474,N_3207,N_3173);
xnor U3475 (N_3475,N_3074,N_3046);
nand U3476 (N_3476,N_3079,N_3146);
nand U3477 (N_3477,N_3114,N_3205);
nand U3478 (N_3478,N_3009,N_3008);
nor U3479 (N_3479,N_3039,N_3001);
xor U3480 (N_3480,N_3234,N_3087);
xor U3481 (N_3481,N_3155,N_3023);
and U3482 (N_3482,N_3207,N_3014);
xor U3483 (N_3483,N_3051,N_3167);
nor U3484 (N_3484,N_3156,N_3170);
and U3485 (N_3485,N_3068,N_3015);
or U3486 (N_3486,N_3117,N_3151);
nand U3487 (N_3487,N_3135,N_3069);
xnor U3488 (N_3488,N_3065,N_3060);
nor U3489 (N_3489,N_3007,N_3181);
nor U3490 (N_3490,N_3124,N_3016);
nor U3491 (N_3491,N_3225,N_3021);
nand U3492 (N_3492,N_3065,N_3241);
or U3493 (N_3493,N_3169,N_3130);
xnor U3494 (N_3494,N_3028,N_3153);
or U3495 (N_3495,N_3209,N_3053);
nand U3496 (N_3496,N_3200,N_3071);
xnor U3497 (N_3497,N_3232,N_3057);
or U3498 (N_3498,N_3024,N_3200);
nor U3499 (N_3499,N_3177,N_3110);
nor U3500 (N_3500,N_3355,N_3432);
nand U3501 (N_3501,N_3368,N_3361);
and U3502 (N_3502,N_3283,N_3378);
and U3503 (N_3503,N_3291,N_3344);
or U3504 (N_3504,N_3294,N_3350);
nand U3505 (N_3505,N_3251,N_3308);
and U3506 (N_3506,N_3440,N_3424);
and U3507 (N_3507,N_3477,N_3299);
xor U3508 (N_3508,N_3262,N_3447);
or U3509 (N_3509,N_3326,N_3281);
nor U3510 (N_3510,N_3445,N_3489);
and U3511 (N_3511,N_3254,N_3336);
or U3512 (N_3512,N_3339,N_3307);
or U3513 (N_3513,N_3453,N_3464);
nand U3514 (N_3514,N_3474,N_3498);
nand U3515 (N_3515,N_3250,N_3439);
nand U3516 (N_3516,N_3471,N_3373);
nand U3517 (N_3517,N_3412,N_3438);
xor U3518 (N_3518,N_3315,N_3332);
and U3519 (N_3519,N_3260,N_3274);
xnor U3520 (N_3520,N_3351,N_3385);
nand U3521 (N_3521,N_3257,N_3382);
nor U3522 (N_3522,N_3311,N_3414);
nand U3523 (N_3523,N_3337,N_3296);
nand U3524 (N_3524,N_3401,N_3395);
or U3525 (N_3525,N_3463,N_3347);
nor U3526 (N_3526,N_3313,N_3287);
or U3527 (N_3527,N_3425,N_3333);
or U3528 (N_3528,N_3300,N_3486);
nor U3529 (N_3529,N_3276,N_3429);
and U3530 (N_3530,N_3431,N_3420);
nand U3531 (N_3531,N_3263,N_3318);
xnor U3532 (N_3532,N_3467,N_3292);
nand U3533 (N_3533,N_3269,N_3319);
nand U3534 (N_3534,N_3383,N_3356);
or U3535 (N_3535,N_3266,N_3271);
nand U3536 (N_3536,N_3265,N_3314);
or U3537 (N_3537,N_3327,N_3341);
and U3538 (N_3538,N_3367,N_3279);
nor U3539 (N_3539,N_3436,N_3478);
nand U3540 (N_3540,N_3444,N_3258);
and U3541 (N_3541,N_3365,N_3499);
xor U3542 (N_3542,N_3446,N_3277);
and U3543 (N_3543,N_3402,N_3349);
nor U3544 (N_3544,N_3480,N_3405);
nand U3545 (N_3545,N_3305,N_3255);
and U3546 (N_3546,N_3370,N_3363);
xnor U3547 (N_3547,N_3415,N_3253);
nand U3548 (N_3548,N_3470,N_3297);
nor U3549 (N_3549,N_3304,N_3324);
and U3550 (N_3550,N_3495,N_3423);
nand U3551 (N_3551,N_3298,N_3461);
and U3552 (N_3552,N_3472,N_3309);
and U3553 (N_3553,N_3353,N_3384);
nor U3554 (N_3554,N_3290,N_3452);
and U3555 (N_3555,N_3497,N_3413);
or U3556 (N_3556,N_3375,N_3458);
or U3557 (N_3557,N_3273,N_3462);
nand U3558 (N_3558,N_3264,N_3479);
and U3559 (N_3559,N_3427,N_3342);
and U3560 (N_3560,N_3496,N_3450);
or U3561 (N_3561,N_3357,N_3302);
or U3562 (N_3562,N_3391,N_3387);
and U3563 (N_3563,N_3459,N_3451);
xnor U3564 (N_3564,N_3380,N_3312);
nor U3565 (N_3565,N_3282,N_3270);
or U3566 (N_3566,N_3389,N_3417);
nand U3567 (N_3567,N_3331,N_3485);
nand U3568 (N_3568,N_3488,N_3376);
xnor U3569 (N_3569,N_3284,N_3293);
nand U3570 (N_3570,N_3448,N_3466);
xnor U3571 (N_3571,N_3289,N_3460);
nor U3572 (N_3572,N_3483,N_3275);
or U3573 (N_3573,N_3360,N_3456);
xnor U3574 (N_3574,N_3487,N_3411);
nand U3575 (N_3575,N_3386,N_3403);
and U3576 (N_3576,N_3267,N_3381);
nor U3577 (N_3577,N_3371,N_3404);
xor U3578 (N_3578,N_3406,N_3278);
nor U3579 (N_3579,N_3388,N_3493);
and U3580 (N_3580,N_3494,N_3465);
xnor U3581 (N_3581,N_3330,N_3390);
nand U3582 (N_3582,N_3256,N_3397);
and U3583 (N_3583,N_3320,N_3329);
nand U3584 (N_3584,N_3379,N_3408);
nand U3585 (N_3585,N_3449,N_3338);
and U3586 (N_3586,N_3426,N_3377);
nand U3587 (N_3587,N_3484,N_3399);
nand U3588 (N_3588,N_3469,N_3334);
or U3589 (N_3589,N_3328,N_3435);
and U3590 (N_3590,N_3345,N_3325);
and U3591 (N_3591,N_3372,N_3354);
nor U3592 (N_3592,N_3346,N_3396);
and U3593 (N_3593,N_3321,N_3393);
and U3594 (N_3594,N_3457,N_3407);
and U3595 (N_3595,N_3316,N_3335);
or U3596 (N_3596,N_3392,N_3416);
or U3597 (N_3597,N_3482,N_3418);
and U3598 (N_3598,N_3285,N_3419);
nand U3599 (N_3599,N_3476,N_3366);
xnor U3600 (N_3600,N_3394,N_3455);
nor U3601 (N_3601,N_3428,N_3303);
xor U3602 (N_3602,N_3442,N_3410);
or U3603 (N_3603,N_3286,N_3288);
xor U3604 (N_3604,N_3369,N_3362);
or U3605 (N_3605,N_3490,N_3492);
and U3606 (N_3606,N_3261,N_3443);
and U3607 (N_3607,N_3310,N_3468);
and U3608 (N_3608,N_3343,N_3473);
or U3609 (N_3609,N_3434,N_3359);
and U3610 (N_3610,N_3340,N_3430);
nand U3611 (N_3611,N_3322,N_3374);
nor U3612 (N_3612,N_3268,N_3400);
and U3613 (N_3613,N_3280,N_3252);
or U3614 (N_3614,N_3437,N_3348);
xnor U3615 (N_3615,N_3306,N_3454);
nor U3616 (N_3616,N_3441,N_3421);
nand U3617 (N_3617,N_3481,N_3409);
and U3618 (N_3618,N_3422,N_3433);
and U3619 (N_3619,N_3323,N_3358);
nand U3620 (N_3620,N_3475,N_3364);
and U3621 (N_3621,N_3317,N_3398);
and U3622 (N_3622,N_3491,N_3301);
nand U3623 (N_3623,N_3352,N_3259);
nor U3624 (N_3624,N_3295,N_3272);
xor U3625 (N_3625,N_3378,N_3383);
and U3626 (N_3626,N_3480,N_3494);
xnor U3627 (N_3627,N_3344,N_3346);
and U3628 (N_3628,N_3407,N_3464);
nand U3629 (N_3629,N_3392,N_3413);
nor U3630 (N_3630,N_3376,N_3300);
xnor U3631 (N_3631,N_3333,N_3372);
and U3632 (N_3632,N_3361,N_3330);
and U3633 (N_3633,N_3274,N_3383);
nor U3634 (N_3634,N_3494,N_3336);
nor U3635 (N_3635,N_3498,N_3288);
or U3636 (N_3636,N_3383,N_3350);
nand U3637 (N_3637,N_3382,N_3481);
nor U3638 (N_3638,N_3379,N_3456);
nand U3639 (N_3639,N_3350,N_3384);
nor U3640 (N_3640,N_3466,N_3346);
and U3641 (N_3641,N_3270,N_3420);
or U3642 (N_3642,N_3335,N_3321);
nand U3643 (N_3643,N_3251,N_3290);
nor U3644 (N_3644,N_3390,N_3392);
xnor U3645 (N_3645,N_3373,N_3286);
nor U3646 (N_3646,N_3387,N_3372);
xnor U3647 (N_3647,N_3321,N_3368);
xnor U3648 (N_3648,N_3482,N_3289);
and U3649 (N_3649,N_3496,N_3360);
nand U3650 (N_3650,N_3347,N_3442);
nand U3651 (N_3651,N_3322,N_3345);
or U3652 (N_3652,N_3486,N_3462);
and U3653 (N_3653,N_3432,N_3284);
or U3654 (N_3654,N_3354,N_3470);
and U3655 (N_3655,N_3400,N_3316);
or U3656 (N_3656,N_3296,N_3478);
nand U3657 (N_3657,N_3312,N_3467);
nand U3658 (N_3658,N_3351,N_3313);
or U3659 (N_3659,N_3419,N_3290);
nand U3660 (N_3660,N_3327,N_3306);
and U3661 (N_3661,N_3284,N_3462);
nor U3662 (N_3662,N_3365,N_3330);
or U3663 (N_3663,N_3400,N_3330);
or U3664 (N_3664,N_3326,N_3412);
xnor U3665 (N_3665,N_3377,N_3318);
nor U3666 (N_3666,N_3308,N_3436);
nor U3667 (N_3667,N_3493,N_3326);
xnor U3668 (N_3668,N_3449,N_3272);
or U3669 (N_3669,N_3382,N_3478);
and U3670 (N_3670,N_3478,N_3404);
and U3671 (N_3671,N_3292,N_3312);
xor U3672 (N_3672,N_3423,N_3489);
nor U3673 (N_3673,N_3402,N_3335);
nor U3674 (N_3674,N_3363,N_3350);
nor U3675 (N_3675,N_3367,N_3253);
xor U3676 (N_3676,N_3401,N_3432);
nand U3677 (N_3677,N_3276,N_3383);
xor U3678 (N_3678,N_3359,N_3253);
or U3679 (N_3679,N_3258,N_3396);
nor U3680 (N_3680,N_3441,N_3381);
and U3681 (N_3681,N_3406,N_3487);
nand U3682 (N_3682,N_3380,N_3395);
and U3683 (N_3683,N_3459,N_3262);
nor U3684 (N_3684,N_3268,N_3267);
xnor U3685 (N_3685,N_3329,N_3442);
and U3686 (N_3686,N_3480,N_3495);
xor U3687 (N_3687,N_3309,N_3328);
or U3688 (N_3688,N_3266,N_3267);
nand U3689 (N_3689,N_3498,N_3263);
or U3690 (N_3690,N_3418,N_3256);
or U3691 (N_3691,N_3254,N_3433);
nor U3692 (N_3692,N_3395,N_3496);
and U3693 (N_3693,N_3458,N_3363);
xor U3694 (N_3694,N_3399,N_3498);
nand U3695 (N_3695,N_3411,N_3455);
and U3696 (N_3696,N_3496,N_3251);
and U3697 (N_3697,N_3432,N_3352);
nor U3698 (N_3698,N_3278,N_3412);
xor U3699 (N_3699,N_3417,N_3343);
nand U3700 (N_3700,N_3373,N_3495);
or U3701 (N_3701,N_3427,N_3481);
xnor U3702 (N_3702,N_3438,N_3328);
nor U3703 (N_3703,N_3276,N_3256);
or U3704 (N_3704,N_3252,N_3315);
xnor U3705 (N_3705,N_3453,N_3435);
nor U3706 (N_3706,N_3336,N_3303);
nor U3707 (N_3707,N_3275,N_3283);
or U3708 (N_3708,N_3353,N_3390);
nand U3709 (N_3709,N_3390,N_3386);
xnor U3710 (N_3710,N_3414,N_3482);
nor U3711 (N_3711,N_3256,N_3465);
nor U3712 (N_3712,N_3388,N_3301);
or U3713 (N_3713,N_3477,N_3368);
nand U3714 (N_3714,N_3491,N_3472);
and U3715 (N_3715,N_3498,N_3339);
nor U3716 (N_3716,N_3318,N_3351);
xor U3717 (N_3717,N_3299,N_3463);
and U3718 (N_3718,N_3251,N_3452);
xor U3719 (N_3719,N_3389,N_3415);
xnor U3720 (N_3720,N_3418,N_3298);
and U3721 (N_3721,N_3405,N_3287);
xor U3722 (N_3722,N_3471,N_3394);
or U3723 (N_3723,N_3492,N_3397);
and U3724 (N_3724,N_3434,N_3390);
nor U3725 (N_3725,N_3440,N_3353);
nand U3726 (N_3726,N_3250,N_3415);
nor U3727 (N_3727,N_3309,N_3491);
xnor U3728 (N_3728,N_3433,N_3286);
xor U3729 (N_3729,N_3262,N_3310);
nand U3730 (N_3730,N_3334,N_3389);
xnor U3731 (N_3731,N_3412,N_3257);
and U3732 (N_3732,N_3352,N_3262);
and U3733 (N_3733,N_3271,N_3470);
and U3734 (N_3734,N_3359,N_3439);
xor U3735 (N_3735,N_3285,N_3396);
and U3736 (N_3736,N_3475,N_3456);
nand U3737 (N_3737,N_3421,N_3449);
or U3738 (N_3738,N_3275,N_3361);
xor U3739 (N_3739,N_3341,N_3253);
or U3740 (N_3740,N_3479,N_3436);
nand U3741 (N_3741,N_3304,N_3341);
nand U3742 (N_3742,N_3344,N_3301);
and U3743 (N_3743,N_3263,N_3429);
xor U3744 (N_3744,N_3420,N_3376);
xnor U3745 (N_3745,N_3475,N_3469);
nand U3746 (N_3746,N_3368,N_3424);
xnor U3747 (N_3747,N_3292,N_3388);
xnor U3748 (N_3748,N_3279,N_3424);
nor U3749 (N_3749,N_3440,N_3435);
nor U3750 (N_3750,N_3685,N_3611);
xnor U3751 (N_3751,N_3501,N_3584);
xor U3752 (N_3752,N_3721,N_3609);
or U3753 (N_3753,N_3671,N_3698);
nor U3754 (N_3754,N_3612,N_3733);
nor U3755 (N_3755,N_3608,N_3749);
nor U3756 (N_3756,N_3617,N_3505);
nor U3757 (N_3757,N_3578,N_3666);
nor U3758 (N_3758,N_3732,N_3709);
nand U3759 (N_3759,N_3623,N_3688);
nor U3760 (N_3760,N_3618,N_3695);
and U3761 (N_3761,N_3659,N_3509);
nor U3762 (N_3762,N_3634,N_3529);
nand U3763 (N_3763,N_3678,N_3518);
or U3764 (N_3764,N_3651,N_3516);
and U3765 (N_3765,N_3726,N_3592);
and U3766 (N_3766,N_3711,N_3670);
nand U3767 (N_3767,N_3632,N_3548);
nor U3768 (N_3768,N_3504,N_3631);
nand U3769 (N_3769,N_3537,N_3664);
nand U3770 (N_3770,N_3534,N_3697);
nand U3771 (N_3771,N_3649,N_3579);
or U3772 (N_3772,N_3627,N_3638);
xnor U3773 (N_3773,N_3636,N_3644);
and U3774 (N_3774,N_3737,N_3715);
and U3775 (N_3775,N_3707,N_3563);
nand U3776 (N_3776,N_3693,N_3681);
and U3777 (N_3777,N_3589,N_3716);
xor U3778 (N_3778,N_3637,N_3720);
xnor U3779 (N_3779,N_3536,N_3561);
nand U3780 (N_3780,N_3524,N_3574);
nand U3781 (N_3781,N_3710,N_3519);
nand U3782 (N_3782,N_3729,N_3610);
xor U3783 (N_3783,N_3656,N_3541);
or U3784 (N_3784,N_3645,N_3723);
and U3785 (N_3785,N_3567,N_3547);
nor U3786 (N_3786,N_3503,N_3740);
or U3787 (N_3787,N_3582,N_3641);
nor U3788 (N_3788,N_3511,N_3619);
nand U3789 (N_3789,N_3706,N_3701);
nand U3790 (N_3790,N_3564,N_3620);
or U3791 (N_3791,N_3735,N_3602);
nand U3792 (N_3792,N_3559,N_3665);
nor U3793 (N_3793,N_3662,N_3731);
xnor U3794 (N_3794,N_3590,N_3722);
or U3795 (N_3795,N_3633,N_3672);
and U3796 (N_3796,N_3521,N_3531);
xor U3797 (N_3797,N_3585,N_3580);
or U3798 (N_3798,N_3552,N_3684);
and U3799 (N_3799,N_3725,N_3605);
and U3800 (N_3800,N_3570,N_3679);
or U3801 (N_3801,N_3667,N_3680);
xnor U3802 (N_3802,N_3593,N_3745);
and U3803 (N_3803,N_3703,N_3748);
nor U3804 (N_3804,N_3522,N_3639);
nand U3805 (N_3805,N_3513,N_3557);
or U3806 (N_3806,N_3507,N_3560);
nand U3807 (N_3807,N_3538,N_3738);
nor U3808 (N_3808,N_3652,N_3646);
and U3809 (N_3809,N_3586,N_3601);
xor U3810 (N_3810,N_3626,N_3699);
or U3811 (N_3811,N_3571,N_3588);
nor U3812 (N_3812,N_3500,N_3525);
xor U3813 (N_3813,N_3654,N_3515);
and U3814 (N_3814,N_3746,N_3643);
or U3815 (N_3815,N_3668,N_3742);
nand U3816 (N_3816,N_3717,N_3677);
nand U3817 (N_3817,N_3714,N_3724);
or U3818 (N_3818,N_3628,N_3675);
nor U3819 (N_3819,N_3747,N_3517);
nand U3820 (N_3820,N_3520,N_3676);
nand U3821 (N_3821,N_3708,N_3658);
xor U3822 (N_3822,N_3514,N_3566);
and U3823 (N_3823,N_3527,N_3744);
nor U3824 (N_3824,N_3572,N_3663);
nand U3825 (N_3825,N_3562,N_3583);
and U3826 (N_3826,N_3647,N_3568);
and U3827 (N_3827,N_3549,N_3615);
and U3828 (N_3828,N_3545,N_3630);
or U3829 (N_3829,N_3616,N_3719);
or U3830 (N_3830,N_3535,N_3607);
and U3831 (N_3831,N_3542,N_3606);
xnor U3832 (N_3832,N_3543,N_3603);
nor U3833 (N_3833,N_3621,N_3591);
nand U3834 (N_3834,N_3624,N_3739);
nor U3835 (N_3835,N_3712,N_3506);
nor U3836 (N_3836,N_3650,N_3625);
nand U3837 (N_3837,N_3532,N_3508);
and U3838 (N_3838,N_3727,N_3598);
nor U3839 (N_3839,N_3730,N_3686);
xnor U3840 (N_3840,N_3648,N_3596);
or U3841 (N_3841,N_3687,N_3673);
xnor U3842 (N_3842,N_3526,N_3704);
xnor U3843 (N_3843,N_3683,N_3700);
xnor U3844 (N_3844,N_3657,N_3594);
or U3845 (N_3845,N_3551,N_3736);
nor U3846 (N_3846,N_3705,N_3622);
nor U3847 (N_3847,N_3573,N_3692);
nand U3848 (N_3848,N_3661,N_3595);
nand U3849 (N_3849,N_3682,N_3597);
nor U3850 (N_3850,N_3523,N_3604);
nand U3851 (N_3851,N_3556,N_3614);
nand U3852 (N_3852,N_3533,N_3635);
xnor U3853 (N_3853,N_3528,N_3530);
nand U3854 (N_3854,N_3669,N_3553);
xor U3855 (N_3855,N_3576,N_3581);
xnor U3856 (N_3856,N_3743,N_3696);
and U3857 (N_3857,N_3629,N_3558);
xor U3858 (N_3858,N_3539,N_3540);
nand U3859 (N_3859,N_3689,N_3655);
xor U3860 (N_3860,N_3599,N_3550);
nand U3861 (N_3861,N_3613,N_3728);
nor U3862 (N_3862,N_3702,N_3569);
nand U3863 (N_3863,N_3555,N_3674);
or U3864 (N_3864,N_3713,N_3642);
nand U3865 (N_3865,N_3734,N_3544);
or U3866 (N_3866,N_3546,N_3718);
or U3867 (N_3867,N_3512,N_3653);
or U3868 (N_3868,N_3600,N_3640);
nand U3869 (N_3869,N_3502,N_3694);
xor U3870 (N_3870,N_3660,N_3691);
or U3871 (N_3871,N_3510,N_3565);
nor U3872 (N_3872,N_3587,N_3575);
nor U3873 (N_3873,N_3554,N_3690);
nor U3874 (N_3874,N_3577,N_3741);
and U3875 (N_3875,N_3745,N_3517);
nor U3876 (N_3876,N_3636,N_3630);
nand U3877 (N_3877,N_3633,N_3735);
and U3878 (N_3878,N_3674,N_3690);
and U3879 (N_3879,N_3525,N_3609);
nand U3880 (N_3880,N_3504,N_3547);
nor U3881 (N_3881,N_3703,N_3606);
xor U3882 (N_3882,N_3641,N_3561);
xnor U3883 (N_3883,N_3693,N_3651);
nor U3884 (N_3884,N_3613,N_3524);
nand U3885 (N_3885,N_3671,N_3654);
nor U3886 (N_3886,N_3506,N_3552);
xnor U3887 (N_3887,N_3718,N_3502);
nand U3888 (N_3888,N_3607,N_3739);
or U3889 (N_3889,N_3645,N_3572);
and U3890 (N_3890,N_3667,N_3656);
nand U3891 (N_3891,N_3501,N_3546);
nand U3892 (N_3892,N_3527,N_3528);
and U3893 (N_3893,N_3570,N_3704);
or U3894 (N_3894,N_3655,N_3685);
nand U3895 (N_3895,N_3690,N_3669);
and U3896 (N_3896,N_3649,N_3705);
nor U3897 (N_3897,N_3725,N_3571);
xor U3898 (N_3898,N_3657,N_3587);
nand U3899 (N_3899,N_3559,N_3610);
nor U3900 (N_3900,N_3694,N_3545);
and U3901 (N_3901,N_3562,N_3642);
or U3902 (N_3902,N_3577,N_3605);
nand U3903 (N_3903,N_3660,N_3613);
xnor U3904 (N_3904,N_3733,N_3718);
and U3905 (N_3905,N_3697,N_3613);
and U3906 (N_3906,N_3536,N_3717);
and U3907 (N_3907,N_3684,N_3605);
nor U3908 (N_3908,N_3582,N_3654);
and U3909 (N_3909,N_3706,N_3608);
or U3910 (N_3910,N_3622,N_3665);
and U3911 (N_3911,N_3621,N_3647);
and U3912 (N_3912,N_3556,N_3733);
or U3913 (N_3913,N_3669,N_3748);
nor U3914 (N_3914,N_3534,N_3574);
or U3915 (N_3915,N_3504,N_3619);
nor U3916 (N_3916,N_3625,N_3579);
or U3917 (N_3917,N_3591,N_3570);
nor U3918 (N_3918,N_3539,N_3614);
xnor U3919 (N_3919,N_3600,N_3611);
xnor U3920 (N_3920,N_3685,N_3669);
xor U3921 (N_3921,N_3607,N_3745);
or U3922 (N_3922,N_3559,N_3554);
xnor U3923 (N_3923,N_3692,N_3554);
nor U3924 (N_3924,N_3509,N_3517);
nor U3925 (N_3925,N_3528,N_3645);
xor U3926 (N_3926,N_3685,N_3734);
nand U3927 (N_3927,N_3581,N_3554);
nor U3928 (N_3928,N_3687,N_3524);
nor U3929 (N_3929,N_3562,N_3545);
xor U3930 (N_3930,N_3509,N_3648);
xnor U3931 (N_3931,N_3598,N_3738);
and U3932 (N_3932,N_3523,N_3503);
or U3933 (N_3933,N_3522,N_3620);
xor U3934 (N_3934,N_3634,N_3695);
nor U3935 (N_3935,N_3514,N_3576);
and U3936 (N_3936,N_3657,N_3533);
xor U3937 (N_3937,N_3673,N_3667);
nor U3938 (N_3938,N_3563,N_3617);
xor U3939 (N_3939,N_3717,N_3636);
nor U3940 (N_3940,N_3693,N_3695);
nand U3941 (N_3941,N_3693,N_3701);
or U3942 (N_3942,N_3629,N_3638);
xor U3943 (N_3943,N_3617,N_3561);
or U3944 (N_3944,N_3661,N_3601);
and U3945 (N_3945,N_3720,N_3516);
nor U3946 (N_3946,N_3676,N_3625);
and U3947 (N_3947,N_3667,N_3548);
and U3948 (N_3948,N_3580,N_3637);
or U3949 (N_3949,N_3578,N_3598);
or U3950 (N_3950,N_3681,N_3515);
and U3951 (N_3951,N_3630,N_3622);
xor U3952 (N_3952,N_3657,N_3670);
nand U3953 (N_3953,N_3571,N_3520);
or U3954 (N_3954,N_3592,N_3589);
nor U3955 (N_3955,N_3643,N_3514);
nand U3956 (N_3956,N_3546,N_3547);
or U3957 (N_3957,N_3705,N_3730);
nor U3958 (N_3958,N_3687,N_3515);
or U3959 (N_3959,N_3517,N_3531);
xor U3960 (N_3960,N_3661,N_3549);
xnor U3961 (N_3961,N_3665,N_3627);
nor U3962 (N_3962,N_3625,N_3541);
or U3963 (N_3963,N_3524,N_3632);
or U3964 (N_3964,N_3690,N_3640);
nand U3965 (N_3965,N_3625,N_3538);
and U3966 (N_3966,N_3612,N_3629);
nand U3967 (N_3967,N_3604,N_3710);
xor U3968 (N_3968,N_3553,N_3717);
or U3969 (N_3969,N_3654,N_3559);
and U3970 (N_3970,N_3611,N_3578);
xnor U3971 (N_3971,N_3551,N_3694);
and U3972 (N_3972,N_3660,N_3536);
xnor U3973 (N_3973,N_3651,N_3625);
nor U3974 (N_3974,N_3675,N_3571);
nor U3975 (N_3975,N_3678,N_3708);
nand U3976 (N_3976,N_3514,N_3730);
nand U3977 (N_3977,N_3675,N_3594);
or U3978 (N_3978,N_3539,N_3558);
nor U3979 (N_3979,N_3542,N_3706);
nand U3980 (N_3980,N_3730,N_3510);
nor U3981 (N_3981,N_3706,N_3636);
and U3982 (N_3982,N_3510,N_3710);
or U3983 (N_3983,N_3560,N_3669);
nand U3984 (N_3984,N_3588,N_3597);
nor U3985 (N_3985,N_3642,N_3578);
and U3986 (N_3986,N_3737,N_3695);
nor U3987 (N_3987,N_3521,N_3747);
xor U3988 (N_3988,N_3712,N_3736);
nor U3989 (N_3989,N_3539,N_3646);
nand U3990 (N_3990,N_3576,N_3569);
or U3991 (N_3991,N_3511,N_3671);
nand U3992 (N_3992,N_3593,N_3535);
nand U3993 (N_3993,N_3544,N_3599);
and U3994 (N_3994,N_3613,N_3584);
xnor U3995 (N_3995,N_3597,N_3642);
nand U3996 (N_3996,N_3620,N_3669);
or U3997 (N_3997,N_3705,N_3522);
or U3998 (N_3998,N_3567,N_3626);
xor U3999 (N_3999,N_3747,N_3727);
nor U4000 (N_4000,N_3977,N_3961);
nor U4001 (N_4001,N_3768,N_3985);
xor U4002 (N_4002,N_3852,N_3923);
xor U4003 (N_4003,N_3878,N_3998);
xnor U4004 (N_4004,N_3834,N_3838);
xor U4005 (N_4005,N_3787,N_3924);
nand U4006 (N_4006,N_3771,N_3839);
and U4007 (N_4007,N_3916,N_3811);
or U4008 (N_4008,N_3910,N_3782);
or U4009 (N_4009,N_3992,N_3821);
nand U4010 (N_4010,N_3769,N_3765);
nor U4011 (N_4011,N_3796,N_3883);
nor U4012 (N_4012,N_3843,N_3766);
xnor U4013 (N_4013,N_3802,N_3779);
or U4014 (N_4014,N_3778,N_3988);
and U4015 (N_4015,N_3812,N_3795);
nand U4016 (N_4016,N_3845,N_3814);
nor U4017 (N_4017,N_3897,N_3900);
and U4018 (N_4018,N_3783,N_3776);
or U4019 (N_4019,N_3790,N_3848);
and U4020 (N_4020,N_3904,N_3996);
or U4021 (N_4021,N_3939,N_3835);
and U4022 (N_4022,N_3840,N_3865);
nand U4023 (N_4023,N_3946,N_3829);
or U4024 (N_4024,N_3938,N_3793);
xnor U4025 (N_4025,N_3979,N_3945);
xor U4026 (N_4026,N_3906,N_3804);
or U4027 (N_4027,N_3826,N_3911);
nand U4028 (N_4028,N_3944,N_3841);
nand U4029 (N_4029,N_3907,N_3857);
and U4030 (N_4030,N_3917,N_3750);
nor U4031 (N_4031,N_3993,N_3899);
xnor U4032 (N_4032,N_3858,N_3866);
nor U4033 (N_4033,N_3958,N_3886);
nand U4034 (N_4034,N_3825,N_3764);
or U4035 (N_4035,N_3797,N_3850);
or U4036 (N_4036,N_3894,N_3934);
nand U4037 (N_4037,N_3752,N_3922);
or U4038 (N_4038,N_3891,N_3846);
nor U4039 (N_4039,N_3849,N_3994);
and U4040 (N_4040,N_3855,N_3966);
and U4041 (N_4041,N_3935,N_3827);
xnor U4042 (N_4042,N_3931,N_3833);
nand U4043 (N_4043,N_3959,N_3819);
nor U4044 (N_4044,N_3963,N_3936);
or U4045 (N_4045,N_3862,N_3842);
and U4046 (N_4046,N_3785,N_3892);
nand U4047 (N_4047,N_3851,N_3844);
and U4048 (N_4048,N_3759,N_3962);
and U4049 (N_4049,N_3948,N_3805);
or U4050 (N_4050,N_3763,N_3896);
xor U4051 (N_4051,N_3880,N_3755);
xor U4052 (N_4052,N_3960,N_3984);
and U4053 (N_4053,N_3953,N_3928);
nand U4054 (N_4054,N_3895,N_3952);
and U4055 (N_4055,N_3786,N_3893);
nand U4056 (N_4056,N_3915,N_3762);
nor U4057 (N_4057,N_3818,N_3887);
and U4058 (N_4058,N_3942,N_3918);
nor U4059 (N_4059,N_3903,N_3999);
or U4060 (N_4060,N_3968,N_3919);
or U4061 (N_4061,N_3940,N_3986);
or U4062 (N_4062,N_3920,N_3908);
nand U4063 (N_4063,N_3863,N_3973);
or U4064 (N_4064,N_3773,N_3974);
xnor U4065 (N_4065,N_3875,N_3753);
nand U4066 (N_4066,N_3925,N_3800);
or U4067 (N_4067,N_3969,N_3861);
or U4068 (N_4068,N_3751,N_3912);
nor U4069 (N_4069,N_3921,N_3820);
and U4070 (N_4070,N_3777,N_3799);
xnor U4071 (N_4071,N_3997,N_3815);
xor U4072 (N_4072,N_3975,N_3930);
xnor U4073 (N_4073,N_3830,N_3901);
or U4074 (N_4074,N_3964,N_3980);
nor U4075 (N_4075,N_3956,N_3869);
or U4076 (N_4076,N_3831,N_3864);
nand U4077 (N_4077,N_3913,N_3954);
or U4078 (N_4078,N_3853,N_3832);
nor U4079 (N_4079,N_3767,N_3784);
nand U4080 (N_4080,N_3976,N_3837);
and U4081 (N_4081,N_3972,N_3882);
or U4082 (N_4082,N_3859,N_3932);
and U4083 (N_4083,N_3775,N_3788);
nor U4084 (N_4084,N_3951,N_3965);
nor U4085 (N_4085,N_3889,N_3909);
nor U4086 (N_4086,N_3879,N_3868);
xnor U4087 (N_4087,N_3967,N_3824);
and U4088 (N_4088,N_3890,N_3823);
nand U4089 (N_4089,N_3983,N_3789);
xor U4090 (N_4090,N_3822,N_3981);
or U4091 (N_4091,N_3754,N_3885);
nor U4092 (N_4092,N_3806,N_3949);
and U4093 (N_4093,N_3808,N_3876);
or U4094 (N_4094,N_3854,N_3933);
nand U4095 (N_4095,N_3982,N_3888);
or U4096 (N_4096,N_3860,N_3794);
nor U4097 (N_4097,N_3877,N_3770);
or U4098 (N_4098,N_3757,N_3809);
and U4099 (N_4099,N_3873,N_3943);
xor U4100 (N_4100,N_3991,N_3937);
nor U4101 (N_4101,N_3871,N_3929);
xor U4102 (N_4102,N_3947,N_3872);
nor U4103 (N_4103,N_3971,N_3989);
xor U4104 (N_4104,N_3898,N_3791);
and U4105 (N_4105,N_3798,N_3902);
or U4106 (N_4106,N_3970,N_3870);
or U4107 (N_4107,N_3810,N_3758);
or U4108 (N_4108,N_3817,N_3836);
xor U4109 (N_4109,N_3828,N_3856);
nor U4110 (N_4110,N_3760,N_3990);
nand U4111 (N_4111,N_3995,N_3761);
xor U4112 (N_4112,N_3950,N_3884);
nand U4113 (N_4113,N_3941,N_3927);
nor U4114 (N_4114,N_3780,N_3781);
and U4115 (N_4115,N_3847,N_3774);
nor U4116 (N_4116,N_3955,N_3813);
xor U4117 (N_4117,N_3816,N_3987);
and U4118 (N_4118,N_3926,N_3874);
nand U4119 (N_4119,N_3792,N_3756);
and U4120 (N_4120,N_3807,N_3881);
and U4121 (N_4121,N_3914,N_3867);
nand U4122 (N_4122,N_3978,N_3905);
nor U4123 (N_4123,N_3957,N_3772);
xor U4124 (N_4124,N_3801,N_3803);
or U4125 (N_4125,N_3846,N_3911);
nand U4126 (N_4126,N_3890,N_3780);
or U4127 (N_4127,N_3977,N_3754);
and U4128 (N_4128,N_3982,N_3812);
or U4129 (N_4129,N_3879,N_3839);
and U4130 (N_4130,N_3954,N_3930);
xor U4131 (N_4131,N_3765,N_3902);
or U4132 (N_4132,N_3782,N_3792);
or U4133 (N_4133,N_3872,N_3927);
nor U4134 (N_4134,N_3752,N_3977);
nor U4135 (N_4135,N_3896,N_3887);
nor U4136 (N_4136,N_3754,N_3937);
xnor U4137 (N_4137,N_3946,N_3995);
or U4138 (N_4138,N_3847,N_3814);
nor U4139 (N_4139,N_3750,N_3815);
or U4140 (N_4140,N_3781,N_3824);
xor U4141 (N_4141,N_3804,N_3963);
and U4142 (N_4142,N_3801,N_3894);
xor U4143 (N_4143,N_3922,N_3994);
nor U4144 (N_4144,N_3926,N_3950);
nand U4145 (N_4145,N_3849,N_3764);
nand U4146 (N_4146,N_3866,N_3750);
and U4147 (N_4147,N_3829,N_3792);
nand U4148 (N_4148,N_3931,N_3821);
nor U4149 (N_4149,N_3824,N_3994);
xor U4150 (N_4150,N_3832,N_3973);
or U4151 (N_4151,N_3941,N_3946);
and U4152 (N_4152,N_3979,N_3835);
xnor U4153 (N_4153,N_3787,N_3993);
and U4154 (N_4154,N_3940,N_3762);
or U4155 (N_4155,N_3888,N_3824);
xnor U4156 (N_4156,N_3801,N_3909);
or U4157 (N_4157,N_3812,N_3797);
or U4158 (N_4158,N_3869,N_3855);
xor U4159 (N_4159,N_3836,N_3938);
xnor U4160 (N_4160,N_3879,N_3836);
or U4161 (N_4161,N_3961,N_3823);
or U4162 (N_4162,N_3998,N_3967);
and U4163 (N_4163,N_3945,N_3929);
or U4164 (N_4164,N_3979,N_3843);
xnor U4165 (N_4165,N_3878,N_3925);
nand U4166 (N_4166,N_3891,N_3929);
nor U4167 (N_4167,N_3758,N_3840);
and U4168 (N_4168,N_3846,N_3984);
or U4169 (N_4169,N_3974,N_3765);
or U4170 (N_4170,N_3813,N_3913);
nor U4171 (N_4171,N_3911,N_3960);
xnor U4172 (N_4172,N_3830,N_3754);
xnor U4173 (N_4173,N_3811,N_3976);
nor U4174 (N_4174,N_3916,N_3859);
nand U4175 (N_4175,N_3898,N_3892);
and U4176 (N_4176,N_3915,N_3848);
and U4177 (N_4177,N_3754,N_3911);
nor U4178 (N_4178,N_3844,N_3999);
nand U4179 (N_4179,N_3860,N_3864);
and U4180 (N_4180,N_3956,N_3789);
or U4181 (N_4181,N_3782,N_3767);
or U4182 (N_4182,N_3759,N_3978);
and U4183 (N_4183,N_3879,N_3913);
xnor U4184 (N_4184,N_3801,N_3979);
or U4185 (N_4185,N_3955,N_3928);
and U4186 (N_4186,N_3818,N_3793);
nor U4187 (N_4187,N_3828,N_3925);
nand U4188 (N_4188,N_3849,N_3845);
nor U4189 (N_4189,N_3933,N_3800);
xor U4190 (N_4190,N_3965,N_3847);
xnor U4191 (N_4191,N_3938,N_3873);
nand U4192 (N_4192,N_3820,N_3914);
or U4193 (N_4193,N_3950,N_3991);
and U4194 (N_4194,N_3865,N_3943);
nand U4195 (N_4195,N_3785,N_3762);
and U4196 (N_4196,N_3875,N_3918);
xnor U4197 (N_4197,N_3910,N_3948);
nor U4198 (N_4198,N_3879,N_3896);
and U4199 (N_4199,N_3959,N_3971);
xor U4200 (N_4200,N_3815,N_3926);
nand U4201 (N_4201,N_3950,N_3988);
or U4202 (N_4202,N_3916,N_3882);
or U4203 (N_4203,N_3790,N_3776);
and U4204 (N_4204,N_3851,N_3843);
and U4205 (N_4205,N_3763,N_3982);
or U4206 (N_4206,N_3852,N_3996);
and U4207 (N_4207,N_3905,N_3980);
nor U4208 (N_4208,N_3893,N_3984);
xnor U4209 (N_4209,N_3832,N_3829);
or U4210 (N_4210,N_3904,N_3847);
nor U4211 (N_4211,N_3896,N_3823);
nor U4212 (N_4212,N_3776,N_3822);
nand U4213 (N_4213,N_3870,N_3945);
nor U4214 (N_4214,N_3887,N_3875);
nor U4215 (N_4215,N_3794,N_3841);
xor U4216 (N_4216,N_3849,N_3827);
or U4217 (N_4217,N_3878,N_3971);
and U4218 (N_4218,N_3907,N_3919);
nor U4219 (N_4219,N_3842,N_3889);
xor U4220 (N_4220,N_3889,N_3989);
or U4221 (N_4221,N_3785,N_3965);
xor U4222 (N_4222,N_3839,N_3893);
nand U4223 (N_4223,N_3780,N_3803);
xor U4224 (N_4224,N_3759,N_3795);
xor U4225 (N_4225,N_3976,N_3826);
nor U4226 (N_4226,N_3862,N_3915);
and U4227 (N_4227,N_3920,N_3756);
nor U4228 (N_4228,N_3767,N_3822);
or U4229 (N_4229,N_3750,N_3895);
nand U4230 (N_4230,N_3907,N_3793);
xnor U4231 (N_4231,N_3840,N_3790);
nor U4232 (N_4232,N_3870,N_3779);
xor U4233 (N_4233,N_3891,N_3918);
or U4234 (N_4234,N_3973,N_3981);
xnor U4235 (N_4235,N_3812,N_3752);
and U4236 (N_4236,N_3899,N_3793);
nor U4237 (N_4237,N_3892,N_3890);
or U4238 (N_4238,N_3812,N_3833);
and U4239 (N_4239,N_3995,N_3899);
and U4240 (N_4240,N_3988,N_3932);
and U4241 (N_4241,N_3824,N_3974);
and U4242 (N_4242,N_3750,N_3814);
nand U4243 (N_4243,N_3814,N_3978);
nand U4244 (N_4244,N_3780,N_3985);
xnor U4245 (N_4245,N_3750,N_3766);
xnor U4246 (N_4246,N_3903,N_3941);
nor U4247 (N_4247,N_3912,N_3902);
and U4248 (N_4248,N_3937,N_3843);
or U4249 (N_4249,N_3977,N_3878);
nor U4250 (N_4250,N_4027,N_4029);
nand U4251 (N_4251,N_4216,N_4016);
nor U4252 (N_4252,N_4189,N_4075);
nor U4253 (N_4253,N_4170,N_4060);
xor U4254 (N_4254,N_4091,N_4121);
and U4255 (N_4255,N_4167,N_4102);
or U4256 (N_4256,N_4058,N_4095);
or U4257 (N_4257,N_4061,N_4206);
and U4258 (N_4258,N_4153,N_4071);
or U4259 (N_4259,N_4145,N_4136);
nor U4260 (N_4260,N_4238,N_4147);
and U4261 (N_4261,N_4126,N_4118);
xnor U4262 (N_4262,N_4059,N_4222);
or U4263 (N_4263,N_4096,N_4213);
or U4264 (N_4264,N_4179,N_4092);
xnor U4265 (N_4265,N_4039,N_4152);
nand U4266 (N_4266,N_4001,N_4119);
nor U4267 (N_4267,N_4233,N_4084);
nand U4268 (N_4268,N_4127,N_4031);
and U4269 (N_4269,N_4134,N_4020);
and U4270 (N_4270,N_4174,N_4228);
or U4271 (N_4271,N_4181,N_4205);
and U4272 (N_4272,N_4176,N_4011);
or U4273 (N_4273,N_4028,N_4239);
nor U4274 (N_4274,N_4115,N_4249);
and U4275 (N_4275,N_4040,N_4108);
or U4276 (N_4276,N_4191,N_4101);
nand U4277 (N_4277,N_4246,N_4122);
nor U4278 (N_4278,N_4229,N_4244);
xnor U4279 (N_4279,N_4225,N_4094);
nor U4280 (N_4280,N_4187,N_4175);
and U4281 (N_4281,N_4237,N_4166);
or U4282 (N_4282,N_4182,N_4073);
or U4283 (N_4283,N_4074,N_4018);
and U4284 (N_4284,N_4218,N_4232);
nand U4285 (N_4285,N_4105,N_4009);
nor U4286 (N_4286,N_4143,N_4034);
or U4287 (N_4287,N_4100,N_4186);
and U4288 (N_4288,N_4211,N_4087);
nor U4289 (N_4289,N_4159,N_4109);
nand U4290 (N_4290,N_4204,N_4188);
nand U4291 (N_4291,N_4046,N_4043);
nand U4292 (N_4292,N_4190,N_4000);
and U4293 (N_4293,N_4064,N_4215);
nor U4294 (N_4294,N_4066,N_4088);
nand U4295 (N_4295,N_4098,N_4002);
and U4296 (N_4296,N_4192,N_4015);
and U4297 (N_4297,N_4234,N_4163);
xnor U4298 (N_4298,N_4055,N_4199);
nand U4299 (N_4299,N_4132,N_4014);
xnor U4300 (N_4300,N_4086,N_4035);
or U4301 (N_4301,N_4097,N_4005);
nand U4302 (N_4302,N_4128,N_4135);
xor U4303 (N_4303,N_4236,N_4223);
and U4304 (N_4304,N_4248,N_4082);
xnor U4305 (N_4305,N_4053,N_4036);
and U4306 (N_4306,N_4154,N_4090);
nor U4307 (N_4307,N_4026,N_4124);
xor U4308 (N_4308,N_4150,N_4070);
or U4309 (N_4309,N_4183,N_4054);
nand U4310 (N_4310,N_4010,N_4019);
and U4311 (N_4311,N_4072,N_4169);
nor U4312 (N_4312,N_4042,N_4068);
nand U4313 (N_4313,N_4220,N_4133);
nand U4314 (N_4314,N_4139,N_4138);
nand U4315 (N_4315,N_4079,N_4045);
nor U4316 (N_4316,N_4103,N_4080);
nor U4317 (N_4317,N_4196,N_4117);
nand U4318 (N_4318,N_4243,N_4226);
or U4319 (N_4319,N_4208,N_4202);
or U4320 (N_4320,N_4231,N_4038);
xnor U4321 (N_4321,N_4116,N_4160);
or U4322 (N_4322,N_4203,N_4207);
and U4323 (N_4323,N_4173,N_4024);
or U4324 (N_4324,N_4155,N_4217);
or U4325 (N_4325,N_4111,N_4164);
or U4326 (N_4326,N_4230,N_4104);
nor U4327 (N_4327,N_4149,N_4065);
xor U4328 (N_4328,N_4047,N_4180);
xnor U4329 (N_4329,N_4006,N_4227);
or U4330 (N_4330,N_4242,N_4235);
xnor U4331 (N_4331,N_4157,N_4200);
and U4332 (N_4332,N_4158,N_4184);
xor U4333 (N_4333,N_4113,N_4161);
nand U4334 (N_4334,N_4131,N_4067);
xnor U4335 (N_4335,N_4221,N_4051);
or U4336 (N_4336,N_4032,N_4037);
xor U4337 (N_4337,N_4156,N_4168);
nand U4338 (N_4338,N_4089,N_4052);
or U4339 (N_4339,N_4165,N_4195);
nand U4340 (N_4340,N_4114,N_4146);
nand U4341 (N_4341,N_4081,N_4044);
and U4342 (N_4342,N_4178,N_4110);
xnor U4343 (N_4343,N_4030,N_4201);
and U4344 (N_4344,N_4224,N_4106);
and U4345 (N_4345,N_4214,N_4093);
nor U4346 (N_4346,N_4099,N_4025);
and U4347 (N_4347,N_4172,N_4033);
nor U4348 (N_4348,N_4197,N_4137);
nor U4349 (N_4349,N_4023,N_4012);
nor U4350 (N_4350,N_4007,N_4241);
nor U4351 (N_4351,N_4129,N_4247);
and U4352 (N_4352,N_4008,N_4085);
xnor U4353 (N_4353,N_4198,N_4050);
nand U4354 (N_4354,N_4077,N_4140);
or U4355 (N_4355,N_4076,N_4107);
nor U4356 (N_4356,N_4078,N_4013);
nor U4357 (N_4357,N_4062,N_4022);
and U4358 (N_4358,N_4057,N_4240);
nor U4359 (N_4359,N_4063,N_4083);
and U4360 (N_4360,N_4120,N_4049);
or U4361 (N_4361,N_4017,N_4162);
xnor U4362 (N_4362,N_4209,N_4056);
nor U4363 (N_4363,N_4151,N_4003);
xor U4364 (N_4364,N_4123,N_4219);
and U4365 (N_4365,N_4193,N_4004);
nor U4366 (N_4366,N_4048,N_4142);
nor U4367 (N_4367,N_4112,N_4177);
nor U4368 (N_4368,N_4125,N_4130);
xor U4369 (N_4369,N_4141,N_4212);
nand U4370 (N_4370,N_4041,N_4148);
and U4371 (N_4371,N_4194,N_4245);
nand U4372 (N_4372,N_4171,N_4069);
or U4373 (N_4373,N_4144,N_4210);
and U4374 (N_4374,N_4021,N_4185);
or U4375 (N_4375,N_4118,N_4179);
and U4376 (N_4376,N_4218,N_4031);
xnor U4377 (N_4377,N_4092,N_4077);
nor U4378 (N_4378,N_4032,N_4150);
xnor U4379 (N_4379,N_4116,N_4094);
nor U4380 (N_4380,N_4090,N_4078);
and U4381 (N_4381,N_4161,N_4041);
or U4382 (N_4382,N_4087,N_4050);
nor U4383 (N_4383,N_4056,N_4131);
and U4384 (N_4384,N_4145,N_4119);
and U4385 (N_4385,N_4068,N_4145);
xnor U4386 (N_4386,N_4138,N_4151);
and U4387 (N_4387,N_4145,N_4183);
or U4388 (N_4388,N_4099,N_4194);
nor U4389 (N_4389,N_4148,N_4237);
xnor U4390 (N_4390,N_4127,N_4115);
or U4391 (N_4391,N_4245,N_4136);
or U4392 (N_4392,N_4208,N_4088);
or U4393 (N_4393,N_4221,N_4042);
nand U4394 (N_4394,N_4234,N_4016);
nand U4395 (N_4395,N_4008,N_4080);
xor U4396 (N_4396,N_4102,N_4067);
nand U4397 (N_4397,N_4105,N_4212);
xor U4398 (N_4398,N_4218,N_4052);
and U4399 (N_4399,N_4110,N_4047);
xnor U4400 (N_4400,N_4069,N_4223);
xnor U4401 (N_4401,N_4217,N_4176);
and U4402 (N_4402,N_4159,N_4213);
xnor U4403 (N_4403,N_4138,N_4176);
and U4404 (N_4404,N_4001,N_4162);
and U4405 (N_4405,N_4145,N_4231);
nor U4406 (N_4406,N_4156,N_4058);
or U4407 (N_4407,N_4112,N_4170);
xor U4408 (N_4408,N_4238,N_4172);
xnor U4409 (N_4409,N_4162,N_4249);
or U4410 (N_4410,N_4066,N_4044);
nor U4411 (N_4411,N_4249,N_4125);
nand U4412 (N_4412,N_4188,N_4178);
nand U4413 (N_4413,N_4148,N_4223);
nand U4414 (N_4414,N_4240,N_4110);
nor U4415 (N_4415,N_4175,N_4044);
and U4416 (N_4416,N_4181,N_4097);
nor U4417 (N_4417,N_4207,N_4169);
nor U4418 (N_4418,N_4023,N_4040);
nand U4419 (N_4419,N_4193,N_4175);
nor U4420 (N_4420,N_4189,N_4138);
nor U4421 (N_4421,N_4097,N_4146);
and U4422 (N_4422,N_4131,N_4124);
or U4423 (N_4423,N_4075,N_4078);
nand U4424 (N_4424,N_4155,N_4038);
or U4425 (N_4425,N_4144,N_4082);
nand U4426 (N_4426,N_4043,N_4012);
and U4427 (N_4427,N_4217,N_4207);
and U4428 (N_4428,N_4130,N_4174);
and U4429 (N_4429,N_4061,N_4142);
nand U4430 (N_4430,N_4060,N_4000);
nand U4431 (N_4431,N_4232,N_4004);
nor U4432 (N_4432,N_4124,N_4057);
nor U4433 (N_4433,N_4088,N_4148);
nor U4434 (N_4434,N_4134,N_4206);
xnor U4435 (N_4435,N_4010,N_4138);
or U4436 (N_4436,N_4206,N_4198);
or U4437 (N_4437,N_4244,N_4141);
or U4438 (N_4438,N_4050,N_4047);
and U4439 (N_4439,N_4236,N_4148);
nor U4440 (N_4440,N_4067,N_4063);
xnor U4441 (N_4441,N_4090,N_4202);
nand U4442 (N_4442,N_4013,N_4154);
nor U4443 (N_4443,N_4025,N_4095);
xor U4444 (N_4444,N_4157,N_4068);
or U4445 (N_4445,N_4175,N_4176);
nand U4446 (N_4446,N_4151,N_4154);
and U4447 (N_4447,N_4103,N_4057);
xnor U4448 (N_4448,N_4050,N_4076);
or U4449 (N_4449,N_4136,N_4104);
and U4450 (N_4450,N_4019,N_4072);
xor U4451 (N_4451,N_4244,N_4078);
xnor U4452 (N_4452,N_4099,N_4122);
and U4453 (N_4453,N_4064,N_4074);
and U4454 (N_4454,N_4212,N_4168);
nand U4455 (N_4455,N_4150,N_4046);
or U4456 (N_4456,N_4173,N_4153);
nor U4457 (N_4457,N_4047,N_4031);
and U4458 (N_4458,N_4092,N_4111);
or U4459 (N_4459,N_4041,N_4111);
or U4460 (N_4460,N_4106,N_4171);
xor U4461 (N_4461,N_4171,N_4132);
nor U4462 (N_4462,N_4172,N_4008);
nand U4463 (N_4463,N_4157,N_4029);
and U4464 (N_4464,N_4108,N_4197);
xnor U4465 (N_4465,N_4211,N_4214);
nand U4466 (N_4466,N_4029,N_4218);
or U4467 (N_4467,N_4070,N_4097);
xor U4468 (N_4468,N_4111,N_4038);
and U4469 (N_4469,N_4228,N_4055);
nand U4470 (N_4470,N_4131,N_4104);
xnor U4471 (N_4471,N_4221,N_4096);
nand U4472 (N_4472,N_4217,N_4215);
and U4473 (N_4473,N_4171,N_4092);
nand U4474 (N_4474,N_4180,N_4128);
xnor U4475 (N_4475,N_4152,N_4147);
and U4476 (N_4476,N_4136,N_4072);
or U4477 (N_4477,N_4097,N_4179);
nand U4478 (N_4478,N_4092,N_4204);
nor U4479 (N_4479,N_4194,N_4130);
nor U4480 (N_4480,N_4183,N_4097);
or U4481 (N_4481,N_4211,N_4219);
nand U4482 (N_4482,N_4204,N_4035);
and U4483 (N_4483,N_4018,N_4183);
and U4484 (N_4484,N_4053,N_4241);
or U4485 (N_4485,N_4112,N_4215);
and U4486 (N_4486,N_4158,N_4189);
nor U4487 (N_4487,N_4169,N_4239);
nand U4488 (N_4488,N_4097,N_4132);
nand U4489 (N_4489,N_4057,N_4018);
or U4490 (N_4490,N_4058,N_4133);
nand U4491 (N_4491,N_4156,N_4003);
and U4492 (N_4492,N_4089,N_4009);
nand U4493 (N_4493,N_4169,N_4050);
nand U4494 (N_4494,N_4205,N_4115);
and U4495 (N_4495,N_4114,N_4220);
and U4496 (N_4496,N_4024,N_4201);
nand U4497 (N_4497,N_4014,N_4125);
and U4498 (N_4498,N_4161,N_4153);
nor U4499 (N_4499,N_4215,N_4116);
nand U4500 (N_4500,N_4398,N_4479);
nor U4501 (N_4501,N_4489,N_4435);
or U4502 (N_4502,N_4270,N_4422);
and U4503 (N_4503,N_4363,N_4366);
nor U4504 (N_4504,N_4325,N_4261);
xnor U4505 (N_4505,N_4466,N_4378);
nand U4506 (N_4506,N_4319,N_4362);
and U4507 (N_4507,N_4394,N_4475);
nor U4508 (N_4508,N_4365,N_4294);
nor U4509 (N_4509,N_4462,N_4258);
nor U4510 (N_4510,N_4382,N_4295);
or U4511 (N_4511,N_4379,N_4340);
or U4512 (N_4512,N_4293,N_4367);
and U4513 (N_4513,N_4472,N_4337);
and U4514 (N_4514,N_4455,N_4368);
nand U4515 (N_4515,N_4432,N_4411);
xnor U4516 (N_4516,N_4463,N_4491);
nand U4517 (N_4517,N_4300,N_4361);
nor U4518 (N_4518,N_4331,N_4346);
nand U4519 (N_4519,N_4381,N_4391);
or U4520 (N_4520,N_4452,N_4454);
xor U4521 (N_4521,N_4495,N_4306);
nor U4522 (N_4522,N_4480,N_4269);
or U4523 (N_4523,N_4288,N_4339);
xor U4524 (N_4524,N_4471,N_4444);
xnor U4525 (N_4525,N_4460,N_4441);
nor U4526 (N_4526,N_4344,N_4449);
nor U4527 (N_4527,N_4386,N_4286);
xor U4528 (N_4528,N_4470,N_4302);
nand U4529 (N_4529,N_4349,N_4324);
and U4530 (N_4530,N_4404,N_4254);
and U4531 (N_4531,N_4267,N_4473);
or U4532 (N_4532,N_4275,N_4464);
and U4533 (N_4533,N_4438,N_4264);
nor U4534 (N_4534,N_4279,N_4380);
nand U4535 (N_4535,N_4373,N_4289);
and U4536 (N_4536,N_4451,N_4375);
nor U4537 (N_4537,N_4414,N_4350);
and U4538 (N_4538,N_4447,N_4303);
or U4539 (N_4539,N_4299,N_4371);
and U4540 (N_4540,N_4320,N_4416);
nand U4541 (N_4541,N_4421,N_4469);
xnor U4542 (N_4542,N_4351,N_4332);
nand U4543 (N_4543,N_4252,N_4429);
nand U4544 (N_4544,N_4266,N_4282);
nand U4545 (N_4545,N_4392,N_4476);
or U4546 (N_4546,N_4403,N_4496);
and U4547 (N_4547,N_4374,N_4376);
or U4548 (N_4548,N_4317,N_4327);
xor U4549 (N_4549,N_4256,N_4312);
nor U4550 (N_4550,N_4385,N_4314);
nand U4551 (N_4551,N_4304,N_4413);
and U4552 (N_4552,N_4310,N_4263);
xor U4553 (N_4553,N_4355,N_4396);
or U4554 (N_4554,N_4410,N_4418);
nor U4555 (N_4555,N_4387,N_4415);
xor U4556 (N_4556,N_4364,N_4399);
or U4557 (N_4557,N_4492,N_4445);
or U4558 (N_4558,N_4250,N_4326);
xor U4559 (N_4559,N_4490,N_4305);
or U4560 (N_4560,N_4271,N_4297);
or U4561 (N_4561,N_4285,N_4276);
or U4562 (N_4562,N_4329,N_4458);
nand U4563 (N_4563,N_4383,N_4465);
xnor U4564 (N_4564,N_4442,N_4430);
nand U4565 (N_4565,N_4352,N_4301);
nor U4566 (N_4566,N_4348,N_4417);
nor U4567 (N_4567,N_4420,N_4409);
and U4568 (N_4568,N_4393,N_4281);
xor U4569 (N_4569,N_4482,N_4316);
nand U4570 (N_4570,N_4359,N_4321);
nand U4571 (N_4571,N_4298,N_4401);
nor U4572 (N_4572,N_4265,N_4290);
nor U4573 (N_4573,N_4426,N_4456);
or U4574 (N_4574,N_4347,N_4330);
or U4575 (N_4575,N_4397,N_4284);
or U4576 (N_4576,N_4313,N_4311);
and U4577 (N_4577,N_4487,N_4259);
xnor U4578 (N_4578,N_4273,N_4283);
xnor U4579 (N_4579,N_4453,N_4253);
or U4580 (N_4580,N_4354,N_4333);
and U4581 (N_4581,N_4488,N_4272);
or U4582 (N_4582,N_4296,N_4424);
xor U4583 (N_4583,N_4372,N_4450);
or U4584 (N_4584,N_4408,N_4307);
and U4585 (N_4585,N_4274,N_4474);
nor U4586 (N_4586,N_4431,N_4443);
xnor U4587 (N_4587,N_4309,N_4497);
nand U4588 (N_4588,N_4322,N_4377);
or U4589 (N_4589,N_4437,N_4434);
and U4590 (N_4590,N_4423,N_4477);
xnor U4591 (N_4591,N_4356,N_4440);
and U4592 (N_4592,N_4268,N_4459);
and U4593 (N_4593,N_4419,N_4483);
or U4594 (N_4594,N_4433,N_4448);
or U4595 (N_4595,N_4478,N_4323);
or U4596 (N_4596,N_4494,N_4315);
xnor U4597 (N_4597,N_4278,N_4407);
nand U4598 (N_4598,N_4498,N_4342);
and U4599 (N_4599,N_4338,N_4395);
nor U4600 (N_4600,N_4428,N_4360);
xor U4601 (N_4601,N_4389,N_4357);
nor U4602 (N_4602,N_4336,N_4390);
and U4603 (N_4603,N_4427,N_4493);
or U4604 (N_4604,N_4260,N_4277);
or U4605 (N_4605,N_4406,N_4353);
nand U4606 (N_4606,N_4499,N_4439);
or U4607 (N_4607,N_4280,N_4484);
or U4608 (N_4608,N_4345,N_4369);
and U4609 (N_4609,N_4328,N_4402);
nor U4610 (N_4610,N_4425,N_4468);
nor U4611 (N_4611,N_4251,N_4308);
nor U4612 (N_4612,N_4412,N_4467);
or U4613 (N_4613,N_4405,N_4318);
nor U4614 (N_4614,N_4255,N_4400);
or U4615 (N_4615,N_4358,N_4461);
and U4616 (N_4616,N_4370,N_4292);
or U4617 (N_4617,N_4262,N_4486);
nor U4618 (N_4618,N_4388,N_4343);
nor U4619 (N_4619,N_4334,N_4287);
and U4620 (N_4620,N_4384,N_4291);
xnor U4621 (N_4621,N_4436,N_4485);
xor U4622 (N_4622,N_4335,N_4457);
xnor U4623 (N_4623,N_4481,N_4341);
nor U4624 (N_4624,N_4257,N_4446);
nor U4625 (N_4625,N_4389,N_4289);
nand U4626 (N_4626,N_4442,N_4283);
nor U4627 (N_4627,N_4262,N_4368);
xnor U4628 (N_4628,N_4317,N_4391);
and U4629 (N_4629,N_4278,N_4454);
xor U4630 (N_4630,N_4452,N_4380);
or U4631 (N_4631,N_4316,N_4423);
or U4632 (N_4632,N_4494,N_4359);
nor U4633 (N_4633,N_4431,N_4292);
nand U4634 (N_4634,N_4268,N_4396);
nor U4635 (N_4635,N_4356,N_4315);
and U4636 (N_4636,N_4280,N_4439);
or U4637 (N_4637,N_4460,N_4341);
or U4638 (N_4638,N_4307,N_4279);
or U4639 (N_4639,N_4389,N_4392);
xnor U4640 (N_4640,N_4449,N_4396);
or U4641 (N_4641,N_4434,N_4276);
nor U4642 (N_4642,N_4422,N_4278);
nor U4643 (N_4643,N_4408,N_4409);
nand U4644 (N_4644,N_4483,N_4322);
or U4645 (N_4645,N_4251,N_4456);
or U4646 (N_4646,N_4471,N_4355);
and U4647 (N_4647,N_4396,N_4414);
xor U4648 (N_4648,N_4258,N_4478);
or U4649 (N_4649,N_4347,N_4363);
or U4650 (N_4650,N_4442,N_4439);
and U4651 (N_4651,N_4263,N_4368);
nor U4652 (N_4652,N_4365,N_4290);
nand U4653 (N_4653,N_4378,N_4476);
nor U4654 (N_4654,N_4320,N_4259);
nor U4655 (N_4655,N_4438,N_4308);
nand U4656 (N_4656,N_4250,N_4475);
nand U4657 (N_4657,N_4312,N_4311);
or U4658 (N_4658,N_4468,N_4333);
nand U4659 (N_4659,N_4355,N_4348);
and U4660 (N_4660,N_4449,N_4339);
nand U4661 (N_4661,N_4252,N_4392);
and U4662 (N_4662,N_4437,N_4371);
xnor U4663 (N_4663,N_4282,N_4438);
nor U4664 (N_4664,N_4385,N_4320);
nand U4665 (N_4665,N_4272,N_4285);
xnor U4666 (N_4666,N_4405,N_4429);
nand U4667 (N_4667,N_4491,N_4379);
nor U4668 (N_4668,N_4307,N_4250);
nor U4669 (N_4669,N_4311,N_4441);
xnor U4670 (N_4670,N_4303,N_4442);
nor U4671 (N_4671,N_4360,N_4498);
or U4672 (N_4672,N_4374,N_4279);
xnor U4673 (N_4673,N_4491,N_4457);
and U4674 (N_4674,N_4495,N_4327);
nand U4675 (N_4675,N_4481,N_4469);
and U4676 (N_4676,N_4478,N_4383);
and U4677 (N_4677,N_4314,N_4379);
xor U4678 (N_4678,N_4324,N_4306);
nor U4679 (N_4679,N_4446,N_4370);
and U4680 (N_4680,N_4465,N_4412);
nand U4681 (N_4681,N_4396,N_4336);
and U4682 (N_4682,N_4455,N_4481);
and U4683 (N_4683,N_4276,N_4266);
and U4684 (N_4684,N_4347,N_4343);
or U4685 (N_4685,N_4377,N_4427);
xnor U4686 (N_4686,N_4304,N_4352);
or U4687 (N_4687,N_4273,N_4322);
xnor U4688 (N_4688,N_4430,N_4407);
xor U4689 (N_4689,N_4380,N_4333);
or U4690 (N_4690,N_4376,N_4494);
or U4691 (N_4691,N_4337,N_4452);
nor U4692 (N_4692,N_4422,N_4288);
and U4693 (N_4693,N_4279,N_4333);
and U4694 (N_4694,N_4445,N_4417);
or U4695 (N_4695,N_4427,N_4307);
xor U4696 (N_4696,N_4269,N_4435);
or U4697 (N_4697,N_4299,N_4446);
nand U4698 (N_4698,N_4476,N_4467);
xor U4699 (N_4699,N_4489,N_4476);
nor U4700 (N_4700,N_4287,N_4370);
xor U4701 (N_4701,N_4328,N_4442);
xor U4702 (N_4702,N_4329,N_4478);
or U4703 (N_4703,N_4454,N_4359);
nand U4704 (N_4704,N_4253,N_4494);
and U4705 (N_4705,N_4440,N_4340);
nand U4706 (N_4706,N_4477,N_4388);
or U4707 (N_4707,N_4347,N_4450);
or U4708 (N_4708,N_4316,N_4461);
nand U4709 (N_4709,N_4404,N_4350);
or U4710 (N_4710,N_4272,N_4473);
xor U4711 (N_4711,N_4490,N_4350);
nor U4712 (N_4712,N_4259,N_4466);
or U4713 (N_4713,N_4342,N_4414);
or U4714 (N_4714,N_4399,N_4265);
nand U4715 (N_4715,N_4332,N_4273);
nand U4716 (N_4716,N_4497,N_4314);
nor U4717 (N_4717,N_4399,N_4452);
nand U4718 (N_4718,N_4285,N_4280);
nand U4719 (N_4719,N_4478,N_4453);
nand U4720 (N_4720,N_4360,N_4302);
xnor U4721 (N_4721,N_4258,N_4404);
and U4722 (N_4722,N_4386,N_4435);
nor U4723 (N_4723,N_4497,N_4499);
and U4724 (N_4724,N_4323,N_4495);
nor U4725 (N_4725,N_4427,N_4354);
nand U4726 (N_4726,N_4450,N_4471);
xnor U4727 (N_4727,N_4262,N_4250);
nand U4728 (N_4728,N_4478,N_4456);
and U4729 (N_4729,N_4369,N_4375);
xor U4730 (N_4730,N_4325,N_4328);
nand U4731 (N_4731,N_4367,N_4429);
or U4732 (N_4732,N_4461,N_4269);
nand U4733 (N_4733,N_4453,N_4493);
nor U4734 (N_4734,N_4427,N_4413);
or U4735 (N_4735,N_4383,N_4423);
nor U4736 (N_4736,N_4460,N_4423);
nor U4737 (N_4737,N_4485,N_4492);
xor U4738 (N_4738,N_4430,N_4408);
and U4739 (N_4739,N_4466,N_4261);
and U4740 (N_4740,N_4280,N_4358);
and U4741 (N_4741,N_4412,N_4329);
or U4742 (N_4742,N_4363,N_4344);
or U4743 (N_4743,N_4321,N_4281);
nand U4744 (N_4744,N_4486,N_4369);
nor U4745 (N_4745,N_4334,N_4476);
or U4746 (N_4746,N_4359,N_4283);
nor U4747 (N_4747,N_4435,N_4345);
xnor U4748 (N_4748,N_4407,N_4378);
nor U4749 (N_4749,N_4318,N_4382);
nor U4750 (N_4750,N_4549,N_4583);
and U4751 (N_4751,N_4627,N_4626);
nand U4752 (N_4752,N_4609,N_4538);
and U4753 (N_4753,N_4636,N_4648);
or U4754 (N_4754,N_4713,N_4742);
xnor U4755 (N_4755,N_4666,N_4630);
nand U4756 (N_4756,N_4574,N_4502);
nand U4757 (N_4757,N_4619,N_4646);
nor U4758 (N_4758,N_4537,N_4731);
nor U4759 (N_4759,N_4696,N_4661);
and U4760 (N_4760,N_4730,N_4718);
xnor U4761 (N_4761,N_4726,N_4504);
nand U4762 (N_4762,N_4519,N_4680);
xor U4763 (N_4763,N_4584,N_4581);
nor U4764 (N_4764,N_4640,N_4684);
nand U4765 (N_4765,N_4709,N_4722);
nor U4766 (N_4766,N_4653,N_4501);
or U4767 (N_4767,N_4605,N_4539);
or U4768 (N_4768,N_4566,N_4523);
and U4769 (N_4769,N_4591,N_4725);
and U4770 (N_4770,N_4582,N_4513);
and U4771 (N_4771,N_4589,N_4535);
nand U4772 (N_4772,N_4520,N_4724);
and U4773 (N_4773,N_4531,N_4647);
xor U4774 (N_4774,N_4565,N_4685);
nor U4775 (N_4775,N_4576,N_4559);
and U4776 (N_4776,N_4500,N_4623);
nand U4777 (N_4777,N_4708,N_4712);
or U4778 (N_4778,N_4515,N_4701);
nand U4779 (N_4779,N_4541,N_4606);
and U4780 (N_4780,N_4675,N_4747);
xnor U4781 (N_4781,N_4621,N_4598);
nor U4782 (N_4782,N_4620,N_4649);
and U4783 (N_4783,N_4643,N_4656);
nor U4784 (N_4784,N_4737,N_4560);
xnor U4785 (N_4785,N_4509,N_4664);
nand U4786 (N_4786,N_4704,N_4600);
nor U4787 (N_4787,N_4614,N_4608);
or U4788 (N_4788,N_4575,N_4690);
nand U4789 (N_4789,N_4544,N_4668);
or U4790 (N_4790,N_4602,N_4601);
xnor U4791 (N_4791,N_4551,N_4728);
and U4792 (N_4792,N_4596,N_4545);
or U4793 (N_4793,N_4667,N_4510);
and U4794 (N_4794,N_4683,N_4610);
nor U4795 (N_4795,N_4739,N_4514);
xor U4796 (N_4796,N_4613,N_4695);
or U4797 (N_4797,N_4716,N_4700);
xnor U4798 (N_4798,N_4736,N_4632);
or U4799 (N_4799,N_4705,N_4590);
xnor U4800 (N_4800,N_4554,N_4748);
xnor U4801 (N_4801,N_4518,N_4524);
or U4802 (N_4802,N_4522,N_4593);
xnor U4803 (N_4803,N_4548,N_4727);
nor U4804 (N_4804,N_4557,N_4563);
xor U4805 (N_4805,N_4687,N_4585);
nor U4806 (N_4806,N_4635,N_4660);
and U4807 (N_4807,N_4542,N_4677);
and U4808 (N_4808,N_4703,N_4633);
nand U4809 (N_4809,N_4597,N_4517);
nor U4810 (N_4810,N_4707,N_4672);
nor U4811 (N_4811,N_4503,N_4568);
and U4812 (N_4812,N_4719,N_4592);
and U4813 (N_4813,N_4611,N_4603);
xor U4814 (N_4814,N_4612,N_4670);
xor U4815 (N_4815,N_4629,N_4564);
or U4816 (N_4816,N_4512,N_4587);
xnor U4817 (N_4817,N_4655,N_4644);
nand U4818 (N_4818,N_4580,N_4735);
nor U4819 (N_4819,N_4671,N_4599);
or U4820 (N_4820,N_4749,N_4658);
nor U4821 (N_4821,N_4721,N_4521);
or U4822 (N_4822,N_4579,N_4546);
xor U4823 (N_4823,N_4540,N_4723);
and U4824 (N_4824,N_4536,N_4665);
and U4825 (N_4825,N_4673,N_4622);
nor U4826 (N_4826,N_4654,N_4552);
and U4827 (N_4827,N_4691,N_4604);
and U4828 (N_4828,N_4530,N_4637);
nand U4829 (N_4829,N_4689,N_4738);
or U4830 (N_4830,N_4692,N_4697);
xor U4831 (N_4831,N_4516,N_4714);
nand U4832 (N_4832,N_4642,N_4676);
or U4833 (N_4833,N_4717,N_4631);
or U4834 (N_4834,N_4688,N_4645);
nor U4835 (N_4835,N_4650,N_4618);
or U4836 (N_4836,N_4659,N_4570);
xor U4837 (N_4837,N_4543,N_4741);
xnor U4838 (N_4838,N_4625,N_4533);
xor U4839 (N_4839,N_4594,N_4720);
xor U4840 (N_4840,N_4569,N_4639);
and U4841 (N_4841,N_4553,N_4617);
and U4842 (N_4842,N_4527,N_4556);
xnor U4843 (N_4843,N_4662,N_4744);
nand U4844 (N_4844,N_4550,N_4555);
nand U4845 (N_4845,N_4508,N_4710);
nor U4846 (N_4846,N_4669,N_4711);
nand U4847 (N_4847,N_4706,N_4595);
nor U4848 (N_4848,N_4562,N_4682);
or U4849 (N_4849,N_4578,N_4624);
nand U4850 (N_4850,N_4526,N_4734);
or U4851 (N_4851,N_4715,N_4686);
and U4852 (N_4852,N_4693,N_4586);
and U4853 (N_4853,N_4634,N_4740);
or U4854 (N_4854,N_4641,N_4615);
and U4855 (N_4855,N_4507,N_4505);
xor U4856 (N_4856,N_4607,N_4674);
nand U4857 (N_4857,N_4572,N_4529);
nand U4858 (N_4858,N_4506,N_4532);
xor U4859 (N_4859,N_4694,N_4681);
nor U4860 (N_4860,N_4573,N_4547);
or U4861 (N_4861,N_4679,N_4588);
and U4862 (N_4862,N_4571,N_4743);
or U4863 (N_4863,N_4616,N_4534);
and U4864 (N_4864,N_4651,N_4577);
or U4865 (N_4865,N_4528,N_4628);
xnor U4866 (N_4866,N_4663,N_4733);
xnor U4867 (N_4867,N_4746,N_4729);
xor U4868 (N_4868,N_4561,N_4732);
nand U4869 (N_4869,N_4699,N_4702);
nor U4870 (N_4870,N_4638,N_4567);
or U4871 (N_4871,N_4698,N_4525);
xor U4872 (N_4872,N_4678,N_4657);
xor U4873 (N_4873,N_4558,N_4511);
nand U4874 (N_4874,N_4745,N_4652);
nor U4875 (N_4875,N_4686,N_4625);
nand U4876 (N_4876,N_4545,N_4634);
and U4877 (N_4877,N_4717,N_4739);
and U4878 (N_4878,N_4709,N_4654);
and U4879 (N_4879,N_4589,N_4746);
nand U4880 (N_4880,N_4605,N_4520);
nand U4881 (N_4881,N_4647,N_4594);
or U4882 (N_4882,N_4589,N_4583);
nor U4883 (N_4883,N_4570,N_4679);
nor U4884 (N_4884,N_4663,N_4619);
nor U4885 (N_4885,N_4560,N_4665);
nor U4886 (N_4886,N_4555,N_4507);
or U4887 (N_4887,N_4657,N_4718);
nand U4888 (N_4888,N_4717,N_4506);
and U4889 (N_4889,N_4516,N_4603);
xor U4890 (N_4890,N_4736,N_4649);
or U4891 (N_4891,N_4649,N_4692);
or U4892 (N_4892,N_4739,N_4695);
and U4893 (N_4893,N_4684,N_4622);
nand U4894 (N_4894,N_4746,N_4707);
or U4895 (N_4895,N_4660,N_4562);
or U4896 (N_4896,N_4578,N_4641);
or U4897 (N_4897,N_4615,N_4633);
and U4898 (N_4898,N_4737,N_4644);
nor U4899 (N_4899,N_4616,N_4632);
or U4900 (N_4900,N_4511,N_4623);
and U4901 (N_4901,N_4689,N_4573);
xnor U4902 (N_4902,N_4681,N_4706);
xnor U4903 (N_4903,N_4592,N_4577);
and U4904 (N_4904,N_4651,N_4684);
and U4905 (N_4905,N_4725,N_4555);
nand U4906 (N_4906,N_4706,N_4606);
xnor U4907 (N_4907,N_4560,N_4598);
and U4908 (N_4908,N_4535,N_4607);
nor U4909 (N_4909,N_4500,N_4689);
nand U4910 (N_4910,N_4741,N_4596);
nor U4911 (N_4911,N_4687,N_4559);
nor U4912 (N_4912,N_4550,N_4540);
xor U4913 (N_4913,N_4577,N_4578);
nand U4914 (N_4914,N_4736,N_4708);
nor U4915 (N_4915,N_4658,N_4540);
or U4916 (N_4916,N_4511,N_4715);
nor U4917 (N_4917,N_4543,N_4624);
or U4918 (N_4918,N_4572,N_4580);
and U4919 (N_4919,N_4623,N_4602);
or U4920 (N_4920,N_4662,N_4501);
xor U4921 (N_4921,N_4730,N_4542);
xor U4922 (N_4922,N_4670,N_4625);
or U4923 (N_4923,N_4740,N_4701);
nand U4924 (N_4924,N_4559,N_4728);
xor U4925 (N_4925,N_4727,N_4741);
and U4926 (N_4926,N_4525,N_4652);
or U4927 (N_4927,N_4507,N_4700);
nor U4928 (N_4928,N_4587,N_4700);
nor U4929 (N_4929,N_4509,N_4739);
nand U4930 (N_4930,N_4661,N_4620);
nand U4931 (N_4931,N_4643,N_4562);
nand U4932 (N_4932,N_4562,N_4671);
or U4933 (N_4933,N_4694,N_4516);
nor U4934 (N_4934,N_4698,N_4733);
and U4935 (N_4935,N_4603,N_4673);
nor U4936 (N_4936,N_4613,N_4519);
or U4937 (N_4937,N_4636,N_4710);
and U4938 (N_4938,N_4532,N_4681);
nor U4939 (N_4939,N_4500,N_4546);
nor U4940 (N_4940,N_4724,N_4679);
or U4941 (N_4941,N_4544,N_4739);
or U4942 (N_4942,N_4723,N_4515);
nand U4943 (N_4943,N_4620,N_4591);
xor U4944 (N_4944,N_4588,N_4512);
nand U4945 (N_4945,N_4530,N_4546);
nor U4946 (N_4946,N_4608,N_4615);
and U4947 (N_4947,N_4522,N_4544);
and U4948 (N_4948,N_4656,N_4607);
nand U4949 (N_4949,N_4539,N_4589);
or U4950 (N_4950,N_4567,N_4657);
and U4951 (N_4951,N_4569,N_4703);
or U4952 (N_4952,N_4647,N_4579);
and U4953 (N_4953,N_4715,N_4739);
or U4954 (N_4954,N_4690,N_4595);
and U4955 (N_4955,N_4738,N_4589);
and U4956 (N_4956,N_4627,N_4605);
nor U4957 (N_4957,N_4671,N_4693);
xor U4958 (N_4958,N_4668,N_4658);
and U4959 (N_4959,N_4742,N_4567);
nor U4960 (N_4960,N_4702,N_4533);
or U4961 (N_4961,N_4598,N_4676);
or U4962 (N_4962,N_4722,N_4569);
xnor U4963 (N_4963,N_4571,N_4620);
and U4964 (N_4964,N_4601,N_4715);
or U4965 (N_4965,N_4640,N_4570);
nor U4966 (N_4966,N_4706,N_4561);
xnor U4967 (N_4967,N_4720,N_4733);
nand U4968 (N_4968,N_4526,N_4682);
nor U4969 (N_4969,N_4560,N_4540);
xnor U4970 (N_4970,N_4748,N_4637);
nand U4971 (N_4971,N_4532,N_4609);
or U4972 (N_4972,N_4730,N_4550);
and U4973 (N_4973,N_4608,N_4622);
or U4974 (N_4974,N_4622,N_4566);
nor U4975 (N_4975,N_4581,N_4639);
nor U4976 (N_4976,N_4540,N_4630);
nor U4977 (N_4977,N_4673,N_4533);
and U4978 (N_4978,N_4678,N_4601);
xnor U4979 (N_4979,N_4515,N_4731);
or U4980 (N_4980,N_4657,N_4569);
xnor U4981 (N_4981,N_4620,N_4672);
nor U4982 (N_4982,N_4604,N_4525);
xor U4983 (N_4983,N_4635,N_4503);
xor U4984 (N_4984,N_4666,N_4566);
xor U4985 (N_4985,N_4686,N_4653);
and U4986 (N_4986,N_4505,N_4687);
and U4987 (N_4987,N_4714,N_4697);
nor U4988 (N_4988,N_4685,N_4635);
nand U4989 (N_4989,N_4642,N_4582);
nand U4990 (N_4990,N_4501,N_4504);
xnor U4991 (N_4991,N_4738,N_4655);
and U4992 (N_4992,N_4707,N_4572);
or U4993 (N_4993,N_4720,N_4506);
nand U4994 (N_4994,N_4549,N_4510);
and U4995 (N_4995,N_4650,N_4558);
and U4996 (N_4996,N_4606,N_4655);
nand U4997 (N_4997,N_4647,N_4733);
nor U4998 (N_4998,N_4547,N_4545);
nor U4999 (N_4999,N_4564,N_4547);
and U5000 (N_5000,N_4964,N_4871);
nand U5001 (N_5001,N_4764,N_4886);
or U5002 (N_5002,N_4856,N_4754);
xnor U5003 (N_5003,N_4908,N_4905);
or U5004 (N_5004,N_4831,N_4922);
xnor U5005 (N_5005,N_4877,N_4775);
nor U5006 (N_5006,N_4891,N_4809);
nand U5007 (N_5007,N_4954,N_4950);
nor U5008 (N_5008,N_4949,N_4766);
nor U5009 (N_5009,N_4872,N_4857);
xor U5010 (N_5010,N_4889,N_4923);
nand U5011 (N_5011,N_4821,N_4795);
nand U5012 (N_5012,N_4878,N_4783);
nor U5013 (N_5013,N_4892,N_4909);
nor U5014 (N_5014,N_4761,N_4890);
or U5015 (N_5015,N_4963,N_4934);
xor U5016 (N_5016,N_4976,N_4753);
nand U5017 (N_5017,N_4815,N_4958);
nand U5018 (N_5018,N_4813,N_4803);
xor U5019 (N_5019,N_4789,N_4942);
and U5020 (N_5020,N_4893,N_4854);
nor U5021 (N_5021,N_4990,N_4955);
nand U5022 (N_5022,N_4796,N_4822);
or U5023 (N_5023,N_4818,N_4769);
xnor U5024 (N_5024,N_4919,N_4842);
and U5025 (N_5025,N_4910,N_4814);
nand U5026 (N_5026,N_4888,N_4838);
xnor U5027 (N_5027,N_4907,N_4972);
xor U5028 (N_5028,N_4758,N_4782);
and U5029 (N_5029,N_4962,N_4874);
nor U5030 (N_5030,N_4985,N_4757);
and U5031 (N_5031,N_4866,N_4847);
and U5032 (N_5032,N_4793,N_4810);
xor U5033 (N_5033,N_4875,N_4873);
or U5034 (N_5034,N_4924,N_4816);
nand U5035 (N_5035,N_4956,N_4846);
and U5036 (N_5036,N_4997,N_4841);
xor U5037 (N_5037,N_4975,N_4953);
nor U5038 (N_5038,N_4869,N_4999);
nor U5039 (N_5039,N_4863,N_4870);
nor U5040 (N_5040,N_4802,N_4834);
xor U5041 (N_5041,N_4798,N_4767);
and U5042 (N_5042,N_4849,N_4836);
nand U5043 (N_5043,N_4974,N_4931);
nand U5044 (N_5044,N_4845,N_4968);
and U5045 (N_5045,N_4765,N_4797);
nor U5046 (N_5046,N_4933,N_4884);
or U5047 (N_5047,N_4947,N_4938);
and U5048 (N_5048,N_4926,N_4925);
nand U5049 (N_5049,N_4763,N_4986);
nor U5050 (N_5050,N_4832,N_4952);
and U5051 (N_5051,N_4996,N_4858);
nand U5052 (N_5052,N_4887,N_4799);
nand U5053 (N_5053,N_4776,N_4983);
and U5054 (N_5054,N_4973,N_4855);
xnor U5055 (N_5055,N_4794,N_4751);
xnor U5056 (N_5056,N_4957,N_4801);
xnor U5057 (N_5057,N_4928,N_4839);
xnor U5058 (N_5058,N_4921,N_4773);
nor U5059 (N_5059,N_4808,N_4840);
nand U5060 (N_5060,N_4807,N_4786);
xor U5061 (N_5061,N_4812,N_4937);
xor U5062 (N_5062,N_4768,N_4774);
or U5063 (N_5063,N_4800,N_4959);
or U5064 (N_5064,N_4916,N_4880);
or U5065 (N_5065,N_4904,N_4784);
or U5066 (N_5066,N_4785,N_4790);
or U5067 (N_5067,N_4897,N_4804);
and U5068 (N_5068,N_4970,N_4939);
nor U5069 (N_5069,N_4759,N_4932);
nor U5070 (N_5070,N_4762,N_4912);
nor U5071 (N_5071,N_4966,N_4779);
and U5072 (N_5072,N_4876,N_4824);
nor U5073 (N_5073,N_4825,N_4944);
nor U5074 (N_5074,N_4971,N_4778);
and U5075 (N_5075,N_4965,N_4830);
and U5076 (N_5076,N_4998,N_4993);
nand U5077 (N_5077,N_4755,N_4752);
or U5078 (N_5078,N_4899,N_4982);
nand U5079 (N_5079,N_4867,N_4935);
nand U5080 (N_5080,N_4991,N_4852);
xor U5081 (N_5081,N_4918,N_4981);
nand U5082 (N_5082,N_4920,N_4994);
or U5083 (N_5083,N_4930,N_4819);
or U5084 (N_5084,N_4817,N_4850);
or U5085 (N_5085,N_4969,N_4929);
and U5086 (N_5086,N_4960,N_4977);
and U5087 (N_5087,N_4980,N_4978);
xor U5088 (N_5088,N_4948,N_4914);
nor U5089 (N_5089,N_4760,N_4826);
or U5090 (N_5090,N_4946,N_4806);
nand U5091 (N_5091,N_4860,N_4805);
nor U5092 (N_5092,N_4859,N_4777);
or U5093 (N_5093,N_4750,N_4936);
nand U5094 (N_5094,N_4895,N_4791);
xnor U5095 (N_5095,N_4792,N_4979);
or U5096 (N_5096,N_4882,N_4833);
nor U5097 (N_5097,N_4848,N_4829);
and U5098 (N_5098,N_4992,N_4772);
or U5099 (N_5099,N_4828,N_4835);
xnor U5100 (N_5100,N_4898,N_4896);
or U5101 (N_5101,N_4940,N_4881);
xnor U5102 (N_5102,N_4901,N_4915);
nor U5103 (N_5103,N_4943,N_4913);
nand U5104 (N_5104,N_4811,N_4781);
nor U5105 (N_5105,N_4823,N_4883);
and U5106 (N_5106,N_4906,N_4902);
nor U5107 (N_5107,N_4961,N_4868);
nor U5108 (N_5108,N_4820,N_4756);
xnor U5109 (N_5109,N_4843,N_4780);
and U5110 (N_5110,N_4837,N_4844);
and U5111 (N_5111,N_4885,N_4879);
and U5112 (N_5112,N_4911,N_4851);
and U5113 (N_5113,N_4900,N_4984);
or U5114 (N_5114,N_4827,N_4861);
and U5115 (N_5115,N_4987,N_4788);
nor U5116 (N_5116,N_4951,N_4917);
or U5117 (N_5117,N_4787,N_4941);
nor U5118 (N_5118,N_4903,N_4967);
or U5119 (N_5119,N_4862,N_4853);
and U5120 (N_5120,N_4894,N_4770);
or U5121 (N_5121,N_4927,N_4864);
and U5122 (N_5122,N_4988,N_4865);
or U5123 (N_5123,N_4995,N_4945);
nand U5124 (N_5124,N_4771,N_4989);
xnor U5125 (N_5125,N_4852,N_4857);
nor U5126 (N_5126,N_4845,N_4859);
or U5127 (N_5127,N_4874,N_4901);
or U5128 (N_5128,N_4799,N_4993);
xnor U5129 (N_5129,N_4937,N_4855);
or U5130 (N_5130,N_4838,N_4891);
xnor U5131 (N_5131,N_4987,N_4996);
nand U5132 (N_5132,N_4929,N_4964);
or U5133 (N_5133,N_4826,N_4945);
nor U5134 (N_5134,N_4929,N_4801);
nor U5135 (N_5135,N_4973,N_4856);
xnor U5136 (N_5136,N_4883,N_4969);
xor U5137 (N_5137,N_4785,N_4942);
and U5138 (N_5138,N_4778,N_4801);
or U5139 (N_5139,N_4768,N_4887);
nand U5140 (N_5140,N_4899,N_4986);
and U5141 (N_5141,N_4899,N_4801);
or U5142 (N_5142,N_4833,N_4772);
nand U5143 (N_5143,N_4880,N_4945);
nor U5144 (N_5144,N_4832,N_4925);
nor U5145 (N_5145,N_4993,N_4972);
nor U5146 (N_5146,N_4892,N_4834);
nand U5147 (N_5147,N_4903,N_4794);
nor U5148 (N_5148,N_4932,N_4893);
or U5149 (N_5149,N_4773,N_4814);
nand U5150 (N_5150,N_4983,N_4789);
or U5151 (N_5151,N_4943,N_4938);
nand U5152 (N_5152,N_4923,N_4816);
and U5153 (N_5153,N_4814,N_4956);
nor U5154 (N_5154,N_4858,N_4864);
xnor U5155 (N_5155,N_4903,N_4899);
or U5156 (N_5156,N_4997,N_4820);
nor U5157 (N_5157,N_4945,N_4764);
or U5158 (N_5158,N_4809,N_4907);
or U5159 (N_5159,N_4838,N_4856);
and U5160 (N_5160,N_4855,N_4965);
nand U5161 (N_5161,N_4841,N_4784);
and U5162 (N_5162,N_4962,N_4925);
nand U5163 (N_5163,N_4769,N_4788);
nor U5164 (N_5164,N_4835,N_4988);
xnor U5165 (N_5165,N_4767,N_4857);
nor U5166 (N_5166,N_4919,N_4870);
or U5167 (N_5167,N_4846,N_4884);
nor U5168 (N_5168,N_4900,N_4757);
and U5169 (N_5169,N_4763,N_4828);
nand U5170 (N_5170,N_4892,N_4875);
nand U5171 (N_5171,N_4794,N_4979);
and U5172 (N_5172,N_4823,N_4804);
and U5173 (N_5173,N_4813,N_4858);
and U5174 (N_5174,N_4773,N_4791);
and U5175 (N_5175,N_4812,N_4873);
nor U5176 (N_5176,N_4942,N_4881);
nand U5177 (N_5177,N_4868,N_4969);
and U5178 (N_5178,N_4750,N_4794);
nor U5179 (N_5179,N_4902,N_4755);
and U5180 (N_5180,N_4920,N_4926);
or U5181 (N_5181,N_4920,N_4953);
xor U5182 (N_5182,N_4870,N_4878);
xnor U5183 (N_5183,N_4920,N_4793);
xnor U5184 (N_5184,N_4919,N_4907);
nor U5185 (N_5185,N_4806,N_4939);
xnor U5186 (N_5186,N_4990,N_4894);
xnor U5187 (N_5187,N_4862,N_4762);
xnor U5188 (N_5188,N_4935,N_4918);
or U5189 (N_5189,N_4835,N_4841);
or U5190 (N_5190,N_4859,N_4908);
nand U5191 (N_5191,N_4986,N_4800);
or U5192 (N_5192,N_4865,N_4933);
nand U5193 (N_5193,N_4945,N_4770);
xor U5194 (N_5194,N_4772,N_4968);
and U5195 (N_5195,N_4791,N_4913);
and U5196 (N_5196,N_4809,N_4892);
and U5197 (N_5197,N_4847,N_4885);
xor U5198 (N_5198,N_4826,N_4847);
xor U5199 (N_5199,N_4973,N_4890);
and U5200 (N_5200,N_4847,N_4936);
or U5201 (N_5201,N_4787,N_4833);
nand U5202 (N_5202,N_4873,N_4805);
nor U5203 (N_5203,N_4957,N_4983);
or U5204 (N_5204,N_4873,N_4872);
nor U5205 (N_5205,N_4917,N_4836);
nand U5206 (N_5206,N_4915,N_4916);
and U5207 (N_5207,N_4792,N_4940);
or U5208 (N_5208,N_4971,N_4888);
xor U5209 (N_5209,N_4816,N_4836);
xnor U5210 (N_5210,N_4802,N_4839);
nand U5211 (N_5211,N_4934,N_4793);
and U5212 (N_5212,N_4892,N_4975);
or U5213 (N_5213,N_4772,N_4997);
nor U5214 (N_5214,N_4814,N_4912);
nand U5215 (N_5215,N_4926,N_4826);
or U5216 (N_5216,N_4937,N_4801);
or U5217 (N_5217,N_4861,N_4776);
nor U5218 (N_5218,N_4783,N_4991);
or U5219 (N_5219,N_4775,N_4852);
or U5220 (N_5220,N_4946,N_4905);
nand U5221 (N_5221,N_4810,N_4796);
xor U5222 (N_5222,N_4791,N_4756);
and U5223 (N_5223,N_4829,N_4891);
xor U5224 (N_5224,N_4849,N_4812);
and U5225 (N_5225,N_4895,N_4889);
and U5226 (N_5226,N_4812,N_4915);
nand U5227 (N_5227,N_4920,N_4818);
nor U5228 (N_5228,N_4768,N_4923);
or U5229 (N_5229,N_4753,N_4778);
or U5230 (N_5230,N_4838,N_4901);
nand U5231 (N_5231,N_4806,N_4816);
or U5232 (N_5232,N_4919,N_4882);
xnor U5233 (N_5233,N_4945,N_4964);
or U5234 (N_5234,N_4852,N_4978);
or U5235 (N_5235,N_4795,N_4894);
nand U5236 (N_5236,N_4826,N_4934);
nand U5237 (N_5237,N_4866,N_4958);
xor U5238 (N_5238,N_4819,N_4921);
or U5239 (N_5239,N_4815,N_4869);
or U5240 (N_5240,N_4883,N_4973);
and U5241 (N_5241,N_4892,N_4811);
and U5242 (N_5242,N_4793,N_4868);
xnor U5243 (N_5243,N_4983,N_4813);
and U5244 (N_5244,N_4953,N_4905);
or U5245 (N_5245,N_4983,N_4950);
or U5246 (N_5246,N_4843,N_4985);
and U5247 (N_5247,N_4912,N_4801);
and U5248 (N_5248,N_4914,N_4908);
and U5249 (N_5249,N_4842,N_4984);
xor U5250 (N_5250,N_5210,N_5067);
nor U5251 (N_5251,N_5023,N_5055);
xnor U5252 (N_5252,N_5083,N_5170);
nor U5253 (N_5253,N_5179,N_5020);
and U5254 (N_5254,N_5006,N_5040);
and U5255 (N_5255,N_5019,N_5117);
nand U5256 (N_5256,N_5120,N_5014);
nand U5257 (N_5257,N_5143,N_5072);
nand U5258 (N_5258,N_5176,N_5090);
and U5259 (N_5259,N_5193,N_5198);
or U5260 (N_5260,N_5099,N_5241);
nand U5261 (N_5261,N_5025,N_5157);
nand U5262 (N_5262,N_5042,N_5121);
nor U5263 (N_5263,N_5208,N_5249);
nor U5264 (N_5264,N_5026,N_5008);
or U5265 (N_5265,N_5203,N_5087);
xor U5266 (N_5266,N_5235,N_5105);
or U5267 (N_5267,N_5244,N_5243);
and U5268 (N_5268,N_5155,N_5205);
and U5269 (N_5269,N_5147,N_5233);
xor U5270 (N_5270,N_5237,N_5015);
or U5271 (N_5271,N_5005,N_5052);
and U5272 (N_5272,N_5148,N_5082);
xor U5273 (N_5273,N_5166,N_5225);
and U5274 (N_5274,N_5207,N_5064);
and U5275 (N_5275,N_5038,N_5194);
nor U5276 (N_5276,N_5178,N_5065);
and U5277 (N_5277,N_5124,N_5118);
xnor U5278 (N_5278,N_5007,N_5130);
nor U5279 (N_5279,N_5238,N_5127);
or U5280 (N_5280,N_5114,N_5131);
and U5281 (N_5281,N_5151,N_5200);
and U5282 (N_5282,N_5069,N_5141);
nor U5283 (N_5283,N_5165,N_5076);
nor U5284 (N_5284,N_5220,N_5097);
or U5285 (N_5285,N_5027,N_5214);
nor U5286 (N_5286,N_5041,N_5000);
nor U5287 (N_5287,N_5231,N_5183);
and U5288 (N_5288,N_5144,N_5016);
xor U5289 (N_5289,N_5248,N_5240);
or U5290 (N_5290,N_5091,N_5011);
nand U5291 (N_5291,N_5095,N_5122);
and U5292 (N_5292,N_5145,N_5169);
or U5293 (N_5293,N_5092,N_5163);
nor U5294 (N_5294,N_5236,N_5223);
and U5295 (N_5295,N_5104,N_5196);
and U5296 (N_5296,N_5195,N_5232);
and U5297 (N_5297,N_5197,N_5229);
or U5298 (N_5298,N_5212,N_5078);
nor U5299 (N_5299,N_5132,N_5051);
nor U5300 (N_5300,N_5224,N_5174);
nand U5301 (N_5301,N_5149,N_5164);
xnor U5302 (N_5302,N_5204,N_5128);
or U5303 (N_5303,N_5219,N_5033);
or U5304 (N_5304,N_5031,N_5209);
xnor U5305 (N_5305,N_5086,N_5044);
nand U5306 (N_5306,N_5084,N_5039);
nand U5307 (N_5307,N_5032,N_5162);
and U5308 (N_5308,N_5070,N_5075);
nand U5309 (N_5309,N_5180,N_5085);
or U5310 (N_5310,N_5109,N_5213);
xor U5311 (N_5311,N_5049,N_5211);
or U5312 (N_5312,N_5227,N_5160);
nand U5313 (N_5313,N_5079,N_5138);
xor U5314 (N_5314,N_5187,N_5036);
xnor U5315 (N_5315,N_5071,N_5061);
nand U5316 (N_5316,N_5159,N_5247);
nand U5317 (N_5317,N_5246,N_5140);
nor U5318 (N_5318,N_5010,N_5022);
xor U5319 (N_5319,N_5002,N_5106);
nand U5320 (N_5320,N_5139,N_5074);
and U5321 (N_5321,N_5116,N_5185);
xor U5322 (N_5322,N_5034,N_5102);
nand U5323 (N_5323,N_5024,N_5012);
or U5324 (N_5324,N_5046,N_5045);
or U5325 (N_5325,N_5242,N_5060);
or U5326 (N_5326,N_5217,N_5215);
and U5327 (N_5327,N_5234,N_5030);
or U5328 (N_5328,N_5062,N_5172);
and U5329 (N_5329,N_5088,N_5150);
nor U5330 (N_5330,N_5056,N_5161);
nand U5331 (N_5331,N_5158,N_5037);
nor U5332 (N_5332,N_5003,N_5201);
xor U5333 (N_5333,N_5054,N_5188);
or U5334 (N_5334,N_5081,N_5068);
or U5335 (N_5335,N_5101,N_5021);
nor U5336 (N_5336,N_5050,N_5129);
xnor U5337 (N_5337,N_5047,N_5216);
and U5338 (N_5338,N_5222,N_5103);
nor U5339 (N_5339,N_5199,N_5137);
nand U5340 (N_5340,N_5107,N_5018);
nand U5341 (N_5341,N_5228,N_5221);
nor U5342 (N_5342,N_5152,N_5202);
nand U5343 (N_5343,N_5191,N_5035);
nor U5344 (N_5344,N_5134,N_5156);
nand U5345 (N_5345,N_5245,N_5029);
nand U5346 (N_5346,N_5230,N_5017);
xor U5347 (N_5347,N_5094,N_5119);
xor U5348 (N_5348,N_5048,N_5175);
or U5349 (N_5349,N_5080,N_5108);
or U5350 (N_5350,N_5136,N_5028);
nand U5351 (N_5351,N_5123,N_5186);
nand U5352 (N_5352,N_5053,N_5177);
or U5353 (N_5353,N_5115,N_5192);
nand U5354 (N_5354,N_5135,N_5063);
or U5355 (N_5355,N_5146,N_5112);
and U5356 (N_5356,N_5206,N_5043);
and U5357 (N_5357,N_5167,N_5142);
xnor U5358 (N_5358,N_5182,N_5066);
nor U5359 (N_5359,N_5004,N_5189);
or U5360 (N_5360,N_5181,N_5057);
xnor U5361 (N_5361,N_5089,N_5058);
and U5362 (N_5362,N_5133,N_5168);
and U5363 (N_5363,N_5154,N_5153);
or U5364 (N_5364,N_5125,N_5001);
or U5365 (N_5365,N_5073,N_5226);
nand U5366 (N_5366,N_5239,N_5098);
nor U5367 (N_5367,N_5013,N_5077);
nor U5368 (N_5368,N_5096,N_5218);
or U5369 (N_5369,N_5171,N_5190);
nor U5370 (N_5370,N_5173,N_5111);
nor U5371 (N_5371,N_5009,N_5126);
nand U5372 (N_5372,N_5110,N_5113);
or U5373 (N_5373,N_5093,N_5059);
or U5374 (N_5374,N_5184,N_5100);
nand U5375 (N_5375,N_5128,N_5152);
xnor U5376 (N_5376,N_5214,N_5011);
or U5377 (N_5377,N_5204,N_5134);
nand U5378 (N_5378,N_5080,N_5117);
nor U5379 (N_5379,N_5162,N_5087);
xnor U5380 (N_5380,N_5173,N_5010);
and U5381 (N_5381,N_5229,N_5060);
nand U5382 (N_5382,N_5005,N_5136);
xor U5383 (N_5383,N_5013,N_5218);
xor U5384 (N_5384,N_5113,N_5177);
and U5385 (N_5385,N_5142,N_5164);
or U5386 (N_5386,N_5054,N_5000);
xnor U5387 (N_5387,N_5142,N_5035);
and U5388 (N_5388,N_5059,N_5167);
and U5389 (N_5389,N_5125,N_5185);
nor U5390 (N_5390,N_5153,N_5249);
nand U5391 (N_5391,N_5015,N_5156);
and U5392 (N_5392,N_5061,N_5126);
or U5393 (N_5393,N_5183,N_5130);
nand U5394 (N_5394,N_5120,N_5103);
nor U5395 (N_5395,N_5029,N_5116);
xnor U5396 (N_5396,N_5093,N_5146);
xnor U5397 (N_5397,N_5191,N_5140);
and U5398 (N_5398,N_5059,N_5235);
nand U5399 (N_5399,N_5218,N_5123);
xnor U5400 (N_5400,N_5232,N_5055);
nor U5401 (N_5401,N_5020,N_5197);
or U5402 (N_5402,N_5131,N_5154);
nor U5403 (N_5403,N_5107,N_5092);
nand U5404 (N_5404,N_5248,N_5191);
and U5405 (N_5405,N_5122,N_5069);
xor U5406 (N_5406,N_5110,N_5238);
or U5407 (N_5407,N_5234,N_5085);
xnor U5408 (N_5408,N_5105,N_5102);
nor U5409 (N_5409,N_5224,N_5062);
and U5410 (N_5410,N_5225,N_5200);
and U5411 (N_5411,N_5064,N_5104);
or U5412 (N_5412,N_5088,N_5165);
or U5413 (N_5413,N_5064,N_5248);
nand U5414 (N_5414,N_5199,N_5015);
or U5415 (N_5415,N_5086,N_5027);
nand U5416 (N_5416,N_5088,N_5092);
nor U5417 (N_5417,N_5194,N_5077);
nor U5418 (N_5418,N_5071,N_5217);
or U5419 (N_5419,N_5133,N_5169);
and U5420 (N_5420,N_5089,N_5104);
nor U5421 (N_5421,N_5018,N_5125);
nand U5422 (N_5422,N_5200,N_5165);
xnor U5423 (N_5423,N_5039,N_5025);
or U5424 (N_5424,N_5113,N_5155);
nand U5425 (N_5425,N_5243,N_5196);
and U5426 (N_5426,N_5202,N_5132);
xnor U5427 (N_5427,N_5219,N_5018);
and U5428 (N_5428,N_5030,N_5015);
or U5429 (N_5429,N_5156,N_5032);
nand U5430 (N_5430,N_5060,N_5160);
nor U5431 (N_5431,N_5187,N_5136);
xnor U5432 (N_5432,N_5221,N_5165);
xor U5433 (N_5433,N_5023,N_5038);
or U5434 (N_5434,N_5158,N_5099);
nor U5435 (N_5435,N_5189,N_5180);
nor U5436 (N_5436,N_5093,N_5015);
xor U5437 (N_5437,N_5013,N_5038);
xnor U5438 (N_5438,N_5231,N_5088);
and U5439 (N_5439,N_5154,N_5106);
nor U5440 (N_5440,N_5058,N_5108);
nor U5441 (N_5441,N_5047,N_5211);
xor U5442 (N_5442,N_5127,N_5131);
nor U5443 (N_5443,N_5158,N_5188);
nor U5444 (N_5444,N_5208,N_5218);
xnor U5445 (N_5445,N_5047,N_5193);
xnor U5446 (N_5446,N_5233,N_5048);
and U5447 (N_5447,N_5066,N_5056);
nor U5448 (N_5448,N_5047,N_5097);
or U5449 (N_5449,N_5209,N_5108);
and U5450 (N_5450,N_5173,N_5051);
and U5451 (N_5451,N_5155,N_5154);
and U5452 (N_5452,N_5118,N_5082);
or U5453 (N_5453,N_5217,N_5015);
and U5454 (N_5454,N_5221,N_5019);
xor U5455 (N_5455,N_5182,N_5026);
nor U5456 (N_5456,N_5018,N_5114);
or U5457 (N_5457,N_5207,N_5106);
nand U5458 (N_5458,N_5067,N_5174);
nand U5459 (N_5459,N_5087,N_5075);
and U5460 (N_5460,N_5197,N_5048);
xor U5461 (N_5461,N_5148,N_5239);
nand U5462 (N_5462,N_5237,N_5193);
nand U5463 (N_5463,N_5164,N_5095);
and U5464 (N_5464,N_5004,N_5027);
and U5465 (N_5465,N_5215,N_5031);
nand U5466 (N_5466,N_5171,N_5098);
or U5467 (N_5467,N_5199,N_5112);
xor U5468 (N_5468,N_5021,N_5105);
or U5469 (N_5469,N_5196,N_5061);
and U5470 (N_5470,N_5011,N_5064);
nand U5471 (N_5471,N_5070,N_5044);
or U5472 (N_5472,N_5081,N_5055);
nand U5473 (N_5473,N_5091,N_5019);
nand U5474 (N_5474,N_5165,N_5023);
nor U5475 (N_5475,N_5165,N_5019);
or U5476 (N_5476,N_5117,N_5103);
and U5477 (N_5477,N_5174,N_5117);
nand U5478 (N_5478,N_5106,N_5237);
and U5479 (N_5479,N_5238,N_5056);
xor U5480 (N_5480,N_5073,N_5044);
or U5481 (N_5481,N_5195,N_5093);
nand U5482 (N_5482,N_5152,N_5055);
xor U5483 (N_5483,N_5031,N_5237);
or U5484 (N_5484,N_5224,N_5244);
nor U5485 (N_5485,N_5148,N_5141);
nor U5486 (N_5486,N_5138,N_5235);
nand U5487 (N_5487,N_5029,N_5191);
nor U5488 (N_5488,N_5041,N_5175);
nor U5489 (N_5489,N_5004,N_5041);
and U5490 (N_5490,N_5160,N_5029);
and U5491 (N_5491,N_5041,N_5157);
xnor U5492 (N_5492,N_5242,N_5076);
and U5493 (N_5493,N_5074,N_5097);
nand U5494 (N_5494,N_5229,N_5032);
and U5495 (N_5495,N_5117,N_5110);
xor U5496 (N_5496,N_5056,N_5052);
and U5497 (N_5497,N_5098,N_5130);
and U5498 (N_5498,N_5053,N_5045);
or U5499 (N_5499,N_5000,N_5242);
or U5500 (N_5500,N_5480,N_5279);
nor U5501 (N_5501,N_5398,N_5306);
nor U5502 (N_5502,N_5460,N_5317);
and U5503 (N_5503,N_5369,N_5436);
nor U5504 (N_5504,N_5463,N_5324);
nor U5505 (N_5505,N_5293,N_5473);
xnor U5506 (N_5506,N_5377,N_5411);
xnor U5507 (N_5507,N_5419,N_5337);
nand U5508 (N_5508,N_5359,N_5255);
nor U5509 (N_5509,N_5310,N_5435);
and U5510 (N_5510,N_5385,N_5413);
and U5511 (N_5511,N_5472,N_5296);
xor U5512 (N_5512,N_5388,N_5394);
nor U5513 (N_5513,N_5384,N_5489);
nand U5514 (N_5514,N_5259,N_5260);
nand U5515 (N_5515,N_5499,N_5367);
nand U5516 (N_5516,N_5266,N_5361);
nor U5517 (N_5517,N_5358,N_5275);
nor U5518 (N_5518,N_5465,N_5481);
xnor U5519 (N_5519,N_5373,N_5360);
xnor U5520 (N_5520,N_5332,N_5378);
nor U5521 (N_5521,N_5458,N_5392);
xnor U5522 (N_5522,N_5366,N_5469);
and U5523 (N_5523,N_5300,N_5417);
nor U5524 (N_5524,N_5423,N_5298);
or U5525 (N_5525,N_5487,N_5406);
xor U5526 (N_5526,N_5280,N_5407);
nor U5527 (N_5527,N_5292,N_5386);
xor U5528 (N_5528,N_5431,N_5414);
nand U5529 (N_5529,N_5402,N_5250);
nor U5530 (N_5530,N_5405,N_5322);
xor U5531 (N_5531,N_5486,N_5420);
nor U5532 (N_5532,N_5331,N_5342);
xor U5533 (N_5533,N_5316,N_5273);
or U5534 (N_5534,N_5461,N_5440);
or U5535 (N_5535,N_5447,N_5395);
nor U5536 (N_5536,N_5299,N_5258);
and U5537 (N_5537,N_5430,N_5443);
nand U5538 (N_5538,N_5454,N_5383);
nand U5539 (N_5539,N_5329,N_5297);
nand U5540 (N_5540,N_5305,N_5446);
nand U5541 (N_5541,N_5401,N_5451);
xor U5542 (N_5542,N_5362,N_5294);
nand U5543 (N_5543,N_5415,N_5477);
nand U5544 (N_5544,N_5285,N_5380);
nand U5545 (N_5545,N_5277,N_5476);
nor U5546 (N_5546,N_5283,N_5326);
xnor U5547 (N_5547,N_5276,N_5301);
xor U5548 (N_5548,N_5488,N_5456);
xnor U5549 (N_5549,N_5320,N_5421);
xnor U5550 (N_5550,N_5475,N_5351);
xnor U5551 (N_5551,N_5271,N_5448);
nand U5552 (N_5552,N_5374,N_5341);
nand U5553 (N_5553,N_5496,N_5468);
nor U5554 (N_5554,N_5399,N_5453);
nor U5555 (N_5555,N_5335,N_5262);
or U5556 (N_5556,N_5495,N_5363);
xor U5557 (N_5557,N_5368,N_5343);
xor U5558 (N_5558,N_5340,N_5311);
nor U5559 (N_5559,N_5325,N_5330);
and U5560 (N_5560,N_5287,N_5349);
and U5561 (N_5561,N_5467,N_5295);
nor U5562 (N_5562,N_5483,N_5452);
or U5563 (N_5563,N_5408,N_5357);
xor U5564 (N_5564,N_5323,N_5432);
xnor U5565 (N_5565,N_5354,N_5434);
xnor U5566 (N_5566,N_5409,N_5444);
and U5567 (N_5567,N_5304,N_5410);
nor U5568 (N_5568,N_5286,N_5345);
nand U5569 (N_5569,N_5390,N_5485);
xnor U5570 (N_5570,N_5265,N_5284);
and U5571 (N_5571,N_5272,N_5381);
xor U5572 (N_5572,N_5313,N_5352);
and U5573 (N_5573,N_5397,N_5437);
xnor U5574 (N_5574,N_5338,N_5466);
or U5575 (N_5575,N_5427,N_5375);
nand U5576 (N_5576,N_5391,N_5334);
and U5577 (N_5577,N_5492,N_5319);
xnor U5578 (N_5578,N_5416,N_5382);
nor U5579 (N_5579,N_5470,N_5474);
nor U5580 (N_5580,N_5404,N_5387);
or U5581 (N_5581,N_5498,N_5424);
nor U5582 (N_5582,N_5425,N_5252);
and U5583 (N_5583,N_5493,N_5263);
and U5584 (N_5584,N_5318,N_5364);
nand U5585 (N_5585,N_5312,N_5457);
xnor U5586 (N_5586,N_5308,N_5471);
xnor U5587 (N_5587,N_5355,N_5251);
and U5588 (N_5588,N_5274,N_5288);
nor U5589 (N_5589,N_5339,N_5309);
nand U5590 (N_5590,N_5455,N_5356);
and U5591 (N_5591,N_5422,N_5433);
xnor U5592 (N_5592,N_5303,N_5261);
or U5593 (N_5593,N_5450,N_5281);
and U5594 (N_5594,N_5464,N_5438);
xor U5595 (N_5595,N_5462,N_5327);
nand U5596 (N_5596,N_5365,N_5257);
or U5597 (N_5597,N_5442,N_5479);
xnor U5598 (N_5598,N_5459,N_5441);
xnor U5599 (N_5599,N_5403,N_5346);
nand U5600 (N_5600,N_5291,N_5445);
or U5601 (N_5601,N_5268,N_5328);
or U5602 (N_5602,N_5321,N_5426);
and U5603 (N_5603,N_5302,N_5400);
nor U5604 (N_5604,N_5333,N_5267);
or U5605 (N_5605,N_5497,N_5484);
nor U5606 (N_5606,N_5379,N_5270);
nor U5607 (N_5607,N_5253,N_5307);
nand U5608 (N_5608,N_5269,N_5439);
nand U5609 (N_5609,N_5347,N_5336);
xnor U5610 (N_5610,N_5353,N_5482);
nand U5611 (N_5611,N_5344,N_5372);
or U5612 (N_5612,N_5289,N_5282);
or U5613 (N_5613,N_5490,N_5264);
nand U5614 (N_5614,N_5314,N_5376);
and U5615 (N_5615,N_5315,N_5290);
nor U5616 (N_5616,N_5412,N_5478);
nand U5617 (N_5617,N_5418,N_5254);
nor U5618 (N_5618,N_5494,N_5371);
xnor U5619 (N_5619,N_5393,N_5396);
or U5620 (N_5620,N_5428,N_5389);
nand U5621 (N_5621,N_5350,N_5256);
and U5622 (N_5622,N_5348,N_5278);
xnor U5623 (N_5623,N_5449,N_5429);
xor U5624 (N_5624,N_5370,N_5491);
nand U5625 (N_5625,N_5382,N_5492);
or U5626 (N_5626,N_5271,N_5462);
or U5627 (N_5627,N_5466,N_5350);
nor U5628 (N_5628,N_5307,N_5291);
xnor U5629 (N_5629,N_5379,N_5352);
or U5630 (N_5630,N_5464,N_5254);
nor U5631 (N_5631,N_5336,N_5441);
xnor U5632 (N_5632,N_5264,N_5463);
nand U5633 (N_5633,N_5443,N_5412);
xor U5634 (N_5634,N_5259,N_5326);
and U5635 (N_5635,N_5396,N_5476);
or U5636 (N_5636,N_5400,N_5419);
nand U5637 (N_5637,N_5491,N_5341);
or U5638 (N_5638,N_5402,N_5455);
nand U5639 (N_5639,N_5440,N_5324);
and U5640 (N_5640,N_5342,N_5420);
or U5641 (N_5641,N_5486,N_5450);
xor U5642 (N_5642,N_5257,N_5357);
xnor U5643 (N_5643,N_5275,N_5435);
or U5644 (N_5644,N_5453,N_5297);
xor U5645 (N_5645,N_5333,N_5424);
and U5646 (N_5646,N_5289,N_5312);
or U5647 (N_5647,N_5409,N_5428);
and U5648 (N_5648,N_5407,N_5467);
nor U5649 (N_5649,N_5297,N_5318);
xnor U5650 (N_5650,N_5358,N_5430);
or U5651 (N_5651,N_5312,N_5470);
xnor U5652 (N_5652,N_5399,N_5470);
nand U5653 (N_5653,N_5359,N_5459);
and U5654 (N_5654,N_5295,N_5383);
xor U5655 (N_5655,N_5481,N_5499);
and U5656 (N_5656,N_5379,N_5288);
or U5657 (N_5657,N_5354,N_5414);
xnor U5658 (N_5658,N_5307,N_5484);
and U5659 (N_5659,N_5418,N_5268);
nand U5660 (N_5660,N_5305,N_5377);
and U5661 (N_5661,N_5337,N_5460);
or U5662 (N_5662,N_5397,N_5428);
xor U5663 (N_5663,N_5473,N_5374);
nor U5664 (N_5664,N_5313,N_5287);
and U5665 (N_5665,N_5472,N_5447);
and U5666 (N_5666,N_5390,N_5458);
xor U5667 (N_5667,N_5390,N_5357);
and U5668 (N_5668,N_5299,N_5383);
and U5669 (N_5669,N_5435,N_5430);
xnor U5670 (N_5670,N_5402,N_5435);
or U5671 (N_5671,N_5291,N_5367);
nor U5672 (N_5672,N_5381,N_5327);
nand U5673 (N_5673,N_5411,N_5495);
and U5674 (N_5674,N_5342,N_5381);
and U5675 (N_5675,N_5332,N_5353);
nand U5676 (N_5676,N_5303,N_5495);
nand U5677 (N_5677,N_5390,N_5322);
nand U5678 (N_5678,N_5435,N_5458);
nand U5679 (N_5679,N_5458,N_5402);
nand U5680 (N_5680,N_5425,N_5450);
nor U5681 (N_5681,N_5422,N_5390);
or U5682 (N_5682,N_5288,N_5449);
nor U5683 (N_5683,N_5423,N_5378);
xor U5684 (N_5684,N_5392,N_5317);
nand U5685 (N_5685,N_5397,N_5290);
nand U5686 (N_5686,N_5447,N_5291);
nor U5687 (N_5687,N_5253,N_5347);
and U5688 (N_5688,N_5262,N_5339);
and U5689 (N_5689,N_5358,N_5435);
nand U5690 (N_5690,N_5439,N_5293);
nand U5691 (N_5691,N_5441,N_5349);
or U5692 (N_5692,N_5387,N_5367);
nand U5693 (N_5693,N_5301,N_5420);
nor U5694 (N_5694,N_5439,N_5386);
xor U5695 (N_5695,N_5257,N_5311);
nor U5696 (N_5696,N_5322,N_5289);
xor U5697 (N_5697,N_5470,N_5353);
or U5698 (N_5698,N_5431,N_5437);
or U5699 (N_5699,N_5493,N_5489);
nand U5700 (N_5700,N_5269,N_5392);
nor U5701 (N_5701,N_5268,N_5290);
nand U5702 (N_5702,N_5367,N_5410);
and U5703 (N_5703,N_5469,N_5281);
xor U5704 (N_5704,N_5444,N_5265);
xor U5705 (N_5705,N_5267,N_5440);
xor U5706 (N_5706,N_5309,N_5324);
nor U5707 (N_5707,N_5366,N_5322);
or U5708 (N_5708,N_5255,N_5329);
nand U5709 (N_5709,N_5494,N_5349);
xor U5710 (N_5710,N_5254,N_5318);
xnor U5711 (N_5711,N_5340,N_5482);
nand U5712 (N_5712,N_5435,N_5484);
nor U5713 (N_5713,N_5386,N_5257);
or U5714 (N_5714,N_5353,N_5460);
nand U5715 (N_5715,N_5489,N_5357);
nor U5716 (N_5716,N_5457,N_5354);
xnor U5717 (N_5717,N_5250,N_5268);
nor U5718 (N_5718,N_5253,N_5496);
xor U5719 (N_5719,N_5443,N_5396);
nor U5720 (N_5720,N_5326,N_5461);
xnor U5721 (N_5721,N_5267,N_5335);
or U5722 (N_5722,N_5382,N_5495);
nand U5723 (N_5723,N_5290,N_5429);
or U5724 (N_5724,N_5428,N_5419);
nor U5725 (N_5725,N_5413,N_5463);
nor U5726 (N_5726,N_5410,N_5423);
or U5727 (N_5727,N_5429,N_5412);
or U5728 (N_5728,N_5422,N_5449);
and U5729 (N_5729,N_5332,N_5443);
or U5730 (N_5730,N_5358,N_5250);
and U5731 (N_5731,N_5484,N_5282);
nor U5732 (N_5732,N_5357,N_5454);
and U5733 (N_5733,N_5268,N_5285);
and U5734 (N_5734,N_5364,N_5461);
or U5735 (N_5735,N_5334,N_5469);
nand U5736 (N_5736,N_5412,N_5469);
nand U5737 (N_5737,N_5470,N_5308);
nand U5738 (N_5738,N_5478,N_5278);
or U5739 (N_5739,N_5295,N_5476);
nor U5740 (N_5740,N_5499,N_5296);
nor U5741 (N_5741,N_5434,N_5298);
nor U5742 (N_5742,N_5306,N_5297);
and U5743 (N_5743,N_5300,N_5294);
and U5744 (N_5744,N_5280,N_5257);
or U5745 (N_5745,N_5439,N_5379);
xnor U5746 (N_5746,N_5307,N_5405);
nand U5747 (N_5747,N_5446,N_5387);
nor U5748 (N_5748,N_5416,N_5436);
or U5749 (N_5749,N_5384,N_5362);
and U5750 (N_5750,N_5681,N_5731);
and U5751 (N_5751,N_5601,N_5569);
nor U5752 (N_5752,N_5613,N_5512);
or U5753 (N_5753,N_5534,N_5561);
and U5754 (N_5754,N_5598,N_5684);
and U5755 (N_5755,N_5522,N_5573);
nand U5756 (N_5756,N_5640,N_5648);
xor U5757 (N_5757,N_5695,N_5609);
or U5758 (N_5758,N_5662,N_5585);
nor U5759 (N_5759,N_5541,N_5708);
nor U5760 (N_5760,N_5641,N_5603);
xnor U5761 (N_5761,N_5549,N_5700);
and U5762 (N_5762,N_5553,N_5679);
or U5763 (N_5763,N_5527,N_5721);
nor U5764 (N_5764,N_5545,N_5652);
xnor U5765 (N_5765,N_5654,N_5665);
nand U5766 (N_5766,N_5516,N_5574);
or U5767 (N_5767,N_5607,N_5659);
nor U5768 (N_5768,N_5529,N_5517);
and U5769 (N_5769,N_5515,N_5719);
nand U5770 (N_5770,N_5732,N_5745);
and U5771 (N_5771,N_5686,N_5507);
nand U5772 (N_5772,N_5744,N_5646);
nor U5773 (N_5773,N_5728,N_5670);
nor U5774 (N_5774,N_5502,N_5590);
nand U5775 (N_5775,N_5701,N_5581);
nor U5776 (N_5776,N_5589,N_5599);
or U5777 (N_5777,N_5558,N_5644);
nand U5778 (N_5778,N_5597,N_5666);
nor U5779 (N_5779,N_5693,N_5530);
nor U5780 (N_5780,N_5746,N_5632);
xnor U5781 (N_5781,N_5702,N_5595);
and U5782 (N_5782,N_5618,N_5559);
nand U5783 (N_5783,N_5657,N_5532);
nand U5784 (N_5784,N_5593,N_5658);
nor U5785 (N_5785,N_5564,N_5536);
xnor U5786 (N_5786,N_5544,N_5624);
xor U5787 (N_5787,N_5500,N_5735);
xnor U5788 (N_5788,N_5741,N_5738);
nand U5789 (N_5789,N_5661,N_5716);
or U5790 (N_5790,N_5503,N_5547);
xor U5791 (N_5791,N_5623,N_5672);
nand U5792 (N_5792,N_5637,N_5582);
or U5793 (N_5793,N_5694,N_5577);
or U5794 (N_5794,N_5629,N_5604);
or U5795 (N_5795,N_5718,N_5570);
or U5796 (N_5796,N_5696,N_5643);
and U5797 (N_5797,N_5625,N_5552);
and U5798 (N_5798,N_5705,N_5505);
xor U5799 (N_5799,N_5563,N_5578);
or U5800 (N_5800,N_5556,N_5683);
and U5801 (N_5801,N_5689,N_5636);
and U5802 (N_5802,N_5667,N_5656);
or U5803 (N_5803,N_5639,N_5733);
xnor U5804 (N_5804,N_5687,N_5592);
nand U5805 (N_5805,N_5523,N_5554);
and U5806 (N_5806,N_5680,N_5571);
nor U5807 (N_5807,N_5633,N_5566);
nor U5808 (N_5808,N_5538,N_5533);
xor U5809 (N_5809,N_5734,N_5596);
nor U5810 (N_5810,N_5727,N_5535);
and U5811 (N_5811,N_5676,N_5651);
nor U5812 (N_5812,N_5675,N_5707);
and U5813 (N_5813,N_5520,N_5551);
and U5814 (N_5814,N_5720,N_5740);
nand U5815 (N_5815,N_5514,N_5504);
xor U5816 (N_5816,N_5614,N_5717);
and U5817 (N_5817,N_5638,N_5587);
and U5818 (N_5818,N_5616,N_5671);
xnor U5819 (N_5819,N_5580,N_5749);
and U5820 (N_5820,N_5704,N_5560);
nor U5821 (N_5821,N_5612,N_5691);
and U5822 (N_5822,N_5736,N_5511);
or U5823 (N_5823,N_5678,N_5540);
and U5824 (N_5824,N_5711,N_5610);
or U5825 (N_5825,N_5508,N_5567);
nor U5826 (N_5826,N_5615,N_5631);
or U5827 (N_5827,N_5699,N_5660);
nand U5828 (N_5828,N_5521,N_5725);
and U5829 (N_5829,N_5748,N_5509);
or U5830 (N_5830,N_5579,N_5576);
and U5831 (N_5831,N_5747,N_5682);
nor U5832 (N_5832,N_5690,N_5605);
nor U5833 (N_5833,N_5621,N_5645);
nand U5834 (N_5834,N_5626,N_5739);
nand U5835 (N_5835,N_5594,N_5584);
or U5836 (N_5836,N_5557,N_5712);
nand U5837 (N_5837,N_5548,N_5531);
xnor U5838 (N_5838,N_5674,N_5519);
xnor U5839 (N_5839,N_5726,N_5600);
xor U5840 (N_5840,N_5526,N_5510);
nand U5841 (N_5841,N_5528,N_5642);
or U5842 (N_5842,N_5550,N_5542);
or U5843 (N_5843,N_5518,N_5630);
nand U5844 (N_5844,N_5685,N_5591);
xor U5845 (N_5845,N_5627,N_5714);
nor U5846 (N_5846,N_5663,N_5524);
nand U5847 (N_5847,N_5668,N_5664);
nor U5848 (N_5848,N_5724,N_5713);
nand U5849 (N_5849,N_5619,N_5655);
xor U5850 (N_5850,N_5647,N_5562);
xor U5851 (N_5851,N_5543,N_5617);
nor U5852 (N_5852,N_5635,N_5634);
and U5853 (N_5853,N_5698,N_5608);
xnor U5854 (N_5854,N_5688,N_5653);
nand U5855 (N_5855,N_5703,N_5730);
nand U5856 (N_5856,N_5715,N_5706);
nand U5857 (N_5857,N_5546,N_5677);
or U5858 (N_5858,N_5537,N_5649);
or U5859 (N_5859,N_5710,N_5628);
or U5860 (N_5860,N_5723,N_5565);
and U5861 (N_5861,N_5743,N_5692);
or U5862 (N_5862,N_5669,N_5709);
nand U5863 (N_5863,N_5697,N_5539);
xnor U5864 (N_5864,N_5742,N_5506);
xnor U5865 (N_5865,N_5568,N_5620);
nor U5866 (N_5866,N_5737,N_5622);
and U5867 (N_5867,N_5650,N_5583);
nand U5868 (N_5868,N_5673,N_5588);
xor U5869 (N_5869,N_5729,N_5606);
and U5870 (N_5870,N_5586,N_5722);
and U5871 (N_5871,N_5575,N_5525);
nor U5872 (N_5872,N_5611,N_5572);
and U5873 (N_5873,N_5555,N_5501);
xnor U5874 (N_5874,N_5513,N_5602);
xor U5875 (N_5875,N_5563,N_5635);
nand U5876 (N_5876,N_5649,N_5564);
nand U5877 (N_5877,N_5596,N_5580);
or U5878 (N_5878,N_5578,N_5542);
nor U5879 (N_5879,N_5529,N_5736);
nand U5880 (N_5880,N_5632,N_5713);
nor U5881 (N_5881,N_5616,N_5642);
or U5882 (N_5882,N_5589,N_5652);
nand U5883 (N_5883,N_5711,N_5647);
nand U5884 (N_5884,N_5707,N_5583);
and U5885 (N_5885,N_5598,N_5613);
or U5886 (N_5886,N_5695,N_5749);
and U5887 (N_5887,N_5555,N_5553);
nand U5888 (N_5888,N_5612,N_5613);
xnor U5889 (N_5889,N_5678,N_5562);
or U5890 (N_5890,N_5689,N_5542);
xnor U5891 (N_5891,N_5534,N_5615);
or U5892 (N_5892,N_5660,N_5719);
xnor U5893 (N_5893,N_5607,N_5564);
and U5894 (N_5894,N_5587,N_5578);
or U5895 (N_5895,N_5555,N_5748);
and U5896 (N_5896,N_5550,N_5731);
nor U5897 (N_5897,N_5509,N_5565);
nand U5898 (N_5898,N_5558,N_5718);
and U5899 (N_5899,N_5560,N_5588);
nor U5900 (N_5900,N_5711,N_5656);
or U5901 (N_5901,N_5646,N_5618);
nor U5902 (N_5902,N_5682,N_5644);
xnor U5903 (N_5903,N_5520,N_5729);
or U5904 (N_5904,N_5602,N_5712);
nor U5905 (N_5905,N_5637,N_5726);
or U5906 (N_5906,N_5605,N_5711);
nor U5907 (N_5907,N_5670,N_5562);
and U5908 (N_5908,N_5667,N_5583);
and U5909 (N_5909,N_5501,N_5744);
xnor U5910 (N_5910,N_5624,N_5702);
or U5911 (N_5911,N_5674,N_5616);
nor U5912 (N_5912,N_5684,N_5661);
and U5913 (N_5913,N_5593,N_5712);
xor U5914 (N_5914,N_5744,N_5599);
and U5915 (N_5915,N_5720,N_5556);
xor U5916 (N_5916,N_5572,N_5634);
xnor U5917 (N_5917,N_5624,N_5607);
and U5918 (N_5918,N_5705,N_5513);
nor U5919 (N_5919,N_5672,N_5683);
xor U5920 (N_5920,N_5735,N_5641);
or U5921 (N_5921,N_5551,N_5543);
or U5922 (N_5922,N_5514,N_5623);
and U5923 (N_5923,N_5602,N_5569);
and U5924 (N_5924,N_5748,N_5623);
or U5925 (N_5925,N_5667,N_5603);
and U5926 (N_5926,N_5509,N_5632);
and U5927 (N_5927,N_5647,N_5535);
nand U5928 (N_5928,N_5553,N_5623);
and U5929 (N_5929,N_5740,N_5525);
xnor U5930 (N_5930,N_5546,N_5649);
xnor U5931 (N_5931,N_5722,N_5524);
xor U5932 (N_5932,N_5652,N_5724);
xor U5933 (N_5933,N_5707,N_5502);
and U5934 (N_5934,N_5687,N_5501);
or U5935 (N_5935,N_5684,N_5536);
xnor U5936 (N_5936,N_5597,N_5615);
xnor U5937 (N_5937,N_5572,N_5710);
or U5938 (N_5938,N_5658,N_5699);
or U5939 (N_5939,N_5624,N_5525);
xor U5940 (N_5940,N_5668,N_5551);
and U5941 (N_5941,N_5606,N_5648);
nor U5942 (N_5942,N_5575,N_5511);
xor U5943 (N_5943,N_5638,N_5598);
and U5944 (N_5944,N_5620,N_5691);
and U5945 (N_5945,N_5551,N_5501);
nand U5946 (N_5946,N_5636,N_5665);
and U5947 (N_5947,N_5705,N_5515);
nor U5948 (N_5948,N_5562,N_5617);
nor U5949 (N_5949,N_5550,N_5562);
xor U5950 (N_5950,N_5604,N_5617);
nand U5951 (N_5951,N_5731,N_5687);
or U5952 (N_5952,N_5543,N_5672);
nor U5953 (N_5953,N_5721,N_5620);
nor U5954 (N_5954,N_5525,N_5683);
and U5955 (N_5955,N_5744,N_5526);
or U5956 (N_5956,N_5643,N_5707);
nor U5957 (N_5957,N_5545,N_5744);
nand U5958 (N_5958,N_5572,N_5601);
and U5959 (N_5959,N_5548,N_5500);
and U5960 (N_5960,N_5579,N_5596);
or U5961 (N_5961,N_5546,N_5556);
or U5962 (N_5962,N_5661,N_5745);
nand U5963 (N_5963,N_5568,N_5642);
and U5964 (N_5964,N_5640,N_5738);
nor U5965 (N_5965,N_5518,N_5735);
xnor U5966 (N_5966,N_5577,N_5711);
or U5967 (N_5967,N_5616,N_5648);
and U5968 (N_5968,N_5677,N_5560);
xor U5969 (N_5969,N_5516,N_5682);
xor U5970 (N_5970,N_5562,N_5566);
nand U5971 (N_5971,N_5726,N_5503);
or U5972 (N_5972,N_5725,N_5581);
xor U5973 (N_5973,N_5719,N_5538);
nor U5974 (N_5974,N_5693,N_5676);
nand U5975 (N_5975,N_5732,N_5586);
or U5976 (N_5976,N_5685,N_5635);
xor U5977 (N_5977,N_5726,N_5745);
and U5978 (N_5978,N_5749,N_5633);
nand U5979 (N_5979,N_5715,N_5628);
xnor U5980 (N_5980,N_5552,N_5501);
nand U5981 (N_5981,N_5618,N_5593);
or U5982 (N_5982,N_5651,N_5626);
nor U5983 (N_5983,N_5601,N_5587);
nor U5984 (N_5984,N_5652,N_5634);
nand U5985 (N_5985,N_5571,N_5648);
nor U5986 (N_5986,N_5558,N_5578);
nand U5987 (N_5987,N_5672,N_5574);
and U5988 (N_5988,N_5651,N_5679);
xnor U5989 (N_5989,N_5600,N_5674);
nand U5990 (N_5990,N_5681,N_5577);
xnor U5991 (N_5991,N_5587,N_5561);
xnor U5992 (N_5992,N_5656,N_5567);
nor U5993 (N_5993,N_5559,N_5696);
nor U5994 (N_5994,N_5531,N_5729);
nor U5995 (N_5995,N_5597,N_5685);
xor U5996 (N_5996,N_5592,N_5669);
and U5997 (N_5997,N_5676,N_5571);
nor U5998 (N_5998,N_5516,N_5551);
nor U5999 (N_5999,N_5675,N_5599);
xnor U6000 (N_6000,N_5961,N_5953);
xnor U6001 (N_6001,N_5956,N_5775);
or U6002 (N_6002,N_5812,N_5874);
nand U6003 (N_6003,N_5935,N_5912);
nand U6004 (N_6004,N_5862,N_5978);
or U6005 (N_6005,N_5921,N_5859);
or U6006 (N_6006,N_5801,N_5960);
and U6007 (N_6007,N_5815,N_5906);
and U6008 (N_6008,N_5922,N_5800);
nand U6009 (N_6009,N_5831,N_5780);
xnor U6010 (N_6010,N_5808,N_5883);
and U6011 (N_6011,N_5901,N_5911);
or U6012 (N_6012,N_5963,N_5943);
or U6013 (N_6013,N_5990,N_5931);
and U6014 (N_6014,N_5904,N_5849);
xnor U6015 (N_6015,N_5851,N_5798);
or U6016 (N_6016,N_5987,N_5973);
and U6017 (N_6017,N_5971,N_5794);
nor U6018 (N_6018,N_5942,N_5864);
and U6019 (N_6019,N_5882,N_5790);
nor U6020 (N_6020,N_5785,N_5970);
nor U6021 (N_6021,N_5755,N_5784);
and U6022 (N_6022,N_5880,N_5870);
nor U6023 (N_6023,N_5842,N_5934);
xor U6024 (N_6024,N_5804,N_5757);
and U6025 (N_6025,N_5892,N_5781);
nand U6026 (N_6026,N_5758,N_5772);
or U6027 (N_6027,N_5991,N_5827);
or U6028 (N_6028,N_5786,N_5825);
nand U6029 (N_6029,N_5795,N_5857);
and U6030 (N_6030,N_5760,N_5899);
nand U6031 (N_6031,N_5975,N_5951);
and U6032 (N_6032,N_5823,N_5998);
nor U6033 (N_6033,N_5944,N_5837);
and U6034 (N_6034,N_5791,N_5787);
and U6035 (N_6035,N_5872,N_5850);
nor U6036 (N_6036,N_5910,N_5806);
or U6037 (N_6037,N_5750,N_5796);
or U6038 (N_6038,N_5836,N_5923);
xnor U6039 (N_6039,N_5869,N_5832);
xor U6040 (N_6040,N_5926,N_5834);
nand U6041 (N_6041,N_5913,N_5879);
nand U6042 (N_6042,N_5939,N_5838);
nor U6043 (N_6043,N_5887,N_5845);
nand U6044 (N_6044,N_5949,N_5771);
xor U6045 (N_6045,N_5860,N_5875);
and U6046 (N_6046,N_5813,N_5829);
nand U6047 (N_6047,N_5828,N_5803);
xor U6048 (N_6048,N_5756,N_5855);
or U6049 (N_6049,N_5936,N_5843);
and U6050 (N_6050,N_5933,N_5778);
nand U6051 (N_6051,N_5995,N_5809);
xnor U6052 (N_6052,N_5927,N_5821);
xor U6053 (N_6053,N_5774,N_5788);
nand U6054 (N_6054,N_5988,N_5805);
nor U6055 (N_6055,N_5985,N_5969);
nor U6056 (N_6056,N_5903,N_5773);
nand U6057 (N_6057,N_5799,N_5884);
nor U6058 (N_6058,N_5908,N_5897);
nand U6059 (N_6059,N_5830,N_5852);
and U6060 (N_6060,N_5885,N_5776);
xor U6061 (N_6061,N_5810,N_5802);
and U6062 (N_6062,N_5958,N_5753);
nor U6063 (N_6063,N_5817,N_5811);
xnor U6064 (N_6064,N_5853,N_5950);
nor U6065 (N_6065,N_5766,N_5767);
nor U6066 (N_6066,N_5765,N_5962);
xnor U6067 (N_6067,N_5976,N_5881);
nor U6068 (N_6068,N_5866,N_5814);
nor U6069 (N_6069,N_5997,N_5972);
or U6070 (N_6070,N_5768,N_5863);
or U6071 (N_6071,N_5777,N_5977);
nand U6072 (N_6072,N_5994,N_5779);
xnor U6073 (N_6073,N_5986,N_5820);
nand U6074 (N_6074,N_5873,N_5981);
nor U6075 (N_6075,N_5854,N_5941);
xnor U6076 (N_6076,N_5751,N_5876);
and U6077 (N_6077,N_5856,N_5797);
nand U6078 (N_6078,N_5782,N_5848);
and U6079 (N_6079,N_5844,N_5819);
xnor U6080 (N_6080,N_5917,N_5871);
nor U6081 (N_6081,N_5920,N_5992);
and U6082 (N_6082,N_5763,N_5867);
nor U6083 (N_6083,N_5861,N_5916);
nand U6084 (N_6084,N_5930,N_5937);
xor U6085 (N_6085,N_5957,N_5764);
xnor U6086 (N_6086,N_5964,N_5816);
and U6087 (N_6087,N_5902,N_5974);
xor U6088 (N_6088,N_5979,N_5858);
xnor U6089 (N_6089,N_5919,N_5865);
and U6090 (N_6090,N_5952,N_5839);
and U6091 (N_6091,N_5868,N_5891);
nor U6092 (N_6092,N_5754,N_5993);
and U6093 (N_6093,N_5968,N_5841);
and U6094 (N_6094,N_5807,N_5761);
or U6095 (N_6095,N_5905,N_5955);
xnor U6096 (N_6096,N_5940,N_5762);
xor U6097 (N_6097,N_5954,N_5965);
xnor U6098 (N_6098,N_5890,N_5938);
xnor U6099 (N_6099,N_5929,N_5792);
and U6100 (N_6100,N_5984,N_5928);
or U6101 (N_6101,N_5886,N_5915);
xor U6102 (N_6102,N_5999,N_5983);
xnor U6103 (N_6103,N_5840,N_5980);
xor U6104 (N_6104,N_5966,N_5833);
xnor U6105 (N_6105,N_5877,N_5759);
nand U6106 (N_6106,N_5889,N_5996);
xor U6107 (N_6107,N_5925,N_5789);
or U6108 (N_6108,N_5900,N_5909);
nor U6109 (N_6109,N_5894,N_5895);
or U6110 (N_6110,N_5924,N_5822);
xor U6111 (N_6111,N_5826,N_5918);
or U6112 (N_6112,N_5959,N_5898);
nor U6113 (N_6113,N_5893,N_5989);
and U6114 (N_6114,N_5907,N_5932);
xnor U6115 (N_6115,N_5752,N_5770);
and U6116 (N_6116,N_5947,N_5946);
nand U6117 (N_6117,N_5888,N_5948);
nand U6118 (N_6118,N_5846,N_5835);
xnor U6119 (N_6119,N_5824,N_5914);
nand U6120 (N_6120,N_5878,N_5896);
and U6121 (N_6121,N_5945,N_5847);
and U6122 (N_6122,N_5793,N_5769);
xnor U6123 (N_6123,N_5818,N_5982);
nor U6124 (N_6124,N_5967,N_5783);
nor U6125 (N_6125,N_5985,N_5787);
nand U6126 (N_6126,N_5961,N_5791);
and U6127 (N_6127,N_5824,N_5866);
nor U6128 (N_6128,N_5804,N_5839);
or U6129 (N_6129,N_5911,N_5915);
or U6130 (N_6130,N_5771,N_5750);
and U6131 (N_6131,N_5889,N_5970);
nor U6132 (N_6132,N_5989,N_5906);
nor U6133 (N_6133,N_5912,N_5798);
nor U6134 (N_6134,N_5947,N_5948);
nand U6135 (N_6135,N_5780,N_5852);
xnor U6136 (N_6136,N_5948,N_5807);
or U6137 (N_6137,N_5764,N_5977);
nor U6138 (N_6138,N_5968,N_5895);
nor U6139 (N_6139,N_5922,N_5945);
nand U6140 (N_6140,N_5793,N_5962);
nor U6141 (N_6141,N_5944,N_5828);
or U6142 (N_6142,N_5851,N_5837);
or U6143 (N_6143,N_5934,N_5768);
nand U6144 (N_6144,N_5751,N_5986);
nor U6145 (N_6145,N_5823,N_5861);
and U6146 (N_6146,N_5765,N_5810);
xnor U6147 (N_6147,N_5804,N_5901);
and U6148 (N_6148,N_5838,N_5798);
nor U6149 (N_6149,N_5905,N_5920);
and U6150 (N_6150,N_5947,N_5949);
nor U6151 (N_6151,N_5959,N_5916);
nor U6152 (N_6152,N_5778,N_5777);
xor U6153 (N_6153,N_5844,N_5814);
or U6154 (N_6154,N_5920,N_5970);
nor U6155 (N_6155,N_5849,N_5984);
xnor U6156 (N_6156,N_5932,N_5892);
nor U6157 (N_6157,N_5983,N_5763);
nor U6158 (N_6158,N_5861,N_5909);
nor U6159 (N_6159,N_5759,N_5799);
nand U6160 (N_6160,N_5903,N_5899);
nor U6161 (N_6161,N_5970,N_5786);
and U6162 (N_6162,N_5909,N_5956);
and U6163 (N_6163,N_5867,N_5881);
or U6164 (N_6164,N_5809,N_5956);
and U6165 (N_6165,N_5770,N_5996);
and U6166 (N_6166,N_5787,N_5764);
nand U6167 (N_6167,N_5900,N_5791);
or U6168 (N_6168,N_5959,N_5754);
and U6169 (N_6169,N_5868,N_5906);
or U6170 (N_6170,N_5957,N_5797);
nand U6171 (N_6171,N_5848,N_5905);
nand U6172 (N_6172,N_5868,N_5950);
xor U6173 (N_6173,N_5954,N_5815);
and U6174 (N_6174,N_5953,N_5966);
or U6175 (N_6175,N_5938,N_5837);
nand U6176 (N_6176,N_5868,N_5804);
and U6177 (N_6177,N_5776,N_5994);
xor U6178 (N_6178,N_5983,N_5790);
nor U6179 (N_6179,N_5848,N_5934);
and U6180 (N_6180,N_5997,N_5968);
xor U6181 (N_6181,N_5807,N_5840);
nand U6182 (N_6182,N_5972,N_5953);
xnor U6183 (N_6183,N_5962,N_5784);
or U6184 (N_6184,N_5991,N_5917);
and U6185 (N_6185,N_5972,N_5804);
nor U6186 (N_6186,N_5996,N_5952);
nor U6187 (N_6187,N_5794,N_5942);
and U6188 (N_6188,N_5928,N_5856);
and U6189 (N_6189,N_5872,N_5821);
and U6190 (N_6190,N_5976,N_5788);
nor U6191 (N_6191,N_5956,N_5929);
nor U6192 (N_6192,N_5868,N_5867);
xnor U6193 (N_6193,N_5851,N_5985);
nand U6194 (N_6194,N_5828,N_5897);
nand U6195 (N_6195,N_5754,N_5780);
and U6196 (N_6196,N_5770,N_5884);
and U6197 (N_6197,N_5990,N_5773);
and U6198 (N_6198,N_5847,N_5764);
nor U6199 (N_6199,N_5949,N_5795);
and U6200 (N_6200,N_5980,N_5977);
or U6201 (N_6201,N_5852,N_5928);
nand U6202 (N_6202,N_5963,N_5885);
nor U6203 (N_6203,N_5764,N_5981);
nand U6204 (N_6204,N_5955,N_5992);
and U6205 (N_6205,N_5859,N_5881);
or U6206 (N_6206,N_5932,N_5952);
nand U6207 (N_6207,N_5940,N_5840);
nand U6208 (N_6208,N_5980,N_5850);
or U6209 (N_6209,N_5893,N_5836);
xnor U6210 (N_6210,N_5874,N_5796);
and U6211 (N_6211,N_5840,N_5966);
xor U6212 (N_6212,N_5805,N_5802);
xnor U6213 (N_6213,N_5811,N_5781);
nor U6214 (N_6214,N_5916,N_5999);
nor U6215 (N_6215,N_5771,N_5883);
xor U6216 (N_6216,N_5930,N_5894);
xor U6217 (N_6217,N_5847,N_5896);
xnor U6218 (N_6218,N_5923,N_5999);
or U6219 (N_6219,N_5919,N_5878);
or U6220 (N_6220,N_5921,N_5858);
or U6221 (N_6221,N_5785,N_5969);
or U6222 (N_6222,N_5932,N_5854);
and U6223 (N_6223,N_5782,N_5835);
nor U6224 (N_6224,N_5770,N_5851);
or U6225 (N_6225,N_5758,N_5912);
nor U6226 (N_6226,N_5840,N_5925);
xnor U6227 (N_6227,N_5992,N_5952);
xnor U6228 (N_6228,N_5918,N_5916);
or U6229 (N_6229,N_5796,N_5959);
or U6230 (N_6230,N_5766,N_5984);
nand U6231 (N_6231,N_5812,N_5969);
and U6232 (N_6232,N_5755,N_5993);
and U6233 (N_6233,N_5777,N_5863);
or U6234 (N_6234,N_5865,N_5825);
or U6235 (N_6235,N_5977,N_5892);
xnor U6236 (N_6236,N_5863,N_5996);
and U6237 (N_6237,N_5822,N_5813);
nor U6238 (N_6238,N_5960,N_5907);
and U6239 (N_6239,N_5884,N_5756);
or U6240 (N_6240,N_5961,N_5967);
and U6241 (N_6241,N_5801,N_5858);
nand U6242 (N_6242,N_5919,N_5869);
nor U6243 (N_6243,N_5865,N_5942);
or U6244 (N_6244,N_5933,N_5813);
xnor U6245 (N_6245,N_5761,N_5913);
or U6246 (N_6246,N_5794,N_5919);
and U6247 (N_6247,N_5915,N_5909);
nand U6248 (N_6248,N_5828,N_5895);
nand U6249 (N_6249,N_5891,N_5888);
nand U6250 (N_6250,N_6035,N_6024);
nand U6251 (N_6251,N_6169,N_6080);
nor U6252 (N_6252,N_6245,N_6060);
nor U6253 (N_6253,N_6020,N_6138);
xnor U6254 (N_6254,N_6010,N_6246);
or U6255 (N_6255,N_6063,N_6027);
nor U6256 (N_6256,N_6102,N_6036);
or U6257 (N_6257,N_6054,N_6176);
nor U6258 (N_6258,N_6047,N_6104);
nor U6259 (N_6259,N_6200,N_6195);
xnor U6260 (N_6260,N_6073,N_6199);
and U6261 (N_6261,N_6014,N_6099);
nor U6262 (N_6262,N_6235,N_6037);
nand U6263 (N_6263,N_6136,N_6057);
nor U6264 (N_6264,N_6107,N_6013);
nor U6265 (N_6265,N_6189,N_6091);
nor U6266 (N_6266,N_6053,N_6124);
and U6267 (N_6267,N_6148,N_6188);
and U6268 (N_6268,N_6103,N_6179);
xor U6269 (N_6269,N_6230,N_6227);
and U6270 (N_6270,N_6074,N_6117);
xnor U6271 (N_6271,N_6064,N_6134);
and U6272 (N_6272,N_6108,N_6133);
and U6273 (N_6273,N_6127,N_6056);
and U6274 (N_6274,N_6113,N_6183);
or U6275 (N_6275,N_6168,N_6070);
nor U6276 (N_6276,N_6210,N_6086);
and U6277 (N_6277,N_6238,N_6211);
xnor U6278 (N_6278,N_6129,N_6203);
nor U6279 (N_6279,N_6042,N_6198);
nor U6280 (N_6280,N_6118,N_6029);
or U6281 (N_6281,N_6193,N_6130);
or U6282 (N_6282,N_6110,N_6028);
nand U6283 (N_6283,N_6084,N_6039);
and U6284 (N_6284,N_6085,N_6007);
nand U6285 (N_6285,N_6098,N_6018);
and U6286 (N_6286,N_6165,N_6043);
and U6287 (N_6287,N_6159,N_6034);
nand U6288 (N_6288,N_6229,N_6213);
and U6289 (N_6289,N_6067,N_6212);
or U6290 (N_6290,N_6071,N_6019);
or U6291 (N_6291,N_6033,N_6061);
and U6292 (N_6292,N_6208,N_6106);
nand U6293 (N_6293,N_6248,N_6204);
xor U6294 (N_6294,N_6144,N_6224);
and U6295 (N_6295,N_6149,N_6012);
and U6296 (N_6296,N_6145,N_6160);
nor U6297 (N_6297,N_6236,N_6177);
xor U6298 (N_6298,N_6031,N_6146);
nor U6299 (N_6299,N_6194,N_6058);
nor U6300 (N_6300,N_6123,N_6231);
nand U6301 (N_6301,N_6017,N_6062);
or U6302 (N_6302,N_6178,N_6038);
nand U6303 (N_6303,N_6205,N_6202);
xor U6304 (N_6304,N_6240,N_6087);
or U6305 (N_6305,N_6089,N_6002);
nor U6306 (N_6306,N_6175,N_6082);
xnor U6307 (N_6307,N_6217,N_6097);
xnor U6308 (N_6308,N_6155,N_6090);
nand U6309 (N_6309,N_6164,N_6201);
xor U6310 (N_6310,N_6121,N_6030);
nand U6311 (N_6311,N_6192,N_6166);
and U6312 (N_6312,N_6100,N_6214);
xnor U6313 (N_6313,N_6125,N_6132);
nand U6314 (N_6314,N_6172,N_6190);
and U6315 (N_6315,N_6156,N_6044);
nand U6316 (N_6316,N_6109,N_6243);
and U6317 (N_6317,N_6112,N_6167);
nor U6318 (N_6318,N_6093,N_6218);
xnor U6319 (N_6319,N_6216,N_6120);
nor U6320 (N_6320,N_6055,N_6131);
or U6321 (N_6321,N_6000,N_6143);
nand U6322 (N_6322,N_6076,N_6242);
nor U6323 (N_6323,N_6069,N_6151);
or U6324 (N_6324,N_6048,N_6187);
xnor U6325 (N_6325,N_6225,N_6094);
or U6326 (N_6326,N_6185,N_6171);
nor U6327 (N_6327,N_6079,N_6157);
nand U6328 (N_6328,N_6158,N_6173);
nand U6329 (N_6329,N_6220,N_6186);
nand U6330 (N_6330,N_6050,N_6182);
or U6331 (N_6331,N_6081,N_6162);
nand U6332 (N_6332,N_6170,N_6105);
and U6333 (N_6333,N_6150,N_6226);
nor U6334 (N_6334,N_6249,N_6234);
or U6335 (N_6335,N_6068,N_6114);
and U6336 (N_6336,N_6009,N_6075);
or U6337 (N_6337,N_6241,N_6041);
and U6338 (N_6338,N_6021,N_6004);
and U6339 (N_6339,N_6119,N_6239);
or U6340 (N_6340,N_6152,N_6139);
xnor U6341 (N_6341,N_6046,N_6045);
nor U6342 (N_6342,N_6015,N_6059);
or U6343 (N_6343,N_6092,N_6008);
or U6344 (N_6344,N_6122,N_6161);
nor U6345 (N_6345,N_6244,N_6222);
xnor U6346 (N_6346,N_6101,N_6040);
or U6347 (N_6347,N_6181,N_6128);
xor U6348 (N_6348,N_6126,N_6072);
nand U6349 (N_6349,N_6215,N_6233);
nor U6350 (N_6350,N_6174,N_6016);
nand U6351 (N_6351,N_6232,N_6221);
and U6352 (N_6352,N_6025,N_6223);
nand U6353 (N_6353,N_6209,N_6196);
or U6354 (N_6354,N_6206,N_6111);
nand U6355 (N_6355,N_6078,N_6163);
nor U6356 (N_6356,N_6207,N_6077);
and U6357 (N_6357,N_6154,N_6247);
and U6358 (N_6358,N_6147,N_6153);
or U6359 (N_6359,N_6237,N_6066);
nor U6360 (N_6360,N_6228,N_6011);
or U6361 (N_6361,N_6180,N_6137);
nor U6362 (N_6362,N_6096,N_6191);
or U6363 (N_6363,N_6135,N_6219);
nor U6364 (N_6364,N_6049,N_6023);
and U6365 (N_6365,N_6083,N_6116);
xnor U6366 (N_6366,N_6197,N_6006);
nand U6367 (N_6367,N_6140,N_6051);
or U6368 (N_6368,N_6065,N_6032);
or U6369 (N_6369,N_6142,N_6115);
and U6370 (N_6370,N_6052,N_6005);
nor U6371 (N_6371,N_6022,N_6003);
and U6372 (N_6372,N_6095,N_6088);
nor U6373 (N_6373,N_6026,N_6141);
and U6374 (N_6374,N_6184,N_6001);
nand U6375 (N_6375,N_6194,N_6097);
nand U6376 (N_6376,N_6173,N_6222);
xnor U6377 (N_6377,N_6175,N_6144);
nand U6378 (N_6378,N_6018,N_6131);
nor U6379 (N_6379,N_6180,N_6135);
xor U6380 (N_6380,N_6002,N_6135);
nor U6381 (N_6381,N_6118,N_6156);
nor U6382 (N_6382,N_6083,N_6132);
nand U6383 (N_6383,N_6016,N_6136);
or U6384 (N_6384,N_6112,N_6023);
or U6385 (N_6385,N_6099,N_6053);
xnor U6386 (N_6386,N_6069,N_6248);
nor U6387 (N_6387,N_6235,N_6234);
xor U6388 (N_6388,N_6015,N_6011);
xor U6389 (N_6389,N_6074,N_6045);
xnor U6390 (N_6390,N_6214,N_6135);
or U6391 (N_6391,N_6184,N_6131);
xnor U6392 (N_6392,N_6095,N_6104);
or U6393 (N_6393,N_6067,N_6102);
xor U6394 (N_6394,N_6202,N_6197);
and U6395 (N_6395,N_6204,N_6030);
nor U6396 (N_6396,N_6083,N_6113);
and U6397 (N_6397,N_6116,N_6048);
nor U6398 (N_6398,N_6165,N_6202);
or U6399 (N_6399,N_6103,N_6011);
and U6400 (N_6400,N_6244,N_6154);
or U6401 (N_6401,N_6090,N_6086);
xor U6402 (N_6402,N_6186,N_6066);
or U6403 (N_6403,N_6136,N_6006);
xor U6404 (N_6404,N_6051,N_6208);
nor U6405 (N_6405,N_6072,N_6043);
xnor U6406 (N_6406,N_6147,N_6134);
nor U6407 (N_6407,N_6204,N_6116);
nor U6408 (N_6408,N_6073,N_6015);
or U6409 (N_6409,N_6189,N_6102);
xnor U6410 (N_6410,N_6008,N_6236);
nand U6411 (N_6411,N_6028,N_6038);
nor U6412 (N_6412,N_6221,N_6095);
nand U6413 (N_6413,N_6043,N_6157);
xor U6414 (N_6414,N_6127,N_6208);
nand U6415 (N_6415,N_6169,N_6182);
and U6416 (N_6416,N_6014,N_6064);
xor U6417 (N_6417,N_6062,N_6117);
or U6418 (N_6418,N_6098,N_6180);
xor U6419 (N_6419,N_6239,N_6234);
nand U6420 (N_6420,N_6211,N_6124);
nor U6421 (N_6421,N_6081,N_6056);
xnor U6422 (N_6422,N_6198,N_6080);
nand U6423 (N_6423,N_6134,N_6088);
and U6424 (N_6424,N_6015,N_6051);
or U6425 (N_6425,N_6149,N_6132);
xor U6426 (N_6426,N_6058,N_6146);
nor U6427 (N_6427,N_6099,N_6050);
xor U6428 (N_6428,N_6050,N_6008);
xor U6429 (N_6429,N_6024,N_6077);
xnor U6430 (N_6430,N_6233,N_6218);
nor U6431 (N_6431,N_6020,N_6240);
and U6432 (N_6432,N_6111,N_6055);
or U6433 (N_6433,N_6046,N_6152);
and U6434 (N_6434,N_6017,N_6170);
and U6435 (N_6435,N_6202,N_6041);
or U6436 (N_6436,N_6050,N_6180);
nand U6437 (N_6437,N_6102,N_6211);
nand U6438 (N_6438,N_6192,N_6093);
or U6439 (N_6439,N_6144,N_6054);
or U6440 (N_6440,N_6138,N_6187);
and U6441 (N_6441,N_6200,N_6005);
xor U6442 (N_6442,N_6055,N_6191);
or U6443 (N_6443,N_6139,N_6144);
or U6444 (N_6444,N_6231,N_6192);
xnor U6445 (N_6445,N_6142,N_6003);
or U6446 (N_6446,N_6138,N_6240);
or U6447 (N_6447,N_6178,N_6193);
xnor U6448 (N_6448,N_6100,N_6175);
or U6449 (N_6449,N_6021,N_6209);
and U6450 (N_6450,N_6135,N_6051);
or U6451 (N_6451,N_6029,N_6045);
and U6452 (N_6452,N_6164,N_6230);
or U6453 (N_6453,N_6100,N_6119);
nand U6454 (N_6454,N_6224,N_6218);
and U6455 (N_6455,N_6107,N_6126);
and U6456 (N_6456,N_6199,N_6075);
and U6457 (N_6457,N_6239,N_6095);
xor U6458 (N_6458,N_6219,N_6016);
nand U6459 (N_6459,N_6209,N_6109);
or U6460 (N_6460,N_6204,N_6154);
xnor U6461 (N_6461,N_6040,N_6218);
nand U6462 (N_6462,N_6157,N_6213);
nor U6463 (N_6463,N_6183,N_6074);
nand U6464 (N_6464,N_6110,N_6197);
nor U6465 (N_6465,N_6054,N_6136);
or U6466 (N_6466,N_6215,N_6078);
or U6467 (N_6467,N_6241,N_6019);
or U6468 (N_6468,N_6224,N_6024);
or U6469 (N_6469,N_6232,N_6029);
or U6470 (N_6470,N_6024,N_6062);
or U6471 (N_6471,N_6173,N_6050);
or U6472 (N_6472,N_6206,N_6062);
or U6473 (N_6473,N_6202,N_6069);
or U6474 (N_6474,N_6129,N_6152);
xor U6475 (N_6475,N_6012,N_6159);
or U6476 (N_6476,N_6180,N_6002);
or U6477 (N_6477,N_6054,N_6050);
or U6478 (N_6478,N_6190,N_6038);
nor U6479 (N_6479,N_6007,N_6038);
nor U6480 (N_6480,N_6118,N_6079);
and U6481 (N_6481,N_6013,N_6003);
or U6482 (N_6482,N_6062,N_6210);
and U6483 (N_6483,N_6168,N_6119);
or U6484 (N_6484,N_6207,N_6192);
nand U6485 (N_6485,N_6207,N_6210);
nand U6486 (N_6486,N_6221,N_6013);
or U6487 (N_6487,N_6065,N_6237);
and U6488 (N_6488,N_6127,N_6118);
and U6489 (N_6489,N_6179,N_6230);
xnor U6490 (N_6490,N_6215,N_6222);
and U6491 (N_6491,N_6176,N_6078);
xnor U6492 (N_6492,N_6211,N_6012);
or U6493 (N_6493,N_6217,N_6102);
nor U6494 (N_6494,N_6007,N_6122);
or U6495 (N_6495,N_6096,N_6181);
nor U6496 (N_6496,N_6041,N_6162);
or U6497 (N_6497,N_6142,N_6043);
xor U6498 (N_6498,N_6148,N_6055);
xnor U6499 (N_6499,N_6171,N_6216);
and U6500 (N_6500,N_6251,N_6275);
nand U6501 (N_6501,N_6285,N_6295);
or U6502 (N_6502,N_6305,N_6441);
and U6503 (N_6503,N_6298,N_6374);
or U6504 (N_6504,N_6420,N_6489);
xor U6505 (N_6505,N_6453,N_6299);
nor U6506 (N_6506,N_6437,N_6421);
nor U6507 (N_6507,N_6325,N_6381);
nand U6508 (N_6508,N_6485,N_6432);
or U6509 (N_6509,N_6266,N_6483);
xor U6510 (N_6510,N_6292,N_6418);
and U6511 (N_6511,N_6277,N_6486);
nor U6512 (N_6512,N_6480,N_6397);
and U6513 (N_6513,N_6326,N_6354);
or U6514 (N_6514,N_6372,N_6276);
nor U6515 (N_6515,N_6355,N_6384);
nor U6516 (N_6516,N_6308,N_6312);
and U6517 (N_6517,N_6368,N_6382);
nand U6518 (N_6518,N_6495,N_6461);
and U6519 (N_6519,N_6451,N_6423);
or U6520 (N_6520,N_6282,N_6329);
or U6521 (N_6521,N_6393,N_6405);
and U6522 (N_6522,N_6287,N_6466);
or U6523 (N_6523,N_6396,N_6264);
or U6524 (N_6524,N_6359,N_6265);
or U6525 (N_6525,N_6336,N_6296);
nand U6526 (N_6526,N_6400,N_6457);
and U6527 (N_6527,N_6255,N_6438);
and U6528 (N_6528,N_6452,N_6320);
or U6529 (N_6529,N_6449,N_6297);
nor U6530 (N_6530,N_6278,N_6450);
nor U6531 (N_6531,N_6318,N_6306);
xnor U6532 (N_6532,N_6410,N_6430);
nand U6533 (N_6533,N_6250,N_6256);
and U6534 (N_6534,N_6479,N_6447);
xnor U6535 (N_6535,N_6472,N_6484);
nor U6536 (N_6536,N_6362,N_6494);
nand U6537 (N_6537,N_6470,N_6402);
nand U6538 (N_6538,N_6401,N_6353);
and U6539 (N_6539,N_6390,N_6434);
nor U6540 (N_6540,N_6291,N_6375);
or U6541 (N_6541,N_6379,N_6414);
nand U6542 (N_6542,N_6398,N_6428);
nor U6543 (N_6543,N_6263,N_6476);
and U6544 (N_6544,N_6268,N_6411);
or U6545 (N_6545,N_6314,N_6464);
and U6546 (N_6546,N_6475,N_6334);
nor U6547 (N_6547,N_6459,N_6313);
nor U6548 (N_6548,N_6280,N_6377);
nand U6549 (N_6549,N_6339,N_6348);
xor U6550 (N_6550,N_6487,N_6433);
and U6551 (N_6551,N_6492,N_6253);
nor U6552 (N_6552,N_6272,N_6356);
or U6553 (N_6553,N_6462,N_6360);
nand U6554 (N_6554,N_6436,N_6262);
and U6555 (N_6555,N_6407,N_6482);
or U6556 (N_6556,N_6254,N_6286);
xnor U6557 (N_6557,N_6281,N_6274);
nor U6558 (N_6558,N_6269,N_6399);
or U6559 (N_6559,N_6271,N_6456);
nand U6560 (N_6560,N_6363,N_6454);
and U6561 (N_6561,N_6257,N_6311);
nand U6562 (N_6562,N_6419,N_6388);
and U6563 (N_6563,N_6303,N_6258);
nand U6564 (N_6564,N_6427,N_6370);
or U6565 (N_6565,N_6369,N_6367);
nand U6566 (N_6566,N_6469,N_6301);
nor U6567 (N_6567,N_6499,N_6378);
xnor U6568 (N_6568,N_6289,N_6424);
or U6569 (N_6569,N_6332,N_6488);
and U6570 (N_6570,N_6284,N_6273);
xor U6571 (N_6571,N_6394,N_6290);
and U6572 (N_6572,N_6321,N_6327);
nand U6573 (N_6573,N_6279,N_6358);
nand U6574 (N_6574,N_6365,N_6435);
nor U6575 (N_6575,N_6267,N_6490);
nor U6576 (N_6576,N_6352,N_6431);
or U6577 (N_6577,N_6309,N_6463);
xor U6578 (N_6578,N_6330,N_6448);
xor U6579 (N_6579,N_6404,N_6337);
xor U6580 (N_6580,N_6491,N_6371);
xor U6581 (N_6581,N_6455,N_6444);
and U6582 (N_6582,N_6304,N_6347);
and U6583 (N_6583,N_6425,N_6468);
nand U6584 (N_6584,N_6350,N_6366);
and U6585 (N_6585,N_6364,N_6345);
and U6586 (N_6586,N_6416,N_6260);
nand U6587 (N_6587,N_6252,N_6458);
xor U6588 (N_6588,N_6460,N_6440);
nand U6589 (N_6589,N_6387,N_6412);
xor U6590 (N_6590,N_6317,N_6323);
and U6591 (N_6591,N_6315,N_6391);
xnor U6592 (N_6592,N_6341,N_6288);
and U6593 (N_6593,N_6259,N_6413);
nor U6594 (N_6594,N_6471,N_6346);
or U6595 (N_6595,N_6392,N_6389);
xnor U6596 (N_6596,N_6328,N_6331);
nor U6597 (N_6597,N_6373,N_6349);
xor U6598 (N_6598,N_6409,N_6442);
nor U6599 (N_6599,N_6338,N_6351);
or U6600 (N_6600,N_6333,N_6498);
nor U6601 (N_6601,N_6294,N_6376);
or U6602 (N_6602,N_6403,N_6300);
and U6603 (N_6603,N_6322,N_6474);
xnor U6604 (N_6604,N_6385,N_6261);
xnor U6605 (N_6605,N_6283,N_6310);
xnor U6606 (N_6606,N_6383,N_6406);
nor U6607 (N_6607,N_6342,N_6429);
or U6608 (N_6608,N_6497,N_6344);
nor U6609 (N_6609,N_6324,N_6446);
or U6610 (N_6610,N_6496,N_6415);
or U6611 (N_6611,N_6439,N_6386);
nand U6612 (N_6612,N_6493,N_6293);
xor U6613 (N_6613,N_6467,N_6417);
xnor U6614 (N_6614,N_6340,N_6307);
xor U6615 (N_6615,N_6380,N_6361);
nand U6616 (N_6616,N_6477,N_6408);
nor U6617 (N_6617,N_6473,N_6443);
and U6618 (N_6618,N_6481,N_6465);
or U6619 (N_6619,N_6357,N_6335);
and U6620 (N_6620,N_6445,N_6316);
and U6621 (N_6621,N_6302,N_6422);
xor U6622 (N_6622,N_6343,N_6426);
and U6623 (N_6623,N_6395,N_6478);
nand U6624 (N_6624,N_6319,N_6270);
xor U6625 (N_6625,N_6286,N_6469);
nand U6626 (N_6626,N_6331,N_6402);
nor U6627 (N_6627,N_6365,N_6251);
and U6628 (N_6628,N_6348,N_6483);
xor U6629 (N_6629,N_6287,N_6325);
xnor U6630 (N_6630,N_6326,N_6411);
and U6631 (N_6631,N_6497,N_6408);
nor U6632 (N_6632,N_6440,N_6307);
nor U6633 (N_6633,N_6400,N_6435);
xnor U6634 (N_6634,N_6387,N_6298);
nor U6635 (N_6635,N_6310,N_6466);
xnor U6636 (N_6636,N_6250,N_6336);
xnor U6637 (N_6637,N_6307,N_6428);
and U6638 (N_6638,N_6300,N_6463);
nor U6639 (N_6639,N_6406,N_6367);
and U6640 (N_6640,N_6368,N_6362);
or U6641 (N_6641,N_6315,N_6483);
and U6642 (N_6642,N_6355,N_6434);
nor U6643 (N_6643,N_6499,N_6468);
xnor U6644 (N_6644,N_6379,N_6480);
nand U6645 (N_6645,N_6306,N_6328);
or U6646 (N_6646,N_6252,N_6469);
nand U6647 (N_6647,N_6330,N_6438);
xnor U6648 (N_6648,N_6286,N_6463);
or U6649 (N_6649,N_6406,N_6446);
and U6650 (N_6650,N_6304,N_6377);
xnor U6651 (N_6651,N_6337,N_6299);
nor U6652 (N_6652,N_6414,N_6312);
xnor U6653 (N_6653,N_6435,N_6465);
nor U6654 (N_6654,N_6296,N_6286);
or U6655 (N_6655,N_6391,N_6304);
or U6656 (N_6656,N_6336,N_6315);
xor U6657 (N_6657,N_6491,N_6280);
xnor U6658 (N_6658,N_6286,N_6486);
and U6659 (N_6659,N_6478,N_6495);
and U6660 (N_6660,N_6438,N_6388);
and U6661 (N_6661,N_6273,N_6436);
nor U6662 (N_6662,N_6281,N_6442);
or U6663 (N_6663,N_6308,N_6444);
nor U6664 (N_6664,N_6283,N_6397);
or U6665 (N_6665,N_6326,N_6449);
nand U6666 (N_6666,N_6311,N_6457);
nor U6667 (N_6667,N_6368,N_6435);
and U6668 (N_6668,N_6261,N_6281);
and U6669 (N_6669,N_6403,N_6450);
and U6670 (N_6670,N_6256,N_6474);
nor U6671 (N_6671,N_6362,N_6419);
nor U6672 (N_6672,N_6439,N_6457);
and U6673 (N_6673,N_6282,N_6413);
xnor U6674 (N_6674,N_6307,N_6492);
and U6675 (N_6675,N_6303,N_6466);
or U6676 (N_6676,N_6261,N_6362);
nand U6677 (N_6677,N_6443,N_6399);
and U6678 (N_6678,N_6396,N_6381);
nor U6679 (N_6679,N_6310,N_6366);
or U6680 (N_6680,N_6300,N_6433);
nand U6681 (N_6681,N_6489,N_6433);
nor U6682 (N_6682,N_6321,N_6423);
xor U6683 (N_6683,N_6251,N_6485);
nand U6684 (N_6684,N_6366,N_6499);
and U6685 (N_6685,N_6459,N_6411);
nor U6686 (N_6686,N_6373,N_6482);
or U6687 (N_6687,N_6357,N_6367);
and U6688 (N_6688,N_6429,N_6396);
nor U6689 (N_6689,N_6468,N_6387);
or U6690 (N_6690,N_6447,N_6481);
nand U6691 (N_6691,N_6439,N_6484);
or U6692 (N_6692,N_6312,N_6324);
nor U6693 (N_6693,N_6275,N_6259);
nand U6694 (N_6694,N_6426,N_6328);
xnor U6695 (N_6695,N_6292,N_6261);
nand U6696 (N_6696,N_6411,N_6458);
nand U6697 (N_6697,N_6497,N_6416);
nand U6698 (N_6698,N_6308,N_6353);
or U6699 (N_6699,N_6318,N_6474);
and U6700 (N_6700,N_6456,N_6304);
xor U6701 (N_6701,N_6373,N_6439);
nand U6702 (N_6702,N_6427,N_6280);
xor U6703 (N_6703,N_6319,N_6430);
or U6704 (N_6704,N_6362,N_6316);
nor U6705 (N_6705,N_6262,N_6398);
nor U6706 (N_6706,N_6414,N_6318);
nor U6707 (N_6707,N_6330,N_6291);
xor U6708 (N_6708,N_6425,N_6255);
and U6709 (N_6709,N_6342,N_6331);
nor U6710 (N_6710,N_6311,N_6327);
xor U6711 (N_6711,N_6300,N_6414);
xor U6712 (N_6712,N_6496,N_6349);
or U6713 (N_6713,N_6445,N_6283);
and U6714 (N_6714,N_6427,N_6372);
nand U6715 (N_6715,N_6276,N_6423);
nor U6716 (N_6716,N_6486,N_6491);
xnor U6717 (N_6717,N_6297,N_6496);
and U6718 (N_6718,N_6387,N_6380);
nand U6719 (N_6719,N_6399,N_6252);
or U6720 (N_6720,N_6391,N_6370);
nand U6721 (N_6721,N_6269,N_6351);
nor U6722 (N_6722,N_6390,N_6328);
nor U6723 (N_6723,N_6341,N_6457);
nor U6724 (N_6724,N_6484,N_6311);
nor U6725 (N_6725,N_6264,N_6420);
xnor U6726 (N_6726,N_6468,N_6380);
xnor U6727 (N_6727,N_6267,N_6299);
nand U6728 (N_6728,N_6452,N_6318);
and U6729 (N_6729,N_6371,N_6494);
and U6730 (N_6730,N_6480,N_6324);
nor U6731 (N_6731,N_6274,N_6309);
or U6732 (N_6732,N_6422,N_6263);
and U6733 (N_6733,N_6300,N_6424);
or U6734 (N_6734,N_6256,N_6416);
nor U6735 (N_6735,N_6405,N_6497);
xor U6736 (N_6736,N_6414,N_6485);
or U6737 (N_6737,N_6344,N_6375);
and U6738 (N_6738,N_6401,N_6323);
xnor U6739 (N_6739,N_6413,N_6312);
xnor U6740 (N_6740,N_6254,N_6389);
nand U6741 (N_6741,N_6460,N_6295);
and U6742 (N_6742,N_6444,N_6434);
xnor U6743 (N_6743,N_6456,N_6489);
or U6744 (N_6744,N_6353,N_6260);
and U6745 (N_6745,N_6294,N_6488);
and U6746 (N_6746,N_6256,N_6466);
xnor U6747 (N_6747,N_6383,N_6417);
and U6748 (N_6748,N_6413,N_6264);
nand U6749 (N_6749,N_6480,N_6272);
nand U6750 (N_6750,N_6617,N_6630);
xnor U6751 (N_6751,N_6669,N_6585);
xor U6752 (N_6752,N_6627,N_6736);
xor U6753 (N_6753,N_6650,N_6705);
or U6754 (N_6754,N_6599,N_6571);
and U6755 (N_6755,N_6634,N_6730);
or U6756 (N_6756,N_6653,N_6671);
and U6757 (N_6757,N_6636,N_6525);
and U6758 (N_6758,N_6731,N_6518);
or U6759 (N_6759,N_6555,N_6519);
xnor U6760 (N_6760,N_6664,N_6602);
or U6761 (N_6761,N_6714,N_6743);
nand U6762 (N_6762,N_6575,N_6741);
or U6763 (N_6763,N_6713,N_6722);
xnor U6764 (N_6764,N_6564,N_6594);
xor U6765 (N_6765,N_6694,N_6607);
or U6766 (N_6766,N_6689,N_6666);
nand U6767 (N_6767,N_6549,N_6582);
xnor U6768 (N_6768,N_6605,N_6560);
xor U6769 (N_6769,N_6572,N_6632);
xor U6770 (N_6770,N_6719,N_6576);
or U6771 (N_6771,N_6639,N_6744);
nand U6772 (N_6772,N_6547,N_6672);
or U6773 (N_6773,N_6701,N_6651);
nand U6774 (N_6774,N_6502,N_6723);
and U6775 (N_6775,N_6610,N_6558);
nand U6776 (N_6776,N_6531,N_6579);
or U6777 (N_6777,N_6727,N_6684);
and U6778 (N_6778,N_6643,N_6615);
nand U6779 (N_6779,N_6748,N_6539);
and U6780 (N_6780,N_6712,N_6516);
nand U6781 (N_6781,N_6633,N_6655);
nand U6782 (N_6782,N_6606,N_6552);
and U6783 (N_6783,N_6667,N_6526);
nand U6784 (N_6784,N_6604,N_6514);
nor U6785 (N_6785,N_6556,N_6640);
xnor U6786 (N_6786,N_6674,N_6749);
nor U6787 (N_6787,N_6698,N_6663);
nor U6788 (N_6788,N_6624,N_6532);
or U6789 (N_6789,N_6500,N_6670);
or U6790 (N_6790,N_6533,N_6535);
or U6791 (N_6791,N_6562,N_6520);
or U6792 (N_6792,N_6740,N_6563);
or U6793 (N_6793,N_6517,N_6692);
nor U6794 (N_6794,N_6746,N_6595);
xor U6795 (N_6795,N_6638,N_6676);
nand U6796 (N_6796,N_6534,N_6616);
xor U6797 (N_6797,N_6631,N_6561);
xnor U6798 (N_6798,N_6578,N_6551);
or U6799 (N_6799,N_6611,N_6721);
nor U6800 (N_6800,N_6512,N_6598);
nand U6801 (N_6801,N_6629,N_6681);
xor U6802 (N_6802,N_6662,N_6680);
and U6803 (N_6803,N_6695,N_6503);
and U6804 (N_6804,N_6589,N_6554);
and U6805 (N_6805,N_6691,N_6635);
nor U6806 (N_6806,N_6711,N_6718);
nand U6807 (N_6807,N_6577,N_6506);
nor U6808 (N_6808,N_6557,N_6726);
xnor U6809 (N_6809,N_6592,N_6702);
nand U6810 (N_6810,N_6528,N_6548);
and U6811 (N_6811,N_6536,N_6673);
xnor U6812 (N_6812,N_6515,N_6724);
xor U6813 (N_6813,N_6546,N_6679);
or U6814 (N_6814,N_6739,N_6693);
xnor U6815 (N_6815,N_6686,N_6742);
or U6816 (N_6816,N_6527,N_6593);
nand U6817 (N_6817,N_6618,N_6600);
or U6818 (N_6818,N_6745,N_6568);
nand U6819 (N_6819,N_6657,N_6541);
xnor U6820 (N_6820,N_6504,N_6696);
nand U6821 (N_6821,N_6675,N_6738);
nand U6822 (N_6822,N_6687,N_6603);
nand U6823 (N_6823,N_6507,N_6710);
or U6824 (N_6824,N_6737,N_6508);
xnor U6825 (N_6825,N_6647,N_6732);
nand U6826 (N_6826,N_6588,N_6580);
or U6827 (N_6827,N_6522,N_6747);
and U6828 (N_6828,N_6716,N_6637);
nor U6829 (N_6829,N_6553,N_6708);
and U6830 (N_6830,N_6682,N_6614);
and U6831 (N_6831,N_6537,N_6715);
nand U6832 (N_6832,N_6645,N_6609);
or U6833 (N_6833,N_6646,N_6725);
or U6834 (N_6834,N_6521,N_6626);
or U6835 (N_6835,N_6510,N_6658);
nor U6836 (N_6836,N_6612,N_6620);
nor U6837 (N_6837,N_6623,N_6613);
xor U6838 (N_6838,N_6591,N_6688);
nor U6839 (N_6839,N_6733,N_6720);
xor U6840 (N_6840,N_6540,N_6573);
or U6841 (N_6841,N_6567,N_6608);
xor U6842 (N_6842,N_6704,N_6513);
nand U6843 (N_6843,N_6735,N_6685);
or U6844 (N_6844,N_6717,N_6511);
nor U6845 (N_6845,N_6690,N_6734);
nand U6846 (N_6846,N_6501,N_6699);
nor U6847 (N_6847,N_6559,N_6574);
xor U6848 (N_6848,N_6706,N_6583);
or U6849 (N_6849,N_6703,N_6625);
or U6850 (N_6850,N_6709,N_6729);
and U6851 (N_6851,N_6545,N_6728);
xnor U6852 (N_6852,N_6581,N_6542);
or U6853 (N_6853,N_6707,N_6544);
nor U6854 (N_6854,N_6509,N_6524);
nor U6855 (N_6855,N_6530,N_6621);
or U6856 (N_6856,N_6697,N_6628);
or U6857 (N_6857,N_6622,N_6543);
or U6858 (N_6858,N_6590,N_6566);
xor U6859 (N_6859,N_6660,N_6678);
or U6860 (N_6860,N_6654,N_6586);
nand U6861 (N_6861,N_6649,N_6656);
or U6862 (N_6862,N_6601,N_6661);
xnor U6863 (N_6863,N_6683,N_6529);
xnor U6864 (N_6864,N_6565,N_6648);
nand U6865 (N_6865,N_6505,N_6569);
xnor U6866 (N_6866,N_6587,N_6597);
nand U6867 (N_6867,N_6700,N_6584);
or U6868 (N_6868,N_6619,N_6550);
xnor U6869 (N_6869,N_6668,N_6642);
and U6870 (N_6870,N_6665,N_6596);
and U6871 (N_6871,N_6641,N_6677);
xnor U6872 (N_6872,N_6659,N_6644);
xnor U6873 (N_6873,N_6538,N_6652);
and U6874 (N_6874,N_6570,N_6523);
nor U6875 (N_6875,N_6658,N_6640);
nor U6876 (N_6876,N_6712,N_6667);
nand U6877 (N_6877,N_6575,N_6647);
nor U6878 (N_6878,N_6516,N_6575);
xnor U6879 (N_6879,N_6688,N_6618);
and U6880 (N_6880,N_6501,N_6639);
xnor U6881 (N_6881,N_6702,N_6534);
xor U6882 (N_6882,N_6681,N_6670);
nor U6883 (N_6883,N_6713,N_6620);
and U6884 (N_6884,N_6667,N_6621);
nand U6885 (N_6885,N_6685,N_6694);
nor U6886 (N_6886,N_6542,N_6563);
nor U6887 (N_6887,N_6568,N_6666);
xor U6888 (N_6888,N_6518,N_6559);
nand U6889 (N_6889,N_6590,N_6620);
nand U6890 (N_6890,N_6642,N_6628);
or U6891 (N_6891,N_6553,N_6711);
and U6892 (N_6892,N_6687,N_6568);
or U6893 (N_6893,N_6673,N_6514);
and U6894 (N_6894,N_6681,N_6646);
nor U6895 (N_6895,N_6583,N_6520);
or U6896 (N_6896,N_6717,N_6682);
or U6897 (N_6897,N_6666,N_6515);
nor U6898 (N_6898,N_6692,N_6721);
and U6899 (N_6899,N_6542,N_6570);
nor U6900 (N_6900,N_6661,N_6548);
nand U6901 (N_6901,N_6579,N_6749);
or U6902 (N_6902,N_6594,N_6734);
or U6903 (N_6903,N_6681,N_6549);
or U6904 (N_6904,N_6653,N_6718);
nor U6905 (N_6905,N_6745,N_6554);
or U6906 (N_6906,N_6659,N_6672);
and U6907 (N_6907,N_6665,N_6675);
xor U6908 (N_6908,N_6669,N_6546);
nor U6909 (N_6909,N_6518,N_6736);
nand U6910 (N_6910,N_6552,N_6699);
and U6911 (N_6911,N_6726,N_6670);
and U6912 (N_6912,N_6714,N_6594);
xnor U6913 (N_6913,N_6554,N_6661);
or U6914 (N_6914,N_6691,N_6500);
or U6915 (N_6915,N_6747,N_6541);
or U6916 (N_6916,N_6515,N_6550);
and U6917 (N_6917,N_6661,N_6694);
nand U6918 (N_6918,N_6645,N_6701);
or U6919 (N_6919,N_6573,N_6506);
xnor U6920 (N_6920,N_6608,N_6715);
or U6921 (N_6921,N_6624,N_6620);
xnor U6922 (N_6922,N_6556,N_6540);
xor U6923 (N_6923,N_6743,N_6544);
and U6924 (N_6924,N_6742,N_6745);
xor U6925 (N_6925,N_6554,N_6587);
xnor U6926 (N_6926,N_6525,N_6711);
nand U6927 (N_6927,N_6684,N_6622);
and U6928 (N_6928,N_6678,N_6689);
and U6929 (N_6929,N_6718,N_6603);
nor U6930 (N_6930,N_6564,N_6727);
xnor U6931 (N_6931,N_6596,N_6526);
and U6932 (N_6932,N_6575,N_6611);
xnor U6933 (N_6933,N_6504,N_6628);
xnor U6934 (N_6934,N_6506,N_6539);
nand U6935 (N_6935,N_6719,N_6525);
nor U6936 (N_6936,N_6517,N_6553);
nand U6937 (N_6937,N_6542,N_6735);
and U6938 (N_6938,N_6500,N_6540);
xor U6939 (N_6939,N_6740,N_6594);
nor U6940 (N_6940,N_6748,N_6584);
nand U6941 (N_6941,N_6615,N_6635);
and U6942 (N_6942,N_6638,N_6646);
xnor U6943 (N_6943,N_6592,N_6591);
xnor U6944 (N_6944,N_6510,N_6518);
xnor U6945 (N_6945,N_6568,N_6549);
nand U6946 (N_6946,N_6678,N_6703);
xnor U6947 (N_6947,N_6575,N_6621);
nor U6948 (N_6948,N_6546,N_6569);
nand U6949 (N_6949,N_6544,N_6655);
nor U6950 (N_6950,N_6529,N_6534);
nand U6951 (N_6951,N_6741,N_6728);
and U6952 (N_6952,N_6618,N_6748);
nand U6953 (N_6953,N_6599,N_6686);
nand U6954 (N_6954,N_6697,N_6642);
or U6955 (N_6955,N_6541,N_6715);
and U6956 (N_6956,N_6616,N_6605);
nor U6957 (N_6957,N_6672,N_6668);
xnor U6958 (N_6958,N_6503,N_6659);
or U6959 (N_6959,N_6529,N_6695);
and U6960 (N_6960,N_6540,N_6699);
nand U6961 (N_6961,N_6573,N_6711);
or U6962 (N_6962,N_6667,N_6726);
and U6963 (N_6963,N_6738,N_6598);
xnor U6964 (N_6964,N_6528,N_6514);
xor U6965 (N_6965,N_6742,N_6530);
xor U6966 (N_6966,N_6528,N_6627);
xnor U6967 (N_6967,N_6604,N_6744);
and U6968 (N_6968,N_6604,N_6692);
and U6969 (N_6969,N_6641,N_6729);
nor U6970 (N_6970,N_6579,N_6734);
and U6971 (N_6971,N_6742,N_6510);
and U6972 (N_6972,N_6629,N_6514);
xor U6973 (N_6973,N_6567,N_6605);
xnor U6974 (N_6974,N_6707,N_6502);
nand U6975 (N_6975,N_6685,N_6729);
nand U6976 (N_6976,N_6628,N_6685);
nand U6977 (N_6977,N_6701,N_6646);
nand U6978 (N_6978,N_6697,N_6545);
or U6979 (N_6979,N_6610,N_6559);
nand U6980 (N_6980,N_6733,N_6686);
and U6981 (N_6981,N_6594,N_6666);
nand U6982 (N_6982,N_6543,N_6637);
or U6983 (N_6983,N_6652,N_6518);
xor U6984 (N_6984,N_6519,N_6668);
xor U6985 (N_6985,N_6725,N_6597);
xnor U6986 (N_6986,N_6700,N_6608);
or U6987 (N_6987,N_6687,N_6564);
nor U6988 (N_6988,N_6513,N_6599);
nand U6989 (N_6989,N_6645,N_6743);
or U6990 (N_6990,N_6504,N_6595);
and U6991 (N_6991,N_6714,N_6689);
and U6992 (N_6992,N_6737,N_6657);
xor U6993 (N_6993,N_6681,N_6590);
xnor U6994 (N_6994,N_6739,N_6575);
nor U6995 (N_6995,N_6578,N_6658);
and U6996 (N_6996,N_6584,N_6635);
nor U6997 (N_6997,N_6585,N_6717);
nand U6998 (N_6998,N_6743,N_6713);
xor U6999 (N_6999,N_6615,N_6695);
and U7000 (N_7000,N_6929,N_6964);
nand U7001 (N_7001,N_6957,N_6809);
and U7002 (N_7002,N_6870,N_6765);
or U7003 (N_7003,N_6879,N_6769);
nor U7004 (N_7004,N_6935,N_6807);
nand U7005 (N_7005,N_6992,N_6944);
xor U7006 (N_7006,N_6753,N_6886);
nor U7007 (N_7007,N_6919,N_6988);
nor U7008 (N_7008,N_6812,N_6789);
nand U7009 (N_7009,N_6810,N_6827);
xor U7010 (N_7010,N_6772,N_6797);
or U7011 (N_7011,N_6926,N_6760);
xnor U7012 (N_7012,N_6750,N_6984);
and U7013 (N_7013,N_6793,N_6791);
nor U7014 (N_7014,N_6841,N_6761);
nor U7015 (N_7015,N_6792,N_6854);
nor U7016 (N_7016,N_6806,N_6999);
nand U7017 (N_7017,N_6971,N_6861);
nor U7018 (N_7018,N_6853,N_6848);
or U7019 (N_7019,N_6826,N_6947);
or U7020 (N_7020,N_6986,N_6802);
xor U7021 (N_7021,N_6784,N_6990);
or U7022 (N_7022,N_6815,N_6909);
and U7023 (N_7023,N_6759,N_6887);
xor U7024 (N_7024,N_6950,N_6923);
xor U7025 (N_7025,N_6906,N_6951);
nor U7026 (N_7026,N_6920,N_6946);
nor U7027 (N_7027,N_6890,N_6832);
nand U7028 (N_7028,N_6775,N_6771);
xnor U7029 (N_7029,N_6875,N_6766);
or U7030 (N_7030,N_6777,N_6849);
nor U7031 (N_7031,N_6869,N_6911);
or U7032 (N_7032,N_6884,N_6788);
nor U7033 (N_7033,N_6994,N_6997);
nand U7034 (N_7034,N_6805,N_6872);
nand U7035 (N_7035,N_6939,N_6837);
and U7036 (N_7036,N_6758,N_6823);
nand U7037 (N_7037,N_6836,N_6995);
and U7038 (N_7038,N_6907,N_6843);
nor U7039 (N_7039,N_6770,N_6976);
xnor U7040 (N_7040,N_6891,N_6813);
nand U7041 (N_7041,N_6794,N_6779);
xnor U7042 (N_7042,N_6928,N_6897);
nand U7043 (N_7043,N_6780,N_6968);
xor U7044 (N_7044,N_6817,N_6859);
xor U7045 (N_7045,N_6961,N_6960);
and U7046 (N_7046,N_6931,N_6956);
nand U7047 (N_7047,N_6987,N_6844);
nand U7048 (N_7048,N_6889,N_6996);
and U7049 (N_7049,N_6851,N_6959);
nor U7050 (N_7050,N_6800,N_6916);
or U7051 (N_7051,N_6965,N_6894);
xnor U7052 (N_7052,N_6822,N_6940);
nand U7053 (N_7053,N_6821,N_6958);
xnor U7054 (N_7054,N_6852,N_6803);
xor U7055 (N_7055,N_6868,N_6764);
and U7056 (N_7056,N_6846,N_6795);
nor U7057 (N_7057,N_6828,N_6834);
xnor U7058 (N_7058,N_6966,N_6787);
and U7059 (N_7059,N_6902,N_6867);
nor U7060 (N_7060,N_6820,N_6838);
xor U7061 (N_7061,N_6754,N_6918);
or U7062 (N_7062,N_6901,N_6979);
and U7063 (N_7063,N_6782,N_6845);
or U7064 (N_7064,N_6858,N_6757);
and U7065 (N_7065,N_6924,N_6917);
nor U7066 (N_7066,N_6932,N_6967);
or U7067 (N_7067,N_6831,N_6899);
xnor U7068 (N_7068,N_6922,N_6840);
and U7069 (N_7069,N_6762,N_6989);
nor U7070 (N_7070,N_6808,N_6752);
or U7071 (N_7071,N_6895,N_6903);
nor U7072 (N_7072,N_6914,N_6991);
or U7073 (N_7073,N_6949,N_6880);
xor U7074 (N_7074,N_6892,N_6835);
and U7075 (N_7075,N_6921,N_6915);
xnor U7076 (N_7076,N_6755,N_6977);
or U7077 (N_7077,N_6927,N_6871);
nor U7078 (N_7078,N_6980,N_6814);
and U7079 (N_7079,N_6839,N_6930);
nor U7080 (N_7080,N_6978,N_6981);
nor U7081 (N_7081,N_6877,N_6860);
and U7082 (N_7082,N_6898,N_6774);
or U7083 (N_7083,N_6824,N_6882);
or U7084 (N_7084,N_6847,N_6819);
and U7085 (N_7085,N_6778,N_6799);
nand U7086 (N_7086,N_6955,N_6751);
or U7087 (N_7087,N_6982,N_6829);
xnor U7088 (N_7088,N_6876,N_6934);
nand U7089 (N_7089,N_6963,N_6796);
or U7090 (N_7090,N_6970,N_6904);
and U7091 (N_7091,N_6938,N_6865);
nor U7092 (N_7092,N_6900,N_6833);
nor U7093 (N_7093,N_6825,N_6790);
nand U7094 (N_7094,N_6972,N_6804);
and U7095 (N_7095,N_6786,N_6888);
nand U7096 (N_7096,N_6945,N_6767);
or U7097 (N_7097,N_6975,N_6811);
nand U7098 (N_7098,N_6842,N_6783);
xor U7099 (N_7099,N_6893,N_6856);
nand U7100 (N_7100,N_6905,N_6948);
or U7101 (N_7101,N_6941,N_6885);
nand U7102 (N_7102,N_6913,N_6974);
or U7103 (N_7103,N_6933,N_6763);
nor U7104 (N_7104,N_6862,N_6943);
or U7105 (N_7105,N_6925,N_6942);
and U7106 (N_7106,N_6768,N_6855);
nand U7107 (N_7107,N_6883,N_6818);
nand U7108 (N_7108,N_6969,N_6857);
nand U7109 (N_7109,N_6816,N_6954);
and U7110 (N_7110,N_6998,N_6936);
xnor U7111 (N_7111,N_6896,N_6756);
or U7112 (N_7112,N_6985,N_6773);
and U7113 (N_7113,N_6973,N_6781);
nand U7114 (N_7114,N_6952,N_6785);
nand U7115 (N_7115,N_6983,N_6910);
xnor U7116 (N_7116,N_6830,N_6962);
nor U7117 (N_7117,N_6850,N_6878);
nor U7118 (N_7118,N_6798,N_6864);
or U7119 (N_7119,N_6912,N_6881);
or U7120 (N_7120,N_6874,N_6908);
and U7121 (N_7121,N_6873,N_6866);
and U7122 (N_7122,N_6953,N_6993);
xor U7123 (N_7123,N_6863,N_6776);
and U7124 (N_7124,N_6937,N_6801);
nor U7125 (N_7125,N_6951,N_6789);
nand U7126 (N_7126,N_6959,N_6847);
or U7127 (N_7127,N_6805,N_6893);
nor U7128 (N_7128,N_6977,N_6911);
nand U7129 (N_7129,N_6785,N_6971);
nand U7130 (N_7130,N_6761,N_6935);
xor U7131 (N_7131,N_6933,N_6937);
xnor U7132 (N_7132,N_6982,N_6802);
and U7133 (N_7133,N_6822,N_6955);
xor U7134 (N_7134,N_6909,N_6995);
or U7135 (N_7135,N_6793,N_6889);
and U7136 (N_7136,N_6849,N_6984);
xnor U7137 (N_7137,N_6960,N_6987);
nand U7138 (N_7138,N_6833,N_6765);
or U7139 (N_7139,N_6785,N_6900);
and U7140 (N_7140,N_6830,N_6818);
xor U7141 (N_7141,N_6973,N_6861);
nor U7142 (N_7142,N_6949,N_6943);
xor U7143 (N_7143,N_6870,N_6975);
or U7144 (N_7144,N_6956,N_6846);
and U7145 (N_7145,N_6945,N_6878);
xnor U7146 (N_7146,N_6979,N_6912);
or U7147 (N_7147,N_6867,N_6877);
or U7148 (N_7148,N_6864,N_6832);
xor U7149 (N_7149,N_6962,N_6794);
nand U7150 (N_7150,N_6758,N_6877);
nand U7151 (N_7151,N_6868,N_6966);
and U7152 (N_7152,N_6904,N_6957);
or U7153 (N_7153,N_6762,N_6924);
nor U7154 (N_7154,N_6772,N_6751);
and U7155 (N_7155,N_6967,N_6799);
or U7156 (N_7156,N_6991,N_6976);
xor U7157 (N_7157,N_6888,N_6942);
and U7158 (N_7158,N_6897,N_6892);
nor U7159 (N_7159,N_6804,N_6924);
and U7160 (N_7160,N_6858,N_6896);
xnor U7161 (N_7161,N_6763,N_6780);
or U7162 (N_7162,N_6893,N_6757);
or U7163 (N_7163,N_6858,N_6913);
or U7164 (N_7164,N_6994,N_6756);
or U7165 (N_7165,N_6997,N_6905);
nor U7166 (N_7166,N_6854,N_6815);
xnor U7167 (N_7167,N_6870,N_6886);
or U7168 (N_7168,N_6813,N_6865);
xor U7169 (N_7169,N_6952,N_6915);
and U7170 (N_7170,N_6796,N_6942);
and U7171 (N_7171,N_6948,N_6953);
nand U7172 (N_7172,N_6751,N_6909);
nor U7173 (N_7173,N_6881,N_6849);
nand U7174 (N_7174,N_6870,N_6821);
and U7175 (N_7175,N_6996,N_6909);
and U7176 (N_7176,N_6804,N_6951);
nor U7177 (N_7177,N_6974,N_6979);
and U7178 (N_7178,N_6971,N_6915);
or U7179 (N_7179,N_6840,N_6847);
nor U7180 (N_7180,N_6929,N_6895);
xor U7181 (N_7181,N_6929,N_6957);
nor U7182 (N_7182,N_6784,N_6889);
and U7183 (N_7183,N_6993,N_6770);
nand U7184 (N_7184,N_6987,N_6962);
xnor U7185 (N_7185,N_6910,N_6979);
or U7186 (N_7186,N_6823,N_6858);
xor U7187 (N_7187,N_6984,N_6801);
and U7188 (N_7188,N_6836,N_6962);
xor U7189 (N_7189,N_6916,N_6963);
nor U7190 (N_7190,N_6944,N_6812);
nor U7191 (N_7191,N_6914,N_6948);
or U7192 (N_7192,N_6989,N_6903);
and U7193 (N_7193,N_6957,N_6980);
and U7194 (N_7194,N_6800,N_6988);
nor U7195 (N_7195,N_6761,N_6933);
nor U7196 (N_7196,N_6998,N_6974);
nor U7197 (N_7197,N_6871,N_6804);
xnor U7198 (N_7198,N_6873,N_6784);
xnor U7199 (N_7199,N_6863,N_6860);
nand U7200 (N_7200,N_6844,N_6806);
and U7201 (N_7201,N_6891,N_6981);
and U7202 (N_7202,N_6882,N_6903);
nor U7203 (N_7203,N_6863,N_6932);
or U7204 (N_7204,N_6812,N_6906);
and U7205 (N_7205,N_6812,N_6896);
nor U7206 (N_7206,N_6970,N_6808);
or U7207 (N_7207,N_6790,N_6887);
and U7208 (N_7208,N_6862,N_6796);
xor U7209 (N_7209,N_6844,N_6814);
nand U7210 (N_7210,N_6752,N_6943);
xnor U7211 (N_7211,N_6808,N_6996);
nand U7212 (N_7212,N_6799,N_6802);
or U7213 (N_7213,N_6988,N_6802);
and U7214 (N_7214,N_6814,N_6973);
xnor U7215 (N_7215,N_6939,N_6901);
xor U7216 (N_7216,N_6802,N_6969);
nand U7217 (N_7217,N_6887,N_6846);
and U7218 (N_7218,N_6971,N_6843);
xor U7219 (N_7219,N_6861,N_6815);
and U7220 (N_7220,N_6900,N_6832);
xnor U7221 (N_7221,N_6878,N_6821);
or U7222 (N_7222,N_6887,N_6894);
or U7223 (N_7223,N_6803,N_6850);
and U7224 (N_7224,N_6840,N_6855);
xor U7225 (N_7225,N_6998,N_6829);
or U7226 (N_7226,N_6964,N_6867);
or U7227 (N_7227,N_6884,N_6969);
nand U7228 (N_7228,N_6830,N_6758);
and U7229 (N_7229,N_6751,N_6865);
or U7230 (N_7230,N_6832,N_6819);
and U7231 (N_7231,N_6793,N_6945);
xnor U7232 (N_7232,N_6823,N_6886);
xnor U7233 (N_7233,N_6816,N_6814);
nor U7234 (N_7234,N_6796,N_6865);
or U7235 (N_7235,N_6750,N_6824);
nor U7236 (N_7236,N_6950,N_6844);
xnor U7237 (N_7237,N_6796,N_6765);
or U7238 (N_7238,N_6915,N_6767);
nor U7239 (N_7239,N_6962,N_6960);
nor U7240 (N_7240,N_6764,N_6950);
nand U7241 (N_7241,N_6770,N_6853);
nand U7242 (N_7242,N_6922,N_6755);
nor U7243 (N_7243,N_6887,N_6967);
and U7244 (N_7244,N_6842,N_6768);
nand U7245 (N_7245,N_6910,N_6765);
nor U7246 (N_7246,N_6993,N_6871);
xor U7247 (N_7247,N_6774,N_6931);
xnor U7248 (N_7248,N_6803,N_6805);
nand U7249 (N_7249,N_6814,N_6757);
and U7250 (N_7250,N_7106,N_7104);
or U7251 (N_7251,N_7172,N_7050);
xor U7252 (N_7252,N_7158,N_7100);
nor U7253 (N_7253,N_7135,N_7054);
nor U7254 (N_7254,N_7101,N_7161);
and U7255 (N_7255,N_7218,N_7208);
nor U7256 (N_7256,N_7030,N_7143);
nor U7257 (N_7257,N_7006,N_7204);
or U7258 (N_7258,N_7185,N_7011);
xnor U7259 (N_7259,N_7098,N_7159);
and U7260 (N_7260,N_7224,N_7141);
nand U7261 (N_7261,N_7035,N_7225);
or U7262 (N_7262,N_7083,N_7057);
and U7263 (N_7263,N_7007,N_7245);
and U7264 (N_7264,N_7013,N_7133);
nor U7265 (N_7265,N_7021,N_7240);
nor U7266 (N_7266,N_7226,N_7053);
nor U7267 (N_7267,N_7210,N_7125);
nor U7268 (N_7268,N_7191,N_7199);
nor U7269 (N_7269,N_7183,N_7156);
or U7270 (N_7270,N_7086,N_7154);
nor U7271 (N_7271,N_7081,N_7031);
nor U7272 (N_7272,N_7248,N_7150);
nand U7273 (N_7273,N_7008,N_7120);
nand U7274 (N_7274,N_7169,N_7058);
and U7275 (N_7275,N_7038,N_7062);
or U7276 (N_7276,N_7137,N_7134);
xor U7277 (N_7277,N_7155,N_7034);
nand U7278 (N_7278,N_7142,N_7138);
nor U7279 (N_7279,N_7244,N_7197);
nor U7280 (N_7280,N_7139,N_7052);
nand U7281 (N_7281,N_7063,N_7201);
xnor U7282 (N_7282,N_7099,N_7166);
nor U7283 (N_7283,N_7236,N_7109);
nand U7284 (N_7284,N_7198,N_7164);
xor U7285 (N_7285,N_7088,N_7193);
and U7286 (N_7286,N_7091,N_7069);
and U7287 (N_7287,N_7196,N_7033);
nand U7288 (N_7288,N_7115,N_7237);
nor U7289 (N_7289,N_7176,N_7149);
and U7290 (N_7290,N_7160,N_7130);
nor U7291 (N_7291,N_7174,N_7184);
nand U7292 (N_7292,N_7114,N_7206);
nor U7293 (N_7293,N_7005,N_7173);
or U7294 (N_7294,N_7020,N_7129);
or U7295 (N_7295,N_7107,N_7014);
nor U7296 (N_7296,N_7221,N_7162);
or U7297 (N_7297,N_7039,N_7077);
nand U7298 (N_7298,N_7064,N_7165);
and U7299 (N_7299,N_7093,N_7140);
xnor U7300 (N_7300,N_7222,N_7235);
or U7301 (N_7301,N_7178,N_7227);
nand U7302 (N_7302,N_7095,N_7232);
and U7303 (N_7303,N_7202,N_7131);
and U7304 (N_7304,N_7027,N_7238);
or U7305 (N_7305,N_7118,N_7096);
nor U7306 (N_7306,N_7084,N_7042);
and U7307 (N_7307,N_7068,N_7200);
or U7308 (N_7308,N_7016,N_7059);
nand U7309 (N_7309,N_7079,N_7103);
xor U7310 (N_7310,N_7110,N_7246);
nand U7311 (N_7311,N_7239,N_7056);
or U7312 (N_7312,N_7070,N_7074);
or U7313 (N_7313,N_7217,N_7180);
xor U7314 (N_7314,N_7076,N_7182);
or U7315 (N_7315,N_7247,N_7010);
or U7316 (N_7316,N_7157,N_7085);
or U7317 (N_7317,N_7051,N_7177);
or U7318 (N_7318,N_7097,N_7209);
or U7319 (N_7319,N_7094,N_7188);
xnor U7320 (N_7320,N_7080,N_7044);
xor U7321 (N_7321,N_7168,N_7211);
and U7322 (N_7322,N_7040,N_7117);
or U7323 (N_7323,N_7127,N_7049);
or U7324 (N_7324,N_7144,N_7223);
or U7325 (N_7325,N_7065,N_7102);
xnor U7326 (N_7326,N_7151,N_7136);
xor U7327 (N_7327,N_7075,N_7009);
nor U7328 (N_7328,N_7055,N_7214);
nor U7329 (N_7329,N_7229,N_7195);
nand U7330 (N_7330,N_7167,N_7181);
nor U7331 (N_7331,N_7028,N_7041);
or U7332 (N_7332,N_7219,N_7171);
and U7333 (N_7333,N_7153,N_7243);
nand U7334 (N_7334,N_7124,N_7216);
nand U7335 (N_7335,N_7128,N_7190);
nand U7336 (N_7336,N_7192,N_7152);
or U7337 (N_7337,N_7163,N_7090);
xnor U7338 (N_7338,N_7022,N_7105);
nor U7339 (N_7339,N_7024,N_7126);
and U7340 (N_7340,N_7148,N_7003);
nand U7341 (N_7341,N_7203,N_7002);
nand U7342 (N_7342,N_7072,N_7233);
nor U7343 (N_7343,N_7170,N_7078);
xor U7344 (N_7344,N_7234,N_7228);
nand U7345 (N_7345,N_7045,N_7205);
and U7346 (N_7346,N_7186,N_7231);
nor U7347 (N_7347,N_7037,N_7123);
xor U7348 (N_7348,N_7018,N_7089);
or U7349 (N_7349,N_7046,N_7121);
or U7350 (N_7350,N_7215,N_7061);
nand U7351 (N_7351,N_7249,N_7146);
and U7352 (N_7352,N_7119,N_7189);
nand U7353 (N_7353,N_7017,N_7000);
xnor U7354 (N_7354,N_7015,N_7012);
and U7355 (N_7355,N_7147,N_7113);
nand U7356 (N_7356,N_7019,N_7087);
nand U7357 (N_7357,N_7066,N_7029);
xor U7358 (N_7358,N_7145,N_7047);
and U7359 (N_7359,N_7111,N_7179);
or U7360 (N_7360,N_7067,N_7213);
nand U7361 (N_7361,N_7043,N_7108);
xor U7362 (N_7362,N_7025,N_7048);
or U7363 (N_7363,N_7220,N_7230);
or U7364 (N_7364,N_7207,N_7001);
or U7365 (N_7365,N_7092,N_7023);
nand U7366 (N_7366,N_7212,N_7032);
and U7367 (N_7367,N_7132,N_7082);
nand U7368 (N_7368,N_7073,N_7241);
nor U7369 (N_7369,N_7116,N_7242);
and U7370 (N_7370,N_7004,N_7036);
nand U7371 (N_7371,N_7175,N_7112);
nor U7372 (N_7372,N_7026,N_7060);
nor U7373 (N_7373,N_7194,N_7187);
or U7374 (N_7374,N_7071,N_7122);
xnor U7375 (N_7375,N_7129,N_7057);
xor U7376 (N_7376,N_7235,N_7233);
and U7377 (N_7377,N_7202,N_7066);
xor U7378 (N_7378,N_7099,N_7006);
nor U7379 (N_7379,N_7226,N_7001);
or U7380 (N_7380,N_7223,N_7041);
or U7381 (N_7381,N_7064,N_7189);
nand U7382 (N_7382,N_7211,N_7149);
xor U7383 (N_7383,N_7168,N_7223);
and U7384 (N_7384,N_7010,N_7039);
xor U7385 (N_7385,N_7016,N_7240);
or U7386 (N_7386,N_7070,N_7009);
and U7387 (N_7387,N_7246,N_7183);
or U7388 (N_7388,N_7057,N_7179);
nand U7389 (N_7389,N_7092,N_7210);
nand U7390 (N_7390,N_7207,N_7006);
nor U7391 (N_7391,N_7242,N_7113);
or U7392 (N_7392,N_7039,N_7029);
xnor U7393 (N_7393,N_7139,N_7099);
nor U7394 (N_7394,N_7155,N_7126);
nand U7395 (N_7395,N_7211,N_7174);
nor U7396 (N_7396,N_7017,N_7164);
xor U7397 (N_7397,N_7173,N_7136);
xnor U7398 (N_7398,N_7140,N_7077);
nand U7399 (N_7399,N_7165,N_7162);
xnor U7400 (N_7400,N_7193,N_7121);
or U7401 (N_7401,N_7232,N_7190);
xor U7402 (N_7402,N_7065,N_7196);
and U7403 (N_7403,N_7248,N_7098);
or U7404 (N_7404,N_7083,N_7195);
nor U7405 (N_7405,N_7189,N_7091);
nor U7406 (N_7406,N_7036,N_7186);
or U7407 (N_7407,N_7071,N_7202);
nor U7408 (N_7408,N_7211,N_7109);
and U7409 (N_7409,N_7062,N_7101);
and U7410 (N_7410,N_7178,N_7019);
xnor U7411 (N_7411,N_7193,N_7161);
nor U7412 (N_7412,N_7114,N_7170);
nand U7413 (N_7413,N_7163,N_7158);
or U7414 (N_7414,N_7101,N_7239);
nor U7415 (N_7415,N_7061,N_7123);
or U7416 (N_7416,N_7088,N_7046);
and U7417 (N_7417,N_7209,N_7238);
xnor U7418 (N_7418,N_7178,N_7115);
nand U7419 (N_7419,N_7107,N_7042);
nand U7420 (N_7420,N_7207,N_7053);
xor U7421 (N_7421,N_7158,N_7187);
xor U7422 (N_7422,N_7000,N_7138);
or U7423 (N_7423,N_7222,N_7027);
nor U7424 (N_7424,N_7053,N_7008);
nand U7425 (N_7425,N_7170,N_7196);
or U7426 (N_7426,N_7086,N_7164);
and U7427 (N_7427,N_7127,N_7167);
nand U7428 (N_7428,N_7209,N_7099);
and U7429 (N_7429,N_7053,N_7166);
and U7430 (N_7430,N_7004,N_7137);
and U7431 (N_7431,N_7160,N_7179);
or U7432 (N_7432,N_7084,N_7040);
or U7433 (N_7433,N_7208,N_7223);
nor U7434 (N_7434,N_7204,N_7078);
nand U7435 (N_7435,N_7108,N_7085);
or U7436 (N_7436,N_7154,N_7167);
xnor U7437 (N_7437,N_7021,N_7067);
nand U7438 (N_7438,N_7144,N_7090);
nand U7439 (N_7439,N_7101,N_7043);
nor U7440 (N_7440,N_7078,N_7201);
or U7441 (N_7441,N_7175,N_7061);
nor U7442 (N_7442,N_7170,N_7026);
nor U7443 (N_7443,N_7240,N_7161);
xor U7444 (N_7444,N_7082,N_7174);
or U7445 (N_7445,N_7142,N_7184);
nand U7446 (N_7446,N_7041,N_7235);
and U7447 (N_7447,N_7066,N_7027);
or U7448 (N_7448,N_7171,N_7212);
nor U7449 (N_7449,N_7130,N_7243);
nor U7450 (N_7450,N_7213,N_7191);
and U7451 (N_7451,N_7137,N_7120);
xor U7452 (N_7452,N_7159,N_7029);
nand U7453 (N_7453,N_7148,N_7238);
nor U7454 (N_7454,N_7021,N_7198);
or U7455 (N_7455,N_7078,N_7007);
xnor U7456 (N_7456,N_7141,N_7215);
and U7457 (N_7457,N_7210,N_7155);
and U7458 (N_7458,N_7021,N_7119);
nand U7459 (N_7459,N_7120,N_7247);
or U7460 (N_7460,N_7077,N_7088);
xor U7461 (N_7461,N_7221,N_7242);
nor U7462 (N_7462,N_7085,N_7064);
or U7463 (N_7463,N_7187,N_7123);
and U7464 (N_7464,N_7092,N_7021);
nor U7465 (N_7465,N_7124,N_7241);
nor U7466 (N_7466,N_7074,N_7135);
and U7467 (N_7467,N_7088,N_7054);
xor U7468 (N_7468,N_7239,N_7022);
nand U7469 (N_7469,N_7149,N_7033);
nand U7470 (N_7470,N_7051,N_7124);
nand U7471 (N_7471,N_7035,N_7219);
and U7472 (N_7472,N_7048,N_7003);
and U7473 (N_7473,N_7122,N_7046);
xnor U7474 (N_7474,N_7117,N_7153);
nand U7475 (N_7475,N_7092,N_7192);
and U7476 (N_7476,N_7186,N_7200);
or U7477 (N_7477,N_7047,N_7095);
xnor U7478 (N_7478,N_7000,N_7159);
nor U7479 (N_7479,N_7229,N_7113);
and U7480 (N_7480,N_7225,N_7055);
and U7481 (N_7481,N_7154,N_7163);
nand U7482 (N_7482,N_7038,N_7057);
nand U7483 (N_7483,N_7062,N_7247);
or U7484 (N_7484,N_7242,N_7182);
nor U7485 (N_7485,N_7180,N_7189);
or U7486 (N_7486,N_7208,N_7241);
and U7487 (N_7487,N_7185,N_7148);
nand U7488 (N_7488,N_7245,N_7092);
nor U7489 (N_7489,N_7165,N_7006);
nand U7490 (N_7490,N_7161,N_7244);
nand U7491 (N_7491,N_7247,N_7171);
nand U7492 (N_7492,N_7086,N_7018);
nor U7493 (N_7493,N_7092,N_7100);
xnor U7494 (N_7494,N_7216,N_7028);
nor U7495 (N_7495,N_7046,N_7160);
nor U7496 (N_7496,N_7125,N_7025);
nor U7497 (N_7497,N_7052,N_7150);
nor U7498 (N_7498,N_7063,N_7089);
nor U7499 (N_7499,N_7135,N_7200);
xnor U7500 (N_7500,N_7408,N_7413);
nand U7501 (N_7501,N_7466,N_7252);
nor U7502 (N_7502,N_7419,N_7324);
or U7503 (N_7503,N_7457,N_7328);
xnor U7504 (N_7504,N_7436,N_7311);
nor U7505 (N_7505,N_7287,N_7274);
or U7506 (N_7506,N_7381,N_7327);
nand U7507 (N_7507,N_7367,N_7269);
nand U7508 (N_7508,N_7499,N_7319);
and U7509 (N_7509,N_7388,N_7470);
xor U7510 (N_7510,N_7437,N_7478);
nor U7511 (N_7511,N_7486,N_7275);
xor U7512 (N_7512,N_7348,N_7286);
xor U7513 (N_7513,N_7268,N_7317);
nand U7514 (N_7514,N_7353,N_7409);
nor U7515 (N_7515,N_7488,N_7341);
and U7516 (N_7516,N_7318,N_7435);
nor U7517 (N_7517,N_7425,N_7359);
xor U7518 (N_7518,N_7471,N_7371);
nand U7519 (N_7519,N_7451,N_7309);
and U7520 (N_7520,N_7326,N_7279);
xor U7521 (N_7521,N_7422,N_7360);
or U7522 (N_7522,N_7362,N_7494);
nor U7523 (N_7523,N_7391,N_7469);
or U7524 (N_7524,N_7401,N_7480);
or U7525 (N_7525,N_7496,N_7423);
or U7526 (N_7526,N_7293,N_7482);
nand U7527 (N_7527,N_7263,N_7330);
nor U7528 (N_7528,N_7373,N_7399);
nand U7529 (N_7529,N_7390,N_7261);
and U7530 (N_7530,N_7389,N_7334);
or U7531 (N_7531,N_7410,N_7257);
and U7532 (N_7532,N_7403,N_7283);
xor U7533 (N_7533,N_7355,N_7262);
or U7534 (N_7534,N_7400,N_7464);
nand U7535 (N_7535,N_7430,N_7481);
xor U7536 (N_7536,N_7461,N_7377);
xor U7537 (N_7537,N_7431,N_7375);
xor U7538 (N_7538,N_7404,N_7402);
nor U7539 (N_7539,N_7485,N_7380);
or U7540 (N_7540,N_7296,N_7254);
or U7541 (N_7541,N_7297,N_7492);
nor U7542 (N_7542,N_7284,N_7427);
nor U7543 (N_7543,N_7312,N_7426);
and U7544 (N_7544,N_7331,N_7428);
or U7545 (N_7545,N_7365,N_7384);
and U7546 (N_7546,N_7290,N_7343);
nor U7547 (N_7547,N_7259,N_7383);
nand U7548 (N_7548,N_7446,N_7369);
nand U7549 (N_7549,N_7442,N_7421);
xor U7550 (N_7550,N_7253,N_7445);
nand U7551 (N_7551,N_7372,N_7434);
nor U7552 (N_7552,N_7250,N_7260);
or U7553 (N_7553,N_7288,N_7352);
xnor U7554 (N_7554,N_7474,N_7278);
or U7555 (N_7555,N_7354,N_7285);
and U7556 (N_7556,N_7452,N_7345);
nor U7557 (N_7557,N_7497,N_7438);
or U7558 (N_7558,N_7306,N_7270);
and U7559 (N_7559,N_7484,N_7475);
nor U7560 (N_7560,N_7366,N_7387);
nor U7561 (N_7561,N_7294,N_7405);
or U7562 (N_7562,N_7289,N_7357);
or U7563 (N_7563,N_7465,N_7460);
nor U7564 (N_7564,N_7467,N_7455);
and U7565 (N_7565,N_7376,N_7258);
nor U7566 (N_7566,N_7271,N_7472);
or U7567 (N_7567,N_7418,N_7313);
xor U7568 (N_7568,N_7379,N_7448);
nand U7569 (N_7569,N_7468,N_7479);
nor U7570 (N_7570,N_7358,N_7412);
or U7571 (N_7571,N_7351,N_7364);
nor U7572 (N_7572,N_7397,N_7315);
or U7573 (N_7573,N_7440,N_7483);
or U7574 (N_7574,N_7363,N_7450);
nor U7575 (N_7575,N_7338,N_7382);
xnor U7576 (N_7576,N_7310,N_7308);
nand U7577 (N_7577,N_7251,N_7429);
nor U7578 (N_7578,N_7420,N_7255);
nor U7579 (N_7579,N_7498,N_7356);
xor U7580 (N_7580,N_7307,N_7265);
nor U7581 (N_7581,N_7264,N_7323);
nor U7582 (N_7582,N_7361,N_7444);
and U7583 (N_7583,N_7304,N_7347);
nor U7584 (N_7584,N_7414,N_7407);
or U7585 (N_7585,N_7490,N_7473);
xnor U7586 (N_7586,N_7280,N_7267);
or U7587 (N_7587,N_7322,N_7456);
and U7588 (N_7588,N_7394,N_7300);
or U7589 (N_7589,N_7487,N_7491);
nand U7590 (N_7590,N_7392,N_7339);
nor U7591 (N_7591,N_7370,N_7476);
nand U7592 (N_7592,N_7337,N_7374);
xor U7593 (N_7593,N_7276,N_7329);
xor U7594 (N_7594,N_7333,N_7325);
and U7595 (N_7595,N_7349,N_7305);
nand U7596 (N_7596,N_7459,N_7298);
and U7597 (N_7597,N_7411,N_7477);
and U7598 (N_7598,N_7454,N_7385);
nor U7599 (N_7599,N_7439,N_7432);
and U7600 (N_7600,N_7299,N_7443);
xor U7601 (N_7601,N_7441,N_7314);
and U7602 (N_7602,N_7350,N_7332);
and U7603 (N_7603,N_7344,N_7340);
nand U7604 (N_7604,N_7463,N_7256);
and U7605 (N_7605,N_7406,N_7266);
nor U7606 (N_7606,N_7281,N_7273);
nor U7607 (N_7607,N_7282,N_7395);
nand U7608 (N_7608,N_7316,N_7424);
nand U7609 (N_7609,N_7462,N_7302);
nor U7610 (N_7610,N_7396,N_7447);
nor U7611 (N_7611,N_7393,N_7458);
nand U7612 (N_7612,N_7321,N_7453);
or U7613 (N_7613,N_7378,N_7303);
nor U7614 (N_7614,N_7415,N_7346);
and U7615 (N_7615,N_7277,N_7368);
xor U7616 (N_7616,N_7398,N_7386);
xor U7617 (N_7617,N_7495,N_7416);
or U7618 (N_7618,N_7320,N_7291);
xnor U7619 (N_7619,N_7433,N_7272);
nor U7620 (N_7620,N_7342,N_7292);
and U7621 (N_7621,N_7336,N_7295);
xor U7622 (N_7622,N_7493,N_7489);
nand U7623 (N_7623,N_7449,N_7417);
nand U7624 (N_7624,N_7335,N_7301);
or U7625 (N_7625,N_7303,N_7307);
or U7626 (N_7626,N_7280,N_7393);
nand U7627 (N_7627,N_7293,N_7274);
nand U7628 (N_7628,N_7411,N_7263);
or U7629 (N_7629,N_7466,N_7434);
nor U7630 (N_7630,N_7268,N_7411);
nor U7631 (N_7631,N_7365,N_7343);
or U7632 (N_7632,N_7469,N_7448);
nor U7633 (N_7633,N_7460,N_7464);
and U7634 (N_7634,N_7473,N_7286);
xnor U7635 (N_7635,N_7444,N_7362);
or U7636 (N_7636,N_7350,N_7289);
nor U7637 (N_7637,N_7339,N_7342);
xor U7638 (N_7638,N_7480,N_7354);
xnor U7639 (N_7639,N_7384,N_7287);
xnor U7640 (N_7640,N_7301,N_7267);
xnor U7641 (N_7641,N_7265,N_7346);
or U7642 (N_7642,N_7398,N_7310);
nor U7643 (N_7643,N_7343,N_7262);
nand U7644 (N_7644,N_7419,N_7272);
and U7645 (N_7645,N_7257,N_7255);
and U7646 (N_7646,N_7379,N_7461);
or U7647 (N_7647,N_7466,N_7322);
nand U7648 (N_7648,N_7383,N_7421);
and U7649 (N_7649,N_7460,N_7309);
nand U7650 (N_7650,N_7367,N_7276);
and U7651 (N_7651,N_7269,N_7355);
or U7652 (N_7652,N_7475,N_7393);
or U7653 (N_7653,N_7464,N_7427);
and U7654 (N_7654,N_7365,N_7333);
nand U7655 (N_7655,N_7354,N_7433);
xor U7656 (N_7656,N_7301,N_7399);
or U7657 (N_7657,N_7496,N_7466);
and U7658 (N_7658,N_7363,N_7325);
nor U7659 (N_7659,N_7413,N_7456);
xor U7660 (N_7660,N_7324,N_7313);
or U7661 (N_7661,N_7304,N_7418);
nor U7662 (N_7662,N_7290,N_7333);
nand U7663 (N_7663,N_7307,N_7453);
xnor U7664 (N_7664,N_7314,N_7300);
nor U7665 (N_7665,N_7256,N_7413);
nor U7666 (N_7666,N_7407,N_7413);
or U7667 (N_7667,N_7424,N_7398);
xnor U7668 (N_7668,N_7435,N_7449);
xor U7669 (N_7669,N_7264,N_7448);
xnor U7670 (N_7670,N_7332,N_7475);
xnor U7671 (N_7671,N_7397,N_7311);
or U7672 (N_7672,N_7312,N_7446);
and U7673 (N_7673,N_7430,N_7493);
xnor U7674 (N_7674,N_7467,N_7405);
and U7675 (N_7675,N_7390,N_7347);
or U7676 (N_7676,N_7324,N_7387);
xor U7677 (N_7677,N_7300,N_7349);
and U7678 (N_7678,N_7397,N_7494);
and U7679 (N_7679,N_7312,N_7325);
xnor U7680 (N_7680,N_7454,N_7354);
nand U7681 (N_7681,N_7352,N_7256);
xnor U7682 (N_7682,N_7260,N_7273);
and U7683 (N_7683,N_7334,N_7274);
and U7684 (N_7684,N_7494,N_7476);
nor U7685 (N_7685,N_7458,N_7374);
nand U7686 (N_7686,N_7427,N_7310);
nor U7687 (N_7687,N_7264,N_7301);
xor U7688 (N_7688,N_7304,N_7446);
xor U7689 (N_7689,N_7495,N_7460);
and U7690 (N_7690,N_7250,N_7326);
and U7691 (N_7691,N_7350,N_7269);
nor U7692 (N_7692,N_7470,N_7460);
nor U7693 (N_7693,N_7430,N_7394);
xnor U7694 (N_7694,N_7444,N_7420);
and U7695 (N_7695,N_7437,N_7269);
or U7696 (N_7696,N_7454,N_7468);
and U7697 (N_7697,N_7424,N_7439);
xor U7698 (N_7698,N_7320,N_7279);
nand U7699 (N_7699,N_7471,N_7415);
or U7700 (N_7700,N_7464,N_7407);
nor U7701 (N_7701,N_7415,N_7281);
xnor U7702 (N_7702,N_7462,N_7251);
nor U7703 (N_7703,N_7267,N_7492);
xor U7704 (N_7704,N_7304,N_7476);
nand U7705 (N_7705,N_7347,N_7362);
and U7706 (N_7706,N_7478,N_7304);
or U7707 (N_7707,N_7334,N_7301);
and U7708 (N_7708,N_7483,N_7280);
nand U7709 (N_7709,N_7261,N_7383);
or U7710 (N_7710,N_7498,N_7302);
nand U7711 (N_7711,N_7401,N_7286);
or U7712 (N_7712,N_7452,N_7367);
nand U7713 (N_7713,N_7368,N_7460);
xnor U7714 (N_7714,N_7480,N_7293);
nor U7715 (N_7715,N_7370,N_7313);
nor U7716 (N_7716,N_7284,N_7301);
xor U7717 (N_7717,N_7319,N_7308);
nor U7718 (N_7718,N_7404,N_7488);
nand U7719 (N_7719,N_7359,N_7376);
nand U7720 (N_7720,N_7476,N_7336);
xor U7721 (N_7721,N_7283,N_7401);
or U7722 (N_7722,N_7391,N_7429);
or U7723 (N_7723,N_7485,N_7318);
and U7724 (N_7724,N_7419,N_7367);
nand U7725 (N_7725,N_7358,N_7279);
and U7726 (N_7726,N_7413,N_7324);
nand U7727 (N_7727,N_7307,N_7355);
or U7728 (N_7728,N_7401,N_7327);
nor U7729 (N_7729,N_7474,N_7451);
or U7730 (N_7730,N_7454,N_7485);
nor U7731 (N_7731,N_7460,N_7371);
xor U7732 (N_7732,N_7265,N_7291);
nor U7733 (N_7733,N_7279,N_7338);
or U7734 (N_7734,N_7323,N_7250);
and U7735 (N_7735,N_7437,N_7301);
nand U7736 (N_7736,N_7255,N_7495);
nand U7737 (N_7737,N_7373,N_7405);
xor U7738 (N_7738,N_7331,N_7257);
xor U7739 (N_7739,N_7369,N_7322);
or U7740 (N_7740,N_7287,N_7305);
and U7741 (N_7741,N_7429,N_7375);
nor U7742 (N_7742,N_7462,N_7316);
nand U7743 (N_7743,N_7255,N_7332);
xnor U7744 (N_7744,N_7410,N_7359);
nor U7745 (N_7745,N_7354,N_7327);
nor U7746 (N_7746,N_7308,N_7268);
nand U7747 (N_7747,N_7265,N_7323);
xnor U7748 (N_7748,N_7362,N_7283);
nand U7749 (N_7749,N_7446,N_7344);
and U7750 (N_7750,N_7601,N_7636);
nor U7751 (N_7751,N_7522,N_7500);
nor U7752 (N_7752,N_7611,N_7688);
and U7753 (N_7753,N_7538,N_7729);
and U7754 (N_7754,N_7677,N_7526);
xor U7755 (N_7755,N_7719,N_7617);
and U7756 (N_7756,N_7562,N_7706);
and U7757 (N_7757,N_7702,N_7598);
or U7758 (N_7758,N_7564,N_7687);
xor U7759 (N_7759,N_7614,N_7684);
or U7760 (N_7760,N_7673,N_7672);
xnor U7761 (N_7761,N_7698,N_7704);
and U7762 (N_7762,N_7667,N_7615);
nand U7763 (N_7763,N_7735,N_7543);
xor U7764 (N_7764,N_7693,N_7519);
nand U7765 (N_7765,N_7658,N_7738);
and U7766 (N_7766,N_7559,N_7514);
xnor U7767 (N_7767,N_7690,N_7714);
xor U7768 (N_7768,N_7717,N_7548);
and U7769 (N_7769,N_7647,N_7661);
nand U7770 (N_7770,N_7572,N_7744);
nand U7771 (N_7771,N_7648,N_7604);
or U7772 (N_7772,N_7554,N_7711);
xnor U7773 (N_7773,N_7534,N_7718);
xnor U7774 (N_7774,N_7613,N_7509);
or U7775 (N_7775,N_7629,N_7682);
xnor U7776 (N_7776,N_7565,N_7708);
xor U7777 (N_7777,N_7701,N_7523);
nor U7778 (N_7778,N_7571,N_7511);
or U7779 (N_7779,N_7664,N_7622);
nand U7780 (N_7780,N_7624,N_7605);
nand U7781 (N_7781,N_7640,N_7692);
xnor U7782 (N_7782,N_7505,N_7639);
or U7783 (N_7783,N_7743,N_7533);
and U7784 (N_7784,N_7644,N_7635);
and U7785 (N_7785,N_7650,N_7691);
nor U7786 (N_7786,N_7528,N_7535);
nor U7787 (N_7787,N_7678,N_7620);
xor U7788 (N_7788,N_7632,N_7726);
nand U7789 (N_7789,N_7663,N_7730);
xnor U7790 (N_7790,N_7707,N_7740);
nor U7791 (N_7791,N_7686,N_7521);
xor U7792 (N_7792,N_7699,N_7563);
nor U7793 (N_7793,N_7723,N_7587);
and U7794 (N_7794,N_7558,N_7728);
or U7795 (N_7795,N_7651,N_7621);
and U7796 (N_7796,N_7733,N_7749);
xnor U7797 (N_7797,N_7515,N_7585);
and U7798 (N_7798,N_7731,N_7676);
nor U7799 (N_7799,N_7713,N_7502);
or U7800 (N_7800,N_7685,N_7659);
nand U7801 (N_7801,N_7506,N_7649);
or U7802 (N_7802,N_7697,N_7627);
nand U7803 (N_7803,N_7679,N_7507);
xnor U7804 (N_7804,N_7748,N_7705);
xnor U7805 (N_7805,N_7584,N_7517);
nand U7806 (N_7806,N_7670,N_7724);
and U7807 (N_7807,N_7736,N_7588);
xor U7808 (N_7808,N_7669,N_7510);
and U7809 (N_7809,N_7737,N_7680);
nor U7810 (N_7810,N_7568,N_7583);
or U7811 (N_7811,N_7579,N_7671);
nand U7812 (N_7812,N_7630,N_7596);
nor U7813 (N_7813,N_7549,N_7634);
or U7814 (N_7814,N_7550,N_7745);
xnor U7815 (N_7815,N_7683,N_7626);
xnor U7816 (N_7816,N_7665,N_7712);
xor U7817 (N_7817,N_7551,N_7504);
nor U7818 (N_7818,N_7646,N_7594);
xnor U7819 (N_7819,N_7715,N_7518);
or U7820 (N_7820,N_7542,N_7552);
or U7821 (N_7821,N_7536,N_7734);
nor U7822 (N_7822,N_7592,N_7586);
or U7823 (N_7823,N_7516,N_7593);
nand U7824 (N_7824,N_7603,N_7591);
xnor U7825 (N_7825,N_7747,N_7581);
nand U7826 (N_7826,N_7531,N_7657);
xor U7827 (N_7827,N_7694,N_7606);
and U7828 (N_7828,N_7580,N_7637);
or U7829 (N_7829,N_7545,N_7600);
nor U7830 (N_7830,N_7501,N_7681);
and U7831 (N_7831,N_7546,N_7557);
and U7832 (N_7832,N_7520,N_7556);
and U7833 (N_7833,N_7577,N_7631);
nand U7834 (N_7834,N_7595,N_7638);
or U7835 (N_7835,N_7527,N_7727);
or U7836 (N_7836,N_7643,N_7721);
or U7837 (N_7837,N_7709,N_7503);
nor U7838 (N_7838,N_7739,N_7625);
xor U7839 (N_7839,N_7662,N_7566);
and U7840 (N_7840,N_7652,N_7530);
nand U7841 (N_7841,N_7513,N_7720);
and U7842 (N_7842,N_7696,N_7532);
xor U7843 (N_7843,N_7578,N_7524);
or U7844 (N_7844,N_7674,N_7540);
xnor U7845 (N_7845,N_7508,N_7619);
nor U7846 (N_7846,N_7675,N_7716);
nor U7847 (N_7847,N_7741,N_7618);
and U7848 (N_7848,N_7746,N_7666);
and U7849 (N_7849,N_7576,N_7512);
and U7850 (N_7850,N_7612,N_7725);
or U7851 (N_7851,N_7529,N_7633);
or U7852 (N_7852,N_7573,N_7539);
nor U7853 (N_7853,N_7547,N_7668);
nor U7854 (N_7854,N_7616,N_7608);
xor U7855 (N_7855,N_7544,N_7645);
xor U7856 (N_7856,N_7689,N_7653);
or U7857 (N_7857,N_7574,N_7610);
nor U7858 (N_7858,N_7628,N_7655);
or U7859 (N_7859,N_7700,N_7555);
and U7860 (N_7860,N_7537,N_7569);
and U7861 (N_7861,N_7722,N_7541);
or U7862 (N_7862,N_7732,N_7607);
nor U7863 (N_7863,N_7597,N_7560);
or U7864 (N_7864,N_7602,N_7742);
nand U7865 (N_7865,N_7570,N_7695);
xor U7866 (N_7866,N_7575,N_7654);
or U7867 (N_7867,N_7710,N_7641);
nor U7868 (N_7868,N_7656,N_7590);
and U7869 (N_7869,N_7525,N_7553);
xnor U7870 (N_7870,N_7660,N_7599);
xnor U7871 (N_7871,N_7589,N_7567);
xnor U7872 (N_7872,N_7623,N_7561);
and U7873 (N_7873,N_7582,N_7609);
xor U7874 (N_7874,N_7642,N_7703);
nor U7875 (N_7875,N_7675,N_7598);
xnor U7876 (N_7876,N_7529,N_7712);
and U7877 (N_7877,N_7503,N_7548);
nand U7878 (N_7878,N_7659,N_7669);
xor U7879 (N_7879,N_7572,N_7679);
nor U7880 (N_7880,N_7586,N_7551);
nor U7881 (N_7881,N_7627,N_7688);
nand U7882 (N_7882,N_7660,N_7639);
and U7883 (N_7883,N_7728,N_7594);
xnor U7884 (N_7884,N_7587,N_7667);
nor U7885 (N_7885,N_7677,N_7672);
xor U7886 (N_7886,N_7702,N_7575);
and U7887 (N_7887,N_7630,N_7574);
nand U7888 (N_7888,N_7669,N_7584);
nand U7889 (N_7889,N_7605,N_7507);
and U7890 (N_7890,N_7679,N_7519);
xor U7891 (N_7891,N_7593,N_7652);
and U7892 (N_7892,N_7580,N_7582);
xor U7893 (N_7893,N_7503,N_7532);
xor U7894 (N_7894,N_7583,N_7746);
nand U7895 (N_7895,N_7529,N_7622);
xor U7896 (N_7896,N_7544,N_7699);
xnor U7897 (N_7897,N_7694,N_7638);
nor U7898 (N_7898,N_7718,N_7732);
and U7899 (N_7899,N_7585,N_7680);
or U7900 (N_7900,N_7580,N_7666);
nand U7901 (N_7901,N_7602,N_7651);
xnor U7902 (N_7902,N_7729,N_7508);
nand U7903 (N_7903,N_7627,N_7741);
xnor U7904 (N_7904,N_7634,N_7542);
xor U7905 (N_7905,N_7650,N_7562);
xnor U7906 (N_7906,N_7627,N_7554);
nand U7907 (N_7907,N_7641,N_7725);
xnor U7908 (N_7908,N_7614,N_7601);
or U7909 (N_7909,N_7531,N_7721);
or U7910 (N_7910,N_7663,N_7678);
xnor U7911 (N_7911,N_7749,N_7734);
xnor U7912 (N_7912,N_7741,N_7559);
and U7913 (N_7913,N_7602,N_7513);
nand U7914 (N_7914,N_7593,N_7506);
and U7915 (N_7915,N_7527,N_7506);
xor U7916 (N_7916,N_7588,N_7711);
nor U7917 (N_7917,N_7513,N_7705);
and U7918 (N_7918,N_7533,N_7584);
and U7919 (N_7919,N_7599,N_7511);
xor U7920 (N_7920,N_7529,N_7636);
xnor U7921 (N_7921,N_7501,N_7541);
xnor U7922 (N_7922,N_7542,N_7709);
xor U7923 (N_7923,N_7685,N_7621);
and U7924 (N_7924,N_7524,N_7615);
nor U7925 (N_7925,N_7520,N_7631);
nand U7926 (N_7926,N_7642,N_7687);
nand U7927 (N_7927,N_7651,N_7633);
and U7928 (N_7928,N_7567,N_7696);
xor U7929 (N_7929,N_7722,N_7688);
nor U7930 (N_7930,N_7535,N_7613);
nor U7931 (N_7931,N_7679,N_7634);
nand U7932 (N_7932,N_7661,N_7531);
nor U7933 (N_7933,N_7722,N_7668);
or U7934 (N_7934,N_7508,N_7655);
xor U7935 (N_7935,N_7505,N_7699);
and U7936 (N_7936,N_7564,N_7668);
nor U7937 (N_7937,N_7525,N_7579);
nor U7938 (N_7938,N_7601,N_7723);
xor U7939 (N_7939,N_7717,N_7530);
nand U7940 (N_7940,N_7696,N_7569);
nor U7941 (N_7941,N_7515,N_7691);
nand U7942 (N_7942,N_7610,N_7696);
xor U7943 (N_7943,N_7585,N_7749);
or U7944 (N_7944,N_7674,N_7619);
nand U7945 (N_7945,N_7724,N_7732);
nor U7946 (N_7946,N_7562,N_7564);
or U7947 (N_7947,N_7514,N_7568);
or U7948 (N_7948,N_7588,N_7727);
nand U7949 (N_7949,N_7523,N_7597);
nor U7950 (N_7950,N_7524,N_7661);
and U7951 (N_7951,N_7700,N_7725);
xor U7952 (N_7952,N_7709,N_7567);
xnor U7953 (N_7953,N_7572,N_7522);
nor U7954 (N_7954,N_7552,N_7688);
nand U7955 (N_7955,N_7659,N_7697);
nor U7956 (N_7956,N_7609,N_7666);
xnor U7957 (N_7957,N_7707,N_7579);
nand U7958 (N_7958,N_7721,N_7520);
or U7959 (N_7959,N_7557,N_7664);
and U7960 (N_7960,N_7597,N_7672);
and U7961 (N_7961,N_7631,N_7642);
or U7962 (N_7962,N_7730,N_7538);
xnor U7963 (N_7963,N_7634,N_7741);
xor U7964 (N_7964,N_7657,N_7640);
nor U7965 (N_7965,N_7721,N_7686);
nor U7966 (N_7966,N_7737,N_7719);
nand U7967 (N_7967,N_7524,N_7710);
nor U7968 (N_7968,N_7530,N_7566);
nor U7969 (N_7969,N_7679,N_7671);
nand U7970 (N_7970,N_7690,N_7675);
nand U7971 (N_7971,N_7719,N_7538);
or U7972 (N_7972,N_7615,N_7662);
nor U7973 (N_7973,N_7690,N_7657);
xor U7974 (N_7974,N_7675,N_7655);
and U7975 (N_7975,N_7663,N_7529);
and U7976 (N_7976,N_7525,N_7522);
xnor U7977 (N_7977,N_7694,N_7739);
or U7978 (N_7978,N_7561,N_7730);
or U7979 (N_7979,N_7621,N_7679);
nand U7980 (N_7980,N_7668,N_7725);
and U7981 (N_7981,N_7584,N_7612);
nor U7982 (N_7982,N_7634,N_7704);
xor U7983 (N_7983,N_7628,N_7692);
and U7984 (N_7984,N_7609,N_7550);
or U7985 (N_7985,N_7598,N_7553);
xnor U7986 (N_7986,N_7676,N_7721);
or U7987 (N_7987,N_7634,N_7536);
nor U7988 (N_7988,N_7541,N_7583);
or U7989 (N_7989,N_7709,N_7604);
nand U7990 (N_7990,N_7505,N_7701);
or U7991 (N_7991,N_7733,N_7746);
nand U7992 (N_7992,N_7742,N_7711);
xor U7993 (N_7993,N_7628,N_7519);
and U7994 (N_7994,N_7671,N_7591);
nand U7995 (N_7995,N_7513,N_7713);
nor U7996 (N_7996,N_7711,N_7545);
xnor U7997 (N_7997,N_7679,N_7655);
or U7998 (N_7998,N_7691,N_7657);
and U7999 (N_7999,N_7621,N_7501);
or U8000 (N_8000,N_7814,N_7992);
or U8001 (N_8001,N_7918,N_7855);
nand U8002 (N_8002,N_7877,N_7803);
or U8003 (N_8003,N_7982,N_7836);
nand U8004 (N_8004,N_7808,N_7797);
nand U8005 (N_8005,N_7965,N_7755);
nor U8006 (N_8006,N_7779,N_7997);
and U8007 (N_8007,N_7975,N_7981);
xor U8008 (N_8008,N_7765,N_7969);
nor U8009 (N_8009,N_7781,N_7957);
or U8010 (N_8010,N_7782,N_7769);
nand U8011 (N_8011,N_7931,N_7860);
or U8012 (N_8012,N_7942,N_7810);
and U8013 (N_8013,N_7928,N_7983);
or U8014 (N_8014,N_7921,N_7955);
and U8015 (N_8015,N_7880,N_7909);
and U8016 (N_8016,N_7937,N_7932);
or U8017 (N_8017,N_7904,N_7787);
and U8018 (N_8018,N_7775,N_7919);
nand U8019 (N_8019,N_7973,N_7999);
nor U8020 (N_8020,N_7913,N_7883);
xnor U8021 (N_8021,N_7758,N_7795);
and U8022 (N_8022,N_7944,N_7876);
or U8023 (N_8023,N_7867,N_7771);
xnor U8024 (N_8024,N_7900,N_7933);
nor U8025 (N_8025,N_7946,N_7766);
and U8026 (N_8026,N_7784,N_7839);
or U8027 (N_8027,N_7798,N_7847);
nor U8028 (N_8028,N_7953,N_7911);
xnor U8029 (N_8029,N_7948,N_7993);
or U8030 (N_8030,N_7772,N_7927);
or U8031 (N_8031,N_7789,N_7812);
and U8032 (N_8032,N_7967,N_7988);
xor U8033 (N_8033,N_7793,N_7972);
nor U8034 (N_8034,N_7892,N_7936);
nor U8035 (N_8035,N_7869,N_7773);
nor U8036 (N_8036,N_7974,N_7903);
and U8037 (N_8037,N_7970,N_7785);
nand U8038 (N_8038,N_7873,N_7846);
and U8039 (N_8039,N_7825,N_7833);
or U8040 (N_8040,N_7934,N_7998);
nor U8041 (N_8041,N_7802,N_7882);
and U8042 (N_8042,N_7905,N_7887);
nor U8043 (N_8043,N_7895,N_7837);
or U8044 (N_8044,N_7767,N_7954);
nand U8045 (N_8045,N_7757,N_7906);
xor U8046 (N_8046,N_7929,N_7759);
xor U8047 (N_8047,N_7991,N_7939);
or U8048 (N_8048,N_7786,N_7870);
xnor U8049 (N_8049,N_7813,N_7897);
and U8050 (N_8050,N_7807,N_7894);
xnor U8051 (N_8051,N_7801,N_7985);
nor U8052 (N_8052,N_7893,N_7899);
nor U8053 (N_8053,N_7861,N_7852);
xor U8054 (N_8054,N_7823,N_7886);
xor U8055 (N_8055,N_7960,N_7878);
xor U8056 (N_8056,N_7820,N_7842);
nor U8057 (N_8057,N_7764,N_7831);
and U8058 (N_8058,N_7815,N_7940);
nor U8059 (N_8059,N_7912,N_7995);
xnor U8060 (N_8060,N_7834,N_7824);
xor U8061 (N_8061,N_7752,N_7865);
xor U8062 (N_8062,N_7851,N_7858);
or U8063 (N_8063,N_7818,N_7874);
nand U8064 (N_8064,N_7863,N_7956);
xnor U8065 (N_8065,N_7753,N_7788);
and U8066 (N_8066,N_7796,N_7838);
and U8067 (N_8067,N_7854,N_7890);
or U8068 (N_8068,N_7862,N_7952);
nor U8069 (N_8069,N_7829,N_7941);
or U8070 (N_8070,N_7857,N_7989);
nor U8071 (N_8071,N_7935,N_7968);
and U8072 (N_8072,N_7938,N_7920);
and U8073 (N_8073,N_7971,N_7791);
and U8074 (N_8074,N_7907,N_7875);
nand U8075 (N_8075,N_7868,N_7783);
or U8076 (N_8076,N_7827,N_7884);
nand U8077 (N_8077,N_7891,N_7819);
and U8078 (N_8078,N_7996,N_7950);
nand U8079 (N_8079,N_7864,N_7966);
nor U8080 (N_8080,N_7790,N_7843);
or U8081 (N_8081,N_7915,N_7849);
or U8082 (N_8082,N_7770,N_7848);
or U8083 (N_8083,N_7964,N_7751);
nor U8084 (N_8084,N_7879,N_7816);
and U8085 (N_8085,N_7821,N_7961);
nor U8086 (N_8086,N_7871,N_7925);
xnor U8087 (N_8087,N_7830,N_7845);
xor U8088 (N_8088,N_7959,N_7951);
and U8089 (N_8089,N_7976,N_7898);
nand U8090 (N_8090,N_7756,N_7805);
or U8091 (N_8091,N_7853,N_7979);
xor U8092 (N_8092,N_7910,N_7914);
nand U8093 (N_8093,N_7943,N_7872);
and U8094 (N_8094,N_7844,N_7866);
or U8095 (N_8095,N_7908,N_7841);
nor U8096 (N_8096,N_7822,N_7922);
nor U8097 (N_8097,N_7828,N_7809);
xnor U8098 (N_8098,N_7840,N_7859);
nand U8099 (N_8099,N_7792,N_7977);
and U8100 (N_8100,N_7888,N_7949);
and U8101 (N_8101,N_7761,N_7924);
xor U8102 (N_8102,N_7901,N_7962);
and U8103 (N_8103,N_7835,N_7923);
nand U8104 (N_8104,N_7776,N_7806);
nor U8105 (N_8105,N_7763,N_7804);
xnor U8106 (N_8106,N_7889,N_7754);
and U8107 (N_8107,N_7832,N_7826);
nand U8108 (N_8108,N_7980,N_7850);
and U8109 (N_8109,N_7986,N_7800);
xor U8110 (N_8110,N_7947,N_7987);
xor U8111 (N_8111,N_7926,N_7990);
xor U8112 (N_8112,N_7885,N_7774);
or U8113 (N_8113,N_7902,N_7958);
nor U8114 (N_8114,N_7777,N_7963);
nand U8115 (N_8115,N_7856,N_7945);
nand U8116 (N_8116,N_7799,N_7762);
xor U8117 (N_8117,N_7817,N_7896);
nand U8118 (N_8118,N_7930,N_7978);
and U8119 (N_8119,N_7811,N_7794);
and U8120 (N_8120,N_7780,N_7768);
xnor U8121 (N_8121,N_7760,N_7984);
nand U8122 (N_8122,N_7916,N_7917);
nor U8123 (N_8123,N_7778,N_7994);
nor U8124 (N_8124,N_7881,N_7750);
xnor U8125 (N_8125,N_7943,N_7876);
nand U8126 (N_8126,N_7956,N_7949);
and U8127 (N_8127,N_7993,N_7882);
xor U8128 (N_8128,N_7949,N_7937);
or U8129 (N_8129,N_7991,N_7850);
or U8130 (N_8130,N_7852,N_7873);
and U8131 (N_8131,N_7775,N_7756);
xnor U8132 (N_8132,N_7891,N_7765);
xnor U8133 (N_8133,N_7906,N_7873);
nand U8134 (N_8134,N_7917,N_7993);
nand U8135 (N_8135,N_7795,N_7790);
and U8136 (N_8136,N_7858,N_7968);
or U8137 (N_8137,N_7758,N_7866);
nand U8138 (N_8138,N_7935,N_7949);
xor U8139 (N_8139,N_7989,N_7983);
xnor U8140 (N_8140,N_7813,N_7995);
nor U8141 (N_8141,N_7785,N_7755);
or U8142 (N_8142,N_7895,N_7973);
or U8143 (N_8143,N_7855,N_7972);
or U8144 (N_8144,N_7901,N_7998);
nor U8145 (N_8145,N_7913,N_7936);
nor U8146 (N_8146,N_7787,N_7953);
and U8147 (N_8147,N_7917,N_7786);
or U8148 (N_8148,N_7867,N_7994);
xor U8149 (N_8149,N_7988,N_7927);
or U8150 (N_8150,N_7761,N_7938);
nand U8151 (N_8151,N_7768,N_7937);
or U8152 (N_8152,N_7793,N_7943);
xor U8153 (N_8153,N_7762,N_7866);
xnor U8154 (N_8154,N_7839,N_7918);
or U8155 (N_8155,N_7919,N_7819);
nand U8156 (N_8156,N_7923,N_7876);
xnor U8157 (N_8157,N_7853,N_7895);
nor U8158 (N_8158,N_7944,N_7925);
xnor U8159 (N_8159,N_7839,N_7763);
nand U8160 (N_8160,N_7982,N_7940);
nand U8161 (N_8161,N_7754,N_7907);
nand U8162 (N_8162,N_7920,N_7933);
xor U8163 (N_8163,N_7896,N_7824);
or U8164 (N_8164,N_7834,N_7836);
nand U8165 (N_8165,N_7905,N_7835);
and U8166 (N_8166,N_7856,N_7988);
or U8167 (N_8167,N_7841,N_7793);
nor U8168 (N_8168,N_7756,N_7764);
or U8169 (N_8169,N_7792,N_7827);
nor U8170 (N_8170,N_7800,N_7752);
nand U8171 (N_8171,N_7751,N_7836);
or U8172 (N_8172,N_7814,N_7940);
or U8173 (N_8173,N_7939,N_7990);
or U8174 (N_8174,N_7793,N_7873);
and U8175 (N_8175,N_7952,N_7852);
or U8176 (N_8176,N_7911,N_7791);
and U8177 (N_8177,N_7853,N_7850);
nand U8178 (N_8178,N_7837,N_7828);
xnor U8179 (N_8179,N_7828,N_7967);
or U8180 (N_8180,N_7953,N_7847);
or U8181 (N_8181,N_7884,N_7833);
nand U8182 (N_8182,N_7869,N_7845);
and U8183 (N_8183,N_7843,N_7989);
xnor U8184 (N_8184,N_7869,N_7927);
and U8185 (N_8185,N_7953,N_7755);
and U8186 (N_8186,N_7779,N_7836);
nand U8187 (N_8187,N_7891,N_7822);
and U8188 (N_8188,N_7841,N_7871);
nor U8189 (N_8189,N_7942,N_7983);
xor U8190 (N_8190,N_7795,N_7811);
xor U8191 (N_8191,N_7797,N_7864);
xnor U8192 (N_8192,N_7934,N_7930);
nor U8193 (N_8193,N_7932,N_7833);
xnor U8194 (N_8194,N_7822,N_7879);
xor U8195 (N_8195,N_7874,N_7838);
nand U8196 (N_8196,N_7788,N_7825);
nor U8197 (N_8197,N_7773,N_7944);
or U8198 (N_8198,N_7844,N_7948);
and U8199 (N_8199,N_7777,N_7908);
nand U8200 (N_8200,N_7870,N_7965);
nand U8201 (N_8201,N_7836,N_7977);
nor U8202 (N_8202,N_7958,N_7819);
nand U8203 (N_8203,N_7754,N_7938);
xor U8204 (N_8204,N_7982,N_7758);
or U8205 (N_8205,N_7899,N_7900);
nand U8206 (N_8206,N_7960,N_7785);
nor U8207 (N_8207,N_7928,N_7948);
nand U8208 (N_8208,N_7959,N_7831);
and U8209 (N_8209,N_7937,N_7991);
nand U8210 (N_8210,N_7764,N_7869);
and U8211 (N_8211,N_7765,N_7904);
nor U8212 (N_8212,N_7876,N_7906);
or U8213 (N_8213,N_7863,N_7777);
nor U8214 (N_8214,N_7780,N_7879);
nand U8215 (N_8215,N_7868,N_7751);
nand U8216 (N_8216,N_7765,N_7987);
and U8217 (N_8217,N_7762,N_7940);
or U8218 (N_8218,N_7857,N_7999);
and U8219 (N_8219,N_7836,N_7839);
xor U8220 (N_8220,N_7926,N_7946);
and U8221 (N_8221,N_7842,N_7956);
or U8222 (N_8222,N_7827,N_7946);
nor U8223 (N_8223,N_7804,N_7815);
and U8224 (N_8224,N_7911,N_7934);
nor U8225 (N_8225,N_7922,N_7930);
xnor U8226 (N_8226,N_7878,N_7935);
xnor U8227 (N_8227,N_7813,N_7934);
xnor U8228 (N_8228,N_7996,N_7876);
nand U8229 (N_8229,N_7916,N_7819);
nand U8230 (N_8230,N_7934,N_7952);
nand U8231 (N_8231,N_7922,N_7844);
and U8232 (N_8232,N_7878,N_7765);
or U8233 (N_8233,N_7853,N_7847);
nand U8234 (N_8234,N_7972,N_7820);
or U8235 (N_8235,N_7812,N_7800);
and U8236 (N_8236,N_7941,N_7958);
and U8237 (N_8237,N_7950,N_7879);
nor U8238 (N_8238,N_7980,N_7940);
nor U8239 (N_8239,N_7979,N_7968);
nor U8240 (N_8240,N_7936,N_7966);
nand U8241 (N_8241,N_7875,N_7766);
nand U8242 (N_8242,N_7860,N_7784);
or U8243 (N_8243,N_7901,N_7910);
nand U8244 (N_8244,N_7922,N_7842);
and U8245 (N_8245,N_7821,N_7868);
xor U8246 (N_8246,N_7774,N_7900);
nand U8247 (N_8247,N_7935,N_7789);
xor U8248 (N_8248,N_7949,N_7963);
or U8249 (N_8249,N_7777,N_7801);
nor U8250 (N_8250,N_8178,N_8222);
nand U8251 (N_8251,N_8232,N_8139);
and U8252 (N_8252,N_8208,N_8237);
nand U8253 (N_8253,N_8064,N_8205);
nor U8254 (N_8254,N_8090,N_8000);
xnor U8255 (N_8255,N_8249,N_8078);
nand U8256 (N_8256,N_8083,N_8246);
xor U8257 (N_8257,N_8218,N_8063);
nand U8258 (N_8258,N_8120,N_8239);
nand U8259 (N_8259,N_8019,N_8115);
or U8260 (N_8260,N_8045,N_8032);
xor U8261 (N_8261,N_8065,N_8085);
and U8262 (N_8262,N_8073,N_8013);
or U8263 (N_8263,N_8099,N_8056);
nor U8264 (N_8264,N_8068,N_8102);
nand U8265 (N_8265,N_8195,N_8125);
and U8266 (N_8266,N_8191,N_8159);
or U8267 (N_8267,N_8118,N_8135);
nor U8268 (N_8268,N_8214,N_8132);
and U8269 (N_8269,N_8180,N_8247);
nor U8270 (N_8270,N_8052,N_8058);
nand U8271 (N_8271,N_8174,N_8213);
nor U8272 (N_8272,N_8110,N_8181);
or U8273 (N_8273,N_8012,N_8016);
and U8274 (N_8274,N_8037,N_8154);
and U8275 (N_8275,N_8034,N_8241);
nand U8276 (N_8276,N_8179,N_8164);
nand U8277 (N_8277,N_8224,N_8106);
or U8278 (N_8278,N_8201,N_8143);
xor U8279 (N_8279,N_8057,N_8113);
xor U8280 (N_8280,N_8217,N_8119);
or U8281 (N_8281,N_8131,N_8226);
or U8282 (N_8282,N_8039,N_8146);
nor U8283 (N_8283,N_8108,N_8163);
or U8284 (N_8284,N_8173,N_8008);
xor U8285 (N_8285,N_8194,N_8089);
nor U8286 (N_8286,N_8026,N_8053);
xnor U8287 (N_8287,N_8169,N_8192);
nand U8288 (N_8288,N_8041,N_8002);
or U8289 (N_8289,N_8055,N_8081);
and U8290 (N_8290,N_8087,N_8242);
and U8291 (N_8291,N_8104,N_8022);
and U8292 (N_8292,N_8031,N_8123);
xnor U8293 (N_8293,N_8162,N_8015);
nand U8294 (N_8294,N_8138,N_8040);
xnor U8295 (N_8295,N_8095,N_8185);
and U8296 (N_8296,N_8235,N_8018);
or U8297 (N_8297,N_8049,N_8170);
and U8298 (N_8298,N_8175,N_8137);
and U8299 (N_8299,N_8003,N_8133);
xnor U8300 (N_8300,N_8079,N_8004);
xor U8301 (N_8301,N_8197,N_8209);
xnor U8302 (N_8302,N_8212,N_8062);
and U8303 (N_8303,N_8007,N_8144);
nor U8304 (N_8304,N_8027,N_8070);
or U8305 (N_8305,N_8029,N_8060);
nor U8306 (N_8306,N_8158,N_8109);
or U8307 (N_8307,N_8005,N_8066);
and U8308 (N_8308,N_8204,N_8076);
or U8309 (N_8309,N_8184,N_8020);
nand U8310 (N_8310,N_8152,N_8199);
and U8311 (N_8311,N_8088,N_8200);
nor U8312 (N_8312,N_8077,N_8025);
and U8313 (N_8313,N_8189,N_8091);
or U8314 (N_8314,N_8219,N_8134);
nor U8315 (N_8315,N_8117,N_8047);
xnor U8316 (N_8316,N_8238,N_8156);
xor U8317 (N_8317,N_8236,N_8030);
nand U8318 (N_8318,N_8054,N_8202);
and U8319 (N_8319,N_8017,N_8033);
xor U8320 (N_8320,N_8101,N_8096);
xor U8321 (N_8321,N_8050,N_8142);
nand U8322 (N_8322,N_8067,N_8231);
or U8323 (N_8323,N_8245,N_8248);
or U8324 (N_8324,N_8177,N_8021);
or U8325 (N_8325,N_8098,N_8121);
nor U8326 (N_8326,N_8084,N_8234);
or U8327 (N_8327,N_8105,N_8075);
xnor U8328 (N_8328,N_8230,N_8190);
or U8329 (N_8329,N_8176,N_8072);
or U8330 (N_8330,N_8046,N_8042);
or U8331 (N_8331,N_8048,N_8207);
nor U8332 (N_8332,N_8182,N_8086);
or U8333 (N_8333,N_8233,N_8127);
and U8334 (N_8334,N_8206,N_8043);
nand U8335 (N_8335,N_8129,N_8069);
or U8336 (N_8336,N_8116,N_8186);
or U8337 (N_8337,N_8168,N_8059);
or U8338 (N_8338,N_8010,N_8225);
xor U8339 (N_8339,N_8097,N_8211);
xor U8340 (N_8340,N_8128,N_8051);
or U8341 (N_8341,N_8220,N_8240);
xor U8342 (N_8342,N_8183,N_8215);
or U8343 (N_8343,N_8130,N_8023);
xor U8344 (N_8344,N_8122,N_8161);
and U8345 (N_8345,N_8153,N_8140);
nand U8346 (N_8346,N_8011,N_8093);
nor U8347 (N_8347,N_8193,N_8223);
nor U8348 (N_8348,N_8229,N_8111);
nor U8349 (N_8349,N_8114,N_8074);
and U8350 (N_8350,N_8035,N_8126);
or U8351 (N_8351,N_8082,N_8221);
or U8352 (N_8352,N_8001,N_8172);
nor U8353 (N_8353,N_8107,N_8149);
nor U8354 (N_8354,N_8187,N_8014);
nor U8355 (N_8355,N_8036,N_8210);
or U8356 (N_8356,N_8228,N_8203);
xor U8357 (N_8357,N_8094,N_8165);
nor U8358 (N_8358,N_8150,N_8044);
nor U8359 (N_8359,N_8028,N_8244);
and U8360 (N_8360,N_8071,N_8147);
nand U8361 (N_8361,N_8167,N_8006);
and U8362 (N_8362,N_8141,N_8009);
nand U8363 (N_8363,N_8151,N_8160);
or U8364 (N_8364,N_8092,N_8024);
nor U8365 (N_8365,N_8196,N_8155);
nand U8366 (N_8366,N_8198,N_8171);
or U8367 (N_8367,N_8061,N_8124);
and U8368 (N_8368,N_8112,N_8243);
nor U8369 (N_8369,N_8080,N_8100);
nor U8370 (N_8370,N_8136,N_8227);
and U8371 (N_8371,N_8188,N_8166);
nand U8372 (N_8372,N_8145,N_8157);
nor U8373 (N_8373,N_8148,N_8103);
xnor U8374 (N_8374,N_8038,N_8216);
or U8375 (N_8375,N_8057,N_8031);
and U8376 (N_8376,N_8167,N_8176);
xor U8377 (N_8377,N_8093,N_8236);
or U8378 (N_8378,N_8003,N_8033);
nand U8379 (N_8379,N_8167,N_8152);
xor U8380 (N_8380,N_8144,N_8020);
nand U8381 (N_8381,N_8062,N_8241);
or U8382 (N_8382,N_8033,N_8108);
and U8383 (N_8383,N_8149,N_8135);
xnor U8384 (N_8384,N_8144,N_8023);
nor U8385 (N_8385,N_8010,N_8040);
nand U8386 (N_8386,N_8090,N_8225);
or U8387 (N_8387,N_8056,N_8114);
or U8388 (N_8388,N_8096,N_8216);
or U8389 (N_8389,N_8074,N_8142);
xnor U8390 (N_8390,N_8040,N_8102);
xor U8391 (N_8391,N_8188,N_8143);
nor U8392 (N_8392,N_8176,N_8004);
xor U8393 (N_8393,N_8078,N_8028);
or U8394 (N_8394,N_8046,N_8198);
nor U8395 (N_8395,N_8070,N_8211);
nor U8396 (N_8396,N_8014,N_8202);
or U8397 (N_8397,N_8227,N_8055);
and U8398 (N_8398,N_8124,N_8179);
nor U8399 (N_8399,N_8219,N_8100);
nor U8400 (N_8400,N_8248,N_8236);
nand U8401 (N_8401,N_8057,N_8184);
or U8402 (N_8402,N_8191,N_8145);
nand U8403 (N_8403,N_8003,N_8234);
xnor U8404 (N_8404,N_8023,N_8024);
nor U8405 (N_8405,N_8158,N_8015);
nor U8406 (N_8406,N_8217,N_8160);
or U8407 (N_8407,N_8157,N_8130);
and U8408 (N_8408,N_8041,N_8071);
nor U8409 (N_8409,N_8079,N_8016);
or U8410 (N_8410,N_8003,N_8120);
and U8411 (N_8411,N_8147,N_8222);
nor U8412 (N_8412,N_8018,N_8099);
nand U8413 (N_8413,N_8235,N_8104);
or U8414 (N_8414,N_8149,N_8060);
xor U8415 (N_8415,N_8208,N_8082);
nand U8416 (N_8416,N_8060,N_8011);
nand U8417 (N_8417,N_8223,N_8030);
nand U8418 (N_8418,N_8230,N_8118);
xor U8419 (N_8419,N_8222,N_8056);
nand U8420 (N_8420,N_8101,N_8013);
and U8421 (N_8421,N_8192,N_8081);
or U8422 (N_8422,N_8131,N_8080);
nand U8423 (N_8423,N_8158,N_8081);
xor U8424 (N_8424,N_8187,N_8139);
and U8425 (N_8425,N_8121,N_8223);
nand U8426 (N_8426,N_8169,N_8143);
nor U8427 (N_8427,N_8170,N_8059);
nor U8428 (N_8428,N_8033,N_8050);
nor U8429 (N_8429,N_8067,N_8189);
or U8430 (N_8430,N_8209,N_8065);
nand U8431 (N_8431,N_8149,N_8226);
nor U8432 (N_8432,N_8213,N_8010);
xnor U8433 (N_8433,N_8174,N_8061);
xnor U8434 (N_8434,N_8129,N_8009);
nand U8435 (N_8435,N_8135,N_8236);
nor U8436 (N_8436,N_8107,N_8105);
and U8437 (N_8437,N_8158,N_8204);
nor U8438 (N_8438,N_8165,N_8191);
xor U8439 (N_8439,N_8249,N_8219);
nor U8440 (N_8440,N_8080,N_8128);
nand U8441 (N_8441,N_8024,N_8073);
xor U8442 (N_8442,N_8017,N_8179);
nand U8443 (N_8443,N_8182,N_8124);
nand U8444 (N_8444,N_8244,N_8083);
xor U8445 (N_8445,N_8002,N_8166);
nor U8446 (N_8446,N_8141,N_8149);
or U8447 (N_8447,N_8139,N_8241);
or U8448 (N_8448,N_8120,N_8152);
xor U8449 (N_8449,N_8102,N_8088);
or U8450 (N_8450,N_8118,N_8180);
or U8451 (N_8451,N_8089,N_8058);
nand U8452 (N_8452,N_8022,N_8037);
xor U8453 (N_8453,N_8114,N_8080);
nand U8454 (N_8454,N_8188,N_8038);
or U8455 (N_8455,N_8193,N_8115);
and U8456 (N_8456,N_8223,N_8140);
or U8457 (N_8457,N_8172,N_8107);
nand U8458 (N_8458,N_8018,N_8200);
or U8459 (N_8459,N_8235,N_8192);
nand U8460 (N_8460,N_8248,N_8228);
and U8461 (N_8461,N_8006,N_8111);
nor U8462 (N_8462,N_8006,N_8199);
or U8463 (N_8463,N_8113,N_8085);
nand U8464 (N_8464,N_8210,N_8209);
nor U8465 (N_8465,N_8039,N_8055);
nor U8466 (N_8466,N_8110,N_8225);
and U8467 (N_8467,N_8148,N_8075);
xor U8468 (N_8468,N_8125,N_8110);
or U8469 (N_8469,N_8027,N_8211);
and U8470 (N_8470,N_8218,N_8085);
nor U8471 (N_8471,N_8125,N_8141);
nand U8472 (N_8472,N_8169,N_8043);
nand U8473 (N_8473,N_8162,N_8178);
and U8474 (N_8474,N_8091,N_8007);
nand U8475 (N_8475,N_8235,N_8075);
and U8476 (N_8476,N_8120,N_8070);
xor U8477 (N_8477,N_8203,N_8191);
nor U8478 (N_8478,N_8039,N_8219);
nand U8479 (N_8479,N_8125,N_8153);
xor U8480 (N_8480,N_8238,N_8074);
and U8481 (N_8481,N_8077,N_8195);
and U8482 (N_8482,N_8049,N_8089);
nand U8483 (N_8483,N_8153,N_8036);
nand U8484 (N_8484,N_8083,N_8131);
nor U8485 (N_8485,N_8028,N_8232);
xnor U8486 (N_8486,N_8086,N_8089);
nand U8487 (N_8487,N_8206,N_8062);
or U8488 (N_8488,N_8035,N_8187);
xor U8489 (N_8489,N_8160,N_8044);
nor U8490 (N_8490,N_8213,N_8102);
xor U8491 (N_8491,N_8066,N_8055);
nand U8492 (N_8492,N_8065,N_8055);
xnor U8493 (N_8493,N_8004,N_8055);
nand U8494 (N_8494,N_8174,N_8161);
and U8495 (N_8495,N_8235,N_8236);
nor U8496 (N_8496,N_8114,N_8174);
or U8497 (N_8497,N_8095,N_8073);
nand U8498 (N_8498,N_8057,N_8038);
nand U8499 (N_8499,N_8128,N_8094);
or U8500 (N_8500,N_8455,N_8345);
nand U8501 (N_8501,N_8483,N_8318);
nand U8502 (N_8502,N_8374,N_8261);
nor U8503 (N_8503,N_8356,N_8252);
and U8504 (N_8504,N_8383,N_8382);
xnor U8505 (N_8505,N_8404,N_8451);
and U8506 (N_8506,N_8341,N_8293);
nand U8507 (N_8507,N_8322,N_8365);
nor U8508 (N_8508,N_8277,N_8364);
nand U8509 (N_8509,N_8308,N_8371);
nand U8510 (N_8510,N_8271,N_8388);
and U8511 (N_8511,N_8448,N_8367);
and U8512 (N_8512,N_8454,N_8408);
nand U8513 (N_8513,N_8427,N_8332);
xor U8514 (N_8514,N_8311,N_8310);
xor U8515 (N_8515,N_8424,N_8285);
nor U8516 (N_8516,N_8411,N_8436);
nor U8517 (N_8517,N_8279,N_8290);
nand U8518 (N_8518,N_8428,N_8385);
xnor U8519 (N_8519,N_8409,N_8460);
nand U8520 (N_8520,N_8278,N_8340);
xnor U8521 (N_8521,N_8349,N_8346);
and U8522 (N_8522,N_8302,N_8420);
and U8523 (N_8523,N_8276,N_8353);
or U8524 (N_8524,N_8257,N_8274);
nand U8525 (N_8525,N_8369,N_8312);
and U8526 (N_8526,N_8434,N_8399);
or U8527 (N_8527,N_8272,N_8260);
nor U8528 (N_8528,N_8498,N_8425);
xor U8529 (N_8529,N_8407,N_8415);
nor U8530 (N_8530,N_8284,N_8363);
and U8531 (N_8531,N_8360,N_8323);
or U8532 (N_8532,N_8444,N_8389);
or U8533 (N_8533,N_8354,N_8289);
and U8534 (N_8534,N_8485,N_8372);
nor U8535 (N_8535,N_8307,N_8362);
or U8536 (N_8536,N_8273,N_8343);
nor U8537 (N_8537,N_8496,N_8432);
nor U8538 (N_8538,N_8294,N_8442);
nand U8539 (N_8539,N_8440,N_8291);
and U8540 (N_8540,N_8426,N_8412);
or U8541 (N_8541,N_8472,N_8446);
nor U8542 (N_8542,N_8377,N_8480);
nor U8543 (N_8543,N_8392,N_8326);
nand U8544 (N_8544,N_8300,N_8282);
xor U8545 (N_8545,N_8469,N_8431);
or U8546 (N_8546,N_8250,N_8286);
or U8547 (N_8547,N_8430,N_8380);
and U8548 (N_8548,N_8254,N_8378);
and U8549 (N_8549,N_8330,N_8334);
xor U8550 (N_8550,N_8418,N_8479);
and U8551 (N_8551,N_8296,N_8410);
and U8552 (N_8552,N_8394,N_8456);
and U8553 (N_8553,N_8297,N_8347);
nor U8554 (N_8554,N_8459,N_8406);
or U8555 (N_8555,N_8268,N_8488);
and U8556 (N_8556,N_8466,N_8379);
nand U8557 (N_8557,N_8361,N_8251);
and U8558 (N_8558,N_8309,N_8338);
or U8559 (N_8559,N_8405,N_8495);
nand U8560 (N_8560,N_8355,N_8450);
nand U8561 (N_8561,N_8384,N_8475);
xor U8562 (N_8562,N_8484,N_8489);
xor U8563 (N_8563,N_8333,N_8373);
xor U8564 (N_8564,N_8449,N_8281);
xor U8565 (N_8565,N_8470,N_8481);
xnor U8566 (N_8566,N_8299,N_8462);
nand U8567 (N_8567,N_8437,N_8453);
nand U8568 (N_8568,N_8403,N_8357);
nand U8569 (N_8569,N_8468,N_8387);
or U8570 (N_8570,N_8329,N_8391);
nand U8571 (N_8571,N_8263,N_8352);
nand U8572 (N_8572,N_8256,N_8315);
and U8573 (N_8573,N_8473,N_8381);
nor U8574 (N_8574,N_8267,N_8313);
nand U8575 (N_8575,N_8401,N_8370);
or U8576 (N_8576,N_8283,N_8325);
or U8577 (N_8577,N_8266,N_8348);
or U8578 (N_8578,N_8328,N_8350);
nand U8579 (N_8579,N_8270,N_8482);
and U8580 (N_8580,N_8474,N_8331);
xnor U8581 (N_8581,N_8393,N_8429);
xnor U8582 (N_8582,N_8464,N_8397);
nor U8583 (N_8583,N_8417,N_8258);
and U8584 (N_8584,N_8478,N_8452);
nand U8585 (N_8585,N_8265,N_8320);
nand U8586 (N_8586,N_8317,N_8376);
and U8587 (N_8587,N_8324,N_8262);
nor U8588 (N_8588,N_8390,N_8447);
xor U8589 (N_8589,N_8337,N_8327);
and U8590 (N_8590,N_8269,N_8366);
nor U8591 (N_8591,N_8416,N_8301);
xnor U8592 (N_8592,N_8264,N_8344);
xor U8593 (N_8593,N_8467,N_8493);
xnor U8594 (N_8594,N_8303,N_8458);
nor U8595 (N_8595,N_8435,N_8491);
and U8596 (N_8596,N_8477,N_8295);
nor U8597 (N_8597,N_8463,N_8499);
or U8598 (N_8598,N_8487,N_8413);
nor U8599 (N_8599,N_8321,N_8457);
or U8600 (N_8600,N_8398,N_8396);
nand U8601 (N_8601,N_8445,N_8359);
or U8602 (N_8602,N_8386,N_8465);
xor U8603 (N_8603,N_8492,N_8486);
nand U8604 (N_8604,N_8422,N_8305);
and U8605 (N_8605,N_8368,N_8443);
nor U8606 (N_8606,N_8438,N_8306);
or U8607 (N_8607,N_8402,N_8395);
nor U8608 (N_8608,N_8423,N_8414);
nor U8609 (N_8609,N_8441,N_8497);
xor U8610 (N_8610,N_8433,N_8490);
xor U8611 (N_8611,N_8253,N_8471);
xnor U8612 (N_8612,N_8314,N_8419);
and U8613 (N_8613,N_8304,N_8298);
and U8614 (N_8614,N_8292,N_8358);
nor U8615 (N_8615,N_8494,N_8319);
xnor U8616 (N_8616,N_8259,N_8280);
xnor U8617 (N_8617,N_8461,N_8351);
and U8618 (N_8618,N_8476,N_8342);
xor U8619 (N_8619,N_8288,N_8439);
and U8620 (N_8620,N_8375,N_8339);
or U8621 (N_8621,N_8400,N_8255);
nor U8622 (N_8622,N_8336,N_8335);
or U8623 (N_8623,N_8287,N_8316);
xnor U8624 (N_8624,N_8275,N_8421);
nor U8625 (N_8625,N_8442,N_8349);
and U8626 (N_8626,N_8304,N_8441);
nand U8627 (N_8627,N_8390,N_8291);
or U8628 (N_8628,N_8440,N_8340);
or U8629 (N_8629,N_8492,N_8471);
xnor U8630 (N_8630,N_8312,N_8302);
nor U8631 (N_8631,N_8469,N_8335);
nor U8632 (N_8632,N_8433,N_8323);
nor U8633 (N_8633,N_8498,N_8408);
nor U8634 (N_8634,N_8300,N_8421);
nand U8635 (N_8635,N_8264,N_8302);
xnor U8636 (N_8636,N_8330,N_8400);
nor U8637 (N_8637,N_8265,N_8338);
or U8638 (N_8638,N_8409,N_8463);
or U8639 (N_8639,N_8440,N_8404);
nor U8640 (N_8640,N_8329,N_8375);
nand U8641 (N_8641,N_8323,N_8294);
or U8642 (N_8642,N_8494,N_8481);
and U8643 (N_8643,N_8265,N_8417);
nor U8644 (N_8644,N_8477,N_8489);
or U8645 (N_8645,N_8410,N_8487);
and U8646 (N_8646,N_8262,N_8317);
or U8647 (N_8647,N_8400,N_8271);
or U8648 (N_8648,N_8445,N_8321);
nand U8649 (N_8649,N_8464,N_8461);
nand U8650 (N_8650,N_8401,N_8394);
nor U8651 (N_8651,N_8411,N_8443);
or U8652 (N_8652,N_8349,N_8499);
or U8653 (N_8653,N_8460,N_8300);
and U8654 (N_8654,N_8397,N_8499);
or U8655 (N_8655,N_8414,N_8458);
nor U8656 (N_8656,N_8338,N_8436);
and U8657 (N_8657,N_8456,N_8310);
xnor U8658 (N_8658,N_8484,N_8363);
and U8659 (N_8659,N_8382,N_8388);
nor U8660 (N_8660,N_8309,N_8284);
or U8661 (N_8661,N_8320,N_8309);
and U8662 (N_8662,N_8338,N_8382);
nor U8663 (N_8663,N_8270,N_8396);
xnor U8664 (N_8664,N_8383,N_8430);
or U8665 (N_8665,N_8409,N_8264);
nand U8666 (N_8666,N_8250,N_8259);
or U8667 (N_8667,N_8305,N_8304);
nand U8668 (N_8668,N_8409,N_8393);
xor U8669 (N_8669,N_8353,N_8420);
or U8670 (N_8670,N_8409,N_8288);
or U8671 (N_8671,N_8255,N_8408);
and U8672 (N_8672,N_8274,N_8323);
and U8673 (N_8673,N_8482,N_8259);
nor U8674 (N_8674,N_8360,N_8270);
nor U8675 (N_8675,N_8325,N_8447);
nand U8676 (N_8676,N_8390,N_8373);
nand U8677 (N_8677,N_8446,N_8380);
xnor U8678 (N_8678,N_8332,N_8348);
or U8679 (N_8679,N_8493,N_8271);
nor U8680 (N_8680,N_8305,N_8464);
and U8681 (N_8681,N_8377,N_8264);
or U8682 (N_8682,N_8272,N_8341);
nand U8683 (N_8683,N_8391,N_8337);
nor U8684 (N_8684,N_8449,N_8380);
xnor U8685 (N_8685,N_8292,N_8300);
xor U8686 (N_8686,N_8449,N_8438);
nor U8687 (N_8687,N_8334,N_8438);
or U8688 (N_8688,N_8481,N_8297);
and U8689 (N_8689,N_8304,N_8259);
or U8690 (N_8690,N_8453,N_8438);
or U8691 (N_8691,N_8476,N_8373);
nand U8692 (N_8692,N_8383,N_8287);
or U8693 (N_8693,N_8347,N_8487);
and U8694 (N_8694,N_8402,N_8359);
nand U8695 (N_8695,N_8289,N_8453);
xnor U8696 (N_8696,N_8469,N_8455);
nor U8697 (N_8697,N_8347,N_8489);
xnor U8698 (N_8698,N_8347,N_8395);
xnor U8699 (N_8699,N_8458,N_8334);
nor U8700 (N_8700,N_8365,N_8346);
or U8701 (N_8701,N_8303,N_8401);
nand U8702 (N_8702,N_8381,N_8489);
nand U8703 (N_8703,N_8374,N_8322);
or U8704 (N_8704,N_8422,N_8462);
and U8705 (N_8705,N_8277,N_8286);
nor U8706 (N_8706,N_8416,N_8459);
nand U8707 (N_8707,N_8449,N_8347);
nor U8708 (N_8708,N_8493,N_8475);
xor U8709 (N_8709,N_8380,N_8404);
xnor U8710 (N_8710,N_8358,N_8300);
xnor U8711 (N_8711,N_8405,N_8316);
or U8712 (N_8712,N_8410,N_8485);
nand U8713 (N_8713,N_8476,N_8280);
nand U8714 (N_8714,N_8302,N_8261);
xor U8715 (N_8715,N_8466,N_8331);
or U8716 (N_8716,N_8261,N_8498);
nor U8717 (N_8717,N_8312,N_8394);
nand U8718 (N_8718,N_8313,N_8497);
and U8719 (N_8719,N_8311,N_8396);
nor U8720 (N_8720,N_8329,N_8295);
or U8721 (N_8721,N_8393,N_8430);
nand U8722 (N_8722,N_8356,N_8343);
nor U8723 (N_8723,N_8294,N_8413);
nor U8724 (N_8724,N_8435,N_8415);
or U8725 (N_8725,N_8454,N_8417);
and U8726 (N_8726,N_8325,N_8340);
nand U8727 (N_8727,N_8265,N_8363);
and U8728 (N_8728,N_8438,N_8282);
xor U8729 (N_8729,N_8277,N_8390);
nor U8730 (N_8730,N_8419,N_8369);
and U8731 (N_8731,N_8273,N_8333);
nand U8732 (N_8732,N_8257,N_8322);
nand U8733 (N_8733,N_8462,N_8273);
xnor U8734 (N_8734,N_8293,N_8307);
nand U8735 (N_8735,N_8335,N_8490);
nand U8736 (N_8736,N_8481,N_8308);
xnor U8737 (N_8737,N_8452,N_8258);
xnor U8738 (N_8738,N_8273,N_8459);
or U8739 (N_8739,N_8499,N_8460);
nand U8740 (N_8740,N_8425,N_8402);
nand U8741 (N_8741,N_8428,N_8292);
or U8742 (N_8742,N_8284,N_8432);
xor U8743 (N_8743,N_8295,N_8298);
or U8744 (N_8744,N_8411,N_8495);
and U8745 (N_8745,N_8350,N_8449);
and U8746 (N_8746,N_8471,N_8318);
or U8747 (N_8747,N_8330,N_8358);
and U8748 (N_8748,N_8423,N_8452);
and U8749 (N_8749,N_8303,N_8379);
xor U8750 (N_8750,N_8663,N_8573);
nand U8751 (N_8751,N_8654,N_8690);
nand U8752 (N_8752,N_8568,N_8622);
nand U8753 (N_8753,N_8714,N_8546);
or U8754 (N_8754,N_8574,N_8708);
or U8755 (N_8755,N_8631,N_8628);
nor U8756 (N_8756,N_8544,N_8731);
and U8757 (N_8757,N_8534,N_8600);
nand U8758 (N_8758,N_8715,N_8704);
or U8759 (N_8759,N_8709,N_8548);
nor U8760 (N_8760,N_8543,N_8612);
xnor U8761 (N_8761,N_8618,N_8555);
nand U8762 (N_8762,N_8685,N_8525);
or U8763 (N_8763,N_8660,N_8640);
nor U8764 (N_8764,N_8577,N_8616);
or U8765 (N_8765,N_8566,N_8695);
or U8766 (N_8766,N_8535,N_8641);
and U8767 (N_8767,N_8581,N_8729);
or U8768 (N_8768,N_8559,N_8686);
and U8769 (N_8769,N_8648,N_8739);
xor U8770 (N_8770,N_8516,N_8747);
nor U8771 (N_8771,N_8677,N_8716);
nor U8772 (N_8772,N_8596,N_8643);
nor U8773 (N_8773,N_8599,N_8552);
xnor U8774 (N_8774,N_8736,N_8586);
nand U8775 (N_8775,N_8579,N_8684);
and U8776 (N_8776,N_8523,N_8683);
nand U8777 (N_8777,N_8692,N_8706);
xnor U8778 (N_8778,N_8570,N_8567);
or U8779 (N_8779,N_8733,N_8623);
or U8780 (N_8780,N_8730,N_8538);
or U8781 (N_8781,N_8594,N_8595);
nor U8782 (N_8782,N_8531,N_8504);
and U8783 (N_8783,N_8703,N_8565);
nand U8784 (N_8784,N_8657,N_8537);
xnor U8785 (N_8785,N_8593,N_8655);
xnor U8786 (N_8786,N_8532,N_8591);
nand U8787 (N_8787,N_8673,N_8607);
nand U8788 (N_8788,N_8509,N_8521);
xnor U8789 (N_8789,N_8652,N_8676);
or U8790 (N_8790,N_8678,N_8584);
xor U8791 (N_8791,N_8635,N_8512);
nor U8792 (N_8792,N_8514,N_8545);
or U8793 (N_8793,N_8557,N_8642);
and U8794 (N_8794,N_8634,N_8601);
xnor U8795 (N_8795,N_8675,N_8734);
or U8796 (N_8796,N_8681,N_8705);
and U8797 (N_8797,N_8513,N_8728);
nand U8798 (N_8798,N_8667,N_8721);
nor U8799 (N_8799,N_8710,N_8614);
or U8800 (N_8800,N_8542,N_8701);
and U8801 (N_8801,N_8645,N_8719);
or U8802 (N_8802,N_8503,N_8603);
and U8803 (N_8803,N_8587,N_8602);
and U8804 (N_8804,N_8670,N_8554);
and U8805 (N_8805,N_8556,N_8528);
xnor U8806 (N_8806,N_8687,N_8679);
xor U8807 (N_8807,N_8621,N_8533);
nand U8808 (N_8808,N_8627,N_8529);
or U8809 (N_8809,N_8562,N_8735);
and U8810 (N_8810,N_8625,N_8725);
and U8811 (N_8811,N_8638,N_8620);
and U8812 (N_8812,N_8629,N_8720);
nor U8813 (N_8813,N_8507,N_8696);
xor U8814 (N_8814,N_8632,N_8576);
and U8815 (N_8815,N_8724,N_8742);
nand U8816 (N_8816,N_8658,N_8630);
and U8817 (N_8817,N_8501,N_8726);
or U8818 (N_8818,N_8646,N_8605);
or U8819 (N_8819,N_8745,N_8617);
nand U8820 (N_8820,N_8526,N_8547);
or U8821 (N_8821,N_8502,N_8589);
nor U8822 (N_8822,N_8519,N_8740);
nand U8823 (N_8823,N_8590,N_8737);
or U8824 (N_8824,N_8606,N_8610);
nor U8825 (N_8825,N_8717,N_8624);
nor U8826 (N_8826,N_8613,N_8636);
nand U8827 (N_8827,N_8553,N_8572);
nand U8828 (N_8828,N_8699,N_8522);
and U8829 (N_8829,N_8539,N_8609);
nor U8830 (N_8830,N_8588,N_8671);
xnor U8831 (N_8831,N_8580,N_8651);
nand U8832 (N_8832,N_8649,N_8561);
xnor U8833 (N_8833,N_8664,N_8639);
xor U8834 (N_8834,N_8650,N_8707);
nand U8835 (N_8835,N_8540,N_8647);
nor U8836 (N_8836,N_8691,N_8694);
nor U8837 (N_8837,N_8541,N_8672);
or U8838 (N_8838,N_8558,N_8511);
and U8839 (N_8839,N_8702,N_8530);
nand U8840 (N_8840,N_8659,N_8712);
or U8841 (N_8841,N_8551,N_8656);
and U8842 (N_8842,N_8536,N_8585);
nand U8843 (N_8843,N_8563,N_8680);
nand U8844 (N_8844,N_8688,N_8718);
nor U8845 (N_8845,N_8619,N_8744);
and U8846 (N_8846,N_8722,N_8527);
and U8847 (N_8847,N_8741,N_8746);
xnor U8848 (N_8848,N_8592,N_8711);
xnor U8849 (N_8849,N_8682,N_8578);
or U8850 (N_8850,N_8550,N_8698);
or U8851 (N_8851,N_8611,N_8723);
and U8852 (N_8852,N_8506,N_8669);
and U8853 (N_8853,N_8571,N_8560);
or U8854 (N_8854,N_8515,N_8524);
nand U8855 (N_8855,N_8564,N_8626);
and U8856 (N_8856,N_8665,N_8713);
and U8857 (N_8857,N_8582,N_8604);
nand U8858 (N_8858,N_8517,N_8732);
nor U8859 (N_8859,N_8661,N_8697);
xor U8860 (N_8860,N_8743,N_8644);
or U8861 (N_8861,N_8615,N_8637);
nor U8862 (N_8862,N_8738,N_8727);
xor U8863 (N_8863,N_8518,N_8569);
and U8864 (N_8864,N_8689,N_8505);
nand U8865 (N_8865,N_8674,N_8597);
nand U8866 (N_8866,N_8693,N_8700);
xnor U8867 (N_8867,N_8653,N_8508);
xor U8868 (N_8868,N_8662,N_8749);
xor U8869 (N_8869,N_8520,N_8549);
and U8870 (N_8870,N_8575,N_8598);
nand U8871 (N_8871,N_8500,N_8583);
or U8872 (N_8872,N_8668,N_8666);
nand U8873 (N_8873,N_8510,N_8748);
xor U8874 (N_8874,N_8608,N_8633);
nor U8875 (N_8875,N_8561,N_8679);
nor U8876 (N_8876,N_8555,N_8665);
or U8877 (N_8877,N_8719,N_8550);
and U8878 (N_8878,N_8749,N_8637);
or U8879 (N_8879,N_8528,N_8606);
and U8880 (N_8880,N_8660,N_8724);
nand U8881 (N_8881,N_8689,N_8642);
or U8882 (N_8882,N_8659,N_8662);
xnor U8883 (N_8883,N_8726,N_8525);
and U8884 (N_8884,N_8705,N_8526);
nor U8885 (N_8885,N_8691,N_8505);
nor U8886 (N_8886,N_8573,N_8591);
nand U8887 (N_8887,N_8743,N_8610);
nor U8888 (N_8888,N_8648,N_8534);
xor U8889 (N_8889,N_8645,N_8501);
nand U8890 (N_8890,N_8709,N_8634);
or U8891 (N_8891,N_8552,N_8676);
nor U8892 (N_8892,N_8742,N_8560);
nand U8893 (N_8893,N_8512,N_8667);
xor U8894 (N_8894,N_8536,N_8586);
nand U8895 (N_8895,N_8693,N_8638);
nand U8896 (N_8896,N_8526,N_8674);
and U8897 (N_8897,N_8655,N_8596);
xor U8898 (N_8898,N_8747,N_8698);
xnor U8899 (N_8899,N_8624,N_8555);
and U8900 (N_8900,N_8533,N_8697);
nor U8901 (N_8901,N_8726,N_8628);
or U8902 (N_8902,N_8644,N_8510);
and U8903 (N_8903,N_8664,N_8650);
xnor U8904 (N_8904,N_8657,N_8615);
nor U8905 (N_8905,N_8662,N_8631);
xnor U8906 (N_8906,N_8694,N_8522);
nor U8907 (N_8907,N_8560,N_8559);
xor U8908 (N_8908,N_8566,N_8685);
or U8909 (N_8909,N_8654,N_8559);
nand U8910 (N_8910,N_8504,N_8721);
and U8911 (N_8911,N_8577,N_8501);
xor U8912 (N_8912,N_8671,N_8737);
nand U8913 (N_8913,N_8513,N_8592);
xnor U8914 (N_8914,N_8719,N_8644);
xor U8915 (N_8915,N_8536,N_8518);
nor U8916 (N_8916,N_8686,N_8733);
nor U8917 (N_8917,N_8502,N_8543);
or U8918 (N_8918,N_8586,N_8533);
nor U8919 (N_8919,N_8698,N_8512);
and U8920 (N_8920,N_8607,N_8578);
nand U8921 (N_8921,N_8691,N_8557);
and U8922 (N_8922,N_8547,N_8648);
and U8923 (N_8923,N_8713,N_8599);
xor U8924 (N_8924,N_8562,N_8689);
nor U8925 (N_8925,N_8744,N_8617);
xor U8926 (N_8926,N_8690,N_8589);
nor U8927 (N_8927,N_8532,N_8533);
nor U8928 (N_8928,N_8583,N_8726);
nand U8929 (N_8929,N_8724,N_8706);
and U8930 (N_8930,N_8685,N_8693);
nor U8931 (N_8931,N_8659,N_8520);
nor U8932 (N_8932,N_8669,N_8642);
xnor U8933 (N_8933,N_8598,N_8665);
and U8934 (N_8934,N_8554,N_8631);
xnor U8935 (N_8935,N_8543,N_8577);
nor U8936 (N_8936,N_8593,N_8553);
nor U8937 (N_8937,N_8728,N_8643);
xnor U8938 (N_8938,N_8701,N_8519);
or U8939 (N_8939,N_8596,N_8540);
nor U8940 (N_8940,N_8587,N_8574);
nand U8941 (N_8941,N_8641,N_8676);
and U8942 (N_8942,N_8602,N_8551);
nand U8943 (N_8943,N_8724,N_8616);
and U8944 (N_8944,N_8639,N_8732);
and U8945 (N_8945,N_8546,N_8547);
or U8946 (N_8946,N_8601,N_8741);
and U8947 (N_8947,N_8708,N_8589);
xor U8948 (N_8948,N_8564,N_8716);
nor U8949 (N_8949,N_8605,N_8711);
and U8950 (N_8950,N_8644,N_8608);
nand U8951 (N_8951,N_8739,N_8735);
and U8952 (N_8952,N_8690,N_8580);
nor U8953 (N_8953,N_8713,N_8679);
or U8954 (N_8954,N_8544,N_8672);
xnor U8955 (N_8955,N_8561,N_8536);
nand U8956 (N_8956,N_8562,N_8733);
and U8957 (N_8957,N_8647,N_8719);
or U8958 (N_8958,N_8531,N_8712);
and U8959 (N_8959,N_8629,N_8613);
nand U8960 (N_8960,N_8642,N_8501);
nor U8961 (N_8961,N_8590,N_8537);
nand U8962 (N_8962,N_8731,N_8682);
nand U8963 (N_8963,N_8605,N_8638);
and U8964 (N_8964,N_8640,N_8630);
or U8965 (N_8965,N_8746,N_8538);
nand U8966 (N_8966,N_8548,N_8617);
xnor U8967 (N_8967,N_8734,N_8511);
xor U8968 (N_8968,N_8546,N_8502);
nand U8969 (N_8969,N_8624,N_8725);
or U8970 (N_8970,N_8549,N_8527);
nor U8971 (N_8971,N_8742,N_8740);
and U8972 (N_8972,N_8652,N_8726);
xnor U8973 (N_8973,N_8561,N_8735);
nand U8974 (N_8974,N_8613,N_8581);
and U8975 (N_8975,N_8711,N_8732);
xor U8976 (N_8976,N_8515,N_8674);
or U8977 (N_8977,N_8662,N_8677);
nand U8978 (N_8978,N_8520,N_8710);
and U8979 (N_8979,N_8611,N_8637);
and U8980 (N_8980,N_8710,N_8693);
and U8981 (N_8981,N_8513,N_8591);
or U8982 (N_8982,N_8621,N_8746);
or U8983 (N_8983,N_8534,N_8660);
nor U8984 (N_8984,N_8606,N_8599);
or U8985 (N_8985,N_8639,N_8613);
xnor U8986 (N_8986,N_8744,N_8528);
or U8987 (N_8987,N_8663,N_8562);
nand U8988 (N_8988,N_8628,N_8699);
and U8989 (N_8989,N_8565,N_8688);
or U8990 (N_8990,N_8712,N_8569);
and U8991 (N_8991,N_8698,N_8517);
nand U8992 (N_8992,N_8557,N_8540);
nor U8993 (N_8993,N_8569,N_8546);
and U8994 (N_8994,N_8615,N_8672);
nand U8995 (N_8995,N_8651,N_8502);
and U8996 (N_8996,N_8572,N_8684);
nor U8997 (N_8997,N_8652,N_8566);
nor U8998 (N_8998,N_8521,N_8562);
or U8999 (N_8999,N_8525,N_8631);
or U9000 (N_9000,N_8959,N_8938);
or U9001 (N_9001,N_8752,N_8870);
or U9002 (N_9002,N_8765,N_8824);
xnor U9003 (N_9003,N_8978,N_8966);
and U9004 (N_9004,N_8964,N_8796);
nand U9005 (N_9005,N_8857,N_8916);
nand U9006 (N_9006,N_8905,N_8887);
nor U9007 (N_9007,N_8790,N_8853);
and U9008 (N_9008,N_8903,N_8823);
and U9009 (N_9009,N_8838,N_8846);
nor U9010 (N_9010,N_8795,N_8917);
nor U9011 (N_9011,N_8979,N_8991);
xnor U9012 (N_9012,N_8884,N_8788);
and U9013 (N_9013,N_8922,N_8802);
or U9014 (N_9014,N_8815,N_8866);
or U9015 (N_9015,N_8986,N_8821);
or U9016 (N_9016,N_8988,N_8750);
or U9017 (N_9017,N_8924,N_8950);
or U9018 (N_9018,N_8787,N_8931);
xnor U9019 (N_9019,N_8832,N_8890);
and U9020 (N_9020,N_8797,N_8904);
nor U9021 (N_9021,N_8892,N_8830);
nor U9022 (N_9022,N_8920,N_8847);
nand U9023 (N_9023,N_8804,N_8818);
nand U9024 (N_9024,N_8994,N_8987);
nand U9025 (N_9025,N_8912,N_8863);
and U9026 (N_9026,N_8961,N_8755);
nand U9027 (N_9027,N_8980,N_8780);
or U9028 (N_9028,N_8955,N_8913);
and U9029 (N_9029,N_8899,N_8864);
nand U9030 (N_9030,N_8807,N_8891);
and U9031 (N_9031,N_8897,N_8845);
nand U9032 (N_9032,N_8881,N_8948);
or U9033 (N_9033,N_8839,N_8969);
nand U9034 (N_9034,N_8810,N_8825);
xnor U9035 (N_9035,N_8927,N_8761);
or U9036 (N_9036,N_8910,N_8889);
nand U9037 (N_9037,N_8935,N_8990);
nand U9038 (N_9038,N_8783,N_8933);
xor U9039 (N_9039,N_8768,N_8770);
nor U9040 (N_9040,N_8858,N_8972);
or U9041 (N_9041,N_8967,N_8831);
nand U9042 (N_9042,N_8751,N_8968);
xor U9043 (N_9043,N_8827,N_8775);
nand U9044 (N_9044,N_8936,N_8883);
xnor U9045 (N_9045,N_8940,N_8896);
xor U9046 (N_9046,N_8976,N_8840);
xnor U9047 (N_9047,N_8970,N_8753);
and U9048 (N_9048,N_8957,N_8981);
and U9049 (N_9049,N_8833,N_8829);
or U9050 (N_9050,N_8929,N_8814);
xor U9051 (N_9051,N_8805,N_8996);
xor U9052 (N_9052,N_8756,N_8867);
and U9053 (N_9053,N_8777,N_8862);
nor U9054 (N_9054,N_8868,N_8850);
xnor U9055 (N_9055,N_8811,N_8882);
or U9056 (N_9056,N_8836,N_8963);
xor U9057 (N_9057,N_8949,N_8791);
or U9058 (N_9058,N_8928,N_8789);
or U9059 (N_9059,N_8914,N_8943);
and U9060 (N_9060,N_8906,N_8794);
xor U9061 (N_9061,N_8997,N_8817);
and U9062 (N_9062,N_8806,N_8934);
nor U9063 (N_9063,N_8769,N_8983);
xor U9064 (N_9064,N_8757,N_8834);
xnor U9065 (N_9065,N_8860,N_8918);
and U9066 (N_9066,N_8841,N_8809);
nand U9067 (N_9067,N_8872,N_8898);
nand U9068 (N_9068,N_8992,N_8848);
nor U9069 (N_9069,N_8871,N_8953);
and U9070 (N_9070,N_8946,N_8754);
or U9071 (N_9071,N_8982,N_8902);
nand U9072 (N_9072,N_8861,N_8798);
and U9073 (N_9073,N_8965,N_8793);
xor U9074 (N_9074,N_8971,N_8820);
nand U9075 (N_9075,N_8958,N_8975);
xnor U9076 (N_9076,N_8759,N_8855);
or U9077 (N_9077,N_8803,N_8995);
nand U9078 (N_9078,N_8886,N_8763);
xnor U9079 (N_9079,N_8799,N_8937);
xnor U9080 (N_9080,N_8911,N_8771);
nor U9081 (N_9081,N_8888,N_8962);
xor U9082 (N_9082,N_8942,N_8900);
nand U9083 (N_9083,N_8837,N_8915);
or U9084 (N_9084,N_8784,N_8973);
and U9085 (N_9085,N_8843,N_8852);
xor U9086 (N_9086,N_8859,N_8951);
xnor U9087 (N_9087,N_8776,N_8813);
nand U9088 (N_9088,N_8781,N_8842);
and U9089 (N_9089,N_8774,N_8812);
and U9090 (N_9090,N_8879,N_8926);
or U9091 (N_9091,N_8954,N_8873);
nand U9092 (N_9092,N_8800,N_8849);
or U9093 (N_9093,N_8782,N_8826);
or U9094 (N_9094,N_8909,N_8808);
xor U9095 (N_9095,N_8944,N_8939);
nand U9096 (N_9096,N_8894,N_8977);
nor U9097 (N_9097,N_8758,N_8792);
nor U9098 (N_9098,N_8851,N_8773);
xor U9099 (N_9099,N_8772,N_8941);
or U9100 (N_9100,N_8878,N_8844);
or U9101 (N_9101,N_8766,N_8778);
nor U9102 (N_9102,N_8786,N_8801);
and U9103 (N_9103,N_8760,N_8856);
nand U9104 (N_9104,N_8998,N_8764);
or U9105 (N_9105,N_8785,N_8932);
or U9106 (N_9106,N_8989,N_8876);
xor U9107 (N_9107,N_8923,N_8999);
or U9108 (N_9108,N_8880,N_8819);
nor U9109 (N_9109,N_8895,N_8919);
nor U9110 (N_9110,N_8822,N_8762);
nor U9111 (N_9111,N_8835,N_8947);
and U9112 (N_9112,N_8875,N_8767);
xor U9113 (N_9113,N_8956,N_8877);
xor U9114 (N_9114,N_8893,N_8993);
xor U9115 (N_9115,N_8952,N_8930);
or U9116 (N_9116,N_8945,N_8816);
nand U9117 (N_9117,N_8960,N_8854);
xor U9118 (N_9118,N_8984,N_8779);
xor U9119 (N_9119,N_8885,N_8907);
nand U9120 (N_9120,N_8921,N_8985);
nand U9121 (N_9121,N_8901,N_8869);
and U9122 (N_9122,N_8908,N_8974);
or U9123 (N_9123,N_8925,N_8828);
xor U9124 (N_9124,N_8865,N_8874);
nand U9125 (N_9125,N_8942,N_8787);
xor U9126 (N_9126,N_8879,N_8832);
nand U9127 (N_9127,N_8809,N_8757);
or U9128 (N_9128,N_8932,N_8938);
nor U9129 (N_9129,N_8956,N_8826);
or U9130 (N_9130,N_8956,N_8973);
and U9131 (N_9131,N_8842,N_8808);
nand U9132 (N_9132,N_8940,N_8751);
and U9133 (N_9133,N_8967,N_8919);
nand U9134 (N_9134,N_8800,N_8979);
or U9135 (N_9135,N_8802,N_8936);
and U9136 (N_9136,N_8942,N_8774);
or U9137 (N_9137,N_8850,N_8983);
xor U9138 (N_9138,N_8751,N_8887);
nor U9139 (N_9139,N_8771,N_8867);
xnor U9140 (N_9140,N_8866,N_8919);
or U9141 (N_9141,N_8855,N_8935);
xnor U9142 (N_9142,N_8803,N_8950);
nand U9143 (N_9143,N_8916,N_8940);
and U9144 (N_9144,N_8866,N_8880);
or U9145 (N_9145,N_8774,N_8979);
nor U9146 (N_9146,N_8949,N_8969);
and U9147 (N_9147,N_8918,N_8893);
nand U9148 (N_9148,N_8983,N_8758);
nand U9149 (N_9149,N_8812,N_8986);
nor U9150 (N_9150,N_8802,N_8982);
nand U9151 (N_9151,N_8982,N_8809);
xor U9152 (N_9152,N_8775,N_8830);
or U9153 (N_9153,N_8960,N_8770);
nand U9154 (N_9154,N_8769,N_8919);
or U9155 (N_9155,N_8794,N_8806);
xnor U9156 (N_9156,N_8941,N_8912);
xnor U9157 (N_9157,N_8918,N_8856);
nor U9158 (N_9158,N_8975,N_8905);
nor U9159 (N_9159,N_8811,N_8919);
and U9160 (N_9160,N_8909,N_8821);
xor U9161 (N_9161,N_8842,N_8902);
or U9162 (N_9162,N_8830,N_8803);
nand U9163 (N_9163,N_8900,N_8903);
nor U9164 (N_9164,N_8908,N_8750);
nand U9165 (N_9165,N_8822,N_8926);
and U9166 (N_9166,N_8878,N_8816);
and U9167 (N_9167,N_8904,N_8830);
xor U9168 (N_9168,N_8812,N_8813);
or U9169 (N_9169,N_8844,N_8975);
and U9170 (N_9170,N_8847,N_8869);
xnor U9171 (N_9171,N_8876,N_8756);
nand U9172 (N_9172,N_8767,N_8986);
nor U9173 (N_9173,N_8764,N_8934);
xnor U9174 (N_9174,N_8901,N_8935);
nand U9175 (N_9175,N_8936,N_8781);
and U9176 (N_9176,N_8803,N_8762);
nand U9177 (N_9177,N_8829,N_8996);
xnor U9178 (N_9178,N_8801,N_8797);
nor U9179 (N_9179,N_8939,N_8893);
and U9180 (N_9180,N_8831,N_8924);
nand U9181 (N_9181,N_8969,N_8850);
and U9182 (N_9182,N_8938,N_8948);
xnor U9183 (N_9183,N_8900,N_8925);
nor U9184 (N_9184,N_8818,N_8933);
or U9185 (N_9185,N_8851,N_8845);
xnor U9186 (N_9186,N_8797,N_8906);
and U9187 (N_9187,N_8788,N_8999);
and U9188 (N_9188,N_8820,N_8904);
xnor U9189 (N_9189,N_8924,N_8913);
and U9190 (N_9190,N_8750,N_8902);
xnor U9191 (N_9191,N_8983,N_8837);
and U9192 (N_9192,N_8937,N_8808);
and U9193 (N_9193,N_8922,N_8784);
or U9194 (N_9194,N_8890,N_8752);
nand U9195 (N_9195,N_8789,N_8893);
nor U9196 (N_9196,N_8936,N_8969);
and U9197 (N_9197,N_8791,N_8942);
nor U9198 (N_9198,N_8755,N_8971);
nor U9199 (N_9199,N_8988,N_8830);
and U9200 (N_9200,N_8899,N_8901);
nand U9201 (N_9201,N_8834,N_8841);
nand U9202 (N_9202,N_8774,N_8835);
or U9203 (N_9203,N_8937,N_8942);
nand U9204 (N_9204,N_8795,N_8900);
nor U9205 (N_9205,N_8936,N_8756);
xor U9206 (N_9206,N_8811,N_8771);
nand U9207 (N_9207,N_8867,N_8872);
nor U9208 (N_9208,N_8938,N_8861);
nand U9209 (N_9209,N_8760,N_8758);
nor U9210 (N_9210,N_8835,N_8846);
xnor U9211 (N_9211,N_8828,N_8907);
xor U9212 (N_9212,N_8758,N_8923);
or U9213 (N_9213,N_8913,N_8948);
or U9214 (N_9214,N_8791,N_8758);
or U9215 (N_9215,N_8912,N_8879);
xor U9216 (N_9216,N_8803,N_8789);
nand U9217 (N_9217,N_8911,N_8941);
nor U9218 (N_9218,N_8992,N_8995);
or U9219 (N_9219,N_8813,N_8852);
or U9220 (N_9220,N_8867,N_8948);
nand U9221 (N_9221,N_8774,N_8960);
nor U9222 (N_9222,N_8897,N_8756);
nor U9223 (N_9223,N_8939,N_8789);
xnor U9224 (N_9224,N_8946,N_8988);
or U9225 (N_9225,N_8919,N_8934);
and U9226 (N_9226,N_8811,N_8926);
nor U9227 (N_9227,N_8889,N_8965);
nand U9228 (N_9228,N_8831,N_8777);
nand U9229 (N_9229,N_8772,N_8916);
nand U9230 (N_9230,N_8976,N_8985);
or U9231 (N_9231,N_8915,N_8751);
nand U9232 (N_9232,N_8956,N_8797);
xnor U9233 (N_9233,N_8868,N_8941);
nor U9234 (N_9234,N_8751,N_8877);
or U9235 (N_9235,N_8961,N_8845);
or U9236 (N_9236,N_8931,N_8838);
xor U9237 (N_9237,N_8808,N_8831);
nand U9238 (N_9238,N_8927,N_8780);
nor U9239 (N_9239,N_8928,N_8823);
nor U9240 (N_9240,N_8941,N_8946);
or U9241 (N_9241,N_8886,N_8812);
nand U9242 (N_9242,N_8789,N_8783);
nand U9243 (N_9243,N_8786,N_8965);
nor U9244 (N_9244,N_8977,N_8857);
nand U9245 (N_9245,N_8934,N_8921);
or U9246 (N_9246,N_8750,N_8916);
and U9247 (N_9247,N_8951,N_8887);
and U9248 (N_9248,N_8828,N_8764);
nand U9249 (N_9249,N_8768,N_8806);
nor U9250 (N_9250,N_9154,N_9119);
xnor U9251 (N_9251,N_9141,N_9082);
nand U9252 (N_9252,N_9213,N_9179);
and U9253 (N_9253,N_9078,N_9035);
nand U9254 (N_9254,N_9135,N_9232);
nor U9255 (N_9255,N_9240,N_9113);
nor U9256 (N_9256,N_9199,N_9087);
xor U9257 (N_9257,N_9060,N_9027);
nor U9258 (N_9258,N_9166,N_9136);
nand U9259 (N_9259,N_9129,N_9067);
and U9260 (N_9260,N_9002,N_9244);
or U9261 (N_9261,N_9152,N_9132);
nor U9262 (N_9262,N_9045,N_9009);
xnor U9263 (N_9263,N_9193,N_9014);
xor U9264 (N_9264,N_9163,N_9085);
nor U9265 (N_9265,N_9249,N_9194);
and U9266 (N_9266,N_9025,N_9076);
nand U9267 (N_9267,N_9040,N_9219);
or U9268 (N_9268,N_9112,N_9061);
nor U9269 (N_9269,N_9241,N_9050);
nand U9270 (N_9270,N_9070,N_9042);
nand U9271 (N_9271,N_9115,N_9097);
or U9272 (N_9272,N_9168,N_9186);
or U9273 (N_9273,N_9195,N_9030);
nand U9274 (N_9274,N_9073,N_9142);
nand U9275 (N_9275,N_9234,N_9124);
and U9276 (N_9276,N_9196,N_9075);
nor U9277 (N_9277,N_9008,N_9150);
xor U9278 (N_9278,N_9096,N_9077);
and U9279 (N_9279,N_9043,N_9010);
or U9280 (N_9280,N_9182,N_9031);
nand U9281 (N_9281,N_9224,N_9012);
xnor U9282 (N_9282,N_9208,N_9211);
and U9283 (N_9283,N_9047,N_9165);
nand U9284 (N_9284,N_9210,N_9004);
and U9285 (N_9285,N_9086,N_9094);
xnor U9286 (N_9286,N_9079,N_9206);
and U9287 (N_9287,N_9198,N_9169);
xnor U9288 (N_9288,N_9083,N_9226);
or U9289 (N_9289,N_9118,N_9049);
or U9290 (N_9290,N_9170,N_9181);
nand U9291 (N_9291,N_9120,N_9156);
or U9292 (N_9292,N_9029,N_9177);
and U9293 (N_9293,N_9055,N_9143);
nand U9294 (N_9294,N_9091,N_9233);
or U9295 (N_9295,N_9236,N_9242);
or U9296 (N_9296,N_9167,N_9039);
nor U9297 (N_9297,N_9011,N_9157);
or U9298 (N_9298,N_9117,N_9140);
or U9299 (N_9299,N_9158,N_9056);
and U9300 (N_9300,N_9229,N_9122);
or U9301 (N_9301,N_9048,N_9053);
and U9302 (N_9302,N_9172,N_9064);
and U9303 (N_9303,N_9081,N_9066);
and U9304 (N_9304,N_9243,N_9051);
and U9305 (N_9305,N_9036,N_9088);
xnor U9306 (N_9306,N_9028,N_9247);
or U9307 (N_9307,N_9099,N_9024);
nor U9308 (N_9308,N_9216,N_9190);
or U9309 (N_9309,N_9217,N_9006);
xor U9310 (N_9310,N_9175,N_9022);
nand U9311 (N_9311,N_9018,N_9130);
xor U9312 (N_9312,N_9220,N_9218);
nand U9313 (N_9313,N_9200,N_9000);
xor U9314 (N_9314,N_9069,N_9215);
nor U9315 (N_9315,N_9013,N_9245);
nor U9316 (N_9316,N_9105,N_9209);
and U9317 (N_9317,N_9071,N_9133);
or U9318 (N_9318,N_9100,N_9180);
nor U9319 (N_9319,N_9178,N_9107);
nor U9320 (N_9320,N_9202,N_9015);
nor U9321 (N_9321,N_9225,N_9041);
nor U9322 (N_9322,N_9020,N_9212);
or U9323 (N_9323,N_9222,N_9093);
nor U9324 (N_9324,N_9111,N_9161);
xnor U9325 (N_9325,N_9235,N_9110);
and U9326 (N_9326,N_9034,N_9058);
nor U9327 (N_9327,N_9054,N_9159);
nor U9328 (N_9328,N_9204,N_9080);
xnor U9329 (N_9329,N_9095,N_9173);
and U9330 (N_9330,N_9231,N_9023);
and U9331 (N_9331,N_9189,N_9021);
or U9332 (N_9332,N_9038,N_9003);
and U9333 (N_9333,N_9155,N_9148);
or U9334 (N_9334,N_9104,N_9139);
or U9335 (N_9335,N_9188,N_9065);
nand U9336 (N_9336,N_9239,N_9185);
nor U9337 (N_9337,N_9123,N_9151);
nand U9338 (N_9338,N_9033,N_9074);
and U9339 (N_9339,N_9171,N_9203);
or U9340 (N_9340,N_9214,N_9164);
or U9341 (N_9341,N_9153,N_9126);
xnor U9342 (N_9342,N_9187,N_9090);
nand U9343 (N_9343,N_9052,N_9059);
nor U9344 (N_9344,N_9138,N_9089);
nor U9345 (N_9345,N_9005,N_9197);
and U9346 (N_9346,N_9191,N_9192);
nand U9347 (N_9347,N_9230,N_9062);
xor U9348 (N_9348,N_9037,N_9121);
nand U9349 (N_9349,N_9145,N_9174);
nor U9350 (N_9350,N_9246,N_9221);
or U9351 (N_9351,N_9044,N_9127);
and U9352 (N_9352,N_9101,N_9223);
nand U9353 (N_9353,N_9092,N_9184);
xor U9354 (N_9354,N_9001,N_9134);
xor U9355 (N_9355,N_9207,N_9084);
xnor U9356 (N_9356,N_9114,N_9228);
xnor U9357 (N_9357,N_9019,N_9046);
nor U9358 (N_9358,N_9125,N_9237);
nand U9359 (N_9359,N_9103,N_9109);
or U9360 (N_9360,N_9147,N_9144);
nor U9361 (N_9361,N_9205,N_9201);
nand U9362 (N_9362,N_9162,N_9026);
and U9363 (N_9363,N_9063,N_9072);
nand U9364 (N_9364,N_9007,N_9102);
and U9365 (N_9365,N_9227,N_9098);
or U9366 (N_9366,N_9183,N_9116);
nor U9367 (N_9367,N_9248,N_9068);
nor U9368 (N_9368,N_9108,N_9057);
or U9369 (N_9369,N_9032,N_9128);
or U9370 (N_9370,N_9131,N_9016);
nor U9371 (N_9371,N_9137,N_9146);
and U9372 (N_9372,N_9017,N_9149);
and U9373 (N_9373,N_9160,N_9176);
and U9374 (N_9374,N_9106,N_9238);
xor U9375 (N_9375,N_9191,N_9045);
nand U9376 (N_9376,N_9228,N_9005);
and U9377 (N_9377,N_9142,N_9074);
nor U9378 (N_9378,N_9063,N_9152);
nor U9379 (N_9379,N_9160,N_9104);
nand U9380 (N_9380,N_9141,N_9238);
nand U9381 (N_9381,N_9187,N_9203);
nor U9382 (N_9382,N_9224,N_9227);
or U9383 (N_9383,N_9204,N_9249);
and U9384 (N_9384,N_9020,N_9045);
or U9385 (N_9385,N_9212,N_9053);
nor U9386 (N_9386,N_9058,N_9145);
or U9387 (N_9387,N_9210,N_9098);
and U9388 (N_9388,N_9139,N_9182);
nor U9389 (N_9389,N_9222,N_9244);
and U9390 (N_9390,N_9031,N_9079);
nor U9391 (N_9391,N_9000,N_9206);
and U9392 (N_9392,N_9208,N_9195);
or U9393 (N_9393,N_9146,N_9085);
and U9394 (N_9394,N_9160,N_9015);
or U9395 (N_9395,N_9054,N_9132);
nor U9396 (N_9396,N_9090,N_9234);
nand U9397 (N_9397,N_9052,N_9173);
xor U9398 (N_9398,N_9076,N_9017);
or U9399 (N_9399,N_9195,N_9063);
xor U9400 (N_9400,N_9079,N_9220);
xor U9401 (N_9401,N_9095,N_9062);
or U9402 (N_9402,N_9065,N_9183);
xor U9403 (N_9403,N_9184,N_9149);
xnor U9404 (N_9404,N_9044,N_9231);
nand U9405 (N_9405,N_9129,N_9032);
nand U9406 (N_9406,N_9209,N_9020);
xnor U9407 (N_9407,N_9112,N_9050);
or U9408 (N_9408,N_9113,N_9048);
and U9409 (N_9409,N_9136,N_9118);
xor U9410 (N_9410,N_9187,N_9174);
nor U9411 (N_9411,N_9052,N_9011);
nor U9412 (N_9412,N_9197,N_9208);
and U9413 (N_9413,N_9245,N_9106);
nand U9414 (N_9414,N_9174,N_9212);
nand U9415 (N_9415,N_9162,N_9161);
nand U9416 (N_9416,N_9077,N_9057);
and U9417 (N_9417,N_9077,N_9234);
or U9418 (N_9418,N_9113,N_9001);
and U9419 (N_9419,N_9098,N_9129);
nor U9420 (N_9420,N_9160,N_9142);
nor U9421 (N_9421,N_9103,N_9193);
nor U9422 (N_9422,N_9058,N_9064);
nor U9423 (N_9423,N_9045,N_9032);
nand U9424 (N_9424,N_9236,N_9225);
and U9425 (N_9425,N_9152,N_9182);
or U9426 (N_9426,N_9036,N_9027);
nand U9427 (N_9427,N_9074,N_9140);
and U9428 (N_9428,N_9083,N_9232);
and U9429 (N_9429,N_9010,N_9190);
and U9430 (N_9430,N_9085,N_9225);
nor U9431 (N_9431,N_9207,N_9225);
nor U9432 (N_9432,N_9231,N_9060);
nor U9433 (N_9433,N_9089,N_9010);
and U9434 (N_9434,N_9107,N_9104);
or U9435 (N_9435,N_9086,N_9024);
nand U9436 (N_9436,N_9219,N_9248);
nor U9437 (N_9437,N_9014,N_9092);
or U9438 (N_9438,N_9188,N_9115);
and U9439 (N_9439,N_9066,N_9133);
nand U9440 (N_9440,N_9228,N_9020);
and U9441 (N_9441,N_9045,N_9227);
nand U9442 (N_9442,N_9189,N_9243);
nor U9443 (N_9443,N_9155,N_9074);
or U9444 (N_9444,N_9197,N_9105);
nor U9445 (N_9445,N_9032,N_9088);
and U9446 (N_9446,N_9144,N_9167);
nand U9447 (N_9447,N_9176,N_9246);
nor U9448 (N_9448,N_9102,N_9016);
or U9449 (N_9449,N_9097,N_9017);
nand U9450 (N_9450,N_9105,N_9137);
xor U9451 (N_9451,N_9203,N_9131);
nand U9452 (N_9452,N_9226,N_9125);
nand U9453 (N_9453,N_9243,N_9144);
and U9454 (N_9454,N_9243,N_9034);
nand U9455 (N_9455,N_9249,N_9239);
and U9456 (N_9456,N_9072,N_9102);
nand U9457 (N_9457,N_9215,N_9107);
and U9458 (N_9458,N_9219,N_9118);
nor U9459 (N_9459,N_9134,N_9085);
nand U9460 (N_9460,N_9002,N_9050);
and U9461 (N_9461,N_9063,N_9248);
nand U9462 (N_9462,N_9075,N_9074);
or U9463 (N_9463,N_9197,N_9058);
or U9464 (N_9464,N_9233,N_9141);
nand U9465 (N_9465,N_9134,N_9058);
or U9466 (N_9466,N_9003,N_9090);
and U9467 (N_9467,N_9188,N_9137);
or U9468 (N_9468,N_9189,N_9064);
or U9469 (N_9469,N_9015,N_9186);
xnor U9470 (N_9470,N_9029,N_9063);
nor U9471 (N_9471,N_9240,N_9131);
nand U9472 (N_9472,N_9201,N_9066);
nor U9473 (N_9473,N_9175,N_9152);
and U9474 (N_9474,N_9078,N_9033);
xnor U9475 (N_9475,N_9204,N_9179);
or U9476 (N_9476,N_9078,N_9094);
and U9477 (N_9477,N_9089,N_9220);
and U9478 (N_9478,N_9002,N_9098);
nand U9479 (N_9479,N_9091,N_9086);
nand U9480 (N_9480,N_9055,N_9099);
or U9481 (N_9481,N_9180,N_9059);
nor U9482 (N_9482,N_9130,N_9029);
or U9483 (N_9483,N_9066,N_9064);
nor U9484 (N_9484,N_9124,N_9243);
xor U9485 (N_9485,N_9114,N_9037);
nor U9486 (N_9486,N_9156,N_9189);
nand U9487 (N_9487,N_9188,N_9012);
or U9488 (N_9488,N_9122,N_9144);
nor U9489 (N_9489,N_9176,N_9015);
nor U9490 (N_9490,N_9160,N_9025);
and U9491 (N_9491,N_9162,N_9124);
xnor U9492 (N_9492,N_9218,N_9191);
nand U9493 (N_9493,N_9112,N_9192);
nand U9494 (N_9494,N_9029,N_9073);
and U9495 (N_9495,N_9187,N_9078);
xor U9496 (N_9496,N_9115,N_9144);
nand U9497 (N_9497,N_9044,N_9087);
nand U9498 (N_9498,N_9101,N_9099);
or U9499 (N_9499,N_9072,N_9210);
and U9500 (N_9500,N_9461,N_9297);
nor U9501 (N_9501,N_9299,N_9463);
and U9502 (N_9502,N_9376,N_9497);
nand U9503 (N_9503,N_9320,N_9306);
or U9504 (N_9504,N_9250,N_9340);
or U9505 (N_9505,N_9490,N_9401);
or U9506 (N_9506,N_9296,N_9454);
xor U9507 (N_9507,N_9305,N_9325);
xor U9508 (N_9508,N_9479,N_9397);
nand U9509 (N_9509,N_9272,N_9267);
nand U9510 (N_9510,N_9334,N_9378);
and U9511 (N_9511,N_9315,N_9492);
and U9512 (N_9512,N_9390,N_9486);
or U9513 (N_9513,N_9285,N_9482);
nand U9514 (N_9514,N_9287,N_9438);
xor U9515 (N_9515,N_9258,N_9485);
xnor U9516 (N_9516,N_9350,N_9295);
nor U9517 (N_9517,N_9427,N_9270);
nand U9518 (N_9518,N_9435,N_9333);
nor U9519 (N_9519,N_9478,N_9256);
or U9520 (N_9520,N_9382,N_9304);
or U9521 (N_9521,N_9419,N_9418);
nor U9522 (N_9522,N_9434,N_9493);
nand U9523 (N_9523,N_9322,N_9355);
or U9524 (N_9524,N_9269,N_9293);
or U9525 (N_9525,N_9360,N_9459);
xor U9526 (N_9526,N_9465,N_9458);
and U9527 (N_9527,N_9303,N_9271);
or U9528 (N_9528,N_9341,N_9375);
xnor U9529 (N_9529,N_9289,N_9354);
and U9530 (N_9530,N_9346,N_9424);
nor U9531 (N_9531,N_9327,N_9413);
xor U9532 (N_9532,N_9426,N_9409);
nand U9533 (N_9533,N_9311,N_9398);
nor U9534 (N_9534,N_9301,N_9282);
xor U9535 (N_9535,N_9336,N_9453);
xnor U9536 (N_9536,N_9488,N_9276);
or U9537 (N_9537,N_9475,N_9395);
nand U9538 (N_9538,N_9281,N_9323);
and U9539 (N_9539,N_9348,N_9474);
and U9540 (N_9540,N_9286,N_9337);
nor U9541 (N_9541,N_9288,N_9481);
or U9542 (N_9542,N_9432,N_9344);
and U9543 (N_9543,N_9469,N_9464);
nor U9544 (N_9544,N_9471,N_9472);
nand U9545 (N_9545,N_9477,N_9406);
and U9546 (N_9546,N_9410,N_9319);
or U9547 (N_9547,N_9266,N_9415);
xor U9548 (N_9548,N_9317,N_9483);
nand U9549 (N_9549,N_9309,N_9407);
xnor U9550 (N_9550,N_9430,N_9447);
nor U9551 (N_9551,N_9396,N_9405);
nor U9552 (N_9552,N_9314,N_9455);
or U9553 (N_9553,N_9496,N_9357);
and U9554 (N_9554,N_9274,N_9391);
xnor U9555 (N_9555,N_9307,N_9462);
nor U9556 (N_9556,N_9313,N_9489);
xnor U9557 (N_9557,N_9416,N_9362);
xor U9558 (N_9558,N_9300,N_9470);
nor U9559 (N_9559,N_9252,N_9425);
xor U9560 (N_9560,N_9429,N_9371);
and U9561 (N_9561,N_9253,N_9403);
nor U9562 (N_9562,N_9491,N_9468);
and U9563 (N_9563,N_9411,N_9291);
nor U9564 (N_9564,N_9329,N_9404);
xor U9565 (N_9565,N_9321,N_9440);
nand U9566 (N_9566,N_9265,N_9417);
nor U9567 (N_9567,N_9484,N_9412);
nor U9568 (N_9568,N_9308,N_9449);
xor U9569 (N_9569,N_9456,N_9251);
nand U9570 (N_9570,N_9367,N_9294);
or U9571 (N_9571,N_9448,N_9358);
and U9572 (N_9572,N_9431,N_9439);
xor U9573 (N_9573,N_9373,N_9298);
or U9574 (N_9574,N_9441,N_9264);
nor U9575 (N_9575,N_9437,N_9275);
and U9576 (N_9576,N_9364,N_9380);
xor U9577 (N_9577,N_9460,N_9273);
nand U9578 (N_9578,N_9332,N_9399);
and U9579 (N_9579,N_9292,N_9389);
and U9580 (N_9580,N_9339,N_9284);
or U9581 (N_9581,N_9283,N_9318);
nand U9582 (N_9582,N_9259,N_9347);
and U9583 (N_9583,N_9324,N_9342);
or U9584 (N_9584,N_9352,N_9445);
or U9585 (N_9585,N_9343,N_9423);
xnor U9586 (N_9586,N_9451,N_9383);
nand U9587 (N_9587,N_9302,N_9280);
and U9588 (N_9588,N_9495,N_9457);
nor U9589 (N_9589,N_9494,N_9385);
nor U9590 (N_9590,N_9372,N_9436);
or U9591 (N_9591,N_9349,N_9330);
nor U9592 (N_9592,N_9310,N_9254);
nor U9593 (N_9593,N_9408,N_9366);
xor U9594 (N_9594,N_9277,N_9498);
nand U9595 (N_9595,N_9255,N_9331);
or U9596 (N_9596,N_9368,N_9466);
or U9597 (N_9597,N_9290,N_9421);
xnor U9598 (N_9598,N_9351,N_9369);
or U9599 (N_9599,N_9381,N_9261);
or U9600 (N_9600,N_9420,N_9386);
nor U9601 (N_9601,N_9388,N_9402);
and U9602 (N_9602,N_9363,N_9268);
nor U9603 (N_9603,N_9326,N_9353);
and U9604 (N_9604,N_9476,N_9361);
xor U9605 (N_9605,N_9356,N_9278);
xnor U9606 (N_9606,N_9257,N_9328);
and U9607 (N_9607,N_9473,N_9392);
xnor U9608 (N_9608,N_9452,N_9487);
or U9609 (N_9609,N_9480,N_9365);
xnor U9610 (N_9610,N_9433,N_9359);
nand U9611 (N_9611,N_9377,N_9316);
and U9612 (N_9612,N_9387,N_9374);
xor U9613 (N_9613,N_9338,N_9370);
and U9614 (N_9614,N_9260,N_9422);
nor U9615 (N_9615,N_9428,N_9444);
xnor U9616 (N_9616,N_9467,N_9414);
nand U9617 (N_9617,N_9263,N_9499);
and U9618 (N_9618,N_9450,N_9393);
nor U9619 (N_9619,N_9384,N_9400);
xnor U9620 (N_9620,N_9345,N_9279);
or U9621 (N_9621,N_9335,N_9443);
and U9622 (N_9622,N_9312,N_9394);
or U9623 (N_9623,N_9442,N_9446);
xor U9624 (N_9624,N_9262,N_9379);
xor U9625 (N_9625,N_9263,N_9269);
and U9626 (N_9626,N_9393,N_9361);
and U9627 (N_9627,N_9350,N_9368);
nor U9628 (N_9628,N_9435,N_9290);
and U9629 (N_9629,N_9329,N_9461);
nor U9630 (N_9630,N_9393,N_9422);
xor U9631 (N_9631,N_9254,N_9297);
nand U9632 (N_9632,N_9334,N_9455);
and U9633 (N_9633,N_9443,N_9357);
nand U9634 (N_9634,N_9396,N_9388);
nor U9635 (N_9635,N_9437,N_9293);
xnor U9636 (N_9636,N_9440,N_9445);
nor U9637 (N_9637,N_9444,N_9409);
nand U9638 (N_9638,N_9275,N_9494);
nor U9639 (N_9639,N_9282,N_9250);
nor U9640 (N_9640,N_9408,N_9377);
nand U9641 (N_9641,N_9433,N_9259);
xnor U9642 (N_9642,N_9332,N_9360);
or U9643 (N_9643,N_9386,N_9301);
nor U9644 (N_9644,N_9457,N_9259);
and U9645 (N_9645,N_9277,N_9280);
or U9646 (N_9646,N_9476,N_9315);
or U9647 (N_9647,N_9473,N_9378);
nand U9648 (N_9648,N_9413,N_9467);
and U9649 (N_9649,N_9435,N_9339);
xor U9650 (N_9650,N_9286,N_9401);
and U9651 (N_9651,N_9477,N_9270);
xnor U9652 (N_9652,N_9442,N_9461);
nand U9653 (N_9653,N_9461,N_9439);
nand U9654 (N_9654,N_9255,N_9289);
and U9655 (N_9655,N_9415,N_9286);
xnor U9656 (N_9656,N_9428,N_9479);
nor U9657 (N_9657,N_9455,N_9403);
and U9658 (N_9658,N_9440,N_9448);
xnor U9659 (N_9659,N_9349,N_9285);
xnor U9660 (N_9660,N_9360,N_9280);
nor U9661 (N_9661,N_9321,N_9346);
xor U9662 (N_9662,N_9479,N_9331);
nor U9663 (N_9663,N_9404,N_9319);
nor U9664 (N_9664,N_9434,N_9460);
or U9665 (N_9665,N_9292,N_9341);
nor U9666 (N_9666,N_9296,N_9451);
nor U9667 (N_9667,N_9391,N_9460);
nand U9668 (N_9668,N_9465,N_9368);
nor U9669 (N_9669,N_9487,N_9440);
xnor U9670 (N_9670,N_9401,N_9489);
xor U9671 (N_9671,N_9344,N_9437);
nand U9672 (N_9672,N_9250,N_9354);
xor U9673 (N_9673,N_9469,N_9409);
nand U9674 (N_9674,N_9299,N_9276);
xnor U9675 (N_9675,N_9324,N_9318);
xnor U9676 (N_9676,N_9276,N_9314);
nor U9677 (N_9677,N_9440,N_9300);
and U9678 (N_9678,N_9267,N_9447);
xnor U9679 (N_9679,N_9354,N_9468);
and U9680 (N_9680,N_9331,N_9478);
or U9681 (N_9681,N_9433,N_9311);
and U9682 (N_9682,N_9485,N_9284);
and U9683 (N_9683,N_9396,N_9486);
and U9684 (N_9684,N_9467,N_9268);
xnor U9685 (N_9685,N_9373,N_9275);
nor U9686 (N_9686,N_9389,N_9495);
nor U9687 (N_9687,N_9461,N_9253);
or U9688 (N_9688,N_9268,N_9453);
xor U9689 (N_9689,N_9372,N_9342);
nor U9690 (N_9690,N_9376,N_9251);
nand U9691 (N_9691,N_9478,N_9329);
xor U9692 (N_9692,N_9307,N_9435);
or U9693 (N_9693,N_9437,N_9273);
or U9694 (N_9694,N_9392,N_9424);
and U9695 (N_9695,N_9400,N_9444);
and U9696 (N_9696,N_9358,N_9371);
nor U9697 (N_9697,N_9302,N_9408);
nor U9698 (N_9698,N_9487,N_9398);
or U9699 (N_9699,N_9402,N_9449);
or U9700 (N_9700,N_9313,N_9491);
nor U9701 (N_9701,N_9256,N_9485);
and U9702 (N_9702,N_9440,N_9411);
nand U9703 (N_9703,N_9447,N_9458);
or U9704 (N_9704,N_9252,N_9275);
nor U9705 (N_9705,N_9344,N_9333);
or U9706 (N_9706,N_9478,N_9447);
and U9707 (N_9707,N_9258,N_9427);
nor U9708 (N_9708,N_9434,N_9311);
or U9709 (N_9709,N_9321,N_9271);
xor U9710 (N_9710,N_9360,N_9480);
xnor U9711 (N_9711,N_9375,N_9498);
or U9712 (N_9712,N_9308,N_9294);
or U9713 (N_9713,N_9402,N_9315);
nand U9714 (N_9714,N_9253,N_9383);
xnor U9715 (N_9715,N_9421,N_9349);
xor U9716 (N_9716,N_9305,N_9487);
nand U9717 (N_9717,N_9462,N_9429);
nand U9718 (N_9718,N_9292,N_9446);
xnor U9719 (N_9719,N_9394,N_9380);
nor U9720 (N_9720,N_9402,N_9494);
or U9721 (N_9721,N_9418,N_9392);
nand U9722 (N_9722,N_9258,N_9428);
or U9723 (N_9723,N_9301,N_9399);
xor U9724 (N_9724,N_9277,N_9455);
or U9725 (N_9725,N_9473,N_9323);
nand U9726 (N_9726,N_9459,N_9280);
xor U9727 (N_9727,N_9364,N_9465);
or U9728 (N_9728,N_9250,N_9267);
xnor U9729 (N_9729,N_9265,N_9491);
xnor U9730 (N_9730,N_9464,N_9383);
or U9731 (N_9731,N_9317,N_9295);
xnor U9732 (N_9732,N_9439,N_9258);
nor U9733 (N_9733,N_9333,N_9354);
or U9734 (N_9734,N_9396,N_9364);
xor U9735 (N_9735,N_9450,N_9403);
nor U9736 (N_9736,N_9359,N_9448);
or U9737 (N_9737,N_9380,N_9379);
nand U9738 (N_9738,N_9462,N_9467);
nand U9739 (N_9739,N_9338,N_9362);
nand U9740 (N_9740,N_9445,N_9420);
xnor U9741 (N_9741,N_9279,N_9346);
or U9742 (N_9742,N_9280,N_9367);
and U9743 (N_9743,N_9369,N_9414);
or U9744 (N_9744,N_9470,N_9375);
or U9745 (N_9745,N_9271,N_9493);
nor U9746 (N_9746,N_9457,N_9291);
and U9747 (N_9747,N_9474,N_9440);
nor U9748 (N_9748,N_9469,N_9394);
nor U9749 (N_9749,N_9422,N_9295);
nor U9750 (N_9750,N_9600,N_9533);
xor U9751 (N_9751,N_9625,N_9611);
or U9752 (N_9752,N_9677,N_9730);
nand U9753 (N_9753,N_9716,N_9728);
or U9754 (N_9754,N_9603,N_9699);
and U9755 (N_9755,N_9586,N_9678);
nand U9756 (N_9756,N_9626,N_9594);
nor U9757 (N_9757,N_9584,N_9717);
nand U9758 (N_9758,N_9577,N_9534);
xor U9759 (N_9759,N_9617,N_9688);
xnor U9760 (N_9760,N_9602,N_9620);
nand U9761 (N_9761,N_9524,N_9519);
nand U9762 (N_9762,N_9543,N_9606);
xor U9763 (N_9763,N_9559,N_9502);
and U9764 (N_9764,N_9647,N_9578);
nor U9765 (N_9765,N_9618,N_9684);
or U9766 (N_9766,N_9651,N_9595);
or U9767 (N_9767,N_9644,N_9707);
or U9768 (N_9768,N_9746,N_9573);
xnor U9769 (N_9769,N_9547,N_9633);
nand U9770 (N_9770,N_9650,N_9562);
or U9771 (N_9771,N_9747,N_9657);
nand U9772 (N_9772,N_9557,N_9561);
or U9773 (N_9773,N_9662,N_9675);
and U9774 (N_9774,N_9663,N_9552);
and U9775 (N_9775,N_9504,N_9530);
or U9776 (N_9776,N_9637,N_9575);
nand U9777 (N_9777,N_9631,N_9668);
and U9778 (N_9778,N_9743,N_9583);
xnor U9779 (N_9779,N_9599,N_9683);
or U9780 (N_9780,N_9567,N_9674);
and U9781 (N_9781,N_9740,N_9541);
nand U9782 (N_9782,N_9540,N_9679);
xor U9783 (N_9783,N_9601,N_9741);
nor U9784 (N_9784,N_9640,N_9658);
nor U9785 (N_9785,N_9642,N_9635);
or U9786 (N_9786,N_9682,N_9616);
nor U9787 (N_9787,N_9520,N_9729);
nor U9788 (N_9788,N_9627,N_9694);
and U9789 (N_9789,N_9597,N_9564);
nor U9790 (N_9790,N_9558,N_9693);
nor U9791 (N_9791,N_9739,N_9697);
and U9792 (N_9792,N_9610,N_9514);
or U9793 (N_9793,N_9588,N_9548);
nor U9794 (N_9794,N_9749,N_9538);
xor U9795 (N_9795,N_9585,N_9571);
nor U9796 (N_9796,N_9560,N_9596);
nand U9797 (N_9797,N_9748,N_9680);
nor U9798 (N_9798,N_9580,N_9581);
nand U9799 (N_9799,N_9632,N_9732);
xor U9800 (N_9800,N_9576,N_9654);
nor U9801 (N_9801,N_9593,N_9612);
xnor U9802 (N_9802,N_9726,N_9526);
xor U9803 (N_9803,N_9572,N_9676);
or U9804 (N_9804,N_9673,N_9702);
nand U9805 (N_9805,N_9645,N_9661);
and U9806 (N_9806,N_9700,N_9745);
nand U9807 (N_9807,N_9665,N_9698);
or U9808 (N_9808,N_9686,N_9568);
nand U9809 (N_9809,N_9629,N_9511);
or U9810 (N_9810,N_9685,N_9725);
or U9811 (N_9811,N_9681,N_9727);
nor U9812 (N_9812,N_9720,N_9609);
nor U9813 (N_9813,N_9744,N_9554);
and U9814 (N_9814,N_9701,N_9638);
xnor U9815 (N_9815,N_9639,N_9653);
xor U9816 (N_9816,N_9721,N_9656);
or U9817 (N_9817,N_9523,N_9643);
nand U9818 (N_9818,N_9710,N_9624);
or U9819 (N_9819,N_9592,N_9501);
and U9820 (N_9820,N_9672,N_9510);
xnor U9821 (N_9821,N_9659,N_9590);
nor U9822 (N_9822,N_9605,N_9536);
nand U9823 (N_9823,N_9566,N_9508);
nor U9824 (N_9824,N_9634,N_9544);
xnor U9825 (N_9825,N_9551,N_9515);
nand U9826 (N_9826,N_9742,N_9733);
xnor U9827 (N_9827,N_9591,N_9655);
nand U9828 (N_9828,N_9549,N_9630);
or U9829 (N_9829,N_9512,N_9509);
nand U9830 (N_9830,N_9722,N_9516);
or U9831 (N_9831,N_9587,N_9545);
nand U9832 (N_9832,N_9715,N_9604);
nand U9833 (N_9833,N_9503,N_9731);
or U9834 (N_9834,N_9667,N_9670);
xnor U9835 (N_9835,N_9703,N_9527);
and U9836 (N_9836,N_9531,N_9705);
nand U9837 (N_9837,N_9718,N_9695);
and U9838 (N_9838,N_9692,N_9507);
or U9839 (N_9839,N_9724,N_9706);
xor U9840 (N_9840,N_9712,N_9619);
xnor U9841 (N_9841,N_9652,N_9529);
xnor U9842 (N_9842,N_9649,N_9579);
xor U9843 (N_9843,N_9521,N_9737);
nor U9844 (N_9844,N_9608,N_9704);
xor U9845 (N_9845,N_9723,N_9734);
or U9846 (N_9846,N_9607,N_9505);
and U9847 (N_9847,N_9528,N_9691);
or U9848 (N_9848,N_9621,N_9539);
xnor U9849 (N_9849,N_9708,N_9613);
or U9850 (N_9850,N_9736,N_9532);
and U9851 (N_9851,N_9711,N_9696);
or U9852 (N_9852,N_9537,N_9628);
nand U9853 (N_9853,N_9666,N_9689);
xor U9854 (N_9854,N_9570,N_9660);
or U9855 (N_9855,N_9555,N_9735);
or U9856 (N_9856,N_9506,N_9589);
xor U9857 (N_9857,N_9669,N_9569);
and U9858 (N_9858,N_9615,N_9500);
and U9859 (N_9859,N_9565,N_9687);
nor U9860 (N_9860,N_9574,N_9614);
and U9861 (N_9861,N_9553,N_9522);
xor U9862 (N_9862,N_9622,N_9671);
and U9863 (N_9863,N_9542,N_9641);
xnor U9864 (N_9864,N_9517,N_9714);
and U9865 (N_9865,N_9623,N_9738);
and U9866 (N_9866,N_9582,N_9664);
xnor U9867 (N_9867,N_9563,N_9709);
xnor U9868 (N_9868,N_9636,N_9518);
nand U9869 (N_9869,N_9646,N_9648);
xnor U9870 (N_9870,N_9550,N_9535);
nand U9871 (N_9871,N_9513,N_9556);
and U9872 (N_9872,N_9690,N_9719);
and U9873 (N_9873,N_9546,N_9713);
nor U9874 (N_9874,N_9525,N_9598);
nor U9875 (N_9875,N_9577,N_9640);
and U9876 (N_9876,N_9697,N_9674);
xor U9877 (N_9877,N_9726,N_9642);
or U9878 (N_9878,N_9588,N_9534);
nand U9879 (N_9879,N_9687,N_9710);
nor U9880 (N_9880,N_9591,N_9529);
nor U9881 (N_9881,N_9560,N_9648);
and U9882 (N_9882,N_9523,N_9516);
and U9883 (N_9883,N_9560,N_9740);
or U9884 (N_9884,N_9689,N_9582);
nand U9885 (N_9885,N_9603,N_9690);
xnor U9886 (N_9886,N_9654,N_9598);
nor U9887 (N_9887,N_9503,N_9514);
nand U9888 (N_9888,N_9737,N_9623);
or U9889 (N_9889,N_9608,N_9639);
or U9890 (N_9890,N_9657,N_9537);
and U9891 (N_9891,N_9648,N_9577);
or U9892 (N_9892,N_9651,N_9619);
nor U9893 (N_9893,N_9604,N_9663);
nor U9894 (N_9894,N_9522,N_9608);
nand U9895 (N_9895,N_9519,N_9533);
and U9896 (N_9896,N_9505,N_9644);
or U9897 (N_9897,N_9647,N_9562);
nor U9898 (N_9898,N_9618,N_9699);
nor U9899 (N_9899,N_9522,N_9582);
and U9900 (N_9900,N_9739,N_9534);
nand U9901 (N_9901,N_9576,N_9706);
nor U9902 (N_9902,N_9704,N_9607);
nand U9903 (N_9903,N_9601,N_9615);
and U9904 (N_9904,N_9594,N_9617);
or U9905 (N_9905,N_9595,N_9690);
and U9906 (N_9906,N_9663,N_9626);
or U9907 (N_9907,N_9603,N_9583);
and U9908 (N_9908,N_9529,N_9561);
xor U9909 (N_9909,N_9690,N_9673);
nor U9910 (N_9910,N_9624,N_9738);
or U9911 (N_9911,N_9719,N_9662);
and U9912 (N_9912,N_9567,N_9692);
and U9913 (N_9913,N_9680,N_9530);
or U9914 (N_9914,N_9672,N_9507);
and U9915 (N_9915,N_9543,N_9519);
xnor U9916 (N_9916,N_9592,N_9546);
nand U9917 (N_9917,N_9537,N_9514);
nor U9918 (N_9918,N_9513,N_9696);
xor U9919 (N_9919,N_9624,N_9509);
nand U9920 (N_9920,N_9540,N_9694);
nor U9921 (N_9921,N_9710,N_9640);
or U9922 (N_9922,N_9575,N_9683);
nand U9923 (N_9923,N_9748,N_9726);
nand U9924 (N_9924,N_9553,N_9727);
nor U9925 (N_9925,N_9690,N_9713);
and U9926 (N_9926,N_9696,N_9560);
xnor U9927 (N_9927,N_9632,N_9628);
xnor U9928 (N_9928,N_9721,N_9598);
nand U9929 (N_9929,N_9713,N_9700);
and U9930 (N_9930,N_9538,N_9699);
nor U9931 (N_9931,N_9636,N_9680);
xnor U9932 (N_9932,N_9541,N_9707);
nor U9933 (N_9933,N_9557,N_9671);
nand U9934 (N_9934,N_9518,N_9574);
nor U9935 (N_9935,N_9675,N_9740);
or U9936 (N_9936,N_9665,N_9745);
or U9937 (N_9937,N_9630,N_9569);
and U9938 (N_9938,N_9708,N_9565);
xnor U9939 (N_9939,N_9515,N_9608);
xor U9940 (N_9940,N_9602,N_9730);
xor U9941 (N_9941,N_9510,N_9625);
nand U9942 (N_9942,N_9609,N_9699);
xor U9943 (N_9943,N_9511,N_9619);
and U9944 (N_9944,N_9624,N_9611);
or U9945 (N_9945,N_9673,N_9534);
nor U9946 (N_9946,N_9742,N_9518);
or U9947 (N_9947,N_9609,N_9639);
nor U9948 (N_9948,N_9633,N_9734);
nor U9949 (N_9949,N_9568,N_9617);
and U9950 (N_9950,N_9643,N_9613);
nand U9951 (N_9951,N_9508,N_9638);
nor U9952 (N_9952,N_9741,N_9553);
xor U9953 (N_9953,N_9641,N_9670);
or U9954 (N_9954,N_9501,N_9523);
and U9955 (N_9955,N_9585,N_9653);
nor U9956 (N_9956,N_9500,N_9503);
or U9957 (N_9957,N_9734,N_9558);
and U9958 (N_9958,N_9608,N_9564);
nor U9959 (N_9959,N_9551,N_9613);
xor U9960 (N_9960,N_9514,N_9654);
or U9961 (N_9961,N_9581,N_9657);
xnor U9962 (N_9962,N_9590,N_9503);
nor U9963 (N_9963,N_9651,N_9679);
and U9964 (N_9964,N_9557,N_9618);
and U9965 (N_9965,N_9561,N_9673);
xnor U9966 (N_9966,N_9656,N_9623);
or U9967 (N_9967,N_9578,N_9718);
nand U9968 (N_9968,N_9702,N_9500);
or U9969 (N_9969,N_9727,N_9623);
xnor U9970 (N_9970,N_9590,N_9699);
and U9971 (N_9971,N_9704,N_9708);
nand U9972 (N_9972,N_9628,N_9588);
and U9973 (N_9973,N_9721,N_9596);
xor U9974 (N_9974,N_9719,N_9738);
nand U9975 (N_9975,N_9724,N_9570);
or U9976 (N_9976,N_9600,N_9608);
nand U9977 (N_9977,N_9723,N_9580);
nand U9978 (N_9978,N_9664,N_9727);
or U9979 (N_9979,N_9600,N_9635);
and U9980 (N_9980,N_9702,N_9661);
xor U9981 (N_9981,N_9736,N_9744);
or U9982 (N_9982,N_9673,N_9584);
nand U9983 (N_9983,N_9541,N_9659);
or U9984 (N_9984,N_9679,N_9583);
or U9985 (N_9985,N_9539,N_9712);
nor U9986 (N_9986,N_9583,N_9706);
xnor U9987 (N_9987,N_9532,N_9606);
or U9988 (N_9988,N_9675,N_9733);
or U9989 (N_9989,N_9693,N_9588);
or U9990 (N_9990,N_9582,N_9683);
nand U9991 (N_9991,N_9626,N_9743);
or U9992 (N_9992,N_9575,N_9590);
or U9993 (N_9993,N_9507,N_9638);
xor U9994 (N_9994,N_9549,N_9687);
and U9995 (N_9995,N_9517,N_9585);
nand U9996 (N_9996,N_9661,N_9641);
or U9997 (N_9997,N_9697,N_9546);
nor U9998 (N_9998,N_9618,N_9616);
nor U9999 (N_9999,N_9580,N_9716);
nor U10000 (N_10000,N_9975,N_9799);
xor U10001 (N_10001,N_9938,N_9961);
and U10002 (N_10002,N_9841,N_9875);
nor U10003 (N_10003,N_9974,N_9944);
or U10004 (N_10004,N_9930,N_9942);
nor U10005 (N_10005,N_9805,N_9919);
or U10006 (N_10006,N_9801,N_9834);
nand U10007 (N_10007,N_9885,N_9889);
nor U10008 (N_10008,N_9920,N_9782);
or U10009 (N_10009,N_9852,N_9802);
nor U10010 (N_10010,N_9814,N_9902);
xor U10011 (N_10011,N_9916,N_9973);
nand U10012 (N_10012,N_9810,N_9999);
nor U10013 (N_10013,N_9987,N_9827);
nor U10014 (N_10014,N_9767,N_9878);
and U10015 (N_10015,N_9756,N_9934);
xnor U10016 (N_10016,N_9797,N_9849);
nand U10017 (N_10017,N_9762,N_9850);
and U10018 (N_10018,N_9845,N_9868);
nor U10019 (N_10019,N_9857,N_9812);
nand U10020 (N_10020,N_9867,N_9753);
xnor U10021 (N_10021,N_9925,N_9958);
and U10022 (N_10022,N_9828,N_9754);
and U10023 (N_10023,N_9906,N_9811);
nand U10024 (N_10024,N_9790,N_9766);
xor U10025 (N_10025,N_9793,N_9819);
and U10026 (N_10026,N_9905,N_9968);
and U10027 (N_10027,N_9864,N_9768);
nand U10028 (N_10028,N_9788,N_9763);
xnor U10029 (N_10029,N_9877,N_9806);
or U10030 (N_10030,N_9879,N_9794);
nand U10031 (N_10031,N_9836,N_9899);
and U10032 (N_10032,N_9777,N_9912);
and U10033 (N_10033,N_9853,N_9984);
xnor U10034 (N_10034,N_9903,N_9921);
xnor U10035 (N_10035,N_9796,N_9838);
nor U10036 (N_10036,N_9952,N_9821);
xor U10037 (N_10037,N_9943,N_9817);
nor U10038 (N_10038,N_9994,N_9893);
nand U10039 (N_10039,N_9967,N_9989);
and U10040 (N_10040,N_9783,N_9960);
xnor U10041 (N_10041,N_9829,N_9991);
and U10042 (N_10042,N_9996,N_9846);
nand U10043 (N_10043,N_9964,N_9923);
or U10044 (N_10044,N_9939,N_9954);
nand U10045 (N_10045,N_9992,N_9972);
and U10046 (N_10046,N_9894,N_9804);
and U10047 (N_10047,N_9800,N_9949);
or U10048 (N_10048,N_9976,N_9755);
or U10049 (N_10049,N_9966,N_9824);
xor U10050 (N_10050,N_9781,N_9775);
nor U10051 (N_10051,N_9859,N_9924);
and U10052 (N_10052,N_9854,N_9888);
nor U10053 (N_10053,N_9915,N_9891);
or U10054 (N_10054,N_9953,N_9890);
xor U10055 (N_10055,N_9978,N_9844);
nor U10056 (N_10056,N_9896,N_9917);
and U10057 (N_10057,N_9951,N_9780);
nand U10058 (N_10058,N_9981,N_9870);
and U10059 (N_10059,N_9956,N_9881);
and U10060 (N_10060,N_9757,N_9932);
and U10061 (N_10061,N_9820,N_9998);
nor U10062 (N_10062,N_9760,N_9892);
and U10063 (N_10063,N_9803,N_9988);
nand U10064 (N_10064,N_9933,N_9818);
and U10065 (N_10065,N_9936,N_9770);
nand U10066 (N_10066,N_9959,N_9927);
xor U10067 (N_10067,N_9970,N_9761);
nor U10068 (N_10068,N_9928,N_9895);
or U10069 (N_10069,N_9937,N_9779);
nor U10070 (N_10070,N_9901,N_9839);
or U10071 (N_10071,N_9861,N_9985);
xor U10072 (N_10072,N_9983,N_9813);
nand U10073 (N_10073,N_9913,N_9969);
xnor U10074 (N_10074,N_9977,N_9869);
or U10075 (N_10075,N_9830,N_9882);
or U10076 (N_10076,N_9764,N_9995);
nor U10077 (N_10077,N_9855,N_9833);
and U10078 (N_10078,N_9826,N_9858);
xor U10079 (N_10079,N_9909,N_9871);
nand U10080 (N_10080,N_9897,N_9886);
and U10081 (N_10081,N_9789,N_9947);
or U10082 (N_10082,N_9898,N_9798);
or U10083 (N_10083,N_9786,N_9950);
and U10084 (N_10084,N_9856,N_9872);
nor U10085 (N_10085,N_9776,N_9940);
nand U10086 (N_10086,N_9843,N_9908);
and U10087 (N_10087,N_9945,N_9965);
xor U10088 (N_10088,N_9948,N_9980);
or U10089 (N_10089,N_9807,N_9941);
xor U10090 (N_10090,N_9946,N_9955);
or U10091 (N_10091,N_9785,N_9840);
nand U10092 (N_10092,N_9935,N_9929);
or U10093 (N_10093,N_9904,N_9831);
or U10094 (N_10094,N_9884,N_9758);
and U10095 (N_10095,N_9832,N_9808);
nor U10096 (N_10096,N_9860,N_9863);
nand U10097 (N_10097,N_9848,N_9751);
nor U10098 (N_10098,N_9752,N_9862);
and U10099 (N_10099,N_9979,N_9769);
or U10100 (N_10100,N_9911,N_9792);
nand U10101 (N_10101,N_9880,N_9865);
nor U10102 (N_10102,N_9922,N_9866);
or U10103 (N_10103,N_9963,N_9993);
nand U10104 (N_10104,N_9765,N_9962);
or U10105 (N_10105,N_9784,N_9822);
and U10106 (N_10106,N_9750,N_9900);
or U10107 (N_10107,N_9971,N_9982);
nand U10108 (N_10108,N_9787,N_9825);
nor U10109 (N_10109,N_9997,N_9774);
xnor U10110 (N_10110,N_9778,N_9918);
or U10111 (N_10111,N_9809,N_9847);
nor U10112 (N_10112,N_9772,N_9986);
and U10113 (N_10113,N_9837,N_9823);
nor U10114 (N_10114,N_9883,N_9759);
nor U10115 (N_10115,N_9771,N_9815);
xor U10116 (N_10116,N_9931,N_9887);
nand U10117 (N_10117,N_9876,N_9795);
or U10118 (N_10118,N_9835,N_9874);
and U10119 (N_10119,N_9791,N_9851);
or U10120 (N_10120,N_9842,N_9926);
nand U10121 (N_10121,N_9907,N_9873);
and U10122 (N_10122,N_9990,N_9816);
or U10123 (N_10123,N_9914,N_9773);
nor U10124 (N_10124,N_9910,N_9957);
xnor U10125 (N_10125,N_9983,N_9881);
nor U10126 (N_10126,N_9901,N_9829);
and U10127 (N_10127,N_9916,N_9869);
or U10128 (N_10128,N_9845,N_9878);
nor U10129 (N_10129,N_9795,N_9836);
and U10130 (N_10130,N_9916,N_9992);
xor U10131 (N_10131,N_9775,N_9798);
or U10132 (N_10132,N_9984,N_9772);
xor U10133 (N_10133,N_9826,N_9935);
nor U10134 (N_10134,N_9804,N_9888);
or U10135 (N_10135,N_9899,N_9751);
xnor U10136 (N_10136,N_9777,N_9961);
and U10137 (N_10137,N_9903,N_9861);
nand U10138 (N_10138,N_9932,N_9853);
and U10139 (N_10139,N_9919,N_9895);
nand U10140 (N_10140,N_9935,N_9836);
or U10141 (N_10141,N_9913,N_9758);
xor U10142 (N_10142,N_9846,N_9963);
xor U10143 (N_10143,N_9825,N_9762);
xor U10144 (N_10144,N_9872,N_9824);
nor U10145 (N_10145,N_9773,N_9871);
nor U10146 (N_10146,N_9941,N_9822);
and U10147 (N_10147,N_9791,N_9963);
xnor U10148 (N_10148,N_9798,N_9808);
nor U10149 (N_10149,N_9812,N_9829);
xor U10150 (N_10150,N_9877,N_9934);
or U10151 (N_10151,N_9759,N_9999);
nor U10152 (N_10152,N_9766,N_9813);
xnor U10153 (N_10153,N_9834,N_9998);
nor U10154 (N_10154,N_9903,N_9817);
xnor U10155 (N_10155,N_9894,N_9936);
xor U10156 (N_10156,N_9878,N_9858);
xnor U10157 (N_10157,N_9936,N_9853);
nor U10158 (N_10158,N_9845,N_9961);
nor U10159 (N_10159,N_9865,N_9882);
or U10160 (N_10160,N_9873,N_9946);
nand U10161 (N_10161,N_9909,N_9861);
xnor U10162 (N_10162,N_9996,N_9872);
xnor U10163 (N_10163,N_9753,N_9871);
nor U10164 (N_10164,N_9770,N_9785);
nor U10165 (N_10165,N_9923,N_9861);
nor U10166 (N_10166,N_9878,N_9881);
xnor U10167 (N_10167,N_9837,N_9954);
nand U10168 (N_10168,N_9964,N_9823);
and U10169 (N_10169,N_9774,N_9924);
nand U10170 (N_10170,N_9786,N_9932);
nor U10171 (N_10171,N_9976,N_9920);
xnor U10172 (N_10172,N_9762,N_9827);
or U10173 (N_10173,N_9809,N_9941);
xnor U10174 (N_10174,N_9886,N_9758);
nand U10175 (N_10175,N_9878,N_9980);
nand U10176 (N_10176,N_9820,N_9890);
or U10177 (N_10177,N_9949,N_9874);
xnor U10178 (N_10178,N_9951,N_9819);
and U10179 (N_10179,N_9876,N_9830);
and U10180 (N_10180,N_9777,N_9874);
and U10181 (N_10181,N_9798,N_9960);
nand U10182 (N_10182,N_9756,N_9992);
xor U10183 (N_10183,N_9868,N_9750);
and U10184 (N_10184,N_9987,N_9941);
nand U10185 (N_10185,N_9882,N_9808);
nand U10186 (N_10186,N_9864,N_9790);
nand U10187 (N_10187,N_9866,N_9963);
nor U10188 (N_10188,N_9972,N_9750);
nor U10189 (N_10189,N_9770,N_9792);
and U10190 (N_10190,N_9996,N_9966);
or U10191 (N_10191,N_9786,N_9839);
and U10192 (N_10192,N_9889,N_9989);
or U10193 (N_10193,N_9864,N_9828);
xor U10194 (N_10194,N_9973,N_9821);
and U10195 (N_10195,N_9791,N_9883);
nor U10196 (N_10196,N_9972,N_9878);
and U10197 (N_10197,N_9897,N_9955);
xnor U10198 (N_10198,N_9819,N_9776);
nand U10199 (N_10199,N_9880,N_9962);
and U10200 (N_10200,N_9768,N_9957);
or U10201 (N_10201,N_9967,N_9984);
xor U10202 (N_10202,N_9808,N_9973);
nor U10203 (N_10203,N_9872,N_9932);
nor U10204 (N_10204,N_9905,N_9886);
and U10205 (N_10205,N_9750,N_9962);
nor U10206 (N_10206,N_9764,N_9872);
xnor U10207 (N_10207,N_9784,N_9858);
nor U10208 (N_10208,N_9892,N_9903);
and U10209 (N_10209,N_9755,N_9882);
or U10210 (N_10210,N_9760,N_9849);
xor U10211 (N_10211,N_9852,N_9810);
nand U10212 (N_10212,N_9948,N_9876);
nand U10213 (N_10213,N_9896,N_9864);
or U10214 (N_10214,N_9828,N_9856);
nand U10215 (N_10215,N_9771,N_9817);
xor U10216 (N_10216,N_9799,N_9879);
and U10217 (N_10217,N_9895,N_9923);
nand U10218 (N_10218,N_9994,N_9832);
or U10219 (N_10219,N_9802,N_9888);
xor U10220 (N_10220,N_9797,N_9858);
or U10221 (N_10221,N_9938,N_9903);
nor U10222 (N_10222,N_9914,N_9792);
or U10223 (N_10223,N_9801,N_9776);
or U10224 (N_10224,N_9795,N_9993);
nor U10225 (N_10225,N_9755,N_9993);
nand U10226 (N_10226,N_9971,N_9831);
nand U10227 (N_10227,N_9850,N_9957);
or U10228 (N_10228,N_9873,N_9903);
and U10229 (N_10229,N_9949,N_9917);
nor U10230 (N_10230,N_9971,N_9943);
nor U10231 (N_10231,N_9928,N_9939);
nor U10232 (N_10232,N_9875,N_9899);
nor U10233 (N_10233,N_9996,N_9949);
and U10234 (N_10234,N_9909,N_9915);
nand U10235 (N_10235,N_9825,N_9875);
and U10236 (N_10236,N_9964,N_9999);
and U10237 (N_10237,N_9942,N_9803);
nand U10238 (N_10238,N_9778,N_9936);
and U10239 (N_10239,N_9795,N_9999);
or U10240 (N_10240,N_9885,N_9908);
or U10241 (N_10241,N_9946,N_9898);
nor U10242 (N_10242,N_9923,N_9995);
nand U10243 (N_10243,N_9763,N_9880);
or U10244 (N_10244,N_9923,N_9829);
nand U10245 (N_10245,N_9853,N_9776);
or U10246 (N_10246,N_9764,N_9956);
nor U10247 (N_10247,N_9758,N_9833);
nor U10248 (N_10248,N_9993,N_9990);
nand U10249 (N_10249,N_9764,N_9757);
and U10250 (N_10250,N_10230,N_10111);
xnor U10251 (N_10251,N_10050,N_10033);
xor U10252 (N_10252,N_10051,N_10044);
nand U10253 (N_10253,N_10196,N_10185);
or U10254 (N_10254,N_10120,N_10208);
xor U10255 (N_10255,N_10153,N_10147);
or U10256 (N_10256,N_10123,N_10133);
nand U10257 (N_10257,N_10092,N_10002);
or U10258 (N_10258,N_10020,N_10014);
or U10259 (N_10259,N_10069,N_10118);
nor U10260 (N_10260,N_10030,N_10248);
or U10261 (N_10261,N_10209,N_10138);
nand U10262 (N_10262,N_10204,N_10059);
nand U10263 (N_10263,N_10135,N_10056);
nand U10264 (N_10264,N_10088,N_10075);
and U10265 (N_10265,N_10239,N_10145);
and U10266 (N_10266,N_10124,N_10184);
nand U10267 (N_10267,N_10049,N_10099);
nand U10268 (N_10268,N_10001,N_10043);
nand U10269 (N_10269,N_10160,N_10005);
nand U10270 (N_10270,N_10172,N_10127);
nor U10271 (N_10271,N_10095,N_10202);
or U10272 (N_10272,N_10187,N_10188);
nand U10273 (N_10273,N_10213,N_10175);
or U10274 (N_10274,N_10164,N_10074);
and U10275 (N_10275,N_10183,N_10119);
xnor U10276 (N_10276,N_10212,N_10057);
nand U10277 (N_10277,N_10094,N_10086);
nor U10278 (N_10278,N_10042,N_10149);
nor U10279 (N_10279,N_10129,N_10136);
or U10280 (N_10280,N_10079,N_10078);
nor U10281 (N_10281,N_10067,N_10190);
xnor U10282 (N_10282,N_10226,N_10235);
nand U10283 (N_10283,N_10199,N_10217);
and U10284 (N_10284,N_10016,N_10017);
xor U10285 (N_10285,N_10089,N_10162);
nand U10286 (N_10286,N_10060,N_10132);
nor U10287 (N_10287,N_10211,N_10058);
xor U10288 (N_10288,N_10003,N_10077);
and U10289 (N_10289,N_10180,N_10008);
nand U10290 (N_10290,N_10143,N_10206);
nor U10291 (N_10291,N_10018,N_10122);
nor U10292 (N_10292,N_10223,N_10219);
nand U10293 (N_10293,N_10152,N_10216);
or U10294 (N_10294,N_10197,N_10195);
and U10295 (N_10295,N_10110,N_10103);
nor U10296 (N_10296,N_10177,N_10080);
and U10297 (N_10297,N_10072,N_10054);
nand U10298 (N_10298,N_10065,N_10245);
or U10299 (N_10299,N_10171,N_10186);
xor U10300 (N_10300,N_10224,N_10198);
nor U10301 (N_10301,N_10243,N_10036);
xnor U10302 (N_10302,N_10159,N_10125);
or U10303 (N_10303,N_10109,N_10131);
nor U10304 (N_10304,N_10112,N_10169);
xor U10305 (N_10305,N_10105,N_10144);
and U10306 (N_10306,N_10038,N_10128);
xnor U10307 (N_10307,N_10182,N_10146);
xnor U10308 (N_10308,N_10007,N_10221);
or U10309 (N_10309,N_10222,N_10022);
nand U10310 (N_10310,N_10139,N_10247);
nand U10311 (N_10311,N_10170,N_10200);
or U10312 (N_10312,N_10238,N_10240);
nor U10313 (N_10313,N_10141,N_10249);
nand U10314 (N_10314,N_10142,N_10040);
or U10315 (N_10315,N_10168,N_10228);
xor U10316 (N_10316,N_10047,N_10066);
xor U10317 (N_10317,N_10004,N_10039);
nand U10318 (N_10318,N_10013,N_10166);
or U10319 (N_10319,N_10009,N_10082);
xor U10320 (N_10320,N_10207,N_10097);
xnor U10321 (N_10321,N_10041,N_10052);
nor U10322 (N_10322,N_10130,N_10062);
xor U10323 (N_10323,N_10148,N_10178);
nand U10324 (N_10324,N_10117,N_10242);
and U10325 (N_10325,N_10012,N_10090);
xor U10326 (N_10326,N_10241,N_10157);
or U10327 (N_10327,N_10192,N_10023);
or U10328 (N_10328,N_10061,N_10179);
and U10329 (N_10329,N_10068,N_10244);
nand U10330 (N_10330,N_10234,N_10091);
or U10331 (N_10331,N_10071,N_10011);
nand U10332 (N_10332,N_10140,N_10096);
xor U10333 (N_10333,N_10076,N_10167);
nor U10334 (N_10334,N_10031,N_10246);
nor U10335 (N_10335,N_10215,N_10165);
and U10336 (N_10336,N_10102,N_10218);
xor U10337 (N_10337,N_10137,N_10121);
nor U10338 (N_10338,N_10113,N_10045);
nor U10339 (N_10339,N_10024,N_10227);
nand U10340 (N_10340,N_10154,N_10114);
nor U10341 (N_10341,N_10237,N_10010);
xnor U10342 (N_10342,N_10176,N_10034);
nand U10343 (N_10343,N_10116,N_10070);
and U10344 (N_10344,N_10189,N_10063);
and U10345 (N_10345,N_10150,N_10236);
and U10346 (N_10346,N_10087,N_10028);
xnor U10347 (N_10347,N_10193,N_10232);
xnor U10348 (N_10348,N_10084,N_10104);
nor U10349 (N_10349,N_10134,N_10201);
or U10350 (N_10350,N_10181,N_10015);
nor U10351 (N_10351,N_10194,N_10098);
or U10352 (N_10352,N_10225,N_10115);
nor U10353 (N_10353,N_10026,N_10053);
nor U10354 (N_10354,N_10083,N_10233);
nand U10355 (N_10355,N_10229,N_10163);
xor U10356 (N_10356,N_10100,N_10027);
and U10357 (N_10357,N_10126,N_10073);
xor U10358 (N_10358,N_10029,N_10032);
or U10359 (N_10359,N_10220,N_10156);
nand U10360 (N_10360,N_10006,N_10107);
nor U10361 (N_10361,N_10158,N_10093);
or U10362 (N_10362,N_10037,N_10048);
nand U10363 (N_10363,N_10191,N_10025);
or U10364 (N_10364,N_10231,N_10108);
nand U10365 (N_10365,N_10085,N_10021);
nor U10366 (N_10366,N_10173,N_10046);
nor U10367 (N_10367,N_10210,N_10106);
and U10368 (N_10368,N_10000,N_10035);
nand U10369 (N_10369,N_10155,N_10055);
xnor U10370 (N_10370,N_10064,N_10214);
nor U10371 (N_10371,N_10203,N_10161);
nand U10372 (N_10372,N_10205,N_10151);
or U10373 (N_10373,N_10174,N_10101);
and U10374 (N_10374,N_10019,N_10081);
nor U10375 (N_10375,N_10023,N_10168);
xnor U10376 (N_10376,N_10177,N_10184);
or U10377 (N_10377,N_10146,N_10142);
or U10378 (N_10378,N_10153,N_10037);
xor U10379 (N_10379,N_10125,N_10247);
nor U10380 (N_10380,N_10043,N_10223);
xnor U10381 (N_10381,N_10172,N_10235);
or U10382 (N_10382,N_10199,N_10122);
and U10383 (N_10383,N_10085,N_10084);
nor U10384 (N_10384,N_10143,N_10168);
xor U10385 (N_10385,N_10207,N_10028);
and U10386 (N_10386,N_10025,N_10071);
nor U10387 (N_10387,N_10061,N_10176);
and U10388 (N_10388,N_10165,N_10009);
nand U10389 (N_10389,N_10181,N_10190);
and U10390 (N_10390,N_10045,N_10092);
nor U10391 (N_10391,N_10220,N_10193);
nand U10392 (N_10392,N_10160,N_10051);
nand U10393 (N_10393,N_10148,N_10187);
xor U10394 (N_10394,N_10020,N_10174);
nor U10395 (N_10395,N_10136,N_10081);
and U10396 (N_10396,N_10058,N_10065);
and U10397 (N_10397,N_10051,N_10125);
and U10398 (N_10398,N_10124,N_10133);
nor U10399 (N_10399,N_10076,N_10103);
or U10400 (N_10400,N_10061,N_10034);
xnor U10401 (N_10401,N_10042,N_10089);
nor U10402 (N_10402,N_10177,N_10233);
or U10403 (N_10403,N_10001,N_10170);
and U10404 (N_10404,N_10128,N_10244);
xor U10405 (N_10405,N_10045,N_10231);
nand U10406 (N_10406,N_10243,N_10227);
xor U10407 (N_10407,N_10223,N_10107);
and U10408 (N_10408,N_10219,N_10084);
or U10409 (N_10409,N_10030,N_10097);
and U10410 (N_10410,N_10241,N_10100);
or U10411 (N_10411,N_10209,N_10118);
or U10412 (N_10412,N_10023,N_10105);
or U10413 (N_10413,N_10032,N_10100);
xor U10414 (N_10414,N_10028,N_10029);
nand U10415 (N_10415,N_10239,N_10226);
nor U10416 (N_10416,N_10156,N_10169);
xnor U10417 (N_10417,N_10224,N_10107);
and U10418 (N_10418,N_10025,N_10034);
or U10419 (N_10419,N_10023,N_10094);
xnor U10420 (N_10420,N_10226,N_10067);
and U10421 (N_10421,N_10000,N_10079);
or U10422 (N_10422,N_10244,N_10010);
nor U10423 (N_10423,N_10050,N_10205);
or U10424 (N_10424,N_10214,N_10233);
and U10425 (N_10425,N_10081,N_10113);
or U10426 (N_10426,N_10189,N_10096);
nor U10427 (N_10427,N_10198,N_10003);
nand U10428 (N_10428,N_10066,N_10051);
xor U10429 (N_10429,N_10232,N_10189);
or U10430 (N_10430,N_10248,N_10059);
or U10431 (N_10431,N_10172,N_10205);
and U10432 (N_10432,N_10026,N_10166);
xnor U10433 (N_10433,N_10127,N_10226);
nand U10434 (N_10434,N_10086,N_10218);
nor U10435 (N_10435,N_10231,N_10090);
nor U10436 (N_10436,N_10154,N_10151);
and U10437 (N_10437,N_10054,N_10045);
nor U10438 (N_10438,N_10078,N_10095);
and U10439 (N_10439,N_10149,N_10162);
and U10440 (N_10440,N_10107,N_10195);
xnor U10441 (N_10441,N_10181,N_10066);
xnor U10442 (N_10442,N_10086,N_10024);
and U10443 (N_10443,N_10070,N_10158);
nor U10444 (N_10444,N_10209,N_10045);
xnor U10445 (N_10445,N_10208,N_10058);
nor U10446 (N_10446,N_10010,N_10026);
and U10447 (N_10447,N_10206,N_10118);
nor U10448 (N_10448,N_10161,N_10036);
nor U10449 (N_10449,N_10075,N_10027);
or U10450 (N_10450,N_10019,N_10051);
xnor U10451 (N_10451,N_10178,N_10124);
nand U10452 (N_10452,N_10119,N_10153);
or U10453 (N_10453,N_10073,N_10179);
and U10454 (N_10454,N_10012,N_10154);
and U10455 (N_10455,N_10109,N_10163);
nor U10456 (N_10456,N_10168,N_10086);
and U10457 (N_10457,N_10053,N_10219);
nor U10458 (N_10458,N_10093,N_10134);
nand U10459 (N_10459,N_10162,N_10083);
nand U10460 (N_10460,N_10205,N_10044);
nor U10461 (N_10461,N_10012,N_10196);
nand U10462 (N_10462,N_10014,N_10034);
and U10463 (N_10463,N_10193,N_10120);
nand U10464 (N_10464,N_10096,N_10172);
and U10465 (N_10465,N_10108,N_10111);
nand U10466 (N_10466,N_10045,N_10121);
nand U10467 (N_10467,N_10227,N_10064);
or U10468 (N_10468,N_10017,N_10159);
xnor U10469 (N_10469,N_10096,N_10000);
nor U10470 (N_10470,N_10179,N_10199);
or U10471 (N_10471,N_10022,N_10033);
and U10472 (N_10472,N_10008,N_10232);
nor U10473 (N_10473,N_10075,N_10041);
nand U10474 (N_10474,N_10067,N_10154);
xnor U10475 (N_10475,N_10083,N_10243);
or U10476 (N_10476,N_10215,N_10042);
nor U10477 (N_10477,N_10145,N_10017);
xnor U10478 (N_10478,N_10120,N_10020);
nand U10479 (N_10479,N_10016,N_10091);
and U10480 (N_10480,N_10226,N_10084);
nand U10481 (N_10481,N_10038,N_10054);
xnor U10482 (N_10482,N_10019,N_10147);
nand U10483 (N_10483,N_10069,N_10212);
xor U10484 (N_10484,N_10027,N_10076);
nor U10485 (N_10485,N_10032,N_10026);
nand U10486 (N_10486,N_10118,N_10216);
nor U10487 (N_10487,N_10016,N_10243);
nor U10488 (N_10488,N_10083,N_10108);
xor U10489 (N_10489,N_10132,N_10211);
or U10490 (N_10490,N_10008,N_10052);
xnor U10491 (N_10491,N_10051,N_10136);
or U10492 (N_10492,N_10102,N_10060);
or U10493 (N_10493,N_10139,N_10008);
nand U10494 (N_10494,N_10215,N_10074);
xnor U10495 (N_10495,N_10202,N_10101);
and U10496 (N_10496,N_10157,N_10044);
xor U10497 (N_10497,N_10009,N_10196);
nand U10498 (N_10498,N_10100,N_10095);
nor U10499 (N_10499,N_10238,N_10119);
nor U10500 (N_10500,N_10315,N_10418);
nand U10501 (N_10501,N_10329,N_10391);
xor U10502 (N_10502,N_10368,N_10478);
xnor U10503 (N_10503,N_10288,N_10486);
or U10504 (N_10504,N_10392,N_10449);
nor U10505 (N_10505,N_10408,N_10476);
xnor U10506 (N_10506,N_10432,N_10356);
or U10507 (N_10507,N_10345,N_10436);
or U10508 (N_10508,N_10459,N_10370);
nor U10509 (N_10509,N_10265,N_10362);
nand U10510 (N_10510,N_10493,N_10332);
and U10511 (N_10511,N_10429,N_10499);
xnor U10512 (N_10512,N_10498,N_10317);
and U10513 (N_10513,N_10266,N_10427);
or U10514 (N_10514,N_10341,N_10277);
or U10515 (N_10515,N_10294,N_10325);
or U10516 (N_10516,N_10286,N_10346);
nand U10517 (N_10517,N_10250,N_10333);
or U10518 (N_10518,N_10335,N_10412);
or U10519 (N_10519,N_10393,N_10423);
or U10520 (N_10520,N_10416,N_10401);
xor U10521 (N_10521,N_10428,N_10483);
and U10522 (N_10522,N_10275,N_10377);
nor U10523 (N_10523,N_10293,N_10276);
nor U10524 (N_10524,N_10470,N_10330);
nand U10525 (N_10525,N_10420,N_10338);
nor U10526 (N_10526,N_10361,N_10384);
xnor U10527 (N_10527,N_10474,N_10425);
and U10528 (N_10528,N_10475,N_10487);
and U10529 (N_10529,N_10347,N_10430);
and U10530 (N_10530,N_10343,N_10355);
nor U10531 (N_10531,N_10394,N_10446);
and U10532 (N_10532,N_10326,N_10410);
xor U10533 (N_10533,N_10278,N_10259);
and U10534 (N_10534,N_10385,N_10299);
and U10535 (N_10535,N_10448,N_10337);
or U10536 (N_10536,N_10441,N_10365);
xnor U10537 (N_10537,N_10484,N_10285);
and U10538 (N_10538,N_10477,N_10389);
nand U10539 (N_10539,N_10331,N_10291);
xnor U10540 (N_10540,N_10379,N_10296);
nand U10541 (N_10541,N_10352,N_10454);
nor U10542 (N_10542,N_10434,N_10464);
and U10543 (N_10543,N_10468,N_10471);
or U10544 (N_10544,N_10473,N_10450);
and U10545 (N_10545,N_10466,N_10262);
nand U10546 (N_10546,N_10463,N_10460);
nand U10547 (N_10547,N_10282,N_10403);
nor U10548 (N_10548,N_10458,N_10271);
nor U10549 (N_10549,N_10342,N_10426);
nor U10550 (N_10550,N_10386,N_10437);
and U10551 (N_10551,N_10388,N_10268);
xnor U10552 (N_10552,N_10407,N_10311);
and U10553 (N_10553,N_10455,N_10322);
xnor U10554 (N_10554,N_10283,N_10297);
nand U10555 (N_10555,N_10435,N_10415);
nor U10556 (N_10556,N_10324,N_10480);
and U10557 (N_10557,N_10387,N_10414);
xnor U10558 (N_10558,N_10479,N_10372);
xnor U10559 (N_10559,N_10264,N_10327);
and U10560 (N_10560,N_10358,N_10287);
nor U10561 (N_10561,N_10371,N_10316);
nand U10562 (N_10562,N_10251,N_10263);
and U10563 (N_10563,N_10279,N_10318);
nand U10564 (N_10564,N_10398,N_10395);
and U10565 (N_10565,N_10462,N_10301);
nand U10566 (N_10566,N_10252,N_10363);
nand U10567 (N_10567,N_10310,N_10349);
and U10568 (N_10568,N_10472,N_10453);
xnor U10569 (N_10569,N_10490,N_10273);
or U10570 (N_10570,N_10314,N_10456);
nor U10571 (N_10571,N_10360,N_10492);
nand U10572 (N_10572,N_10469,N_10439);
xor U10573 (N_10573,N_10397,N_10376);
nand U10574 (N_10574,N_10298,N_10440);
nor U10575 (N_10575,N_10381,N_10400);
xor U10576 (N_10576,N_10421,N_10438);
or U10577 (N_10577,N_10290,N_10417);
nor U10578 (N_10578,N_10442,N_10411);
xnor U10579 (N_10579,N_10405,N_10399);
and U10580 (N_10580,N_10339,N_10481);
or U10581 (N_10581,N_10323,N_10353);
nor U10582 (N_10582,N_10382,N_10305);
and U10583 (N_10583,N_10366,N_10419);
and U10584 (N_10584,N_10380,N_10289);
and U10585 (N_10585,N_10467,N_10304);
and U10586 (N_10586,N_10452,N_10485);
nor U10587 (N_10587,N_10320,N_10375);
nand U10588 (N_10588,N_10257,N_10261);
xor U10589 (N_10589,N_10433,N_10396);
nand U10590 (N_10590,N_10284,N_10351);
and U10591 (N_10591,N_10367,N_10280);
and U10592 (N_10592,N_10302,N_10445);
and U10593 (N_10593,N_10359,N_10390);
nand U10594 (N_10594,N_10336,N_10269);
nor U10595 (N_10595,N_10409,N_10319);
nand U10596 (N_10596,N_10413,N_10496);
nand U10597 (N_10597,N_10422,N_10424);
nand U10598 (N_10598,N_10321,N_10369);
and U10599 (N_10599,N_10334,N_10497);
nand U10600 (N_10600,N_10383,N_10451);
nor U10601 (N_10601,N_10313,N_10488);
xnor U10602 (N_10602,N_10443,N_10274);
and U10603 (N_10603,N_10309,N_10364);
or U10604 (N_10604,N_10495,N_10489);
xor U10605 (N_10605,N_10373,N_10431);
and U10606 (N_10606,N_10260,N_10465);
nand U10607 (N_10607,N_10402,N_10300);
and U10608 (N_10608,N_10295,N_10374);
or U10609 (N_10609,N_10491,N_10357);
xor U10610 (N_10610,N_10406,N_10328);
nor U10611 (N_10611,N_10258,N_10281);
nor U10612 (N_10612,N_10303,N_10267);
nor U10613 (N_10613,N_10308,N_10457);
nand U10614 (N_10614,N_10354,N_10344);
nor U10615 (N_10615,N_10270,N_10378);
nand U10616 (N_10616,N_10350,N_10348);
xnor U10617 (N_10617,N_10272,N_10447);
nand U10618 (N_10618,N_10253,N_10494);
and U10619 (N_10619,N_10292,N_10307);
xnor U10620 (N_10620,N_10256,N_10461);
and U10621 (N_10621,N_10255,N_10444);
and U10622 (N_10622,N_10254,N_10482);
xnor U10623 (N_10623,N_10404,N_10340);
nor U10624 (N_10624,N_10306,N_10312);
or U10625 (N_10625,N_10286,N_10365);
and U10626 (N_10626,N_10451,N_10454);
and U10627 (N_10627,N_10359,N_10415);
nor U10628 (N_10628,N_10421,N_10369);
xnor U10629 (N_10629,N_10350,N_10316);
nor U10630 (N_10630,N_10329,N_10355);
xor U10631 (N_10631,N_10388,N_10497);
and U10632 (N_10632,N_10305,N_10332);
or U10633 (N_10633,N_10351,N_10253);
or U10634 (N_10634,N_10329,N_10447);
xor U10635 (N_10635,N_10401,N_10288);
or U10636 (N_10636,N_10454,N_10339);
nor U10637 (N_10637,N_10443,N_10411);
or U10638 (N_10638,N_10442,N_10401);
xor U10639 (N_10639,N_10283,N_10457);
nand U10640 (N_10640,N_10487,N_10428);
nand U10641 (N_10641,N_10322,N_10368);
xor U10642 (N_10642,N_10405,N_10348);
xnor U10643 (N_10643,N_10462,N_10312);
and U10644 (N_10644,N_10260,N_10286);
nor U10645 (N_10645,N_10499,N_10350);
nand U10646 (N_10646,N_10456,N_10454);
and U10647 (N_10647,N_10494,N_10307);
nand U10648 (N_10648,N_10498,N_10264);
xor U10649 (N_10649,N_10332,N_10460);
and U10650 (N_10650,N_10405,N_10420);
or U10651 (N_10651,N_10489,N_10290);
xor U10652 (N_10652,N_10300,N_10369);
nand U10653 (N_10653,N_10320,N_10287);
and U10654 (N_10654,N_10407,N_10269);
nor U10655 (N_10655,N_10390,N_10354);
xor U10656 (N_10656,N_10352,N_10322);
xor U10657 (N_10657,N_10310,N_10363);
nor U10658 (N_10658,N_10298,N_10361);
nand U10659 (N_10659,N_10498,N_10258);
or U10660 (N_10660,N_10406,N_10334);
nor U10661 (N_10661,N_10403,N_10471);
nor U10662 (N_10662,N_10329,N_10424);
or U10663 (N_10663,N_10498,N_10466);
and U10664 (N_10664,N_10372,N_10394);
nand U10665 (N_10665,N_10291,N_10452);
and U10666 (N_10666,N_10415,N_10257);
and U10667 (N_10667,N_10378,N_10386);
nand U10668 (N_10668,N_10364,N_10275);
nor U10669 (N_10669,N_10309,N_10347);
xor U10670 (N_10670,N_10351,N_10391);
nand U10671 (N_10671,N_10297,N_10315);
nand U10672 (N_10672,N_10316,N_10458);
nor U10673 (N_10673,N_10375,N_10264);
xnor U10674 (N_10674,N_10367,N_10294);
and U10675 (N_10675,N_10361,N_10463);
or U10676 (N_10676,N_10384,N_10401);
xnor U10677 (N_10677,N_10472,N_10336);
nor U10678 (N_10678,N_10400,N_10493);
and U10679 (N_10679,N_10474,N_10437);
nand U10680 (N_10680,N_10458,N_10464);
or U10681 (N_10681,N_10318,N_10473);
nand U10682 (N_10682,N_10416,N_10300);
nand U10683 (N_10683,N_10339,N_10312);
nor U10684 (N_10684,N_10399,N_10478);
nor U10685 (N_10685,N_10358,N_10437);
or U10686 (N_10686,N_10251,N_10427);
nor U10687 (N_10687,N_10301,N_10457);
and U10688 (N_10688,N_10388,N_10252);
xnor U10689 (N_10689,N_10460,N_10398);
or U10690 (N_10690,N_10331,N_10270);
or U10691 (N_10691,N_10375,N_10302);
nand U10692 (N_10692,N_10306,N_10429);
and U10693 (N_10693,N_10291,N_10409);
nand U10694 (N_10694,N_10260,N_10309);
nor U10695 (N_10695,N_10284,N_10387);
nor U10696 (N_10696,N_10286,N_10253);
or U10697 (N_10697,N_10293,N_10487);
xor U10698 (N_10698,N_10478,N_10301);
or U10699 (N_10699,N_10305,N_10470);
xnor U10700 (N_10700,N_10377,N_10467);
xor U10701 (N_10701,N_10432,N_10475);
xnor U10702 (N_10702,N_10464,N_10480);
xnor U10703 (N_10703,N_10282,N_10354);
xnor U10704 (N_10704,N_10467,N_10341);
and U10705 (N_10705,N_10481,N_10261);
and U10706 (N_10706,N_10257,N_10339);
nand U10707 (N_10707,N_10498,N_10262);
xor U10708 (N_10708,N_10254,N_10332);
nor U10709 (N_10709,N_10483,N_10400);
nand U10710 (N_10710,N_10344,N_10331);
or U10711 (N_10711,N_10250,N_10270);
or U10712 (N_10712,N_10388,N_10446);
or U10713 (N_10713,N_10250,N_10300);
xnor U10714 (N_10714,N_10389,N_10356);
xor U10715 (N_10715,N_10373,N_10266);
xor U10716 (N_10716,N_10274,N_10394);
nor U10717 (N_10717,N_10285,N_10416);
and U10718 (N_10718,N_10380,N_10370);
and U10719 (N_10719,N_10472,N_10348);
nor U10720 (N_10720,N_10261,N_10367);
nand U10721 (N_10721,N_10491,N_10370);
and U10722 (N_10722,N_10392,N_10393);
and U10723 (N_10723,N_10411,N_10363);
nand U10724 (N_10724,N_10469,N_10480);
or U10725 (N_10725,N_10275,N_10336);
xor U10726 (N_10726,N_10308,N_10288);
and U10727 (N_10727,N_10355,N_10250);
and U10728 (N_10728,N_10374,N_10424);
or U10729 (N_10729,N_10477,N_10469);
nor U10730 (N_10730,N_10295,N_10492);
and U10731 (N_10731,N_10348,N_10493);
and U10732 (N_10732,N_10283,N_10271);
or U10733 (N_10733,N_10301,N_10300);
and U10734 (N_10734,N_10434,N_10369);
or U10735 (N_10735,N_10486,N_10275);
xor U10736 (N_10736,N_10468,N_10276);
nand U10737 (N_10737,N_10313,N_10375);
nor U10738 (N_10738,N_10259,N_10291);
nand U10739 (N_10739,N_10307,N_10353);
nor U10740 (N_10740,N_10425,N_10298);
and U10741 (N_10741,N_10438,N_10399);
or U10742 (N_10742,N_10314,N_10380);
and U10743 (N_10743,N_10383,N_10446);
nor U10744 (N_10744,N_10446,N_10380);
nor U10745 (N_10745,N_10323,N_10257);
nand U10746 (N_10746,N_10484,N_10460);
nand U10747 (N_10747,N_10473,N_10296);
xor U10748 (N_10748,N_10368,N_10401);
nand U10749 (N_10749,N_10328,N_10323);
and U10750 (N_10750,N_10690,N_10572);
and U10751 (N_10751,N_10501,N_10540);
nand U10752 (N_10752,N_10625,N_10581);
nor U10753 (N_10753,N_10552,N_10638);
or U10754 (N_10754,N_10648,N_10574);
xnor U10755 (N_10755,N_10582,N_10708);
nand U10756 (N_10756,N_10643,N_10590);
nand U10757 (N_10757,N_10507,N_10509);
nand U10758 (N_10758,N_10709,N_10530);
xor U10759 (N_10759,N_10550,N_10706);
nor U10760 (N_10760,N_10697,N_10533);
or U10761 (N_10761,N_10506,N_10615);
xnor U10762 (N_10762,N_10724,N_10662);
and U10763 (N_10763,N_10603,N_10632);
or U10764 (N_10764,N_10541,N_10680);
xnor U10765 (N_10765,N_10576,N_10585);
or U10766 (N_10766,N_10570,N_10536);
xor U10767 (N_10767,N_10639,N_10735);
or U10768 (N_10768,N_10586,N_10503);
and U10769 (N_10769,N_10640,N_10727);
or U10770 (N_10770,N_10584,N_10636);
nand U10771 (N_10771,N_10723,N_10525);
nand U10772 (N_10772,N_10717,N_10558);
nand U10773 (N_10773,N_10655,N_10623);
and U10774 (N_10774,N_10677,N_10654);
or U10775 (N_10775,N_10544,N_10634);
nor U10776 (N_10776,N_10714,N_10721);
xor U10777 (N_10777,N_10742,N_10713);
nor U10778 (N_10778,N_10518,N_10641);
and U10779 (N_10779,N_10629,N_10539);
nand U10780 (N_10780,N_10599,N_10656);
xor U10781 (N_10781,N_10602,N_10542);
nand U10782 (N_10782,N_10524,N_10588);
and U10783 (N_10783,N_10606,N_10647);
nand U10784 (N_10784,N_10598,N_10601);
xnor U10785 (N_10785,N_10664,N_10517);
or U10786 (N_10786,N_10705,N_10611);
and U10787 (N_10787,N_10521,N_10534);
or U10788 (N_10788,N_10748,N_10616);
nor U10789 (N_10789,N_10538,N_10564);
and U10790 (N_10790,N_10665,N_10736);
xnor U10791 (N_10791,N_10644,N_10734);
nor U10792 (N_10792,N_10679,N_10627);
nor U10793 (N_10793,N_10729,N_10553);
and U10794 (N_10794,N_10650,N_10513);
nand U10795 (N_10795,N_10591,N_10694);
and U10796 (N_10796,N_10711,N_10562);
and U10797 (N_10797,N_10739,N_10673);
xnor U10798 (N_10798,N_10569,N_10749);
xnor U10799 (N_10799,N_10670,N_10699);
nand U10800 (N_10800,N_10519,N_10728);
nor U10801 (N_10801,N_10698,N_10566);
nor U10802 (N_10802,N_10686,N_10658);
or U10803 (N_10803,N_10504,N_10505);
or U10804 (N_10804,N_10743,N_10747);
nand U10805 (N_10805,N_10689,N_10737);
nor U10806 (N_10806,N_10692,N_10730);
nand U10807 (N_10807,N_10551,N_10637);
xor U10808 (N_10808,N_10710,N_10520);
xnor U10809 (N_10809,N_10666,N_10612);
xor U10810 (N_10810,N_10614,N_10510);
and U10811 (N_10811,N_10703,N_10583);
and U10812 (N_10812,N_10682,N_10657);
nor U10813 (N_10813,N_10617,N_10594);
and U10814 (N_10814,N_10568,N_10701);
nand U10815 (N_10815,N_10565,N_10577);
xnor U10816 (N_10816,N_10628,N_10516);
nor U10817 (N_10817,N_10635,N_10649);
xor U10818 (N_10818,N_10702,N_10738);
nor U10819 (N_10819,N_10653,N_10652);
or U10820 (N_10820,N_10555,N_10684);
or U10821 (N_10821,N_10545,N_10529);
nand U10822 (N_10822,N_10531,N_10608);
nand U10823 (N_10823,N_10587,N_10549);
nor U10824 (N_10824,N_10722,N_10676);
nand U10825 (N_10825,N_10600,N_10595);
xnor U10826 (N_10826,N_10597,N_10579);
nand U10827 (N_10827,N_10573,N_10700);
nor U10828 (N_10828,N_10620,N_10546);
or U10829 (N_10829,N_10548,N_10712);
and U10830 (N_10830,N_10661,N_10646);
or U10831 (N_10831,N_10526,N_10688);
nand U10832 (N_10832,N_10642,N_10695);
nor U10833 (N_10833,N_10651,N_10745);
nand U10834 (N_10834,N_10718,N_10500);
xnor U10835 (N_10835,N_10733,N_10511);
nor U10836 (N_10836,N_10523,N_10619);
xnor U10837 (N_10837,N_10561,N_10502);
and U10838 (N_10838,N_10535,N_10557);
and U10839 (N_10839,N_10685,N_10740);
nand U10840 (N_10840,N_10580,N_10589);
nand U10841 (N_10841,N_10626,N_10659);
or U10842 (N_10842,N_10571,N_10575);
nand U10843 (N_10843,N_10528,N_10527);
or U10844 (N_10844,N_10508,N_10522);
nand U10845 (N_10845,N_10674,N_10693);
nor U10846 (N_10846,N_10567,N_10687);
or U10847 (N_10847,N_10744,N_10630);
or U10848 (N_10848,N_10725,N_10681);
or U10849 (N_10849,N_10609,N_10715);
and U10850 (N_10850,N_10691,N_10645);
and U10851 (N_10851,N_10618,N_10547);
xor U10852 (N_10852,N_10675,N_10683);
nor U10853 (N_10853,N_10593,N_10512);
or U10854 (N_10854,N_10543,N_10678);
xor U10855 (N_10855,N_10720,N_10671);
or U10856 (N_10856,N_10605,N_10672);
xor U10857 (N_10857,N_10704,N_10631);
and U10858 (N_10858,N_10604,N_10667);
and U10859 (N_10859,N_10559,N_10554);
nor U10860 (N_10860,N_10563,N_10560);
nor U10861 (N_10861,N_10622,N_10633);
nor U10862 (N_10862,N_10707,N_10624);
and U10863 (N_10863,N_10741,N_10610);
xnor U10864 (N_10864,N_10663,N_10592);
and U10865 (N_10865,N_10746,N_10613);
or U10866 (N_10866,N_10578,N_10596);
or U10867 (N_10867,N_10514,N_10556);
or U10868 (N_10868,N_10731,N_10607);
nand U10869 (N_10869,N_10532,N_10660);
nand U10870 (N_10870,N_10515,N_10669);
and U10871 (N_10871,N_10719,N_10537);
nand U10872 (N_10872,N_10726,N_10732);
nor U10873 (N_10873,N_10668,N_10696);
and U10874 (N_10874,N_10716,N_10621);
nor U10875 (N_10875,N_10723,N_10732);
xnor U10876 (N_10876,N_10736,N_10658);
nor U10877 (N_10877,N_10667,N_10678);
or U10878 (N_10878,N_10577,N_10732);
and U10879 (N_10879,N_10540,N_10537);
nand U10880 (N_10880,N_10602,N_10562);
nor U10881 (N_10881,N_10556,N_10530);
and U10882 (N_10882,N_10528,N_10694);
xor U10883 (N_10883,N_10503,N_10654);
and U10884 (N_10884,N_10546,N_10734);
nor U10885 (N_10885,N_10610,N_10720);
nor U10886 (N_10886,N_10729,N_10749);
and U10887 (N_10887,N_10658,N_10587);
nand U10888 (N_10888,N_10720,N_10708);
xnor U10889 (N_10889,N_10524,N_10614);
or U10890 (N_10890,N_10681,N_10747);
or U10891 (N_10891,N_10610,N_10691);
nor U10892 (N_10892,N_10747,N_10505);
and U10893 (N_10893,N_10500,N_10667);
nor U10894 (N_10894,N_10663,N_10748);
and U10895 (N_10895,N_10583,N_10684);
or U10896 (N_10896,N_10547,N_10647);
and U10897 (N_10897,N_10715,N_10668);
nor U10898 (N_10898,N_10581,N_10601);
or U10899 (N_10899,N_10565,N_10585);
and U10900 (N_10900,N_10599,N_10654);
or U10901 (N_10901,N_10727,N_10623);
nor U10902 (N_10902,N_10525,N_10720);
xnor U10903 (N_10903,N_10645,N_10618);
and U10904 (N_10904,N_10693,N_10507);
and U10905 (N_10905,N_10747,N_10617);
or U10906 (N_10906,N_10582,N_10603);
or U10907 (N_10907,N_10607,N_10570);
nand U10908 (N_10908,N_10610,N_10667);
nor U10909 (N_10909,N_10698,N_10639);
and U10910 (N_10910,N_10696,N_10741);
nor U10911 (N_10911,N_10739,N_10690);
and U10912 (N_10912,N_10708,N_10709);
or U10913 (N_10913,N_10542,N_10539);
xor U10914 (N_10914,N_10660,N_10718);
nand U10915 (N_10915,N_10677,N_10712);
nand U10916 (N_10916,N_10634,N_10728);
and U10917 (N_10917,N_10736,N_10732);
nand U10918 (N_10918,N_10608,N_10515);
nand U10919 (N_10919,N_10528,N_10703);
xor U10920 (N_10920,N_10706,N_10605);
nor U10921 (N_10921,N_10690,N_10676);
or U10922 (N_10922,N_10651,N_10553);
or U10923 (N_10923,N_10550,N_10686);
and U10924 (N_10924,N_10694,N_10685);
xor U10925 (N_10925,N_10711,N_10694);
and U10926 (N_10926,N_10706,N_10592);
nand U10927 (N_10927,N_10655,N_10701);
nand U10928 (N_10928,N_10701,N_10623);
and U10929 (N_10929,N_10569,N_10521);
and U10930 (N_10930,N_10656,N_10713);
nand U10931 (N_10931,N_10577,N_10605);
or U10932 (N_10932,N_10534,N_10589);
or U10933 (N_10933,N_10681,N_10542);
xor U10934 (N_10934,N_10614,N_10727);
nand U10935 (N_10935,N_10682,N_10560);
nor U10936 (N_10936,N_10652,N_10672);
or U10937 (N_10937,N_10556,N_10732);
nor U10938 (N_10938,N_10663,N_10747);
xnor U10939 (N_10939,N_10534,N_10564);
or U10940 (N_10940,N_10746,N_10553);
or U10941 (N_10941,N_10655,N_10616);
nand U10942 (N_10942,N_10531,N_10650);
nand U10943 (N_10943,N_10691,N_10537);
and U10944 (N_10944,N_10646,N_10592);
or U10945 (N_10945,N_10617,N_10585);
xor U10946 (N_10946,N_10673,N_10588);
and U10947 (N_10947,N_10698,N_10660);
nor U10948 (N_10948,N_10516,N_10533);
xor U10949 (N_10949,N_10542,N_10609);
nor U10950 (N_10950,N_10700,N_10500);
or U10951 (N_10951,N_10666,N_10525);
xnor U10952 (N_10952,N_10693,N_10653);
or U10953 (N_10953,N_10615,N_10718);
and U10954 (N_10954,N_10666,N_10738);
and U10955 (N_10955,N_10600,N_10579);
nor U10956 (N_10956,N_10545,N_10744);
nor U10957 (N_10957,N_10739,N_10678);
nor U10958 (N_10958,N_10532,N_10526);
nand U10959 (N_10959,N_10722,N_10662);
xor U10960 (N_10960,N_10593,N_10709);
xnor U10961 (N_10961,N_10739,N_10694);
xnor U10962 (N_10962,N_10744,N_10731);
and U10963 (N_10963,N_10680,N_10617);
or U10964 (N_10964,N_10645,N_10524);
and U10965 (N_10965,N_10669,N_10536);
and U10966 (N_10966,N_10676,N_10715);
and U10967 (N_10967,N_10727,N_10609);
nor U10968 (N_10968,N_10599,N_10740);
nand U10969 (N_10969,N_10635,N_10530);
and U10970 (N_10970,N_10607,N_10561);
nor U10971 (N_10971,N_10508,N_10703);
and U10972 (N_10972,N_10598,N_10642);
nor U10973 (N_10973,N_10713,N_10545);
and U10974 (N_10974,N_10701,N_10578);
or U10975 (N_10975,N_10619,N_10725);
and U10976 (N_10976,N_10612,N_10600);
or U10977 (N_10977,N_10627,N_10548);
or U10978 (N_10978,N_10683,N_10609);
xor U10979 (N_10979,N_10553,N_10556);
nand U10980 (N_10980,N_10685,N_10591);
and U10981 (N_10981,N_10566,N_10575);
or U10982 (N_10982,N_10681,N_10660);
nand U10983 (N_10983,N_10686,N_10589);
or U10984 (N_10984,N_10547,N_10553);
nand U10985 (N_10985,N_10625,N_10614);
nor U10986 (N_10986,N_10515,N_10566);
nand U10987 (N_10987,N_10581,N_10735);
nor U10988 (N_10988,N_10740,N_10501);
or U10989 (N_10989,N_10669,N_10565);
nor U10990 (N_10990,N_10675,N_10612);
nor U10991 (N_10991,N_10697,N_10725);
nor U10992 (N_10992,N_10609,N_10637);
xnor U10993 (N_10993,N_10566,N_10505);
xnor U10994 (N_10994,N_10680,N_10724);
or U10995 (N_10995,N_10698,N_10517);
or U10996 (N_10996,N_10717,N_10638);
nand U10997 (N_10997,N_10726,N_10700);
and U10998 (N_10998,N_10627,N_10582);
and U10999 (N_10999,N_10644,N_10685);
xor U11000 (N_11000,N_10874,N_10796);
and U11001 (N_11001,N_10888,N_10802);
nor U11002 (N_11002,N_10880,N_10928);
or U11003 (N_11003,N_10850,N_10933);
xnor U11004 (N_11004,N_10955,N_10757);
and U11005 (N_11005,N_10985,N_10975);
xor U11006 (N_11006,N_10769,N_10962);
nand U11007 (N_11007,N_10766,N_10792);
or U11008 (N_11008,N_10924,N_10949);
nand U11009 (N_11009,N_10883,N_10900);
nor U11010 (N_11010,N_10828,N_10848);
and U11011 (N_11011,N_10812,N_10965);
nand U11012 (N_11012,N_10830,N_10979);
nand U11013 (N_11013,N_10760,N_10956);
xor U11014 (N_11014,N_10842,N_10972);
xor U11015 (N_11015,N_10896,N_10978);
nand U11016 (N_11016,N_10858,N_10932);
xnor U11017 (N_11017,N_10934,N_10783);
xor U11018 (N_11018,N_10815,N_10887);
and U11019 (N_11019,N_10867,N_10870);
nand U11020 (N_11020,N_10776,N_10810);
nand U11021 (N_11021,N_10881,N_10781);
nor U11022 (N_11022,N_10770,N_10831);
nor U11023 (N_11023,N_10948,N_10753);
xnor U11024 (N_11024,N_10889,N_10897);
nand U11025 (N_11025,N_10873,N_10790);
and U11026 (N_11026,N_10895,N_10921);
xnor U11027 (N_11027,N_10782,N_10763);
nor U11028 (N_11028,N_10931,N_10761);
nand U11029 (N_11029,N_10898,N_10829);
xor U11030 (N_11030,N_10785,N_10989);
or U11031 (N_11031,N_10798,N_10862);
xor U11032 (N_11032,N_10852,N_10847);
and U11033 (N_11033,N_10800,N_10846);
xor U11034 (N_11034,N_10859,N_10856);
nand U11035 (N_11035,N_10839,N_10968);
and U11036 (N_11036,N_10801,N_10843);
xnor U11037 (N_11037,N_10899,N_10768);
and U11038 (N_11038,N_10803,N_10772);
xor U11039 (N_11039,N_10857,N_10844);
nor U11040 (N_11040,N_10779,N_10984);
or U11041 (N_11041,N_10780,N_10868);
or U11042 (N_11042,N_10995,N_10990);
nand U11043 (N_11043,N_10777,N_10959);
xnor U11044 (N_11044,N_10907,N_10891);
xnor U11045 (N_11045,N_10944,N_10811);
nand U11046 (N_11046,N_10813,N_10799);
and U11047 (N_11047,N_10835,N_10987);
xnor U11048 (N_11048,N_10967,N_10894);
xnor U11049 (N_11049,N_10863,N_10855);
nor U11050 (N_11050,N_10974,N_10774);
nor U11051 (N_11051,N_10939,N_10946);
nor U11052 (N_11052,N_10814,N_10773);
xor U11053 (N_11053,N_10824,N_10901);
and U11054 (N_11054,N_10877,N_10791);
xor U11055 (N_11055,N_10998,N_10886);
or U11056 (N_11056,N_10952,N_10903);
nor U11057 (N_11057,N_10795,N_10993);
nor U11058 (N_11058,N_10820,N_10927);
xor U11059 (N_11059,N_10919,N_10970);
and U11060 (N_11060,N_10971,N_10958);
nand U11061 (N_11061,N_10935,N_10864);
xor U11062 (N_11062,N_10892,N_10929);
xor U11063 (N_11063,N_10884,N_10953);
and U11064 (N_11064,N_10960,N_10797);
or U11065 (N_11065,N_10941,N_10821);
nor U11066 (N_11066,N_10966,N_10909);
or U11067 (N_11067,N_10784,N_10983);
nor U11068 (N_11068,N_10926,N_10876);
or U11069 (N_11069,N_10977,N_10865);
nor U11070 (N_11070,N_10992,N_10938);
nand U11071 (N_11071,N_10923,N_10860);
or U11072 (N_11072,N_10794,N_10981);
or U11073 (N_11073,N_10823,N_10908);
xor U11074 (N_11074,N_10912,N_10775);
and U11075 (N_11075,N_10837,N_10818);
and U11076 (N_11076,N_10754,N_10942);
xor U11077 (N_11077,N_10872,N_10804);
xor U11078 (N_11078,N_10765,N_10756);
nand U11079 (N_11079,N_10841,N_10825);
nor U11080 (N_11080,N_10902,N_10991);
nand U11081 (N_11081,N_10882,N_10916);
nand U11082 (N_11082,N_10854,N_10982);
nor U11083 (N_11083,N_10875,N_10964);
xor U11084 (N_11084,N_10890,N_10937);
nand U11085 (N_11085,N_10996,N_10834);
xnor U11086 (N_11086,N_10771,N_10807);
nand U11087 (N_11087,N_10969,N_10920);
nor U11088 (N_11088,N_10751,N_10904);
xnor U11089 (N_11089,N_10866,N_10925);
nor U11090 (N_11090,N_10947,N_10893);
and U11091 (N_11091,N_10879,N_10819);
or U11092 (N_11092,N_10914,N_10806);
and U11093 (N_11093,N_10915,N_10758);
nor U11094 (N_11094,N_10833,N_10869);
nand U11095 (N_11095,N_10845,N_10849);
nand U11096 (N_11096,N_10913,N_10822);
or U11097 (N_11097,N_10805,N_10809);
or U11098 (N_11098,N_10954,N_10861);
xor U11099 (N_11099,N_10817,N_10945);
or U11100 (N_11100,N_10762,N_10840);
xor U11101 (N_11101,N_10940,N_10816);
and U11102 (N_11102,N_10905,N_10911);
and U11103 (N_11103,N_10788,N_10853);
nand U11104 (N_11104,N_10999,N_10750);
nor U11105 (N_11105,N_10997,N_10767);
nand U11106 (N_11106,N_10917,N_10918);
and U11107 (N_11107,N_10826,N_10943);
xor U11108 (N_11108,N_10910,N_10961);
xnor U11109 (N_11109,N_10838,N_10980);
and U11110 (N_11110,N_10759,N_10930);
and U11111 (N_11111,N_10789,N_10885);
nor U11112 (N_11112,N_10936,N_10808);
xnor U11113 (N_11113,N_10786,N_10994);
nor U11114 (N_11114,N_10963,N_10973);
or U11115 (N_11115,N_10957,N_10778);
and U11116 (N_11116,N_10851,N_10906);
and U11117 (N_11117,N_10922,N_10976);
xnor U11118 (N_11118,N_10836,N_10950);
and U11119 (N_11119,N_10764,N_10986);
or U11120 (N_11120,N_10871,N_10878);
or U11121 (N_11121,N_10988,N_10832);
and U11122 (N_11122,N_10787,N_10951);
nor U11123 (N_11123,N_10755,N_10793);
and U11124 (N_11124,N_10752,N_10827);
nand U11125 (N_11125,N_10756,N_10839);
xnor U11126 (N_11126,N_10774,N_10859);
or U11127 (N_11127,N_10903,N_10917);
or U11128 (N_11128,N_10794,N_10993);
xnor U11129 (N_11129,N_10784,N_10976);
nand U11130 (N_11130,N_10770,N_10754);
or U11131 (N_11131,N_10975,N_10879);
xnor U11132 (N_11132,N_10994,N_10773);
nor U11133 (N_11133,N_10963,N_10790);
or U11134 (N_11134,N_10891,N_10758);
xnor U11135 (N_11135,N_10879,N_10954);
xor U11136 (N_11136,N_10959,N_10971);
or U11137 (N_11137,N_10773,N_10799);
xnor U11138 (N_11138,N_10936,N_10948);
nor U11139 (N_11139,N_10821,N_10795);
xnor U11140 (N_11140,N_10795,N_10884);
or U11141 (N_11141,N_10898,N_10801);
or U11142 (N_11142,N_10943,N_10871);
xor U11143 (N_11143,N_10823,N_10836);
or U11144 (N_11144,N_10775,N_10942);
nand U11145 (N_11145,N_10870,N_10882);
xnor U11146 (N_11146,N_10826,N_10873);
nand U11147 (N_11147,N_10885,N_10930);
and U11148 (N_11148,N_10819,N_10977);
xor U11149 (N_11149,N_10980,N_10824);
nor U11150 (N_11150,N_10988,N_10922);
or U11151 (N_11151,N_10998,N_10775);
xor U11152 (N_11152,N_10867,N_10991);
xor U11153 (N_11153,N_10853,N_10780);
nand U11154 (N_11154,N_10845,N_10882);
xor U11155 (N_11155,N_10994,N_10776);
nand U11156 (N_11156,N_10755,N_10759);
nand U11157 (N_11157,N_10826,N_10860);
or U11158 (N_11158,N_10770,N_10792);
or U11159 (N_11159,N_10758,N_10841);
nand U11160 (N_11160,N_10930,N_10998);
nor U11161 (N_11161,N_10851,N_10809);
nor U11162 (N_11162,N_10788,N_10845);
nand U11163 (N_11163,N_10791,N_10961);
xor U11164 (N_11164,N_10942,N_10835);
nor U11165 (N_11165,N_10765,N_10956);
nand U11166 (N_11166,N_10788,N_10773);
or U11167 (N_11167,N_10869,N_10758);
nand U11168 (N_11168,N_10811,N_10757);
and U11169 (N_11169,N_10814,N_10770);
nand U11170 (N_11170,N_10850,N_10761);
xor U11171 (N_11171,N_10862,N_10966);
or U11172 (N_11172,N_10905,N_10899);
nor U11173 (N_11173,N_10777,N_10913);
nand U11174 (N_11174,N_10950,N_10867);
xor U11175 (N_11175,N_10773,N_10968);
nand U11176 (N_11176,N_10986,N_10846);
and U11177 (N_11177,N_10990,N_10880);
nor U11178 (N_11178,N_10856,N_10828);
and U11179 (N_11179,N_10968,N_10751);
and U11180 (N_11180,N_10855,N_10989);
xnor U11181 (N_11181,N_10930,N_10952);
nand U11182 (N_11182,N_10984,N_10862);
or U11183 (N_11183,N_10861,N_10755);
nor U11184 (N_11184,N_10943,N_10763);
xor U11185 (N_11185,N_10856,N_10862);
nor U11186 (N_11186,N_10995,N_10755);
xor U11187 (N_11187,N_10758,N_10787);
or U11188 (N_11188,N_10863,N_10968);
and U11189 (N_11189,N_10953,N_10799);
or U11190 (N_11190,N_10789,N_10751);
and U11191 (N_11191,N_10830,N_10995);
and U11192 (N_11192,N_10868,N_10898);
and U11193 (N_11193,N_10821,N_10839);
nor U11194 (N_11194,N_10812,N_10762);
or U11195 (N_11195,N_10996,N_10924);
xor U11196 (N_11196,N_10913,N_10792);
xor U11197 (N_11197,N_10776,N_10812);
or U11198 (N_11198,N_10902,N_10938);
xor U11199 (N_11199,N_10755,N_10986);
and U11200 (N_11200,N_10864,N_10816);
nor U11201 (N_11201,N_10801,N_10922);
nor U11202 (N_11202,N_10902,N_10776);
xnor U11203 (N_11203,N_10906,N_10898);
and U11204 (N_11204,N_10944,N_10925);
nand U11205 (N_11205,N_10915,N_10859);
and U11206 (N_11206,N_10836,N_10812);
and U11207 (N_11207,N_10925,N_10847);
nor U11208 (N_11208,N_10915,N_10794);
nor U11209 (N_11209,N_10778,N_10939);
xor U11210 (N_11210,N_10850,N_10800);
xor U11211 (N_11211,N_10808,N_10872);
nand U11212 (N_11212,N_10775,N_10761);
xor U11213 (N_11213,N_10931,N_10915);
nor U11214 (N_11214,N_10830,N_10944);
nand U11215 (N_11215,N_10987,N_10831);
or U11216 (N_11216,N_10825,N_10974);
or U11217 (N_11217,N_10971,N_10881);
nand U11218 (N_11218,N_10832,N_10985);
xnor U11219 (N_11219,N_10884,N_10984);
nor U11220 (N_11220,N_10866,N_10960);
xor U11221 (N_11221,N_10865,N_10896);
xnor U11222 (N_11222,N_10993,N_10838);
nor U11223 (N_11223,N_10990,N_10792);
nor U11224 (N_11224,N_10802,N_10980);
nand U11225 (N_11225,N_10895,N_10781);
xnor U11226 (N_11226,N_10833,N_10755);
or U11227 (N_11227,N_10809,N_10918);
nor U11228 (N_11228,N_10980,N_10911);
nor U11229 (N_11229,N_10979,N_10983);
nor U11230 (N_11230,N_10842,N_10834);
and U11231 (N_11231,N_10843,N_10814);
xnor U11232 (N_11232,N_10803,N_10855);
xnor U11233 (N_11233,N_10827,N_10831);
nand U11234 (N_11234,N_10923,N_10869);
or U11235 (N_11235,N_10824,N_10777);
nand U11236 (N_11236,N_10897,N_10928);
nor U11237 (N_11237,N_10763,N_10907);
nor U11238 (N_11238,N_10811,N_10794);
xor U11239 (N_11239,N_10907,N_10830);
nand U11240 (N_11240,N_10966,N_10959);
nand U11241 (N_11241,N_10955,N_10920);
and U11242 (N_11242,N_10947,N_10961);
nor U11243 (N_11243,N_10911,N_10916);
nand U11244 (N_11244,N_10894,N_10991);
or U11245 (N_11245,N_10956,N_10942);
nand U11246 (N_11246,N_10793,N_10932);
xnor U11247 (N_11247,N_10855,N_10779);
nor U11248 (N_11248,N_10860,N_10789);
nor U11249 (N_11249,N_10784,N_10877);
xor U11250 (N_11250,N_11187,N_11124);
nor U11251 (N_11251,N_11155,N_11189);
nor U11252 (N_11252,N_11144,N_11142);
xor U11253 (N_11253,N_11059,N_11070);
or U11254 (N_11254,N_11015,N_11139);
nor U11255 (N_11255,N_11169,N_11052);
and U11256 (N_11256,N_11249,N_11137);
nand U11257 (N_11257,N_11192,N_11111);
or U11258 (N_11258,N_11042,N_11082);
nand U11259 (N_11259,N_11162,N_11109);
xor U11260 (N_11260,N_11180,N_11181);
nor U11261 (N_11261,N_11227,N_11229);
nor U11262 (N_11262,N_11079,N_11034);
nor U11263 (N_11263,N_11226,N_11153);
or U11264 (N_11264,N_11117,N_11010);
nor U11265 (N_11265,N_11081,N_11014);
and U11266 (N_11266,N_11149,N_11237);
nor U11267 (N_11267,N_11131,N_11043);
xnor U11268 (N_11268,N_11132,N_11016);
xnor U11269 (N_11269,N_11176,N_11200);
xor U11270 (N_11270,N_11185,N_11217);
nor U11271 (N_11271,N_11094,N_11133);
and U11272 (N_11272,N_11221,N_11123);
or U11273 (N_11273,N_11173,N_11106);
xor U11274 (N_11274,N_11045,N_11074);
nor U11275 (N_11275,N_11158,N_11108);
xor U11276 (N_11276,N_11012,N_11211);
or U11277 (N_11277,N_11178,N_11222);
nor U11278 (N_11278,N_11190,N_11095);
or U11279 (N_11279,N_11234,N_11213);
nor U11280 (N_11280,N_11056,N_11191);
or U11281 (N_11281,N_11138,N_11107);
xnor U11282 (N_11282,N_11125,N_11186);
or U11283 (N_11283,N_11203,N_11143);
nor U11284 (N_11284,N_11001,N_11044);
nand U11285 (N_11285,N_11188,N_11002);
and U11286 (N_11286,N_11197,N_11161);
or U11287 (N_11287,N_11023,N_11099);
xor U11288 (N_11288,N_11090,N_11013);
nor U11289 (N_11289,N_11242,N_11089);
nand U11290 (N_11290,N_11129,N_11019);
nand U11291 (N_11291,N_11174,N_11201);
xor U11292 (N_11292,N_11195,N_11146);
and U11293 (N_11293,N_11062,N_11047);
xnor U11294 (N_11294,N_11136,N_11127);
and U11295 (N_11295,N_11245,N_11119);
nand U11296 (N_11296,N_11154,N_11036);
and U11297 (N_11297,N_11147,N_11061);
xor U11298 (N_11298,N_11057,N_11055);
and U11299 (N_11299,N_11071,N_11004);
or U11300 (N_11300,N_11128,N_11210);
and U11301 (N_11301,N_11168,N_11038);
nor U11302 (N_11302,N_11228,N_11075);
xor U11303 (N_11303,N_11026,N_11215);
nand U11304 (N_11304,N_11231,N_11170);
nand U11305 (N_11305,N_11140,N_11239);
nand U11306 (N_11306,N_11204,N_11166);
and U11307 (N_11307,N_11098,N_11148);
xnor U11308 (N_11308,N_11066,N_11091);
nor U11309 (N_11309,N_11084,N_11244);
nor U11310 (N_11310,N_11165,N_11087);
nand U11311 (N_11311,N_11150,N_11223);
nor U11312 (N_11312,N_11048,N_11134);
and U11313 (N_11313,N_11024,N_11093);
xor U11314 (N_11314,N_11039,N_11029);
and U11315 (N_11315,N_11105,N_11060);
nand U11316 (N_11316,N_11163,N_11198);
xor U11317 (N_11317,N_11214,N_11145);
nand U11318 (N_11318,N_11160,N_11141);
nand U11319 (N_11319,N_11116,N_11050);
nor U11320 (N_11320,N_11104,N_11021);
xor U11321 (N_11321,N_11018,N_11085);
and U11322 (N_11322,N_11120,N_11035);
nand U11323 (N_11323,N_11063,N_11088);
and U11324 (N_11324,N_11030,N_11248);
nor U11325 (N_11325,N_11103,N_11046);
nor U11326 (N_11326,N_11218,N_11232);
nor U11327 (N_11327,N_11022,N_11003);
or U11328 (N_11328,N_11041,N_11179);
xnor U11329 (N_11329,N_11025,N_11073);
nand U11330 (N_11330,N_11101,N_11207);
and U11331 (N_11331,N_11183,N_11097);
nand U11332 (N_11332,N_11194,N_11112);
or U11333 (N_11333,N_11216,N_11064);
nand U11334 (N_11334,N_11065,N_11224);
nor U11335 (N_11335,N_11076,N_11028);
xor U11336 (N_11336,N_11156,N_11159);
xor U11337 (N_11337,N_11114,N_11080);
xor U11338 (N_11338,N_11037,N_11121);
nand U11339 (N_11339,N_11020,N_11077);
nor U11340 (N_11340,N_11072,N_11096);
nor U11341 (N_11341,N_11040,N_11017);
nor U11342 (N_11342,N_11068,N_11051);
xnor U11343 (N_11343,N_11122,N_11102);
xnor U11344 (N_11344,N_11175,N_11113);
xnor U11345 (N_11345,N_11135,N_11157);
and U11346 (N_11346,N_11193,N_11058);
xor U11347 (N_11347,N_11199,N_11177);
xnor U11348 (N_11348,N_11196,N_11007);
or U11349 (N_11349,N_11049,N_11205);
nand U11350 (N_11350,N_11115,N_11184);
nor U11351 (N_11351,N_11083,N_11126);
nand U11352 (N_11352,N_11247,N_11219);
nand U11353 (N_11353,N_11118,N_11092);
or U11354 (N_11354,N_11208,N_11078);
nand U11355 (N_11355,N_11009,N_11006);
nor U11356 (N_11356,N_11220,N_11067);
nor U11357 (N_11357,N_11152,N_11053);
xnor U11358 (N_11358,N_11011,N_11172);
or U11359 (N_11359,N_11171,N_11225);
xor U11360 (N_11360,N_11241,N_11240);
and U11361 (N_11361,N_11054,N_11212);
nand U11362 (N_11362,N_11243,N_11151);
or U11363 (N_11363,N_11236,N_11167);
nor U11364 (N_11364,N_11032,N_11182);
or U11365 (N_11365,N_11000,N_11202);
or U11366 (N_11366,N_11110,N_11209);
xor U11367 (N_11367,N_11033,N_11230);
and U11368 (N_11368,N_11005,N_11206);
or U11369 (N_11369,N_11233,N_11086);
xor U11370 (N_11370,N_11027,N_11235);
or U11371 (N_11371,N_11130,N_11100);
nand U11372 (N_11372,N_11238,N_11069);
nor U11373 (N_11373,N_11031,N_11164);
nor U11374 (N_11374,N_11008,N_11246);
and U11375 (N_11375,N_11217,N_11160);
nand U11376 (N_11376,N_11011,N_11173);
nor U11377 (N_11377,N_11028,N_11020);
xor U11378 (N_11378,N_11182,N_11068);
and U11379 (N_11379,N_11093,N_11180);
xnor U11380 (N_11380,N_11130,N_11121);
or U11381 (N_11381,N_11183,N_11238);
xnor U11382 (N_11382,N_11182,N_11135);
nor U11383 (N_11383,N_11093,N_11199);
xnor U11384 (N_11384,N_11050,N_11040);
and U11385 (N_11385,N_11220,N_11235);
nor U11386 (N_11386,N_11177,N_11032);
and U11387 (N_11387,N_11021,N_11190);
nand U11388 (N_11388,N_11198,N_11233);
and U11389 (N_11389,N_11131,N_11045);
or U11390 (N_11390,N_11041,N_11034);
xor U11391 (N_11391,N_11047,N_11074);
or U11392 (N_11392,N_11235,N_11001);
nor U11393 (N_11393,N_11131,N_11034);
xnor U11394 (N_11394,N_11210,N_11180);
xnor U11395 (N_11395,N_11113,N_11194);
nand U11396 (N_11396,N_11072,N_11201);
xor U11397 (N_11397,N_11146,N_11056);
xnor U11398 (N_11398,N_11164,N_11061);
xor U11399 (N_11399,N_11199,N_11124);
or U11400 (N_11400,N_11208,N_11181);
nor U11401 (N_11401,N_11196,N_11179);
xor U11402 (N_11402,N_11175,N_11225);
xnor U11403 (N_11403,N_11193,N_11233);
nor U11404 (N_11404,N_11024,N_11189);
and U11405 (N_11405,N_11247,N_11060);
nand U11406 (N_11406,N_11034,N_11099);
xnor U11407 (N_11407,N_11037,N_11026);
nand U11408 (N_11408,N_11132,N_11229);
or U11409 (N_11409,N_11199,N_11006);
nor U11410 (N_11410,N_11050,N_11231);
nor U11411 (N_11411,N_11227,N_11084);
nand U11412 (N_11412,N_11087,N_11011);
nor U11413 (N_11413,N_11241,N_11053);
nand U11414 (N_11414,N_11072,N_11198);
or U11415 (N_11415,N_11131,N_11150);
and U11416 (N_11416,N_11014,N_11232);
and U11417 (N_11417,N_11041,N_11144);
and U11418 (N_11418,N_11227,N_11009);
nand U11419 (N_11419,N_11052,N_11001);
nand U11420 (N_11420,N_11118,N_11020);
nor U11421 (N_11421,N_11025,N_11056);
and U11422 (N_11422,N_11087,N_11052);
or U11423 (N_11423,N_11060,N_11027);
or U11424 (N_11424,N_11125,N_11078);
nor U11425 (N_11425,N_11187,N_11205);
xnor U11426 (N_11426,N_11147,N_11030);
nor U11427 (N_11427,N_11061,N_11175);
nor U11428 (N_11428,N_11155,N_11135);
or U11429 (N_11429,N_11155,N_11148);
or U11430 (N_11430,N_11176,N_11249);
xnor U11431 (N_11431,N_11072,N_11066);
nand U11432 (N_11432,N_11026,N_11210);
or U11433 (N_11433,N_11247,N_11128);
nand U11434 (N_11434,N_11243,N_11185);
or U11435 (N_11435,N_11241,N_11043);
and U11436 (N_11436,N_11186,N_11083);
nand U11437 (N_11437,N_11037,N_11174);
nand U11438 (N_11438,N_11146,N_11223);
and U11439 (N_11439,N_11243,N_11123);
or U11440 (N_11440,N_11139,N_11026);
nor U11441 (N_11441,N_11026,N_11219);
nor U11442 (N_11442,N_11178,N_11121);
or U11443 (N_11443,N_11097,N_11028);
or U11444 (N_11444,N_11082,N_11017);
nand U11445 (N_11445,N_11078,N_11021);
nor U11446 (N_11446,N_11073,N_11118);
nand U11447 (N_11447,N_11154,N_11156);
or U11448 (N_11448,N_11247,N_11035);
nor U11449 (N_11449,N_11109,N_11203);
or U11450 (N_11450,N_11017,N_11139);
xor U11451 (N_11451,N_11132,N_11103);
xnor U11452 (N_11452,N_11081,N_11101);
and U11453 (N_11453,N_11121,N_11029);
xor U11454 (N_11454,N_11222,N_11183);
nand U11455 (N_11455,N_11045,N_11032);
and U11456 (N_11456,N_11086,N_11202);
xor U11457 (N_11457,N_11130,N_11206);
or U11458 (N_11458,N_11221,N_11104);
or U11459 (N_11459,N_11029,N_11024);
or U11460 (N_11460,N_11093,N_11096);
nand U11461 (N_11461,N_11115,N_11122);
or U11462 (N_11462,N_11167,N_11041);
nor U11463 (N_11463,N_11193,N_11057);
and U11464 (N_11464,N_11153,N_11051);
nand U11465 (N_11465,N_11226,N_11172);
or U11466 (N_11466,N_11188,N_11027);
xnor U11467 (N_11467,N_11222,N_11062);
nor U11468 (N_11468,N_11248,N_11008);
xor U11469 (N_11469,N_11077,N_11110);
and U11470 (N_11470,N_11067,N_11094);
or U11471 (N_11471,N_11116,N_11127);
and U11472 (N_11472,N_11003,N_11208);
xor U11473 (N_11473,N_11110,N_11107);
nor U11474 (N_11474,N_11174,N_11004);
nor U11475 (N_11475,N_11249,N_11181);
nor U11476 (N_11476,N_11248,N_11202);
and U11477 (N_11477,N_11126,N_11228);
nor U11478 (N_11478,N_11031,N_11131);
nand U11479 (N_11479,N_11177,N_11176);
xnor U11480 (N_11480,N_11113,N_11101);
nor U11481 (N_11481,N_11224,N_11069);
nand U11482 (N_11482,N_11020,N_11074);
and U11483 (N_11483,N_11058,N_11041);
or U11484 (N_11484,N_11201,N_11054);
nand U11485 (N_11485,N_11182,N_11230);
nor U11486 (N_11486,N_11071,N_11154);
or U11487 (N_11487,N_11186,N_11198);
or U11488 (N_11488,N_11075,N_11150);
nor U11489 (N_11489,N_11064,N_11205);
nor U11490 (N_11490,N_11213,N_11079);
nand U11491 (N_11491,N_11248,N_11245);
nor U11492 (N_11492,N_11135,N_11126);
or U11493 (N_11493,N_11023,N_11180);
nand U11494 (N_11494,N_11243,N_11114);
xnor U11495 (N_11495,N_11186,N_11240);
nand U11496 (N_11496,N_11218,N_11164);
xor U11497 (N_11497,N_11077,N_11143);
or U11498 (N_11498,N_11129,N_11128);
and U11499 (N_11499,N_11115,N_11049);
and U11500 (N_11500,N_11304,N_11468);
or U11501 (N_11501,N_11305,N_11393);
and U11502 (N_11502,N_11269,N_11499);
nor U11503 (N_11503,N_11358,N_11367);
and U11504 (N_11504,N_11282,N_11364);
nand U11505 (N_11505,N_11251,N_11397);
or U11506 (N_11506,N_11497,N_11326);
xnor U11507 (N_11507,N_11341,N_11257);
and U11508 (N_11508,N_11403,N_11265);
nand U11509 (N_11509,N_11391,N_11441);
xnor U11510 (N_11510,N_11431,N_11464);
nor U11511 (N_11511,N_11267,N_11261);
and U11512 (N_11512,N_11423,N_11365);
or U11513 (N_11513,N_11357,N_11350);
or U11514 (N_11514,N_11334,N_11417);
and U11515 (N_11515,N_11458,N_11498);
xor U11516 (N_11516,N_11467,N_11487);
nand U11517 (N_11517,N_11363,N_11321);
and U11518 (N_11518,N_11409,N_11413);
and U11519 (N_11519,N_11308,N_11402);
or U11520 (N_11520,N_11454,N_11366);
nor U11521 (N_11521,N_11325,N_11399);
and U11522 (N_11522,N_11395,N_11340);
and U11523 (N_11523,N_11448,N_11408);
xor U11524 (N_11524,N_11373,N_11262);
xor U11525 (N_11525,N_11436,N_11411);
nor U11526 (N_11526,N_11488,N_11300);
nand U11527 (N_11527,N_11432,N_11404);
nor U11528 (N_11528,N_11465,N_11478);
and U11529 (N_11529,N_11359,N_11461);
nor U11530 (N_11530,N_11283,N_11443);
and U11531 (N_11531,N_11285,N_11361);
xor U11532 (N_11532,N_11276,N_11485);
nand U11533 (N_11533,N_11462,N_11424);
nor U11534 (N_11534,N_11456,N_11306);
nor U11535 (N_11535,N_11475,N_11290);
nand U11536 (N_11536,N_11375,N_11319);
or U11537 (N_11537,N_11287,N_11278);
and U11538 (N_11538,N_11444,N_11386);
nand U11539 (N_11539,N_11253,N_11320);
nor U11540 (N_11540,N_11442,N_11437);
or U11541 (N_11541,N_11400,N_11260);
and U11542 (N_11542,N_11451,N_11296);
or U11543 (N_11543,N_11310,N_11491);
and U11544 (N_11544,N_11303,N_11299);
nor U11545 (N_11545,N_11470,N_11472);
or U11546 (N_11546,N_11414,N_11463);
nor U11547 (N_11547,N_11396,N_11473);
nand U11548 (N_11548,N_11494,N_11374);
and U11549 (N_11549,N_11314,N_11279);
xor U11550 (N_11550,N_11312,N_11309);
and U11551 (N_11551,N_11422,N_11415);
and U11552 (N_11552,N_11425,N_11383);
nor U11553 (N_11553,N_11493,N_11480);
and U11554 (N_11554,N_11412,N_11410);
or U11555 (N_11555,N_11457,N_11489);
or U11556 (N_11556,N_11370,N_11484);
nand U11557 (N_11557,N_11297,N_11416);
and U11558 (N_11558,N_11378,N_11483);
nand U11559 (N_11559,N_11335,N_11281);
nand U11560 (N_11560,N_11254,N_11496);
or U11561 (N_11561,N_11407,N_11250);
nor U11562 (N_11562,N_11460,N_11455);
nor U11563 (N_11563,N_11259,N_11268);
nand U11564 (N_11564,N_11384,N_11471);
and U11565 (N_11565,N_11405,N_11330);
nor U11566 (N_11566,N_11434,N_11353);
nor U11567 (N_11567,N_11392,N_11453);
xnor U11568 (N_11568,N_11495,N_11270);
and U11569 (N_11569,N_11430,N_11286);
nor U11570 (N_11570,N_11284,N_11387);
or U11571 (N_11571,N_11302,N_11377);
nand U11572 (N_11572,N_11349,N_11332);
and U11573 (N_11573,N_11371,N_11311);
nor U11574 (N_11574,N_11433,N_11427);
and U11575 (N_11575,N_11333,N_11394);
nor U11576 (N_11576,N_11295,N_11482);
xnor U11577 (N_11577,N_11360,N_11362);
nand U11578 (N_11578,N_11338,N_11490);
and U11579 (N_11579,N_11273,N_11420);
nor U11580 (N_11580,N_11301,N_11264);
nor U11581 (N_11581,N_11385,N_11271);
nor U11582 (N_11582,N_11318,N_11439);
and U11583 (N_11583,N_11351,N_11336);
xnor U11584 (N_11584,N_11298,N_11292);
nor U11585 (N_11585,N_11354,N_11401);
xor U11586 (N_11586,N_11263,N_11342);
xnor U11587 (N_11587,N_11258,N_11376);
nand U11588 (N_11588,N_11328,N_11315);
xnor U11589 (N_11589,N_11343,N_11438);
and U11590 (N_11590,N_11355,N_11380);
xor U11591 (N_11591,N_11452,N_11347);
nand U11592 (N_11592,N_11346,N_11313);
nand U11593 (N_11593,N_11449,N_11293);
nor U11594 (N_11594,N_11288,N_11345);
or U11595 (N_11595,N_11450,N_11289);
nand U11596 (N_11596,N_11469,N_11419);
nor U11597 (N_11597,N_11479,N_11481);
or U11598 (N_11598,N_11274,N_11322);
xor U11599 (N_11599,N_11317,N_11428);
xor U11600 (N_11600,N_11372,N_11388);
xnor U11601 (N_11601,N_11382,N_11277);
and U11602 (N_11602,N_11406,N_11323);
or U11603 (N_11603,N_11348,N_11356);
nor U11604 (N_11604,N_11256,N_11369);
and U11605 (N_11605,N_11418,N_11255);
nor U11606 (N_11606,N_11344,N_11492);
nand U11607 (N_11607,N_11389,N_11316);
or U11608 (N_11608,N_11474,N_11280);
and U11609 (N_11609,N_11294,N_11331);
and U11610 (N_11610,N_11291,N_11275);
nor U11611 (N_11611,N_11379,N_11307);
nor U11612 (N_11612,N_11435,N_11459);
or U11613 (N_11613,N_11329,N_11368);
nand U11614 (N_11614,N_11440,N_11447);
and U11615 (N_11615,N_11429,N_11252);
nor U11616 (N_11616,N_11352,N_11327);
and U11617 (N_11617,N_11266,N_11486);
and U11618 (N_11618,N_11381,N_11476);
nand U11619 (N_11619,N_11477,N_11426);
xor U11620 (N_11620,N_11337,N_11339);
nor U11621 (N_11621,N_11445,N_11390);
nand U11622 (N_11622,N_11324,N_11272);
and U11623 (N_11623,N_11421,N_11446);
nand U11624 (N_11624,N_11398,N_11466);
nand U11625 (N_11625,N_11404,N_11316);
nor U11626 (N_11626,N_11468,N_11459);
xnor U11627 (N_11627,N_11479,N_11290);
nand U11628 (N_11628,N_11453,N_11344);
or U11629 (N_11629,N_11489,N_11383);
xor U11630 (N_11630,N_11400,N_11490);
and U11631 (N_11631,N_11420,N_11339);
and U11632 (N_11632,N_11459,N_11284);
nor U11633 (N_11633,N_11493,N_11399);
or U11634 (N_11634,N_11417,N_11393);
nand U11635 (N_11635,N_11320,N_11321);
or U11636 (N_11636,N_11473,N_11250);
or U11637 (N_11637,N_11476,N_11423);
nor U11638 (N_11638,N_11439,N_11360);
or U11639 (N_11639,N_11334,N_11499);
and U11640 (N_11640,N_11498,N_11387);
and U11641 (N_11641,N_11338,N_11309);
nand U11642 (N_11642,N_11405,N_11452);
xor U11643 (N_11643,N_11430,N_11257);
and U11644 (N_11644,N_11291,N_11448);
xor U11645 (N_11645,N_11472,N_11336);
nand U11646 (N_11646,N_11274,N_11427);
and U11647 (N_11647,N_11446,N_11392);
nand U11648 (N_11648,N_11472,N_11291);
nand U11649 (N_11649,N_11336,N_11428);
nor U11650 (N_11650,N_11423,N_11276);
nand U11651 (N_11651,N_11336,N_11402);
nor U11652 (N_11652,N_11314,N_11400);
nand U11653 (N_11653,N_11482,N_11253);
or U11654 (N_11654,N_11447,N_11446);
xor U11655 (N_11655,N_11467,N_11300);
or U11656 (N_11656,N_11396,N_11349);
or U11657 (N_11657,N_11459,N_11286);
xor U11658 (N_11658,N_11258,N_11413);
and U11659 (N_11659,N_11405,N_11327);
nand U11660 (N_11660,N_11385,N_11470);
xnor U11661 (N_11661,N_11366,N_11452);
or U11662 (N_11662,N_11400,N_11416);
or U11663 (N_11663,N_11468,N_11450);
or U11664 (N_11664,N_11493,N_11428);
and U11665 (N_11665,N_11284,N_11382);
xnor U11666 (N_11666,N_11414,N_11396);
or U11667 (N_11667,N_11492,N_11430);
xnor U11668 (N_11668,N_11382,N_11372);
or U11669 (N_11669,N_11416,N_11272);
nand U11670 (N_11670,N_11298,N_11344);
nand U11671 (N_11671,N_11290,N_11396);
nor U11672 (N_11672,N_11340,N_11365);
or U11673 (N_11673,N_11385,N_11406);
xnor U11674 (N_11674,N_11412,N_11288);
xor U11675 (N_11675,N_11420,N_11284);
and U11676 (N_11676,N_11413,N_11459);
xnor U11677 (N_11677,N_11346,N_11341);
and U11678 (N_11678,N_11259,N_11482);
nor U11679 (N_11679,N_11492,N_11268);
nor U11680 (N_11680,N_11285,N_11253);
or U11681 (N_11681,N_11382,N_11338);
and U11682 (N_11682,N_11392,N_11299);
and U11683 (N_11683,N_11482,N_11498);
and U11684 (N_11684,N_11268,N_11462);
nand U11685 (N_11685,N_11316,N_11350);
nor U11686 (N_11686,N_11427,N_11422);
and U11687 (N_11687,N_11446,N_11490);
nor U11688 (N_11688,N_11477,N_11483);
nand U11689 (N_11689,N_11426,N_11311);
xor U11690 (N_11690,N_11437,N_11457);
or U11691 (N_11691,N_11324,N_11259);
nand U11692 (N_11692,N_11354,N_11309);
or U11693 (N_11693,N_11276,N_11250);
nor U11694 (N_11694,N_11325,N_11439);
nor U11695 (N_11695,N_11281,N_11428);
xnor U11696 (N_11696,N_11335,N_11339);
or U11697 (N_11697,N_11302,N_11331);
nor U11698 (N_11698,N_11443,N_11337);
nand U11699 (N_11699,N_11420,N_11471);
or U11700 (N_11700,N_11457,N_11384);
nand U11701 (N_11701,N_11365,N_11486);
and U11702 (N_11702,N_11482,N_11313);
nand U11703 (N_11703,N_11407,N_11455);
nor U11704 (N_11704,N_11361,N_11391);
xor U11705 (N_11705,N_11438,N_11325);
and U11706 (N_11706,N_11461,N_11410);
xnor U11707 (N_11707,N_11314,N_11484);
nand U11708 (N_11708,N_11257,N_11348);
nand U11709 (N_11709,N_11427,N_11383);
or U11710 (N_11710,N_11447,N_11258);
nand U11711 (N_11711,N_11461,N_11371);
xnor U11712 (N_11712,N_11379,N_11298);
and U11713 (N_11713,N_11397,N_11312);
nand U11714 (N_11714,N_11331,N_11266);
and U11715 (N_11715,N_11353,N_11279);
nor U11716 (N_11716,N_11312,N_11493);
or U11717 (N_11717,N_11473,N_11411);
xor U11718 (N_11718,N_11285,N_11321);
nand U11719 (N_11719,N_11332,N_11294);
nand U11720 (N_11720,N_11278,N_11477);
nand U11721 (N_11721,N_11280,N_11476);
or U11722 (N_11722,N_11384,N_11441);
nand U11723 (N_11723,N_11335,N_11367);
or U11724 (N_11724,N_11481,N_11467);
nor U11725 (N_11725,N_11349,N_11466);
and U11726 (N_11726,N_11466,N_11411);
or U11727 (N_11727,N_11251,N_11374);
and U11728 (N_11728,N_11291,N_11443);
nor U11729 (N_11729,N_11315,N_11334);
or U11730 (N_11730,N_11472,N_11456);
nor U11731 (N_11731,N_11428,N_11398);
xnor U11732 (N_11732,N_11343,N_11347);
nand U11733 (N_11733,N_11431,N_11324);
nor U11734 (N_11734,N_11275,N_11494);
nor U11735 (N_11735,N_11457,N_11258);
and U11736 (N_11736,N_11486,N_11426);
nor U11737 (N_11737,N_11317,N_11309);
xnor U11738 (N_11738,N_11289,N_11496);
and U11739 (N_11739,N_11418,N_11291);
or U11740 (N_11740,N_11423,N_11329);
xnor U11741 (N_11741,N_11483,N_11415);
nor U11742 (N_11742,N_11346,N_11415);
xor U11743 (N_11743,N_11345,N_11253);
xor U11744 (N_11744,N_11339,N_11360);
nor U11745 (N_11745,N_11320,N_11427);
nor U11746 (N_11746,N_11324,N_11278);
or U11747 (N_11747,N_11293,N_11482);
xnor U11748 (N_11748,N_11372,N_11341);
and U11749 (N_11749,N_11448,N_11407);
or U11750 (N_11750,N_11518,N_11685);
and U11751 (N_11751,N_11660,N_11700);
nor U11752 (N_11752,N_11571,N_11636);
and U11753 (N_11753,N_11505,N_11572);
xnor U11754 (N_11754,N_11525,N_11677);
nand U11755 (N_11755,N_11510,N_11578);
or U11756 (N_11756,N_11520,N_11729);
nand U11757 (N_11757,N_11611,N_11604);
xnor U11758 (N_11758,N_11720,N_11621);
xor U11759 (N_11759,N_11693,N_11589);
xnor U11760 (N_11760,N_11575,N_11674);
xnor U11761 (N_11761,N_11620,N_11561);
nand U11762 (N_11762,N_11539,N_11509);
nor U11763 (N_11763,N_11570,N_11635);
xor U11764 (N_11764,N_11567,N_11516);
and U11765 (N_11765,N_11629,N_11634);
and U11766 (N_11766,N_11647,N_11601);
and U11767 (N_11767,N_11632,N_11627);
xor U11768 (N_11768,N_11569,N_11663);
nand U11769 (N_11769,N_11603,N_11612);
nor U11770 (N_11770,N_11545,N_11557);
and U11771 (N_11771,N_11594,N_11548);
nand U11772 (N_11772,N_11556,N_11513);
and U11773 (N_11773,N_11640,N_11686);
xor U11774 (N_11774,N_11695,N_11623);
nor U11775 (N_11775,N_11533,N_11559);
or U11776 (N_11776,N_11746,N_11566);
nand U11777 (N_11777,N_11667,N_11590);
nand U11778 (N_11778,N_11526,N_11535);
or U11779 (N_11779,N_11669,N_11713);
xnor U11780 (N_11780,N_11717,N_11564);
or U11781 (N_11781,N_11645,N_11684);
or U11782 (N_11782,N_11642,N_11732);
nand U11783 (N_11783,N_11507,N_11501);
or U11784 (N_11784,N_11678,N_11527);
nor U11785 (N_11785,N_11692,N_11522);
nor U11786 (N_11786,N_11641,N_11740);
nand U11787 (N_11787,N_11600,N_11551);
nor U11788 (N_11788,N_11748,N_11698);
and U11789 (N_11789,N_11679,N_11649);
and U11790 (N_11790,N_11715,N_11552);
and U11791 (N_11791,N_11710,N_11585);
nor U11792 (N_11792,N_11653,N_11714);
nand U11793 (N_11793,N_11719,N_11579);
xor U11794 (N_11794,N_11689,N_11741);
and U11795 (N_11795,N_11705,N_11616);
and U11796 (N_11796,N_11697,N_11565);
and U11797 (N_11797,N_11736,N_11614);
xor U11798 (N_11798,N_11680,N_11576);
nor U11799 (N_11799,N_11630,N_11506);
and U11800 (N_11800,N_11671,N_11596);
xnor U11801 (N_11801,N_11721,N_11595);
xor U11802 (N_11802,N_11665,N_11696);
nand U11803 (N_11803,N_11704,N_11711);
nand U11804 (N_11804,N_11703,N_11592);
nand U11805 (N_11805,N_11555,N_11706);
nor U11806 (N_11806,N_11724,N_11744);
and U11807 (N_11807,N_11659,N_11519);
and U11808 (N_11808,N_11615,N_11568);
nand U11809 (N_11809,N_11581,N_11666);
xor U11810 (N_11810,N_11587,N_11699);
and U11811 (N_11811,N_11728,N_11718);
or U11812 (N_11812,N_11544,N_11707);
xor U11813 (N_11813,N_11676,N_11633);
nor U11814 (N_11814,N_11738,N_11530);
or U11815 (N_11815,N_11747,N_11608);
nor U11816 (N_11816,N_11625,N_11673);
and U11817 (N_11817,N_11577,N_11500);
or U11818 (N_11818,N_11716,N_11683);
nor U11819 (N_11819,N_11584,N_11737);
and U11820 (N_11820,N_11708,N_11504);
xor U11821 (N_11821,N_11722,N_11543);
nor U11822 (N_11822,N_11681,N_11534);
nand U11823 (N_11823,N_11605,N_11538);
nand U11824 (N_11824,N_11658,N_11515);
nor U11825 (N_11825,N_11588,N_11661);
or U11826 (N_11826,N_11512,N_11687);
xor U11827 (N_11827,N_11610,N_11537);
nor U11828 (N_11828,N_11524,N_11734);
or U11829 (N_11829,N_11550,N_11726);
nor U11830 (N_11830,N_11531,N_11591);
or U11831 (N_11831,N_11624,N_11709);
or U11832 (N_11832,N_11514,N_11691);
and U11833 (N_11833,N_11563,N_11743);
nand U11834 (N_11834,N_11739,N_11668);
nor U11835 (N_11835,N_11725,N_11637);
or U11836 (N_11836,N_11727,N_11656);
xor U11837 (N_11837,N_11517,N_11688);
nor U11838 (N_11838,N_11597,N_11626);
or U11839 (N_11839,N_11731,N_11502);
xor U11840 (N_11840,N_11733,N_11593);
nor U11841 (N_11841,N_11554,N_11558);
nor U11842 (N_11842,N_11638,N_11583);
or U11843 (N_11843,N_11639,N_11723);
xnor U11844 (N_11844,N_11646,N_11690);
nand U11845 (N_11845,N_11602,N_11682);
and U11846 (N_11846,N_11523,N_11609);
xnor U11847 (N_11847,N_11618,N_11546);
xnor U11848 (N_11848,N_11655,N_11650);
or U11849 (N_11849,N_11654,N_11701);
or U11850 (N_11850,N_11712,N_11619);
xor U11851 (N_11851,N_11670,N_11622);
and U11852 (N_11852,N_11573,N_11528);
and U11853 (N_11853,N_11606,N_11617);
or U11854 (N_11854,N_11730,N_11742);
and U11855 (N_11855,N_11613,N_11529);
xor U11856 (N_11856,N_11511,N_11652);
xor U11857 (N_11857,N_11749,N_11657);
nor U11858 (N_11858,N_11503,N_11745);
nor U11859 (N_11859,N_11648,N_11508);
or U11860 (N_11860,N_11547,N_11664);
or U11861 (N_11861,N_11702,N_11651);
xnor U11862 (N_11862,N_11599,N_11562);
and U11863 (N_11863,N_11580,N_11607);
nand U11864 (N_11864,N_11549,N_11598);
xnor U11865 (N_11865,N_11644,N_11675);
nand U11866 (N_11866,N_11662,N_11574);
or U11867 (N_11867,N_11540,N_11582);
xnor U11868 (N_11868,N_11631,N_11643);
nor U11869 (N_11869,N_11541,N_11532);
nand U11870 (N_11870,N_11542,N_11628);
nor U11871 (N_11871,N_11553,N_11536);
nor U11872 (N_11872,N_11735,N_11521);
nor U11873 (N_11873,N_11672,N_11586);
and U11874 (N_11874,N_11560,N_11694);
or U11875 (N_11875,N_11584,N_11553);
and U11876 (N_11876,N_11699,N_11559);
xnor U11877 (N_11877,N_11661,N_11701);
nand U11878 (N_11878,N_11518,N_11613);
or U11879 (N_11879,N_11733,N_11723);
or U11880 (N_11880,N_11561,N_11549);
and U11881 (N_11881,N_11642,N_11581);
or U11882 (N_11882,N_11576,N_11711);
xor U11883 (N_11883,N_11654,N_11658);
nand U11884 (N_11884,N_11626,N_11674);
nor U11885 (N_11885,N_11675,N_11587);
or U11886 (N_11886,N_11668,N_11586);
nor U11887 (N_11887,N_11706,N_11539);
and U11888 (N_11888,N_11645,N_11710);
or U11889 (N_11889,N_11567,N_11728);
nand U11890 (N_11890,N_11544,N_11597);
nor U11891 (N_11891,N_11739,N_11629);
nor U11892 (N_11892,N_11632,N_11586);
and U11893 (N_11893,N_11628,N_11598);
and U11894 (N_11894,N_11538,N_11582);
and U11895 (N_11895,N_11619,N_11562);
nor U11896 (N_11896,N_11577,N_11705);
nor U11897 (N_11897,N_11607,N_11645);
nor U11898 (N_11898,N_11540,N_11601);
xor U11899 (N_11899,N_11541,N_11699);
and U11900 (N_11900,N_11536,N_11679);
and U11901 (N_11901,N_11625,N_11676);
and U11902 (N_11902,N_11650,N_11519);
and U11903 (N_11903,N_11563,N_11714);
xor U11904 (N_11904,N_11656,N_11706);
or U11905 (N_11905,N_11680,N_11577);
nor U11906 (N_11906,N_11520,N_11656);
nor U11907 (N_11907,N_11740,N_11645);
nand U11908 (N_11908,N_11678,N_11646);
or U11909 (N_11909,N_11541,N_11571);
xor U11910 (N_11910,N_11729,N_11672);
or U11911 (N_11911,N_11530,N_11647);
nor U11912 (N_11912,N_11593,N_11512);
nand U11913 (N_11913,N_11647,N_11582);
or U11914 (N_11914,N_11658,N_11604);
or U11915 (N_11915,N_11640,N_11732);
or U11916 (N_11916,N_11633,N_11610);
nand U11917 (N_11917,N_11708,N_11698);
nand U11918 (N_11918,N_11569,N_11588);
or U11919 (N_11919,N_11508,N_11742);
nand U11920 (N_11920,N_11533,N_11652);
xnor U11921 (N_11921,N_11535,N_11585);
or U11922 (N_11922,N_11536,N_11666);
xor U11923 (N_11923,N_11681,N_11531);
nand U11924 (N_11924,N_11594,N_11696);
nor U11925 (N_11925,N_11543,N_11653);
nor U11926 (N_11926,N_11505,N_11592);
and U11927 (N_11927,N_11565,N_11719);
xor U11928 (N_11928,N_11581,N_11730);
or U11929 (N_11929,N_11697,N_11654);
nand U11930 (N_11930,N_11620,N_11744);
and U11931 (N_11931,N_11653,N_11538);
xor U11932 (N_11932,N_11734,N_11597);
and U11933 (N_11933,N_11594,N_11699);
nor U11934 (N_11934,N_11667,N_11641);
or U11935 (N_11935,N_11601,N_11714);
nor U11936 (N_11936,N_11586,N_11513);
and U11937 (N_11937,N_11607,N_11726);
or U11938 (N_11938,N_11674,N_11591);
xor U11939 (N_11939,N_11700,N_11541);
xor U11940 (N_11940,N_11509,N_11553);
or U11941 (N_11941,N_11541,N_11662);
or U11942 (N_11942,N_11683,N_11523);
nor U11943 (N_11943,N_11550,N_11500);
xnor U11944 (N_11944,N_11681,N_11623);
xor U11945 (N_11945,N_11591,N_11512);
nand U11946 (N_11946,N_11707,N_11702);
or U11947 (N_11947,N_11520,N_11748);
nor U11948 (N_11948,N_11686,N_11564);
xnor U11949 (N_11949,N_11737,N_11601);
or U11950 (N_11950,N_11596,N_11527);
xor U11951 (N_11951,N_11567,N_11690);
and U11952 (N_11952,N_11505,N_11685);
nand U11953 (N_11953,N_11519,N_11661);
xor U11954 (N_11954,N_11637,N_11722);
or U11955 (N_11955,N_11684,N_11578);
xnor U11956 (N_11956,N_11528,N_11613);
xnor U11957 (N_11957,N_11632,N_11509);
and U11958 (N_11958,N_11610,N_11580);
or U11959 (N_11959,N_11692,N_11722);
nand U11960 (N_11960,N_11573,N_11613);
or U11961 (N_11961,N_11700,N_11527);
nor U11962 (N_11962,N_11551,N_11626);
nor U11963 (N_11963,N_11583,N_11546);
or U11964 (N_11964,N_11680,N_11604);
and U11965 (N_11965,N_11510,N_11676);
nor U11966 (N_11966,N_11600,N_11579);
and U11967 (N_11967,N_11507,N_11584);
and U11968 (N_11968,N_11513,N_11524);
nand U11969 (N_11969,N_11585,N_11681);
nand U11970 (N_11970,N_11649,N_11662);
and U11971 (N_11971,N_11748,N_11727);
nand U11972 (N_11972,N_11532,N_11633);
nand U11973 (N_11973,N_11737,N_11682);
and U11974 (N_11974,N_11512,N_11638);
nor U11975 (N_11975,N_11712,N_11545);
nand U11976 (N_11976,N_11604,N_11551);
nand U11977 (N_11977,N_11523,N_11700);
nor U11978 (N_11978,N_11559,N_11689);
and U11979 (N_11979,N_11599,N_11616);
xnor U11980 (N_11980,N_11616,N_11620);
nor U11981 (N_11981,N_11607,N_11606);
nand U11982 (N_11982,N_11523,N_11549);
nand U11983 (N_11983,N_11637,N_11609);
or U11984 (N_11984,N_11635,N_11537);
and U11985 (N_11985,N_11701,N_11510);
nor U11986 (N_11986,N_11582,N_11607);
nor U11987 (N_11987,N_11682,N_11558);
or U11988 (N_11988,N_11729,N_11601);
nor U11989 (N_11989,N_11614,N_11716);
xnor U11990 (N_11990,N_11734,N_11649);
and U11991 (N_11991,N_11598,N_11742);
nor U11992 (N_11992,N_11716,N_11505);
and U11993 (N_11993,N_11601,N_11684);
or U11994 (N_11994,N_11575,N_11549);
and U11995 (N_11995,N_11717,N_11652);
and U11996 (N_11996,N_11571,N_11672);
xor U11997 (N_11997,N_11733,N_11501);
xor U11998 (N_11998,N_11524,N_11709);
or U11999 (N_11999,N_11731,N_11709);
and U12000 (N_12000,N_11828,N_11984);
or U12001 (N_12001,N_11813,N_11802);
xor U12002 (N_12002,N_11810,N_11833);
nand U12003 (N_12003,N_11988,N_11985);
nor U12004 (N_12004,N_11896,N_11788);
xnor U12005 (N_12005,N_11950,N_11934);
xor U12006 (N_12006,N_11768,N_11811);
and U12007 (N_12007,N_11889,N_11752);
or U12008 (N_12008,N_11754,N_11904);
or U12009 (N_12009,N_11977,N_11852);
and U12010 (N_12010,N_11817,N_11758);
or U12011 (N_12011,N_11910,N_11829);
xnor U12012 (N_12012,N_11793,N_11875);
or U12013 (N_12013,N_11902,N_11860);
and U12014 (N_12014,N_11916,N_11960);
xnor U12015 (N_12015,N_11967,N_11929);
or U12016 (N_12016,N_11812,N_11785);
or U12017 (N_12017,N_11803,N_11994);
xnor U12018 (N_12018,N_11932,N_11789);
nor U12019 (N_12019,N_11830,N_11972);
nand U12020 (N_12020,N_11771,N_11973);
nor U12021 (N_12021,N_11907,N_11770);
nor U12022 (N_12022,N_11931,N_11870);
or U12023 (N_12023,N_11766,N_11757);
and U12024 (N_12024,N_11790,N_11877);
nand U12025 (N_12025,N_11952,N_11781);
xnor U12026 (N_12026,N_11996,N_11814);
xor U12027 (N_12027,N_11778,N_11943);
nor U12028 (N_12028,N_11968,N_11762);
or U12029 (N_12029,N_11843,N_11981);
nor U12030 (N_12030,N_11854,N_11782);
xor U12031 (N_12031,N_11888,N_11837);
or U12032 (N_12032,N_11964,N_11826);
nor U12033 (N_12033,N_11901,N_11897);
nor U12034 (N_12034,N_11962,N_11776);
nor U12035 (N_12035,N_11940,N_11992);
nor U12036 (N_12036,N_11918,N_11956);
xnor U12037 (N_12037,N_11945,N_11874);
and U12038 (N_12038,N_11755,N_11818);
or U12039 (N_12039,N_11947,N_11844);
xor U12040 (N_12040,N_11795,N_11941);
nor U12041 (N_12041,N_11991,N_11938);
or U12042 (N_12042,N_11961,N_11989);
nand U12043 (N_12043,N_11857,N_11753);
xor U12044 (N_12044,N_11908,N_11851);
xnor U12045 (N_12045,N_11796,N_11858);
xnor U12046 (N_12046,N_11775,N_11825);
nand U12047 (N_12047,N_11871,N_11765);
nand U12048 (N_12048,N_11800,N_11784);
nand U12049 (N_12049,N_11832,N_11933);
nor U12050 (N_12050,N_11998,N_11944);
xnor U12051 (N_12051,N_11999,N_11884);
and U12052 (N_12052,N_11773,N_11866);
nand U12053 (N_12053,N_11921,N_11926);
and U12054 (N_12054,N_11986,N_11850);
xnor U12055 (N_12055,N_11979,N_11808);
or U12056 (N_12056,N_11935,N_11970);
nand U12057 (N_12057,N_11848,N_11946);
xnor U12058 (N_12058,N_11914,N_11925);
nand U12059 (N_12059,N_11867,N_11879);
nor U12060 (N_12060,N_11792,N_11899);
nor U12061 (N_12061,N_11955,N_11807);
nor U12062 (N_12062,N_11764,N_11855);
nor U12063 (N_12063,N_11783,N_11797);
and U12064 (N_12064,N_11868,N_11791);
or U12065 (N_12065,N_11786,N_11856);
and U12066 (N_12066,N_11835,N_11975);
nor U12067 (N_12067,N_11815,N_11769);
xnor U12068 (N_12068,N_11898,N_11920);
nand U12069 (N_12069,N_11980,N_11903);
nand U12070 (N_12070,N_11767,N_11834);
nor U12071 (N_12071,N_11913,N_11772);
and U12072 (N_12072,N_11824,N_11982);
or U12073 (N_12073,N_11862,N_11993);
or U12074 (N_12074,N_11891,N_11930);
and U12075 (N_12075,N_11959,N_11819);
and U12076 (N_12076,N_11839,N_11777);
nor U12077 (N_12077,N_11780,N_11948);
nor U12078 (N_12078,N_11936,N_11847);
nand U12079 (N_12079,N_11804,N_11997);
or U12080 (N_12080,N_11756,N_11823);
nand U12081 (N_12081,N_11774,N_11845);
or U12082 (N_12082,N_11881,N_11840);
xnor U12083 (N_12083,N_11987,N_11859);
xor U12084 (N_12084,N_11954,N_11882);
nor U12085 (N_12085,N_11760,N_11895);
nand U12086 (N_12086,N_11939,N_11915);
nor U12087 (N_12087,N_11893,N_11953);
nand U12088 (N_12088,N_11969,N_11836);
or U12089 (N_12089,N_11861,N_11806);
nor U12090 (N_12090,N_11876,N_11827);
nor U12091 (N_12091,N_11849,N_11809);
and U12092 (N_12092,N_11917,N_11957);
nand U12093 (N_12093,N_11872,N_11923);
nor U12094 (N_12094,N_11798,N_11846);
or U12095 (N_12095,N_11937,N_11942);
and U12096 (N_12096,N_11906,N_11822);
and U12097 (N_12097,N_11900,N_11878);
and U12098 (N_12098,N_11842,N_11787);
xnor U12099 (N_12099,N_11863,N_11909);
xnor U12100 (N_12100,N_11966,N_11759);
nand U12101 (N_12101,N_11761,N_11750);
xor U12102 (N_12102,N_11873,N_11922);
nand U12103 (N_12103,N_11949,N_11838);
nand U12104 (N_12104,N_11864,N_11885);
xnor U12105 (N_12105,N_11794,N_11971);
and U12106 (N_12106,N_11865,N_11912);
and U12107 (N_12107,N_11958,N_11751);
xor U12108 (N_12108,N_11919,N_11983);
or U12109 (N_12109,N_11894,N_11805);
xor U12110 (N_12110,N_11841,N_11963);
and U12111 (N_12111,N_11990,N_11974);
nand U12112 (N_12112,N_11831,N_11965);
or U12113 (N_12113,N_11880,N_11927);
nand U12114 (N_12114,N_11911,N_11821);
xnor U12115 (N_12115,N_11924,N_11886);
nand U12116 (N_12116,N_11799,N_11890);
nor U12117 (N_12117,N_11816,N_11976);
nand U12118 (N_12118,N_11978,N_11801);
nor U12119 (N_12119,N_11951,N_11779);
xor U12120 (N_12120,N_11820,N_11928);
or U12121 (N_12121,N_11869,N_11763);
and U12122 (N_12122,N_11892,N_11887);
and U12123 (N_12123,N_11995,N_11905);
nor U12124 (N_12124,N_11883,N_11853);
nor U12125 (N_12125,N_11876,N_11891);
nand U12126 (N_12126,N_11881,N_11786);
xnor U12127 (N_12127,N_11849,N_11922);
and U12128 (N_12128,N_11938,N_11825);
and U12129 (N_12129,N_11790,N_11932);
nand U12130 (N_12130,N_11949,N_11811);
nor U12131 (N_12131,N_11925,N_11983);
nor U12132 (N_12132,N_11888,N_11982);
xnor U12133 (N_12133,N_11753,N_11889);
xor U12134 (N_12134,N_11961,N_11840);
nand U12135 (N_12135,N_11967,N_11991);
xor U12136 (N_12136,N_11762,N_11886);
nand U12137 (N_12137,N_11813,N_11773);
nand U12138 (N_12138,N_11885,N_11974);
or U12139 (N_12139,N_11789,N_11785);
nor U12140 (N_12140,N_11810,N_11836);
or U12141 (N_12141,N_11928,N_11983);
nand U12142 (N_12142,N_11832,N_11773);
and U12143 (N_12143,N_11984,N_11838);
xnor U12144 (N_12144,N_11932,N_11951);
xor U12145 (N_12145,N_11849,N_11907);
and U12146 (N_12146,N_11785,N_11915);
and U12147 (N_12147,N_11896,N_11795);
and U12148 (N_12148,N_11806,N_11833);
nor U12149 (N_12149,N_11921,N_11938);
nand U12150 (N_12150,N_11763,N_11837);
or U12151 (N_12151,N_11897,N_11965);
or U12152 (N_12152,N_11953,N_11832);
nor U12153 (N_12153,N_11996,N_11842);
and U12154 (N_12154,N_11798,N_11757);
xnor U12155 (N_12155,N_11935,N_11817);
nand U12156 (N_12156,N_11886,N_11957);
nor U12157 (N_12157,N_11752,N_11893);
or U12158 (N_12158,N_11987,N_11992);
or U12159 (N_12159,N_11958,N_11999);
xor U12160 (N_12160,N_11927,N_11918);
or U12161 (N_12161,N_11911,N_11963);
or U12162 (N_12162,N_11867,N_11863);
nor U12163 (N_12163,N_11939,N_11831);
xnor U12164 (N_12164,N_11798,N_11781);
or U12165 (N_12165,N_11908,N_11757);
and U12166 (N_12166,N_11838,N_11812);
nand U12167 (N_12167,N_11782,N_11977);
or U12168 (N_12168,N_11785,N_11866);
nand U12169 (N_12169,N_11828,N_11853);
or U12170 (N_12170,N_11912,N_11994);
or U12171 (N_12171,N_11917,N_11999);
nor U12172 (N_12172,N_11861,N_11912);
or U12173 (N_12173,N_11970,N_11861);
or U12174 (N_12174,N_11751,N_11790);
or U12175 (N_12175,N_11962,N_11821);
nand U12176 (N_12176,N_11811,N_11765);
and U12177 (N_12177,N_11965,N_11917);
nor U12178 (N_12178,N_11859,N_11915);
nor U12179 (N_12179,N_11884,N_11882);
nand U12180 (N_12180,N_11894,N_11804);
or U12181 (N_12181,N_11964,N_11938);
xor U12182 (N_12182,N_11935,N_11867);
xnor U12183 (N_12183,N_11951,N_11900);
nor U12184 (N_12184,N_11800,N_11755);
nor U12185 (N_12185,N_11811,N_11896);
or U12186 (N_12186,N_11770,N_11988);
or U12187 (N_12187,N_11780,N_11929);
and U12188 (N_12188,N_11842,N_11908);
or U12189 (N_12189,N_11920,N_11829);
xor U12190 (N_12190,N_11769,N_11862);
and U12191 (N_12191,N_11817,N_11762);
nor U12192 (N_12192,N_11978,N_11923);
xnor U12193 (N_12193,N_11892,N_11977);
or U12194 (N_12194,N_11835,N_11804);
or U12195 (N_12195,N_11935,N_11963);
nand U12196 (N_12196,N_11811,N_11802);
nand U12197 (N_12197,N_11880,N_11903);
nor U12198 (N_12198,N_11794,N_11936);
and U12199 (N_12199,N_11864,N_11844);
nand U12200 (N_12200,N_11978,N_11908);
or U12201 (N_12201,N_11805,N_11964);
or U12202 (N_12202,N_11903,N_11949);
xnor U12203 (N_12203,N_11958,N_11895);
or U12204 (N_12204,N_11894,N_11995);
nand U12205 (N_12205,N_11791,N_11925);
nor U12206 (N_12206,N_11803,N_11981);
xor U12207 (N_12207,N_11861,N_11924);
nand U12208 (N_12208,N_11898,N_11939);
nor U12209 (N_12209,N_11975,N_11793);
xor U12210 (N_12210,N_11847,N_11809);
nand U12211 (N_12211,N_11876,N_11819);
xor U12212 (N_12212,N_11976,N_11871);
xnor U12213 (N_12213,N_11765,N_11849);
xnor U12214 (N_12214,N_11761,N_11937);
xnor U12215 (N_12215,N_11859,N_11949);
or U12216 (N_12216,N_11848,N_11936);
nor U12217 (N_12217,N_11774,N_11881);
nor U12218 (N_12218,N_11907,N_11929);
or U12219 (N_12219,N_11934,N_11807);
nor U12220 (N_12220,N_11781,N_11978);
or U12221 (N_12221,N_11941,N_11986);
nor U12222 (N_12222,N_11974,N_11955);
xnor U12223 (N_12223,N_11932,N_11833);
and U12224 (N_12224,N_11802,N_11856);
xnor U12225 (N_12225,N_11883,N_11932);
xnor U12226 (N_12226,N_11774,N_11799);
nor U12227 (N_12227,N_11957,N_11899);
and U12228 (N_12228,N_11773,N_11892);
and U12229 (N_12229,N_11945,N_11893);
or U12230 (N_12230,N_11932,N_11888);
and U12231 (N_12231,N_11865,N_11920);
or U12232 (N_12232,N_11791,N_11920);
or U12233 (N_12233,N_11855,N_11858);
nand U12234 (N_12234,N_11969,N_11838);
xnor U12235 (N_12235,N_11859,N_11952);
or U12236 (N_12236,N_11912,N_11849);
xnor U12237 (N_12237,N_11950,N_11968);
nand U12238 (N_12238,N_11846,N_11976);
and U12239 (N_12239,N_11888,N_11894);
xor U12240 (N_12240,N_11782,N_11889);
nor U12241 (N_12241,N_11758,N_11901);
or U12242 (N_12242,N_11843,N_11815);
xnor U12243 (N_12243,N_11939,N_11813);
and U12244 (N_12244,N_11943,N_11869);
nand U12245 (N_12245,N_11910,N_11891);
nand U12246 (N_12246,N_11809,N_11878);
nand U12247 (N_12247,N_11782,N_11823);
nand U12248 (N_12248,N_11759,N_11810);
or U12249 (N_12249,N_11953,N_11919);
xnor U12250 (N_12250,N_12181,N_12213);
and U12251 (N_12251,N_12003,N_12145);
or U12252 (N_12252,N_12004,N_12130);
xor U12253 (N_12253,N_12067,N_12140);
and U12254 (N_12254,N_12209,N_12185);
nand U12255 (N_12255,N_12195,N_12034);
or U12256 (N_12256,N_12191,N_12187);
nor U12257 (N_12257,N_12246,N_12066);
xor U12258 (N_12258,N_12126,N_12135);
nand U12259 (N_12259,N_12098,N_12042);
and U12260 (N_12260,N_12232,N_12089);
or U12261 (N_12261,N_12204,N_12163);
or U12262 (N_12262,N_12044,N_12026);
or U12263 (N_12263,N_12104,N_12106);
and U12264 (N_12264,N_12116,N_12202);
xnor U12265 (N_12265,N_12031,N_12219);
xnor U12266 (N_12266,N_12162,N_12223);
nor U12267 (N_12267,N_12028,N_12109);
xor U12268 (N_12268,N_12080,N_12012);
and U12269 (N_12269,N_12088,N_12176);
nand U12270 (N_12270,N_12009,N_12069);
nor U12271 (N_12271,N_12236,N_12240);
nand U12272 (N_12272,N_12074,N_12085);
and U12273 (N_12273,N_12148,N_12239);
or U12274 (N_12274,N_12041,N_12039);
nor U12275 (N_12275,N_12090,N_12238);
nor U12276 (N_12276,N_12179,N_12072);
xnor U12277 (N_12277,N_12171,N_12128);
xor U12278 (N_12278,N_12220,N_12013);
xnor U12279 (N_12279,N_12062,N_12097);
and U12280 (N_12280,N_12065,N_12131);
xnor U12281 (N_12281,N_12092,N_12078);
or U12282 (N_12282,N_12211,N_12083);
or U12283 (N_12283,N_12235,N_12134);
nand U12284 (N_12284,N_12226,N_12188);
nor U12285 (N_12285,N_12010,N_12054);
and U12286 (N_12286,N_12076,N_12112);
nor U12287 (N_12287,N_12198,N_12111);
and U12288 (N_12288,N_12032,N_12049);
and U12289 (N_12289,N_12151,N_12170);
or U12290 (N_12290,N_12186,N_12201);
xor U12291 (N_12291,N_12189,N_12047);
nand U12292 (N_12292,N_12053,N_12021);
nor U12293 (N_12293,N_12190,N_12212);
nor U12294 (N_12294,N_12160,N_12007);
and U12295 (N_12295,N_12124,N_12183);
xnor U12296 (N_12296,N_12167,N_12114);
and U12297 (N_12297,N_12046,N_12052);
xor U12298 (N_12298,N_12045,N_12147);
and U12299 (N_12299,N_12203,N_12159);
xor U12300 (N_12300,N_12113,N_12022);
nand U12301 (N_12301,N_12018,N_12178);
nor U12302 (N_12302,N_12118,N_12197);
xnor U12303 (N_12303,N_12117,N_12155);
and U12304 (N_12304,N_12180,N_12081);
nor U12305 (N_12305,N_12165,N_12144);
and U12306 (N_12306,N_12127,N_12023);
nor U12307 (N_12307,N_12218,N_12000);
or U12308 (N_12308,N_12017,N_12196);
nand U12309 (N_12309,N_12115,N_12107);
nand U12310 (N_12310,N_12184,N_12095);
xor U12311 (N_12311,N_12227,N_12174);
or U12312 (N_12312,N_12156,N_12101);
and U12313 (N_12313,N_12057,N_12099);
and U12314 (N_12314,N_12093,N_12030);
nor U12315 (N_12315,N_12139,N_12241);
or U12316 (N_12316,N_12002,N_12175);
nor U12317 (N_12317,N_12122,N_12207);
nor U12318 (N_12318,N_12172,N_12234);
nand U12319 (N_12319,N_12233,N_12216);
nand U12320 (N_12320,N_12094,N_12150);
nand U12321 (N_12321,N_12105,N_12051);
xnor U12322 (N_12322,N_12091,N_12169);
nor U12323 (N_12323,N_12079,N_12217);
xor U12324 (N_12324,N_12068,N_12225);
nor U12325 (N_12325,N_12016,N_12006);
nor U12326 (N_12326,N_12152,N_12164);
or U12327 (N_12327,N_12177,N_12027);
and U12328 (N_12328,N_12020,N_12073);
and U12329 (N_12329,N_12029,N_12025);
nand U12330 (N_12330,N_12103,N_12230);
nand U12331 (N_12331,N_12214,N_12096);
nor U12332 (N_12332,N_12129,N_12108);
and U12333 (N_12333,N_12064,N_12193);
and U12334 (N_12334,N_12200,N_12199);
nand U12335 (N_12335,N_12100,N_12245);
and U12336 (N_12336,N_12137,N_12149);
nor U12337 (N_12337,N_12194,N_12157);
nand U12338 (N_12338,N_12014,N_12206);
xor U12339 (N_12339,N_12132,N_12119);
nor U12340 (N_12340,N_12229,N_12120);
or U12341 (N_12341,N_12125,N_12055);
or U12342 (N_12342,N_12138,N_12048);
and U12343 (N_12343,N_12221,N_12102);
and U12344 (N_12344,N_12075,N_12036);
or U12345 (N_12345,N_12024,N_12154);
and U12346 (N_12346,N_12237,N_12244);
nor U12347 (N_12347,N_12033,N_12243);
and U12348 (N_12348,N_12146,N_12224);
nand U12349 (N_12349,N_12192,N_12222);
nor U12350 (N_12350,N_12038,N_12037);
and U12351 (N_12351,N_12248,N_12208);
nor U12352 (N_12352,N_12158,N_12123);
nor U12353 (N_12353,N_12153,N_12228);
xor U12354 (N_12354,N_12015,N_12070);
or U12355 (N_12355,N_12063,N_12058);
xor U12356 (N_12356,N_12242,N_12173);
and U12357 (N_12357,N_12143,N_12077);
and U12358 (N_12358,N_12161,N_12136);
nor U12359 (N_12359,N_12168,N_12050);
nand U12360 (N_12360,N_12001,N_12008);
nor U12361 (N_12361,N_12110,N_12082);
nand U12362 (N_12362,N_12059,N_12205);
xnor U12363 (N_12363,N_12056,N_12060);
nor U12364 (N_12364,N_12182,N_12141);
nand U12365 (N_12365,N_12086,N_12133);
and U12366 (N_12366,N_12061,N_12231);
xor U12367 (N_12367,N_12121,N_12210);
nor U12368 (N_12368,N_12035,N_12071);
and U12369 (N_12369,N_12084,N_12019);
xor U12370 (N_12370,N_12005,N_12043);
and U12371 (N_12371,N_12011,N_12142);
nor U12372 (N_12372,N_12166,N_12087);
nor U12373 (N_12373,N_12215,N_12247);
xor U12374 (N_12374,N_12040,N_12249);
nor U12375 (N_12375,N_12177,N_12166);
nor U12376 (N_12376,N_12014,N_12211);
and U12377 (N_12377,N_12204,N_12164);
or U12378 (N_12378,N_12022,N_12087);
or U12379 (N_12379,N_12168,N_12134);
xnor U12380 (N_12380,N_12168,N_12081);
or U12381 (N_12381,N_12073,N_12168);
nor U12382 (N_12382,N_12130,N_12079);
xor U12383 (N_12383,N_12120,N_12207);
nor U12384 (N_12384,N_12105,N_12056);
and U12385 (N_12385,N_12051,N_12007);
or U12386 (N_12386,N_12091,N_12125);
nand U12387 (N_12387,N_12211,N_12019);
xnor U12388 (N_12388,N_12068,N_12166);
or U12389 (N_12389,N_12079,N_12221);
and U12390 (N_12390,N_12025,N_12051);
nand U12391 (N_12391,N_12215,N_12079);
nand U12392 (N_12392,N_12075,N_12110);
or U12393 (N_12393,N_12139,N_12216);
xnor U12394 (N_12394,N_12100,N_12012);
nand U12395 (N_12395,N_12061,N_12032);
or U12396 (N_12396,N_12172,N_12090);
nor U12397 (N_12397,N_12063,N_12038);
xor U12398 (N_12398,N_12116,N_12122);
and U12399 (N_12399,N_12204,N_12144);
nand U12400 (N_12400,N_12126,N_12238);
or U12401 (N_12401,N_12024,N_12192);
nand U12402 (N_12402,N_12046,N_12173);
nor U12403 (N_12403,N_12079,N_12125);
nand U12404 (N_12404,N_12082,N_12117);
or U12405 (N_12405,N_12212,N_12145);
and U12406 (N_12406,N_12025,N_12091);
xor U12407 (N_12407,N_12144,N_12058);
nor U12408 (N_12408,N_12038,N_12072);
or U12409 (N_12409,N_12219,N_12126);
nor U12410 (N_12410,N_12238,N_12004);
or U12411 (N_12411,N_12164,N_12120);
or U12412 (N_12412,N_12188,N_12156);
nand U12413 (N_12413,N_12249,N_12075);
xor U12414 (N_12414,N_12072,N_12093);
nand U12415 (N_12415,N_12190,N_12013);
nor U12416 (N_12416,N_12030,N_12218);
and U12417 (N_12417,N_12120,N_12069);
nor U12418 (N_12418,N_12135,N_12168);
xnor U12419 (N_12419,N_12172,N_12032);
nand U12420 (N_12420,N_12125,N_12059);
xnor U12421 (N_12421,N_12187,N_12021);
and U12422 (N_12422,N_12151,N_12021);
nor U12423 (N_12423,N_12160,N_12214);
nor U12424 (N_12424,N_12134,N_12187);
xor U12425 (N_12425,N_12245,N_12153);
or U12426 (N_12426,N_12140,N_12178);
nand U12427 (N_12427,N_12128,N_12232);
nand U12428 (N_12428,N_12133,N_12176);
xnor U12429 (N_12429,N_12088,N_12059);
nand U12430 (N_12430,N_12022,N_12238);
or U12431 (N_12431,N_12135,N_12136);
nand U12432 (N_12432,N_12232,N_12217);
nor U12433 (N_12433,N_12140,N_12119);
xnor U12434 (N_12434,N_12193,N_12063);
xnor U12435 (N_12435,N_12004,N_12075);
or U12436 (N_12436,N_12210,N_12079);
xnor U12437 (N_12437,N_12077,N_12099);
nand U12438 (N_12438,N_12002,N_12005);
and U12439 (N_12439,N_12137,N_12135);
and U12440 (N_12440,N_12236,N_12156);
nand U12441 (N_12441,N_12042,N_12004);
or U12442 (N_12442,N_12136,N_12149);
nor U12443 (N_12443,N_12247,N_12031);
and U12444 (N_12444,N_12079,N_12050);
or U12445 (N_12445,N_12046,N_12032);
nand U12446 (N_12446,N_12204,N_12090);
xnor U12447 (N_12447,N_12200,N_12186);
xnor U12448 (N_12448,N_12237,N_12226);
nor U12449 (N_12449,N_12088,N_12146);
xor U12450 (N_12450,N_12104,N_12078);
and U12451 (N_12451,N_12245,N_12146);
xnor U12452 (N_12452,N_12246,N_12138);
nand U12453 (N_12453,N_12213,N_12039);
xor U12454 (N_12454,N_12248,N_12070);
nand U12455 (N_12455,N_12153,N_12146);
and U12456 (N_12456,N_12048,N_12080);
nor U12457 (N_12457,N_12060,N_12176);
and U12458 (N_12458,N_12000,N_12088);
nor U12459 (N_12459,N_12006,N_12138);
and U12460 (N_12460,N_12017,N_12013);
or U12461 (N_12461,N_12071,N_12205);
nor U12462 (N_12462,N_12115,N_12110);
nor U12463 (N_12463,N_12007,N_12150);
or U12464 (N_12464,N_12031,N_12063);
nor U12465 (N_12465,N_12041,N_12159);
and U12466 (N_12466,N_12130,N_12048);
or U12467 (N_12467,N_12067,N_12137);
nand U12468 (N_12468,N_12092,N_12169);
and U12469 (N_12469,N_12216,N_12173);
or U12470 (N_12470,N_12019,N_12244);
nor U12471 (N_12471,N_12046,N_12043);
and U12472 (N_12472,N_12183,N_12011);
nand U12473 (N_12473,N_12108,N_12118);
nor U12474 (N_12474,N_12100,N_12196);
xnor U12475 (N_12475,N_12112,N_12053);
nor U12476 (N_12476,N_12004,N_12132);
nor U12477 (N_12477,N_12132,N_12071);
nand U12478 (N_12478,N_12062,N_12125);
nor U12479 (N_12479,N_12066,N_12069);
nand U12480 (N_12480,N_12196,N_12134);
xnor U12481 (N_12481,N_12066,N_12106);
nand U12482 (N_12482,N_12178,N_12047);
or U12483 (N_12483,N_12229,N_12053);
or U12484 (N_12484,N_12181,N_12228);
xor U12485 (N_12485,N_12090,N_12069);
or U12486 (N_12486,N_12067,N_12216);
xor U12487 (N_12487,N_12094,N_12011);
or U12488 (N_12488,N_12229,N_12223);
nand U12489 (N_12489,N_12188,N_12209);
nand U12490 (N_12490,N_12112,N_12065);
nand U12491 (N_12491,N_12210,N_12185);
xor U12492 (N_12492,N_12046,N_12191);
nand U12493 (N_12493,N_12123,N_12079);
or U12494 (N_12494,N_12029,N_12016);
or U12495 (N_12495,N_12128,N_12220);
and U12496 (N_12496,N_12131,N_12072);
nand U12497 (N_12497,N_12151,N_12004);
xnor U12498 (N_12498,N_12038,N_12092);
nand U12499 (N_12499,N_12216,N_12181);
nand U12500 (N_12500,N_12422,N_12394);
nor U12501 (N_12501,N_12399,N_12270);
and U12502 (N_12502,N_12352,N_12419);
xor U12503 (N_12503,N_12273,N_12427);
nand U12504 (N_12504,N_12357,N_12483);
and U12505 (N_12505,N_12250,N_12263);
nand U12506 (N_12506,N_12374,N_12449);
xor U12507 (N_12507,N_12356,N_12283);
and U12508 (N_12508,N_12271,N_12319);
and U12509 (N_12509,N_12269,N_12308);
and U12510 (N_12510,N_12292,N_12439);
xor U12511 (N_12511,N_12497,N_12408);
nor U12512 (N_12512,N_12280,N_12454);
xnor U12513 (N_12513,N_12418,N_12462);
nand U12514 (N_12514,N_12295,N_12274);
xnor U12515 (N_12515,N_12383,N_12254);
and U12516 (N_12516,N_12488,N_12404);
or U12517 (N_12517,N_12477,N_12317);
nor U12518 (N_12518,N_12298,N_12407);
nor U12519 (N_12519,N_12337,N_12458);
and U12520 (N_12520,N_12397,N_12370);
or U12521 (N_12521,N_12387,N_12428);
nand U12522 (N_12522,N_12431,N_12421);
or U12523 (N_12523,N_12380,N_12349);
and U12524 (N_12524,N_12359,N_12345);
and U12525 (N_12525,N_12293,N_12262);
nor U12526 (N_12526,N_12360,N_12276);
nor U12527 (N_12527,N_12331,N_12266);
nor U12528 (N_12528,N_12253,N_12303);
xnor U12529 (N_12529,N_12368,N_12480);
nand U12530 (N_12530,N_12320,N_12289);
nand U12531 (N_12531,N_12414,N_12347);
xor U12532 (N_12532,N_12464,N_12410);
and U12533 (N_12533,N_12491,N_12259);
or U12534 (N_12534,N_12378,N_12469);
and U12535 (N_12535,N_12287,N_12300);
and U12536 (N_12536,N_12382,N_12297);
nor U12537 (N_12537,N_12369,N_12455);
nor U12538 (N_12538,N_12323,N_12470);
or U12539 (N_12539,N_12321,N_12342);
and U12540 (N_12540,N_12318,N_12492);
and U12541 (N_12541,N_12456,N_12351);
and U12542 (N_12542,N_12487,N_12395);
or U12543 (N_12543,N_12364,N_12485);
and U12544 (N_12544,N_12405,N_12344);
nor U12545 (N_12545,N_12481,N_12251);
and U12546 (N_12546,N_12437,N_12446);
or U12547 (N_12547,N_12332,N_12438);
nor U12548 (N_12548,N_12371,N_12328);
xnor U12549 (N_12549,N_12499,N_12482);
xor U12550 (N_12550,N_12416,N_12329);
nand U12551 (N_12551,N_12343,N_12420);
xnor U12552 (N_12552,N_12339,N_12463);
nand U12553 (N_12553,N_12392,N_12363);
and U12554 (N_12554,N_12435,N_12257);
nor U12555 (N_12555,N_12355,N_12286);
nor U12556 (N_12556,N_12285,N_12460);
or U12557 (N_12557,N_12372,N_12284);
xnor U12558 (N_12558,N_12411,N_12278);
nor U12559 (N_12559,N_12451,N_12402);
nand U12560 (N_12560,N_12461,N_12376);
nand U12561 (N_12561,N_12288,N_12468);
and U12562 (N_12562,N_12400,N_12275);
nor U12563 (N_12563,N_12450,N_12322);
nand U12564 (N_12564,N_12327,N_12385);
xnor U12565 (N_12565,N_12401,N_12417);
nor U12566 (N_12566,N_12358,N_12442);
nor U12567 (N_12567,N_12433,N_12265);
and U12568 (N_12568,N_12479,N_12453);
nand U12569 (N_12569,N_12334,N_12466);
nand U12570 (N_12570,N_12436,N_12443);
and U12571 (N_12571,N_12472,N_12448);
nor U12572 (N_12572,N_12389,N_12471);
or U12573 (N_12573,N_12361,N_12350);
xor U12574 (N_12574,N_12252,N_12498);
and U12575 (N_12575,N_12445,N_12313);
nor U12576 (N_12576,N_12365,N_12432);
or U12577 (N_12577,N_12326,N_12452);
xor U12578 (N_12578,N_12425,N_12473);
nand U12579 (N_12579,N_12496,N_12377);
or U12580 (N_12580,N_12316,N_12441);
nor U12581 (N_12581,N_12346,N_12388);
and U12582 (N_12582,N_12306,N_12447);
or U12583 (N_12583,N_12391,N_12340);
and U12584 (N_12584,N_12494,N_12362);
or U12585 (N_12585,N_12426,N_12281);
xor U12586 (N_12586,N_12366,N_12296);
or U12587 (N_12587,N_12413,N_12490);
nand U12588 (N_12588,N_12475,N_12353);
nor U12589 (N_12589,N_12393,N_12379);
and U12590 (N_12590,N_12272,N_12384);
and U12591 (N_12591,N_12336,N_12282);
xor U12592 (N_12592,N_12302,N_12294);
or U12593 (N_12593,N_12310,N_12434);
xnor U12594 (N_12594,N_12312,N_12324);
nand U12595 (N_12595,N_12301,N_12495);
nand U12596 (N_12596,N_12335,N_12423);
or U12597 (N_12597,N_12381,N_12467);
and U12598 (N_12598,N_12279,N_12406);
nor U12599 (N_12599,N_12315,N_12291);
nand U12600 (N_12600,N_12264,N_12489);
nand U12601 (N_12601,N_12299,N_12429);
xnor U12602 (N_12602,N_12354,N_12373);
nor U12603 (N_12603,N_12268,N_12255);
nor U12604 (N_12604,N_12403,N_12261);
nand U12605 (N_12605,N_12256,N_12486);
or U12606 (N_12606,N_12398,N_12277);
xnor U12607 (N_12607,N_12396,N_12290);
or U12608 (N_12608,N_12307,N_12260);
xnor U12609 (N_12609,N_12440,N_12338);
nand U12610 (N_12610,N_12386,N_12412);
or U12611 (N_12611,N_12258,N_12430);
xnor U12612 (N_12612,N_12304,N_12390);
xor U12613 (N_12613,N_12465,N_12333);
or U12614 (N_12614,N_12309,N_12415);
and U12615 (N_12615,N_12330,N_12311);
and U12616 (N_12616,N_12367,N_12267);
nand U12617 (N_12617,N_12478,N_12341);
nand U12618 (N_12618,N_12457,N_12409);
xnor U12619 (N_12619,N_12325,N_12375);
or U12620 (N_12620,N_12476,N_12493);
nand U12621 (N_12621,N_12348,N_12474);
and U12622 (N_12622,N_12444,N_12424);
xor U12623 (N_12623,N_12484,N_12314);
nor U12624 (N_12624,N_12459,N_12305);
nor U12625 (N_12625,N_12264,N_12393);
or U12626 (N_12626,N_12397,N_12469);
and U12627 (N_12627,N_12276,N_12311);
or U12628 (N_12628,N_12455,N_12356);
nand U12629 (N_12629,N_12297,N_12498);
or U12630 (N_12630,N_12310,N_12382);
xor U12631 (N_12631,N_12433,N_12422);
xor U12632 (N_12632,N_12296,N_12283);
nor U12633 (N_12633,N_12438,N_12431);
nor U12634 (N_12634,N_12479,N_12345);
xor U12635 (N_12635,N_12351,N_12288);
and U12636 (N_12636,N_12466,N_12430);
nor U12637 (N_12637,N_12469,N_12260);
nor U12638 (N_12638,N_12453,N_12412);
or U12639 (N_12639,N_12496,N_12439);
nor U12640 (N_12640,N_12358,N_12365);
xor U12641 (N_12641,N_12315,N_12346);
nand U12642 (N_12642,N_12353,N_12268);
xnor U12643 (N_12643,N_12483,N_12275);
and U12644 (N_12644,N_12271,N_12312);
and U12645 (N_12645,N_12333,N_12471);
or U12646 (N_12646,N_12279,N_12402);
and U12647 (N_12647,N_12487,N_12481);
nor U12648 (N_12648,N_12266,N_12395);
xor U12649 (N_12649,N_12495,N_12390);
nor U12650 (N_12650,N_12487,N_12471);
xor U12651 (N_12651,N_12458,N_12370);
and U12652 (N_12652,N_12403,N_12446);
nor U12653 (N_12653,N_12365,N_12385);
and U12654 (N_12654,N_12381,N_12460);
nand U12655 (N_12655,N_12340,N_12387);
xnor U12656 (N_12656,N_12388,N_12351);
and U12657 (N_12657,N_12385,N_12469);
xnor U12658 (N_12658,N_12297,N_12411);
nor U12659 (N_12659,N_12282,N_12497);
nor U12660 (N_12660,N_12255,N_12442);
nor U12661 (N_12661,N_12383,N_12380);
nand U12662 (N_12662,N_12416,N_12335);
nand U12663 (N_12663,N_12420,N_12384);
nor U12664 (N_12664,N_12470,N_12398);
and U12665 (N_12665,N_12420,N_12451);
xor U12666 (N_12666,N_12462,N_12333);
and U12667 (N_12667,N_12307,N_12336);
xnor U12668 (N_12668,N_12498,N_12332);
and U12669 (N_12669,N_12302,N_12317);
or U12670 (N_12670,N_12386,N_12370);
nor U12671 (N_12671,N_12324,N_12487);
xor U12672 (N_12672,N_12393,N_12333);
nor U12673 (N_12673,N_12280,N_12473);
or U12674 (N_12674,N_12287,N_12367);
or U12675 (N_12675,N_12452,N_12273);
or U12676 (N_12676,N_12336,N_12300);
nor U12677 (N_12677,N_12471,N_12266);
nor U12678 (N_12678,N_12387,N_12468);
nand U12679 (N_12679,N_12362,N_12411);
and U12680 (N_12680,N_12443,N_12430);
and U12681 (N_12681,N_12288,N_12441);
or U12682 (N_12682,N_12374,N_12336);
or U12683 (N_12683,N_12346,N_12484);
nand U12684 (N_12684,N_12460,N_12351);
nand U12685 (N_12685,N_12465,N_12327);
nand U12686 (N_12686,N_12462,N_12448);
or U12687 (N_12687,N_12442,N_12253);
nand U12688 (N_12688,N_12452,N_12292);
or U12689 (N_12689,N_12429,N_12353);
nand U12690 (N_12690,N_12313,N_12431);
xnor U12691 (N_12691,N_12285,N_12296);
and U12692 (N_12692,N_12347,N_12296);
or U12693 (N_12693,N_12254,N_12349);
and U12694 (N_12694,N_12480,N_12383);
nor U12695 (N_12695,N_12277,N_12409);
xnor U12696 (N_12696,N_12289,N_12382);
xnor U12697 (N_12697,N_12453,N_12365);
or U12698 (N_12698,N_12407,N_12284);
or U12699 (N_12699,N_12280,N_12403);
nand U12700 (N_12700,N_12495,N_12384);
or U12701 (N_12701,N_12424,N_12277);
or U12702 (N_12702,N_12415,N_12318);
nor U12703 (N_12703,N_12346,N_12262);
nand U12704 (N_12704,N_12314,N_12320);
nor U12705 (N_12705,N_12261,N_12300);
or U12706 (N_12706,N_12371,N_12357);
xnor U12707 (N_12707,N_12256,N_12478);
or U12708 (N_12708,N_12279,N_12360);
nand U12709 (N_12709,N_12324,N_12430);
nor U12710 (N_12710,N_12458,N_12450);
or U12711 (N_12711,N_12406,N_12405);
xor U12712 (N_12712,N_12250,N_12379);
xor U12713 (N_12713,N_12374,N_12342);
or U12714 (N_12714,N_12331,N_12329);
nand U12715 (N_12715,N_12327,N_12473);
xnor U12716 (N_12716,N_12384,N_12446);
or U12717 (N_12717,N_12394,N_12378);
nand U12718 (N_12718,N_12416,N_12284);
or U12719 (N_12719,N_12435,N_12254);
nand U12720 (N_12720,N_12337,N_12269);
and U12721 (N_12721,N_12355,N_12296);
or U12722 (N_12722,N_12281,N_12461);
or U12723 (N_12723,N_12361,N_12445);
nand U12724 (N_12724,N_12472,N_12383);
nor U12725 (N_12725,N_12337,N_12345);
nand U12726 (N_12726,N_12417,N_12330);
nand U12727 (N_12727,N_12265,N_12480);
nand U12728 (N_12728,N_12331,N_12254);
nand U12729 (N_12729,N_12274,N_12422);
and U12730 (N_12730,N_12495,N_12483);
nand U12731 (N_12731,N_12401,N_12294);
xnor U12732 (N_12732,N_12456,N_12459);
nor U12733 (N_12733,N_12485,N_12438);
nand U12734 (N_12734,N_12251,N_12346);
xor U12735 (N_12735,N_12252,N_12481);
or U12736 (N_12736,N_12379,N_12461);
nor U12737 (N_12737,N_12410,N_12393);
xor U12738 (N_12738,N_12388,N_12464);
xor U12739 (N_12739,N_12348,N_12397);
xnor U12740 (N_12740,N_12365,N_12399);
and U12741 (N_12741,N_12286,N_12368);
or U12742 (N_12742,N_12386,N_12266);
nand U12743 (N_12743,N_12401,N_12467);
and U12744 (N_12744,N_12326,N_12498);
xor U12745 (N_12745,N_12281,N_12430);
and U12746 (N_12746,N_12336,N_12455);
xor U12747 (N_12747,N_12449,N_12455);
or U12748 (N_12748,N_12251,N_12297);
xor U12749 (N_12749,N_12349,N_12297);
and U12750 (N_12750,N_12588,N_12689);
xnor U12751 (N_12751,N_12729,N_12611);
or U12752 (N_12752,N_12514,N_12549);
nand U12753 (N_12753,N_12667,N_12688);
nor U12754 (N_12754,N_12746,N_12748);
and U12755 (N_12755,N_12584,N_12663);
nor U12756 (N_12756,N_12525,N_12593);
xor U12757 (N_12757,N_12636,N_12642);
nand U12758 (N_12758,N_12724,N_12595);
or U12759 (N_12759,N_12618,N_12693);
and U12760 (N_12760,N_12606,N_12605);
nand U12761 (N_12761,N_12578,N_12603);
xor U12762 (N_12762,N_12696,N_12576);
and U12763 (N_12763,N_12651,N_12616);
nand U12764 (N_12764,N_12705,N_12528);
or U12765 (N_12765,N_12726,N_12562);
xnor U12766 (N_12766,N_12556,N_12675);
and U12767 (N_12767,N_12735,N_12677);
nand U12768 (N_12768,N_12736,N_12712);
xor U12769 (N_12769,N_12512,N_12644);
and U12770 (N_12770,N_12742,N_12659);
or U12771 (N_12771,N_12565,N_12639);
xor U12772 (N_12772,N_12568,N_12747);
nand U12773 (N_12773,N_12586,N_12721);
and U12774 (N_12774,N_12733,N_12569);
and U12775 (N_12775,N_12602,N_12710);
xor U12776 (N_12776,N_12701,N_12722);
nand U12777 (N_12777,N_12685,N_12535);
or U12778 (N_12778,N_12661,N_12725);
nand U12779 (N_12779,N_12730,N_12620);
xnor U12780 (N_12780,N_12637,N_12655);
nor U12781 (N_12781,N_12518,N_12681);
xor U12782 (N_12782,N_12632,N_12600);
or U12783 (N_12783,N_12613,N_12662);
nor U12784 (N_12784,N_12543,N_12654);
and U12785 (N_12785,N_12591,N_12541);
or U12786 (N_12786,N_12676,N_12523);
or U12787 (N_12787,N_12704,N_12657);
nor U12788 (N_12788,N_12634,N_12739);
nor U12789 (N_12789,N_12660,N_12646);
or U12790 (N_12790,N_12652,N_12515);
and U12791 (N_12791,N_12694,N_12537);
or U12792 (N_12792,N_12577,N_12695);
and U12793 (N_12793,N_12647,N_12626);
xnor U12794 (N_12794,N_12732,N_12737);
nand U12795 (N_12795,N_12589,N_12633);
nand U12796 (N_12796,N_12524,N_12590);
xor U12797 (N_12797,N_12686,N_12740);
or U12798 (N_12798,N_12629,N_12575);
or U12799 (N_12799,N_12580,N_12691);
nand U12800 (N_12800,N_12554,N_12604);
or U12801 (N_12801,N_12664,N_12506);
nand U12802 (N_12802,N_12560,N_12617);
and U12803 (N_12803,N_12643,N_12674);
or U12804 (N_12804,N_12571,N_12526);
xor U12805 (N_12805,N_12731,N_12513);
xnor U12806 (N_12806,N_12745,N_12621);
or U12807 (N_12807,N_12703,N_12517);
nand U12808 (N_12808,N_12608,N_12738);
nor U12809 (N_12809,N_12719,N_12542);
nor U12810 (N_12810,N_12545,N_12572);
nor U12811 (N_12811,N_12532,N_12550);
or U12812 (N_12812,N_12711,N_12610);
nor U12813 (N_12813,N_12708,N_12682);
and U12814 (N_12814,N_12607,N_12640);
or U12815 (N_12815,N_12698,N_12546);
and U12816 (N_12816,N_12509,N_12628);
or U12817 (N_12817,N_12743,N_12507);
nor U12818 (N_12818,N_12744,N_12706);
xnor U12819 (N_12819,N_12622,N_12510);
xnor U12820 (N_12820,N_12692,N_12717);
or U12821 (N_12821,N_12716,N_12631);
xor U12822 (N_12822,N_12531,N_12563);
xnor U12823 (N_12823,N_12653,N_12650);
nand U12824 (N_12824,N_12723,N_12601);
nand U12825 (N_12825,N_12683,N_12567);
nor U12826 (N_12826,N_12552,N_12511);
and U12827 (N_12827,N_12530,N_12641);
or U12828 (N_12828,N_12624,N_12579);
nor U12829 (N_12829,N_12638,N_12714);
nand U12830 (N_12830,N_12697,N_12627);
xor U12831 (N_12831,N_12665,N_12713);
nand U12832 (N_12832,N_12671,N_12678);
or U12833 (N_12833,N_12709,N_12533);
or U12834 (N_12834,N_12645,N_12702);
or U12835 (N_12835,N_12566,N_12548);
nand U12836 (N_12836,N_12596,N_12669);
and U12837 (N_12837,N_12503,N_12551);
and U12838 (N_12838,N_12547,N_12558);
nand U12839 (N_12839,N_12553,N_12619);
nand U12840 (N_12840,N_12504,N_12672);
or U12841 (N_12841,N_12544,N_12540);
nand U12842 (N_12842,N_12522,N_12728);
nor U12843 (N_12843,N_12700,N_12707);
nor U12844 (N_12844,N_12699,N_12559);
or U12845 (N_12845,N_12573,N_12516);
and U12846 (N_12846,N_12670,N_12582);
nor U12847 (N_12847,N_12527,N_12727);
or U12848 (N_12848,N_12720,N_12649);
and U12849 (N_12849,N_12684,N_12521);
and U12850 (N_12850,N_12555,N_12564);
xor U12851 (N_12851,N_12680,N_12718);
nand U12852 (N_12852,N_12598,N_12557);
or U12853 (N_12853,N_12500,N_12570);
nand U12854 (N_12854,N_12561,N_12520);
nand U12855 (N_12855,N_12538,N_12625);
and U12856 (N_12856,N_12581,N_12574);
xor U12857 (N_12857,N_12508,N_12539);
and U12858 (N_12858,N_12648,N_12666);
nor U12859 (N_12859,N_12635,N_12583);
and U12860 (N_12860,N_12609,N_12749);
nand U12861 (N_12861,N_12592,N_12679);
xnor U12862 (N_12862,N_12587,N_12715);
nand U12863 (N_12863,N_12599,N_12594);
xnor U12864 (N_12864,N_12687,N_12630);
and U12865 (N_12865,N_12534,N_12668);
nor U12866 (N_12866,N_12536,N_12623);
xor U12867 (N_12867,N_12673,N_12615);
or U12868 (N_12868,N_12519,N_12585);
and U12869 (N_12869,N_12529,N_12656);
nor U12870 (N_12870,N_12734,N_12505);
and U12871 (N_12871,N_12502,N_12741);
and U12872 (N_12872,N_12501,N_12612);
xnor U12873 (N_12873,N_12658,N_12614);
and U12874 (N_12874,N_12597,N_12690);
and U12875 (N_12875,N_12534,N_12652);
and U12876 (N_12876,N_12621,N_12503);
nor U12877 (N_12877,N_12685,N_12638);
or U12878 (N_12878,N_12521,N_12596);
nor U12879 (N_12879,N_12580,N_12589);
and U12880 (N_12880,N_12602,N_12595);
or U12881 (N_12881,N_12602,N_12611);
xor U12882 (N_12882,N_12695,N_12652);
and U12883 (N_12883,N_12605,N_12537);
or U12884 (N_12884,N_12689,N_12512);
xnor U12885 (N_12885,N_12601,N_12543);
or U12886 (N_12886,N_12749,N_12679);
nand U12887 (N_12887,N_12575,N_12539);
or U12888 (N_12888,N_12538,N_12544);
and U12889 (N_12889,N_12647,N_12639);
and U12890 (N_12890,N_12669,N_12580);
nor U12891 (N_12891,N_12591,N_12636);
or U12892 (N_12892,N_12553,N_12716);
nand U12893 (N_12893,N_12532,N_12677);
nand U12894 (N_12894,N_12618,N_12554);
nand U12895 (N_12895,N_12692,N_12504);
or U12896 (N_12896,N_12730,N_12725);
xor U12897 (N_12897,N_12680,N_12727);
nor U12898 (N_12898,N_12717,N_12652);
or U12899 (N_12899,N_12646,N_12636);
nor U12900 (N_12900,N_12514,N_12640);
and U12901 (N_12901,N_12605,N_12698);
and U12902 (N_12902,N_12746,N_12707);
or U12903 (N_12903,N_12612,N_12564);
nor U12904 (N_12904,N_12554,N_12725);
or U12905 (N_12905,N_12712,N_12536);
nand U12906 (N_12906,N_12658,N_12710);
nand U12907 (N_12907,N_12527,N_12637);
or U12908 (N_12908,N_12593,N_12730);
xnor U12909 (N_12909,N_12627,N_12577);
and U12910 (N_12910,N_12716,N_12738);
nand U12911 (N_12911,N_12725,N_12682);
xnor U12912 (N_12912,N_12682,N_12631);
xor U12913 (N_12913,N_12513,N_12577);
and U12914 (N_12914,N_12741,N_12696);
xnor U12915 (N_12915,N_12509,N_12570);
or U12916 (N_12916,N_12537,N_12668);
xor U12917 (N_12917,N_12647,N_12575);
nand U12918 (N_12918,N_12742,N_12520);
and U12919 (N_12919,N_12699,N_12661);
nor U12920 (N_12920,N_12531,N_12513);
or U12921 (N_12921,N_12746,N_12691);
xor U12922 (N_12922,N_12635,N_12670);
nand U12923 (N_12923,N_12516,N_12739);
xnor U12924 (N_12924,N_12513,N_12501);
and U12925 (N_12925,N_12659,N_12627);
nor U12926 (N_12926,N_12577,N_12674);
and U12927 (N_12927,N_12674,N_12654);
nor U12928 (N_12928,N_12639,N_12609);
nor U12929 (N_12929,N_12670,N_12564);
nand U12930 (N_12930,N_12571,N_12661);
xor U12931 (N_12931,N_12500,N_12521);
and U12932 (N_12932,N_12744,N_12697);
nor U12933 (N_12933,N_12535,N_12624);
and U12934 (N_12934,N_12703,N_12694);
or U12935 (N_12935,N_12689,N_12692);
or U12936 (N_12936,N_12575,N_12598);
xnor U12937 (N_12937,N_12596,N_12748);
nor U12938 (N_12938,N_12738,N_12675);
and U12939 (N_12939,N_12571,N_12543);
nand U12940 (N_12940,N_12627,N_12562);
nand U12941 (N_12941,N_12516,N_12671);
or U12942 (N_12942,N_12597,N_12542);
xor U12943 (N_12943,N_12622,N_12683);
or U12944 (N_12944,N_12690,N_12519);
nand U12945 (N_12945,N_12516,N_12638);
or U12946 (N_12946,N_12674,N_12594);
nor U12947 (N_12947,N_12635,N_12534);
and U12948 (N_12948,N_12718,N_12553);
or U12949 (N_12949,N_12552,N_12549);
nor U12950 (N_12950,N_12639,N_12742);
nand U12951 (N_12951,N_12582,N_12674);
xor U12952 (N_12952,N_12571,N_12501);
or U12953 (N_12953,N_12583,N_12686);
nand U12954 (N_12954,N_12664,N_12626);
and U12955 (N_12955,N_12639,N_12614);
and U12956 (N_12956,N_12597,N_12539);
or U12957 (N_12957,N_12682,N_12582);
or U12958 (N_12958,N_12527,N_12592);
nand U12959 (N_12959,N_12562,N_12532);
and U12960 (N_12960,N_12679,N_12738);
or U12961 (N_12961,N_12540,N_12545);
or U12962 (N_12962,N_12560,N_12589);
or U12963 (N_12963,N_12593,N_12733);
nor U12964 (N_12964,N_12691,N_12519);
and U12965 (N_12965,N_12707,N_12649);
xor U12966 (N_12966,N_12563,N_12717);
xor U12967 (N_12967,N_12746,N_12682);
xnor U12968 (N_12968,N_12617,N_12512);
xor U12969 (N_12969,N_12617,N_12564);
nand U12970 (N_12970,N_12556,N_12651);
and U12971 (N_12971,N_12618,N_12580);
and U12972 (N_12972,N_12521,N_12572);
nor U12973 (N_12973,N_12697,N_12724);
and U12974 (N_12974,N_12727,N_12715);
xor U12975 (N_12975,N_12574,N_12544);
or U12976 (N_12976,N_12606,N_12575);
and U12977 (N_12977,N_12658,N_12728);
nand U12978 (N_12978,N_12690,N_12668);
or U12979 (N_12979,N_12549,N_12656);
xor U12980 (N_12980,N_12743,N_12593);
xnor U12981 (N_12981,N_12552,N_12698);
and U12982 (N_12982,N_12611,N_12559);
nor U12983 (N_12983,N_12582,N_12734);
and U12984 (N_12984,N_12642,N_12740);
nor U12985 (N_12985,N_12545,N_12664);
xor U12986 (N_12986,N_12697,N_12643);
and U12987 (N_12987,N_12575,N_12630);
xnor U12988 (N_12988,N_12638,N_12723);
nand U12989 (N_12989,N_12612,N_12560);
and U12990 (N_12990,N_12674,N_12711);
or U12991 (N_12991,N_12525,N_12502);
nand U12992 (N_12992,N_12590,N_12726);
nor U12993 (N_12993,N_12555,N_12573);
nor U12994 (N_12994,N_12566,N_12611);
xor U12995 (N_12995,N_12505,N_12661);
nor U12996 (N_12996,N_12709,N_12532);
or U12997 (N_12997,N_12650,N_12517);
or U12998 (N_12998,N_12553,N_12698);
xnor U12999 (N_12999,N_12558,N_12576);
or U13000 (N_13000,N_12863,N_12911);
xor U13001 (N_13001,N_12909,N_12905);
nand U13002 (N_13002,N_12804,N_12856);
or U13003 (N_13003,N_12954,N_12774);
xnor U13004 (N_13004,N_12893,N_12845);
or U13005 (N_13005,N_12855,N_12925);
xor U13006 (N_13006,N_12884,N_12952);
or U13007 (N_13007,N_12784,N_12978);
xnor U13008 (N_13008,N_12881,N_12797);
and U13009 (N_13009,N_12995,N_12941);
nor U13010 (N_13010,N_12793,N_12839);
and U13011 (N_13011,N_12788,N_12792);
nor U13012 (N_13012,N_12752,N_12838);
nor U13013 (N_13013,N_12986,N_12970);
nor U13014 (N_13014,N_12853,N_12829);
xor U13015 (N_13015,N_12971,N_12823);
nor U13016 (N_13016,N_12965,N_12922);
nor U13017 (N_13017,N_12948,N_12753);
or U13018 (N_13018,N_12859,N_12757);
nand U13019 (N_13019,N_12787,N_12932);
or U13020 (N_13020,N_12814,N_12754);
and U13021 (N_13021,N_12966,N_12873);
nor U13022 (N_13022,N_12825,N_12848);
xor U13023 (N_13023,N_12773,N_12983);
and U13024 (N_13024,N_12864,N_12815);
or U13025 (N_13025,N_12892,N_12991);
nor U13026 (N_13026,N_12821,N_12960);
or U13027 (N_13027,N_12944,N_12891);
nor U13028 (N_13028,N_12799,N_12979);
nand U13029 (N_13029,N_12877,N_12999);
nand U13030 (N_13030,N_12832,N_12899);
or U13031 (N_13031,N_12876,N_12826);
nand U13032 (N_13032,N_12950,N_12975);
xor U13033 (N_13033,N_12918,N_12834);
and U13034 (N_13034,N_12934,N_12844);
nand U13035 (N_13035,N_12854,N_12920);
nand U13036 (N_13036,N_12997,N_12984);
nand U13037 (N_13037,N_12903,N_12852);
or U13038 (N_13038,N_12946,N_12988);
xor U13039 (N_13039,N_12755,N_12951);
nor U13040 (N_13040,N_12772,N_12926);
or U13041 (N_13041,N_12953,N_12935);
or U13042 (N_13042,N_12769,N_12837);
nor U13043 (N_13043,N_12761,N_12908);
xnor U13044 (N_13044,N_12813,N_12851);
nor U13045 (N_13045,N_12811,N_12849);
and U13046 (N_13046,N_12940,N_12869);
xor U13047 (N_13047,N_12781,N_12827);
nor U13048 (N_13048,N_12820,N_12794);
nand U13049 (N_13049,N_12982,N_12955);
xor U13050 (N_13050,N_12828,N_12961);
nand U13051 (N_13051,N_12969,N_12939);
nand U13052 (N_13052,N_12791,N_12928);
nor U13053 (N_13053,N_12898,N_12850);
nor U13054 (N_13054,N_12783,N_12840);
and U13055 (N_13055,N_12987,N_12846);
xor U13056 (N_13056,N_12880,N_12830);
and U13057 (N_13057,N_12980,N_12949);
or U13058 (N_13058,N_12981,N_12902);
or U13059 (N_13059,N_12818,N_12912);
or U13060 (N_13060,N_12930,N_12917);
nor U13061 (N_13061,N_12874,N_12762);
nand U13062 (N_13062,N_12785,N_12861);
xor U13063 (N_13063,N_12998,N_12929);
nand U13064 (N_13064,N_12964,N_12750);
nor U13065 (N_13065,N_12875,N_12759);
xor U13066 (N_13066,N_12809,N_12808);
xnor U13067 (N_13067,N_12947,N_12976);
and U13068 (N_13068,N_12751,N_12802);
or U13069 (N_13069,N_12933,N_12901);
nor U13070 (N_13070,N_12943,N_12870);
nor U13071 (N_13071,N_12882,N_12835);
or U13072 (N_13072,N_12957,N_12879);
and U13073 (N_13073,N_12819,N_12894);
nand U13074 (N_13074,N_12890,N_12779);
and U13075 (N_13075,N_12843,N_12807);
nor U13076 (N_13076,N_12974,N_12765);
nor U13077 (N_13077,N_12790,N_12900);
nor U13078 (N_13078,N_12767,N_12778);
nor U13079 (N_13079,N_12868,N_12841);
and U13080 (N_13080,N_12866,N_12919);
or U13081 (N_13081,N_12914,N_12967);
nor U13082 (N_13082,N_12923,N_12889);
xnor U13083 (N_13083,N_12789,N_12812);
xnor U13084 (N_13084,N_12776,N_12800);
nand U13085 (N_13085,N_12992,N_12915);
or U13086 (N_13086,N_12937,N_12857);
or U13087 (N_13087,N_12885,N_12973);
nand U13088 (N_13088,N_12806,N_12764);
nand U13089 (N_13089,N_12780,N_12878);
or U13090 (N_13090,N_12931,N_12831);
and U13091 (N_13091,N_12886,N_12758);
xor U13092 (N_13092,N_12756,N_12768);
and U13093 (N_13093,N_12993,N_12796);
xor U13094 (N_13094,N_12782,N_12990);
or U13095 (N_13095,N_12836,N_12810);
nand U13096 (N_13096,N_12777,N_12775);
and U13097 (N_13097,N_12824,N_12871);
or U13098 (N_13098,N_12805,N_12883);
nand U13099 (N_13099,N_12972,N_12795);
or U13100 (N_13100,N_12968,N_12858);
nor U13101 (N_13101,N_12766,N_12959);
nor U13102 (N_13102,N_12989,N_12958);
or U13103 (N_13103,N_12996,N_12896);
or U13104 (N_13104,N_12977,N_12803);
and U13105 (N_13105,N_12786,N_12962);
nand U13106 (N_13106,N_12897,N_12895);
xor U13107 (N_13107,N_12942,N_12860);
xnor U13108 (N_13108,N_12910,N_12760);
or U13109 (N_13109,N_12817,N_12801);
xor U13110 (N_13110,N_12816,N_12938);
nand U13111 (N_13111,N_12924,N_12888);
or U13112 (N_13112,N_12956,N_12842);
nand U13113 (N_13113,N_12872,N_12822);
nand U13114 (N_13114,N_12833,N_12936);
xnor U13115 (N_13115,N_12867,N_12771);
and U13116 (N_13116,N_12921,N_12963);
nor U13117 (N_13117,N_12798,N_12913);
nor U13118 (N_13118,N_12862,N_12865);
and U13119 (N_13119,N_12847,N_12985);
and U13120 (N_13120,N_12994,N_12904);
nand U13121 (N_13121,N_12887,N_12927);
nand U13122 (N_13122,N_12763,N_12770);
nor U13123 (N_13123,N_12945,N_12906);
nand U13124 (N_13124,N_12916,N_12907);
nor U13125 (N_13125,N_12927,N_12832);
xnor U13126 (N_13126,N_12768,N_12854);
nand U13127 (N_13127,N_12997,N_12892);
nand U13128 (N_13128,N_12813,N_12773);
and U13129 (N_13129,N_12858,N_12960);
nor U13130 (N_13130,N_12800,N_12769);
nor U13131 (N_13131,N_12847,N_12818);
or U13132 (N_13132,N_12922,N_12796);
nor U13133 (N_13133,N_12929,N_12930);
nor U13134 (N_13134,N_12952,N_12846);
and U13135 (N_13135,N_12984,N_12981);
nor U13136 (N_13136,N_12938,N_12926);
nor U13137 (N_13137,N_12826,N_12866);
xor U13138 (N_13138,N_12778,N_12750);
nand U13139 (N_13139,N_12861,N_12869);
or U13140 (N_13140,N_12835,N_12914);
and U13141 (N_13141,N_12817,N_12824);
nand U13142 (N_13142,N_12798,N_12937);
and U13143 (N_13143,N_12830,N_12788);
nor U13144 (N_13144,N_12866,N_12769);
and U13145 (N_13145,N_12845,N_12991);
or U13146 (N_13146,N_12771,N_12756);
nor U13147 (N_13147,N_12917,N_12811);
and U13148 (N_13148,N_12811,N_12926);
or U13149 (N_13149,N_12884,N_12794);
xnor U13150 (N_13150,N_12772,N_12939);
and U13151 (N_13151,N_12752,N_12889);
nand U13152 (N_13152,N_12823,N_12750);
nand U13153 (N_13153,N_12891,N_12958);
and U13154 (N_13154,N_12943,N_12834);
nor U13155 (N_13155,N_12985,N_12896);
nor U13156 (N_13156,N_12772,N_12837);
or U13157 (N_13157,N_12756,N_12797);
or U13158 (N_13158,N_12987,N_12992);
nor U13159 (N_13159,N_12887,N_12758);
and U13160 (N_13160,N_12959,N_12772);
xor U13161 (N_13161,N_12759,N_12993);
or U13162 (N_13162,N_12927,N_12759);
xor U13163 (N_13163,N_12833,N_12858);
nor U13164 (N_13164,N_12848,N_12846);
nor U13165 (N_13165,N_12950,N_12889);
nor U13166 (N_13166,N_12953,N_12943);
nand U13167 (N_13167,N_12945,N_12860);
nor U13168 (N_13168,N_12860,N_12750);
and U13169 (N_13169,N_12811,N_12951);
nand U13170 (N_13170,N_12810,N_12795);
nor U13171 (N_13171,N_12891,N_12888);
xnor U13172 (N_13172,N_12951,N_12901);
and U13173 (N_13173,N_12819,N_12919);
and U13174 (N_13174,N_12961,N_12959);
nor U13175 (N_13175,N_12872,N_12997);
or U13176 (N_13176,N_12813,N_12767);
nor U13177 (N_13177,N_12759,N_12858);
and U13178 (N_13178,N_12976,N_12872);
nor U13179 (N_13179,N_12776,N_12856);
nand U13180 (N_13180,N_12909,N_12914);
and U13181 (N_13181,N_12967,N_12895);
nor U13182 (N_13182,N_12854,N_12839);
nor U13183 (N_13183,N_12756,N_12791);
and U13184 (N_13184,N_12800,N_12847);
and U13185 (N_13185,N_12943,N_12887);
or U13186 (N_13186,N_12806,N_12795);
nand U13187 (N_13187,N_12900,N_12751);
xor U13188 (N_13188,N_12848,N_12947);
nor U13189 (N_13189,N_12782,N_12894);
and U13190 (N_13190,N_12760,N_12950);
nor U13191 (N_13191,N_12872,N_12906);
xor U13192 (N_13192,N_12924,N_12957);
and U13193 (N_13193,N_12950,N_12971);
nand U13194 (N_13194,N_12888,N_12919);
nor U13195 (N_13195,N_12955,N_12845);
xnor U13196 (N_13196,N_12768,N_12820);
nor U13197 (N_13197,N_12920,N_12896);
or U13198 (N_13198,N_12950,N_12862);
and U13199 (N_13199,N_12776,N_12977);
nand U13200 (N_13200,N_12944,N_12856);
and U13201 (N_13201,N_12864,N_12845);
or U13202 (N_13202,N_12971,N_12802);
nor U13203 (N_13203,N_12938,N_12846);
or U13204 (N_13204,N_12919,N_12777);
nand U13205 (N_13205,N_12889,N_12969);
or U13206 (N_13206,N_12959,N_12758);
and U13207 (N_13207,N_12853,N_12772);
nor U13208 (N_13208,N_12828,N_12895);
xnor U13209 (N_13209,N_12838,N_12902);
nor U13210 (N_13210,N_12769,N_12964);
nand U13211 (N_13211,N_12892,N_12988);
nand U13212 (N_13212,N_12834,N_12843);
and U13213 (N_13213,N_12766,N_12970);
and U13214 (N_13214,N_12927,N_12925);
xor U13215 (N_13215,N_12967,N_12810);
and U13216 (N_13216,N_12751,N_12920);
nor U13217 (N_13217,N_12984,N_12992);
xnor U13218 (N_13218,N_12816,N_12754);
xor U13219 (N_13219,N_12913,N_12972);
xnor U13220 (N_13220,N_12781,N_12838);
xor U13221 (N_13221,N_12930,N_12758);
nor U13222 (N_13222,N_12886,N_12856);
nand U13223 (N_13223,N_12942,N_12885);
xnor U13224 (N_13224,N_12793,N_12982);
or U13225 (N_13225,N_12900,N_12973);
nand U13226 (N_13226,N_12872,N_12981);
or U13227 (N_13227,N_12896,N_12890);
nand U13228 (N_13228,N_12929,N_12921);
xor U13229 (N_13229,N_12964,N_12952);
xnor U13230 (N_13230,N_12807,N_12999);
and U13231 (N_13231,N_12788,N_12905);
nand U13232 (N_13232,N_12815,N_12953);
xor U13233 (N_13233,N_12939,N_12813);
or U13234 (N_13234,N_12913,N_12950);
and U13235 (N_13235,N_12967,N_12821);
nand U13236 (N_13236,N_12984,N_12875);
nand U13237 (N_13237,N_12910,N_12859);
or U13238 (N_13238,N_12929,N_12923);
nand U13239 (N_13239,N_12780,N_12853);
and U13240 (N_13240,N_12931,N_12906);
xor U13241 (N_13241,N_12802,N_12842);
xor U13242 (N_13242,N_12791,N_12945);
or U13243 (N_13243,N_12977,N_12946);
and U13244 (N_13244,N_12826,N_12787);
or U13245 (N_13245,N_12988,N_12807);
xor U13246 (N_13246,N_12835,N_12930);
nand U13247 (N_13247,N_12826,N_12879);
and U13248 (N_13248,N_12974,N_12903);
or U13249 (N_13249,N_12870,N_12810);
nor U13250 (N_13250,N_13241,N_13118);
nor U13251 (N_13251,N_13002,N_13160);
or U13252 (N_13252,N_13050,N_13062);
or U13253 (N_13253,N_13183,N_13012);
or U13254 (N_13254,N_13178,N_13000);
xor U13255 (N_13255,N_13126,N_13122);
or U13256 (N_13256,N_13009,N_13068);
nor U13257 (N_13257,N_13195,N_13100);
nand U13258 (N_13258,N_13010,N_13191);
nor U13259 (N_13259,N_13159,N_13200);
nand U13260 (N_13260,N_13131,N_13161);
or U13261 (N_13261,N_13085,N_13038);
nor U13262 (N_13262,N_13188,N_13235);
and U13263 (N_13263,N_13234,N_13021);
or U13264 (N_13264,N_13049,N_13249);
nand U13265 (N_13265,N_13051,N_13020);
or U13266 (N_13266,N_13084,N_13232);
or U13267 (N_13267,N_13157,N_13201);
nor U13268 (N_13268,N_13153,N_13215);
or U13269 (N_13269,N_13145,N_13179);
or U13270 (N_13270,N_13111,N_13106);
nand U13271 (N_13271,N_13208,N_13031);
xnor U13272 (N_13272,N_13152,N_13142);
nand U13273 (N_13273,N_13203,N_13034);
and U13274 (N_13274,N_13027,N_13086);
or U13275 (N_13275,N_13125,N_13028);
and U13276 (N_13276,N_13121,N_13093);
nand U13277 (N_13277,N_13124,N_13024);
or U13278 (N_13278,N_13040,N_13088);
xor U13279 (N_13279,N_13067,N_13070);
or U13280 (N_13280,N_13025,N_13029);
xor U13281 (N_13281,N_13063,N_13233);
or U13282 (N_13282,N_13081,N_13120);
xnor U13283 (N_13283,N_13218,N_13056);
xor U13284 (N_13284,N_13156,N_13190);
nor U13285 (N_13285,N_13207,N_13102);
or U13286 (N_13286,N_13146,N_13022);
or U13287 (N_13287,N_13026,N_13171);
or U13288 (N_13288,N_13023,N_13047);
xor U13289 (N_13289,N_13054,N_13212);
or U13290 (N_13290,N_13193,N_13003);
nor U13291 (N_13291,N_13032,N_13209);
and U13292 (N_13292,N_13147,N_13065);
nand U13293 (N_13293,N_13238,N_13139);
nor U13294 (N_13294,N_13204,N_13167);
xnor U13295 (N_13295,N_13134,N_13057);
or U13296 (N_13296,N_13089,N_13213);
or U13297 (N_13297,N_13141,N_13177);
xor U13298 (N_13298,N_13035,N_13078);
nand U13299 (N_13299,N_13044,N_13158);
and U13300 (N_13300,N_13189,N_13133);
and U13301 (N_13301,N_13148,N_13059);
and U13302 (N_13302,N_13228,N_13046);
nand U13303 (N_13303,N_13227,N_13237);
and U13304 (N_13304,N_13082,N_13090);
or U13305 (N_13305,N_13137,N_13172);
xnor U13306 (N_13306,N_13008,N_13135);
and U13307 (N_13307,N_13099,N_13069);
xor U13308 (N_13308,N_13229,N_13053);
nor U13309 (N_13309,N_13097,N_13214);
and U13310 (N_13310,N_13168,N_13109);
and U13311 (N_13311,N_13083,N_13030);
and U13312 (N_13312,N_13101,N_13048);
xnor U13313 (N_13313,N_13114,N_13007);
nand U13314 (N_13314,N_13144,N_13011);
and U13315 (N_13315,N_13013,N_13196);
nand U13316 (N_13316,N_13164,N_13066);
or U13317 (N_13317,N_13230,N_13071);
nor U13318 (N_13318,N_13155,N_13150);
nand U13319 (N_13319,N_13197,N_13181);
and U13320 (N_13320,N_13140,N_13154);
and U13321 (N_13321,N_13055,N_13061);
nand U13322 (N_13322,N_13015,N_13246);
nand U13323 (N_13323,N_13166,N_13079);
and U13324 (N_13324,N_13095,N_13143);
and U13325 (N_13325,N_13045,N_13006);
nor U13326 (N_13326,N_13104,N_13187);
or U13327 (N_13327,N_13036,N_13119);
and U13328 (N_13328,N_13018,N_13077);
nand U13329 (N_13329,N_13226,N_13244);
and U13330 (N_13330,N_13091,N_13103);
nor U13331 (N_13331,N_13202,N_13060);
or U13332 (N_13332,N_13001,N_13107);
nand U13333 (N_13333,N_13219,N_13073);
or U13334 (N_13334,N_13064,N_13243);
nor U13335 (N_13335,N_13130,N_13176);
nand U13336 (N_13336,N_13074,N_13217);
and U13337 (N_13337,N_13096,N_13169);
and U13338 (N_13338,N_13245,N_13162);
nand U13339 (N_13339,N_13239,N_13014);
nand U13340 (N_13340,N_13163,N_13129);
xor U13341 (N_13341,N_13185,N_13132);
nor U13342 (N_13342,N_13247,N_13205);
nand U13343 (N_13343,N_13248,N_13043);
or U13344 (N_13344,N_13211,N_13072);
xnor U13345 (N_13345,N_13198,N_13094);
nand U13346 (N_13346,N_13058,N_13165);
nand U13347 (N_13347,N_13223,N_13042);
or U13348 (N_13348,N_13080,N_13184);
xor U13349 (N_13349,N_13149,N_13019);
nand U13350 (N_13350,N_13175,N_13110);
and U13351 (N_13351,N_13174,N_13136);
nor U13352 (N_13352,N_13052,N_13231);
nand U13353 (N_13353,N_13180,N_13127);
nand U13354 (N_13354,N_13098,N_13075);
and U13355 (N_13355,N_13182,N_13087);
xnor U13356 (N_13356,N_13151,N_13092);
and U13357 (N_13357,N_13108,N_13115);
and U13358 (N_13358,N_13220,N_13225);
xor U13359 (N_13359,N_13186,N_13221);
xnor U13360 (N_13360,N_13076,N_13240);
or U13361 (N_13361,N_13222,N_13105);
or U13362 (N_13362,N_13037,N_13117);
nand U13363 (N_13363,N_13113,N_13170);
nand U13364 (N_13364,N_13041,N_13017);
xor U13365 (N_13365,N_13194,N_13199);
or U13366 (N_13366,N_13004,N_13039);
or U13367 (N_13367,N_13173,N_13016);
nor U13368 (N_13368,N_13005,N_13236);
or U13369 (N_13369,N_13138,N_13210);
or U13370 (N_13370,N_13033,N_13192);
nor U13371 (N_13371,N_13116,N_13242);
nor U13372 (N_13372,N_13206,N_13216);
nand U13373 (N_13373,N_13224,N_13123);
nand U13374 (N_13374,N_13112,N_13128);
nor U13375 (N_13375,N_13054,N_13106);
nor U13376 (N_13376,N_13171,N_13229);
or U13377 (N_13377,N_13187,N_13075);
and U13378 (N_13378,N_13118,N_13024);
nor U13379 (N_13379,N_13234,N_13225);
or U13380 (N_13380,N_13184,N_13094);
and U13381 (N_13381,N_13039,N_13152);
or U13382 (N_13382,N_13066,N_13021);
and U13383 (N_13383,N_13200,N_13107);
nand U13384 (N_13384,N_13175,N_13214);
or U13385 (N_13385,N_13069,N_13227);
and U13386 (N_13386,N_13153,N_13044);
nand U13387 (N_13387,N_13013,N_13056);
xor U13388 (N_13388,N_13146,N_13104);
nor U13389 (N_13389,N_13058,N_13160);
or U13390 (N_13390,N_13110,N_13028);
nand U13391 (N_13391,N_13035,N_13183);
nand U13392 (N_13392,N_13081,N_13135);
nand U13393 (N_13393,N_13193,N_13077);
nand U13394 (N_13394,N_13150,N_13247);
and U13395 (N_13395,N_13110,N_13179);
nand U13396 (N_13396,N_13128,N_13036);
or U13397 (N_13397,N_13177,N_13246);
or U13398 (N_13398,N_13082,N_13159);
or U13399 (N_13399,N_13125,N_13031);
nor U13400 (N_13400,N_13204,N_13032);
or U13401 (N_13401,N_13100,N_13029);
nor U13402 (N_13402,N_13013,N_13102);
nor U13403 (N_13403,N_13085,N_13018);
nand U13404 (N_13404,N_13011,N_13008);
nor U13405 (N_13405,N_13047,N_13135);
and U13406 (N_13406,N_13231,N_13211);
and U13407 (N_13407,N_13029,N_13121);
nand U13408 (N_13408,N_13014,N_13210);
nand U13409 (N_13409,N_13193,N_13038);
nor U13410 (N_13410,N_13079,N_13158);
nor U13411 (N_13411,N_13195,N_13162);
and U13412 (N_13412,N_13125,N_13199);
nand U13413 (N_13413,N_13107,N_13050);
nand U13414 (N_13414,N_13157,N_13006);
and U13415 (N_13415,N_13209,N_13021);
and U13416 (N_13416,N_13017,N_13247);
nand U13417 (N_13417,N_13028,N_13029);
xor U13418 (N_13418,N_13027,N_13131);
nand U13419 (N_13419,N_13249,N_13047);
xor U13420 (N_13420,N_13079,N_13017);
nor U13421 (N_13421,N_13246,N_13035);
and U13422 (N_13422,N_13198,N_13089);
and U13423 (N_13423,N_13155,N_13130);
and U13424 (N_13424,N_13043,N_13002);
xnor U13425 (N_13425,N_13095,N_13076);
nor U13426 (N_13426,N_13112,N_13246);
or U13427 (N_13427,N_13228,N_13097);
or U13428 (N_13428,N_13146,N_13212);
xnor U13429 (N_13429,N_13012,N_13176);
and U13430 (N_13430,N_13218,N_13066);
nor U13431 (N_13431,N_13076,N_13217);
and U13432 (N_13432,N_13131,N_13208);
xnor U13433 (N_13433,N_13037,N_13090);
and U13434 (N_13434,N_13094,N_13039);
and U13435 (N_13435,N_13205,N_13038);
and U13436 (N_13436,N_13147,N_13111);
xor U13437 (N_13437,N_13101,N_13147);
nor U13438 (N_13438,N_13247,N_13242);
nand U13439 (N_13439,N_13189,N_13130);
and U13440 (N_13440,N_13229,N_13076);
or U13441 (N_13441,N_13020,N_13063);
or U13442 (N_13442,N_13135,N_13201);
and U13443 (N_13443,N_13126,N_13046);
nor U13444 (N_13444,N_13075,N_13215);
nand U13445 (N_13445,N_13141,N_13155);
xor U13446 (N_13446,N_13157,N_13045);
xnor U13447 (N_13447,N_13152,N_13020);
or U13448 (N_13448,N_13239,N_13191);
nand U13449 (N_13449,N_13105,N_13063);
or U13450 (N_13450,N_13205,N_13102);
nand U13451 (N_13451,N_13208,N_13184);
and U13452 (N_13452,N_13088,N_13083);
or U13453 (N_13453,N_13241,N_13240);
nand U13454 (N_13454,N_13042,N_13079);
nor U13455 (N_13455,N_13128,N_13089);
or U13456 (N_13456,N_13138,N_13098);
or U13457 (N_13457,N_13003,N_13157);
xnor U13458 (N_13458,N_13101,N_13122);
xor U13459 (N_13459,N_13056,N_13132);
or U13460 (N_13460,N_13007,N_13039);
xnor U13461 (N_13461,N_13005,N_13058);
nor U13462 (N_13462,N_13158,N_13011);
and U13463 (N_13463,N_13015,N_13143);
and U13464 (N_13464,N_13124,N_13199);
or U13465 (N_13465,N_13016,N_13188);
nand U13466 (N_13466,N_13191,N_13167);
nand U13467 (N_13467,N_13120,N_13218);
xnor U13468 (N_13468,N_13116,N_13001);
xnor U13469 (N_13469,N_13081,N_13067);
and U13470 (N_13470,N_13114,N_13224);
nor U13471 (N_13471,N_13113,N_13069);
nand U13472 (N_13472,N_13222,N_13183);
nand U13473 (N_13473,N_13219,N_13206);
or U13474 (N_13474,N_13119,N_13108);
nand U13475 (N_13475,N_13248,N_13152);
xor U13476 (N_13476,N_13142,N_13124);
nor U13477 (N_13477,N_13204,N_13180);
nor U13478 (N_13478,N_13096,N_13073);
nor U13479 (N_13479,N_13145,N_13072);
xor U13480 (N_13480,N_13008,N_13162);
xnor U13481 (N_13481,N_13066,N_13237);
xnor U13482 (N_13482,N_13029,N_13249);
and U13483 (N_13483,N_13237,N_13009);
and U13484 (N_13484,N_13207,N_13030);
xor U13485 (N_13485,N_13232,N_13052);
nand U13486 (N_13486,N_13120,N_13073);
and U13487 (N_13487,N_13115,N_13130);
or U13488 (N_13488,N_13240,N_13063);
and U13489 (N_13489,N_13226,N_13109);
xor U13490 (N_13490,N_13093,N_13131);
nand U13491 (N_13491,N_13168,N_13128);
nand U13492 (N_13492,N_13067,N_13024);
nand U13493 (N_13493,N_13011,N_13138);
and U13494 (N_13494,N_13237,N_13232);
and U13495 (N_13495,N_13019,N_13005);
nand U13496 (N_13496,N_13223,N_13230);
nand U13497 (N_13497,N_13014,N_13151);
nor U13498 (N_13498,N_13081,N_13210);
or U13499 (N_13499,N_13202,N_13114);
nor U13500 (N_13500,N_13276,N_13256);
or U13501 (N_13501,N_13293,N_13262);
nor U13502 (N_13502,N_13279,N_13302);
nor U13503 (N_13503,N_13398,N_13266);
nand U13504 (N_13504,N_13362,N_13410);
or U13505 (N_13505,N_13259,N_13318);
xor U13506 (N_13506,N_13379,N_13407);
or U13507 (N_13507,N_13455,N_13476);
nand U13508 (N_13508,N_13359,N_13422);
nand U13509 (N_13509,N_13369,N_13451);
or U13510 (N_13510,N_13340,N_13316);
nand U13511 (N_13511,N_13322,N_13471);
nor U13512 (N_13512,N_13310,N_13389);
or U13513 (N_13513,N_13271,N_13288);
and U13514 (N_13514,N_13339,N_13443);
nor U13515 (N_13515,N_13429,N_13448);
nor U13516 (N_13516,N_13463,N_13433);
or U13517 (N_13517,N_13394,N_13277);
xnor U13518 (N_13518,N_13396,N_13487);
nor U13519 (N_13519,N_13417,N_13481);
xnor U13520 (N_13520,N_13406,N_13352);
or U13521 (N_13521,N_13499,N_13392);
xnor U13522 (N_13522,N_13258,N_13349);
and U13523 (N_13523,N_13364,N_13434);
and U13524 (N_13524,N_13432,N_13368);
nor U13525 (N_13525,N_13409,N_13365);
or U13526 (N_13526,N_13395,N_13405);
nand U13527 (N_13527,N_13336,N_13430);
xnor U13528 (N_13528,N_13294,N_13486);
nand U13529 (N_13529,N_13378,N_13470);
or U13530 (N_13530,N_13263,N_13357);
nand U13531 (N_13531,N_13492,N_13327);
nor U13532 (N_13532,N_13478,N_13411);
xor U13533 (N_13533,N_13458,N_13496);
or U13534 (N_13534,N_13313,N_13418);
xnor U13535 (N_13535,N_13498,N_13402);
xnor U13536 (N_13536,N_13283,N_13298);
and U13537 (N_13537,N_13399,N_13341);
and U13538 (N_13538,N_13356,N_13252);
or U13539 (N_13539,N_13353,N_13388);
nor U13540 (N_13540,N_13255,N_13260);
nor U13541 (N_13541,N_13482,N_13315);
nor U13542 (N_13542,N_13397,N_13329);
nand U13543 (N_13543,N_13377,N_13408);
xor U13544 (N_13544,N_13253,N_13452);
and U13545 (N_13545,N_13366,N_13461);
nand U13546 (N_13546,N_13464,N_13462);
or U13547 (N_13547,N_13424,N_13428);
nand U13548 (N_13548,N_13390,N_13484);
nor U13549 (N_13549,N_13494,N_13449);
nor U13550 (N_13550,N_13441,N_13281);
or U13551 (N_13551,N_13274,N_13337);
nand U13552 (N_13552,N_13420,N_13426);
or U13553 (N_13553,N_13400,N_13342);
nand U13554 (N_13554,N_13438,N_13335);
nor U13555 (N_13555,N_13373,N_13473);
or U13556 (N_13556,N_13250,N_13306);
nand U13557 (N_13557,N_13278,N_13257);
and U13558 (N_13558,N_13325,N_13480);
nand U13559 (N_13559,N_13404,N_13477);
or U13560 (N_13560,N_13334,N_13297);
nand U13561 (N_13561,N_13370,N_13270);
and U13562 (N_13562,N_13305,N_13427);
and U13563 (N_13563,N_13374,N_13344);
and U13564 (N_13564,N_13413,N_13436);
and U13565 (N_13565,N_13483,N_13421);
and U13566 (N_13566,N_13284,N_13382);
nand U13567 (N_13567,N_13360,N_13412);
xnor U13568 (N_13568,N_13460,N_13381);
or U13569 (N_13569,N_13268,N_13350);
or U13570 (N_13570,N_13367,N_13401);
nand U13571 (N_13571,N_13375,N_13273);
and U13572 (N_13572,N_13457,N_13269);
nor U13573 (N_13573,N_13384,N_13431);
and U13574 (N_13574,N_13435,N_13348);
xor U13575 (N_13575,N_13300,N_13456);
xnor U13576 (N_13576,N_13466,N_13376);
and U13577 (N_13577,N_13311,N_13465);
or U13578 (N_13578,N_13346,N_13312);
xnor U13579 (N_13579,N_13459,N_13267);
nand U13580 (N_13580,N_13296,N_13415);
or U13581 (N_13581,N_13425,N_13345);
nor U13582 (N_13582,N_13304,N_13383);
xor U13583 (N_13583,N_13391,N_13272);
nand U13584 (N_13584,N_13468,N_13347);
nor U13585 (N_13585,N_13446,N_13385);
xnor U13586 (N_13586,N_13475,N_13307);
and U13587 (N_13587,N_13488,N_13324);
nor U13588 (N_13588,N_13264,N_13393);
nand U13589 (N_13589,N_13423,N_13491);
xnor U13590 (N_13590,N_13386,N_13387);
nor U13591 (N_13591,N_13380,N_13419);
and U13592 (N_13592,N_13439,N_13447);
xnor U13593 (N_13593,N_13454,N_13343);
xor U13594 (N_13594,N_13354,N_13372);
and U13595 (N_13595,N_13403,N_13437);
and U13596 (N_13596,N_13285,N_13444);
and U13597 (N_13597,N_13363,N_13251);
and U13598 (N_13598,N_13291,N_13295);
and U13599 (N_13599,N_13319,N_13453);
nand U13600 (N_13600,N_13282,N_13314);
or U13601 (N_13601,N_13440,N_13299);
and U13602 (N_13602,N_13289,N_13489);
nand U13603 (N_13603,N_13320,N_13309);
xor U13604 (N_13604,N_13321,N_13414);
and U13605 (N_13605,N_13261,N_13317);
and U13606 (N_13606,N_13287,N_13416);
xnor U13607 (N_13607,N_13371,N_13328);
nand U13608 (N_13608,N_13497,N_13323);
nor U13609 (N_13609,N_13331,N_13301);
or U13610 (N_13610,N_13445,N_13493);
nor U13611 (N_13611,N_13286,N_13265);
nor U13612 (N_13612,N_13450,N_13442);
nor U13613 (N_13613,N_13330,N_13292);
xnor U13614 (N_13614,N_13290,N_13469);
or U13615 (N_13615,N_13308,N_13490);
xnor U13616 (N_13616,N_13485,N_13351);
nand U13617 (N_13617,N_13479,N_13303);
nand U13618 (N_13618,N_13355,N_13326);
nor U13619 (N_13619,N_13275,N_13472);
xor U13620 (N_13620,N_13474,N_13280);
xor U13621 (N_13621,N_13358,N_13332);
and U13622 (N_13622,N_13254,N_13495);
nand U13623 (N_13623,N_13333,N_13361);
nand U13624 (N_13624,N_13467,N_13338);
xnor U13625 (N_13625,N_13392,N_13383);
and U13626 (N_13626,N_13415,N_13250);
and U13627 (N_13627,N_13302,N_13333);
nand U13628 (N_13628,N_13263,N_13418);
xor U13629 (N_13629,N_13441,N_13463);
nor U13630 (N_13630,N_13301,N_13384);
and U13631 (N_13631,N_13258,N_13497);
or U13632 (N_13632,N_13374,N_13475);
nand U13633 (N_13633,N_13439,N_13331);
and U13634 (N_13634,N_13337,N_13499);
nor U13635 (N_13635,N_13296,N_13307);
xnor U13636 (N_13636,N_13407,N_13476);
and U13637 (N_13637,N_13487,N_13307);
nor U13638 (N_13638,N_13469,N_13446);
or U13639 (N_13639,N_13307,N_13370);
xnor U13640 (N_13640,N_13256,N_13481);
or U13641 (N_13641,N_13425,N_13258);
nor U13642 (N_13642,N_13338,N_13447);
or U13643 (N_13643,N_13405,N_13373);
nor U13644 (N_13644,N_13298,N_13413);
nand U13645 (N_13645,N_13262,N_13357);
nor U13646 (N_13646,N_13345,N_13492);
and U13647 (N_13647,N_13359,N_13362);
or U13648 (N_13648,N_13395,N_13257);
and U13649 (N_13649,N_13353,N_13365);
and U13650 (N_13650,N_13399,N_13269);
and U13651 (N_13651,N_13372,N_13428);
xor U13652 (N_13652,N_13375,N_13435);
nand U13653 (N_13653,N_13351,N_13470);
or U13654 (N_13654,N_13482,N_13381);
and U13655 (N_13655,N_13353,N_13349);
or U13656 (N_13656,N_13264,N_13437);
xor U13657 (N_13657,N_13433,N_13275);
xnor U13658 (N_13658,N_13280,N_13440);
and U13659 (N_13659,N_13318,N_13250);
and U13660 (N_13660,N_13447,N_13438);
nand U13661 (N_13661,N_13487,N_13304);
xor U13662 (N_13662,N_13495,N_13294);
nand U13663 (N_13663,N_13264,N_13339);
nor U13664 (N_13664,N_13480,N_13280);
and U13665 (N_13665,N_13294,N_13426);
nor U13666 (N_13666,N_13327,N_13459);
nor U13667 (N_13667,N_13400,N_13403);
and U13668 (N_13668,N_13352,N_13482);
nor U13669 (N_13669,N_13413,N_13268);
nor U13670 (N_13670,N_13339,N_13416);
nor U13671 (N_13671,N_13384,N_13381);
or U13672 (N_13672,N_13253,N_13351);
nand U13673 (N_13673,N_13334,N_13484);
or U13674 (N_13674,N_13383,N_13404);
nor U13675 (N_13675,N_13391,N_13409);
xnor U13676 (N_13676,N_13332,N_13361);
nand U13677 (N_13677,N_13352,N_13403);
and U13678 (N_13678,N_13274,N_13316);
nor U13679 (N_13679,N_13279,N_13288);
nand U13680 (N_13680,N_13289,N_13474);
and U13681 (N_13681,N_13337,N_13425);
and U13682 (N_13682,N_13289,N_13446);
or U13683 (N_13683,N_13269,N_13493);
nor U13684 (N_13684,N_13317,N_13473);
nand U13685 (N_13685,N_13322,N_13254);
and U13686 (N_13686,N_13448,N_13269);
nor U13687 (N_13687,N_13401,N_13278);
and U13688 (N_13688,N_13480,N_13447);
and U13689 (N_13689,N_13294,N_13304);
or U13690 (N_13690,N_13419,N_13328);
nor U13691 (N_13691,N_13443,N_13258);
nor U13692 (N_13692,N_13333,N_13379);
xnor U13693 (N_13693,N_13263,N_13328);
and U13694 (N_13694,N_13362,N_13344);
and U13695 (N_13695,N_13460,N_13327);
nand U13696 (N_13696,N_13427,N_13273);
and U13697 (N_13697,N_13306,N_13332);
and U13698 (N_13698,N_13293,N_13436);
nor U13699 (N_13699,N_13483,N_13481);
or U13700 (N_13700,N_13461,N_13484);
or U13701 (N_13701,N_13285,N_13459);
nor U13702 (N_13702,N_13330,N_13293);
and U13703 (N_13703,N_13430,N_13395);
xnor U13704 (N_13704,N_13341,N_13383);
or U13705 (N_13705,N_13494,N_13303);
xor U13706 (N_13706,N_13447,N_13372);
and U13707 (N_13707,N_13303,N_13436);
xnor U13708 (N_13708,N_13308,N_13495);
nor U13709 (N_13709,N_13336,N_13257);
or U13710 (N_13710,N_13265,N_13459);
nor U13711 (N_13711,N_13303,N_13400);
or U13712 (N_13712,N_13444,N_13402);
or U13713 (N_13713,N_13460,N_13304);
nor U13714 (N_13714,N_13356,N_13253);
nor U13715 (N_13715,N_13415,N_13299);
nor U13716 (N_13716,N_13268,N_13271);
xor U13717 (N_13717,N_13457,N_13452);
and U13718 (N_13718,N_13319,N_13426);
nor U13719 (N_13719,N_13423,N_13386);
nor U13720 (N_13720,N_13382,N_13294);
xor U13721 (N_13721,N_13380,N_13475);
nor U13722 (N_13722,N_13387,N_13319);
nand U13723 (N_13723,N_13338,N_13286);
xnor U13724 (N_13724,N_13254,N_13414);
nor U13725 (N_13725,N_13286,N_13499);
or U13726 (N_13726,N_13318,N_13487);
nor U13727 (N_13727,N_13279,N_13348);
nand U13728 (N_13728,N_13450,N_13324);
nor U13729 (N_13729,N_13333,N_13318);
and U13730 (N_13730,N_13375,N_13424);
xnor U13731 (N_13731,N_13355,N_13254);
or U13732 (N_13732,N_13441,N_13453);
xor U13733 (N_13733,N_13381,N_13401);
xor U13734 (N_13734,N_13369,N_13416);
nand U13735 (N_13735,N_13298,N_13476);
nor U13736 (N_13736,N_13417,N_13488);
nor U13737 (N_13737,N_13285,N_13317);
or U13738 (N_13738,N_13327,N_13256);
nor U13739 (N_13739,N_13453,N_13472);
nand U13740 (N_13740,N_13415,N_13428);
nand U13741 (N_13741,N_13340,N_13260);
nor U13742 (N_13742,N_13376,N_13430);
nand U13743 (N_13743,N_13413,N_13301);
and U13744 (N_13744,N_13262,N_13344);
nand U13745 (N_13745,N_13317,N_13333);
or U13746 (N_13746,N_13455,N_13468);
and U13747 (N_13747,N_13439,N_13301);
xnor U13748 (N_13748,N_13457,N_13273);
nor U13749 (N_13749,N_13303,N_13334);
and U13750 (N_13750,N_13573,N_13746);
nor U13751 (N_13751,N_13611,N_13724);
and U13752 (N_13752,N_13632,N_13668);
nand U13753 (N_13753,N_13650,N_13545);
nand U13754 (N_13754,N_13686,N_13606);
or U13755 (N_13755,N_13639,N_13560);
and U13756 (N_13756,N_13676,N_13648);
xnor U13757 (N_13757,N_13553,N_13695);
nor U13758 (N_13758,N_13587,N_13540);
nand U13759 (N_13759,N_13563,N_13726);
or U13760 (N_13760,N_13674,N_13571);
and U13761 (N_13761,N_13710,N_13514);
xnor U13762 (N_13762,N_13530,N_13538);
nand U13763 (N_13763,N_13511,N_13703);
nor U13764 (N_13764,N_13597,N_13600);
xor U13765 (N_13765,N_13679,N_13578);
nand U13766 (N_13766,N_13633,N_13715);
nor U13767 (N_13767,N_13680,N_13594);
and U13768 (N_13768,N_13512,N_13691);
or U13769 (N_13769,N_13559,N_13651);
or U13770 (N_13770,N_13721,N_13637);
and U13771 (N_13771,N_13670,N_13631);
xnor U13772 (N_13772,N_13604,N_13592);
nor U13773 (N_13773,N_13602,N_13605);
nand U13774 (N_13774,N_13630,N_13687);
and U13775 (N_13775,N_13628,N_13525);
nand U13776 (N_13776,N_13718,N_13623);
nand U13777 (N_13777,N_13515,N_13603);
or U13778 (N_13778,N_13554,N_13655);
and U13779 (N_13779,N_13619,N_13681);
xor U13780 (N_13780,N_13601,N_13504);
or U13781 (N_13781,N_13644,N_13685);
xor U13782 (N_13782,N_13641,N_13636);
or U13783 (N_13783,N_13565,N_13572);
nor U13784 (N_13784,N_13503,N_13555);
nor U13785 (N_13785,N_13656,N_13591);
nand U13786 (N_13786,N_13666,N_13513);
xnor U13787 (N_13787,N_13556,N_13736);
xor U13788 (N_13788,N_13694,N_13742);
or U13789 (N_13789,N_13539,N_13558);
nor U13790 (N_13790,N_13719,N_13716);
nand U13791 (N_13791,N_13502,N_13664);
or U13792 (N_13792,N_13568,N_13708);
and U13793 (N_13793,N_13652,N_13678);
nand U13794 (N_13794,N_13677,N_13642);
nor U13795 (N_13795,N_13638,N_13616);
nand U13796 (N_13796,N_13730,N_13684);
xnor U13797 (N_13797,N_13720,N_13534);
nand U13798 (N_13798,N_13585,N_13582);
and U13799 (N_13799,N_13599,N_13576);
xnor U13800 (N_13800,N_13734,N_13612);
and U13801 (N_13801,N_13618,N_13743);
or U13802 (N_13802,N_13609,N_13693);
and U13803 (N_13803,N_13527,N_13510);
xnor U13804 (N_13804,N_13729,N_13624);
xor U13805 (N_13805,N_13557,N_13627);
and U13806 (N_13806,N_13675,N_13508);
nor U13807 (N_13807,N_13562,N_13712);
nor U13808 (N_13808,N_13598,N_13688);
nor U13809 (N_13809,N_13672,N_13653);
or U13810 (N_13810,N_13584,N_13595);
nand U13811 (N_13811,N_13643,N_13613);
xnor U13812 (N_13812,N_13660,N_13709);
and U13813 (N_13813,N_13564,N_13589);
and U13814 (N_13814,N_13698,N_13745);
and U13815 (N_13815,N_13516,N_13533);
nor U13816 (N_13816,N_13647,N_13546);
nor U13817 (N_13817,N_13583,N_13551);
nor U13818 (N_13818,N_13531,N_13506);
or U13819 (N_13819,N_13741,N_13544);
and U13820 (N_13820,N_13748,N_13532);
nand U13821 (N_13821,N_13661,N_13649);
nor U13822 (N_13822,N_13535,N_13524);
xor U13823 (N_13823,N_13671,N_13588);
xnor U13824 (N_13824,N_13529,N_13728);
or U13825 (N_13825,N_13705,N_13579);
xnor U13826 (N_13826,N_13574,N_13702);
xor U13827 (N_13827,N_13733,N_13581);
and U13828 (N_13828,N_13727,N_13566);
xnor U13829 (N_13829,N_13521,N_13569);
and U13830 (N_13830,N_13629,N_13747);
xnor U13831 (N_13831,N_13500,N_13615);
or U13832 (N_13832,N_13580,N_13586);
or U13833 (N_13833,N_13682,N_13522);
nor U13834 (N_13834,N_13714,N_13704);
or U13835 (N_13835,N_13738,N_13622);
nand U13836 (N_13836,N_13608,N_13593);
nand U13837 (N_13837,N_13725,N_13626);
nand U13838 (N_13838,N_13659,N_13723);
and U13839 (N_13839,N_13662,N_13739);
nand U13840 (N_13840,N_13700,N_13596);
xor U13841 (N_13841,N_13737,N_13614);
xor U13842 (N_13842,N_13732,N_13518);
and U13843 (N_13843,N_13749,N_13634);
and U13844 (N_13844,N_13543,N_13526);
xor U13845 (N_13845,N_13667,N_13706);
xor U13846 (N_13846,N_13713,N_13567);
xor U13847 (N_13847,N_13617,N_13561);
xor U13848 (N_13848,N_13519,N_13520);
and U13849 (N_13849,N_13645,N_13699);
xnor U13850 (N_13850,N_13505,N_13646);
or U13851 (N_13851,N_13590,N_13549);
and U13852 (N_13852,N_13683,N_13707);
nor U13853 (N_13853,N_13552,N_13658);
and U13854 (N_13854,N_13528,N_13547);
and U13855 (N_13855,N_13536,N_13577);
or U13856 (N_13856,N_13735,N_13697);
xor U13857 (N_13857,N_13692,N_13717);
xor U13858 (N_13858,N_13610,N_13625);
xnor U13859 (N_13859,N_13657,N_13690);
or U13860 (N_13860,N_13744,N_13620);
xnor U13861 (N_13861,N_13669,N_13541);
nand U13862 (N_13862,N_13711,N_13517);
xor U13863 (N_13863,N_13509,N_13548);
xor U13864 (N_13864,N_13722,N_13740);
nand U13865 (N_13865,N_13696,N_13550);
xnor U13866 (N_13866,N_13731,N_13640);
xor U13867 (N_13867,N_13542,N_13575);
and U13868 (N_13868,N_13665,N_13570);
xnor U13869 (N_13869,N_13507,N_13635);
and U13870 (N_13870,N_13673,N_13537);
nand U13871 (N_13871,N_13689,N_13621);
and U13872 (N_13872,N_13501,N_13523);
or U13873 (N_13873,N_13607,N_13663);
or U13874 (N_13874,N_13654,N_13701);
xnor U13875 (N_13875,N_13646,N_13652);
and U13876 (N_13876,N_13595,N_13742);
nor U13877 (N_13877,N_13640,N_13660);
nor U13878 (N_13878,N_13502,N_13653);
and U13879 (N_13879,N_13704,N_13574);
nand U13880 (N_13880,N_13703,N_13689);
nor U13881 (N_13881,N_13590,N_13524);
nor U13882 (N_13882,N_13615,N_13596);
or U13883 (N_13883,N_13705,N_13734);
or U13884 (N_13884,N_13694,N_13708);
nand U13885 (N_13885,N_13563,N_13730);
xnor U13886 (N_13886,N_13584,N_13613);
xnor U13887 (N_13887,N_13564,N_13661);
nor U13888 (N_13888,N_13693,N_13543);
xor U13889 (N_13889,N_13714,N_13552);
or U13890 (N_13890,N_13723,N_13559);
nor U13891 (N_13891,N_13724,N_13710);
xor U13892 (N_13892,N_13696,N_13555);
nor U13893 (N_13893,N_13528,N_13642);
xor U13894 (N_13894,N_13542,N_13607);
and U13895 (N_13895,N_13620,N_13533);
or U13896 (N_13896,N_13629,N_13672);
nand U13897 (N_13897,N_13643,N_13609);
or U13898 (N_13898,N_13716,N_13593);
or U13899 (N_13899,N_13548,N_13688);
nand U13900 (N_13900,N_13627,N_13511);
nor U13901 (N_13901,N_13534,N_13700);
or U13902 (N_13902,N_13589,N_13599);
or U13903 (N_13903,N_13714,N_13683);
and U13904 (N_13904,N_13526,N_13590);
xor U13905 (N_13905,N_13690,N_13721);
or U13906 (N_13906,N_13524,N_13647);
nand U13907 (N_13907,N_13564,N_13666);
nor U13908 (N_13908,N_13521,N_13536);
nor U13909 (N_13909,N_13584,N_13580);
nand U13910 (N_13910,N_13561,N_13546);
nand U13911 (N_13911,N_13732,N_13683);
or U13912 (N_13912,N_13654,N_13623);
xnor U13913 (N_13913,N_13655,N_13541);
nand U13914 (N_13914,N_13718,N_13715);
or U13915 (N_13915,N_13730,N_13617);
xnor U13916 (N_13916,N_13657,N_13548);
nor U13917 (N_13917,N_13540,N_13614);
or U13918 (N_13918,N_13636,N_13723);
and U13919 (N_13919,N_13564,N_13582);
xnor U13920 (N_13920,N_13626,N_13620);
and U13921 (N_13921,N_13537,N_13560);
nand U13922 (N_13922,N_13605,N_13666);
xor U13923 (N_13923,N_13706,N_13581);
xnor U13924 (N_13924,N_13503,N_13525);
nand U13925 (N_13925,N_13669,N_13574);
or U13926 (N_13926,N_13521,N_13531);
nor U13927 (N_13927,N_13715,N_13613);
and U13928 (N_13928,N_13516,N_13744);
nand U13929 (N_13929,N_13748,N_13663);
nand U13930 (N_13930,N_13512,N_13681);
or U13931 (N_13931,N_13579,N_13553);
nand U13932 (N_13932,N_13676,N_13597);
nor U13933 (N_13933,N_13649,N_13643);
and U13934 (N_13934,N_13653,N_13530);
nand U13935 (N_13935,N_13600,N_13550);
nor U13936 (N_13936,N_13501,N_13628);
or U13937 (N_13937,N_13644,N_13710);
nor U13938 (N_13938,N_13662,N_13658);
nor U13939 (N_13939,N_13580,N_13671);
and U13940 (N_13940,N_13740,N_13550);
nor U13941 (N_13941,N_13649,N_13537);
or U13942 (N_13942,N_13508,N_13558);
xnor U13943 (N_13943,N_13546,N_13694);
xor U13944 (N_13944,N_13578,N_13748);
and U13945 (N_13945,N_13522,N_13604);
or U13946 (N_13946,N_13648,N_13598);
nand U13947 (N_13947,N_13566,N_13660);
or U13948 (N_13948,N_13577,N_13739);
and U13949 (N_13949,N_13574,N_13693);
nor U13950 (N_13950,N_13555,N_13616);
or U13951 (N_13951,N_13738,N_13696);
nor U13952 (N_13952,N_13714,N_13645);
and U13953 (N_13953,N_13631,N_13501);
and U13954 (N_13954,N_13726,N_13681);
and U13955 (N_13955,N_13545,N_13570);
or U13956 (N_13956,N_13545,N_13554);
or U13957 (N_13957,N_13695,N_13515);
or U13958 (N_13958,N_13509,N_13551);
xnor U13959 (N_13959,N_13527,N_13582);
nand U13960 (N_13960,N_13540,N_13564);
nand U13961 (N_13961,N_13711,N_13728);
xor U13962 (N_13962,N_13741,N_13546);
and U13963 (N_13963,N_13699,N_13679);
or U13964 (N_13964,N_13665,N_13746);
nand U13965 (N_13965,N_13662,N_13652);
or U13966 (N_13966,N_13656,N_13636);
or U13967 (N_13967,N_13528,N_13633);
nand U13968 (N_13968,N_13521,N_13675);
and U13969 (N_13969,N_13617,N_13536);
nor U13970 (N_13970,N_13701,N_13735);
xor U13971 (N_13971,N_13730,N_13670);
and U13972 (N_13972,N_13654,N_13641);
and U13973 (N_13973,N_13565,N_13553);
xnor U13974 (N_13974,N_13500,N_13632);
or U13975 (N_13975,N_13705,N_13654);
nor U13976 (N_13976,N_13598,N_13548);
and U13977 (N_13977,N_13568,N_13598);
nand U13978 (N_13978,N_13676,N_13679);
xnor U13979 (N_13979,N_13616,N_13736);
and U13980 (N_13980,N_13738,N_13694);
nor U13981 (N_13981,N_13698,N_13684);
and U13982 (N_13982,N_13715,N_13711);
or U13983 (N_13983,N_13707,N_13546);
or U13984 (N_13984,N_13565,N_13711);
nor U13985 (N_13985,N_13583,N_13683);
or U13986 (N_13986,N_13679,N_13638);
nor U13987 (N_13987,N_13724,N_13563);
or U13988 (N_13988,N_13619,N_13562);
and U13989 (N_13989,N_13603,N_13729);
and U13990 (N_13990,N_13630,N_13603);
or U13991 (N_13991,N_13525,N_13635);
and U13992 (N_13992,N_13695,N_13599);
nand U13993 (N_13993,N_13619,N_13746);
nand U13994 (N_13994,N_13665,N_13616);
and U13995 (N_13995,N_13615,N_13699);
xnor U13996 (N_13996,N_13561,N_13710);
and U13997 (N_13997,N_13743,N_13704);
and U13998 (N_13998,N_13700,N_13695);
or U13999 (N_13999,N_13507,N_13555);
and U14000 (N_14000,N_13965,N_13770);
xnor U14001 (N_14001,N_13865,N_13940);
nand U14002 (N_14002,N_13946,N_13851);
and U14003 (N_14003,N_13765,N_13885);
xor U14004 (N_14004,N_13760,N_13921);
nor U14005 (N_14005,N_13862,N_13815);
xnor U14006 (N_14006,N_13780,N_13806);
nor U14007 (N_14007,N_13961,N_13874);
nor U14008 (N_14008,N_13769,N_13838);
nor U14009 (N_14009,N_13812,N_13776);
nand U14010 (N_14010,N_13950,N_13848);
and U14011 (N_14011,N_13841,N_13795);
or U14012 (N_14012,N_13933,N_13924);
or U14013 (N_14013,N_13881,N_13980);
xor U14014 (N_14014,N_13916,N_13782);
xor U14015 (N_14015,N_13875,N_13867);
nand U14016 (N_14016,N_13763,N_13797);
nor U14017 (N_14017,N_13873,N_13831);
nand U14018 (N_14018,N_13998,N_13864);
and U14019 (N_14019,N_13988,N_13836);
xor U14020 (N_14020,N_13963,N_13870);
and U14021 (N_14021,N_13788,N_13810);
xor U14022 (N_14022,N_13943,N_13784);
and U14023 (N_14023,N_13796,N_13964);
nor U14024 (N_14024,N_13759,N_13779);
nand U14025 (N_14025,N_13768,N_13798);
nor U14026 (N_14026,N_13775,N_13945);
and U14027 (N_14027,N_13992,N_13813);
nand U14028 (N_14028,N_13846,N_13871);
and U14029 (N_14029,N_13843,N_13897);
xnor U14030 (N_14030,N_13893,N_13982);
xor U14031 (N_14031,N_13755,N_13936);
or U14032 (N_14032,N_13822,N_13842);
and U14033 (N_14033,N_13762,N_13942);
or U14034 (N_14034,N_13777,N_13994);
or U14035 (N_14035,N_13860,N_13772);
nand U14036 (N_14036,N_13958,N_13971);
nor U14037 (N_14037,N_13941,N_13799);
xnor U14038 (N_14038,N_13800,N_13757);
nor U14039 (N_14039,N_13882,N_13935);
and U14040 (N_14040,N_13978,N_13974);
xnor U14041 (N_14041,N_13884,N_13753);
or U14042 (N_14042,N_13837,N_13844);
xnor U14043 (N_14043,N_13787,N_13826);
nor U14044 (N_14044,N_13794,N_13758);
or U14045 (N_14045,N_13944,N_13807);
or U14046 (N_14046,N_13952,N_13754);
or U14047 (N_14047,N_13766,N_13956);
xor U14048 (N_14048,N_13850,N_13931);
xor U14049 (N_14049,N_13825,N_13990);
or U14050 (N_14050,N_13876,N_13898);
or U14051 (N_14051,N_13902,N_13984);
nor U14052 (N_14052,N_13977,N_13805);
nand U14053 (N_14053,N_13814,N_13987);
and U14054 (N_14054,N_13919,N_13986);
xor U14055 (N_14055,N_13764,N_13778);
or U14056 (N_14056,N_13909,N_13802);
nand U14057 (N_14057,N_13995,N_13756);
nand U14058 (N_14058,N_13892,N_13809);
or U14059 (N_14059,N_13811,N_13890);
xor U14060 (N_14060,N_13790,N_13938);
and U14061 (N_14061,N_13966,N_13953);
nand U14062 (N_14062,N_13923,N_13996);
nand U14063 (N_14063,N_13960,N_13915);
nor U14064 (N_14064,N_13821,N_13832);
and U14065 (N_14065,N_13949,N_13959);
nand U14066 (N_14066,N_13951,N_13981);
nand U14067 (N_14067,N_13819,N_13973);
nor U14068 (N_14068,N_13786,N_13818);
nand U14069 (N_14069,N_13816,N_13847);
and U14070 (N_14070,N_13911,N_13857);
or U14071 (N_14071,N_13912,N_13868);
nand U14072 (N_14072,N_13967,N_13771);
nor U14073 (N_14073,N_13792,N_13789);
nor U14074 (N_14074,N_13920,N_13947);
nand U14075 (N_14075,N_13907,N_13918);
nor U14076 (N_14076,N_13983,N_13903);
nand U14077 (N_14077,N_13781,N_13975);
xor U14078 (N_14078,N_13824,N_13999);
nand U14079 (N_14079,N_13979,N_13888);
nor U14080 (N_14080,N_13853,N_13866);
nor U14081 (N_14081,N_13997,N_13877);
nand U14082 (N_14082,N_13828,N_13955);
nand U14083 (N_14083,N_13803,N_13948);
or U14084 (N_14084,N_13937,N_13957);
and U14085 (N_14085,N_13989,N_13991);
and U14086 (N_14086,N_13968,N_13930);
xor U14087 (N_14087,N_13976,N_13904);
xor U14088 (N_14088,N_13849,N_13913);
nor U14089 (N_14089,N_13908,N_13808);
nor U14090 (N_14090,N_13939,N_13905);
or U14091 (N_14091,N_13927,N_13878);
or U14092 (N_14092,N_13889,N_13854);
nand U14093 (N_14093,N_13886,N_13879);
nor U14094 (N_14094,N_13835,N_13985);
nand U14095 (N_14095,N_13751,N_13773);
xnor U14096 (N_14096,N_13926,N_13829);
or U14097 (N_14097,N_13929,N_13767);
xnor U14098 (N_14098,N_13972,N_13954);
and U14099 (N_14099,N_13969,N_13750);
nand U14100 (N_14100,N_13840,N_13925);
and U14101 (N_14101,N_13906,N_13793);
nand U14102 (N_14102,N_13910,N_13839);
or U14103 (N_14103,N_13901,N_13827);
xor U14104 (N_14104,N_13761,N_13830);
nand U14105 (N_14105,N_13863,N_13922);
xnor U14106 (N_14106,N_13833,N_13887);
nand U14107 (N_14107,N_13914,N_13804);
or U14108 (N_14108,N_13900,N_13962);
and U14109 (N_14109,N_13880,N_13823);
nand U14110 (N_14110,N_13858,N_13932);
xor U14111 (N_14111,N_13783,N_13883);
xnor U14112 (N_14112,N_13820,N_13899);
nor U14113 (N_14113,N_13859,N_13895);
nand U14114 (N_14114,N_13861,N_13752);
xor U14115 (N_14115,N_13970,N_13896);
xnor U14116 (N_14116,N_13917,N_13856);
xnor U14117 (N_14117,N_13872,N_13817);
or U14118 (N_14118,N_13934,N_13834);
and U14119 (N_14119,N_13869,N_13774);
and U14120 (N_14120,N_13791,N_13801);
and U14121 (N_14121,N_13894,N_13928);
or U14122 (N_14122,N_13845,N_13993);
or U14123 (N_14123,N_13855,N_13785);
nor U14124 (N_14124,N_13891,N_13852);
nor U14125 (N_14125,N_13800,N_13977);
and U14126 (N_14126,N_13934,N_13863);
and U14127 (N_14127,N_13776,N_13761);
and U14128 (N_14128,N_13835,N_13950);
or U14129 (N_14129,N_13796,N_13942);
nor U14130 (N_14130,N_13789,N_13945);
xor U14131 (N_14131,N_13865,N_13829);
or U14132 (N_14132,N_13951,N_13855);
xor U14133 (N_14133,N_13965,N_13962);
nor U14134 (N_14134,N_13973,N_13922);
nand U14135 (N_14135,N_13872,N_13942);
or U14136 (N_14136,N_13905,N_13750);
and U14137 (N_14137,N_13769,N_13894);
nor U14138 (N_14138,N_13866,N_13796);
nor U14139 (N_14139,N_13785,N_13943);
and U14140 (N_14140,N_13756,N_13986);
and U14141 (N_14141,N_13843,N_13992);
nor U14142 (N_14142,N_13763,N_13801);
xnor U14143 (N_14143,N_13849,N_13872);
nor U14144 (N_14144,N_13981,N_13945);
and U14145 (N_14145,N_13873,N_13862);
nor U14146 (N_14146,N_13841,N_13899);
and U14147 (N_14147,N_13989,N_13941);
nor U14148 (N_14148,N_13942,N_13972);
xnor U14149 (N_14149,N_13902,N_13890);
nor U14150 (N_14150,N_13867,N_13985);
nand U14151 (N_14151,N_13887,N_13808);
nor U14152 (N_14152,N_13835,N_13926);
and U14153 (N_14153,N_13770,N_13891);
nand U14154 (N_14154,N_13942,N_13812);
xnor U14155 (N_14155,N_13987,N_13760);
xnor U14156 (N_14156,N_13904,N_13891);
nand U14157 (N_14157,N_13985,N_13863);
and U14158 (N_14158,N_13974,N_13869);
and U14159 (N_14159,N_13887,N_13960);
or U14160 (N_14160,N_13786,N_13831);
or U14161 (N_14161,N_13819,N_13965);
and U14162 (N_14162,N_13831,N_13921);
nor U14163 (N_14163,N_13882,N_13905);
xor U14164 (N_14164,N_13831,N_13960);
nor U14165 (N_14165,N_13927,N_13804);
nand U14166 (N_14166,N_13753,N_13988);
nor U14167 (N_14167,N_13952,N_13883);
xor U14168 (N_14168,N_13844,N_13755);
or U14169 (N_14169,N_13902,N_13771);
xor U14170 (N_14170,N_13987,N_13941);
nand U14171 (N_14171,N_13944,N_13892);
and U14172 (N_14172,N_13985,N_13876);
or U14173 (N_14173,N_13950,N_13989);
or U14174 (N_14174,N_13888,N_13926);
or U14175 (N_14175,N_13943,N_13768);
nor U14176 (N_14176,N_13877,N_13928);
xnor U14177 (N_14177,N_13806,N_13791);
or U14178 (N_14178,N_13821,N_13793);
xor U14179 (N_14179,N_13938,N_13990);
or U14180 (N_14180,N_13903,N_13817);
or U14181 (N_14181,N_13922,N_13901);
nor U14182 (N_14182,N_13954,N_13987);
nand U14183 (N_14183,N_13817,N_13878);
or U14184 (N_14184,N_13942,N_13947);
nand U14185 (N_14185,N_13788,N_13942);
and U14186 (N_14186,N_13761,N_13919);
xor U14187 (N_14187,N_13767,N_13843);
nand U14188 (N_14188,N_13752,N_13965);
xnor U14189 (N_14189,N_13955,N_13977);
nor U14190 (N_14190,N_13945,N_13826);
or U14191 (N_14191,N_13826,N_13844);
or U14192 (N_14192,N_13987,N_13824);
or U14193 (N_14193,N_13863,N_13956);
nand U14194 (N_14194,N_13895,N_13856);
nor U14195 (N_14195,N_13886,N_13772);
nand U14196 (N_14196,N_13936,N_13751);
nand U14197 (N_14197,N_13986,N_13828);
nor U14198 (N_14198,N_13979,N_13995);
nand U14199 (N_14199,N_13816,N_13820);
nor U14200 (N_14200,N_13786,N_13761);
or U14201 (N_14201,N_13841,N_13785);
and U14202 (N_14202,N_13757,N_13875);
nor U14203 (N_14203,N_13763,N_13750);
nor U14204 (N_14204,N_13887,N_13894);
nor U14205 (N_14205,N_13753,N_13977);
or U14206 (N_14206,N_13861,N_13965);
nand U14207 (N_14207,N_13927,N_13827);
or U14208 (N_14208,N_13831,N_13887);
and U14209 (N_14209,N_13937,N_13916);
xnor U14210 (N_14210,N_13829,N_13759);
and U14211 (N_14211,N_13900,N_13775);
nand U14212 (N_14212,N_13872,N_13823);
nand U14213 (N_14213,N_13984,N_13997);
or U14214 (N_14214,N_13982,N_13895);
and U14215 (N_14215,N_13910,N_13976);
nand U14216 (N_14216,N_13886,N_13832);
nand U14217 (N_14217,N_13804,N_13911);
and U14218 (N_14218,N_13934,N_13914);
nor U14219 (N_14219,N_13871,N_13910);
and U14220 (N_14220,N_13768,N_13950);
nand U14221 (N_14221,N_13846,N_13833);
and U14222 (N_14222,N_13786,N_13777);
and U14223 (N_14223,N_13801,N_13955);
and U14224 (N_14224,N_13835,N_13833);
nand U14225 (N_14225,N_13876,N_13802);
and U14226 (N_14226,N_13992,N_13972);
nor U14227 (N_14227,N_13939,N_13836);
and U14228 (N_14228,N_13937,N_13930);
xnor U14229 (N_14229,N_13855,N_13857);
nand U14230 (N_14230,N_13816,N_13956);
nor U14231 (N_14231,N_13789,N_13922);
nor U14232 (N_14232,N_13844,N_13876);
xnor U14233 (N_14233,N_13799,N_13844);
nand U14234 (N_14234,N_13979,N_13808);
nand U14235 (N_14235,N_13871,N_13872);
and U14236 (N_14236,N_13841,N_13943);
nand U14237 (N_14237,N_13772,N_13968);
and U14238 (N_14238,N_13846,N_13982);
and U14239 (N_14239,N_13914,N_13911);
xor U14240 (N_14240,N_13880,N_13963);
or U14241 (N_14241,N_13902,N_13981);
xnor U14242 (N_14242,N_13900,N_13975);
and U14243 (N_14243,N_13980,N_13800);
and U14244 (N_14244,N_13820,N_13894);
nand U14245 (N_14245,N_13866,N_13919);
nand U14246 (N_14246,N_13982,N_13979);
nor U14247 (N_14247,N_13970,N_13936);
nor U14248 (N_14248,N_13760,N_13968);
nand U14249 (N_14249,N_13945,N_13752);
xnor U14250 (N_14250,N_14026,N_14027);
or U14251 (N_14251,N_14001,N_14040);
or U14252 (N_14252,N_14245,N_14246);
xor U14253 (N_14253,N_14000,N_14158);
and U14254 (N_14254,N_14038,N_14100);
and U14255 (N_14255,N_14183,N_14065);
xor U14256 (N_14256,N_14248,N_14050);
nand U14257 (N_14257,N_14023,N_14204);
xnor U14258 (N_14258,N_14233,N_14003);
nor U14259 (N_14259,N_14066,N_14009);
xnor U14260 (N_14260,N_14051,N_14139);
xnor U14261 (N_14261,N_14157,N_14120);
nand U14262 (N_14262,N_14002,N_14130);
and U14263 (N_14263,N_14240,N_14239);
and U14264 (N_14264,N_14229,N_14166);
and U14265 (N_14265,N_14008,N_14106);
nand U14266 (N_14266,N_14146,N_14102);
nand U14267 (N_14267,N_14016,N_14036);
nand U14268 (N_14268,N_14188,N_14014);
nor U14269 (N_14269,N_14074,N_14127);
nand U14270 (N_14270,N_14237,N_14232);
or U14271 (N_14271,N_14159,N_14125);
nand U14272 (N_14272,N_14230,N_14020);
xnor U14273 (N_14273,N_14241,N_14111);
or U14274 (N_14274,N_14037,N_14156);
nand U14275 (N_14275,N_14175,N_14199);
xor U14276 (N_14276,N_14164,N_14080);
xor U14277 (N_14277,N_14161,N_14035);
and U14278 (N_14278,N_14082,N_14017);
xnor U14279 (N_14279,N_14151,N_14110);
and U14280 (N_14280,N_14076,N_14195);
or U14281 (N_14281,N_14208,N_14162);
xor U14282 (N_14282,N_14062,N_14047);
or U14283 (N_14283,N_14081,N_14079);
nand U14284 (N_14284,N_14011,N_14213);
nor U14285 (N_14285,N_14217,N_14056);
nor U14286 (N_14286,N_14194,N_14238);
or U14287 (N_14287,N_14150,N_14138);
xnor U14288 (N_14288,N_14168,N_14054);
nor U14289 (N_14289,N_14244,N_14090);
nand U14290 (N_14290,N_14083,N_14205);
and U14291 (N_14291,N_14097,N_14179);
and U14292 (N_14292,N_14032,N_14197);
nand U14293 (N_14293,N_14103,N_14227);
nor U14294 (N_14294,N_14222,N_14058);
or U14295 (N_14295,N_14055,N_14072);
xnor U14296 (N_14296,N_14180,N_14142);
nand U14297 (N_14297,N_14006,N_14200);
nor U14298 (N_14298,N_14007,N_14135);
nand U14299 (N_14299,N_14030,N_14028);
nand U14300 (N_14300,N_14021,N_14201);
and U14301 (N_14301,N_14128,N_14123);
xnor U14302 (N_14302,N_14185,N_14202);
nand U14303 (N_14303,N_14184,N_14088);
or U14304 (N_14304,N_14087,N_14243);
xnor U14305 (N_14305,N_14012,N_14061);
and U14306 (N_14306,N_14131,N_14039);
nor U14307 (N_14307,N_14140,N_14013);
nand U14308 (N_14308,N_14078,N_14136);
or U14309 (N_14309,N_14052,N_14219);
or U14310 (N_14310,N_14206,N_14129);
and U14311 (N_14311,N_14094,N_14022);
or U14312 (N_14312,N_14093,N_14109);
nand U14313 (N_14313,N_14145,N_14034);
nand U14314 (N_14314,N_14141,N_14174);
nor U14315 (N_14315,N_14060,N_14203);
nand U14316 (N_14316,N_14095,N_14249);
or U14317 (N_14317,N_14160,N_14215);
xor U14318 (N_14318,N_14212,N_14067);
xnor U14319 (N_14319,N_14228,N_14163);
nand U14320 (N_14320,N_14224,N_14149);
nor U14321 (N_14321,N_14170,N_14075);
nand U14322 (N_14322,N_14225,N_14107);
and U14323 (N_14323,N_14115,N_14105);
nor U14324 (N_14324,N_14133,N_14144);
or U14325 (N_14325,N_14214,N_14010);
xor U14326 (N_14326,N_14031,N_14155);
nand U14327 (N_14327,N_14046,N_14196);
and U14328 (N_14328,N_14193,N_14218);
or U14329 (N_14329,N_14169,N_14167);
nor U14330 (N_14330,N_14033,N_14154);
and U14331 (N_14331,N_14018,N_14064);
xnor U14332 (N_14332,N_14114,N_14121);
nand U14333 (N_14333,N_14041,N_14220);
xnor U14334 (N_14334,N_14070,N_14104);
nor U14335 (N_14335,N_14148,N_14153);
nand U14336 (N_14336,N_14171,N_14019);
nor U14337 (N_14337,N_14084,N_14147);
xnor U14338 (N_14338,N_14053,N_14210);
nand U14339 (N_14339,N_14118,N_14221);
xor U14340 (N_14340,N_14113,N_14057);
and U14341 (N_14341,N_14226,N_14122);
nor U14342 (N_14342,N_14112,N_14043);
nand U14343 (N_14343,N_14181,N_14042);
nand U14344 (N_14344,N_14132,N_14071);
xnor U14345 (N_14345,N_14152,N_14049);
or U14346 (N_14346,N_14077,N_14207);
nand U14347 (N_14347,N_14092,N_14190);
or U14348 (N_14348,N_14247,N_14124);
xnor U14349 (N_14349,N_14048,N_14211);
nor U14350 (N_14350,N_14191,N_14186);
nand U14351 (N_14351,N_14172,N_14223);
xnor U14352 (N_14352,N_14099,N_14089);
and U14353 (N_14353,N_14209,N_14176);
xnor U14354 (N_14354,N_14216,N_14134);
or U14355 (N_14355,N_14004,N_14068);
nand U14356 (N_14356,N_14024,N_14231);
xor U14357 (N_14357,N_14137,N_14073);
or U14358 (N_14358,N_14091,N_14192);
nand U14359 (N_14359,N_14236,N_14173);
or U14360 (N_14360,N_14059,N_14069);
nor U14361 (N_14361,N_14005,N_14085);
and U14362 (N_14362,N_14234,N_14187);
and U14363 (N_14363,N_14117,N_14235);
nand U14364 (N_14364,N_14143,N_14044);
or U14365 (N_14365,N_14242,N_14182);
nor U14366 (N_14366,N_14098,N_14178);
or U14367 (N_14367,N_14119,N_14029);
or U14368 (N_14368,N_14116,N_14096);
nand U14369 (N_14369,N_14108,N_14101);
nand U14370 (N_14370,N_14025,N_14189);
and U14371 (N_14371,N_14165,N_14045);
nor U14372 (N_14372,N_14198,N_14177);
nand U14373 (N_14373,N_14063,N_14015);
and U14374 (N_14374,N_14126,N_14086);
xor U14375 (N_14375,N_14195,N_14175);
and U14376 (N_14376,N_14217,N_14205);
or U14377 (N_14377,N_14132,N_14158);
and U14378 (N_14378,N_14063,N_14159);
and U14379 (N_14379,N_14145,N_14045);
or U14380 (N_14380,N_14245,N_14239);
xnor U14381 (N_14381,N_14202,N_14058);
and U14382 (N_14382,N_14068,N_14138);
and U14383 (N_14383,N_14240,N_14055);
nand U14384 (N_14384,N_14225,N_14224);
nor U14385 (N_14385,N_14058,N_14067);
nand U14386 (N_14386,N_14002,N_14044);
nand U14387 (N_14387,N_14070,N_14170);
nand U14388 (N_14388,N_14093,N_14089);
and U14389 (N_14389,N_14196,N_14198);
xor U14390 (N_14390,N_14133,N_14179);
and U14391 (N_14391,N_14034,N_14015);
nand U14392 (N_14392,N_14078,N_14203);
or U14393 (N_14393,N_14238,N_14210);
xor U14394 (N_14394,N_14053,N_14230);
nand U14395 (N_14395,N_14084,N_14218);
and U14396 (N_14396,N_14030,N_14061);
xnor U14397 (N_14397,N_14117,N_14180);
and U14398 (N_14398,N_14049,N_14217);
or U14399 (N_14399,N_14038,N_14004);
or U14400 (N_14400,N_14083,N_14012);
nor U14401 (N_14401,N_14187,N_14119);
nor U14402 (N_14402,N_14121,N_14050);
nand U14403 (N_14403,N_14020,N_14118);
nor U14404 (N_14404,N_14199,N_14002);
and U14405 (N_14405,N_14017,N_14163);
or U14406 (N_14406,N_14037,N_14194);
nor U14407 (N_14407,N_14208,N_14176);
nand U14408 (N_14408,N_14207,N_14019);
and U14409 (N_14409,N_14058,N_14069);
and U14410 (N_14410,N_14214,N_14190);
xor U14411 (N_14411,N_14114,N_14133);
xor U14412 (N_14412,N_14091,N_14098);
xor U14413 (N_14413,N_14087,N_14125);
nor U14414 (N_14414,N_14161,N_14222);
and U14415 (N_14415,N_14103,N_14019);
xnor U14416 (N_14416,N_14105,N_14008);
or U14417 (N_14417,N_14147,N_14163);
and U14418 (N_14418,N_14188,N_14229);
nor U14419 (N_14419,N_14102,N_14221);
or U14420 (N_14420,N_14045,N_14176);
xnor U14421 (N_14421,N_14154,N_14128);
and U14422 (N_14422,N_14031,N_14070);
nand U14423 (N_14423,N_14034,N_14104);
and U14424 (N_14424,N_14097,N_14138);
nand U14425 (N_14425,N_14117,N_14194);
nand U14426 (N_14426,N_14200,N_14239);
xnor U14427 (N_14427,N_14190,N_14103);
xnor U14428 (N_14428,N_14234,N_14126);
and U14429 (N_14429,N_14030,N_14043);
and U14430 (N_14430,N_14134,N_14107);
xnor U14431 (N_14431,N_14213,N_14185);
nor U14432 (N_14432,N_14042,N_14013);
nor U14433 (N_14433,N_14057,N_14008);
and U14434 (N_14434,N_14240,N_14188);
or U14435 (N_14435,N_14098,N_14001);
xor U14436 (N_14436,N_14048,N_14051);
nand U14437 (N_14437,N_14007,N_14116);
nand U14438 (N_14438,N_14155,N_14230);
nand U14439 (N_14439,N_14003,N_14226);
and U14440 (N_14440,N_14145,N_14174);
nor U14441 (N_14441,N_14114,N_14184);
nand U14442 (N_14442,N_14128,N_14084);
or U14443 (N_14443,N_14230,N_14067);
and U14444 (N_14444,N_14023,N_14020);
xnor U14445 (N_14445,N_14191,N_14181);
and U14446 (N_14446,N_14145,N_14102);
and U14447 (N_14447,N_14068,N_14077);
nor U14448 (N_14448,N_14228,N_14012);
or U14449 (N_14449,N_14123,N_14191);
or U14450 (N_14450,N_14103,N_14142);
and U14451 (N_14451,N_14220,N_14009);
xor U14452 (N_14452,N_14130,N_14049);
nand U14453 (N_14453,N_14235,N_14214);
xnor U14454 (N_14454,N_14181,N_14173);
or U14455 (N_14455,N_14008,N_14163);
and U14456 (N_14456,N_14188,N_14208);
and U14457 (N_14457,N_14104,N_14151);
and U14458 (N_14458,N_14223,N_14221);
xnor U14459 (N_14459,N_14090,N_14057);
xor U14460 (N_14460,N_14248,N_14217);
nor U14461 (N_14461,N_14067,N_14100);
nor U14462 (N_14462,N_14129,N_14216);
and U14463 (N_14463,N_14182,N_14202);
nand U14464 (N_14464,N_14227,N_14079);
nand U14465 (N_14465,N_14097,N_14213);
or U14466 (N_14466,N_14244,N_14037);
nand U14467 (N_14467,N_14173,N_14107);
nand U14468 (N_14468,N_14083,N_14025);
nand U14469 (N_14469,N_14167,N_14079);
or U14470 (N_14470,N_14039,N_14042);
or U14471 (N_14471,N_14208,N_14018);
nor U14472 (N_14472,N_14075,N_14126);
nor U14473 (N_14473,N_14058,N_14103);
and U14474 (N_14474,N_14003,N_14069);
nand U14475 (N_14475,N_14075,N_14082);
nand U14476 (N_14476,N_14084,N_14241);
or U14477 (N_14477,N_14093,N_14049);
and U14478 (N_14478,N_14198,N_14136);
nand U14479 (N_14479,N_14057,N_14018);
or U14480 (N_14480,N_14226,N_14009);
or U14481 (N_14481,N_14136,N_14021);
and U14482 (N_14482,N_14042,N_14142);
or U14483 (N_14483,N_14200,N_14034);
or U14484 (N_14484,N_14059,N_14217);
nor U14485 (N_14485,N_14207,N_14199);
xnor U14486 (N_14486,N_14204,N_14105);
nand U14487 (N_14487,N_14200,N_14007);
or U14488 (N_14488,N_14112,N_14114);
nand U14489 (N_14489,N_14174,N_14040);
or U14490 (N_14490,N_14011,N_14231);
xnor U14491 (N_14491,N_14098,N_14064);
or U14492 (N_14492,N_14184,N_14249);
or U14493 (N_14493,N_14239,N_14126);
nor U14494 (N_14494,N_14020,N_14016);
nand U14495 (N_14495,N_14132,N_14225);
nor U14496 (N_14496,N_14231,N_14052);
and U14497 (N_14497,N_14083,N_14124);
and U14498 (N_14498,N_14219,N_14044);
nor U14499 (N_14499,N_14175,N_14054);
nor U14500 (N_14500,N_14310,N_14450);
xnor U14501 (N_14501,N_14272,N_14344);
nor U14502 (N_14502,N_14297,N_14423);
nor U14503 (N_14503,N_14427,N_14417);
or U14504 (N_14504,N_14313,N_14488);
nor U14505 (N_14505,N_14448,N_14314);
and U14506 (N_14506,N_14452,N_14362);
xnor U14507 (N_14507,N_14279,N_14353);
or U14508 (N_14508,N_14357,N_14393);
or U14509 (N_14509,N_14443,N_14411);
and U14510 (N_14510,N_14253,N_14296);
xnor U14511 (N_14511,N_14375,N_14311);
xnor U14512 (N_14512,N_14390,N_14456);
or U14513 (N_14513,N_14333,N_14460);
xor U14514 (N_14514,N_14259,N_14276);
xor U14515 (N_14515,N_14415,N_14338);
or U14516 (N_14516,N_14435,N_14261);
xor U14517 (N_14517,N_14485,N_14410);
xor U14518 (N_14518,N_14315,N_14336);
and U14519 (N_14519,N_14434,N_14391);
and U14520 (N_14520,N_14422,N_14479);
xor U14521 (N_14521,N_14408,N_14492);
nor U14522 (N_14522,N_14342,N_14358);
xnor U14523 (N_14523,N_14439,N_14378);
and U14524 (N_14524,N_14477,N_14283);
nor U14525 (N_14525,N_14449,N_14286);
and U14526 (N_14526,N_14447,N_14453);
nor U14527 (N_14527,N_14458,N_14473);
or U14528 (N_14528,N_14441,N_14379);
xnor U14529 (N_14529,N_14305,N_14316);
and U14530 (N_14530,N_14429,N_14425);
xor U14531 (N_14531,N_14308,N_14367);
nand U14532 (N_14532,N_14377,N_14294);
xor U14533 (N_14533,N_14468,N_14349);
xnor U14534 (N_14534,N_14476,N_14293);
xnor U14535 (N_14535,N_14494,N_14273);
nor U14536 (N_14536,N_14269,N_14373);
or U14537 (N_14537,N_14480,N_14266);
or U14538 (N_14538,N_14251,N_14376);
and U14539 (N_14539,N_14481,N_14389);
nor U14540 (N_14540,N_14442,N_14304);
nand U14541 (N_14541,N_14351,N_14454);
xnor U14542 (N_14542,N_14312,N_14431);
or U14543 (N_14543,N_14264,N_14356);
nor U14544 (N_14544,N_14256,N_14420);
and U14545 (N_14545,N_14354,N_14385);
nand U14546 (N_14546,N_14307,N_14360);
xor U14547 (N_14547,N_14252,N_14372);
nor U14548 (N_14548,N_14254,N_14430);
and U14549 (N_14549,N_14483,N_14399);
nor U14550 (N_14550,N_14306,N_14370);
or U14551 (N_14551,N_14298,N_14498);
and U14552 (N_14552,N_14486,N_14416);
or U14553 (N_14553,N_14386,N_14278);
nand U14554 (N_14554,N_14255,N_14263);
xnor U14555 (N_14555,N_14405,N_14409);
nor U14556 (N_14556,N_14265,N_14395);
nand U14557 (N_14557,N_14368,N_14328);
and U14558 (N_14558,N_14401,N_14400);
nand U14559 (N_14559,N_14414,N_14499);
nand U14560 (N_14560,N_14406,N_14471);
xnor U14561 (N_14561,N_14365,N_14490);
and U14562 (N_14562,N_14267,N_14484);
or U14563 (N_14563,N_14496,N_14466);
xor U14564 (N_14564,N_14280,N_14436);
xor U14565 (N_14565,N_14418,N_14274);
nor U14566 (N_14566,N_14327,N_14331);
nor U14567 (N_14567,N_14388,N_14432);
or U14568 (N_14568,N_14352,N_14455);
nor U14569 (N_14569,N_14438,N_14285);
xor U14570 (N_14570,N_14318,N_14421);
nor U14571 (N_14571,N_14281,N_14426);
nor U14572 (N_14572,N_14299,N_14482);
and U14573 (N_14573,N_14445,N_14282);
or U14574 (N_14574,N_14369,N_14487);
or U14575 (N_14575,N_14295,N_14364);
nand U14576 (N_14576,N_14433,N_14347);
nand U14577 (N_14577,N_14465,N_14382);
and U14578 (N_14578,N_14384,N_14444);
nand U14579 (N_14579,N_14371,N_14301);
nor U14580 (N_14580,N_14300,N_14497);
xor U14581 (N_14581,N_14330,N_14309);
and U14582 (N_14582,N_14335,N_14459);
or U14583 (N_14583,N_14403,N_14463);
nand U14584 (N_14584,N_14345,N_14341);
or U14585 (N_14585,N_14437,N_14329);
nand U14586 (N_14586,N_14350,N_14260);
or U14587 (N_14587,N_14419,N_14323);
xnor U14588 (N_14588,N_14340,N_14413);
nand U14589 (N_14589,N_14320,N_14287);
and U14590 (N_14590,N_14343,N_14334);
nand U14591 (N_14591,N_14457,N_14493);
or U14592 (N_14592,N_14317,N_14464);
and U14593 (N_14593,N_14398,N_14346);
nand U14594 (N_14594,N_14292,N_14491);
or U14595 (N_14595,N_14363,N_14348);
nand U14596 (N_14596,N_14404,N_14451);
and U14597 (N_14597,N_14470,N_14475);
nor U14598 (N_14598,N_14277,N_14289);
or U14599 (N_14599,N_14284,N_14472);
xnor U14600 (N_14600,N_14489,N_14268);
or U14601 (N_14601,N_14325,N_14339);
nor U14602 (N_14602,N_14397,N_14361);
xor U14603 (N_14603,N_14250,N_14303);
and U14604 (N_14604,N_14467,N_14359);
xor U14605 (N_14605,N_14302,N_14322);
nor U14606 (N_14606,N_14412,N_14258);
nand U14607 (N_14607,N_14461,N_14387);
and U14608 (N_14608,N_14321,N_14440);
xor U14609 (N_14609,N_14478,N_14394);
nor U14610 (N_14610,N_14271,N_14402);
nand U14611 (N_14611,N_14383,N_14270);
nand U14612 (N_14612,N_14291,N_14366);
and U14613 (N_14613,N_14290,N_14462);
nor U14614 (N_14614,N_14262,N_14332);
xnor U14615 (N_14615,N_14374,N_14474);
and U14616 (N_14616,N_14337,N_14257);
or U14617 (N_14617,N_14326,N_14324);
xnor U14618 (N_14618,N_14392,N_14380);
nor U14619 (N_14619,N_14424,N_14469);
nand U14620 (N_14620,N_14319,N_14428);
nand U14621 (N_14621,N_14288,N_14495);
nand U14622 (N_14622,N_14407,N_14446);
or U14623 (N_14623,N_14396,N_14355);
nor U14624 (N_14624,N_14381,N_14275);
or U14625 (N_14625,N_14324,N_14372);
nand U14626 (N_14626,N_14478,N_14447);
nor U14627 (N_14627,N_14297,N_14438);
nor U14628 (N_14628,N_14340,N_14395);
nand U14629 (N_14629,N_14419,N_14293);
nor U14630 (N_14630,N_14389,N_14341);
xor U14631 (N_14631,N_14367,N_14481);
and U14632 (N_14632,N_14265,N_14253);
and U14633 (N_14633,N_14411,N_14307);
nand U14634 (N_14634,N_14353,N_14478);
xor U14635 (N_14635,N_14382,N_14480);
and U14636 (N_14636,N_14321,N_14480);
xor U14637 (N_14637,N_14481,N_14350);
and U14638 (N_14638,N_14397,N_14314);
or U14639 (N_14639,N_14445,N_14358);
xor U14640 (N_14640,N_14356,N_14417);
nand U14641 (N_14641,N_14291,N_14377);
and U14642 (N_14642,N_14295,N_14486);
nand U14643 (N_14643,N_14261,N_14290);
nand U14644 (N_14644,N_14420,N_14301);
and U14645 (N_14645,N_14332,N_14382);
or U14646 (N_14646,N_14379,N_14250);
nor U14647 (N_14647,N_14426,N_14360);
nand U14648 (N_14648,N_14387,N_14342);
or U14649 (N_14649,N_14409,N_14363);
or U14650 (N_14650,N_14432,N_14410);
xnor U14651 (N_14651,N_14464,N_14258);
or U14652 (N_14652,N_14479,N_14296);
or U14653 (N_14653,N_14471,N_14360);
nand U14654 (N_14654,N_14435,N_14346);
or U14655 (N_14655,N_14410,N_14289);
nand U14656 (N_14656,N_14364,N_14379);
nand U14657 (N_14657,N_14303,N_14278);
nand U14658 (N_14658,N_14469,N_14344);
xnor U14659 (N_14659,N_14325,N_14263);
xnor U14660 (N_14660,N_14266,N_14377);
nand U14661 (N_14661,N_14327,N_14381);
and U14662 (N_14662,N_14443,N_14433);
nor U14663 (N_14663,N_14257,N_14381);
and U14664 (N_14664,N_14297,N_14474);
xor U14665 (N_14665,N_14424,N_14413);
nand U14666 (N_14666,N_14298,N_14491);
or U14667 (N_14667,N_14436,N_14310);
and U14668 (N_14668,N_14418,N_14257);
nor U14669 (N_14669,N_14498,N_14434);
nand U14670 (N_14670,N_14445,N_14363);
nor U14671 (N_14671,N_14428,N_14450);
nor U14672 (N_14672,N_14413,N_14266);
nor U14673 (N_14673,N_14410,N_14371);
nand U14674 (N_14674,N_14303,N_14391);
or U14675 (N_14675,N_14385,N_14375);
xnor U14676 (N_14676,N_14459,N_14339);
nand U14677 (N_14677,N_14368,N_14393);
or U14678 (N_14678,N_14450,N_14429);
nor U14679 (N_14679,N_14290,N_14496);
nand U14680 (N_14680,N_14315,N_14478);
and U14681 (N_14681,N_14328,N_14391);
nand U14682 (N_14682,N_14446,N_14431);
xnor U14683 (N_14683,N_14381,N_14365);
or U14684 (N_14684,N_14274,N_14283);
nor U14685 (N_14685,N_14274,N_14368);
or U14686 (N_14686,N_14301,N_14267);
xor U14687 (N_14687,N_14498,N_14323);
xor U14688 (N_14688,N_14258,N_14375);
and U14689 (N_14689,N_14394,N_14491);
nand U14690 (N_14690,N_14495,N_14292);
nor U14691 (N_14691,N_14409,N_14420);
nor U14692 (N_14692,N_14265,N_14463);
xnor U14693 (N_14693,N_14346,N_14464);
and U14694 (N_14694,N_14438,N_14331);
or U14695 (N_14695,N_14359,N_14383);
nand U14696 (N_14696,N_14454,N_14464);
and U14697 (N_14697,N_14303,N_14309);
and U14698 (N_14698,N_14287,N_14347);
xnor U14699 (N_14699,N_14304,N_14317);
or U14700 (N_14700,N_14304,N_14453);
and U14701 (N_14701,N_14353,N_14416);
or U14702 (N_14702,N_14261,N_14483);
or U14703 (N_14703,N_14261,N_14455);
xnor U14704 (N_14704,N_14489,N_14460);
xnor U14705 (N_14705,N_14379,N_14283);
nand U14706 (N_14706,N_14487,N_14442);
nand U14707 (N_14707,N_14363,N_14327);
and U14708 (N_14708,N_14269,N_14390);
or U14709 (N_14709,N_14439,N_14337);
or U14710 (N_14710,N_14351,N_14313);
and U14711 (N_14711,N_14364,N_14292);
nand U14712 (N_14712,N_14333,N_14289);
nor U14713 (N_14713,N_14322,N_14457);
and U14714 (N_14714,N_14292,N_14254);
nand U14715 (N_14715,N_14322,N_14351);
nand U14716 (N_14716,N_14494,N_14487);
nor U14717 (N_14717,N_14408,N_14257);
xnor U14718 (N_14718,N_14284,N_14346);
nand U14719 (N_14719,N_14430,N_14366);
nor U14720 (N_14720,N_14465,N_14295);
nor U14721 (N_14721,N_14380,N_14252);
nor U14722 (N_14722,N_14272,N_14369);
nand U14723 (N_14723,N_14315,N_14394);
and U14724 (N_14724,N_14261,N_14420);
or U14725 (N_14725,N_14347,N_14463);
xnor U14726 (N_14726,N_14407,N_14267);
and U14727 (N_14727,N_14271,N_14451);
xnor U14728 (N_14728,N_14314,N_14279);
or U14729 (N_14729,N_14354,N_14282);
nand U14730 (N_14730,N_14489,N_14331);
xor U14731 (N_14731,N_14347,N_14320);
nand U14732 (N_14732,N_14265,N_14377);
nor U14733 (N_14733,N_14252,N_14434);
and U14734 (N_14734,N_14495,N_14431);
xor U14735 (N_14735,N_14429,N_14331);
nor U14736 (N_14736,N_14421,N_14468);
or U14737 (N_14737,N_14401,N_14467);
or U14738 (N_14738,N_14332,N_14388);
or U14739 (N_14739,N_14368,N_14436);
xor U14740 (N_14740,N_14373,N_14339);
xnor U14741 (N_14741,N_14273,N_14389);
nand U14742 (N_14742,N_14328,N_14324);
xnor U14743 (N_14743,N_14344,N_14307);
xnor U14744 (N_14744,N_14387,N_14315);
nor U14745 (N_14745,N_14380,N_14298);
nor U14746 (N_14746,N_14394,N_14253);
and U14747 (N_14747,N_14429,N_14452);
or U14748 (N_14748,N_14315,N_14426);
nand U14749 (N_14749,N_14315,N_14347);
or U14750 (N_14750,N_14597,N_14748);
xor U14751 (N_14751,N_14673,N_14687);
and U14752 (N_14752,N_14618,N_14532);
xnor U14753 (N_14753,N_14543,N_14645);
nor U14754 (N_14754,N_14571,N_14516);
and U14755 (N_14755,N_14667,N_14518);
nor U14756 (N_14756,N_14739,N_14521);
or U14757 (N_14757,N_14648,N_14575);
or U14758 (N_14758,N_14515,N_14669);
or U14759 (N_14759,N_14555,N_14573);
and U14760 (N_14760,N_14632,N_14698);
nor U14761 (N_14761,N_14599,N_14585);
or U14762 (N_14762,N_14552,N_14732);
xnor U14763 (N_14763,N_14701,N_14694);
and U14764 (N_14764,N_14660,N_14564);
xor U14765 (N_14765,N_14579,N_14595);
and U14766 (N_14766,N_14593,N_14628);
xnor U14767 (N_14767,N_14617,N_14512);
or U14768 (N_14768,N_14592,N_14630);
xor U14769 (N_14769,N_14717,N_14727);
or U14770 (N_14770,N_14554,N_14661);
nor U14771 (N_14771,N_14629,N_14637);
and U14772 (N_14772,N_14635,N_14640);
nand U14773 (N_14773,N_14627,N_14547);
nand U14774 (N_14774,N_14722,N_14605);
and U14775 (N_14775,N_14685,N_14746);
and U14776 (N_14776,N_14590,N_14689);
nor U14777 (N_14777,N_14691,N_14562);
or U14778 (N_14778,N_14638,N_14743);
and U14779 (N_14779,N_14507,N_14613);
xor U14780 (N_14780,N_14559,N_14536);
nand U14781 (N_14781,N_14692,N_14680);
or U14782 (N_14782,N_14504,N_14622);
and U14783 (N_14783,N_14601,N_14671);
nor U14784 (N_14784,N_14744,N_14568);
xor U14785 (N_14785,N_14674,N_14533);
xor U14786 (N_14786,N_14639,N_14738);
or U14787 (N_14787,N_14662,N_14584);
or U14788 (N_14788,N_14610,N_14724);
or U14789 (N_14789,N_14608,N_14656);
and U14790 (N_14790,N_14723,N_14670);
nor U14791 (N_14791,N_14733,N_14578);
xnor U14792 (N_14792,N_14659,N_14587);
nor U14793 (N_14793,N_14567,N_14560);
and U14794 (N_14794,N_14730,N_14545);
nand U14795 (N_14795,N_14588,N_14658);
nor U14796 (N_14796,N_14591,N_14650);
nor U14797 (N_14797,N_14598,N_14594);
nor U14798 (N_14798,N_14557,N_14683);
or U14799 (N_14799,N_14647,N_14527);
nor U14800 (N_14800,N_14528,N_14719);
xor U14801 (N_14801,N_14529,N_14586);
nand U14802 (N_14802,N_14621,N_14684);
nor U14803 (N_14803,N_14700,N_14654);
xnor U14804 (N_14804,N_14542,N_14742);
nand U14805 (N_14805,N_14574,N_14718);
or U14806 (N_14806,N_14693,N_14500);
xor U14807 (N_14807,N_14737,N_14703);
and U14808 (N_14808,N_14537,N_14709);
nor U14809 (N_14809,N_14561,N_14609);
nor U14810 (N_14810,N_14556,N_14634);
or U14811 (N_14811,N_14651,N_14678);
or U14812 (N_14812,N_14710,N_14626);
nor U14813 (N_14813,N_14525,N_14600);
nor U14814 (N_14814,N_14620,N_14688);
nand U14815 (N_14815,N_14524,N_14668);
and U14816 (N_14816,N_14539,N_14704);
and U14817 (N_14817,N_14505,N_14546);
and U14818 (N_14818,N_14679,N_14540);
xor U14819 (N_14819,N_14569,N_14675);
xor U14820 (N_14820,N_14577,N_14713);
or U14821 (N_14821,N_14663,N_14642);
and U14822 (N_14822,N_14501,N_14614);
nand U14823 (N_14823,N_14511,N_14538);
and U14824 (N_14824,N_14548,N_14623);
and U14825 (N_14825,N_14517,N_14535);
nand U14826 (N_14826,N_14696,N_14705);
and U14827 (N_14827,N_14657,N_14697);
xnor U14828 (N_14828,N_14712,N_14558);
and U14829 (N_14829,N_14611,N_14625);
xor U14830 (N_14830,N_14690,N_14513);
or U14831 (N_14831,N_14682,N_14519);
xnor U14832 (N_14832,N_14522,N_14606);
nor U14833 (N_14833,N_14509,N_14503);
nand U14834 (N_14834,N_14716,N_14602);
nand U14835 (N_14835,N_14714,N_14666);
nor U14836 (N_14836,N_14523,N_14665);
xor U14837 (N_14837,N_14583,N_14589);
nor U14838 (N_14838,N_14725,N_14664);
nand U14839 (N_14839,N_14653,N_14646);
xnor U14840 (N_14840,N_14566,N_14550);
xor U14841 (N_14841,N_14576,N_14728);
nand U14842 (N_14842,N_14736,N_14749);
xor U14843 (N_14843,N_14508,N_14715);
nor U14844 (N_14844,N_14652,N_14740);
xnor U14845 (N_14845,N_14551,N_14735);
or U14846 (N_14846,N_14636,N_14530);
or U14847 (N_14847,N_14544,N_14686);
and U14848 (N_14848,N_14570,N_14526);
and U14849 (N_14849,N_14707,N_14506);
or U14850 (N_14850,N_14607,N_14514);
and U14851 (N_14851,N_14582,N_14615);
nand U14852 (N_14852,N_14711,N_14729);
nand U14853 (N_14853,N_14619,N_14624);
and U14854 (N_14854,N_14534,N_14720);
nor U14855 (N_14855,N_14649,N_14731);
nor U14856 (N_14856,N_14531,N_14616);
and U14857 (N_14857,N_14677,N_14641);
xor U14858 (N_14858,N_14672,N_14596);
nand U14859 (N_14859,N_14565,N_14510);
nand U14860 (N_14860,N_14581,N_14695);
and U14861 (N_14861,N_14745,N_14734);
or U14862 (N_14862,N_14541,N_14563);
nor U14863 (N_14863,N_14676,N_14603);
nand U14864 (N_14864,N_14553,N_14502);
or U14865 (N_14865,N_14643,N_14699);
and U14866 (N_14866,N_14702,N_14655);
or U14867 (N_14867,N_14726,N_14520);
xnor U14868 (N_14868,N_14631,N_14708);
or U14869 (N_14869,N_14612,N_14741);
and U14870 (N_14870,N_14747,N_14580);
and U14871 (N_14871,N_14681,N_14706);
nor U14872 (N_14872,N_14572,N_14549);
nor U14873 (N_14873,N_14721,N_14633);
or U14874 (N_14874,N_14644,N_14604);
or U14875 (N_14875,N_14725,N_14502);
nand U14876 (N_14876,N_14656,N_14610);
nand U14877 (N_14877,N_14717,N_14675);
nand U14878 (N_14878,N_14652,N_14674);
nor U14879 (N_14879,N_14699,N_14634);
nor U14880 (N_14880,N_14526,N_14707);
nand U14881 (N_14881,N_14693,N_14605);
xor U14882 (N_14882,N_14528,N_14727);
or U14883 (N_14883,N_14562,N_14702);
or U14884 (N_14884,N_14666,N_14712);
or U14885 (N_14885,N_14549,N_14521);
and U14886 (N_14886,N_14716,N_14508);
nand U14887 (N_14887,N_14547,N_14512);
nor U14888 (N_14888,N_14629,N_14551);
or U14889 (N_14889,N_14672,N_14645);
or U14890 (N_14890,N_14740,N_14603);
xnor U14891 (N_14891,N_14740,N_14634);
or U14892 (N_14892,N_14510,N_14584);
or U14893 (N_14893,N_14581,N_14604);
and U14894 (N_14894,N_14631,N_14672);
nand U14895 (N_14895,N_14512,N_14710);
and U14896 (N_14896,N_14589,N_14637);
xnor U14897 (N_14897,N_14589,N_14554);
nand U14898 (N_14898,N_14517,N_14654);
and U14899 (N_14899,N_14530,N_14716);
and U14900 (N_14900,N_14657,N_14638);
nor U14901 (N_14901,N_14649,N_14739);
and U14902 (N_14902,N_14681,N_14644);
or U14903 (N_14903,N_14681,N_14626);
nand U14904 (N_14904,N_14650,N_14514);
nor U14905 (N_14905,N_14536,N_14701);
nand U14906 (N_14906,N_14544,N_14572);
and U14907 (N_14907,N_14604,N_14584);
nor U14908 (N_14908,N_14631,N_14573);
or U14909 (N_14909,N_14715,N_14563);
and U14910 (N_14910,N_14500,N_14718);
xnor U14911 (N_14911,N_14588,N_14630);
nand U14912 (N_14912,N_14739,N_14683);
or U14913 (N_14913,N_14656,N_14624);
nand U14914 (N_14914,N_14619,N_14676);
and U14915 (N_14915,N_14588,N_14616);
and U14916 (N_14916,N_14676,N_14548);
or U14917 (N_14917,N_14731,N_14692);
nor U14918 (N_14918,N_14529,N_14631);
nand U14919 (N_14919,N_14640,N_14519);
xnor U14920 (N_14920,N_14520,N_14587);
nor U14921 (N_14921,N_14595,N_14628);
nand U14922 (N_14922,N_14548,N_14564);
nor U14923 (N_14923,N_14558,N_14647);
nand U14924 (N_14924,N_14509,N_14621);
nor U14925 (N_14925,N_14553,N_14570);
or U14926 (N_14926,N_14536,N_14620);
xor U14927 (N_14927,N_14719,N_14546);
and U14928 (N_14928,N_14667,N_14544);
and U14929 (N_14929,N_14502,N_14713);
or U14930 (N_14930,N_14530,N_14724);
or U14931 (N_14931,N_14655,N_14544);
or U14932 (N_14932,N_14568,N_14666);
nor U14933 (N_14933,N_14618,N_14742);
nand U14934 (N_14934,N_14544,N_14573);
nor U14935 (N_14935,N_14578,N_14507);
nor U14936 (N_14936,N_14597,N_14589);
nor U14937 (N_14937,N_14708,N_14659);
or U14938 (N_14938,N_14731,N_14723);
xnor U14939 (N_14939,N_14503,N_14746);
xor U14940 (N_14940,N_14578,N_14738);
xor U14941 (N_14941,N_14508,N_14745);
nand U14942 (N_14942,N_14717,N_14633);
or U14943 (N_14943,N_14549,N_14696);
nand U14944 (N_14944,N_14668,N_14641);
nor U14945 (N_14945,N_14597,N_14543);
nor U14946 (N_14946,N_14603,N_14708);
xnor U14947 (N_14947,N_14627,N_14745);
nand U14948 (N_14948,N_14671,N_14605);
or U14949 (N_14949,N_14533,N_14564);
nor U14950 (N_14950,N_14620,N_14531);
or U14951 (N_14951,N_14669,N_14749);
xnor U14952 (N_14952,N_14611,N_14506);
xnor U14953 (N_14953,N_14555,N_14598);
nor U14954 (N_14954,N_14560,N_14616);
nand U14955 (N_14955,N_14575,N_14555);
nor U14956 (N_14956,N_14615,N_14690);
or U14957 (N_14957,N_14680,N_14685);
and U14958 (N_14958,N_14567,N_14531);
nor U14959 (N_14959,N_14617,N_14528);
or U14960 (N_14960,N_14675,N_14508);
or U14961 (N_14961,N_14648,N_14637);
nor U14962 (N_14962,N_14732,N_14705);
or U14963 (N_14963,N_14600,N_14530);
xnor U14964 (N_14964,N_14532,N_14515);
nand U14965 (N_14965,N_14720,N_14570);
and U14966 (N_14966,N_14652,N_14667);
nand U14967 (N_14967,N_14514,N_14510);
or U14968 (N_14968,N_14633,N_14526);
xnor U14969 (N_14969,N_14628,N_14656);
xnor U14970 (N_14970,N_14599,N_14579);
xnor U14971 (N_14971,N_14519,N_14575);
or U14972 (N_14972,N_14640,N_14699);
xor U14973 (N_14973,N_14722,N_14729);
xor U14974 (N_14974,N_14549,N_14707);
or U14975 (N_14975,N_14532,N_14631);
or U14976 (N_14976,N_14561,N_14547);
xnor U14977 (N_14977,N_14528,N_14609);
nand U14978 (N_14978,N_14632,N_14695);
and U14979 (N_14979,N_14596,N_14662);
nand U14980 (N_14980,N_14633,N_14587);
xor U14981 (N_14981,N_14605,N_14586);
nor U14982 (N_14982,N_14625,N_14569);
and U14983 (N_14983,N_14554,N_14515);
xnor U14984 (N_14984,N_14555,N_14504);
or U14985 (N_14985,N_14589,N_14503);
or U14986 (N_14986,N_14668,N_14560);
and U14987 (N_14987,N_14524,N_14516);
nand U14988 (N_14988,N_14528,N_14637);
nand U14989 (N_14989,N_14633,N_14703);
xor U14990 (N_14990,N_14514,N_14528);
or U14991 (N_14991,N_14656,N_14663);
nor U14992 (N_14992,N_14608,N_14563);
and U14993 (N_14993,N_14693,N_14720);
xnor U14994 (N_14994,N_14670,N_14639);
or U14995 (N_14995,N_14721,N_14640);
nand U14996 (N_14996,N_14577,N_14547);
and U14997 (N_14997,N_14694,N_14644);
xor U14998 (N_14998,N_14562,N_14503);
xor U14999 (N_14999,N_14642,N_14720);
and UO_0 (O_0,N_14951,N_14932);
nand UO_1 (O_1,N_14929,N_14906);
and UO_2 (O_2,N_14859,N_14977);
or UO_3 (O_3,N_14769,N_14910);
xor UO_4 (O_4,N_14795,N_14894);
nor UO_5 (O_5,N_14899,N_14781);
nand UO_6 (O_6,N_14927,N_14863);
nor UO_7 (O_7,N_14780,N_14819);
or UO_8 (O_8,N_14760,N_14778);
and UO_9 (O_9,N_14913,N_14771);
nor UO_10 (O_10,N_14980,N_14975);
and UO_11 (O_11,N_14971,N_14855);
nand UO_12 (O_12,N_14974,N_14846);
or UO_13 (O_13,N_14959,N_14821);
and UO_14 (O_14,N_14897,N_14948);
xor UO_15 (O_15,N_14814,N_14753);
nor UO_16 (O_16,N_14824,N_14890);
nor UO_17 (O_17,N_14915,N_14788);
nor UO_18 (O_18,N_14963,N_14923);
or UO_19 (O_19,N_14979,N_14871);
and UO_20 (O_20,N_14793,N_14972);
xnor UO_21 (O_21,N_14849,N_14916);
nand UO_22 (O_22,N_14834,N_14931);
nand UO_23 (O_23,N_14990,N_14961);
xor UO_24 (O_24,N_14955,N_14998);
and UO_25 (O_25,N_14767,N_14904);
xor UO_26 (O_26,N_14988,N_14991);
xor UO_27 (O_27,N_14752,N_14872);
or UO_28 (O_28,N_14909,N_14791);
nor UO_29 (O_29,N_14789,N_14784);
nand UO_30 (O_30,N_14763,N_14861);
xor UO_31 (O_31,N_14981,N_14987);
nor UO_32 (O_32,N_14937,N_14908);
nand UO_33 (O_33,N_14914,N_14919);
nand UO_34 (O_34,N_14857,N_14982);
nor UO_35 (O_35,N_14757,N_14946);
or UO_36 (O_36,N_14842,N_14964);
xnor UO_37 (O_37,N_14833,N_14817);
nand UO_38 (O_38,N_14844,N_14902);
xnor UO_39 (O_39,N_14862,N_14841);
and UO_40 (O_40,N_14802,N_14877);
nand UO_41 (O_41,N_14969,N_14870);
or UO_42 (O_42,N_14815,N_14797);
and UO_43 (O_43,N_14764,N_14756);
or UO_44 (O_44,N_14809,N_14896);
xnor UO_45 (O_45,N_14886,N_14918);
or UO_46 (O_46,N_14792,N_14989);
nor UO_47 (O_47,N_14912,N_14885);
xnor UO_48 (O_48,N_14820,N_14806);
and UO_49 (O_49,N_14776,N_14807);
nor UO_50 (O_50,N_14901,N_14957);
nand UO_51 (O_51,N_14947,N_14852);
or UO_52 (O_52,N_14828,N_14984);
and UO_53 (O_53,N_14958,N_14829);
xnor UO_54 (O_54,N_14926,N_14813);
xor UO_55 (O_55,N_14751,N_14907);
nand UO_56 (O_56,N_14836,N_14935);
xor UO_57 (O_57,N_14920,N_14911);
or UO_58 (O_58,N_14953,N_14892);
nor UO_59 (O_59,N_14798,N_14850);
nand UO_60 (O_60,N_14879,N_14888);
or UO_61 (O_61,N_14876,N_14826);
or UO_62 (O_62,N_14823,N_14925);
nor UO_63 (O_63,N_14867,N_14924);
nand UO_64 (O_64,N_14875,N_14889);
nor UO_65 (O_65,N_14851,N_14801);
or UO_66 (O_66,N_14864,N_14930);
nand UO_67 (O_67,N_14993,N_14996);
xnor UO_68 (O_68,N_14785,N_14754);
nor UO_69 (O_69,N_14810,N_14874);
or UO_70 (O_70,N_14803,N_14856);
and UO_71 (O_71,N_14995,N_14800);
nor UO_72 (O_72,N_14787,N_14816);
nor UO_73 (O_73,N_14811,N_14835);
xor UO_74 (O_74,N_14891,N_14766);
or UO_75 (O_75,N_14860,N_14922);
xor UO_76 (O_76,N_14942,N_14873);
and UO_77 (O_77,N_14950,N_14818);
xnor UO_78 (O_78,N_14962,N_14866);
nand UO_79 (O_79,N_14893,N_14858);
or UO_80 (O_80,N_14822,N_14847);
xnor UO_81 (O_81,N_14887,N_14956);
nor UO_82 (O_82,N_14772,N_14936);
nand UO_83 (O_83,N_14898,N_14978);
nor UO_84 (O_84,N_14884,N_14805);
xor UO_85 (O_85,N_14917,N_14796);
and UO_86 (O_86,N_14999,N_14790);
nor UO_87 (O_87,N_14967,N_14952);
nand UO_88 (O_88,N_14768,N_14944);
nand UO_89 (O_89,N_14994,N_14997);
xnor UO_90 (O_90,N_14779,N_14928);
nor UO_91 (O_91,N_14903,N_14882);
or UO_92 (O_92,N_14848,N_14837);
nor UO_93 (O_93,N_14883,N_14970);
or UO_94 (O_94,N_14869,N_14905);
nor UO_95 (O_95,N_14878,N_14939);
nor UO_96 (O_96,N_14976,N_14825);
or UO_97 (O_97,N_14943,N_14945);
nand UO_98 (O_98,N_14880,N_14949);
nor UO_99 (O_99,N_14966,N_14934);
and UO_100 (O_100,N_14759,N_14960);
nand UO_101 (O_101,N_14831,N_14983);
and UO_102 (O_102,N_14933,N_14765);
nor UO_103 (O_103,N_14808,N_14799);
nor UO_104 (O_104,N_14786,N_14954);
xor UO_105 (O_105,N_14868,N_14986);
nand UO_106 (O_106,N_14865,N_14938);
and UO_107 (O_107,N_14853,N_14783);
nand UO_108 (O_108,N_14992,N_14832);
nand UO_109 (O_109,N_14845,N_14774);
nand UO_110 (O_110,N_14843,N_14900);
nand UO_111 (O_111,N_14777,N_14755);
nor UO_112 (O_112,N_14854,N_14773);
xnor UO_113 (O_113,N_14782,N_14881);
xnor UO_114 (O_114,N_14838,N_14794);
and UO_115 (O_115,N_14968,N_14985);
nor UO_116 (O_116,N_14758,N_14895);
nand UO_117 (O_117,N_14750,N_14761);
and UO_118 (O_118,N_14762,N_14827);
nand UO_119 (O_119,N_14830,N_14812);
and UO_120 (O_120,N_14941,N_14921);
and UO_121 (O_121,N_14965,N_14839);
nand UO_122 (O_122,N_14840,N_14775);
nand UO_123 (O_123,N_14804,N_14770);
xnor UO_124 (O_124,N_14973,N_14940);
or UO_125 (O_125,N_14787,N_14970);
xor UO_126 (O_126,N_14977,N_14885);
nor UO_127 (O_127,N_14778,N_14882);
and UO_128 (O_128,N_14850,N_14945);
or UO_129 (O_129,N_14881,N_14764);
and UO_130 (O_130,N_14817,N_14951);
or UO_131 (O_131,N_14882,N_14967);
xor UO_132 (O_132,N_14914,N_14790);
xor UO_133 (O_133,N_14844,N_14996);
or UO_134 (O_134,N_14892,N_14961);
and UO_135 (O_135,N_14765,N_14834);
and UO_136 (O_136,N_14842,N_14888);
nand UO_137 (O_137,N_14754,N_14884);
nand UO_138 (O_138,N_14752,N_14914);
or UO_139 (O_139,N_14816,N_14927);
nand UO_140 (O_140,N_14764,N_14915);
or UO_141 (O_141,N_14770,N_14829);
nor UO_142 (O_142,N_14930,N_14801);
nand UO_143 (O_143,N_14909,N_14928);
and UO_144 (O_144,N_14750,N_14875);
or UO_145 (O_145,N_14752,N_14770);
xnor UO_146 (O_146,N_14987,N_14833);
nand UO_147 (O_147,N_14840,N_14846);
nor UO_148 (O_148,N_14841,N_14830);
nor UO_149 (O_149,N_14886,N_14812);
nand UO_150 (O_150,N_14845,N_14954);
nor UO_151 (O_151,N_14996,N_14819);
nand UO_152 (O_152,N_14992,N_14849);
or UO_153 (O_153,N_14989,N_14936);
and UO_154 (O_154,N_14920,N_14816);
xor UO_155 (O_155,N_14776,N_14829);
or UO_156 (O_156,N_14865,N_14857);
and UO_157 (O_157,N_14790,N_14975);
nor UO_158 (O_158,N_14949,N_14755);
nor UO_159 (O_159,N_14999,N_14836);
and UO_160 (O_160,N_14982,N_14970);
or UO_161 (O_161,N_14987,N_14784);
or UO_162 (O_162,N_14918,N_14766);
or UO_163 (O_163,N_14876,N_14962);
and UO_164 (O_164,N_14774,N_14811);
or UO_165 (O_165,N_14867,N_14764);
and UO_166 (O_166,N_14999,N_14879);
nor UO_167 (O_167,N_14803,N_14949);
or UO_168 (O_168,N_14832,N_14756);
or UO_169 (O_169,N_14856,N_14816);
nand UO_170 (O_170,N_14805,N_14887);
and UO_171 (O_171,N_14957,N_14891);
or UO_172 (O_172,N_14966,N_14990);
and UO_173 (O_173,N_14859,N_14796);
and UO_174 (O_174,N_14899,N_14850);
and UO_175 (O_175,N_14865,N_14880);
nand UO_176 (O_176,N_14847,N_14941);
nor UO_177 (O_177,N_14987,N_14873);
and UO_178 (O_178,N_14812,N_14964);
nor UO_179 (O_179,N_14956,N_14757);
and UO_180 (O_180,N_14851,N_14904);
nand UO_181 (O_181,N_14907,N_14811);
nand UO_182 (O_182,N_14992,N_14886);
nor UO_183 (O_183,N_14767,N_14795);
or UO_184 (O_184,N_14791,N_14929);
nand UO_185 (O_185,N_14897,N_14893);
nand UO_186 (O_186,N_14889,N_14989);
xnor UO_187 (O_187,N_14925,N_14754);
and UO_188 (O_188,N_14972,N_14931);
or UO_189 (O_189,N_14833,N_14920);
or UO_190 (O_190,N_14800,N_14787);
nand UO_191 (O_191,N_14770,N_14873);
nor UO_192 (O_192,N_14772,N_14788);
and UO_193 (O_193,N_14935,N_14920);
nor UO_194 (O_194,N_14912,N_14770);
nand UO_195 (O_195,N_14796,N_14760);
and UO_196 (O_196,N_14950,N_14903);
and UO_197 (O_197,N_14895,N_14961);
nor UO_198 (O_198,N_14951,N_14786);
and UO_199 (O_199,N_14859,N_14956);
and UO_200 (O_200,N_14971,N_14990);
and UO_201 (O_201,N_14968,N_14815);
and UO_202 (O_202,N_14952,N_14941);
and UO_203 (O_203,N_14910,N_14812);
xnor UO_204 (O_204,N_14871,N_14854);
xor UO_205 (O_205,N_14802,N_14757);
nand UO_206 (O_206,N_14985,N_14925);
nand UO_207 (O_207,N_14971,N_14927);
nor UO_208 (O_208,N_14994,N_14817);
nand UO_209 (O_209,N_14757,N_14788);
or UO_210 (O_210,N_14848,N_14983);
nor UO_211 (O_211,N_14924,N_14758);
nand UO_212 (O_212,N_14916,N_14910);
nand UO_213 (O_213,N_14960,N_14932);
nand UO_214 (O_214,N_14936,N_14807);
nand UO_215 (O_215,N_14994,N_14962);
nand UO_216 (O_216,N_14792,N_14824);
and UO_217 (O_217,N_14936,N_14767);
nor UO_218 (O_218,N_14789,N_14969);
and UO_219 (O_219,N_14811,N_14752);
nand UO_220 (O_220,N_14939,N_14940);
nand UO_221 (O_221,N_14894,N_14900);
nand UO_222 (O_222,N_14813,N_14801);
nand UO_223 (O_223,N_14871,N_14863);
nand UO_224 (O_224,N_14804,N_14936);
nand UO_225 (O_225,N_14897,N_14936);
xor UO_226 (O_226,N_14789,N_14775);
nor UO_227 (O_227,N_14953,N_14752);
and UO_228 (O_228,N_14814,N_14972);
xor UO_229 (O_229,N_14847,N_14815);
nand UO_230 (O_230,N_14781,N_14831);
or UO_231 (O_231,N_14871,N_14813);
and UO_232 (O_232,N_14837,N_14928);
nand UO_233 (O_233,N_14973,N_14818);
nor UO_234 (O_234,N_14950,N_14879);
and UO_235 (O_235,N_14952,N_14883);
nand UO_236 (O_236,N_14960,N_14787);
and UO_237 (O_237,N_14902,N_14879);
nor UO_238 (O_238,N_14973,N_14800);
nor UO_239 (O_239,N_14855,N_14848);
nand UO_240 (O_240,N_14815,N_14962);
nand UO_241 (O_241,N_14942,N_14887);
nand UO_242 (O_242,N_14854,N_14968);
and UO_243 (O_243,N_14973,N_14982);
xnor UO_244 (O_244,N_14758,N_14754);
and UO_245 (O_245,N_14993,N_14810);
nor UO_246 (O_246,N_14904,N_14752);
nand UO_247 (O_247,N_14799,N_14993);
and UO_248 (O_248,N_14960,N_14804);
nor UO_249 (O_249,N_14771,N_14760);
xor UO_250 (O_250,N_14955,N_14915);
and UO_251 (O_251,N_14972,N_14971);
nand UO_252 (O_252,N_14900,N_14803);
and UO_253 (O_253,N_14997,N_14810);
xnor UO_254 (O_254,N_14877,N_14890);
xnor UO_255 (O_255,N_14770,N_14816);
xor UO_256 (O_256,N_14949,N_14829);
nand UO_257 (O_257,N_14750,N_14869);
nor UO_258 (O_258,N_14760,N_14810);
nand UO_259 (O_259,N_14927,N_14773);
nor UO_260 (O_260,N_14862,N_14924);
nor UO_261 (O_261,N_14776,N_14823);
nand UO_262 (O_262,N_14985,N_14953);
nor UO_263 (O_263,N_14970,N_14859);
or UO_264 (O_264,N_14877,N_14942);
nor UO_265 (O_265,N_14777,N_14763);
nor UO_266 (O_266,N_14777,N_14750);
nor UO_267 (O_267,N_14922,N_14989);
xor UO_268 (O_268,N_14896,N_14784);
nand UO_269 (O_269,N_14891,N_14754);
nor UO_270 (O_270,N_14930,N_14755);
nand UO_271 (O_271,N_14948,N_14980);
or UO_272 (O_272,N_14883,N_14899);
xnor UO_273 (O_273,N_14840,N_14899);
or UO_274 (O_274,N_14763,N_14762);
nand UO_275 (O_275,N_14853,N_14880);
xnor UO_276 (O_276,N_14881,N_14759);
nor UO_277 (O_277,N_14878,N_14884);
xnor UO_278 (O_278,N_14944,N_14867);
nand UO_279 (O_279,N_14924,N_14969);
or UO_280 (O_280,N_14869,N_14936);
nor UO_281 (O_281,N_14973,N_14900);
nor UO_282 (O_282,N_14905,N_14833);
nand UO_283 (O_283,N_14919,N_14935);
or UO_284 (O_284,N_14887,N_14792);
nor UO_285 (O_285,N_14935,N_14781);
and UO_286 (O_286,N_14943,N_14825);
xnor UO_287 (O_287,N_14941,N_14926);
and UO_288 (O_288,N_14808,N_14898);
and UO_289 (O_289,N_14819,N_14932);
nand UO_290 (O_290,N_14918,N_14961);
xor UO_291 (O_291,N_14786,N_14850);
nor UO_292 (O_292,N_14894,N_14870);
xnor UO_293 (O_293,N_14836,N_14753);
or UO_294 (O_294,N_14981,N_14957);
nand UO_295 (O_295,N_14970,N_14811);
nand UO_296 (O_296,N_14860,N_14945);
or UO_297 (O_297,N_14810,N_14896);
and UO_298 (O_298,N_14778,N_14812);
nor UO_299 (O_299,N_14933,N_14784);
nand UO_300 (O_300,N_14841,N_14904);
nor UO_301 (O_301,N_14951,N_14996);
xnor UO_302 (O_302,N_14792,N_14944);
nor UO_303 (O_303,N_14818,N_14906);
nor UO_304 (O_304,N_14946,N_14958);
and UO_305 (O_305,N_14779,N_14838);
or UO_306 (O_306,N_14928,N_14861);
nor UO_307 (O_307,N_14848,N_14985);
xnor UO_308 (O_308,N_14835,N_14905);
and UO_309 (O_309,N_14822,N_14986);
and UO_310 (O_310,N_14756,N_14823);
nor UO_311 (O_311,N_14771,N_14884);
nand UO_312 (O_312,N_14797,N_14959);
and UO_313 (O_313,N_14794,N_14970);
nand UO_314 (O_314,N_14800,N_14984);
or UO_315 (O_315,N_14914,N_14840);
nand UO_316 (O_316,N_14773,N_14955);
and UO_317 (O_317,N_14874,N_14798);
nand UO_318 (O_318,N_14833,N_14934);
and UO_319 (O_319,N_14885,N_14811);
or UO_320 (O_320,N_14887,N_14873);
xor UO_321 (O_321,N_14804,N_14889);
and UO_322 (O_322,N_14947,N_14763);
xnor UO_323 (O_323,N_14927,N_14907);
nor UO_324 (O_324,N_14753,N_14756);
nand UO_325 (O_325,N_14987,N_14809);
nand UO_326 (O_326,N_14913,N_14809);
nand UO_327 (O_327,N_14820,N_14826);
and UO_328 (O_328,N_14870,N_14895);
and UO_329 (O_329,N_14865,N_14899);
xnor UO_330 (O_330,N_14776,N_14895);
or UO_331 (O_331,N_14928,N_14871);
nand UO_332 (O_332,N_14788,N_14754);
and UO_333 (O_333,N_14997,N_14978);
nor UO_334 (O_334,N_14961,N_14910);
nor UO_335 (O_335,N_14975,N_14923);
xnor UO_336 (O_336,N_14853,N_14968);
or UO_337 (O_337,N_14784,N_14761);
xnor UO_338 (O_338,N_14760,N_14819);
xnor UO_339 (O_339,N_14850,N_14964);
and UO_340 (O_340,N_14750,N_14768);
or UO_341 (O_341,N_14912,N_14963);
xor UO_342 (O_342,N_14911,N_14935);
and UO_343 (O_343,N_14965,N_14843);
xnor UO_344 (O_344,N_14996,N_14892);
or UO_345 (O_345,N_14838,N_14782);
and UO_346 (O_346,N_14913,N_14911);
nand UO_347 (O_347,N_14854,N_14911);
nand UO_348 (O_348,N_14993,N_14928);
xor UO_349 (O_349,N_14818,N_14801);
xnor UO_350 (O_350,N_14950,N_14881);
xnor UO_351 (O_351,N_14767,N_14991);
and UO_352 (O_352,N_14973,N_14862);
and UO_353 (O_353,N_14888,N_14869);
xnor UO_354 (O_354,N_14876,N_14893);
and UO_355 (O_355,N_14776,N_14864);
nand UO_356 (O_356,N_14880,N_14876);
or UO_357 (O_357,N_14933,N_14965);
nor UO_358 (O_358,N_14984,N_14818);
xnor UO_359 (O_359,N_14860,N_14788);
xor UO_360 (O_360,N_14858,N_14766);
and UO_361 (O_361,N_14838,N_14772);
xnor UO_362 (O_362,N_14857,N_14823);
nor UO_363 (O_363,N_14857,N_14810);
or UO_364 (O_364,N_14759,N_14866);
and UO_365 (O_365,N_14943,N_14979);
nand UO_366 (O_366,N_14855,N_14876);
nor UO_367 (O_367,N_14820,N_14809);
and UO_368 (O_368,N_14990,N_14765);
nand UO_369 (O_369,N_14941,N_14823);
nor UO_370 (O_370,N_14770,N_14773);
and UO_371 (O_371,N_14871,N_14891);
or UO_372 (O_372,N_14931,N_14835);
nand UO_373 (O_373,N_14829,N_14999);
nor UO_374 (O_374,N_14823,N_14855);
nand UO_375 (O_375,N_14783,N_14976);
nor UO_376 (O_376,N_14928,N_14898);
or UO_377 (O_377,N_14995,N_14965);
nand UO_378 (O_378,N_14886,N_14784);
and UO_379 (O_379,N_14906,N_14842);
and UO_380 (O_380,N_14883,N_14796);
and UO_381 (O_381,N_14902,N_14773);
nor UO_382 (O_382,N_14832,N_14882);
nand UO_383 (O_383,N_14960,N_14777);
nand UO_384 (O_384,N_14995,N_14960);
and UO_385 (O_385,N_14949,N_14960);
xor UO_386 (O_386,N_14752,N_14799);
nor UO_387 (O_387,N_14972,N_14801);
nand UO_388 (O_388,N_14776,N_14761);
nor UO_389 (O_389,N_14980,N_14767);
nand UO_390 (O_390,N_14927,N_14946);
and UO_391 (O_391,N_14940,N_14790);
or UO_392 (O_392,N_14820,N_14972);
or UO_393 (O_393,N_14942,N_14959);
nor UO_394 (O_394,N_14821,N_14815);
or UO_395 (O_395,N_14780,N_14971);
and UO_396 (O_396,N_14905,N_14817);
or UO_397 (O_397,N_14984,N_14815);
nand UO_398 (O_398,N_14835,N_14951);
nor UO_399 (O_399,N_14804,N_14938);
and UO_400 (O_400,N_14951,N_14762);
or UO_401 (O_401,N_14930,N_14779);
nand UO_402 (O_402,N_14983,N_14763);
or UO_403 (O_403,N_14952,N_14861);
or UO_404 (O_404,N_14768,N_14973);
nand UO_405 (O_405,N_14945,N_14790);
xnor UO_406 (O_406,N_14969,N_14828);
nor UO_407 (O_407,N_14895,N_14753);
and UO_408 (O_408,N_14966,N_14961);
nor UO_409 (O_409,N_14753,N_14911);
or UO_410 (O_410,N_14933,N_14794);
nor UO_411 (O_411,N_14956,N_14881);
nand UO_412 (O_412,N_14785,N_14833);
and UO_413 (O_413,N_14853,N_14927);
nor UO_414 (O_414,N_14787,N_14754);
xnor UO_415 (O_415,N_14781,N_14969);
nand UO_416 (O_416,N_14786,N_14931);
or UO_417 (O_417,N_14818,N_14798);
or UO_418 (O_418,N_14959,N_14967);
nand UO_419 (O_419,N_14751,N_14818);
nor UO_420 (O_420,N_14844,N_14940);
or UO_421 (O_421,N_14946,N_14900);
or UO_422 (O_422,N_14927,N_14910);
nor UO_423 (O_423,N_14925,N_14966);
nand UO_424 (O_424,N_14787,N_14755);
and UO_425 (O_425,N_14929,N_14981);
nor UO_426 (O_426,N_14971,N_14881);
or UO_427 (O_427,N_14984,N_14759);
nand UO_428 (O_428,N_14919,N_14754);
nor UO_429 (O_429,N_14762,N_14761);
and UO_430 (O_430,N_14918,N_14750);
nand UO_431 (O_431,N_14950,N_14947);
or UO_432 (O_432,N_14831,N_14867);
or UO_433 (O_433,N_14812,N_14897);
and UO_434 (O_434,N_14893,N_14997);
xnor UO_435 (O_435,N_14843,N_14995);
or UO_436 (O_436,N_14952,N_14895);
xor UO_437 (O_437,N_14961,N_14888);
or UO_438 (O_438,N_14928,N_14792);
nand UO_439 (O_439,N_14864,N_14829);
and UO_440 (O_440,N_14927,N_14967);
nand UO_441 (O_441,N_14750,N_14802);
and UO_442 (O_442,N_14973,N_14784);
nand UO_443 (O_443,N_14754,N_14971);
xnor UO_444 (O_444,N_14852,N_14752);
and UO_445 (O_445,N_14918,N_14837);
or UO_446 (O_446,N_14974,N_14836);
nand UO_447 (O_447,N_14862,N_14833);
xor UO_448 (O_448,N_14836,N_14907);
nor UO_449 (O_449,N_14836,N_14968);
and UO_450 (O_450,N_14932,N_14933);
nor UO_451 (O_451,N_14995,N_14952);
or UO_452 (O_452,N_14895,N_14896);
nor UO_453 (O_453,N_14754,N_14857);
xor UO_454 (O_454,N_14954,N_14966);
or UO_455 (O_455,N_14975,N_14958);
xnor UO_456 (O_456,N_14858,N_14876);
and UO_457 (O_457,N_14793,N_14834);
nor UO_458 (O_458,N_14770,N_14967);
or UO_459 (O_459,N_14874,N_14904);
nand UO_460 (O_460,N_14831,N_14886);
or UO_461 (O_461,N_14986,N_14785);
xor UO_462 (O_462,N_14987,N_14856);
or UO_463 (O_463,N_14862,N_14751);
or UO_464 (O_464,N_14851,N_14808);
or UO_465 (O_465,N_14862,N_14759);
and UO_466 (O_466,N_14779,N_14771);
nand UO_467 (O_467,N_14785,N_14834);
and UO_468 (O_468,N_14906,N_14761);
or UO_469 (O_469,N_14775,N_14780);
nand UO_470 (O_470,N_14780,N_14948);
and UO_471 (O_471,N_14961,N_14759);
or UO_472 (O_472,N_14851,N_14906);
nor UO_473 (O_473,N_14957,N_14822);
or UO_474 (O_474,N_14828,N_14852);
nand UO_475 (O_475,N_14996,N_14808);
xnor UO_476 (O_476,N_14825,N_14995);
and UO_477 (O_477,N_14843,N_14775);
xnor UO_478 (O_478,N_14902,N_14778);
xnor UO_479 (O_479,N_14899,N_14763);
nand UO_480 (O_480,N_14921,N_14847);
nand UO_481 (O_481,N_14983,N_14931);
and UO_482 (O_482,N_14816,N_14921);
and UO_483 (O_483,N_14984,N_14825);
or UO_484 (O_484,N_14920,N_14763);
and UO_485 (O_485,N_14992,N_14889);
nand UO_486 (O_486,N_14880,N_14780);
xor UO_487 (O_487,N_14927,N_14824);
and UO_488 (O_488,N_14782,N_14789);
xnor UO_489 (O_489,N_14976,N_14998);
xnor UO_490 (O_490,N_14802,N_14952);
nor UO_491 (O_491,N_14990,N_14924);
or UO_492 (O_492,N_14831,N_14929);
xor UO_493 (O_493,N_14933,N_14895);
nor UO_494 (O_494,N_14815,N_14944);
xnor UO_495 (O_495,N_14771,N_14941);
xor UO_496 (O_496,N_14758,N_14888);
nand UO_497 (O_497,N_14958,N_14991);
and UO_498 (O_498,N_14875,N_14844);
nand UO_499 (O_499,N_14892,N_14882);
or UO_500 (O_500,N_14935,N_14766);
or UO_501 (O_501,N_14936,N_14764);
or UO_502 (O_502,N_14953,N_14940);
nor UO_503 (O_503,N_14990,N_14842);
nor UO_504 (O_504,N_14813,N_14928);
xnor UO_505 (O_505,N_14938,N_14768);
nor UO_506 (O_506,N_14797,N_14897);
xnor UO_507 (O_507,N_14880,N_14784);
nor UO_508 (O_508,N_14750,N_14778);
nand UO_509 (O_509,N_14794,N_14805);
and UO_510 (O_510,N_14984,N_14862);
and UO_511 (O_511,N_14758,N_14809);
nand UO_512 (O_512,N_14905,N_14851);
or UO_513 (O_513,N_14773,N_14972);
nand UO_514 (O_514,N_14938,N_14977);
nand UO_515 (O_515,N_14938,N_14834);
and UO_516 (O_516,N_14761,N_14785);
nor UO_517 (O_517,N_14758,N_14911);
nand UO_518 (O_518,N_14784,N_14751);
nand UO_519 (O_519,N_14952,N_14750);
and UO_520 (O_520,N_14769,N_14803);
nand UO_521 (O_521,N_14791,N_14964);
and UO_522 (O_522,N_14840,N_14908);
and UO_523 (O_523,N_14826,N_14763);
nand UO_524 (O_524,N_14823,N_14950);
and UO_525 (O_525,N_14930,N_14964);
nand UO_526 (O_526,N_14752,N_14935);
and UO_527 (O_527,N_14813,N_14893);
nor UO_528 (O_528,N_14964,N_14974);
and UO_529 (O_529,N_14952,N_14991);
and UO_530 (O_530,N_14944,N_14992);
nand UO_531 (O_531,N_14897,N_14844);
and UO_532 (O_532,N_14844,N_14922);
nor UO_533 (O_533,N_14787,N_14788);
and UO_534 (O_534,N_14818,N_14803);
nand UO_535 (O_535,N_14893,N_14977);
and UO_536 (O_536,N_14900,N_14819);
xnor UO_537 (O_537,N_14771,N_14942);
xnor UO_538 (O_538,N_14860,N_14965);
and UO_539 (O_539,N_14945,N_14952);
xor UO_540 (O_540,N_14933,N_14856);
nor UO_541 (O_541,N_14927,N_14991);
and UO_542 (O_542,N_14916,N_14848);
or UO_543 (O_543,N_14953,N_14918);
and UO_544 (O_544,N_14926,N_14753);
xnor UO_545 (O_545,N_14870,N_14877);
or UO_546 (O_546,N_14906,N_14950);
nor UO_547 (O_547,N_14910,N_14751);
nand UO_548 (O_548,N_14874,N_14855);
nor UO_549 (O_549,N_14919,N_14768);
xor UO_550 (O_550,N_14885,N_14992);
xor UO_551 (O_551,N_14849,N_14755);
xnor UO_552 (O_552,N_14825,N_14961);
or UO_553 (O_553,N_14751,N_14838);
nor UO_554 (O_554,N_14842,N_14898);
nand UO_555 (O_555,N_14903,N_14978);
and UO_556 (O_556,N_14943,N_14861);
xnor UO_557 (O_557,N_14817,N_14920);
nand UO_558 (O_558,N_14812,N_14832);
nand UO_559 (O_559,N_14903,N_14957);
xor UO_560 (O_560,N_14863,N_14872);
xor UO_561 (O_561,N_14758,N_14970);
nor UO_562 (O_562,N_14900,N_14753);
and UO_563 (O_563,N_14948,N_14947);
and UO_564 (O_564,N_14919,N_14810);
nand UO_565 (O_565,N_14877,N_14908);
xnor UO_566 (O_566,N_14945,N_14997);
xor UO_567 (O_567,N_14884,N_14938);
xnor UO_568 (O_568,N_14839,N_14800);
or UO_569 (O_569,N_14944,N_14859);
nand UO_570 (O_570,N_14790,N_14850);
nor UO_571 (O_571,N_14924,N_14857);
xnor UO_572 (O_572,N_14771,N_14765);
xor UO_573 (O_573,N_14895,N_14866);
nor UO_574 (O_574,N_14875,N_14958);
xnor UO_575 (O_575,N_14797,N_14946);
nor UO_576 (O_576,N_14788,N_14881);
or UO_577 (O_577,N_14896,N_14797);
nor UO_578 (O_578,N_14855,N_14968);
nand UO_579 (O_579,N_14979,N_14822);
xor UO_580 (O_580,N_14753,N_14954);
nor UO_581 (O_581,N_14973,N_14972);
and UO_582 (O_582,N_14865,N_14820);
and UO_583 (O_583,N_14856,N_14772);
and UO_584 (O_584,N_14958,N_14813);
and UO_585 (O_585,N_14948,N_14841);
or UO_586 (O_586,N_14839,N_14767);
nor UO_587 (O_587,N_14948,N_14759);
or UO_588 (O_588,N_14806,N_14892);
or UO_589 (O_589,N_14870,N_14991);
and UO_590 (O_590,N_14752,N_14901);
and UO_591 (O_591,N_14885,N_14892);
nand UO_592 (O_592,N_14845,N_14931);
nand UO_593 (O_593,N_14852,N_14994);
and UO_594 (O_594,N_14868,N_14805);
and UO_595 (O_595,N_14996,N_14983);
xor UO_596 (O_596,N_14906,N_14927);
or UO_597 (O_597,N_14878,N_14831);
nor UO_598 (O_598,N_14973,N_14871);
nand UO_599 (O_599,N_14781,N_14965);
xnor UO_600 (O_600,N_14884,N_14974);
xor UO_601 (O_601,N_14819,N_14952);
nor UO_602 (O_602,N_14989,N_14787);
nand UO_603 (O_603,N_14883,N_14938);
and UO_604 (O_604,N_14849,N_14766);
nand UO_605 (O_605,N_14849,N_14986);
or UO_606 (O_606,N_14993,N_14955);
nand UO_607 (O_607,N_14851,N_14817);
or UO_608 (O_608,N_14890,N_14977);
xor UO_609 (O_609,N_14981,N_14918);
xor UO_610 (O_610,N_14992,N_14896);
and UO_611 (O_611,N_14909,N_14837);
xor UO_612 (O_612,N_14904,N_14790);
nor UO_613 (O_613,N_14941,N_14912);
nor UO_614 (O_614,N_14760,N_14754);
and UO_615 (O_615,N_14767,N_14785);
nor UO_616 (O_616,N_14984,N_14983);
xor UO_617 (O_617,N_14753,N_14779);
xor UO_618 (O_618,N_14977,N_14776);
nand UO_619 (O_619,N_14794,N_14965);
nor UO_620 (O_620,N_14960,N_14892);
xnor UO_621 (O_621,N_14837,N_14874);
and UO_622 (O_622,N_14763,N_14931);
nor UO_623 (O_623,N_14806,N_14896);
nand UO_624 (O_624,N_14970,N_14802);
nand UO_625 (O_625,N_14916,N_14803);
nor UO_626 (O_626,N_14993,N_14969);
xor UO_627 (O_627,N_14934,N_14762);
nand UO_628 (O_628,N_14795,N_14940);
xor UO_629 (O_629,N_14967,N_14940);
and UO_630 (O_630,N_14882,N_14891);
xor UO_631 (O_631,N_14838,N_14816);
nor UO_632 (O_632,N_14805,N_14756);
and UO_633 (O_633,N_14987,N_14751);
and UO_634 (O_634,N_14896,N_14917);
and UO_635 (O_635,N_14953,N_14995);
nand UO_636 (O_636,N_14924,N_14935);
and UO_637 (O_637,N_14966,N_14758);
nor UO_638 (O_638,N_14780,N_14917);
nand UO_639 (O_639,N_14978,N_14831);
and UO_640 (O_640,N_14937,N_14899);
nand UO_641 (O_641,N_14848,N_14763);
nand UO_642 (O_642,N_14934,N_14817);
nand UO_643 (O_643,N_14778,N_14864);
nand UO_644 (O_644,N_14790,N_14823);
nor UO_645 (O_645,N_14885,N_14875);
nand UO_646 (O_646,N_14978,N_14982);
xor UO_647 (O_647,N_14956,N_14765);
and UO_648 (O_648,N_14931,N_14963);
nor UO_649 (O_649,N_14850,N_14986);
xor UO_650 (O_650,N_14981,N_14832);
and UO_651 (O_651,N_14882,N_14896);
and UO_652 (O_652,N_14986,N_14791);
nand UO_653 (O_653,N_14891,N_14758);
or UO_654 (O_654,N_14899,N_14910);
and UO_655 (O_655,N_14959,N_14934);
nand UO_656 (O_656,N_14934,N_14819);
or UO_657 (O_657,N_14928,N_14949);
or UO_658 (O_658,N_14815,N_14826);
nor UO_659 (O_659,N_14941,N_14868);
xor UO_660 (O_660,N_14868,N_14983);
xnor UO_661 (O_661,N_14927,N_14911);
and UO_662 (O_662,N_14881,N_14910);
and UO_663 (O_663,N_14890,N_14930);
xor UO_664 (O_664,N_14953,N_14966);
xor UO_665 (O_665,N_14804,N_14753);
xnor UO_666 (O_666,N_14953,N_14860);
nor UO_667 (O_667,N_14904,N_14845);
xor UO_668 (O_668,N_14823,N_14843);
and UO_669 (O_669,N_14848,N_14760);
and UO_670 (O_670,N_14963,N_14773);
nor UO_671 (O_671,N_14921,N_14881);
xnor UO_672 (O_672,N_14965,N_14765);
or UO_673 (O_673,N_14929,N_14787);
or UO_674 (O_674,N_14798,N_14757);
or UO_675 (O_675,N_14760,N_14949);
xor UO_676 (O_676,N_14804,N_14867);
or UO_677 (O_677,N_14782,N_14927);
or UO_678 (O_678,N_14977,N_14814);
or UO_679 (O_679,N_14962,N_14884);
nor UO_680 (O_680,N_14878,N_14791);
nand UO_681 (O_681,N_14821,N_14893);
nor UO_682 (O_682,N_14937,N_14795);
and UO_683 (O_683,N_14971,N_14892);
and UO_684 (O_684,N_14901,N_14809);
nor UO_685 (O_685,N_14856,N_14759);
or UO_686 (O_686,N_14788,N_14832);
xnor UO_687 (O_687,N_14962,N_14761);
nor UO_688 (O_688,N_14957,N_14857);
nand UO_689 (O_689,N_14780,N_14929);
and UO_690 (O_690,N_14904,N_14827);
or UO_691 (O_691,N_14821,N_14885);
or UO_692 (O_692,N_14902,N_14981);
and UO_693 (O_693,N_14901,N_14767);
or UO_694 (O_694,N_14872,N_14934);
or UO_695 (O_695,N_14859,N_14760);
nand UO_696 (O_696,N_14956,N_14930);
nor UO_697 (O_697,N_14978,N_14843);
and UO_698 (O_698,N_14777,N_14783);
nor UO_699 (O_699,N_14769,N_14960);
nor UO_700 (O_700,N_14764,N_14804);
nand UO_701 (O_701,N_14789,N_14760);
nand UO_702 (O_702,N_14942,N_14878);
and UO_703 (O_703,N_14807,N_14989);
and UO_704 (O_704,N_14905,N_14902);
nor UO_705 (O_705,N_14937,N_14909);
and UO_706 (O_706,N_14797,N_14915);
and UO_707 (O_707,N_14888,N_14755);
or UO_708 (O_708,N_14947,N_14819);
nand UO_709 (O_709,N_14893,N_14827);
or UO_710 (O_710,N_14974,N_14976);
and UO_711 (O_711,N_14891,N_14975);
and UO_712 (O_712,N_14993,N_14932);
and UO_713 (O_713,N_14795,N_14902);
or UO_714 (O_714,N_14979,N_14800);
or UO_715 (O_715,N_14828,N_14754);
xor UO_716 (O_716,N_14936,N_14795);
nand UO_717 (O_717,N_14845,N_14889);
and UO_718 (O_718,N_14811,N_14902);
xor UO_719 (O_719,N_14763,N_14757);
and UO_720 (O_720,N_14986,N_14779);
nand UO_721 (O_721,N_14958,N_14793);
xor UO_722 (O_722,N_14806,N_14972);
nor UO_723 (O_723,N_14961,N_14956);
nor UO_724 (O_724,N_14858,N_14867);
and UO_725 (O_725,N_14836,N_14927);
xnor UO_726 (O_726,N_14930,N_14849);
nor UO_727 (O_727,N_14839,N_14821);
nand UO_728 (O_728,N_14798,N_14800);
xnor UO_729 (O_729,N_14967,N_14975);
xor UO_730 (O_730,N_14852,N_14786);
nand UO_731 (O_731,N_14938,N_14826);
xnor UO_732 (O_732,N_14923,N_14897);
or UO_733 (O_733,N_14980,N_14902);
or UO_734 (O_734,N_14868,N_14786);
or UO_735 (O_735,N_14857,N_14981);
nor UO_736 (O_736,N_14980,N_14802);
or UO_737 (O_737,N_14955,N_14928);
xnor UO_738 (O_738,N_14945,N_14821);
and UO_739 (O_739,N_14970,N_14775);
nand UO_740 (O_740,N_14951,N_14858);
nand UO_741 (O_741,N_14889,N_14945);
nor UO_742 (O_742,N_14805,N_14970);
and UO_743 (O_743,N_14982,N_14955);
xnor UO_744 (O_744,N_14882,N_14972);
nor UO_745 (O_745,N_14983,N_14825);
and UO_746 (O_746,N_14793,N_14891);
or UO_747 (O_747,N_14788,N_14837);
xnor UO_748 (O_748,N_14922,N_14893);
nand UO_749 (O_749,N_14888,N_14994);
nand UO_750 (O_750,N_14916,N_14967);
xor UO_751 (O_751,N_14941,N_14826);
xor UO_752 (O_752,N_14930,N_14978);
and UO_753 (O_753,N_14818,N_14846);
xnor UO_754 (O_754,N_14869,N_14973);
xnor UO_755 (O_755,N_14820,N_14903);
nor UO_756 (O_756,N_14907,N_14941);
or UO_757 (O_757,N_14887,N_14948);
and UO_758 (O_758,N_14967,N_14811);
nand UO_759 (O_759,N_14940,N_14932);
nand UO_760 (O_760,N_14799,N_14983);
nand UO_761 (O_761,N_14910,N_14933);
and UO_762 (O_762,N_14929,N_14828);
nor UO_763 (O_763,N_14953,N_14921);
xor UO_764 (O_764,N_14824,N_14903);
and UO_765 (O_765,N_14991,N_14889);
or UO_766 (O_766,N_14986,N_14781);
nand UO_767 (O_767,N_14828,N_14772);
xnor UO_768 (O_768,N_14972,N_14840);
xnor UO_769 (O_769,N_14795,N_14948);
nor UO_770 (O_770,N_14858,N_14977);
xnor UO_771 (O_771,N_14823,N_14871);
xnor UO_772 (O_772,N_14816,N_14951);
and UO_773 (O_773,N_14755,N_14802);
xor UO_774 (O_774,N_14803,N_14890);
and UO_775 (O_775,N_14952,N_14766);
and UO_776 (O_776,N_14764,N_14785);
or UO_777 (O_777,N_14842,N_14772);
nand UO_778 (O_778,N_14825,N_14986);
nand UO_779 (O_779,N_14857,N_14886);
and UO_780 (O_780,N_14771,N_14807);
and UO_781 (O_781,N_14982,N_14831);
and UO_782 (O_782,N_14851,N_14959);
nand UO_783 (O_783,N_14894,N_14912);
or UO_784 (O_784,N_14877,N_14902);
or UO_785 (O_785,N_14783,N_14798);
and UO_786 (O_786,N_14983,N_14935);
xnor UO_787 (O_787,N_14800,N_14983);
nor UO_788 (O_788,N_14898,N_14964);
and UO_789 (O_789,N_14951,N_14852);
and UO_790 (O_790,N_14973,N_14866);
or UO_791 (O_791,N_14857,N_14790);
nor UO_792 (O_792,N_14781,N_14770);
nand UO_793 (O_793,N_14947,N_14987);
xor UO_794 (O_794,N_14858,N_14857);
and UO_795 (O_795,N_14826,N_14993);
and UO_796 (O_796,N_14927,N_14775);
nor UO_797 (O_797,N_14756,N_14924);
xnor UO_798 (O_798,N_14938,N_14828);
or UO_799 (O_799,N_14854,N_14877);
nor UO_800 (O_800,N_14969,N_14757);
nand UO_801 (O_801,N_14853,N_14826);
nand UO_802 (O_802,N_14979,N_14855);
and UO_803 (O_803,N_14828,N_14791);
or UO_804 (O_804,N_14802,N_14851);
nor UO_805 (O_805,N_14875,N_14827);
or UO_806 (O_806,N_14868,N_14965);
nand UO_807 (O_807,N_14906,N_14914);
xor UO_808 (O_808,N_14943,N_14866);
or UO_809 (O_809,N_14757,N_14889);
nand UO_810 (O_810,N_14823,N_14798);
and UO_811 (O_811,N_14869,N_14952);
nand UO_812 (O_812,N_14802,N_14844);
and UO_813 (O_813,N_14768,N_14898);
nor UO_814 (O_814,N_14847,N_14807);
nand UO_815 (O_815,N_14834,N_14866);
nor UO_816 (O_816,N_14820,N_14817);
nor UO_817 (O_817,N_14974,N_14838);
xnor UO_818 (O_818,N_14848,N_14979);
or UO_819 (O_819,N_14983,N_14787);
or UO_820 (O_820,N_14821,N_14966);
or UO_821 (O_821,N_14808,N_14876);
or UO_822 (O_822,N_14766,N_14946);
xor UO_823 (O_823,N_14961,N_14807);
or UO_824 (O_824,N_14928,N_14884);
or UO_825 (O_825,N_14842,N_14902);
xor UO_826 (O_826,N_14819,N_14989);
or UO_827 (O_827,N_14758,N_14822);
nand UO_828 (O_828,N_14755,N_14941);
or UO_829 (O_829,N_14819,N_14817);
xor UO_830 (O_830,N_14816,N_14773);
xor UO_831 (O_831,N_14959,N_14983);
xor UO_832 (O_832,N_14837,N_14763);
and UO_833 (O_833,N_14806,N_14818);
xnor UO_834 (O_834,N_14752,N_14946);
nor UO_835 (O_835,N_14885,N_14778);
nand UO_836 (O_836,N_14821,N_14961);
nor UO_837 (O_837,N_14751,N_14868);
and UO_838 (O_838,N_14996,N_14924);
xnor UO_839 (O_839,N_14916,N_14759);
nand UO_840 (O_840,N_14924,N_14793);
and UO_841 (O_841,N_14888,N_14760);
or UO_842 (O_842,N_14962,N_14783);
or UO_843 (O_843,N_14866,N_14930);
or UO_844 (O_844,N_14966,N_14918);
or UO_845 (O_845,N_14884,N_14933);
nand UO_846 (O_846,N_14998,N_14821);
nor UO_847 (O_847,N_14801,N_14840);
nand UO_848 (O_848,N_14776,N_14909);
nor UO_849 (O_849,N_14942,N_14872);
xor UO_850 (O_850,N_14833,N_14867);
or UO_851 (O_851,N_14862,N_14951);
nor UO_852 (O_852,N_14975,N_14968);
nand UO_853 (O_853,N_14813,N_14984);
nor UO_854 (O_854,N_14763,N_14924);
nand UO_855 (O_855,N_14974,N_14897);
nand UO_856 (O_856,N_14925,N_14763);
or UO_857 (O_857,N_14899,N_14833);
nand UO_858 (O_858,N_14963,N_14755);
or UO_859 (O_859,N_14921,N_14750);
nand UO_860 (O_860,N_14948,N_14825);
or UO_861 (O_861,N_14953,N_14757);
xnor UO_862 (O_862,N_14907,N_14827);
or UO_863 (O_863,N_14824,N_14996);
or UO_864 (O_864,N_14781,N_14862);
nand UO_865 (O_865,N_14848,N_14935);
xor UO_866 (O_866,N_14917,N_14860);
nor UO_867 (O_867,N_14818,N_14951);
xor UO_868 (O_868,N_14871,N_14829);
or UO_869 (O_869,N_14923,N_14796);
or UO_870 (O_870,N_14907,N_14964);
xnor UO_871 (O_871,N_14782,N_14802);
and UO_872 (O_872,N_14994,N_14823);
or UO_873 (O_873,N_14785,N_14952);
or UO_874 (O_874,N_14996,N_14849);
xnor UO_875 (O_875,N_14929,N_14964);
xnor UO_876 (O_876,N_14751,N_14992);
and UO_877 (O_877,N_14782,N_14823);
nand UO_878 (O_878,N_14842,N_14961);
nand UO_879 (O_879,N_14788,N_14978);
nor UO_880 (O_880,N_14835,N_14935);
nand UO_881 (O_881,N_14982,N_14757);
and UO_882 (O_882,N_14867,N_14902);
xor UO_883 (O_883,N_14834,N_14964);
or UO_884 (O_884,N_14984,N_14793);
nor UO_885 (O_885,N_14834,N_14916);
or UO_886 (O_886,N_14765,N_14892);
xor UO_887 (O_887,N_14782,N_14948);
or UO_888 (O_888,N_14928,N_14895);
xor UO_889 (O_889,N_14894,N_14881);
nor UO_890 (O_890,N_14908,N_14927);
nor UO_891 (O_891,N_14911,N_14794);
nor UO_892 (O_892,N_14855,N_14785);
or UO_893 (O_893,N_14891,N_14844);
nand UO_894 (O_894,N_14845,N_14798);
xor UO_895 (O_895,N_14996,N_14757);
xnor UO_896 (O_896,N_14973,N_14849);
or UO_897 (O_897,N_14966,N_14834);
xnor UO_898 (O_898,N_14904,N_14899);
xnor UO_899 (O_899,N_14791,N_14770);
nand UO_900 (O_900,N_14854,N_14789);
or UO_901 (O_901,N_14958,N_14786);
and UO_902 (O_902,N_14968,N_14755);
xor UO_903 (O_903,N_14774,N_14759);
and UO_904 (O_904,N_14876,N_14833);
nor UO_905 (O_905,N_14836,N_14795);
nand UO_906 (O_906,N_14847,N_14899);
nand UO_907 (O_907,N_14895,N_14754);
nor UO_908 (O_908,N_14780,N_14878);
or UO_909 (O_909,N_14915,N_14807);
nor UO_910 (O_910,N_14945,N_14895);
or UO_911 (O_911,N_14806,N_14979);
nand UO_912 (O_912,N_14783,N_14788);
xnor UO_913 (O_913,N_14867,N_14954);
or UO_914 (O_914,N_14780,N_14885);
nor UO_915 (O_915,N_14783,N_14769);
xnor UO_916 (O_916,N_14869,N_14759);
and UO_917 (O_917,N_14924,N_14824);
and UO_918 (O_918,N_14955,N_14945);
and UO_919 (O_919,N_14891,N_14925);
xnor UO_920 (O_920,N_14874,N_14990);
xnor UO_921 (O_921,N_14882,N_14842);
or UO_922 (O_922,N_14922,N_14803);
and UO_923 (O_923,N_14779,N_14754);
nor UO_924 (O_924,N_14940,N_14878);
and UO_925 (O_925,N_14993,N_14816);
xnor UO_926 (O_926,N_14828,N_14796);
xnor UO_927 (O_927,N_14835,N_14893);
xor UO_928 (O_928,N_14911,N_14890);
xor UO_929 (O_929,N_14905,N_14842);
nor UO_930 (O_930,N_14952,N_14924);
xnor UO_931 (O_931,N_14955,N_14879);
and UO_932 (O_932,N_14814,N_14905);
or UO_933 (O_933,N_14820,N_14992);
nand UO_934 (O_934,N_14832,N_14796);
nor UO_935 (O_935,N_14867,N_14960);
and UO_936 (O_936,N_14800,N_14986);
xnor UO_937 (O_937,N_14910,N_14771);
or UO_938 (O_938,N_14822,N_14820);
nor UO_939 (O_939,N_14906,N_14948);
or UO_940 (O_940,N_14834,N_14831);
xor UO_941 (O_941,N_14798,N_14801);
or UO_942 (O_942,N_14822,N_14985);
or UO_943 (O_943,N_14919,N_14761);
or UO_944 (O_944,N_14852,N_14812);
nand UO_945 (O_945,N_14942,N_14810);
or UO_946 (O_946,N_14903,N_14860);
nand UO_947 (O_947,N_14793,N_14941);
and UO_948 (O_948,N_14991,N_14765);
or UO_949 (O_949,N_14975,N_14877);
nor UO_950 (O_950,N_14803,N_14970);
nand UO_951 (O_951,N_14990,N_14802);
nor UO_952 (O_952,N_14993,N_14830);
and UO_953 (O_953,N_14997,N_14856);
xor UO_954 (O_954,N_14858,N_14750);
or UO_955 (O_955,N_14981,N_14970);
nor UO_956 (O_956,N_14923,N_14971);
nor UO_957 (O_957,N_14785,N_14987);
xnor UO_958 (O_958,N_14771,N_14867);
nor UO_959 (O_959,N_14874,N_14846);
nand UO_960 (O_960,N_14899,N_14874);
nand UO_961 (O_961,N_14840,N_14950);
nor UO_962 (O_962,N_14915,N_14953);
or UO_963 (O_963,N_14882,N_14885);
and UO_964 (O_964,N_14804,N_14823);
or UO_965 (O_965,N_14853,N_14936);
or UO_966 (O_966,N_14971,N_14858);
or UO_967 (O_967,N_14893,N_14767);
xor UO_968 (O_968,N_14970,N_14875);
and UO_969 (O_969,N_14952,N_14797);
nand UO_970 (O_970,N_14926,N_14904);
and UO_971 (O_971,N_14952,N_14888);
and UO_972 (O_972,N_14969,N_14989);
xnor UO_973 (O_973,N_14913,N_14839);
or UO_974 (O_974,N_14935,N_14840);
and UO_975 (O_975,N_14752,N_14961);
and UO_976 (O_976,N_14782,N_14855);
and UO_977 (O_977,N_14860,N_14818);
or UO_978 (O_978,N_14788,N_14967);
or UO_979 (O_979,N_14887,N_14901);
nor UO_980 (O_980,N_14851,N_14892);
and UO_981 (O_981,N_14822,N_14834);
or UO_982 (O_982,N_14876,N_14859);
and UO_983 (O_983,N_14827,N_14863);
nand UO_984 (O_984,N_14984,N_14994);
nor UO_985 (O_985,N_14928,N_14938);
and UO_986 (O_986,N_14980,N_14800);
and UO_987 (O_987,N_14981,N_14824);
or UO_988 (O_988,N_14751,N_14926);
xnor UO_989 (O_989,N_14808,N_14895);
nor UO_990 (O_990,N_14825,N_14952);
xor UO_991 (O_991,N_14851,N_14821);
or UO_992 (O_992,N_14947,N_14998);
nor UO_993 (O_993,N_14777,N_14911);
xor UO_994 (O_994,N_14780,N_14857);
xnor UO_995 (O_995,N_14897,N_14996);
or UO_996 (O_996,N_14962,N_14971);
and UO_997 (O_997,N_14771,N_14804);
and UO_998 (O_998,N_14783,N_14916);
nand UO_999 (O_999,N_14988,N_14839);
and UO_1000 (O_1000,N_14756,N_14964);
nor UO_1001 (O_1001,N_14857,N_14866);
xor UO_1002 (O_1002,N_14920,N_14848);
and UO_1003 (O_1003,N_14792,N_14857);
nand UO_1004 (O_1004,N_14754,N_14825);
or UO_1005 (O_1005,N_14751,N_14957);
xnor UO_1006 (O_1006,N_14966,N_14885);
and UO_1007 (O_1007,N_14799,N_14775);
or UO_1008 (O_1008,N_14893,N_14950);
and UO_1009 (O_1009,N_14947,N_14934);
and UO_1010 (O_1010,N_14925,N_14960);
xnor UO_1011 (O_1011,N_14898,N_14904);
and UO_1012 (O_1012,N_14771,N_14846);
nand UO_1013 (O_1013,N_14775,N_14955);
nand UO_1014 (O_1014,N_14965,N_14810);
and UO_1015 (O_1015,N_14820,N_14754);
and UO_1016 (O_1016,N_14908,N_14827);
or UO_1017 (O_1017,N_14864,N_14773);
nor UO_1018 (O_1018,N_14754,N_14985);
or UO_1019 (O_1019,N_14880,N_14890);
or UO_1020 (O_1020,N_14899,N_14757);
or UO_1021 (O_1021,N_14848,N_14955);
xnor UO_1022 (O_1022,N_14937,N_14764);
xnor UO_1023 (O_1023,N_14835,N_14956);
and UO_1024 (O_1024,N_14985,N_14910);
nand UO_1025 (O_1025,N_14841,N_14844);
nor UO_1026 (O_1026,N_14768,N_14979);
xnor UO_1027 (O_1027,N_14872,N_14973);
xnor UO_1028 (O_1028,N_14920,N_14975);
or UO_1029 (O_1029,N_14832,N_14935);
or UO_1030 (O_1030,N_14914,N_14922);
nand UO_1031 (O_1031,N_14811,N_14986);
and UO_1032 (O_1032,N_14999,N_14872);
nand UO_1033 (O_1033,N_14864,N_14862);
nand UO_1034 (O_1034,N_14830,N_14909);
or UO_1035 (O_1035,N_14805,N_14783);
nand UO_1036 (O_1036,N_14827,N_14993);
or UO_1037 (O_1037,N_14802,N_14923);
and UO_1038 (O_1038,N_14837,N_14941);
nor UO_1039 (O_1039,N_14985,N_14758);
nor UO_1040 (O_1040,N_14842,N_14812);
or UO_1041 (O_1041,N_14846,N_14790);
nor UO_1042 (O_1042,N_14751,N_14831);
or UO_1043 (O_1043,N_14994,N_14906);
or UO_1044 (O_1044,N_14934,N_14993);
nor UO_1045 (O_1045,N_14969,N_14877);
nand UO_1046 (O_1046,N_14825,N_14766);
nand UO_1047 (O_1047,N_14964,N_14894);
nor UO_1048 (O_1048,N_14796,N_14825);
nand UO_1049 (O_1049,N_14977,N_14847);
xor UO_1050 (O_1050,N_14957,N_14837);
nand UO_1051 (O_1051,N_14967,N_14895);
nor UO_1052 (O_1052,N_14817,N_14977);
or UO_1053 (O_1053,N_14843,N_14922);
and UO_1054 (O_1054,N_14857,N_14793);
nor UO_1055 (O_1055,N_14865,N_14908);
xor UO_1056 (O_1056,N_14859,N_14846);
nand UO_1057 (O_1057,N_14815,N_14849);
xor UO_1058 (O_1058,N_14850,N_14815);
nand UO_1059 (O_1059,N_14773,N_14822);
nand UO_1060 (O_1060,N_14840,N_14767);
nand UO_1061 (O_1061,N_14851,N_14829);
nand UO_1062 (O_1062,N_14865,N_14992);
or UO_1063 (O_1063,N_14802,N_14936);
nor UO_1064 (O_1064,N_14874,N_14845);
nand UO_1065 (O_1065,N_14984,N_14975);
nor UO_1066 (O_1066,N_14936,N_14851);
nor UO_1067 (O_1067,N_14988,N_14938);
nor UO_1068 (O_1068,N_14842,N_14976);
and UO_1069 (O_1069,N_14872,N_14966);
xor UO_1070 (O_1070,N_14793,N_14959);
and UO_1071 (O_1071,N_14862,N_14882);
and UO_1072 (O_1072,N_14859,N_14785);
nor UO_1073 (O_1073,N_14808,N_14899);
nor UO_1074 (O_1074,N_14901,N_14894);
or UO_1075 (O_1075,N_14883,N_14997);
nor UO_1076 (O_1076,N_14924,N_14946);
and UO_1077 (O_1077,N_14917,N_14755);
or UO_1078 (O_1078,N_14968,N_14861);
nor UO_1079 (O_1079,N_14902,N_14911);
or UO_1080 (O_1080,N_14766,N_14882);
or UO_1081 (O_1081,N_14932,N_14981);
and UO_1082 (O_1082,N_14990,N_14899);
or UO_1083 (O_1083,N_14920,N_14872);
or UO_1084 (O_1084,N_14950,N_14845);
and UO_1085 (O_1085,N_14897,N_14907);
nor UO_1086 (O_1086,N_14975,N_14856);
and UO_1087 (O_1087,N_14973,N_14782);
or UO_1088 (O_1088,N_14955,N_14756);
and UO_1089 (O_1089,N_14865,N_14821);
xnor UO_1090 (O_1090,N_14959,N_14835);
nor UO_1091 (O_1091,N_14898,N_14913);
nor UO_1092 (O_1092,N_14955,N_14890);
nor UO_1093 (O_1093,N_14948,N_14973);
nor UO_1094 (O_1094,N_14762,N_14961);
nor UO_1095 (O_1095,N_14992,N_14843);
nand UO_1096 (O_1096,N_14955,N_14926);
nor UO_1097 (O_1097,N_14974,N_14951);
and UO_1098 (O_1098,N_14968,N_14969);
nor UO_1099 (O_1099,N_14895,N_14940);
nand UO_1100 (O_1100,N_14937,N_14875);
nand UO_1101 (O_1101,N_14957,N_14856);
nand UO_1102 (O_1102,N_14786,N_14878);
nor UO_1103 (O_1103,N_14927,N_14969);
or UO_1104 (O_1104,N_14759,N_14878);
nand UO_1105 (O_1105,N_14770,N_14890);
and UO_1106 (O_1106,N_14927,N_14897);
and UO_1107 (O_1107,N_14751,N_14882);
xor UO_1108 (O_1108,N_14811,N_14891);
nor UO_1109 (O_1109,N_14910,N_14929);
nor UO_1110 (O_1110,N_14962,N_14813);
xor UO_1111 (O_1111,N_14767,N_14908);
and UO_1112 (O_1112,N_14807,N_14825);
nor UO_1113 (O_1113,N_14827,N_14998);
or UO_1114 (O_1114,N_14876,N_14904);
nor UO_1115 (O_1115,N_14876,N_14789);
and UO_1116 (O_1116,N_14840,N_14820);
or UO_1117 (O_1117,N_14829,N_14913);
nor UO_1118 (O_1118,N_14953,N_14821);
nor UO_1119 (O_1119,N_14884,N_14865);
or UO_1120 (O_1120,N_14916,N_14939);
nand UO_1121 (O_1121,N_14795,N_14990);
xnor UO_1122 (O_1122,N_14898,N_14791);
nand UO_1123 (O_1123,N_14870,N_14836);
nand UO_1124 (O_1124,N_14907,N_14968);
and UO_1125 (O_1125,N_14820,N_14973);
xnor UO_1126 (O_1126,N_14810,N_14861);
nand UO_1127 (O_1127,N_14920,N_14987);
or UO_1128 (O_1128,N_14967,N_14855);
nor UO_1129 (O_1129,N_14821,N_14882);
nand UO_1130 (O_1130,N_14932,N_14873);
nand UO_1131 (O_1131,N_14853,N_14852);
or UO_1132 (O_1132,N_14766,N_14774);
nand UO_1133 (O_1133,N_14822,N_14946);
or UO_1134 (O_1134,N_14798,N_14917);
nand UO_1135 (O_1135,N_14986,N_14778);
nor UO_1136 (O_1136,N_14816,N_14803);
and UO_1137 (O_1137,N_14860,N_14912);
xor UO_1138 (O_1138,N_14924,N_14787);
and UO_1139 (O_1139,N_14808,N_14908);
xnor UO_1140 (O_1140,N_14773,N_14751);
xor UO_1141 (O_1141,N_14846,N_14932);
or UO_1142 (O_1142,N_14903,N_14779);
or UO_1143 (O_1143,N_14764,N_14864);
nand UO_1144 (O_1144,N_14761,N_14940);
xor UO_1145 (O_1145,N_14776,N_14998);
xnor UO_1146 (O_1146,N_14755,N_14751);
xor UO_1147 (O_1147,N_14936,N_14854);
xnor UO_1148 (O_1148,N_14767,N_14862);
nor UO_1149 (O_1149,N_14935,N_14809);
nand UO_1150 (O_1150,N_14856,N_14769);
and UO_1151 (O_1151,N_14810,N_14838);
or UO_1152 (O_1152,N_14907,N_14983);
nand UO_1153 (O_1153,N_14816,N_14843);
nor UO_1154 (O_1154,N_14951,N_14967);
nand UO_1155 (O_1155,N_14879,N_14769);
nor UO_1156 (O_1156,N_14770,N_14978);
xnor UO_1157 (O_1157,N_14866,N_14941);
and UO_1158 (O_1158,N_14877,N_14881);
xnor UO_1159 (O_1159,N_14840,N_14880);
or UO_1160 (O_1160,N_14859,N_14926);
nor UO_1161 (O_1161,N_14882,N_14871);
and UO_1162 (O_1162,N_14963,N_14893);
nand UO_1163 (O_1163,N_14951,N_14955);
xnor UO_1164 (O_1164,N_14763,N_14930);
nor UO_1165 (O_1165,N_14967,N_14812);
xnor UO_1166 (O_1166,N_14851,N_14963);
xor UO_1167 (O_1167,N_14888,N_14886);
and UO_1168 (O_1168,N_14814,N_14891);
nand UO_1169 (O_1169,N_14778,N_14889);
or UO_1170 (O_1170,N_14785,N_14933);
and UO_1171 (O_1171,N_14937,N_14891);
nor UO_1172 (O_1172,N_14755,N_14989);
or UO_1173 (O_1173,N_14950,N_14821);
xor UO_1174 (O_1174,N_14758,N_14781);
nor UO_1175 (O_1175,N_14887,N_14994);
nand UO_1176 (O_1176,N_14911,N_14867);
and UO_1177 (O_1177,N_14797,N_14823);
and UO_1178 (O_1178,N_14940,N_14779);
xnor UO_1179 (O_1179,N_14824,N_14768);
or UO_1180 (O_1180,N_14999,N_14903);
nor UO_1181 (O_1181,N_14909,N_14799);
or UO_1182 (O_1182,N_14875,N_14881);
nand UO_1183 (O_1183,N_14920,N_14883);
xor UO_1184 (O_1184,N_14925,N_14858);
and UO_1185 (O_1185,N_14886,N_14843);
nand UO_1186 (O_1186,N_14792,N_14846);
xor UO_1187 (O_1187,N_14873,N_14822);
nand UO_1188 (O_1188,N_14929,N_14939);
or UO_1189 (O_1189,N_14885,N_14753);
or UO_1190 (O_1190,N_14977,N_14933);
xor UO_1191 (O_1191,N_14825,N_14978);
and UO_1192 (O_1192,N_14969,N_14957);
xnor UO_1193 (O_1193,N_14810,N_14835);
or UO_1194 (O_1194,N_14867,N_14806);
and UO_1195 (O_1195,N_14882,N_14872);
xor UO_1196 (O_1196,N_14765,N_14934);
xnor UO_1197 (O_1197,N_14769,N_14815);
nand UO_1198 (O_1198,N_14838,N_14883);
and UO_1199 (O_1199,N_14822,N_14861);
nor UO_1200 (O_1200,N_14782,N_14757);
xnor UO_1201 (O_1201,N_14849,N_14896);
nor UO_1202 (O_1202,N_14771,N_14816);
nor UO_1203 (O_1203,N_14892,N_14988);
nand UO_1204 (O_1204,N_14823,N_14759);
nand UO_1205 (O_1205,N_14910,N_14825);
or UO_1206 (O_1206,N_14832,N_14775);
and UO_1207 (O_1207,N_14787,N_14820);
or UO_1208 (O_1208,N_14790,N_14772);
and UO_1209 (O_1209,N_14821,N_14928);
nor UO_1210 (O_1210,N_14956,N_14784);
nand UO_1211 (O_1211,N_14892,N_14803);
and UO_1212 (O_1212,N_14868,N_14969);
or UO_1213 (O_1213,N_14774,N_14987);
xor UO_1214 (O_1214,N_14961,N_14972);
or UO_1215 (O_1215,N_14949,N_14980);
xor UO_1216 (O_1216,N_14885,N_14923);
or UO_1217 (O_1217,N_14919,N_14947);
nand UO_1218 (O_1218,N_14923,N_14970);
nand UO_1219 (O_1219,N_14961,N_14954);
or UO_1220 (O_1220,N_14997,N_14940);
and UO_1221 (O_1221,N_14909,N_14826);
or UO_1222 (O_1222,N_14886,N_14927);
or UO_1223 (O_1223,N_14836,N_14800);
or UO_1224 (O_1224,N_14922,N_14846);
and UO_1225 (O_1225,N_14815,N_14889);
nor UO_1226 (O_1226,N_14926,N_14877);
xnor UO_1227 (O_1227,N_14998,N_14930);
and UO_1228 (O_1228,N_14776,N_14916);
nand UO_1229 (O_1229,N_14920,N_14986);
xnor UO_1230 (O_1230,N_14863,N_14858);
nor UO_1231 (O_1231,N_14922,N_14979);
and UO_1232 (O_1232,N_14911,N_14782);
xnor UO_1233 (O_1233,N_14811,N_14917);
or UO_1234 (O_1234,N_14871,N_14909);
or UO_1235 (O_1235,N_14824,N_14918);
and UO_1236 (O_1236,N_14958,N_14802);
nand UO_1237 (O_1237,N_14832,N_14839);
nand UO_1238 (O_1238,N_14765,N_14846);
or UO_1239 (O_1239,N_14772,N_14865);
nor UO_1240 (O_1240,N_14797,N_14888);
and UO_1241 (O_1241,N_14788,N_14920);
xnor UO_1242 (O_1242,N_14942,N_14955);
xor UO_1243 (O_1243,N_14798,N_14899);
or UO_1244 (O_1244,N_14994,N_14812);
and UO_1245 (O_1245,N_14757,N_14959);
or UO_1246 (O_1246,N_14936,N_14914);
and UO_1247 (O_1247,N_14992,N_14910);
nor UO_1248 (O_1248,N_14796,N_14875);
xnor UO_1249 (O_1249,N_14995,N_14771);
and UO_1250 (O_1250,N_14898,N_14918);
nand UO_1251 (O_1251,N_14826,N_14782);
nor UO_1252 (O_1252,N_14868,N_14820);
xor UO_1253 (O_1253,N_14980,N_14926);
or UO_1254 (O_1254,N_14828,N_14755);
nor UO_1255 (O_1255,N_14803,N_14889);
xor UO_1256 (O_1256,N_14804,N_14890);
nor UO_1257 (O_1257,N_14920,N_14891);
xnor UO_1258 (O_1258,N_14818,N_14896);
and UO_1259 (O_1259,N_14762,N_14952);
xor UO_1260 (O_1260,N_14985,N_14849);
and UO_1261 (O_1261,N_14770,N_14883);
and UO_1262 (O_1262,N_14899,N_14830);
and UO_1263 (O_1263,N_14846,N_14866);
nand UO_1264 (O_1264,N_14945,N_14875);
or UO_1265 (O_1265,N_14922,N_14970);
xnor UO_1266 (O_1266,N_14895,N_14761);
nand UO_1267 (O_1267,N_14954,N_14995);
or UO_1268 (O_1268,N_14862,N_14964);
nor UO_1269 (O_1269,N_14772,N_14893);
nand UO_1270 (O_1270,N_14984,N_14767);
and UO_1271 (O_1271,N_14908,N_14805);
and UO_1272 (O_1272,N_14946,N_14826);
nor UO_1273 (O_1273,N_14834,N_14873);
or UO_1274 (O_1274,N_14985,N_14774);
nor UO_1275 (O_1275,N_14939,N_14787);
nand UO_1276 (O_1276,N_14864,N_14980);
xnor UO_1277 (O_1277,N_14996,N_14976);
xor UO_1278 (O_1278,N_14892,N_14751);
nand UO_1279 (O_1279,N_14941,N_14872);
xor UO_1280 (O_1280,N_14922,N_14795);
or UO_1281 (O_1281,N_14937,N_14871);
nor UO_1282 (O_1282,N_14851,N_14880);
or UO_1283 (O_1283,N_14976,N_14926);
nor UO_1284 (O_1284,N_14813,N_14993);
or UO_1285 (O_1285,N_14756,N_14906);
nor UO_1286 (O_1286,N_14755,N_14843);
and UO_1287 (O_1287,N_14987,N_14768);
nand UO_1288 (O_1288,N_14818,N_14808);
nor UO_1289 (O_1289,N_14995,N_14984);
nor UO_1290 (O_1290,N_14752,N_14900);
nor UO_1291 (O_1291,N_14821,N_14868);
and UO_1292 (O_1292,N_14953,N_14837);
xor UO_1293 (O_1293,N_14814,N_14997);
nor UO_1294 (O_1294,N_14813,N_14784);
nor UO_1295 (O_1295,N_14962,N_14952);
nand UO_1296 (O_1296,N_14868,N_14866);
or UO_1297 (O_1297,N_14824,N_14994);
and UO_1298 (O_1298,N_14813,N_14883);
and UO_1299 (O_1299,N_14918,N_14888);
or UO_1300 (O_1300,N_14984,N_14978);
nand UO_1301 (O_1301,N_14805,N_14924);
and UO_1302 (O_1302,N_14872,N_14820);
nor UO_1303 (O_1303,N_14801,N_14757);
or UO_1304 (O_1304,N_14878,N_14781);
nand UO_1305 (O_1305,N_14967,N_14885);
xor UO_1306 (O_1306,N_14773,N_14911);
nand UO_1307 (O_1307,N_14985,N_14770);
and UO_1308 (O_1308,N_14783,N_14995);
or UO_1309 (O_1309,N_14844,N_14990);
nand UO_1310 (O_1310,N_14883,N_14823);
nand UO_1311 (O_1311,N_14884,N_14959);
and UO_1312 (O_1312,N_14841,N_14888);
and UO_1313 (O_1313,N_14995,N_14852);
and UO_1314 (O_1314,N_14811,N_14837);
or UO_1315 (O_1315,N_14850,N_14806);
nor UO_1316 (O_1316,N_14974,N_14803);
nand UO_1317 (O_1317,N_14783,N_14982);
nor UO_1318 (O_1318,N_14891,N_14982);
or UO_1319 (O_1319,N_14914,N_14920);
xnor UO_1320 (O_1320,N_14895,N_14983);
or UO_1321 (O_1321,N_14800,N_14913);
and UO_1322 (O_1322,N_14917,N_14822);
and UO_1323 (O_1323,N_14989,N_14804);
nor UO_1324 (O_1324,N_14763,N_14999);
and UO_1325 (O_1325,N_14800,N_14874);
nand UO_1326 (O_1326,N_14881,N_14966);
nor UO_1327 (O_1327,N_14799,N_14827);
nand UO_1328 (O_1328,N_14953,N_14926);
nor UO_1329 (O_1329,N_14899,N_14988);
and UO_1330 (O_1330,N_14866,N_14905);
xor UO_1331 (O_1331,N_14878,N_14924);
nand UO_1332 (O_1332,N_14906,N_14811);
and UO_1333 (O_1333,N_14813,N_14786);
or UO_1334 (O_1334,N_14899,N_14839);
nor UO_1335 (O_1335,N_14872,N_14996);
nor UO_1336 (O_1336,N_14776,N_14947);
nor UO_1337 (O_1337,N_14951,N_14804);
xor UO_1338 (O_1338,N_14823,N_14878);
or UO_1339 (O_1339,N_14769,N_14810);
nor UO_1340 (O_1340,N_14834,N_14867);
xor UO_1341 (O_1341,N_14923,N_14896);
or UO_1342 (O_1342,N_14851,N_14753);
nor UO_1343 (O_1343,N_14776,N_14870);
or UO_1344 (O_1344,N_14848,N_14896);
xor UO_1345 (O_1345,N_14756,N_14843);
nand UO_1346 (O_1346,N_14779,N_14815);
nand UO_1347 (O_1347,N_14986,N_14936);
or UO_1348 (O_1348,N_14863,N_14949);
xor UO_1349 (O_1349,N_14921,N_14789);
nand UO_1350 (O_1350,N_14930,N_14862);
nand UO_1351 (O_1351,N_14831,N_14980);
xor UO_1352 (O_1352,N_14866,N_14784);
xnor UO_1353 (O_1353,N_14889,N_14819);
xor UO_1354 (O_1354,N_14982,N_14889);
and UO_1355 (O_1355,N_14855,N_14993);
and UO_1356 (O_1356,N_14839,N_14961);
xor UO_1357 (O_1357,N_14772,N_14858);
and UO_1358 (O_1358,N_14802,N_14995);
nand UO_1359 (O_1359,N_14981,N_14921);
and UO_1360 (O_1360,N_14945,N_14879);
nor UO_1361 (O_1361,N_14897,N_14813);
xor UO_1362 (O_1362,N_14985,N_14992);
nand UO_1363 (O_1363,N_14891,N_14859);
nand UO_1364 (O_1364,N_14779,N_14793);
xnor UO_1365 (O_1365,N_14783,N_14786);
nand UO_1366 (O_1366,N_14975,N_14926);
nand UO_1367 (O_1367,N_14782,N_14923);
and UO_1368 (O_1368,N_14856,N_14948);
or UO_1369 (O_1369,N_14899,N_14880);
nand UO_1370 (O_1370,N_14996,N_14914);
nor UO_1371 (O_1371,N_14752,N_14764);
nor UO_1372 (O_1372,N_14849,N_14835);
xnor UO_1373 (O_1373,N_14806,N_14776);
and UO_1374 (O_1374,N_14797,N_14961);
and UO_1375 (O_1375,N_14757,N_14846);
xor UO_1376 (O_1376,N_14827,N_14852);
and UO_1377 (O_1377,N_14798,N_14927);
nand UO_1378 (O_1378,N_14768,N_14999);
nor UO_1379 (O_1379,N_14766,N_14965);
nor UO_1380 (O_1380,N_14960,N_14935);
and UO_1381 (O_1381,N_14755,N_14875);
or UO_1382 (O_1382,N_14987,N_14858);
xnor UO_1383 (O_1383,N_14813,N_14987);
or UO_1384 (O_1384,N_14858,N_14773);
and UO_1385 (O_1385,N_14775,N_14918);
xor UO_1386 (O_1386,N_14819,N_14912);
xnor UO_1387 (O_1387,N_14955,N_14824);
or UO_1388 (O_1388,N_14961,N_14805);
nand UO_1389 (O_1389,N_14854,N_14921);
or UO_1390 (O_1390,N_14848,N_14872);
nand UO_1391 (O_1391,N_14859,N_14875);
nand UO_1392 (O_1392,N_14956,N_14854);
and UO_1393 (O_1393,N_14775,N_14796);
xnor UO_1394 (O_1394,N_14994,N_14954);
nor UO_1395 (O_1395,N_14757,N_14916);
xor UO_1396 (O_1396,N_14943,N_14843);
nor UO_1397 (O_1397,N_14855,N_14808);
nor UO_1398 (O_1398,N_14958,N_14821);
nor UO_1399 (O_1399,N_14804,N_14891);
xnor UO_1400 (O_1400,N_14790,N_14901);
xor UO_1401 (O_1401,N_14771,N_14753);
nor UO_1402 (O_1402,N_14843,N_14926);
nand UO_1403 (O_1403,N_14914,N_14957);
or UO_1404 (O_1404,N_14975,N_14991);
nor UO_1405 (O_1405,N_14769,N_14867);
or UO_1406 (O_1406,N_14775,N_14756);
nand UO_1407 (O_1407,N_14831,N_14923);
xnor UO_1408 (O_1408,N_14942,N_14793);
and UO_1409 (O_1409,N_14770,N_14954);
xor UO_1410 (O_1410,N_14866,N_14854);
xor UO_1411 (O_1411,N_14812,N_14948);
nor UO_1412 (O_1412,N_14751,N_14797);
or UO_1413 (O_1413,N_14761,N_14973);
or UO_1414 (O_1414,N_14897,N_14921);
or UO_1415 (O_1415,N_14838,N_14896);
xor UO_1416 (O_1416,N_14860,N_14856);
and UO_1417 (O_1417,N_14835,N_14950);
and UO_1418 (O_1418,N_14988,N_14838);
nand UO_1419 (O_1419,N_14767,N_14934);
nand UO_1420 (O_1420,N_14820,N_14889);
nand UO_1421 (O_1421,N_14994,N_14865);
nand UO_1422 (O_1422,N_14915,N_14778);
nor UO_1423 (O_1423,N_14778,N_14881);
xnor UO_1424 (O_1424,N_14866,N_14827);
nor UO_1425 (O_1425,N_14842,N_14807);
xnor UO_1426 (O_1426,N_14909,N_14910);
nand UO_1427 (O_1427,N_14927,N_14966);
nor UO_1428 (O_1428,N_14930,N_14963);
or UO_1429 (O_1429,N_14969,N_14881);
and UO_1430 (O_1430,N_14873,N_14890);
nor UO_1431 (O_1431,N_14955,N_14751);
and UO_1432 (O_1432,N_14762,N_14813);
nand UO_1433 (O_1433,N_14873,N_14776);
nand UO_1434 (O_1434,N_14915,N_14972);
and UO_1435 (O_1435,N_14782,N_14868);
nand UO_1436 (O_1436,N_14909,N_14894);
nand UO_1437 (O_1437,N_14915,N_14947);
nor UO_1438 (O_1438,N_14871,N_14830);
or UO_1439 (O_1439,N_14838,N_14758);
xor UO_1440 (O_1440,N_14783,N_14885);
and UO_1441 (O_1441,N_14777,N_14782);
xor UO_1442 (O_1442,N_14895,N_14807);
nand UO_1443 (O_1443,N_14771,N_14755);
xnor UO_1444 (O_1444,N_14805,N_14997);
nor UO_1445 (O_1445,N_14934,N_14834);
nor UO_1446 (O_1446,N_14831,N_14877);
xnor UO_1447 (O_1447,N_14754,N_14811);
nand UO_1448 (O_1448,N_14972,N_14750);
nor UO_1449 (O_1449,N_14884,N_14862);
nand UO_1450 (O_1450,N_14931,N_14829);
xor UO_1451 (O_1451,N_14875,N_14979);
nand UO_1452 (O_1452,N_14958,N_14882);
and UO_1453 (O_1453,N_14895,N_14916);
or UO_1454 (O_1454,N_14917,N_14836);
xor UO_1455 (O_1455,N_14843,N_14944);
xor UO_1456 (O_1456,N_14792,N_14940);
nand UO_1457 (O_1457,N_14825,N_14802);
xor UO_1458 (O_1458,N_14927,N_14928);
nor UO_1459 (O_1459,N_14799,N_14844);
nor UO_1460 (O_1460,N_14946,N_14859);
xnor UO_1461 (O_1461,N_14912,N_14832);
or UO_1462 (O_1462,N_14796,N_14961);
xnor UO_1463 (O_1463,N_14850,N_14760);
or UO_1464 (O_1464,N_14847,N_14869);
or UO_1465 (O_1465,N_14795,N_14919);
xor UO_1466 (O_1466,N_14883,N_14947);
or UO_1467 (O_1467,N_14944,N_14905);
nand UO_1468 (O_1468,N_14932,N_14816);
nand UO_1469 (O_1469,N_14870,N_14810);
xor UO_1470 (O_1470,N_14771,N_14994);
nand UO_1471 (O_1471,N_14764,N_14836);
nand UO_1472 (O_1472,N_14950,N_14901);
nand UO_1473 (O_1473,N_14750,N_14780);
or UO_1474 (O_1474,N_14868,N_14992);
nand UO_1475 (O_1475,N_14795,N_14751);
and UO_1476 (O_1476,N_14833,N_14868);
nor UO_1477 (O_1477,N_14957,N_14917);
nand UO_1478 (O_1478,N_14790,N_14892);
nor UO_1479 (O_1479,N_14789,N_14814);
nand UO_1480 (O_1480,N_14941,N_14910);
nor UO_1481 (O_1481,N_14775,N_14800);
nor UO_1482 (O_1482,N_14758,N_14848);
nand UO_1483 (O_1483,N_14947,N_14841);
nor UO_1484 (O_1484,N_14958,N_14963);
nand UO_1485 (O_1485,N_14957,N_14871);
nor UO_1486 (O_1486,N_14813,N_14981);
xnor UO_1487 (O_1487,N_14759,N_14846);
nand UO_1488 (O_1488,N_14861,N_14991);
nand UO_1489 (O_1489,N_14894,N_14810);
nor UO_1490 (O_1490,N_14986,N_14864);
xnor UO_1491 (O_1491,N_14873,N_14991);
or UO_1492 (O_1492,N_14751,N_14948);
and UO_1493 (O_1493,N_14835,N_14825);
or UO_1494 (O_1494,N_14786,N_14907);
or UO_1495 (O_1495,N_14990,N_14817);
nor UO_1496 (O_1496,N_14811,N_14790);
nor UO_1497 (O_1497,N_14876,N_14857);
nand UO_1498 (O_1498,N_14864,N_14963);
nand UO_1499 (O_1499,N_14774,N_14777);
nand UO_1500 (O_1500,N_14885,N_14775);
or UO_1501 (O_1501,N_14875,N_14964);
nand UO_1502 (O_1502,N_14924,N_14923);
and UO_1503 (O_1503,N_14906,N_14843);
and UO_1504 (O_1504,N_14824,N_14786);
nor UO_1505 (O_1505,N_14760,N_14772);
nand UO_1506 (O_1506,N_14991,N_14950);
xor UO_1507 (O_1507,N_14959,N_14965);
or UO_1508 (O_1508,N_14948,N_14813);
nand UO_1509 (O_1509,N_14896,N_14826);
xor UO_1510 (O_1510,N_14959,N_14945);
xnor UO_1511 (O_1511,N_14962,N_14792);
or UO_1512 (O_1512,N_14898,N_14801);
nand UO_1513 (O_1513,N_14878,N_14795);
or UO_1514 (O_1514,N_14765,N_14772);
xor UO_1515 (O_1515,N_14960,N_14795);
xor UO_1516 (O_1516,N_14768,N_14827);
xor UO_1517 (O_1517,N_14787,N_14901);
or UO_1518 (O_1518,N_14914,N_14964);
nand UO_1519 (O_1519,N_14873,N_14857);
xnor UO_1520 (O_1520,N_14845,N_14854);
nor UO_1521 (O_1521,N_14947,N_14927);
or UO_1522 (O_1522,N_14960,N_14811);
or UO_1523 (O_1523,N_14918,N_14817);
xor UO_1524 (O_1524,N_14836,N_14922);
nand UO_1525 (O_1525,N_14873,N_14917);
or UO_1526 (O_1526,N_14758,N_14786);
and UO_1527 (O_1527,N_14807,N_14882);
nor UO_1528 (O_1528,N_14973,N_14875);
and UO_1529 (O_1529,N_14840,N_14924);
nand UO_1530 (O_1530,N_14880,N_14770);
nand UO_1531 (O_1531,N_14989,N_14786);
nor UO_1532 (O_1532,N_14959,N_14921);
and UO_1533 (O_1533,N_14966,N_14900);
nand UO_1534 (O_1534,N_14818,N_14829);
nand UO_1535 (O_1535,N_14864,N_14992);
or UO_1536 (O_1536,N_14933,N_14918);
or UO_1537 (O_1537,N_14923,N_14987);
nand UO_1538 (O_1538,N_14962,N_14825);
nand UO_1539 (O_1539,N_14954,N_14850);
or UO_1540 (O_1540,N_14881,N_14934);
xnor UO_1541 (O_1541,N_14806,N_14938);
and UO_1542 (O_1542,N_14858,N_14759);
or UO_1543 (O_1543,N_14768,N_14764);
nand UO_1544 (O_1544,N_14868,N_14876);
or UO_1545 (O_1545,N_14780,N_14896);
xor UO_1546 (O_1546,N_14822,N_14851);
nand UO_1547 (O_1547,N_14805,N_14881);
and UO_1548 (O_1548,N_14983,N_14775);
xor UO_1549 (O_1549,N_14800,N_14758);
xnor UO_1550 (O_1550,N_14856,N_14844);
nor UO_1551 (O_1551,N_14844,N_14837);
nor UO_1552 (O_1552,N_14874,N_14765);
nand UO_1553 (O_1553,N_14999,N_14786);
or UO_1554 (O_1554,N_14996,N_14940);
and UO_1555 (O_1555,N_14863,N_14829);
and UO_1556 (O_1556,N_14815,N_14950);
nand UO_1557 (O_1557,N_14922,N_14888);
and UO_1558 (O_1558,N_14878,N_14969);
xor UO_1559 (O_1559,N_14953,N_14898);
nor UO_1560 (O_1560,N_14916,N_14965);
nor UO_1561 (O_1561,N_14859,N_14803);
xor UO_1562 (O_1562,N_14955,N_14805);
and UO_1563 (O_1563,N_14958,N_14768);
nor UO_1564 (O_1564,N_14943,N_14788);
xor UO_1565 (O_1565,N_14847,N_14804);
or UO_1566 (O_1566,N_14950,N_14876);
nor UO_1567 (O_1567,N_14782,N_14971);
and UO_1568 (O_1568,N_14829,N_14880);
and UO_1569 (O_1569,N_14768,N_14795);
nand UO_1570 (O_1570,N_14894,N_14950);
nand UO_1571 (O_1571,N_14894,N_14935);
or UO_1572 (O_1572,N_14787,N_14768);
nor UO_1573 (O_1573,N_14896,N_14774);
xor UO_1574 (O_1574,N_14990,N_14750);
and UO_1575 (O_1575,N_14813,N_14976);
or UO_1576 (O_1576,N_14944,N_14788);
xnor UO_1577 (O_1577,N_14834,N_14778);
nand UO_1578 (O_1578,N_14975,N_14885);
nor UO_1579 (O_1579,N_14977,N_14763);
or UO_1580 (O_1580,N_14831,N_14852);
or UO_1581 (O_1581,N_14881,N_14944);
or UO_1582 (O_1582,N_14959,N_14994);
or UO_1583 (O_1583,N_14851,N_14948);
and UO_1584 (O_1584,N_14881,N_14833);
nor UO_1585 (O_1585,N_14968,N_14808);
or UO_1586 (O_1586,N_14802,N_14962);
and UO_1587 (O_1587,N_14863,N_14789);
nand UO_1588 (O_1588,N_14895,N_14904);
nor UO_1589 (O_1589,N_14950,N_14770);
nand UO_1590 (O_1590,N_14771,N_14799);
nor UO_1591 (O_1591,N_14939,N_14849);
xnor UO_1592 (O_1592,N_14932,N_14876);
nand UO_1593 (O_1593,N_14995,N_14810);
or UO_1594 (O_1594,N_14937,N_14786);
and UO_1595 (O_1595,N_14832,N_14766);
or UO_1596 (O_1596,N_14939,N_14760);
nor UO_1597 (O_1597,N_14754,N_14909);
nor UO_1598 (O_1598,N_14964,N_14882);
xnor UO_1599 (O_1599,N_14906,N_14892);
or UO_1600 (O_1600,N_14956,N_14779);
nand UO_1601 (O_1601,N_14902,N_14927);
and UO_1602 (O_1602,N_14947,N_14768);
or UO_1603 (O_1603,N_14961,N_14823);
and UO_1604 (O_1604,N_14830,N_14962);
nor UO_1605 (O_1605,N_14934,N_14864);
xnor UO_1606 (O_1606,N_14931,N_14804);
nor UO_1607 (O_1607,N_14961,N_14928);
xnor UO_1608 (O_1608,N_14920,N_14969);
nor UO_1609 (O_1609,N_14853,N_14836);
xnor UO_1610 (O_1610,N_14931,N_14752);
or UO_1611 (O_1611,N_14906,N_14781);
nor UO_1612 (O_1612,N_14981,N_14931);
or UO_1613 (O_1613,N_14983,N_14807);
nand UO_1614 (O_1614,N_14821,N_14797);
or UO_1615 (O_1615,N_14919,N_14879);
and UO_1616 (O_1616,N_14984,N_14960);
or UO_1617 (O_1617,N_14771,N_14996);
or UO_1618 (O_1618,N_14970,N_14892);
and UO_1619 (O_1619,N_14912,N_14809);
nor UO_1620 (O_1620,N_14824,N_14925);
nor UO_1621 (O_1621,N_14956,N_14939);
nor UO_1622 (O_1622,N_14934,N_14867);
xor UO_1623 (O_1623,N_14908,N_14858);
nor UO_1624 (O_1624,N_14959,N_14848);
and UO_1625 (O_1625,N_14999,N_14898);
nand UO_1626 (O_1626,N_14925,N_14997);
and UO_1627 (O_1627,N_14767,N_14955);
or UO_1628 (O_1628,N_14989,N_14931);
and UO_1629 (O_1629,N_14904,N_14938);
nor UO_1630 (O_1630,N_14828,N_14800);
nor UO_1631 (O_1631,N_14795,N_14891);
nand UO_1632 (O_1632,N_14983,N_14792);
or UO_1633 (O_1633,N_14939,N_14996);
or UO_1634 (O_1634,N_14876,N_14990);
or UO_1635 (O_1635,N_14908,N_14835);
xor UO_1636 (O_1636,N_14908,N_14900);
and UO_1637 (O_1637,N_14750,N_14966);
xor UO_1638 (O_1638,N_14762,N_14857);
xnor UO_1639 (O_1639,N_14848,N_14874);
xor UO_1640 (O_1640,N_14909,N_14806);
or UO_1641 (O_1641,N_14876,N_14975);
nand UO_1642 (O_1642,N_14931,N_14779);
and UO_1643 (O_1643,N_14994,N_14757);
or UO_1644 (O_1644,N_14786,N_14825);
nand UO_1645 (O_1645,N_14922,N_14871);
and UO_1646 (O_1646,N_14798,N_14970);
nand UO_1647 (O_1647,N_14754,N_14860);
nand UO_1648 (O_1648,N_14847,N_14870);
or UO_1649 (O_1649,N_14761,N_14783);
or UO_1650 (O_1650,N_14950,N_14795);
nand UO_1651 (O_1651,N_14877,N_14910);
or UO_1652 (O_1652,N_14819,N_14792);
nor UO_1653 (O_1653,N_14885,N_14968);
and UO_1654 (O_1654,N_14895,N_14939);
xnor UO_1655 (O_1655,N_14750,N_14982);
nor UO_1656 (O_1656,N_14832,N_14953);
and UO_1657 (O_1657,N_14811,N_14847);
and UO_1658 (O_1658,N_14890,N_14918);
nand UO_1659 (O_1659,N_14889,N_14986);
nor UO_1660 (O_1660,N_14884,N_14940);
xnor UO_1661 (O_1661,N_14787,N_14823);
and UO_1662 (O_1662,N_14937,N_14949);
or UO_1663 (O_1663,N_14863,N_14802);
nor UO_1664 (O_1664,N_14802,N_14793);
xor UO_1665 (O_1665,N_14921,N_14957);
nor UO_1666 (O_1666,N_14975,N_14901);
or UO_1667 (O_1667,N_14960,N_14934);
nor UO_1668 (O_1668,N_14868,N_14893);
or UO_1669 (O_1669,N_14826,N_14914);
xor UO_1670 (O_1670,N_14920,N_14818);
or UO_1671 (O_1671,N_14865,N_14933);
nand UO_1672 (O_1672,N_14754,N_14892);
and UO_1673 (O_1673,N_14949,N_14918);
nor UO_1674 (O_1674,N_14930,N_14814);
and UO_1675 (O_1675,N_14965,N_14937);
and UO_1676 (O_1676,N_14803,N_14895);
nor UO_1677 (O_1677,N_14806,N_14837);
or UO_1678 (O_1678,N_14802,N_14967);
nor UO_1679 (O_1679,N_14886,N_14970);
and UO_1680 (O_1680,N_14863,N_14937);
nand UO_1681 (O_1681,N_14786,N_14785);
or UO_1682 (O_1682,N_14977,N_14802);
and UO_1683 (O_1683,N_14873,N_14872);
or UO_1684 (O_1684,N_14877,N_14813);
xnor UO_1685 (O_1685,N_14854,N_14952);
xnor UO_1686 (O_1686,N_14969,N_14875);
or UO_1687 (O_1687,N_14990,N_14811);
nand UO_1688 (O_1688,N_14818,N_14809);
or UO_1689 (O_1689,N_14798,N_14759);
or UO_1690 (O_1690,N_14849,N_14797);
xor UO_1691 (O_1691,N_14755,N_14851);
xnor UO_1692 (O_1692,N_14921,N_14815);
nand UO_1693 (O_1693,N_14964,N_14968);
nand UO_1694 (O_1694,N_14940,N_14959);
or UO_1695 (O_1695,N_14955,N_14851);
xnor UO_1696 (O_1696,N_14852,N_14980);
nor UO_1697 (O_1697,N_14768,N_14813);
nand UO_1698 (O_1698,N_14781,N_14787);
xnor UO_1699 (O_1699,N_14921,N_14826);
or UO_1700 (O_1700,N_14759,N_14777);
xnor UO_1701 (O_1701,N_14751,N_14952);
nor UO_1702 (O_1702,N_14988,N_14835);
or UO_1703 (O_1703,N_14937,N_14987);
or UO_1704 (O_1704,N_14860,N_14904);
or UO_1705 (O_1705,N_14944,N_14836);
or UO_1706 (O_1706,N_14899,N_14892);
nand UO_1707 (O_1707,N_14788,N_14969);
nand UO_1708 (O_1708,N_14756,N_14976);
nand UO_1709 (O_1709,N_14823,N_14813);
nand UO_1710 (O_1710,N_14793,N_14948);
nor UO_1711 (O_1711,N_14966,N_14921);
nor UO_1712 (O_1712,N_14916,N_14987);
or UO_1713 (O_1713,N_14806,N_14784);
xor UO_1714 (O_1714,N_14792,N_14779);
xnor UO_1715 (O_1715,N_14974,N_14778);
or UO_1716 (O_1716,N_14773,N_14857);
nand UO_1717 (O_1717,N_14971,N_14816);
or UO_1718 (O_1718,N_14772,N_14875);
and UO_1719 (O_1719,N_14981,N_14755);
or UO_1720 (O_1720,N_14926,N_14981);
xor UO_1721 (O_1721,N_14988,N_14758);
nor UO_1722 (O_1722,N_14840,N_14761);
nand UO_1723 (O_1723,N_14957,N_14777);
xor UO_1724 (O_1724,N_14998,N_14880);
and UO_1725 (O_1725,N_14882,N_14930);
and UO_1726 (O_1726,N_14923,N_14941);
and UO_1727 (O_1727,N_14812,N_14766);
nor UO_1728 (O_1728,N_14798,N_14960);
nand UO_1729 (O_1729,N_14767,N_14846);
or UO_1730 (O_1730,N_14968,N_14931);
xnor UO_1731 (O_1731,N_14853,N_14900);
and UO_1732 (O_1732,N_14755,N_14922);
or UO_1733 (O_1733,N_14954,N_14891);
nor UO_1734 (O_1734,N_14971,N_14802);
and UO_1735 (O_1735,N_14779,N_14861);
or UO_1736 (O_1736,N_14780,N_14944);
and UO_1737 (O_1737,N_14956,N_14944);
or UO_1738 (O_1738,N_14936,N_14987);
nand UO_1739 (O_1739,N_14897,N_14954);
nor UO_1740 (O_1740,N_14845,N_14827);
or UO_1741 (O_1741,N_14870,N_14941);
and UO_1742 (O_1742,N_14958,N_14973);
or UO_1743 (O_1743,N_14906,N_14769);
nor UO_1744 (O_1744,N_14822,N_14775);
and UO_1745 (O_1745,N_14798,N_14837);
and UO_1746 (O_1746,N_14865,N_14818);
and UO_1747 (O_1747,N_14982,N_14830);
or UO_1748 (O_1748,N_14882,N_14825);
nor UO_1749 (O_1749,N_14953,N_14946);
or UO_1750 (O_1750,N_14977,N_14929);
xor UO_1751 (O_1751,N_14890,N_14978);
nor UO_1752 (O_1752,N_14953,N_14879);
and UO_1753 (O_1753,N_14987,N_14841);
and UO_1754 (O_1754,N_14881,N_14819);
xnor UO_1755 (O_1755,N_14961,N_14795);
xor UO_1756 (O_1756,N_14809,N_14855);
nand UO_1757 (O_1757,N_14777,N_14985);
or UO_1758 (O_1758,N_14776,N_14902);
or UO_1759 (O_1759,N_14918,N_14943);
xor UO_1760 (O_1760,N_14822,N_14762);
or UO_1761 (O_1761,N_14877,N_14769);
nor UO_1762 (O_1762,N_14898,N_14796);
or UO_1763 (O_1763,N_14783,N_14880);
and UO_1764 (O_1764,N_14914,N_14831);
nor UO_1765 (O_1765,N_14866,N_14847);
or UO_1766 (O_1766,N_14866,N_14772);
and UO_1767 (O_1767,N_14783,N_14914);
or UO_1768 (O_1768,N_14855,N_14825);
nor UO_1769 (O_1769,N_14902,N_14787);
xnor UO_1770 (O_1770,N_14961,N_14904);
and UO_1771 (O_1771,N_14903,N_14788);
or UO_1772 (O_1772,N_14829,N_14764);
or UO_1773 (O_1773,N_14953,N_14800);
nor UO_1774 (O_1774,N_14979,N_14836);
nand UO_1775 (O_1775,N_14939,N_14866);
xor UO_1776 (O_1776,N_14797,N_14776);
nand UO_1777 (O_1777,N_14877,N_14937);
and UO_1778 (O_1778,N_14756,N_14944);
nand UO_1779 (O_1779,N_14782,N_14936);
or UO_1780 (O_1780,N_14873,N_14996);
nor UO_1781 (O_1781,N_14886,N_14808);
or UO_1782 (O_1782,N_14836,N_14760);
nor UO_1783 (O_1783,N_14939,N_14817);
or UO_1784 (O_1784,N_14861,N_14938);
and UO_1785 (O_1785,N_14901,N_14819);
or UO_1786 (O_1786,N_14784,N_14824);
and UO_1787 (O_1787,N_14774,N_14960);
xor UO_1788 (O_1788,N_14966,N_14858);
and UO_1789 (O_1789,N_14817,N_14789);
or UO_1790 (O_1790,N_14951,N_14857);
nor UO_1791 (O_1791,N_14816,N_14851);
and UO_1792 (O_1792,N_14984,N_14871);
nand UO_1793 (O_1793,N_14946,N_14991);
or UO_1794 (O_1794,N_14863,N_14760);
nor UO_1795 (O_1795,N_14969,N_14931);
xnor UO_1796 (O_1796,N_14946,N_14800);
nor UO_1797 (O_1797,N_14836,N_14809);
xnor UO_1798 (O_1798,N_14953,N_14803);
nor UO_1799 (O_1799,N_14896,N_14859);
nand UO_1800 (O_1800,N_14934,N_14823);
xnor UO_1801 (O_1801,N_14837,N_14999);
nand UO_1802 (O_1802,N_14872,N_14917);
or UO_1803 (O_1803,N_14905,N_14786);
or UO_1804 (O_1804,N_14753,N_14938);
or UO_1805 (O_1805,N_14846,N_14805);
xnor UO_1806 (O_1806,N_14918,N_14938);
nor UO_1807 (O_1807,N_14989,N_14886);
xor UO_1808 (O_1808,N_14931,N_14782);
and UO_1809 (O_1809,N_14853,N_14804);
nand UO_1810 (O_1810,N_14920,N_14758);
or UO_1811 (O_1811,N_14967,N_14905);
or UO_1812 (O_1812,N_14767,N_14833);
and UO_1813 (O_1813,N_14872,N_14974);
or UO_1814 (O_1814,N_14937,N_14915);
and UO_1815 (O_1815,N_14817,N_14912);
xor UO_1816 (O_1816,N_14975,N_14894);
nand UO_1817 (O_1817,N_14931,N_14926);
nor UO_1818 (O_1818,N_14890,N_14781);
and UO_1819 (O_1819,N_14797,N_14787);
nor UO_1820 (O_1820,N_14985,N_14995);
or UO_1821 (O_1821,N_14889,N_14857);
nor UO_1822 (O_1822,N_14936,N_14765);
or UO_1823 (O_1823,N_14900,N_14983);
nand UO_1824 (O_1824,N_14887,N_14987);
and UO_1825 (O_1825,N_14757,N_14920);
nor UO_1826 (O_1826,N_14805,N_14917);
and UO_1827 (O_1827,N_14834,N_14774);
xor UO_1828 (O_1828,N_14961,N_14967);
and UO_1829 (O_1829,N_14766,N_14942);
nand UO_1830 (O_1830,N_14898,N_14969);
and UO_1831 (O_1831,N_14993,N_14851);
and UO_1832 (O_1832,N_14886,N_14974);
and UO_1833 (O_1833,N_14918,N_14940);
and UO_1834 (O_1834,N_14778,N_14787);
and UO_1835 (O_1835,N_14781,N_14892);
or UO_1836 (O_1836,N_14904,N_14771);
or UO_1837 (O_1837,N_14782,N_14900);
nor UO_1838 (O_1838,N_14785,N_14760);
nor UO_1839 (O_1839,N_14794,N_14934);
xnor UO_1840 (O_1840,N_14916,N_14945);
or UO_1841 (O_1841,N_14881,N_14980);
nor UO_1842 (O_1842,N_14950,N_14865);
nand UO_1843 (O_1843,N_14791,N_14934);
xnor UO_1844 (O_1844,N_14860,N_14911);
and UO_1845 (O_1845,N_14937,N_14927);
or UO_1846 (O_1846,N_14778,N_14894);
or UO_1847 (O_1847,N_14937,N_14872);
nand UO_1848 (O_1848,N_14975,N_14869);
nor UO_1849 (O_1849,N_14810,N_14863);
nor UO_1850 (O_1850,N_14863,N_14839);
xor UO_1851 (O_1851,N_14911,N_14870);
and UO_1852 (O_1852,N_14944,N_14878);
and UO_1853 (O_1853,N_14897,N_14791);
nor UO_1854 (O_1854,N_14965,N_14807);
nor UO_1855 (O_1855,N_14817,N_14992);
nor UO_1856 (O_1856,N_14931,N_14759);
nor UO_1857 (O_1857,N_14986,N_14916);
or UO_1858 (O_1858,N_14823,N_14827);
nand UO_1859 (O_1859,N_14935,N_14768);
and UO_1860 (O_1860,N_14863,N_14832);
nand UO_1861 (O_1861,N_14853,N_14872);
nor UO_1862 (O_1862,N_14770,N_14918);
or UO_1863 (O_1863,N_14798,N_14829);
nor UO_1864 (O_1864,N_14887,N_14892);
nand UO_1865 (O_1865,N_14898,N_14929);
or UO_1866 (O_1866,N_14933,N_14788);
xor UO_1867 (O_1867,N_14927,N_14847);
or UO_1868 (O_1868,N_14957,N_14988);
and UO_1869 (O_1869,N_14970,N_14964);
and UO_1870 (O_1870,N_14798,N_14799);
or UO_1871 (O_1871,N_14872,N_14928);
xnor UO_1872 (O_1872,N_14882,N_14939);
nor UO_1873 (O_1873,N_14921,N_14753);
nand UO_1874 (O_1874,N_14918,N_14828);
nor UO_1875 (O_1875,N_14897,N_14761);
nor UO_1876 (O_1876,N_14847,N_14797);
xor UO_1877 (O_1877,N_14872,N_14772);
nor UO_1878 (O_1878,N_14846,N_14983);
nand UO_1879 (O_1879,N_14891,N_14824);
nand UO_1880 (O_1880,N_14788,N_14765);
xor UO_1881 (O_1881,N_14956,N_14775);
xor UO_1882 (O_1882,N_14989,N_14835);
or UO_1883 (O_1883,N_14794,N_14807);
xor UO_1884 (O_1884,N_14843,N_14891);
and UO_1885 (O_1885,N_14764,N_14885);
or UO_1886 (O_1886,N_14821,N_14866);
or UO_1887 (O_1887,N_14985,N_14795);
xor UO_1888 (O_1888,N_14919,N_14930);
nand UO_1889 (O_1889,N_14863,N_14983);
nand UO_1890 (O_1890,N_14831,N_14964);
xor UO_1891 (O_1891,N_14846,N_14994);
and UO_1892 (O_1892,N_14772,N_14832);
xnor UO_1893 (O_1893,N_14980,N_14977);
and UO_1894 (O_1894,N_14974,N_14966);
nor UO_1895 (O_1895,N_14842,N_14818);
xnor UO_1896 (O_1896,N_14858,N_14762);
and UO_1897 (O_1897,N_14784,N_14919);
and UO_1898 (O_1898,N_14840,N_14931);
nor UO_1899 (O_1899,N_14936,N_14916);
or UO_1900 (O_1900,N_14948,N_14777);
nor UO_1901 (O_1901,N_14920,N_14919);
xor UO_1902 (O_1902,N_14822,N_14961);
or UO_1903 (O_1903,N_14759,N_14991);
or UO_1904 (O_1904,N_14850,N_14752);
or UO_1905 (O_1905,N_14813,N_14847);
xor UO_1906 (O_1906,N_14903,N_14997);
and UO_1907 (O_1907,N_14905,N_14941);
xor UO_1908 (O_1908,N_14867,N_14767);
and UO_1909 (O_1909,N_14771,N_14909);
nor UO_1910 (O_1910,N_14762,N_14921);
or UO_1911 (O_1911,N_14972,N_14921);
and UO_1912 (O_1912,N_14891,N_14886);
and UO_1913 (O_1913,N_14784,N_14955);
nand UO_1914 (O_1914,N_14944,N_14877);
nand UO_1915 (O_1915,N_14832,N_14946);
nor UO_1916 (O_1916,N_14897,N_14856);
or UO_1917 (O_1917,N_14796,N_14984);
nand UO_1918 (O_1918,N_14861,N_14824);
or UO_1919 (O_1919,N_14778,N_14784);
or UO_1920 (O_1920,N_14998,N_14791);
or UO_1921 (O_1921,N_14859,N_14945);
xnor UO_1922 (O_1922,N_14815,N_14805);
nor UO_1923 (O_1923,N_14820,N_14818);
or UO_1924 (O_1924,N_14764,N_14844);
or UO_1925 (O_1925,N_14962,N_14878);
xnor UO_1926 (O_1926,N_14911,N_14944);
xnor UO_1927 (O_1927,N_14838,N_14791);
and UO_1928 (O_1928,N_14769,N_14965);
and UO_1929 (O_1929,N_14810,N_14856);
xnor UO_1930 (O_1930,N_14995,N_14873);
nor UO_1931 (O_1931,N_14817,N_14927);
or UO_1932 (O_1932,N_14915,N_14839);
and UO_1933 (O_1933,N_14927,N_14891);
nor UO_1934 (O_1934,N_14795,N_14871);
xor UO_1935 (O_1935,N_14752,N_14815);
nor UO_1936 (O_1936,N_14786,N_14818);
nand UO_1937 (O_1937,N_14872,N_14781);
or UO_1938 (O_1938,N_14860,N_14862);
or UO_1939 (O_1939,N_14993,N_14989);
and UO_1940 (O_1940,N_14832,N_14866);
and UO_1941 (O_1941,N_14822,N_14849);
and UO_1942 (O_1942,N_14860,N_14805);
and UO_1943 (O_1943,N_14885,N_14807);
nor UO_1944 (O_1944,N_14805,N_14964);
or UO_1945 (O_1945,N_14955,N_14995);
and UO_1946 (O_1946,N_14917,N_14847);
and UO_1947 (O_1947,N_14902,N_14891);
xor UO_1948 (O_1948,N_14945,N_14766);
or UO_1949 (O_1949,N_14751,N_14863);
nor UO_1950 (O_1950,N_14763,N_14845);
and UO_1951 (O_1951,N_14948,N_14956);
nand UO_1952 (O_1952,N_14967,N_14757);
nor UO_1953 (O_1953,N_14886,N_14782);
nand UO_1954 (O_1954,N_14904,N_14795);
nand UO_1955 (O_1955,N_14835,N_14896);
or UO_1956 (O_1956,N_14796,N_14820);
or UO_1957 (O_1957,N_14763,N_14971);
or UO_1958 (O_1958,N_14843,N_14987);
nor UO_1959 (O_1959,N_14907,N_14768);
xnor UO_1960 (O_1960,N_14907,N_14774);
or UO_1961 (O_1961,N_14830,N_14926);
and UO_1962 (O_1962,N_14931,N_14952);
xnor UO_1963 (O_1963,N_14995,N_14874);
and UO_1964 (O_1964,N_14963,N_14924);
or UO_1965 (O_1965,N_14774,N_14971);
nor UO_1966 (O_1966,N_14839,N_14984);
xnor UO_1967 (O_1967,N_14834,N_14773);
nor UO_1968 (O_1968,N_14898,N_14820);
and UO_1969 (O_1969,N_14903,N_14843);
or UO_1970 (O_1970,N_14897,N_14777);
or UO_1971 (O_1971,N_14770,N_14942);
or UO_1972 (O_1972,N_14888,N_14968);
or UO_1973 (O_1973,N_14952,N_14903);
xor UO_1974 (O_1974,N_14955,N_14810);
and UO_1975 (O_1975,N_14851,N_14854);
and UO_1976 (O_1976,N_14934,N_14770);
nand UO_1977 (O_1977,N_14831,N_14910);
and UO_1978 (O_1978,N_14954,N_14962);
xnor UO_1979 (O_1979,N_14769,N_14758);
xor UO_1980 (O_1980,N_14883,N_14789);
nand UO_1981 (O_1981,N_14911,N_14828);
nor UO_1982 (O_1982,N_14763,N_14914);
nor UO_1983 (O_1983,N_14942,N_14958);
nand UO_1984 (O_1984,N_14778,N_14825);
and UO_1985 (O_1985,N_14973,N_14832);
and UO_1986 (O_1986,N_14919,N_14992);
nor UO_1987 (O_1987,N_14838,N_14946);
and UO_1988 (O_1988,N_14968,N_14922);
nand UO_1989 (O_1989,N_14905,N_14933);
xnor UO_1990 (O_1990,N_14881,N_14917);
and UO_1991 (O_1991,N_14782,N_14867);
nor UO_1992 (O_1992,N_14909,N_14804);
xor UO_1993 (O_1993,N_14954,N_14892);
and UO_1994 (O_1994,N_14986,N_14935);
and UO_1995 (O_1995,N_14902,N_14772);
xor UO_1996 (O_1996,N_14810,N_14840);
nor UO_1997 (O_1997,N_14790,N_14889);
nand UO_1998 (O_1998,N_14859,N_14827);
xor UO_1999 (O_1999,N_14759,N_14959);
endmodule