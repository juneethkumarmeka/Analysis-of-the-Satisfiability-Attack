module basic_1000_10000_1500_100_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_128,In_967);
nand U1 (N_1,In_309,In_337);
or U2 (N_2,In_936,In_778);
xor U3 (N_3,In_360,In_501);
or U4 (N_4,In_493,In_849);
or U5 (N_5,In_614,In_41);
nor U6 (N_6,In_701,In_476);
or U7 (N_7,In_974,In_540);
nand U8 (N_8,In_503,In_740);
xor U9 (N_9,In_607,In_66);
or U10 (N_10,In_353,In_277);
nor U11 (N_11,In_755,In_334);
nand U12 (N_12,In_642,In_261);
and U13 (N_13,In_662,In_904);
nand U14 (N_14,In_224,In_997);
or U15 (N_15,In_907,In_706);
nand U16 (N_16,In_980,In_566);
nor U17 (N_17,In_843,In_91);
or U18 (N_18,In_690,In_44);
and U19 (N_19,In_258,In_373);
nand U20 (N_20,In_223,In_657);
xnor U21 (N_21,In_775,In_653);
nand U22 (N_22,In_663,In_20);
and U23 (N_23,In_547,In_754);
and U24 (N_24,In_675,In_921);
nor U25 (N_25,In_227,In_641);
nor U26 (N_26,In_941,In_85);
nor U27 (N_27,In_718,In_576);
nor U28 (N_28,In_589,In_875);
nor U29 (N_29,In_909,In_363);
or U30 (N_30,In_317,In_749);
xnor U31 (N_31,In_435,In_487);
nand U32 (N_32,In_187,In_113);
nor U33 (N_33,In_922,In_463);
and U34 (N_34,In_88,In_715);
nor U35 (N_35,In_957,In_179);
and U36 (N_36,In_897,In_382);
xnor U37 (N_37,In_616,In_838);
and U38 (N_38,In_876,In_119);
or U39 (N_39,In_711,In_863);
xor U40 (N_40,In_573,In_455);
and U41 (N_41,In_162,In_692);
nand U42 (N_42,In_955,In_564);
nand U43 (N_43,In_61,In_206);
nand U44 (N_44,In_6,In_438);
nand U45 (N_45,In_171,In_443);
nor U46 (N_46,In_60,In_143);
nor U47 (N_47,In_504,In_893);
xnor U48 (N_48,In_526,In_31);
or U49 (N_49,In_979,In_43);
or U50 (N_50,In_195,In_857);
or U51 (N_51,In_35,In_599);
xor U52 (N_52,In_0,In_376);
nor U53 (N_53,In_877,In_931);
and U54 (N_54,In_355,In_439);
and U55 (N_55,In_622,In_134);
nor U56 (N_56,In_329,In_627);
nand U57 (N_57,In_82,In_617);
xnor U58 (N_58,In_42,In_318);
and U59 (N_59,In_603,In_252);
or U60 (N_60,In_47,In_530);
xnor U61 (N_61,In_864,In_766);
or U62 (N_62,In_746,In_466);
or U63 (N_63,In_80,In_413);
nand U64 (N_64,In_159,In_770);
or U65 (N_65,In_805,In_968);
nand U66 (N_66,In_279,In_551);
or U67 (N_67,In_804,In_291);
or U68 (N_68,In_668,In_231);
and U69 (N_69,In_519,In_781);
or U70 (N_70,In_685,In_944);
and U71 (N_71,In_584,In_776);
xnor U72 (N_72,In_90,In_570);
or U73 (N_73,In_300,In_483);
or U74 (N_74,In_824,In_216);
and U75 (N_75,In_215,In_816);
and U76 (N_76,In_889,In_76);
nor U77 (N_77,In_544,In_673);
nor U78 (N_78,In_797,In_415);
and U79 (N_79,In_823,In_288);
or U80 (N_80,In_319,In_722);
or U81 (N_81,In_52,In_428);
or U82 (N_82,In_704,In_578);
xor U83 (N_83,In_315,In_490);
nor U84 (N_84,In_624,In_575);
or U85 (N_85,In_267,In_995);
xor U86 (N_86,In_144,In_730);
nor U87 (N_87,In_124,In_537);
xnor U88 (N_88,In_62,In_700);
xor U89 (N_89,In_507,In_266);
or U90 (N_90,In_935,In_946);
or U91 (N_91,In_713,In_422);
nand U92 (N_92,In_157,In_989);
and U93 (N_93,In_965,In_757);
nand U94 (N_94,In_99,In_985);
or U95 (N_95,In_421,In_745);
nor U96 (N_96,In_812,In_939);
nor U97 (N_97,In_908,In_753);
nand U98 (N_98,In_120,In_192);
nand U99 (N_99,In_744,In_556);
xor U100 (N_100,In_901,In_53);
or U101 (N_101,In_238,In_964);
xnor U102 (N_102,In_358,In_664);
xnor U103 (N_103,In_883,In_105);
xor U104 (N_104,N_46,In_264);
or U105 (N_105,N_49,In_869);
and U106 (N_106,N_36,In_139);
nand U107 (N_107,In_170,In_212);
nor U108 (N_108,In_514,In_987);
and U109 (N_109,In_669,In_709);
and U110 (N_110,N_42,In_316);
or U111 (N_111,In_714,In_176);
or U112 (N_112,In_406,In_462);
nor U113 (N_113,In_969,In_445);
xnor U114 (N_114,In_56,In_209);
nand U115 (N_115,In_705,In_188);
nand U116 (N_116,N_69,In_465);
xor U117 (N_117,N_51,In_411);
xnor U118 (N_118,In_178,In_395);
nand U119 (N_119,In_542,In_531);
or U120 (N_120,In_74,In_986);
or U121 (N_121,In_257,In_844);
and U122 (N_122,In_23,N_31);
nand U123 (N_123,In_464,In_879);
or U124 (N_124,In_236,In_506);
and U125 (N_125,In_520,In_761);
or U126 (N_126,In_107,In_423);
xnor U127 (N_127,N_22,In_583);
or U128 (N_128,In_330,In_482);
and U129 (N_129,N_18,In_86);
xnor U130 (N_130,In_436,In_136);
or U131 (N_131,In_480,In_815);
nor U132 (N_132,In_429,In_63);
nor U133 (N_133,N_84,In_882);
nand U134 (N_134,In_220,In_141);
and U135 (N_135,In_574,N_87);
xor U136 (N_136,In_135,In_733);
and U137 (N_137,In_903,In_860);
xor U138 (N_138,In_381,In_517);
nand U139 (N_139,In_446,In_425);
nor U140 (N_140,In_580,In_801);
xnor U141 (N_141,In_920,In_226);
or U142 (N_142,In_160,In_407);
nor U143 (N_143,In_15,In_95);
xor U144 (N_144,In_659,In_453);
nor U145 (N_145,In_509,In_405);
nor U146 (N_146,In_768,In_836);
nand U147 (N_147,In_73,In_481);
or U148 (N_148,In_327,In_630);
nor U149 (N_149,In_606,In_285);
and U150 (N_150,In_132,In_822);
or U151 (N_151,N_2,In_756);
or U152 (N_152,In_270,In_966);
nor U153 (N_153,In_283,N_73);
xor U154 (N_154,In_835,In_803);
xnor U155 (N_155,In_655,In_208);
xnor U156 (N_156,In_568,In_829);
nor U157 (N_157,N_65,In_621);
xor U158 (N_158,In_658,In_281);
nand U159 (N_159,N_60,In_345);
nor U160 (N_160,In_189,In_978);
nor U161 (N_161,In_241,In_271);
and U162 (N_162,In_919,In_456);
or U163 (N_163,In_981,In_728);
nand U164 (N_164,In_100,In_467);
nand U165 (N_165,In_69,N_92);
or U166 (N_166,In_37,In_102);
nor U167 (N_167,In_497,In_249);
nor U168 (N_168,In_856,In_523);
nand U169 (N_169,In_579,In_620);
xor U170 (N_170,In_228,N_4);
xnor U171 (N_171,In_320,In_810);
nor U172 (N_172,In_340,In_555);
xnor U173 (N_173,In_853,In_888);
and U174 (N_174,In_496,In_268);
or U175 (N_175,In_916,In_764);
or U176 (N_176,In_417,N_50);
or U177 (N_177,In_629,In_350);
nand U178 (N_178,In_992,In_654);
xor U179 (N_179,In_612,In_798);
nor U180 (N_180,In_660,N_85);
and U181 (N_181,N_11,In_543);
or U182 (N_182,In_674,In_656);
and U183 (N_183,In_634,In_50);
and U184 (N_184,In_75,In_821);
nor U185 (N_185,In_221,N_86);
xor U186 (N_186,In_211,In_26);
nor U187 (N_187,In_902,In_683);
or U188 (N_188,In_25,In_284);
xnor U189 (N_189,In_806,In_294);
nor U190 (N_190,In_596,In_973);
or U191 (N_191,In_495,In_956);
and U192 (N_192,In_546,In_585);
nand U193 (N_193,In_516,In_48);
nand U194 (N_194,In_870,In_186);
and U195 (N_195,N_54,In_419);
xnor U196 (N_196,In_292,In_293);
and U197 (N_197,N_35,In_457);
nand U198 (N_198,In_813,In_14);
and U199 (N_199,In_959,In_525);
or U200 (N_200,In_247,In_172);
xor U201 (N_201,N_102,In_377);
and U202 (N_202,In_147,In_891);
or U203 (N_203,In_118,In_106);
nor U204 (N_204,In_13,In_528);
and U205 (N_205,In_522,N_74);
xor U206 (N_206,N_41,In_736);
and U207 (N_207,In_1,In_933);
and U208 (N_208,In_945,In_440);
xor U209 (N_209,In_165,N_197);
nand U210 (N_210,N_117,In_881);
xor U211 (N_211,In_923,In_703);
nand U212 (N_212,N_38,In_333);
xor U213 (N_213,In_512,In_286);
nor U214 (N_214,N_157,N_176);
and U215 (N_215,N_194,In_588);
or U216 (N_216,In_800,In_336);
or U217 (N_217,In_866,In_720);
or U218 (N_218,N_58,In_792);
nand U219 (N_219,In_243,In_785);
xnor U220 (N_220,In_689,In_28);
nand U221 (N_221,In_67,In_420);
or U222 (N_222,In_71,N_133);
nor U223 (N_223,In_133,In_845);
nor U224 (N_224,In_508,In_77);
xnor U225 (N_225,In_202,In_153);
and U226 (N_226,In_748,In_511);
nand U227 (N_227,In_650,In_341);
nor U228 (N_228,In_295,In_479);
or U229 (N_229,In_763,In_87);
and U230 (N_230,In_619,In_94);
nand U231 (N_231,In_623,In_587);
nor U232 (N_232,In_983,N_152);
nand U233 (N_233,In_532,In_533);
and U234 (N_234,In_500,In_808);
xor U235 (N_235,N_83,In_724);
xnor U236 (N_236,N_5,In_262);
nand U237 (N_237,In_717,In_193);
nor U238 (N_238,In_488,In_886);
or U239 (N_239,In_324,In_604);
nor U240 (N_240,In_472,In_460);
xor U241 (N_241,In_129,N_137);
xor U242 (N_242,In_638,In_386);
nor U243 (N_243,In_469,N_120);
nor U244 (N_244,N_195,In_510);
nand U245 (N_245,N_128,In_867);
and U246 (N_246,N_90,In_194);
and U247 (N_247,In_311,In_374);
or U248 (N_248,In_737,N_162);
and U249 (N_249,In_789,N_182);
or U250 (N_250,N_160,In_721);
xor U251 (N_251,In_988,In_833);
nand U252 (N_252,In_637,In_930);
nor U253 (N_253,In_237,In_347);
and U254 (N_254,In_938,In_915);
nor U255 (N_255,In_834,In_93);
xor U256 (N_256,N_139,In_552);
and U257 (N_257,In_592,In_72);
nor U258 (N_258,In_416,N_81);
nor U259 (N_259,In_890,In_926);
nand U260 (N_260,N_122,N_172);
and U261 (N_261,In_557,In_962);
nand U262 (N_262,In_30,In_458);
xor U263 (N_263,In_851,In_847);
or U264 (N_264,In_648,In_747);
and U265 (N_265,In_898,In_68);
xnor U266 (N_266,In_577,In_858);
or U267 (N_267,In_788,In_447);
xnor U268 (N_268,N_13,N_169);
xnor U269 (N_269,In_723,In_871);
or U270 (N_270,In_36,In_913);
and U271 (N_271,In_426,In_151);
nand U272 (N_272,N_184,In_832);
or U273 (N_273,In_280,In_260);
and U274 (N_274,N_193,In_357);
or U275 (N_275,In_887,In_4);
nor U276 (N_276,In_950,In_613);
or U277 (N_277,In_352,N_12);
and U278 (N_278,In_647,N_91);
nor U279 (N_279,In_937,In_394);
and U280 (N_280,In_644,In_817);
xor U281 (N_281,N_75,In_802);
or U282 (N_282,In_49,In_301);
nor U283 (N_283,In_632,In_9);
nand U284 (N_284,In_678,In_168);
and U285 (N_285,In_59,In_492);
xnor U286 (N_286,In_993,N_94);
and U287 (N_287,In_651,In_862);
and U288 (N_288,In_914,In_254);
and U289 (N_289,In_786,In_433);
nor U290 (N_290,In_475,In_399);
nand U291 (N_291,In_698,In_750);
and U292 (N_292,In_84,In_96);
and U293 (N_293,N_143,In_716);
nand U294 (N_294,In_625,N_174);
nor U295 (N_295,N_10,In_586);
nand U296 (N_296,In_296,In_773);
and U297 (N_297,N_1,N_98);
nor U298 (N_298,In_640,In_297);
and U299 (N_299,In_32,In_972);
xnor U300 (N_300,In_470,N_263);
nor U301 (N_301,In_672,N_254);
nor U302 (N_302,In_951,N_97);
xor U303 (N_303,In_807,In_473);
xnor U304 (N_304,In_368,In_484);
xnor U305 (N_305,In_771,In_158);
and U306 (N_306,In_210,In_232);
or U307 (N_307,In_111,In_628);
xnor U308 (N_308,N_181,N_290);
nand U309 (N_309,N_138,In_558);
and U310 (N_310,In_932,N_178);
or U311 (N_311,In_234,In_392);
xor U312 (N_312,In_57,In_767);
or U313 (N_313,N_8,N_222);
xnor U314 (N_314,N_106,In_645);
and U315 (N_315,N_123,In_149);
nand U316 (N_316,N_67,In_38);
xnor U317 (N_317,In_177,N_111);
xor U318 (N_318,In_181,In_200);
nor U319 (N_319,N_141,In_947);
and U320 (N_320,N_32,In_486);
nand U321 (N_321,In_2,N_25);
or U322 (N_322,N_37,N_124);
xnor U323 (N_323,N_244,In_842);
nand U324 (N_324,In_949,In_758);
nand U325 (N_325,In_779,In_454);
nand U326 (N_326,In_375,In_33);
and U327 (N_327,In_554,In_468);
or U328 (N_328,In_404,In_502);
nor U329 (N_329,In_272,In_450);
or U330 (N_330,In_364,In_269);
or U331 (N_331,N_261,N_207);
nand U332 (N_332,N_283,In_975);
and U333 (N_333,In_246,N_223);
or U334 (N_334,N_297,In_852);
nor U335 (N_335,N_72,N_259);
nor U336 (N_336,N_82,In_765);
and U337 (N_337,In_70,In_255);
or U338 (N_338,In_312,In_581);
or U339 (N_339,N_253,In_348);
nor U340 (N_340,In_289,In_342);
nand U341 (N_341,N_24,In_306);
or U342 (N_342,N_226,In_391);
or U343 (N_343,N_14,In_314);
nand U344 (N_344,N_47,N_252);
xor U345 (N_345,N_79,N_295);
nand U346 (N_346,In_150,In_349);
or U347 (N_347,In_710,In_855);
xnor U348 (N_348,N_256,N_258);
nor U349 (N_349,N_21,In_790);
and U350 (N_350,N_232,In_198);
or U351 (N_351,In_225,In_191);
xnor U352 (N_352,N_188,In_796);
xnor U353 (N_353,N_28,N_64);
nand U354 (N_354,N_255,In_524);
nor U355 (N_355,In_250,In_10);
xnor U356 (N_356,N_62,In_777);
nand U357 (N_357,In_811,In_562);
nor U358 (N_358,N_287,N_213);
and U359 (N_359,In_961,In_323);
nor U360 (N_360,In_24,N_156);
nor U361 (N_361,N_291,N_0);
xnor U362 (N_362,In_402,In_365);
nand U363 (N_363,In_505,In_46);
or U364 (N_364,In_884,In_751);
nor U365 (N_365,N_292,In_471);
xnor U366 (N_366,N_245,In_726);
or U367 (N_367,N_148,In_239);
xor U368 (N_368,N_144,In_684);
xnor U369 (N_369,In_741,N_71);
nor U370 (N_370,In_40,In_782);
or U371 (N_371,In_45,In_412);
and U372 (N_372,In_667,N_108);
or U373 (N_373,In_259,In_384);
or U374 (N_374,N_277,N_251);
xnor U375 (N_375,In_990,N_237);
and U376 (N_376,In_18,In_389);
or U377 (N_377,N_228,In_639);
or U378 (N_378,In_708,N_203);
and U379 (N_379,N_170,In_273);
nor U380 (N_380,In_207,In_686);
or U381 (N_381,N_219,In_732);
and U382 (N_382,N_239,In_152);
or U383 (N_383,In_924,In_459);
nand U384 (N_384,In_371,In_928);
or U385 (N_385,In_828,In_98);
nand U386 (N_386,N_149,In_321);
and U387 (N_387,N_250,N_110);
xor U388 (N_388,In_299,In_338);
or U389 (N_389,In_970,In_304);
xnor U390 (N_390,In_122,In_636);
or U391 (N_391,In_991,N_278);
xor U392 (N_392,In_670,In_814);
nor U393 (N_393,N_101,N_44);
nand U394 (N_394,In_276,In_230);
nand U395 (N_395,In_859,In_244);
or U396 (N_396,N_68,N_140);
xor U397 (N_397,In_631,N_167);
or U398 (N_398,N_116,In_848);
or U399 (N_399,In_51,In_489);
or U400 (N_400,N_367,N_201);
or U401 (N_401,In_643,N_381);
and U402 (N_402,N_136,In_372);
or U403 (N_403,In_242,In_680);
nand U404 (N_404,In_665,In_441);
nand U405 (N_405,In_534,In_929);
xnor U406 (N_406,In_560,In_396);
nor U407 (N_407,In_83,In_125);
or U408 (N_408,In_820,In_201);
and U409 (N_409,N_224,N_286);
and U410 (N_410,N_205,N_294);
nor U411 (N_411,In_615,N_389);
or U412 (N_412,In_22,In_335);
nand U413 (N_413,N_374,In_666);
nand U414 (N_414,In_905,N_392);
xor U415 (N_415,N_327,N_177);
and U416 (N_416,In_408,In_769);
and U417 (N_417,In_541,In_245);
xor U418 (N_418,In_954,N_345);
or U419 (N_419,N_88,In_233);
xor U420 (N_420,N_235,N_179);
xor U421 (N_421,In_591,In_403);
nand U422 (N_422,In_203,N_304);
or U423 (N_423,N_293,In_948);
nand U424 (N_424,N_372,In_130);
and U425 (N_425,N_247,In_175);
nand U426 (N_426,In_999,In_205);
or U427 (N_427,N_229,In_952);
nand U428 (N_428,N_6,N_115);
nand U429 (N_429,N_238,In_305);
or U430 (N_430,In_214,N_357);
nand U431 (N_431,In_784,In_12);
or U432 (N_432,In_976,N_164);
and U433 (N_433,N_246,In_894);
xnor U434 (N_434,In_344,N_356);
nand U435 (N_435,N_241,In_608);
nor U436 (N_436,N_302,In_81);
xor U437 (N_437,In_183,In_251);
nand U438 (N_438,In_593,In_166);
nand U439 (N_439,In_16,In_677);
nor U440 (N_440,N_313,N_104);
nor U441 (N_441,N_171,In_444);
nand U442 (N_442,N_121,In_896);
and U443 (N_443,In_248,N_198);
and U444 (N_444,N_383,In_354);
and U445 (N_445,In_11,In_605);
or U446 (N_446,In_64,In_762);
nor U447 (N_447,N_70,In_874);
nor U448 (N_448,N_33,N_29);
nor U449 (N_449,N_388,In_682);
nand U450 (N_450,In_55,N_173);
and U451 (N_451,In_600,N_326);
nor U452 (N_452,In_253,N_394);
xnor U453 (N_453,In_925,N_192);
and U454 (N_454,N_153,In_362);
or U455 (N_455,In_971,N_48);
xor U456 (N_456,N_150,In_671);
xor U457 (N_457,N_234,N_280);
and U458 (N_458,In_691,In_494);
or U459 (N_459,N_270,N_248);
nand U460 (N_460,In_571,In_735);
or U461 (N_461,In_485,In_142);
xnor U462 (N_462,In_731,N_107);
or U463 (N_463,In_256,In_437);
xor U464 (N_464,N_212,N_130);
nor U465 (N_465,In_274,In_114);
nor U466 (N_466,N_257,N_103);
xor U467 (N_467,In_868,In_694);
and U468 (N_468,N_93,In_982);
nor U469 (N_469,N_166,N_366);
nand U470 (N_470,N_307,In_819);
nor U471 (N_471,In_598,N_269);
nor U472 (N_472,In_515,In_21);
and U473 (N_473,N_175,In_567);
xor U474 (N_474,N_3,N_89);
nand U475 (N_475,N_387,In_298);
nand U476 (N_476,N_351,N_373);
xnor U477 (N_477,In_794,N_165);
nand U478 (N_478,In_943,In_182);
or U479 (N_479,In_79,In_760);
and U480 (N_480,In_173,N_40);
and U481 (N_481,N_306,N_320);
xnor U482 (N_482,In_307,N_158);
nor U483 (N_483,In_217,In_213);
or U484 (N_484,N_314,In_388);
xor U485 (N_485,In_934,In_219);
nor U486 (N_486,N_318,N_305);
xor U487 (N_487,In_885,N_66);
nand U488 (N_488,In_958,N_284);
nor U489 (N_489,In_17,In_521);
or U490 (N_490,N_266,N_341);
nor U491 (N_491,N_315,N_19);
or U492 (N_492,N_363,N_159);
or U493 (N_493,N_386,In_313);
nand U494 (N_494,N_114,In_693);
and U495 (N_495,In_89,N_379);
or U496 (N_496,N_183,In_699);
and U497 (N_497,N_322,N_105);
nor U498 (N_498,In_275,In_783);
xor U499 (N_499,In_303,N_303);
xnor U500 (N_500,N_330,In_8);
xor U501 (N_501,In_527,N_63);
nor U502 (N_502,In_795,In_461);
or U503 (N_503,In_652,N_407);
and U504 (N_504,N_488,N_109);
and U505 (N_505,In_618,N_449);
and U506 (N_506,N_384,N_420);
or U507 (N_507,N_99,N_200);
or U508 (N_508,N_23,N_209);
and U509 (N_509,N_397,N_264);
nand U510 (N_510,In_649,In_911);
nand U511 (N_511,N_417,N_344);
nor U512 (N_512,N_456,In_343);
nand U513 (N_513,In_597,In_414);
xor U514 (N_514,N_461,N_249);
nor U515 (N_515,N_355,N_204);
xnor U516 (N_516,In_561,In_799);
xnor U517 (N_517,N_281,In_772);
xnor U518 (N_518,In_553,N_377);
nand U519 (N_519,In_109,N_484);
and U520 (N_520,In_518,In_204);
xnor U521 (N_521,In_190,N_145);
or U522 (N_522,In_559,In_841);
or U523 (N_523,In_854,In_155);
nand U524 (N_524,In_738,N_433);
xor U525 (N_525,In_529,N_190);
xor U526 (N_526,N_419,In_366);
nand U527 (N_527,In_379,In_146);
nand U528 (N_528,In_361,In_601);
xor U529 (N_529,N_448,N_319);
nand U530 (N_530,N_482,In_452);
xor U531 (N_531,N_272,N_275);
and U532 (N_532,N_186,N_180);
nor U533 (N_533,N_78,N_329);
and U534 (N_534,N_494,N_242);
and U535 (N_535,N_55,N_271);
and U536 (N_536,N_437,N_464);
xnor U537 (N_537,In_752,N_442);
or U538 (N_538,In_27,N_360);
and U539 (N_539,N_403,N_323);
or U540 (N_540,N_483,N_395);
or U541 (N_541,In_310,N_478);
nor U542 (N_542,In_290,N_273);
or U543 (N_543,N_473,N_428);
nor U544 (N_544,N_479,N_460);
nor U545 (N_545,N_491,In_103);
xor U546 (N_546,N_471,In_138);
or U547 (N_547,In_827,In_199);
or U548 (N_548,In_610,In_582);
nor U549 (N_549,In_539,In_367);
or U550 (N_550,N_393,N_214);
and U551 (N_551,In_222,In_590);
or U552 (N_552,N_96,N_382);
nor U553 (N_553,N_427,N_230);
xnor U554 (N_554,N_15,N_415);
nand U555 (N_555,In_498,In_397);
or U556 (N_556,N_452,N_369);
or U557 (N_557,N_402,N_470);
xor U558 (N_558,In_826,N_438);
nor U559 (N_559,In_112,N_233);
or U560 (N_560,In_184,N_496);
or U561 (N_561,In_850,In_265);
nor U562 (N_562,N_352,In_19);
nor U563 (N_563,In_148,N_240);
xnor U564 (N_564,N_463,In_942);
xnor U565 (N_565,N_481,In_998);
and U566 (N_566,N_412,In_387);
xor U567 (N_567,In_702,N_455);
nand U568 (N_568,In_984,N_446);
or U569 (N_569,In_695,N_7);
nand U570 (N_570,N_465,In_707);
or U571 (N_571,N_431,In_960);
nand U572 (N_572,In_326,In_563);
or U573 (N_573,N_436,N_414);
nand U574 (N_574,N_95,In_774);
and U575 (N_575,N_267,In_729);
or U576 (N_576,N_466,In_385);
and U577 (N_577,N_161,N_445);
and U578 (N_578,N_359,N_358);
and U579 (N_579,N_225,In_865);
or U580 (N_580,In_131,In_513);
or U581 (N_581,N_340,N_396);
nand U582 (N_582,In_97,N_450);
nand U583 (N_583,N_317,N_185);
nor U584 (N_584,In_351,N_371);
nor U585 (N_585,N_324,In_565);
nor U586 (N_586,N_365,In_878);
nand U587 (N_587,In_535,In_688);
nand U588 (N_588,N_434,N_56);
nor U589 (N_589,N_202,In_895);
nand U590 (N_590,In_156,In_940);
xnor U591 (N_591,N_59,In_263);
nand U592 (N_592,N_426,In_240);
xor U593 (N_593,N_354,In_218);
or U594 (N_594,In_545,In_569);
xnor U595 (N_595,N_135,In_34);
and U596 (N_596,N_211,In_115);
nand U597 (N_597,N_350,N_447);
or U598 (N_598,In_727,N_348);
nand U599 (N_599,In_846,In_370);
or U600 (N_600,N_550,N_52);
nand U601 (N_601,N_499,N_343);
and U602 (N_602,In_549,In_548);
xor U603 (N_603,In_430,In_54);
or U604 (N_604,N_221,N_335);
nor U605 (N_605,In_123,N_333);
or U606 (N_606,N_289,N_592);
nor U607 (N_607,N_332,In_743);
xnor U608 (N_608,In_434,N_416);
or U609 (N_609,In_953,N_537);
and U610 (N_610,N_118,N_574);
nor U611 (N_611,N_288,N_206);
nand U612 (N_612,N_310,N_410);
nor U613 (N_613,In_196,In_451);
nor U614 (N_614,N_312,In_477);
xor U615 (N_615,N_370,N_539);
xnor U616 (N_616,N_508,N_476);
nor U617 (N_617,N_535,N_216);
nand U618 (N_618,N_548,N_154);
nand U619 (N_619,N_580,In_235);
or U620 (N_620,N_505,In_499);
nand U621 (N_621,N_163,N_581);
or U622 (N_622,N_361,N_119);
and U623 (N_623,In_927,In_830);
xnor U624 (N_624,In_409,N_411);
nor U625 (N_625,In_140,In_116);
and U626 (N_626,N_265,In_536);
xor U627 (N_627,N_199,N_525);
nand U628 (N_628,In_229,N_589);
or U629 (N_629,In_594,N_562);
xnor U630 (N_630,N_502,N_391);
or U631 (N_631,N_457,N_495);
or U632 (N_632,In_572,In_912);
or U633 (N_633,N_301,N_486);
nor U634 (N_634,In_393,In_121);
or U635 (N_635,In_154,In_831);
nor U636 (N_636,In_918,N_528);
and U637 (N_637,In_356,In_900);
or U638 (N_638,N_569,N_217);
nor U639 (N_639,In_626,N_274);
nor U640 (N_640,N_339,N_126);
nand U641 (N_641,N_147,N_227);
nor U642 (N_642,N_385,N_53);
nor U643 (N_643,In_424,N_492);
nand U644 (N_644,N_555,In_7);
xor U645 (N_645,N_568,N_493);
and U646 (N_646,N_408,In_635);
or U647 (N_647,N_346,N_527);
xor U648 (N_648,N_585,N_390);
xor U649 (N_649,N_533,N_597);
xor U650 (N_650,N_45,N_547);
and U651 (N_651,In_169,N_511);
xor U652 (N_652,N_467,N_552);
and U653 (N_653,N_298,In_839);
or U654 (N_654,N_524,N_125);
nand U655 (N_655,In_491,N_472);
xnor U656 (N_656,In_633,N_584);
or U657 (N_657,In_996,N_378);
nand U658 (N_658,In_418,N_208);
and U659 (N_659,N_530,In_325);
nand U660 (N_660,N_61,N_262);
or U661 (N_661,N_549,In_679);
nor U662 (N_662,N_563,In_383);
xor U663 (N_663,In_5,In_398);
xor U664 (N_664,N_458,N_595);
nor U665 (N_665,In_676,In_29);
nand U666 (N_666,In_401,In_58);
nand U667 (N_667,In_818,In_78);
and U668 (N_668,N_543,In_101);
and U669 (N_669,In_906,In_39);
nor U670 (N_670,N_362,In_369);
and U671 (N_671,N_328,N_546);
nand U672 (N_672,N_43,N_299);
or U673 (N_673,N_132,N_575);
xor U674 (N_674,N_468,N_338);
or U675 (N_675,In_602,N_497);
xnor U676 (N_676,N_196,N_507);
or U677 (N_677,N_440,N_34);
and U678 (N_678,In_185,In_287);
and U679 (N_679,In_400,N_554);
nand U680 (N_680,In_880,N_331);
nor U681 (N_681,N_435,N_529);
xnor U682 (N_682,N_490,N_430);
and U683 (N_683,N_594,N_316);
xnor U684 (N_684,N_380,N_498);
xnor U685 (N_685,N_588,In_697);
nand U686 (N_686,N_421,In_725);
and U687 (N_687,N_16,In_899);
and U688 (N_688,In_977,N_30);
xnor U689 (N_689,N_308,N_513);
xnor U690 (N_690,N_500,N_542);
nor U691 (N_691,N_134,N_409);
and U692 (N_692,N_586,N_236);
nor U693 (N_693,N_520,In_3);
nand U694 (N_694,N_404,In_550);
nand U695 (N_695,N_276,In_390);
or U696 (N_696,N_510,N_477);
nand U697 (N_697,In_328,In_359);
xnor U698 (N_698,N_325,In_474);
nor U699 (N_699,N_536,N_534);
and U700 (N_700,N_598,N_696);
nor U701 (N_701,N_577,N_422);
or U702 (N_702,N_521,N_131);
nor U703 (N_703,In_595,N_630);
nor U704 (N_704,N_590,N_656);
xnor U705 (N_705,N_652,N_695);
or U706 (N_706,N_560,In_167);
or U707 (N_707,In_332,N_670);
nand U708 (N_708,N_545,N_77);
nand U709 (N_709,N_444,In_432);
xor U710 (N_710,N_375,N_480);
nand U711 (N_711,In_137,N_558);
or U712 (N_712,In_282,N_650);
xnor U713 (N_713,N_429,N_637);
nor U714 (N_714,N_678,N_451);
xnor U715 (N_715,N_618,N_643);
or U716 (N_716,N_337,N_673);
or U717 (N_717,N_635,N_189);
xor U718 (N_718,N_646,N_459);
xnor U719 (N_719,In_380,N_613);
and U720 (N_720,In_180,N_376);
nor U721 (N_721,In_759,N_578);
nand U722 (N_722,In_719,In_410);
or U723 (N_723,N_503,N_565);
or U724 (N_724,N_406,N_516);
nand U725 (N_725,N_698,N_677);
and U726 (N_726,N_614,In_787);
nor U727 (N_727,N_506,N_641);
nor U728 (N_728,In_687,In_892);
nand U729 (N_729,N_443,N_349);
nand U730 (N_730,N_76,In_478);
or U731 (N_731,N_615,N_694);
nor U732 (N_732,N_9,N_666);
nand U733 (N_733,N_601,N_439);
xor U734 (N_734,In_825,N_423);
nor U735 (N_735,N_512,In_611);
and U736 (N_736,N_400,N_605);
xor U737 (N_737,N_300,N_644);
nand U738 (N_738,N_504,In_197);
or U739 (N_739,N_515,In_92);
xor U740 (N_740,In_873,N_675);
nand U741 (N_741,N_285,N_681);
or U742 (N_742,N_693,In_646);
nor U743 (N_743,N_642,N_347);
and U744 (N_744,N_604,In_917);
xnor U745 (N_745,N_654,N_432);
nor U746 (N_746,N_551,N_260);
xnor U747 (N_747,N_669,In_780);
nor U748 (N_748,In_427,N_39);
and U749 (N_749,N_424,N_626);
nor U750 (N_750,In_712,In_110);
and U751 (N_751,N_572,In_837);
or U752 (N_752,N_616,N_663);
xnor U753 (N_753,N_541,N_685);
and U754 (N_754,N_699,In_448);
nor U755 (N_755,N_561,N_628);
or U756 (N_756,In_840,N_342);
xor U757 (N_757,In_161,N_27);
nand U758 (N_758,N_405,In_696);
nand U759 (N_759,N_593,In_174);
nor U760 (N_760,N_268,N_672);
or U761 (N_761,N_631,N_57);
nand U762 (N_762,N_638,N_296);
nand U763 (N_763,N_579,N_688);
nand U764 (N_764,N_676,N_633);
and U765 (N_765,N_453,In_117);
or U766 (N_766,N_519,N_557);
nor U767 (N_767,N_509,N_401);
nor U768 (N_768,In_681,N_573);
nor U769 (N_769,In_793,N_127);
and U770 (N_770,N_334,N_587);
xor U771 (N_771,N_610,N_113);
nor U772 (N_772,N_600,N_647);
and U773 (N_773,N_624,N_576);
nor U774 (N_774,In_302,N_692);
and U775 (N_775,N_485,N_112);
xor U776 (N_776,In_431,N_399);
or U777 (N_777,In_861,N_668);
nand U778 (N_778,N_556,In_661);
or U779 (N_779,N_151,N_566);
nor U780 (N_780,N_648,N_531);
xnor U781 (N_781,In_378,N_475);
and U782 (N_782,N_522,N_691);
and U783 (N_783,N_680,N_609);
or U784 (N_784,N_658,N_526);
xor U785 (N_785,N_311,N_474);
nand U786 (N_786,In_331,N_664);
and U787 (N_787,In_442,N_651);
or U788 (N_788,N_632,N_689);
or U789 (N_789,N_462,N_501);
and U790 (N_790,N_617,N_418);
nand U791 (N_791,N_321,N_454);
or U792 (N_792,N_155,In_145);
nor U793 (N_793,N_636,N_640);
xor U794 (N_794,N_559,N_517);
or U795 (N_795,N_129,N_336);
and U796 (N_796,N_413,N_661);
and U797 (N_797,N_690,N_564);
xnor U798 (N_798,In_127,N_625);
nand U799 (N_799,N_621,N_538);
or U800 (N_800,In_346,In_538);
and U801 (N_801,N_659,N_784);
xnor U802 (N_802,N_719,N_752);
xor U803 (N_803,N_772,N_777);
or U804 (N_804,N_716,N_744);
nand U805 (N_805,N_544,N_758);
xnor U806 (N_806,N_781,In_278);
xnor U807 (N_807,N_710,N_709);
or U808 (N_808,N_364,N_748);
or U809 (N_809,N_210,N_697);
nor U810 (N_810,N_757,N_523);
nand U811 (N_811,N_790,N_570);
and U812 (N_812,In_791,N_794);
nand U813 (N_813,N_775,N_707);
xnor U814 (N_814,N_571,N_674);
or U815 (N_815,N_718,N_623);
xnor U816 (N_816,In_322,N_761);
or U817 (N_817,N_785,N_553);
or U818 (N_818,N_687,N_231);
nor U819 (N_819,N_17,N_567);
nor U820 (N_820,N_671,N_701);
nand U821 (N_821,N_756,N_736);
and U822 (N_822,N_665,N_759);
nor U823 (N_823,N_142,N_26);
nor U824 (N_824,N_662,N_684);
nor U825 (N_825,N_729,N_764);
nor U826 (N_826,N_191,N_80);
xor U827 (N_827,In_963,N_645);
xor U828 (N_828,N_796,N_795);
or U829 (N_829,N_721,N_747);
xnor U830 (N_830,N_789,N_760);
nand U831 (N_831,N_750,N_763);
or U832 (N_832,N_731,N_783);
xnor U833 (N_833,N_682,In_164);
or U834 (N_834,In_308,N_720);
or U835 (N_835,N_611,In_163);
nand U836 (N_836,In_994,N_793);
or U837 (N_837,N_683,N_489);
and U838 (N_838,N_653,N_733);
nand U839 (N_839,N_741,N_778);
xor U840 (N_840,N_742,N_603);
or U841 (N_841,In_339,N_713);
nor U842 (N_842,N_765,N_243);
xor U843 (N_843,N_769,N_591);
nand U844 (N_844,N_606,N_780);
nand U845 (N_845,N_639,N_353);
and U846 (N_846,N_737,N_218);
nor U847 (N_847,N_739,N_187);
or U848 (N_848,N_657,N_622);
nor U849 (N_849,N_368,N_774);
and U850 (N_850,N_732,N_755);
nand U851 (N_851,In_126,N_398);
and U852 (N_852,N_766,In_742);
nor U853 (N_853,N_608,N_667);
nand U854 (N_854,N_704,N_762);
nor U855 (N_855,N_700,In_104);
and U856 (N_856,N_734,N_469);
nor U857 (N_857,N_717,N_771);
xor U858 (N_858,N_168,N_725);
nor U859 (N_859,In_734,N_773);
and U860 (N_860,N_735,N_583);
xnor U861 (N_861,N_749,N_220);
nor U862 (N_862,N_425,N_596);
xor U863 (N_863,N_679,N_703);
xor U864 (N_864,N_787,N_798);
nand U865 (N_865,N_441,In_108);
and U866 (N_866,N_215,N_702);
nand U867 (N_867,In_609,N_282);
nor U868 (N_868,N_612,N_620);
or U869 (N_869,N_532,N_791);
xor U870 (N_870,N_779,N_540);
or U871 (N_871,In_65,N_629);
and U872 (N_872,N_753,N_782);
nor U873 (N_873,N_792,N_599);
nor U874 (N_874,N_518,N_799);
nor U875 (N_875,N_100,N_634);
nor U876 (N_876,In_872,N_582);
nand U877 (N_877,In_809,N_797);
nor U878 (N_878,N_708,N_723);
xor U879 (N_879,N_743,N_146);
nand U880 (N_880,N_724,N_786);
nor U881 (N_881,N_627,N_751);
xnor U882 (N_882,N_715,N_770);
nor U883 (N_883,N_738,N_602);
xor U884 (N_884,N_619,N_649);
and U885 (N_885,In_910,N_722);
or U886 (N_886,N_309,N_727);
or U887 (N_887,N_754,N_660);
and U888 (N_888,N_712,N_776);
or U889 (N_889,N_487,N_730);
nor U890 (N_890,N_607,N_686);
nor U891 (N_891,N_714,N_655);
or U892 (N_892,N_514,N_279);
and U893 (N_893,N_768,N_746);
xnor U894 (N_894,N_767,N_740);
and U895 (N_895,N_20,N_726);
or U896 (N_896,In_739,N_745);
nand U897 (N_897,N_711,N_788);
nand U898 (N_898,N_705,N_728);
nand U899 (N_899,N_706,In_449);
or U900 (N_900,N_898,N_839);
xnor U901 (N_901,N_804,N_824);
nor U902 (N_902,N_849,N_864);
or U903 (N_903,N_831,N_886);
or U904 (N_904,N_883,N_877);
or U905 (N_905,N_829,N_825);
and U906 (N_906,N_867,N_842);
or U907 (N_907,N_894,N_876);
nand U908 (N_908,N_869,N_833);
or U909 (N_909,N_859,N_828);
xor U910 (N_910,N_805,N_812);
or U911 (N_911,N_850,N_857);
xor U912 (N_912,N_899,N_816);
nand U913 (N_913,N_818,N_878);
xor U914 (N_914,N_868,N_826);
and U915 (N_915,N_801,N_808);
or U916 (N_916,N_838,N_881);
and U917 (N_917,N_858,N_897);
and U918 (N_918,N_809,N_884);
xnor U919 (N_919,N_840,N_862);
and U920 (N_920,N_880,N_830);
nand U921 (N_921,N_888,N_810);
and U922 (N_922,N_852,N_861);
nor U923 (N_923,N_855,N_827);
or U924 (N_924,N_800,N_832);
xor U925 (N_925,N_819,N_851);
and U926 (N_926,N_854,N_892);
xor U927 (N_927,N_802,N_807);
xor U928 (N_928,N_896,N_845);
and U929 (N_929,N_860,N_835);
nor U930 (N_930,N_814,N_873);
and U931 (N_931,N_821,N_823);
nor U932 (N_932,N_813,N_872);
and U933 (N_933,N_817,N_846);
nand U934 (N_934,N_887,N_856);
or U935 (N_935,N_866,N_891);
xor U936 (N_936,N_811,N_853);
nand U937 (N_937,N_847,N_885);
nor U938 (N_938,N_890,N_815);
and U939 (N_939,N_865,N_870);
nor U940 (N_940,N_844,N_837);
xnor U941 (N_941,N_895,N_834);
nand U942 (N_942,N_875,N_889);
and U943 (N_943,N_843,N_803);
and U944 (N_944,N_871,N_863);
xor U945 (N_945,N_822,N_874);
nor U946 (N_946,N_836,N_841);
and U947 (N_947,N_893,N_820);
nand U948 (N_948,N_882,N_848);
or U949 (N_949,N_879,N_806);
and U950 (N_950,N_871,N_862);
xnor U951 (N_951,N_883,N_889);
or U952 (N_952,N_874,N_884);
xor U953 (N_953,N_852,N_827);
xnor U954 (N_954,N_864,N_863);
nand U955 (N_955,N_816,N_800);
nand U956 (N_956,N_894,N_829);
and U957 (N_957,N_842,N_847);
nor U958 (N_958,N_854,N_818);
xnor U959 (N_959,N_848,N_854);
or U960 (N_960,N_894,N_859);
nor U961 (N_961,N_801,N_848);
nor U962 (N_962,N_844,N_832);
xor U963 (N_963,N_846,N_830);
or U964 (N_964,N_862,N_819);
nand U965 (N_965,N_884,N_896);
or U966 (N_966,N_866,N_804);
and U967 (N_967,N_893,N_804);
or U968 (N_968,N_805,N_814);
or U969 (N_969,N_898,N_899);
nand U970 (N_970,N_829,N_853);
nand U971 (N_971,N_862,N_808);
and U972 (N_972,N_870,N_809);
xnor U973 (N_973,N_879,N_876);
nand U974 (N_974,N_840,N_891);
nand U975 (N_975,N_851,N_877);
xor U976 (N_976,N_809,N_895);
xnor U977 (N_977,N_892,N_891);
and U978 (N_978,N_892,N_895);
nand U979 (N_979,N_834,N_872);
and U980 (N_980,N_873,N_836);
and U981 (N_981,N_891,N_851);
nand U982 (N_982,N_848,N_857);
nand U983 (N_983,N_873,N_835);
and U984 (N_984,N_837,N_803);
nor U985 (N_985,N_800,N_856);
and U986 (N_986,N_834,N_838);
or U987 (N_987,N_853,N_869);
or U988 (N_988,N_865,N_853);
nor U989 (N_989,N_836,N_827);
nor U990 (N_990,N_890,N_876);
xor U991 (N_991,N_874,N_846);
and U992 (N_992,N_809,N_883);
nand U993 (N_993,N_897,N_873);
nand U994 (N_994,N_881,N_855);
xnor U995 (N_995,N_846,N_893);
and U996 (N_996,N_834,N_871);
xnor U997 (N_997,N_884,N_850);
and U998 (N_998,N_847,N_861);
xor U999 (N_999,N_866,N_820);
or U1000 (N_1000,N_915,N_955);
and U1001 (N_1001,N_921,N_961);
or U1002 (N_1002,N_950,N_986);
xor U1003 (N_1003,N_999,N_907);
nor U1004 (N_1004,N_933,N_948);
and U1005 (N_1005,N_916,N_980);
nor U1006 (N_1006,N_942,N_944);
or U1007 (N_1007,N_919,N_956);
xor U1008 (N_1008,N_993,N_923);
and U1009 (N_1009,N_900,N_924);
and U1010 (N_1010,N_953,N_901);
or U1011 (N_1011,N_977,N_949);
and U1012 (N_1012,N_975,N_913);
nand U1013 (N_1013,N_922,N_947);
nand U1014 (N_1014,N_914,N_940);
and U1015 (N_1015,N_990,N_946);
nand U1016 (N_1016,N_958,N_938);
xnor U1017 (N_1017,N_943,N_952);
and U1018 (N_1018,N_903,N_971);
xnor U1019 (N_1019,N_982,N_935);
xor U1020 (N_1020,N_926,N_967);
and U1021 (N_1021,N_931,N_910);
nand U1022 (N_1022,N_970,N_928);
and U1023 (N_1023,N_945,N_951);
nand U1024 (N_1024,N_965,N_902);
nor U1025 (N_1025,N_941,N_963);
nand U1026 (N_1026,N_912,N_960);
xor U1027 (N_1027,N_905,N_911);
xor U1028 (N_1028,N_964,N_934);
nor U1029 (N_1029,N_962,N_997);
nand U1030 (N_1030,N_937,N_908);
xor U1031 (N_1031,N_917,N_983);
and U1032 (N_1032,N_918,N_976);
and U1033 (N_1033,N_906,N_996);
and U1034 (N_1034,N_909,N_991);
nand U1035 (N_1035,N_979,N_936);
nor U1036 (N_1036,N_957,N_930);
and U1037 (N_1037,N_987,N_981);
nand U1038 (N_1038,N_998,N_954);
and U1039 (N_1039,N_939,N_989);
xnor U1040 (N_1040,N_978,N_969);
nand U1041 (N_1041,N_966,N_972);
or U1042 (N_1042,N_992,N_932);
and U1043 (N_1043,N_995,N_920);
xor U1044 (N_1044,N_973,N_985);
xnor U1045 (N_1045,N_925,N_904);
nor U1046 (N_1046,N_968,N_929);
xor U1047 (N_1047,N_974,N_984);
or U1048 (N_1048,N_959,N_988);
and U1049 (N_1049,N_994,N_927);
nor U1050 (N_1050,N_906,N_952);
nand U1051 (N_1051,N_937,N_955);
nor U1052 (N_1052,N_945,N_908);
or U1053 (N_1053,N_944,N_905);
or U1054 (N_1054,N_904,N_915);
xor U1055 (N_1055,N_940,N_979);
xor U1056 (N_1056,N_930,N_945);
nand U1057 (N_1057,N_939,N_953);
and U1058 (N_1058,N_965,N_912);
nand U1059 (N_1059,N_916,N_932);
nand U1060 (N_1060,N_910,N_921);
or U1061 (N_1061,N_953,N_995);
or U1062 (N_1062,N_987,N_970);
nand U1063 (N_1063,N_935,N_978);
and U1064 (N_1064,N_922,N_923);
xor U1065 (N_1065,N_930,N_935);
xor U1066 (N_1066,N_954,N_942);
nor U1067 (N_1067,N_969,N_992);
or U1068 (N_1068,N_944,N_962);
or U1069 (N_1069,N_928,N_986);
nor U1070 (N_1070,N_959,N_956);
nand U1071 (N_1071,N_938,N_988);
and U1072 (N_1072,N_971,N_935);
xor U1073 (N_1073,N_961,N_986);
and U1074 (N_1074,N_946,N_972);
nor U1075 (N_1075,N_969,N_956);
and U1076 (N_1076,N_981,N_950);
nand U1077 (N_1077,N_938,N_996);
nand U1078 (N_1078,N_911,N_976);
nor U1079 (N_1079,N_905,N_968);
nor U1080 (N_1080,N_908,N_955);
and U1081 (N_1081,N_962,N_994);
and U1082 (N_1082,N_949,N_974);
or U1083 (N_1083,N_971,N_970);
nor U1084 (N_1084,N_974,N_982);
or U1085 (N_1085,N_944,N_981);
and U1086 (N_1086,N_969,N_908);
nor U1087 (N_1087,N_965,N_953);
xnor U1088 (N_1088,N_954,N_930);
or U1089 (N_1089,N_904,N_972);
xor U1090 (N_1090,N_937,N_945);
and U1091 (N_1091,N_980,N_903);
xor U1092 (N_1092,N_925,N_919);
xor U1093 (N_1093,N_985,N_941);
xnor U1094 (N_1094,N_970,N_950);
xnor U1095 (N_1095,N_968,N_981);
nor U1096 (N_1096,N_930,N_953);
xor U1097 (N_1097,N_992,N_961);
nand U1098 (N_1098,N_910,N_915);
and U1099 (N_1099,N_935,N_912);
xor U1100 (N_1100,N_1047,N_1070);
and U1101 (N_1101,N_1049,N_1010);
xnor U1102 (N_1102,N_1090,N_1096);
or U1103 (N_1103,N_1018,N_1005);
nand U1104 (N_1104,N_1022,N_1050);
nand U1105 (N_1105,N_1060,N_1033);
and U1106 (N_1106,N_1081,N_1048);
nand U1107 (N_1107,N_1043,N_1072);
and U1108 (N_1108,N_1020,N_1099);
nand U1109 (N_1109,N_1055,N_1093);
nand U1110 (N_1110,N_1074,N_1059);
xnor U1111 (N_1111,N_1071,N_1003);
and U1112 (N_1112,N_1030,N_1016);
and U1113 (N_1113,N_1008,N_1052);
or U1114 (N_1114,N_1075,N_1067);
or U1115 (N_1115,N_1061,N_1086);
nor U1116 (N_1116,N_1080,N_1021);
xnor U1117 (N_1117,N_1078,N_1007);
and U1118 (N_1118,N_1087,N_1040);
nand U1119 (N_1119,N_1000,N_1051);
and U1120 (N_1120,N_1042,N_1084);
nand U1121 (N_1121,N_1094,N_1097);
xor U1122 (N_1122,N_1006,N_1066);
xnor U1123 (N_1123,N_1058,N_1057);
xnor U1124 (N_1124,N_1009,N_1012);
nand U1125 (N_1125,N_1069,N_1019);
nand U1126 (N_1126,N_1038,N_1098);
or U1127 (N_1127,N_1046,N_1011);
xor U1128 (N_1128,N_1054,N_1013);
and U1129 (N_1129,N_1082,N_1091);
or U1130 (N_1130,N_1024,N_1029);
nor U1131 (N_1131,N_1077,N_1026);
and U1132 (N_1132,N_1031,N_1092);
nand U1133 (N_1133,N_1079,N_1076);
xnor U1134 (N_1134,N_1056,N_1045);
xor U1135 (N_1135,N_1068,N_1089);
nor U1136 (N_1136,N_1032,N_1083);
and U1137 (N_1137,N_1044,N_1036);
xor U1138 (N_1138,N_1063,N_1035);
xnor U1139 (N_1139,N_1088,N_1085);
nor U1140 (N_1140,N_1014,N_1065);
or U1141 (N_1141,N_1017,N_1062);
nor U1142 (N_1142,N_1001,N_1002);
nand U1143 (N_1143,N_1095,N_1004);
xnor U1144 (N_1144,N_1028,N_1034);
nor U1145 (N_1145,N_1053,N_1025);
and U1146 (N_1146,N_1023,N_1027);
xnor U1147 (N_1147,N_1073,N_1064);
nand U1148 (N_1148,N_1041,N_1015);
nand U1149 (N_1149,N_1037,N_1039);
nand U1150 (N_1150,N_1082,N_1008);
and U1151 (N_1151,N_1005,N_1072);
and U1152 (N_1152,N_1001,N_1075);
and U1153 (N_1153,N_1029,N_1018);
nor U1154 (N_1154,N_1061,N_1050);
nand U1155 (N_1155,N_1018,N_1042);
or U1156 (N_1156,N_1000,N_1064);
xor U1157 (N_1157,N_1044,N_1016);
xnor U1158 (N_1158,N_1019,N_1061);
and U1159 (N_1159,N_1045,N_1097);
nor U1160 (N_1160,N_1040,N_1034);
xnor U1161 (N_1161,N_1070,N_1095);
nor U1162 (N_1162,N_1091,N_1042);
or U1163 (N_1163,N_1047,N_1026);
or U1164 (N_1164,N_1018,N_1065);
nor U1165 (N_1165,N_1095,N_1055);
nand U1166 (N_1166,N_1077,N_1015);
and U1167 (N_1167,N_1078,N_1069);
and U1168 (N_1168,N_1097,N_1023);
nor U1169 (N_1169,N_1082,N_1030);
nand U1170 (N_1170,N_1050,N_1031);
or U1171 (N_1171,N_1023,N_1040);
xor U1172 (N_1172,N_1064,N_1043);
xnor U1173 (N_1173,N_1063,N_1057);
or U1174 (N_1174,N_1065,N_1048);
xnor U1175 (N_1175,N_1052,N_1026);
or U1176 (N_1176,N_1042,N_1004);
and U1177 (N_1177,N_1070,N_1043);
nor U1178 (N_1178,N_1066,N_1034);
or U1179 (N_1179,N_1011,N_1096);
nand U1180 (N_1180,N_1071,N_1091);
and U1181 (N_1181,N_1002,N_1009);
and U1182 (N_1182,N_1010,N_1012);
xnor U1183 (N_1183,N_1023,N_1073);
xnor U1184 (N_1184,N_1034,N_1093);
nand U1185 (N_1185,N_1044,N_1055);
or U1186 (N_1186,N_1078,N_1076);
nand U1187 (N_1187,N_1024,N_1022);
or U1188 (N_1188,N_1097,N_1028);
or U1189 (N_1189,N_1038,N_1000);
or U1190 (N_1190,N_1054,N_1001);
nor U1191 (N_1191,N_1000,N_1040);
nor U1192 (N_1192,N_1075,N_1087);
or U1193 (N_1193,N_1072,N_1027);
and U1194 (N_1194,N_1022,N_1014);
xnor U1195 (N_1195,N_1057,N_1056);
nor U1196 (N_1196,N_1006,N_1005);
or U1197 (N_1197,N_1075,N_1083);
and U1198 (N_1198,N_1018,N_1052);
or U1199 (N_1199,N_1017,N_1039);
or U1200 (N_1200,N_1166,N_1188);
nand U1201 (N_1201,N_1139,N_1113);
nand U1202 (N_1202,N_1187,N_1158);
xnor U1203 (N_1203,N_1138,N_1198);
nor U1204 (N_1204,N_1143,N_1102);
xnor U1205 (N_1205,N_1167,N_1150);
or U1206 (N_1206,N_1119,N_1127);
xnor U1207 (N_1207,N_1152,N_1115);
or U1208 (N_1208,N_1109,N_1145);
or U1209 (N_1209,N_1177,N_1103);
and U1210 (N_1210,N_1137,N_1156);
and U1211 (N_1211,N_1122,N_1140);
nor U1212 (N_1212,N_1142,N_1165);
nand U1213 (N_1213,N_1141,N_1106);
or U1214 (N_1214,N_1136,N_1163);
and U1215 (N_1215,N_1154,N_1120);
and U1216 (N_1216,N_1101,N_1172);
or U1217 (N_1217,N_1147,N_1124);
nand U1218 (N_1218,N_1125,N_1105);
or U1219 (N_1219,N_1182,N_1161);
xor U1220 (N_1220,N_1118,N_1195);
xor U1221 (N_1221,N_1174,N_1117);
nor U1222 (N_1222,N_1170,N_1185);
or U1223 (N_1223,N_1173,N_1151);
or U1224 (N_1224,N_1107,N_1199);
nor U1225 (N_1225,N_1155,N_1162);
or U1226 (N_1226,N_1111,N_1160);
or U1227 (N_1227,N_1178,N_1169);
and U1228 (N_1228,N_1153,N_1130);
and U1229 (N_1229,N_1128,N_1104);
or U1230 (N_1230,N_1126,N_1186);
or U1231 (N_1231,N_1175,N_1123);
or U1232 (N_1232,N_1181,N_1164);
and U1233 (N_1233,N_1132,N_1191);
or U1234 (N_1234,N_1179,N_1189);
and U1235 (N_1235,N_1197,N_1100);
and U1236 (N_1236,N_1148,N_1133);
xnor U1237 (N_1237,N_1171,N_1146);
or U1238 (N_1238,N_1194,N_1149);
nor U1239 (N_1239,N_1129,N_1131);
and U1240 (N_1240,N_1144,N_1112);
and U1241 (N_1241,N_1157,N_1159);
xor U1242 (N_1242,N_1168,N_1121);
and U1243 (N_1243,N_1135,N_1183);
nor U1244 (N_1244,N_1114,N_1192);
nor U1245 (N_1245,N_1110,N_1184);
nor U1246 (N_1246,N_1193,N_1180);
or U1247 (N_1247,N_1116,N_1196);
xor U1248 (N_1248,N_1108,N_1190);
and U1249 (N_1249,N_1134,N_1176);
nor U1250 (N_1250,N_1162,N_1193);
nor U1251 (N_1251,N_1134,N_1105);
nor U1252 (N_1252,N_1168,N_1164);
xnor U1253 (N_1253,N_1158,N_1195);
nor U1254 (N_1254,N_1151,N_1128);
and U1255 (N_1255,N_1119,N_1132);
or U1256 (N_1256,N_1196,N_1120);
or U1257 (N_1257,N_1140,N_1133);
or U1258 (N_1258,N_1151,N_1143);
or U1259 (N_1259,N_1143,N_1167);
nor U1260 (N_1260,N_1169,N_1158);
xor U1261 (N_1261,N_1188,N_1191);
and U1262 (N_1262,N_1102,N_1119);
or U1263 (N_1263,N_1194,N_1117);
nor U1264 (N_1264,N_1150,N_1126);
xnor U1265 (N_1265,N_1119,N_1164);
and U1266 (N_1266,N_1119,N_1175);
nor U1267 (N_1267,N_1184,N_1158);
or U1268 (N_1268,N_1139,N_1105);
or U1269 (N_1269,N_1138,N_1102);
or U1270 (N_1270,N_1105,N_1107);
nor U1271 (N_1271,N_1154,N_1104);
nor U1272 (N_1272,N_1147,N_1152);
and U1273 (N_1273,N_1129,N_1188);
xor U1274 (N_1274,N_1199,N_1148);
xor U1275 (N_1275,N_1186,N_1181);
and U1276 (N_1276,N_1127,N_1125);
and U1277 (N_1277,N_1168,N_1196);
xnor U1278 (N_1278,N_1145,N_1181);
nand U1279 (N_1279,N_1166,N_1118);
nand U1280 (N_1280,N_1157,N_1188);
nor U1281 (N_1281,N_1184,N_1180);
nor U1282 (N_1282,N_1115,N_1124);
xor U1283 (N_1283,N_1119,N_1195);
or U1284 (N_1284,N_1100,N_1124);
xnor U1285 (N_1285,N_1104,N_1196);
nand U1286 (N_1286,N_1161,N_1140);
or U1287 (N_1287,N_1130,N_1113);
xor U1288 (N_1288,N_1184,N_1105);
and U1289 (N_1289,N_1157,N_1186);
or U1290 (N_1290,N_1143,N_1168);
and U1291 (N_1291,N_1174,N_1118);
nor U1292 (N_1292,N_1108,N_1129);
nor U1293 (N_1293,N_1117,N_1149);
or U1294 (N_1294,N_1146,N_1129);
nor U1295 (N_1295,N_1162,N_1117);
or U1296 (N_1296,N_1153,N_1174);
or U1297 (N_1297,N_1110,N_1132);
xor U1298 (N_1298,N_1121,N_1107);
and U1299 (N_1299,N_1164,N_1129);
or U1300 (N_1300,N_1246,N_1219);
or U1301 (N_1301,N_1298,N_1223);
or U1302 (N_1302,N_1277,N_1209);
nor U1303 (N_1303,N_1273,N_1210);
or U1304 (N_1304,N_1220,N_1214);
nor U1305 (N_1305,N_1260,N_1296);
or U1306 (N_1306,N_1287,N_1262);
nand U1307 (N_1307,N_1208,N_1221);
xor U1308 (N_1308,N_1241,N_1263);
nor U1309 (N_1309,N_1268,N_1247);
nor U1310 (N_1310,N_1264,N_1270);
and U1311 (N_1311,N_1293,N_1228);
nand U1312 (N_1312,N_1283,N_1266);
or U1313 (N_1313,N_1267,N_1279);
and U1314 (N_1314,N_1286,N_1227);
or U1315 (N_1315,N_1276,N_1233);
nand U1316 (N_1316,N_1239,N_1207);
xnor U1317 (N_1317,N_1235,N_1280);
and U1318 (N_1318,N_1200,N_1284);
xnor U1319 (N_1319,N_1218,N_1258);
nor U1320 (N_1320,N_1269,N_1244);
xnor U1321 (N_1321,N_1291,N_1259);
nand U1322 (N_1322,N_1242,N_1274);
nand U1323 (N_1323,N_1248,N_1216);
xor U1324 (N_1324,N_1224,N_1295);
nor U1325 (N_1325,N_1297,N_1272);
nor U1326 (N_1326,N_1250,N_1251);
nor U1327 (N_1327,N_1202,N_1236);
or U1328 (N_1328,N_1234,N_1294);
nand U1329 (N_1329,N_1255,N_1261);
nand U1330 (N_1330,N_1225,N_1222);
nand U1331 (N_1331,N_1217,N_1253);
xnor U1332 (N_1332,N_1201,N_1252);
and U1333 (N_1333,N_1240,N_1243);
xor U1334 (N_1334,N_1275,N_1212);
nor U1335 (N_1335,N_1257,N_1292);
and U1336 (N_1336,N_1271,N_1256);
and U1337 (N_1337,N_1278,N_1265);
and U1338 (N_1338,N_1232,N_1204);
or U1339 (N_1339,N_1281,N_1282);
xor U1340 (N_1340,N_1229,N_1203);
xnor U1341 (N_1341,N_1226,N_1289);
nand U1342 (N_1342,N_1206,N_1237);
and U1343 (N_1343,N_1290,N_1231);
nor U1344 (N_1344,N_1249,N_1285);
or U1345 (N_1345,N_1215,N_1254);
xnor U1346 (N_1346,N_1238,N_1230);
or U1347 (N_1347,N_1211,N_1245);
nand U1348 (N_1348,N_1213,N_1288);
nand U1349 (N_1349,N_1205,N_1299);
and U1350 (N_1350,N_1203,N_1219);
nor U1351 (N_1351,N_1292,N_1263);
and U1352 (N_1352,N_1259,N_1283);
xnor U1353 (N_1353,N_1255,N_1294);
xor U1354 (N_1354,N_1203,N_1239);
nand U1355 (N_1355,N_1238,N_1264);
and U1356 (N_1356,N_1285,N_1211);
xnor U1357 (N_1357,N_1266,N_1224);
xor U1358 (N_1358,N_1236,N_1261);
or U1359 (N_1359,N_1232,N_1225);
or U1360 (N_1360,N_1263,N_1278);
nor U1361 (N_1361,N_1295,N_1266);
nor U1362 (N_1362,N_1208,N_1283);
nand U1363 (N_1363,N_1263,N_1230);
nand U1364 (N_1364,N_1205,N_1296);
nor U1365 (N_1365,N_1213,N_1223);
and U1366 (N_1366,N_1211,N_1250);
nand U1367 (N_1367,N_1230,N_1212);
nand U1368 (N_1368,N_1218,N_1217);
xor U1369 (N_1369,N_1238,N_1299);
xnor U1370 (N_1370,N_1226,N_1286);
nor U1371 (N_1371,N_1229,N_1235);
and U1372 (N_1372,N_1212,N_1238);
nor U1373 (N_1373,N_1229,N_1280);
nand U1374 (N_1374,N_1223,N_1296);
and U1375 (N_1375,N_1222,N_1235);
nor U1376 (N_1376,N_1275,N_1297);
and U1377 (N_1377,N_1209,N_1291);
nor U1378 (N_1378,N_1227,N_1229);
or U1379 (N_1379,N_1240,N_1228);
or U1380 (N_1380,N_1225,N_1244);
xor U1381 (N_1381,N_1283,N_1250);
or U1382 (N_1382,N_1231,N_1263);
nor U1383 (N_1383,N_1245,N_1232);
and U1384 (N_1384,N_1237,N_1223);
nand U1385 (N_1385,N_1261,N_1253);
nand U1386 (N_1386,N_1276,N_1242);
nand U1387 (N_1387,N_1235,N_1259);
nor U1388 (N_1388,N_1221,N_1205);
nor U1389 (N_1389,N_1245,N_1291);
or U1390 (N_1390,N_1257,N_1298);
nor U1391 (N_1391,N_1225,N_1240);
or U1392 (N_1392,N_1274,N_1223);
nor U1393 (N_1393,N_1298,N_1274);
nand U1394 (N_1394,N_1293,N_1291);
nand U1395 (N_1395,N_1252,N_1270);
xor U1396 (N_1396,N_1262,N_1271);
or U1397 (N_1397,N_1219,N_1259);
or U1398 (N_1398,N_1244,N_1272);
nand U1399 (N_1399,N_1226,N_1266);
nand U1400 (N_1400,N_1380,N_1362);
xor U1401 (N_1401,N_1328,N_1393);
or U1402 (N_1402,N_1395,N_1320);
nand U1403 (N_1403,N_1340,N_1349);
xor U1404 (N_1404,N_1305,N_1306);
nor U1405 (N_1405,N_1344,N_1327);
xnor U1406 (N_1406,N_1371,N_1365);
xnor U1407 (N_1407,N_1398,N_1309);
and U1408 (N_1408,N_1396,N_1331);
or U1409 (N_1409,N_1308,N_1348);
or U1410 (N_1410,N_1324,N_1303);
or U1411 (N_1411,N_1312,N_1313);
nor U1412 (N_1412,N_1335,N_1321);
or U1413 (N_1413,N_1356,N_1334);
nand U1414 (N_1414,N_1399,N_1373);
xnor U1415 (N_1415,N_1341,N_1366);
and U1416 (N_1416,N_1379,N_1382);
xor U1417 (N_1417,N_1370,N_1311);
nor U1418 (N_1418,N_1372,N_1304);
nand U1419 (N_1419,N_1355,N_1326);
and U1420 (N_1420,N_1315,N_1351);
and U1421 (N_1421,N_1352,N_1364);
nor U1422 (N_1422,N_1363,N_1360);
and U1423 (N_1423,N_1394,N_1397);
and U1424 (N_1424,N_1385,N_1361);
or U1425 (N_1425,N_1376,N_1333);
nor U1426 (N_1426,N_1374,N_1325);
nor U1427 (N_1427,N_1323,N_1336);
nor U1428 (N_1428,N_1337,N_1387);
or U1429 (N_1429,N_1322,N_1353);
or U1430 (N_1430,N_1368,N_1330);
xnor U1431 (N_1431,N_1314,N_1300);
xor U1432 (N_1432,N_1358,N_1392);
nor U1433 (N_1433,N_1329,N_1318);
and U1434 (N_1434,N_1317,N_1350);
nand U1435 (N_1435,N_1338,N_1339);
nor U1436 (N_1436,N_1389,N_1342);
nor U1437 (N_1437,N_1369,N_1378);
nor U1438 (N_1438,N_1390,N_1377);
nand U1439 (N_1439,N_1354,N_1386);
xnor U1440 (N_1440,N_1332,N_1359);
and U1441 (N_1441,N_1391,N_1383);
xor U1442 (N_1442,N_1301,N_1346);
xnor U1443 (N_1443,N_1357,N_1307);
xnor U1444 (N_1444,N_1310,N_1375);
or U1445 (N_1445,N_1343,N_1319);
and U1446 (N_1446,N_1367,N_1316);
nand U1447 (N_1447,N_1388,N_1384);
or U1448 (N_1448,N_1302,N_1345);
nor U1449 (N_1449,N_1381,N_1347);
or U1450 (N_1450,N_1374,N_1330);
xnor U1451 (N_1451,N_1392,N_1321);
and U1452 (N_1452,N_1391,N_1349);
nand U1453 (N_1453,N_1344,N_1351);
and U1454 (N_1454,N_1357,N_1399);
nand U1455 (N_1455,N_1361,N_1335);
or U1456 (N_1456,N_1389,N_1333);
and U1457 (N_1457,N_1338,N_1391);
nand U1458 (N_1458,N_1311,N_1332);
and U1459 (N_1459,N_1326,N_1319);
or U1460 (N_1460,N_1393,N_1348);
or U1461 (N_1461,N_1377,N_1309);
nor U1462 (N_1462,N_1321,N_1391);
nand U1463 (N_1463,N_1392,N_1339);
xor U1464 (N_1464,N_1318,N_1300);
nand U1465 (N_1465,N_1383,N_1354);
or U1466 (N_1466,N_1325,N_1307);
nor U1467 (N_1467,N_1389,N_1319);
or U1468 (N_1468,N_1311,N_1351);
and U1469 (N_1469,N_1361,N_1359);
or U1470 (N_1470,N_1374,N_1304);
and U1471 (N_1471,N_1320,N_1397);
xor U1472 (N_1472,N_1372,N_1379);
xnor U1473 (N_1473,N_1342,N_1372);
nand U1474 (N_1474,N_1363,N_1316);
nor U1475 (N_1475,N_1386,N_1318);
nor U1476 (N_1476,N_1307,N_1320);
or U1477 (N_1477,N_1366,N_1376);
or U1478 (N_1478,N_1332,N_1397);
or U1479 (N_1479,N_1319,N_1338);
xnor U1480 (N_1480,N_1346,N_1331);
or U1481 (N_1481,N_1343,N_1393);
or U1482 (N_1482,N_1376,N_1325);
or U1483 (N_1483,N_1384,N_1316);
or U1484 (N_1484,N_1304,N_1315);
xnor U1485 (N_1485,N_1313,N_1308);
or U1486 (N_1486,N_1396,N_1381);
nor U1487 (N_1487,N_1318,N_1305);
nand U1488 (N_1488,N_1371,N_1391);
xor U1489 (N_1489,N_1352,N_1373);
or U1490 (N_1490,N_1394,N_1347);
nor U1491 (N_1491,N_1396,N_1362);
nand U1492 (N_1492,N_1345,N_1369);
nor U1493 (N_1493,N_1354,N_1361);
and U1494 (N_1494,N_1312,N_1366);
or U1495 (N_1495,N_1343,N_1388);
xnor U1496 (N_1496,N_1334,N_1374);
xor U1497 (N_1497,N_1330,N_1360);
nor U1498 (N_1498,N_1332,N_1305);
and U1499 (N_1499,N_1322,N_1379);
nand U1500 (N_1500,N_1472,N_1404);
nand U1501 (N_1501,N_1468,N_1419);
or U1502 (N_1502,N_1471,N_1497);
and U1503 (N_1503,N_1434,N_1494);
and U1504 (N_1504,N_1403,N_1420);
or U1505 (N_1505,N_1462,N_1492);
and U1506 (N_1506,N_1499,N_1423);
nand U1507 (N_1507,N_1467,N_1456);
nor U1508 (N_1508,N_1482,N_1415);
or U1509 (N_1509,N_1446,N_1422);
nand U1510 (N_1510,N_1491,N_1424);
or U1511 (N_1511,N_1455,N_1433);
nand U1512 (N_1512,N_1493,N_1475);
xor U1513 (N_1513,N_1451,N_1443);
and U1514 (N_1514,N_1410,N_1430);
or U1515 (N_1515,N_1438,N_1486);
nor U1516 (N_1516,N_1448,N_1452);
and U1517 (N_1517,N_1460,N_1425);
or U1518 (N_1518,N_1411,N_1461);
or U1519 (N_1519,N_1477,N_1406);
and U1520 (N_1520,N_1481,N_1436);
and U1521 (N_1521,N_1401,N_1498);
xor U1522 (N_1522,N_1407,N_1484);
nand U1523 (N_1523,N_1400,N_1487);
xnor U1524 (N_1524,N_1429,N_1426);
nand U1525 (N_1525,N_1454,N_1466);
or U1526 (N_1526,N_1457,N_1418);
xnor U1527 (N_1527,N_1495,N_1409);
xor U1528 (N_1528,N_1453,N_1464);
nor U1529 (N_1529,N_1469,N_1444);
and U1530 (N_1530,N_1476,N_1437);
or U1531 (N_1531,N_1450,N_1473);
or U1532 (N_1532,N_1442,N_1459);
and U1533 (N_1533,N_1428,N_1474);
and U1534 (N_1534,N_1490,N_1470);
or U1535 (N_1535,N_1458,N_1445);
nand U1536 (N_1536,N_1447,N_1421);
nor U1537 (N_1537,N_1417,N_1439);
and U1538 (N_1538,N_1416,N_1479);
and U1539 (N_1539,N_1463,N_1427);
nand U1540 (N_1540,N_1465,N_1483);
nand U1541 (N_1541,N_1408,N_1480);
nand U1542 (N_1542,N_1478,N_1440);
or U1543 (N_1543,N_1441,N_1435);
and U1544 (N_1544,N_1413,N_1489);
or U1545 (N_1545,N_1402,N_1488);
and U1546 (N_1546,N_1432,N_1405);
nor U1547 (N_1547,N_1414,N_1496);
nand U1548 (N_1548,N_1412,N_1431);
xor U1549 (N_1549,N_1485,N_1449);
and U1550 (N_1550,N_1459,N_1417);
and U1551 (N_1551,N_1440,N_1442);
and U1552 (N_1552,N_1495,N_1479);
nand U1553 (N_1553,N_1402,N_1492);
nand U1554 (N_1554,N_1420,N_1407);
xnor U1555 (N_1555,N_1440,N_1400);
xnor U1556 (N_1556,N_1413,N_1432);
nand U1557 (N_1557,N_1461,N_1447);
nor U1558 (N_1558,N_1459,N_1430);
nand U1559 (N_1559,N_1442,N_1480);
xor U1560 (N_1560,N_1453,N_1435);
and U1561 (N_1561,N_1413,N_1461);
and U1562 (N_1562,N_1420,N_1455);
xnor U1563 (N_1563,N_1403,N_1469);
or U1564 (N_1564,N_1417,N_1408);
and U1565 (N_1565,N_1488,N_1419);
nand U1566 (N_1566,N_1422,N_1415);
and U1567 (N_1567,N_1440,N_1466);
xnor U1568 (N_1568,N_1452,N_1405);
or U1569 (N_1569,N_1422,N_1418);
nand U1570 (N_1570,N_1498,N_1428);
nor U1571 (N_1571,N_1414,N_1498);
or U1572 (N_1572,N_1418,N_1450);
nand U1573 (N_1573,N_1406,N_1420);
nand U1574 (N_1574,N_1443,N_1485);
xnor U1575 (N_1575,N_1412,N_1423);
nor U1576 (N_1576,N_1431,N_1464);
nor U1577 (N_1577,N_1478,N_1422);
and U1578 (N_1578,N_1415,N_1448);
nor U1579 (N_1579,N_1417,N_1418);
nor U1580 (N_1580,N_1468,N_1433);
nor U1581 (N_1581,N_1471,N_1464);
and U1582 (N_1582,N_1441,N_1408);
xor U1583 (N_1583,N_1408,N_1412);
nor U1584 (N_1584,N_1420,N_1478);
and U1585 (N_1585,N_1405,N_1425);
nor U1586 (N_1586,N_1406,N_1407);
nand U1587 (N_1587,N_1452,N_1422);
nor U1588 (N_1588,N_1443,N_1435);
xor U1589 (N_1589,N_1495,N_1411);
and U1590 (N_1590,N_1482,N_1454);
nand U1591 (N_1591,N_1473,N_1455);
and U1592 (N_1592,N_1435,N_1417);
xor U1593 (N_1593,N_1418,N_1426);
xor U1594 (N_1594,N_1441,N_1413);
nor U1595 (N_1595,N_1438,N_1440);
nand U1596 (N_1596,N_1456,N_1497);
or U1597 (N_1597,N_1442,N_1473);
nor U1598 (N_1598,N_1416,N_1441);
nor U1599 (N_1599,N_1463,N_1402);
nor U1600 (N_1600,N_1596,N_1566);
and U1601 (N_1601,N_1510,N_1586);
xnor U1602 (N_1602,N_1541,N_1551);
or U1603 (N_1603,N_1569,N_1581);
and U1604 (N_1604,N_1574,N_1525);
or U1605 (N_1605,N_1594,N_1502);
xnor U1606 (N_1606,N_1591,N_1550);
and U1607 (N_1607,N_1599,N_1588);
and U1608 (N_1608,N_1504,N_1532);
nand U1609 (N_1609,N_1580,N_1563);
nand U1610 (N_1610,N_1535,N_1547);
nor U1611 (N_1611,N_1568,N_1593);
and U1612 (N_1612,N_1516,N_1571);
and U1613 (N_1613,N_1553,N_1520);
and U1614 (N_1614,N_1543,N_1572);
and U1615 (N_1615,N_1573,N_1511);
nor U1616 (N_1616,N_1555,N_1505);
xor U1617 (N_1617,N_1542,N_1509);
or U1618 (N_1618,N_1592,N_1519);
and U1619 (N_1619,N_1544,N_1552);
and U1620 (N_1620,N_1554,N_1538);
or U1621 (N_1621,N_1597,N_1560);
nor U1622 (N_1622,N_1557,N_1512);
nor U1623 (N_1623,N_1540,N_1575);
nor U1624 (N_1624,N_1503,N_1548);
nor U1625 (N_1625,N_1564,N_1518);
nor U1626 (N_1626,N_1579,N_1545);
nor U1627 (N_1627,N_1549,N_1501);
xor U1628 (N_1628,N_1528,N_1508);
nor U1629 (N_1629,N_1556,N_1590);
and U1630 (N_1630,N_1577,N_1559);
nor U1631 (N_1631,N_1534,N_1558);
xnor U1632 (N_1632,N_1567,N_1526);
or U1633 (N_1633,N_1584,N_1514);
or U1634 (N_1634,N_1570,N_1533);
nor U1635 (N_1635,N_1500,N_1578);
nor U1636 (N_1636,N_1589,N_1587);
nand U1637 (N_1637,N_1576,N_1582);
nor U1638 (N_1638,N_1565,N_1513);
xnor U1639 (N_1639,N_1517,N_1562);
nor U1640 (N_1640,N_1537,N_1529);
or U1641 (N_1641,N_1585,N_1539);
and U1642 (N_1642,N_1561,N_1507);
nor U1643 (N_1643,N_1530,N_1523);
nor U1644 (N_1644,N_1536,N_1583);
and U1645 (N_1645,N_1522,N_1598);
xor U1646 (N_1646,N_1521,N_1506);
nor U1647 (N_1647,N_1527,N_1515);
or U1648 (N_1648,N_1546,N_1531);
xor U1649 (N_1649,N_1595,N_1524);
and U1650 (N_1650,N_1549,N_1537);
xor U1651 (N_1651,N_1517,N_1595);
or U1652 (N_1652,N_1557,N_1569);
and U1653 (N_1653,N_1560,N_1590);
and U1654 (N_1654,N_1535,N_1525);
nand U1655 (N_1655,N_1532,N_1521);
and U1656 (N_1656,N_1557,N_1575);
and U1657 (N_1657,N_1574,N_1521);
and U1658 (N_1658,N_1588,N_1542);
or U1659 (N_1659,N_1564,N_1573);
xnor U1660 (N_1660,N_1583,N_1553);
nand U1661 (N_1661,N_1518,N_1526);
nor U1662 (N_1662,N_1504,N_1529);
xnor U1663 (N_1663,N_1570,N_1559);
nor U1664 (N_1664,N_1587,N_1578);
nand U1665 (N_1665,N_1523,N_1574);
and U1666 (N_1666,N_1513,N_1561);
and U1667 (N_1667,N_1522,N_1505);
nor U1668 (N_1668,N_1500,N_1549);
and U1669 (N_1669,N_1536,N_1571);
xor U1670 (N_1670,N_1588,N_1529);
nor U1671 (N_1671,N_1532,N_1517);
nor U1672 (N_1672,N_1537,N_1522);
nor U1673 (N_1673,N_1555,N_1504);
and U1674 (N_1674,N_1526,N_1530);
nor U1675 (N_1675,N_1500,N_1591);
and U1676 (N_1676,N_1509,N_1574);
and U1677 (N_1677,N_1541,N_1558);
xnor U1678 (N_1678,N_1516,N_1514);
and U1679 (N_1679,N_1543,N_1549);
or U1680 (N_1680,N_1552,N_1561);
or U1681 (N_1681,N_1549,N_1579);
or U1682 (N_1682,N_1596,N_1573);
or U1683 (N_1683,N_1535,N_1599);
xor U1684 (N_1684,N_1557,N_1594);
or U1685 (N_1685,N_1586,N_1569);
or U1686 (N_1686,N_1598,N_1525);
xor U1687 (N_1687,N_1566,N_1525);
nor U1688 (N_1688,N_1524,N_1551);
nor U1689 (N_1689,N_1537,N_1584);
nor U1690 (N_1690,N_1575,N_1589);
nor U1691 (N_1691,N_1553,N_1515);
xor U1692 (N_1692,N_1563,N_1590);
xor U1693 (N_1693,N_1518,N_1549);
nand U1694 (N_1694,N_1512,N_1563);
xor U1695 (N_1695,N_1527,N_1573);
nand U1696 (N_1696,N_1545,N_1553);
and U1697 (N_1697,N_1564,N_1520);
xor U1698 (N_1698,N_1560,N_1541);
xor U1699 (N_1699,N_1596,N_1548);
xor U1700 (N_1700,N_1650,N_1616);
nand U1701 (N_1701,N_1611,N_1600);
nor U1702 (N_1702,N_1601,N_1657);
xnor U1703 (N_1703,N_1617,N_1667);
nand U1704 (N_1704,N_1694,N_1638);
nand U1705 (N_1705,N_1663,N_1665);
xor U1706 (N_1706,N_1634,N_1624);
or U1707 (N_1707,N_1619,N_1675);
xor U1708 (N_1708,N_1692,N_1636);
and U1709 (N_1709,N_1643,N_1699);
or U1710 (N_1710,N_1605,N_1677);
xor U1711 (N_1711,N_1639,N_1632);
or U1712 (N_1712,N_1683,N_1696);
xnor U1713 (N_1713,N_1630,N_1681);
xor U1714 (N_1714,N_1631,N_1620);
nand U1715 (N_1715,N_1664,N_1647);
or U1716 (N_1716,N_1635,N_1658);
or U1717 (N_1717,N_1618,N_1602);
xor U1718 (N_1718,N_1660,N_1613);
and U1719 (N_1719,N_1606,N_1676);
xor U1720 (N_1720,N_1615,N_1673);
nand U1721 (N_1721,N_1689,N_1648);
and U1722 (N_1722,N_1695,N_1644);
and U1723 (N_1723,N_1637,N_1687);
xnor U1724 (N_1724,N_1656,N_1642);
xnor U1725 (N_1725,N_1668,N_1679);
and U1726 (N_1726,N_1672,N_1621);
or U1727 (N_1727,N_1646,N_1623);
or U1728 (N_1728,N_1659,N_1612);
nand U1729 (N_1729,N_1669,N_1609);
or U1730 (N_1730,N_1625,N_1655);
nor U1731 (N_1731,N_1652,N_1671);
and U1732 (N_1732,N_1608,N_1653);
nand U1733 (N_1733,N_1690,N_1654);
nand U1734 (N_1734,N_1649,N_1628);
xnor U1735 (N_1735,N_1622,N_1614);
and U1736 (N_1736,N_1678,N_1686);
nand U1737 (N_1737,N_1645,N_1698);
xor U1738 (N_1738,N_1688,N_1697);
nor U1739 (N_1739,N_1610,N_1607);
or U1740 (N_1740,N_1691,N_1662);
xnor U1741 (N_1741,N_1661,N_1633);
nand U1742 (N_1742,N_1666,N_1684);
and U1743 (N_1743,N_1626,N_1629);
and U1744 (N_1744,N_1640,N_1641);
xnor U1745 (N_1745,N_1693,N_1685);
xor U1746 (N_1746,N_1627,N_1651);
xor U1747 (N_1747,N_1670,N_1604);
nor U1748 (N_1748,N_1603,N_1674);
xor U1749 (N_1749,N_1682,N_1680);
nand U1750 (N_1750,N_1609,N_1652);
or U1751 (N_1751,N_1681,N_1610);
nor U1752 (N_1752,N_1661,N_1686);
nor U1753 (N_1753,N_1687,N_1615);
and U1754 (N_1754,N_1656,N_1661);
nor U1755 (N_1755,N_1685,N_1694);
or U1756 (N_1756,N_1654,N_1640);
xnor U1757 (N_1757,N_1676,N_1671);
or U1758 (N_1758,N_1655,N_1616);
nand U1759 (N_1759,N_1615,N_1657);
nor U1760 (N_1760,N_1646,N_1676);
and U1761 (N_1761,N_1617,N_1644);
and U1762 (N_1762,N_1625,N_1604);
and U1763 (N_1763,N_1694,N_1698);
or U1764 (N_1764,N_1635,N_1630);
xnor U1765 (N_1765,N_1696,N_1661);
xor U1766 (N_1766,N_1651,N_1692);
or U1767 (N_1767,N_1699,N_1606);
nor U1768 (N_1768,N_1645,N_1676);
and U1769 (N_1769,N_1614,N_1617);
xor U1770 (N_1770,N_1623,N_1661);
nand U1771 (N_1771,N_1632,N_1603);
and U1772 (N_1772,N_1639,N_1663);
xor U1773 (N_1773,N_1624,N_1630);
nor U1774 (N_1774,N_1638,N_1699);
nor U1775 (N_1775,N_1698,N_1685);
nand U1776 (N_1776,N_1642,N_1651);
nor U1777 (N_1777,N_1618,N_1616);
nand U1778 (N_1778,N_1604,N_1610);
or U1779 (N_1779,N_1651,N_1625);
or U1780 (N_1780,N_1655,N_1656);
nand U1781 (N_1781,N_1683,N_1686);
nor U1782 (N_1782,N_1663,N_1643);
xor U1783 (N_1783,N_1642,N_1626);
nand U1784 (N_1784,N_1659,N_1605);
or U1785 (N_1785,N_1652,N_1616);
xor U1786 (N_1786,N_1671,N_1609);
and U1787 (N_1787,N_1663,N_1695);
or U1788 (N_1788,N_1680,N_1628);
nor U1789 (N_1789,N_1634,N_1606);
and U1790 (N_1790,N_1671,N_1602);
nor U1791 (N_1791,N_1682,N_1630);
xnor U1792 (N_1792,N_1640,N_1635);
or U1793 (N_1793,N_1653,N_1683);
nor U1794 (N_1794,N_1686,N_1606);
and U1795 (N_1795,N_1648,N_1603);
or U1796 (N_1796,N_1647,N_1608);
xnor U1797 (N_1797,N_1699,N_1620);
nor U1798 (N_1798,N_1611,N_1637);
and U1799 (N_1799,N_1632,N_1649);
and U1800 (N_1800,N_1746,N_1736);
or U1801 (N_1801,N_1725,N_1724);
xnor U1802 (N_1802,N_1704,N_1774);
or U1803 (N_1803,N_1706,N_1701);
xor U1804 (N_1804,N_1723,N_1733);
nand U1805 (N_1805,N_1703,N_1782);
and U1806 (N_1806,N_1790,N_1709);
xor U1807 (N_1807,N_1743,N_1702);
xnor U1808 (N_1808,N_1793,N_1744);
xor U1809 (N_1809,N_1787,N_1776);
or U1810 (N_1810,N_1763,N_1722);
xor U1811 (N_1811,N_1786,N_1758);
and U1812 (N_1812,N_1707,N_1711);
nand U1813 (N_1813,N_1789,N_1796);
xor U1814 (N_1814,N_1767,N_1769);
or U1815 (N_1815,N_1781,N_1757);
nor U1816 (N_1816,N_1764,N_1710);
nor U1817 (N_1817,N_1783,N_1745);
nor U1818 (N_1818,N_1751,N_1700);
or U1819 (N_1819,N_1772,N_1747);
or U1820 (N_1820,N_1729,N_1737);
or U1821 (N_1821,N_1740,N_1770);
nor U1822 (N_1822,N_1752,N_1732);
nor U1823 (N_1823,N_1756,N_1777);
nand U1824 (N_1824,N_1726,N_1731);
and U1825 (N_1825,N_1759,N_1748);
nor U1826 (N_1826,N_1784,N_1753);
or U1827 (N_1827,N_1798,N_1773);
and U1828 (N_1828,N_1791,N_1760);
nor U1829 (N_1829,N_1713,N_1788);
xor U1830 (N_1830,N_1718,N_1761);
or U1831 (N_1831,N_1720,N_1750);
or U1832 (N_1832,N_1727,N_1765);
or U1833 (N_1833,N_1719,N_1741);
nor U1834 (N_1834,N_1794,N_1792);
or U1835 (N_1835,N_1717,N_1766);
and U1836 (N_1836,N_1739,N_1768);
and U1837 (N_1837,N_1778,N_1749);
or U1838 (N_1838,N_1754,N_1721);
nand U1839 (N_1839,N_1738,N_1755);
nor U1840 (N_1840,N_1714,N_1715);
nor U1841 (N_1841,N_1735,N_1708);
or U1842 (N_1842,N_1797,N_1775);
nor U1843 (N_1843,N_1780,N_1795);
or U1844 (N_1844,N_1712,N_1734);
nor U1845 (N_1845,N_1779,N_1716);
nand U1846 (N_1846,N_1705,N_1730);
xor U1847 (N_1847,N_1762,N_1742);
nor U1848 (N_1848,N_1728,N_1771);
or U1849 (N_1849,N_1785,N_1799);
nor U1850 (N_1850,N_1762,N_1794);
xnor U1851 (N_1851,N_1712,N_1713);
nor U1852 (N_1852,N_1725,N_1741);
or U1853 (N_1853,N_1746,N_1738);
and U1854 (N_1854,N_1758,N_1743);
nand U1855 (N_1855,N_1761,N_1798);
nand U1856 (N_1856,N_1702,N_1766);
nand U1857 (N_1857,N_1730,N_1756);
nand U1858 (N_1858,N_1716,N_1741);
or U1859 (N_1859,N_1738,N_1727);
xnor U1860 (N_1860,N_1780,N_1786);
nor U1861 (N_1861,N_1770,N_1746);
and U1862 (N_1862,N_1758,N_1746);
or U1863 (N_1863,N_1765,N_1763);
and U1864 (N_1864,N_1737,N_1784);
xnor U1865 (N_1865,N_1759,N_1719);
nor U1866 (N_1866,N_1761,N_1774);
and U1867 (N_1867,N_1722,N_1760);
xor U1868 (N_1868,N_1702,N_1768);
xor U1869 (N_1869,N_1724,N_1770);
and U1870 (N_1870,N_1775,N_1789);
xor U1871 (N_1871,N_1772,N_1705);
nor U1872 (N_1872,N_1749,N_1760);
xnor U1873 (N_1873,N_1772,N_1766);
nor U1874 (N_1874,N_1732,N_1796);
nand U1875 (N_1875,N_1787,N_1713);
or U1876 (N_1876,N_1779,N_1735);
xnor U1877 (N_1877,N_1774,N_1756);
or U1878 (N_1878,N_1737,N_1751);
nand U1879 (N_1879,N_1761,N_1715);
nand U1880 (N_1880,N_1787,N_1755);
nor U1881 (N_1881,N_1759,N_1700);
nand U1882 (N_1882,N_1755,N_1770);
or U1883 (N_1883,N_1798,N_1794);
and U1884 (N_1884,N_1797,N_1798);
nand U1885 (N_1885,N_1782,N_1724);
nor U1886 (N_1886,N_1790,N_1760);
xor U1887 (N_1887,N_1764,N_1751);
xor U1888 (N_1888,N_1772,N_1710);
and U1889 (N_1889,N_1753,N_1763);
xnor U1890 (N_1890,N_1792,N_1789);
nor U1891 (N_1891,N_1777,N_1726);
and U1892 (N_1892,N_1733,N_1738);
or U1893 (N_1893,N_1786,N_1724);
nand U1894 (N_1894,N_1775,N_1771);
nand U1895 (N_1895,N_1733,N_1792);
and U1896 (N_1896,N_1785,N_1771);
nand U1897 (N_1897,N_1736,N_1744);
xnor U1898 (N_1898,N_1736,N_1721);
or U1899 (N_1899,N_1758,N_1767);
or U1900 (N_1900,N_1855,N_1879);
and U1901 (N_1901,N_1842,N_1846);
nand U1902 (N_1902,N_1825,N_1892);
nand U1903 (N_1903,N_1851,N_1848);
and U1904 (N_1904,N_1841,N_1813);
or U1905 (N_1905,N_1862,N_1861);
or U1906 (N_1906,N_1828,N_1822);
nand U1907 (N_1907,N_1808,N_1865);
xnor U1908 (N_1908,N_1870,N_1845);
nor U1909 (N_1909,N_1849,N_1804);
nand U1910 (N_1910,N_1812,N_1875);
nand U1911 (N_1911,N_1807,N_1885);
nor U1912 (N_1912,N_1884,N_1877);
xor U1913 (N_1913,N_1814,N_1886);
nand U1914 (N_1914,N_1834,N_1881);
or U1915 (N_1915,N_1837,N_1840);
and U1916 (N_1916,N_1850,N_1810);
xnor U1917 (N_1917,N_1817,N_1864);
xnor U1918 (N_1918,N_1836,N_1898);
xor U1919 (N_1919,N_1895,N_1878);
nor U1920 (N_1920,N_1843,N_1889);
nor U1921 (N_1921,N_1867,N_1899);
nand U1922 (N_1922,N_1826,N_1897);
nand U1923 (N_1923,N_1887,N_1830);
nor U1924 (N_1924,N_1815,N_1880);
nor U1925 (N_1925,N_1863,N_1874);
or U1926 (N_1926,N_1882,N_1896);
nand U1927 (N_1927,N_1827,N_1859);
nand U1928 (N_1928,N_1891,N_1833);
or U1929 (N_1929,N_1869,N_1811);
and U1930 (N_1930,N_1858,N_1801);
xnor U1931 (N_1931,N_1866,N_1873);
nand U1932 (N_1932,N_1824,N_1857);
nor U1933 (N_1933,N_1894,N_1802);
nand U1934 (N_1934,N_1809,N_1818);
xor U1935 (N_1935,N_1868,N_1803);
nor U1936 (N_1936,N_1800,N_1872);
nand U1937 (N_1937,N_1806,N_1844);
and U1938 (N_1938,N_1883,N_1860);
or U1939 (N_1939,N_1821,N_1820);
nor U1940 (N_1940,N_1823,N_1838);
nor U1941 (N_1941,N_1847,N_1832);
and U1942 (N_1942,N_1876,N_1871);
or U1943 (N_1943,N_1888,N_1890);
nand U1944 (N_1944,N_1839,N_1854);
or U1945 (N_1945,N_1853,N_1852);
or U1946 (N_1946,N_1819,N_1831);
and U1947 (N_1947,N_1856,N_1829);
xor U1948 (N_1948,N_1805,N_1893);
nand U1949 (N_1949,N_1835,N_1816);
and U1950 (N_1950,N_1881,N_1816);
nand U1951 (N_1951,N_1877,N_1852);
nor U1952 (N_1952,N_1893,N_1858);
nand U1953 (N_1953,N_1884,N_1858);
xnor U1954 (N_1954,N_1835,N_1820);
nand U1955 (N_1955,N_1832,N_1878);
nor U1956 (N_1956,N_1868,N_1879);
xor U1957 (N_1957,N_1885,N_1820);
xor U1958 (N_1958,N_1849,N_1806);
xnor U1959 (N_1959,N_1818,N_1866);
xnor U1960 (N_1960,N_1859,N_1854);
nand U1961 (N_1961,N_1882,N_1843);
xor U1962 (N_1962,N_1837,N_1822);
nor U1963 (N_1963,N_1868,N_1841);
nand U1964 (N_1964,N_1844,N_1878);
or U1965 (N_1965,N_1812,N_1872);
nand U1966 (N_1966,N_1846,N_1818);
and U1967 (N_1967,N_1892,N_1880);
nor U1968 (N_1968,N_1855,N_1827);
nor U1969 (N_1969,N_1811,N_1845);
xor U1970 (N_1970,N_1887,N_1831);
xnor U1971 (N_1971,N_1812,N_1879);
or U1972 (N_1972,N_1893,N_1829);
nand U1973 (N_1973,N_1883,N_1851);
xnor U1974 (N_1974,N_1851,N_1881);
and U1975 (N_1975,N_1813,N_1874);
or U1976 (N_1976,N_1827,N_1839);
nor U1977 (N_1977,N_1833,N_1840);
nand U1978 (N_1978,N_1821,N_1896);
or U1979 (N_1979,N_1825,N_1886);
or U1980 (N_1980,N_1854,N_1811);
xnor U1981 (N_1981,N_1864,N_1867);
or U1982 (N_1982,N_1815,N_1882);
nor U1983 (N_1983,N_1893,N_1859);
and U1984 (N_1984,N_1815,N_1860);
nand U1985 (N_1985,N_1861,N_1883);
and U1986 (N_1986,N_1892,N_1883);
or U1987 (N_1987,N_1882,N_1863);
or U1988 (N_1988,N_1804,N_1866);
and U1989 (N_1989,N_1851,N_1836);
nand U1990 (N_1990,N_1863,N_1861);
and U1991 (N_1991,N_1836,N_1857);
nor U1992 (N_1992,N_1868,N_1852);
nor U1993 (N_1993,N_1830,N_1878);
nand U1994 (N_1994,N_1874,N_1816);
xnor U1995 (N_1995,N_1881,N_1878);
nand U1996 (N_1996,N_1874,N_1868);
nor U1997 (N_1997,N_1839,N_1855);
nor U1998 (N_1998,N_1845,N_1851);
and U1999 (N_1999,N_1872,N_1888);
and U2000 (N_2000,N_1904,N_1988);
and U2001 (N_2001,N_1999,N_1973);
nor U2002 (N_2002,N_1913,N_1911);
or U2003 (N_2003,N_1972,N_1980);
nand U2004 (N_2004,N_1921,N_1953);
and U2005 (N_2005,N_1923,N_1938);
or U2006 (N_2006,N_1984,N_1914);
xor U2007 (N_2007,N_1956,N_1951);
xnor U2008 (N_2008,N_1910,N_1902);
nor U2009 (N_2009,N_1978,N_1982);
nand U2010 (N_2010,N_1907,N_1926);
or U2011 (N_2011,N_1967,N_1995);
nor U2012 (N_2012,N_1935,N_1991);
nand U2013 (N_2013,N_1985,N_1922);
and U2014 (N_2014,N_1976,N_1981);
nand U2015 (N_2015,N_1965,N_1974);
nor U2016 (N_2016,N_1936,N_1954);
xnor U2017 (N_2017,N_1919,N_1942);
and U2018 (N_2018,N_1968,N_1960);
and U2019 (N_2019,N_1949,N_1996);
nor U2020 (N_2020,N_1971,N_1961);
and U2021 (N_2021,N_1916,N_1966);
or U2022 (N_2022,N_1952,N_1920);
or U2023 (N_2023,N_1962,N_1948);
nor U2024 (N_2024,N_1928,N_1941);
nor U2025 (N_2025,N_1934,N_1957);
nand U2026 (N_2026,N_1963,N_1925);
nor U2027 (N_2027,N_1959,N_1931);
or U2028 (N_2028,N_1929,N_1924);
nor U2029 (N_2029,N_1930,N_1946);
nor U2030 (N_2030,N_1908,N_1932);
and U2031 (N_2031,N_1998,N_1986);
nor U2032 (N_2032,N_1917,N_1958);
and U2033 (N_2033,N_1945,N_1950);
and U2034 (N_2034,N_1979,N_1912);
nor U2035 (N_2035,N_1983,N_1947);
and U2036 (N_2036,N_1901,N_1927);
xnor U2037 (N_2037,N_1939,N_1937);
or U2038 (N_2038,N_1906,N_1918);
nand U2039 (N_2039,N_1989,N_1915);
nand U2040 (N_2040,N_1993,N_1994);
nor U2041 (N_2041,N_1964,N_1909);
nor U2042 (N_2042,N_1905,N_1903);
nand U2043 (N_2043,N_1933,N_1940);
nor U2044 (N_2044,N_1943,N_1992);
nor U2045 (N_2045,N_1969,N_1997);
xor U2046 (N_2046,N_1970,N_1987);
nor U2047 (N_2047,N_1990,N_1944);
and U2048 (N_2048,N_1975,N_1977);
and U2049 (N_2049,N_1900,N_1955);
nor U2050 (N_2050,N_1956,N_1948);
and U2051 (N_2051,N_1963,N_1980);
xnor U2052 (N_2052,N_1928,N_1965);
nor U2053 (N_2053,N_1940,N_1979);
and U2054 (N_2054,N_1981,N_1973);
and U2055 (N_2055,N_1918,N_1962);
xnor U2056 (N_2056,N_1979,N_1927);
nor U2057 (N_2057,N_1913,N_1920);
or U2058 (N_2058,N_1975,N_1923);
or U2059 (N_2059,N_1974,N_1991);
nand U2060 (N_2060,N_1956,N_1992);
xnor U2061 (N_2061,N_1927,N_1919);
or U2062 (N_2062,N_1914,N_1912);
xnor U2063 (N_2063,N_1999,N_1960);
and U2064 (N_2064,N_1995,N_1993);
or U2065 (N_2065,N_1957,N_1970);
xor U2066 (N_2066,N_1957,N_1988);
nor U2067 (N_2067,N_1932,N_1939);
nor U2068 (N_2068,N_1953,N_1972);
xnor U2069 (N_2069,N_1902,N_1928);
xnor U2070 (N_2070,N_1907,N_1909);
and U2071 (N_2071,N_1923,N_1968);
nor U2072 (N_2072,N_1987,N_1905);
xnor U2073 (N_2073,N_1970,N_1978);
and U2074 (N_2074,N_1971,N_1920);
and U2075 (N_2075,N_1938,N_1947);
nor U2076 (N_2076,N_1903,N_1932);
nor U2077 (N_2077,N_1973,N_1907);
nor U2078 (N_2078,N_1949,N_1911);
and U2079 (N_2079,N_1906,N_1982);
nor U2080 (N_2080,N_1932,N_1977);
nor U2081 (N_2081,N_1986,N_1901);
and U2082 (N_2082,N_1923,N_1981);
and U2083 (N_2083,N_1924,N_1913);
or U2084 (N_2084,N_1979,N_1948);
nand U2085 (N_2085,N_1992,N_1967);
nand U2086 (N_2086,N_1996,N_1921);
or U2087 (N_2087,N_1916,N_1979);
nand U2088 (N_2088,N_1970,N_1966);
and U2089 (N_2089,N_1999,N_1977);
and U2090 (N_2090,N_1998,N_1930);
or U2091 (N_2091,N_1980,N_1954);
xor U2092 (N_2092,N_1976,N_1990);
nand U2093 (N_2093,N_1936,N_1968);
nand U2094 (N_2094,N_1994,N_1903);
nand U2095 (N_2095,N_1955,N_1968);
and U2096 (N_2096,N_1979,N_1995);
and U2097 (N_2097,N_1991,N_1957);
xor U2098 (N_2098,N_1913,N_1993);
xor U2099 (N_2099,N_1927,N_1907);
or U2100 (N_2100,N_2064,N_2056);
nor U2101 (N_2101,N_2035,N_2019);
or U2102 (N_2102,N_2024,N_2077);
or U2103 (N_2103,N_2055,N_2093);
nand U2104 (N_2104,N_2042,N_2003);
and U2105 (N_2105,N_2052,N_2005);
nor U2106 (N_2106,N_2018,N_2022);
and U2107 (N_2107,N_2058,N_2029);
nor U2108 (N_2108,N_2076,N_2082);
nand U2109 (N_2109,N_2090,N_2075);
nand U2110 (N_2110,N_2095,N_2060);
xnor U2111 (N_2111,N_2021,N_2063);
or U2112 (N_2112,N_2013,N_2047);
and U2113 (N_2113,N_2096,N_2037);
xnor U2114 (N_2114,N_2083,N_2000);
nand U2115 (N_2115,N_2089,N_2034);
xnor U2116 (N_2116,N_2030,N_2009);
nor U2117 (N_2117,N_2010,N_2062);
xnor U2118 (N_2118,N_2080,N_2026);
nor U2119 (N_2119,N_2054,N_2012);
or U2120 (N_2120,N_2065,N_2094);
nand U2121 (N_2121,N_2008,N_2087);
nor U2122 (N_2122,N_2039,N_2023);
xor U2123 (N_2123,N_2044,N_2099);
nand U2124 (N_2124,N_2001,N_2081);
nand U2125 (N_2125,N_2011,N_2086);
nand U2126 (N_2126,N_2006,N_2067);
or U2127 (N_2127,N_2079,N_2051);
nand U2128 (N_2128,N_2040,N_2031);
and U2129 (N_2129,N_2068,N_2057);
nand U2130 (N_2130,N_2069,N_2088);
or U2131 (N_2131,N_2041,N_2091);
nor U2132 (N_2132,N_2061,N_2049);
nor U2133 (N_2133,N_2045,N_2098);
or U2134 (N_2134,N_2073,N_2017);
or U2135 (N_2135,N_2085,N_2007);
or U2136 (N_2136,N_2092,N_2002);
nand U2137 (N_2137,N_2016,N_2074);
and U2138 (N_2138,N_2097,N_2028);
xnor U2139 (N_2139,N_2046,N_2071);
nor U2140 (N_2140,N_2025,N_2070);
nand U2141 (N_2141,N_2053,N_2027);
or U2142 (N_2142,N_2036,N_2059);
and U2143 (N_2143,N_2048,N_2032);
and U2144 (N_2144,N_2043,N_2066);
xnor U2145 (N_2145,N_2050,N_2078);
nor U2146 (N_2146,N_2020,N_2015);
nand U2147 (N_2147,N_2014,N_2072);
xnor U2148 (N_2148,N_2084,N_2004);
nor U2149 (N_2149,N_2033,N_2038);
or U2150 (N_2150,N_2042,N_2011);
xor U2151 (N_2151,N_2045,N_2080);
or U2152 (N_2152,N_2071,N_2057);
xnor U2153 (N_2153,N_2010,N_2038);
and U2154 (N_2154,N_2018,N_2030);
nand U2155 (N_2155,N_2023,N_2075);
or U2156 (N_2156,N_2056,N_2011);
nand U2157 (N_2157,N_2037,N_2036);
xor U2158 (N_2158,N_2035,N_2000);
nor U2159 (N_2159,N_2037,N_2070);
nand U2160 (N_2160,N_2009,N_2031);
xnor U2161 (N_2161,N_2011,N_2070);
and U2162 (N_2162,N_2094,N_2067);
nand U2163 (N_2163,N_2008,N_2051);
xnor U2164 (N_2164,N_2060,N_2087);
nand U2165 (N_2165,N_2023,N_2006);
xnor U2166 (N_2166,N_2036,N_2009);
nand U2167 (N_2167,N_2032,N_2094);
nand U2168 (N_2168,N_2026,N_2079);
or U2169 (N_2169,N_2001,N_2076);
and U2170 (N_2170,N_2026,N_2007);
and U2171 (N_2171,N_2072,N_2019);
xor U2172 (N_2172,N_2087,N_2073);
nor U2173 (N_2173,N_2093,N_2034);
nand U2174 (N_2174,N_2070,N_2056);
nor U2175 (N_2175,N_2000,N_2037);
nor U2176 (N_2176,N_2087,N_2023);
xor U2177 (N_2177,N_2075,N_2088);
xnor U2178 (N_2178,N_2082,N_2041);
xnor U2179 (N_2179,N_2071,N_2025);
or U2180 (N_2180,N_2052,N_2031);
and U2181 (N_2181,N_2061,N_2040);
xnor U2182 (N_2182,N_2021,N_2020);
or U2183 (N_2183,N_2015,N_2030);
and U2184 (N_2184,N_2035,N_2051);
and U2185 (N_2185,N_2028,N_2018);
nor U2186 (N_2186,N_2016,N_2001);
and U2187 (N_2187,N_2081,N_2068);
nor U2188 (N_2188,N_2090,N_2031);
xnor U2189 (N_2189,N_2011,N_2074);
nor U2190 (N_2190,N_2078,N_2026);
and U2191 (N_2191,N_2003,N_2058);
nor U2192 (N_2192,N_2020,N_2027);
nor U2193 (N_2193,N_2045,N_2000);
nor U2194 (N_2194,N_2076,N_2099);
and U2195 (N_2195,N_2056,N_2032);
nand U2196 (N_2196,N_2049,N_2011);
or U2197 (N_2197,N_2095,N_2062);
nand U2198 (N_2198,N_2022,N_2024);
and U2199 (N_2199,N_2048,N_2005);
and U2200 (N_2200,N_2119,N_2186);
and U2201 (N_2201,N_2158,N_2177);
nand U2202 (N_2202,N_2147,N_2194);
or U2203 (N_2203,N_2195,N_2150);
or U2204 (N_2204,N_2159,N_2122);
xnor U2205 (N_2205,N_2130,N_2167);
and U2206 (N_2206,N_2164,N_2107);
xor U2207 (N_2207,N_2187,N_2125);
and U2208 (N_2208,N_2175,N_2189);
nand U2209 (N_2209,N_2115,N_2138);
or U2210 (N_2210,N_2104,N_2131);
xor U2211 (N_2211,N_2139,N_2153);
and U2212 (N_2212,N_2100,N_2149);
nand U2213 (N_2213,N_2113,N_2181);
and U2214 (N_2214,N_2141,N_2182);
or U2215 (N_2215,N_2155,N_2180);
nand U2216 (N_2216,N_2143,N_2156);
and U2217 (N_2217,N_2197,N_2133);
nand U2218 (N_2218,N_2191,N_2116);
and U2219 (N_2219,N_2166,N_2190);
nor U2220 (N_2220,N_2184,N_2126);
or U2221 (N_2221,N_2146,N_2151);
and U2222 (N_2222,N_2185,N_2179);
and U2223 (N_2223,N_2193,N_2171);
and U2224 (N_2224,N_2142,N_2127);
xor U2225 (N_2225,N_2120,N_2148);
or U2226 (N_2226,N_2114,N_2144);
or U2227 (N_2227,N_2165,N_2168);
and U2228 (N_2228,N_2109,N_2110);
or U2229 (N_2229,N_2196,N_2183);
and U2230 (N_2230,N_2198,N_2137);
nor U2231 (N_2231,N_2154,N_2140);
nor U2232 (N_2232,N_2123,N_2136);
xor U2233 (N_2233,N_2169,N_2117);
xor U2234 (N_2234,N_2124,N_2134);
nand U2235 (N_2235,N_2172,N_2192);
xor U2236 (N_2236,N_2163,N_2157);
xnor U2237 (N_2237,N_2188,N_2106);
nand U2238 (N_2238,N_2111,N_2129);
xor U2239 (N_2239,N_2135,N_2176);
nand U2240 (N_2240,N_2108,N_2174);
and U2241 (N_2241,N_2112,N_2118);
nor U2242 (N_2242,N_2170,N_2101);
and U2243 (N_2243,N_2178,N_2132);
nor U2244 (N_2244,N_2105,N_2145);
nor U2245 (N_2245,N_2199,N_2128);
or U2246 (N_2246,N_2160,N_2121);
or U2247 (N_2247,N_2161,N_2152);
nand U2248 (N_2248,N_2173,N_2103);
or U2249 (N_2249,N_2102,N_2162);
nand U2250 (N_2250,N_2185,N_2123);
xor U2251 (N_2251,N_2124,N_2128);
xor U2252 (N_2252,N_2147,N_2197);
nor U2253 (N_2253,N_2184,N_2170);
nor U2254 (N_2254,N_2170,N_2149);
nand U2255 (N_2255,N_2152,N_2191);
and U2256 (N_2256,N_2164,N_2110);
nand U2257 (N_2257,N_2102,N_2126);
or U2258 (N_2258,N_2161,N_2127);
nor U2259 (N_2259,N_2148,N_2198);
nor U2260 (N_2260,N_2100,N_2117);
nand U2261 (N_2261,N_2149,N_2189);
and U2262 (N_2262,N_2155,N_2116);
xnor U2263 (N_2263,N_2190,N_2179);
or U2264 (N_2264,N_2104,N_2187);
or U2265 (N_2265,N_2152,N_2184);
and U2266 (N_2266,N_2190,N_2186);
nand U2267 (N_2267,N_2173,N_2185);
or U2268 (N_2268,N_2144,N_2103);
and U2269 (N_2269,N_2116,N_2184);
nor U2270 (N_2270,N_2121,N_2150);
nor U2271 (N_2271,N_2112,N_2144);
and U2272 (N_2272,N_2160,N_2170);
and U2273 (N_2273,N_2146,N_2142);
or U2274 (N_2274,N_2165,N_2163);
nor U2275 (N_2275,N_2133,N_2147);
nand U2276 (N_2276,N_2125,N_2104);
nand U2277 (N_2277,N_2170,N_2197);
and U2278 (N_2278,N_2157,N_2175);
and U2279 (N_2279,N_2151,N_2133);
xnor U2280 (N_2280,N_2131,N_2101);
nor U2281 (N_2281,N_2103,N_2167);
xor U2282 (N_2282,N_2122,N_2147);
nand U2283 (N_2283,N_2104,N_2133);
or U2284 (N_2284,N_2144,N_2125);
nor U2285 (N_2285,N_2145,N_2173);
nand U2286 (N_2286,N_2148,N_2156);
and U2287 (N_2287,N_2195,N_2136);
and U2288 (N_2288,N_2167,N_2169);
nand U2289 (N_2289,N_2158,N_2166);
xnor U2290 (N_2290,N_2134,N_2149);
xnor U2291 (N_2291,N_2133,N_2167);
nor U2292 (N_2292,N_2131,N_2115);
and U2293 (N_2293,N_2178,N_2173);
or U2294 (N_2294,N_2196,N_2137);
or U2295 (N_2295,N_2116,N_2104);
or U2296 (N_2296,N_2183,N_2124);
nor U2297 (N_2297,N_2154,N_2189);
nor U2298 (N_2298,N_2128,N_2174);
nor U2299 (N_2299,N_2117,N_2177);
xnor U2300 (N_2300,N_2243,N_2204);
nand U2301 (N_2301,N_2276,N_2232);
nand U2302 (N_2302,N_2264,N_2293);
and U2303 (N_2303,N_2258,N_2255);
and U2304 (N_2304,N_2201,N_2205);
nand U2305 (N_2305,N_2228,N_2267);
or U2306 (N_2306,N_2209,N_2288);
xor U2307 (N_2307,N_2286,N_2256);
and U2308 (N_2308,N_2225,N_2274);
and U2309 (N_2309,N_2237,N_2220);
nand U2310 (N_2310,N_2221,N_2259);
or U2311 (N_2311,N_2252,N_2294);
or U2312 (N_2312,N_2226,N_2246);
and U2313 (N_2313,N_2265,N_2291);
nor U2314 (N_2314,N_2257,N_2292);
and U2315 (N_2315,N_2270,N_2290);
xor U2316 (N_2316,N_2296,N_2297);
or U2317 (N_2317,N_2280,N_2240);
and U2318 (N_2318,N_2244,N_2233);
nor U2319 (N_2319,N_2223,N_2238);
or U2320 (N_2320,N_2262,N_2222);
xor U2321 (N_2321,N_2212,N_2211);
or U2322 (N_2322,N_2299,N_2284);
and U2323 (N_2323,N_2208,N_2202);
and U2324 (N_2324,N_2253,N_2279);
nor U2325 (N_2325,N_2250,N_2227);
xnor U2326 (N_2326,N_2295,N_2241);
or U2327 (N_2327,N_2216,N_2218);
and U2328 (N_2328,N_2200,N_2224);
or U2329 (N_2329,N_2247,N_2206);
and U2330 (N_2330,N_2272,N_2245);
and U2331 (N_2331,N_2236,N_2203);
and U2332 (N_2332,N_2254,N_2282);
or U2333 (N_2333,N_2242,N_2213);
and U2334 (N_2334,N_2283,N_2230);
and U2335 (N_2335,N_2281,N_2234);
or U2336 (N_2336,N_2273,N_2249);
and U2337 (N_2337,N_2251,N_2277);
or U2338 (N_2338,N_2214,N_2266);
xnor U2339 (N_2339,N_2268,N_2261);
and U2340 (N_2340,N_2263,N_2275);
or U2341 (N_2341,N_2260,N_2235);
nand U2342 (N_2342,N_2285,N_2271);
or U2343 (N_2343,N_2248,N_2229);
xor U2344 (N_2344,N_2217,N_2207);
or U2345 (N_2345,N_2210,N_2239);
xor U2346 (N_2346,N_2215,N_2269);
or U2347 (N_2347,N_2289,N_2278);
or U2348 (N_2348,N_2219,N_2287);
nor U2349 (N_2349,N_2231,N_2298);
or U2350 (N_2350,N_2212,N_2256);
or U2351 (N_2351,N_2265,N_2281);
nand U2352 (N_2352,N_2283,N_2280);
or U2353 (N_2353,N_2211,N_2229);
nor U2354 (N_2354,N_2240,N_2261);
and U2355 (N_2355,N_2264,N_2263);
xnor U2356 (N_2356,N_2227,N_2225);
nor U2357 (N_2357,N_2216,N_2203);
xor U2358 (N_2358,N_2263,N_2260);
nor U2359 (N_2359,N_2255,N_2280);
or U2360 (N_2360,N_2249,N_2246);
or U2361 (N_2361,N_2207,N_2277);
nor U2362 (N_2362,N_2253,N_2244);
and U2363 (N_2363,N_2298,N_2271);
nand U2364 (N_2364,N_2285,N_2296);
xor U2365 (N_2365,N_2266,N_2276);
or U2366 (N_2366,N_2275,N_2260);
nand U2367 (N_2367,N_2244,N_2256);
xor U2368 (N_2368,N_2260,N_2255);
and U2369 (N_2369,N_2202,N_2290);
and U2370 (N_2370,N_2242,N_2293);
nand U2371 (N_2371,N_2230,N_2279);
or U2372 (N_2372,N_2227,N_2213);
nor U2373 (N_2373,N_2215,N_2202);
and U2374 (N_2374,N_2221,N_2265);
nor U2375 (N_2375,N_2296,N_2278);
nand U2376 (N_2376,N_2287,N_2267);
or U2377 (N_2377,N_2232,N_2225);
nand U2378 (N_2378,N_2248,N_2208);
nand U2379 (N_2379,N_2251,N_2263);
nor U2380 (N_2380,N_2219,N_2231);
nor U2381 (N_2381,N_2208,N_2251);
nor U2382 (N_2382,N_2282,N_2230);
nor U2383 (N_2383,N_2209,N_2281);
or U2384 (N_2384,N_2256,N_2228);
nor U2385 (N_2385,N_2235,N_2215);
nor U2386 (N_2386,N_2283,N_2231);
or U2387 (N_2387,N_2298,N_2277);
nand U2388 (N_2388,N_2259,N_2245);
nor U2389 (N_2389,N_2296,N_2272);
xnor U2390 (N_2390,N_2271,N_2281);
and U2391 (N_2391,N_2241,N_2267);
and U2392 (N_2392,N_2238,N_2274);
nand U2393 (N_2393,N_2248,N_2220);
xnor U2394 (N_2394,N_2269,N_2272);
nor U2395 (N_2395,N_2210,N_2214);
nor U2396 (N_2396,N_2293,N_2204);
or U2397 (N_2397,N_2226,N_2293);
and U2398 (N_2398,N_2277,N_2220);
or U2399 (N_2399,N_2283,N_2263);
xor U2400 (N_2400,N_2381,N_2398);
or U2401 (N_2401,N_2310,N_2370);
xnor U2402 (N_2402,N_2323,N_2383);
xor U2403 (N_2403,N_2371,N_2330);
xnor U2404 (N_2404,N_2338,N_2314);
or U2405 (N_2405,N_2311,N_2334);
or U2406 (N_2406,N_2337,N_2374);
xnor U2407 (N_2407,N_2301,N_2300);
or U2408 (N_2408,N_2304,N_2306);
and U2409 (N_2409,N_2339,N_2366);
nor U2410 (N_2410,N_2351,N_2349);
and U2411 (N_2411,N_2358,N_2361);
nand U2412 (N_2412,N_2396,N_2372);
and U2413 (N_2413,N_2364,N_2382);
or U2414 (N_2414,N_2390,N_2319);
nand U2415 (N_2415,N_2332,N_2388);
and U2416 (N_2416,N_2359,N_2375);
or U2417 (N_2417,N_2324,N_2326);
xnor U2418 (N_2418,N_2340,N_2321);
xor U2419 (N_2419,N_2394,N_2336);
and U2420 (N_2420,N_2362,N_2344);
xnor U2421 (N_2421,N_2377,N_2391);
nor U2422 (N_2422,N_2365,N_2328);
nor U2423 (N_2423,N_2353,N_2376);
nand U2424 (N_2424,N_2352,N_2385);
or U2425 (N_2425,N_2354,N_2393);
nand U2426 (N_2426,N_2342,N_2395);
nand U2427 (N_2427,N_2333,N_2303);
nand U2428 (N_2428,N_2348,N_2360);
nor U2429 (N_2429,N_2302,N_2331);
xnor U2430 (N_2430,N_2350,N_2343);
or U2431 (N_2431,N_2315,N_2346);
nand U2432 (N_2432,N_2378,N_2368);
and U2433 (N_2433,N_2345,N_2355);
xnor U2434 (N_2434,N_2308,N_2399);
nand U2435 (N_2435,N_2318,N_2387);
xor U2436 (N_2436,N_2329,N_2312);
nand U2437 (N_2437,N_2389,N_2325);
xnor U2438 (N_2438,N_2357,N_2320);
and U2439 (N_2439,N_2317,N_2384);
and U2440 (N_2440,N_2307,N_2363);
and U2441 (N_2441,N_2341,N_2386);
nand U2442 (N_2442,N_2367,N_2373);
xnor U2443 (N_2443,N_2327,N_2347);
xor U2444 (N_2444,N_2309,N_2322);
or U2445 (N_2445,N_2380,N_2313);
nand U2446 (N_2446,N_2397,N_2335);
xnor U2447 (N_2447,N_2379,N_2356);
nor U2448 (N_2448,N_2316,N_2305);
or U2449 (N_2449,N_2369,N_2392);
nor U2450 (N_2450,N_2366,N_2318);
and U2451 (N_2451,N_2360,N_2359);
and U2452 (N_2452,N_2344,N_2373);
or U2453 (N_2453,N_2361,N_2337);
nor U2454 (N_2454,N_2350,N_2372);
nor U2455 (N_2455,N_2332,N_2355);
nor U2456 (N_2456,N_2327,N_2348);
or U2457 (N_2457,N_2340,N_2359);
nor U2458 (N_2458,N_2396,N_2325);
nor U2459 (N_2459,N_2352,N_2370);
and U2460 (N_2460,N_2352,N_2357);
xnor U2461 (N_2461,N_2328,N_2371);
nand U2462 (N_2462,N_2384,N_2372);
and U2463 (N_2463,N_2304,N_2362);
and U2464 (N_2464,N_2389,N_2388);
or U2465 (N_2465,N_2384,N_2301);
or U2466 (N_2466,N_2336,N_2346);
xnor U2467 (N_2467,N_2310,N_2317);
nand U2468 (N_2468,N_2321,N_2354);
or U2469 (N_2469,N_2398,N_2316);
or U2470 (N_2470,N_2338,N_2343);
nand U2471 (N_2471,N_2336,N_2390);
or U2472 (N_2472,N_2324,N_2317);
nand U2473 (N_2473,N_2328,N_2325);
or U2474 (N_2474,N_2329,N_2310);
or U2475 (N_2475,N_2376,N_2308);
xnor U2476 (N_2476,N_2372,N_2316);
and U2477 (N_2477,N_2343,N_2325);
nor U2478 (N_2478,N_2348,N_2325);
nor U2479 (N_2479,N_2349,N_2311);
and U2480 (N_2480,N_2350,N_2326);
and U2481 (N_2481,N_2336,N_2387);
or U2482 (N_2482,N_2304,N_2331);
or U2483 (N_2483,N_2377,N_2321);
or U2484 (N_2484,N_2370,N_2323);
nor U2485 (N_2485,N_2325,N_2369);
nor U2486 (N_2486,N_2383,N_2382);
nor U2487 (N_2487,N_2387,N_2366);
xor U2488 (N_2488,N_2318,N_2344);
nand U2489 (N_2489,N_2357,N_2317);
and U2490 (N_2490,N_2323,N_2307);
xnor U2491 (N_2491,N_2361,N_2344);
and U2492 (N_2492,N_2364,N_2371);
and U2493 (N_2493,N_2387,N_2330);
or U2494 (N_2494,N_2325,N_2319);
and U2495 (N_2495,N_2314,N_2367);
nor U2496 (N_2496,N_2366,N_2394);
nor U2497 (N_2497,N_2368,N_2352);
or U2498 (N_2498,N_2334,N_2345);
xor U2499 (N_2499,N_2364,N_2317);
and U2500 (N_2500,N_2418,N_2499);
and U2501 (N_2501,N_2425,N_2464);
and U2502 (N_2502,N_2470,N_2438);
nor U2503 (N_2503,N_2431,N_2454);
nor U2504 (N_2504,N_2463,N_2440);
nor U2505 (N_2505,N_2401,N_2403);
or U2506 (N_2506,N_2430,N_2483);
and U2507 (N_2507,N_2486,N_2495);
xnor U2508 (N_2508,N_2490,N_2406);
xnor U2509 (N_2509,N_2402,N_2481);
xnor U2510 (N_2510,N_2409,N_2459);
nor U2511 (N_2511,N_2484,N_2492);
or U2512 (N_2512,N_2426,N_2491);
nor U2513 (N_2513,N_2493,N_2445);
nor U2514 (N_2514,N_2439,N_2479);
nand U2515 (N_2515,N_2443,N_2434);
nor U2516 (N_2516,N_2482,N_2478);
and U2517 (N_2517,N_2480,N_2474);
and U2518 (N_2518,N_2457,N_2460);
or U2519 (N_2519,N_2451,N_2417);
or U2520 (N_2520,N_2442,N_2407);
xnor U2521 (N_2521,N_2436,N_2446);
or U2522 (N_2522,N_2476,N_2410);
nor U2523 (N_2523,N_2496,N_2461);
nor U2524 (N_2524,N_2494,N_2413);
or U2525 (N_2525,N_2404,N_2412);
or U2526 (N_2526,N_2458,N_2477);
or U2527 (N_2527,N_2466,N_2424);
and U2528 (N_2528,N_2419,N_2468);
nand U2529 (N_2529,N_2415,N_2455);
nand U2530 (N_2530,N_2465,N_2467);
nand U2531 (N_2531,N_2400,N_2449);
nor U2532 (N_2532,N_2456,N_2473);
nor U2533 (N_2533,N_2414,N_2472);
or U2534 (N_2534,N_2444,N_2469);
nor U2535 (N_2535,N_2447,N_2450);
nand U2536 (N_2536,N_2433,N_2497);
and U2537 (N_2537,N_2421,N_2441);
and U2538 (N_2538,N_2475,N_2448);
and U2539 (N_2539,N_2498,N_2452);
xnor U2540 (N_2540,N_2462,N_2429);
nor U2541 (N_2541,N_2453,N_2428);
nor U2542 (N_2542,N_2423,N_2487);
xor U2543 (N_2543,N_2427,N_2411);
and U2544 (N_2544,N_2420,N_2435);
and U2545 (N_2545,N_2416,N_2422);
nor U2546 (N_2546,N_2471,N_2488);
or U2547 (N_2547,N_2432,N_2405);
nor U2548 (N_2548,N_2489,N_2485);
and U2549 (N_2549,N_2437,N_2408);
xnor U2550 (N_2550,N_2469,N_2453);
nor U2551 (N_2551,N_2425,N_2417);
and U2552 (N_2552,N_2495,N_2480);
or U2553 (N_2553,N_2418,N_2415);
nor U2554 (N_2554,N_2400,N_2408);
and U2555 (N_2555,N_2446,N_2460);
nor U2556 (N_2556,N_2472,N_2485);
xor U2557 (N_2557,N_2486,N_2425);
nand U2558 (N_2558,N_2432,N_2434);
or U2559 (N_2559,N_2449,N_2417);
nor U2560 (N_2560,N_2407,N_2477);
and U2561 (N_2561,N_2449,N_2433);
or U2562 (N_2562,N_2475,N_2479);
and U2563 (N_2563,N_2456,N_2406);
nor U2564 (N_2564,N_2480,N_2461);
nand U2565 (N_2565,N_2419,N_2453);
and U2566 (N_2566,N_2421,N_2423);
nor U2567 (N_2567,N_2469,N_2460);
nand U2568 (N_2568,N_2475,N_2404);
or U2569 (N_2569,N_2474,N_2439);
and U2570 (N_2570,N_2480,N_2454);
xnor U2571 (N_2571,N_2418,N_2442);
nand U2572 (N_2572,N_2490,N_2408);
nand U2573 (N_2573,N_2434,N_2469);
or U2574 (N_2574,N_2413,N_2447);
and U2575 (N_2575,N_2470,N_2409);
nand U2576 (N_2576,N_2464,N_2456);
nand U2577 (N_2577,N_2416,N_2424);
xor U2578 (N_2578,N_2441,N_2426);
and U2579 (N_2579,N_2473,N_2422);
xnor U2580 (N_2580,N_2458,N_2496);
and U2581 (N_2581,N_2436,N_2413);
nor U2582 (N_2582,N_2406,N_2442);
and U2583 (N_2583,N_2454,N_2464);
nand U2584 (N_2584,N_2428,N_2436);
xor U2585 (N_2585,N_2470,N_2460);
or U2586 (N_2586,N_2432,N_2420);
and U2587 (N_2587,N_2435,N_2411);
xor U2588 (N_2588,N_2407,N_2488);
nand U2589 (N_2589,N_2411,N_2499);
xnor U2590 (N_2590,N_2402,N_2457);
nand U2591 (N_2591,N_2445,N_2465);
or U2592 (N_2592,N_2449,N_2414);
and U2593 (N_2593,N_2499,N_2434);
xnor U2594 (N_2594,N_2450,N_2415);
or U2595 (N_2595,N_2403,N_2447);
nand U2596 (N_2596,N_2413,N_2475);
nor U2597 (N_2597,N_2491,N_2479);
xor U2598 (N_2598,N_2482,N_2460);
nor U2599 (N_2599,N_2457,N_2465);
nor U2600 (N_2600,N_2549,N_2528);
xor U2601 (N_2601,N_2529,N_2500);
and U2602 (N_2602,N_2540,N_2592);
or U2603 (N_2603,N_2579,N_2565);
nor U2604 (N_2604,N_2596,N_2580);
xor U2605 (N_2605,N_2576,N_2577);
and U2606 (N_2606,N_2575,N_2511);
nand U2607 (N_2607,N_2570,N_2557);
and U2608 (N_2608,N_2525,N_2587);
and U2609 (N_2609,N_2534,N_2518);
nor U2610 (N_2610,N_2526,N_2585);
or U2611 (N_2611,N_2555,N_2550);
nand U2612 (N_2612,N_2598,N_2584);
and U2613 (N_2613,N_2507,N_2535);
nand U2614 (N_2614,N_2501,N_2546);
or U2615 (N_2615,N_2543,N_2566);
nand U2616 (N_2616,N_2508,N_2553);
xor U2617 (N_2617,N_2586,N_2504);
or U2618 (N_2618,N_2520,N_2531);
xor U2619 (N_2619,N_2561,N_2522);
or U2620 (N_2620,N_2558,N_2593);
xnor U2621 (N_2621,N_2527,N_2512);
and U2622 (N_2622,N_2533,N_2559);
nand U2623 (N_2623,N_2541,N_2505);
nor U2624 (N_2624,N_2524,N_2560);
or U2625 (N_2625,N_2530,N_2573);
nand U2626 (N_2626,N_2556,N_2510);
and U2627 (N_2627,N_2581,N_2538);
nor U2628 (N_2628,N_2551,N_2572);
or U2629 (N_2629,N_2554,N_2506);
xnor U2630 (N_2630,N_2599,N_2502);
xnor U2631 (N_2631,N_2563,N_2578);
xnor U2632 (N_2632,N_2583,N_2545);
nor U2633 (N_2633,N_2571,N_2532);
or U2634 (N_2634,N_2536,N_2513);
or U2635 (N_2635,N_2547,N_2537);
xnor U2636 (N_2636,N_2568,N_2567);
nor U2637 (N_2637,N_2509,N_2552);
nand U2638 (N_2638,N_2594,N_2515);
nand U2639 (N_2639,N_2539,N_2595);
nand U2640 (N_2640,N_2523,N_2517);
nand U2641 (N_2641,N_2588,N_2544);
nor U2642 (N_2642,N_2574,N_2503);
nand U2643 (N_2643,N_2589,N_2562);
xor U2644 (N_2644,N_2519,N_2514);
and U2645 (N_2645,N_2591,N_2569);
nand U2646 (N_2646,N_2564,N_2542);
or U2647 (N_2647,N_2548,N_2590);
nor U2648 (N_2648,N_2521,N_2597);
xnor U2649 (N_2649,N_2582,N_2516);
or U2650 (N_2650,N_2564,N_2551);
nand U2651 (N_2651,N_2544,N_2543);
nor U2652 (N_2652,N_2518,N_2557);
or U2653 (N_2653,N_2532,N_2579);
xor U2654 (N_2654,N_2519,N_2543);
xnor U2655 (N_2655,N_2583,N_2538);
nand U2656 (N_2656,N_2508,N_2541);
or U2657 (N_2657,N_2574,N_2592);
and U2658 (N_2658,N_2531,N_2541);
or U2659 (N_2659,N_2567,N_2545);
xor U2660 (N_2660,N_2523,N_2556);
or U2661 (N_2661,N_2567,N_2520);
and U2662 (N_2662,N_2552,N_2550);
xnor U2663 (N_2663,N_2522,N_2506);
nand U2664 (N_2664,N_2551,N_2571);
or U2665 (N_2665,N_2588,N_2561);
nand U2666 (N_2666,N_2540,N_2595);
and U2667 (N_2667,N_2522,N_2503);
or U2668 (N_2668,N_2505,N_2531);
xor U2669 (N_2669,N_2502,N_2588);
nor U2670 (N_2670,N_2530,N_2521);
and U2671 (N_2671,N_2561,N_2546);
nor U2672 (N_2672,N_2579,N_2530);
or U2673 (N_2673,N_2594,N_2527);
or U2674 (N_2674,N_2583,N_2530);
or U2675 (N_2675,N_2559,N_2534);
or U2676 (N_2676,N_2513,N_2520);
nand U2677 (N_2677,N_2503,N_2576);
or U2678 (N_2678,N_2551,N_2518);
nand U2679 (N_2679,N_2507,N_2530);
nand U2680 (N_2680,N_2545,N_2586);
xnor U2681 (N_2681,N_2527,N_2546);
or U2682 (N_2682,N_2527,N_2511);
nand U2683 (N_2683,N_2585,N_2564);
nor U2684 (N_2684,N_2596,N_2531);
and U2685 (N_2685,N_2542,N_2514);
and U2686 (N_2686,N_2587,N_2590);
and U2687 (N_2687,N_2503,N_2533);
and U2688 (N_2688,N_2532,N_2504);
and U2689 (N_2689,N_2514,N_2595);
xnor U2690 (N_2690,N_2518,N_2581);
nor U2691 (N_2691,N_2510,N_2572);
nand U2692 (N_2692,N_2537,N_2578);
and U2693 (N_2693,N_2541,N_2534);
nand U2694 (N_2694,N_2590,N_2592);
nand U2695 (N_2695,N_2515,N_2551);
nor U2696 (N_2696,N_2500,N_2580);
or U2697 (N_2697,N_2506,N_2532);
nand U2698 (N_2698,N_2571,N_2567);
xnor U2699 (N_2699,N_2552,N_2561);
and U2700 (N_2700,N_2621,N_2671);
and U2701 (N_2701,N_2643,N_2633);
nand U2702 (N_2702,N_2661,N_2696);
xnor U2703 (N_2703,N_2601,N_2686);
nand U2704 (N_2704,N_2650,N_2611);
and U2705 (N_2705,N_2695,N_2646);
nor U2706 (N_2706,N_2682,N_2697);
nor U2707 (N_2707,N_2683,N_2612);
nor U2708 (N_2708,N_2631,N_2634);
nand U2709 (N_2709,N_2622,N_2692);
or U2710 (N_2710,N_2641,N_2654);
xor U2711 (N_2711,N_2609,N_2664);
nor U2712 (N_2712,N_2613,N_2626);
nor U2713 (N_2713,N_2665,N_2666);
xor U2714 (N_2714,N_2603,N_2647);
or U2715 (N_2715,N_2606,N_2657);
or U2716 (N_2716,N_2673,N_2649);
or U2717 (N_2717,N_2645,N_2652);
and U2718 (N_2718,N_2639,N_2659);
nand U2719 (N_2719,N_2685,N_2675);
or U2720 (N_2720,N_2687,N_2615);
xnor U2721 (N_2721,N_2637,N_2674);
nand U2722 (N_2722,N_2630,N_2668);
nor U2723 (N_2723,N_2623,N_2635);
nor U2724 (N_2724,N_2690,N_2699);
nor U2725 (N_2725,N_2644,N_2619);
or U2726 (N_2726,N_2655,N_2614);
xnor U2727 (N_2727,N_2625,N_2669);
xor U2728 (N_2728,N_2693,N_2604);
nand U2729 (N_2729,N_2632,N_2627);
or U2730 (N_2730,N_2653,N_2670);
and U2731 (N_2731,N_2642,N_2617);
and U2732 (N_2732,N_2607,N_2676);
xnor U2733 (N_2733,N_2698,N_2629);
nand U2734 (N_2734,N_2648,N_2663);
xor U2735 (N_2735,N_2624,N_2678);
and U2736 (N_2736,N_2684,N_2672);
nand U2737 (N_2737,N_2681,N_2616);
nand U2738 (N_2738,N_2636,N_2600);
or U2739 (N_2739,N_2688,N_2628);
and U2740 (N_2740,N_2660,N_2605);
nor U2741 (N_2741,N_2608,N_2620);
and U2742 (N_2742,N_2610,N_2638);
xor U2743 (N_2743,N_2694,N_2602);
or U2744 (N_2744,N_2691,N_2667);
and U2745 (N_2745,N_2662,N_2651);
xnor U2746 (N_2746,N_2658,N_2640);
nand U2747 (N_2747,N_2680,N_2689);
xnor U2748 (N_2748,N_2677,N_2618);
xor U2749 (N_2749,N_2656,N_2679);
xnor U2750 (N_2750,N_2626,N_2645);
or U2751 (N_2751,N_2620,N_2607);
and U2752 (N_2752,N_2631,N_2649);
nor U2753 (N_2753,N_2663,N_2612);
or U2754 (N_2754,N_2675,N_2608);
nor U2755 (N_2755,N_2683,N_2634);
xor U2756 (N_2756,N_2600,N_2622);
nor U2757 (N_2757,N_2627,N_2691);
nand U2758 (N_2758,N_2639,N_2644);
and U2759 (N_2759,N_2693,N_2641);
nand U2760 (N_2760,N_2618,N_2626);
xnor U2761 (N_2761,N_2667,N_2658);
xor U2762 (N_2762,N_2674,N_2683);
or U2763 (N_2763,N_2637,N_2687);
and U2764 (N_2764,N_2660,N_2613);
nor U2765 (N_2765,N_2641,N_2666);
and U2766 (N_2766,N_2619,N_2606);
and U2767 (N_2767,N_2668,N_2601);
or U2768 (N_2768,N_2695,N_2620);
and U2769 (N_2769,N_2685,N_2630);
xnor U2770 (N_2770,N_2651,N_2642);
xor U2771 (N_2771,N_2685,N_2646);
nand U2772 (N_2772,N_2657,N_2665);
and U2773 (N_2773,N_2635,N_2659);
or U2774 (N_2774,N_2601,N_2627);
and U2775 (N_2775,N_2641,N_2628);
or U2776 (N_2776,N_2629,N_2690);
nand U2777 (N_2777,N_2697,N_2646);
nand U2778 (N_2778,N_2672,N_2636);
nand U2779 (N_2779,N_2679,N_2657);
nor U2780 (N_2780,N_2627,N_2638);
xnor U2781 (N_2781,N_2661,N_2644);
or U2782 (N_2782,N_2624,N_2660);
xnor U2783 (N_2783,N_2695,N_2654);
nand U2784 (N_2784,N_2640,N_2612);
nand U2785 (N_2785,N_2673,N_2645);
nand U2786 (N_2786,N_2636,N_2601);
and U2787 (N_2787,N_2697,N_2698);
nand U2788 (N_2788,N_2610,N_2647);
nand U2789 (N_2789,N_2620,N_2606);
nand U2790 (N_2790,N_2613,N_2698);
and U2791 (N_2791,N_2677,N_2600);
or U2792 (N_2792,N_2614,N_2683);
or U2793 (N_2793,N_2649,N_2667);
nor U2794 (N_2794,N_2675,N_2657);
nor U2795 (N_2795,N_2649,N_2640);
nor U2796 (N_2796,N_2625,N_2631);
nor U2797 (N_2797,N_2640,N_2609);
or U2798 (N_2798,N_2669,N_2697);
xor U2799 (N_2799,N_2619,N_2623);
xnor U2800 (N_2800,N_2717,N_2781);
and U2801 (N_2801,N_2775,N_2746);
nor U2802 (N_2802,N_2701,N_2785);
nand U2803 (N_2803,N_2723,N_2733);
or U2804 (N_2804,N_2742,N_2727);
nand U2805 (N_2805,N_2764,N_2729);
nor U2806 (N_2806,N_2783,N_2740);
xnor U2807 (N_2807,N_2745,N_2782);
and U2808 (N_2808,N_2730,N_2731);
nand U2809 (N_2809,N_2721,N_2744);
nand U2810 (N_2810,N_2741,N_2798);
nor U2811 (N_2811,N_2765,N_2702);
and U2812 (N_2812,N_2753,N_2708);
xor U2813 (N_2813,N_2790,N_2712);
and U2814 (N_2814,N_2734,N_2704);
xnor U2815 (N_2815,N_2786,N_2794);
and U2816 (N_2816,N_2725,N_2792);
or U2817 (N_2817,N_2766,N_2787);
or U2818 (N_2818,N_2796,N_2749);
or U2819 (N_2819,N_2700,N_2750);
xnor U2820 (N_2820,N_2738,N_2779);
nor U2821 (N_2821,N_2706,N_2703);
and U2822 (N_2822,N_2716,N_2732);
or U2823 (N_2823,N_2793,N_2780);
or U2824 (N_2824,N_2756,N_2743);
xnor U2825 (N_2825,N_2713,N_2791);
nor U2826 (N_2826,N_2719,N_2707);
xor U2827 (N_2827,N_2736,N_2772);
and U2828 (N_2828,N_2771,N_2748);
nand U2829 (N_2829,N_2776,N_2751);
xor U2830 (N_2830,N_2760,N_2795);
nand U2831 (N_2831,N_2797,N_2768);
and U2832 (N_2832,N_2763,N_2770);
nand U2833 (N_2833,N_2715,N_2755);
xnor U2834 (N_2834,N_2784,N_2774);
nor U2835 (N_2835,N_2758,N_2752);
xor U2836 (N_2836,N_2767,N_2722);
and U2837 (N_2837,N_2777,N_2711);
xor U2838 (N_2838,N_2778,N_2799);
and U2839 (N_2839,N_2759,N_2773);
nor U2840 (N_2840,N_2718,N_2757);
nand U2841 (N_2841,N_2747,N_2789);
and U2842 (N_2842,N_2769,N_2728);
and U2843 (N_2843,N_2720,N_2754);
nor U2844 (N_2844,N_2739,N_2726);
and U2845 (N_2845,N_2788,N_2735);
and U2846 (N_2846,N_2737,N_2709);
nor U2847 (N_2847,N_2710,N_2724);
and U2848 (N_2848,N_2705,N_2762);
xor U2849 (N_2849,N_2761,N_2714);
nand U2850 (N_2850,N_2757,N_2756);
xnor U2851 (N_2851,N_2780,N_2782);
nor U2852 (N_2852,N_2774,N_2720);
nor U2853 (N_2853,N_2754,N_2768);
or U2854 (N_2854,N_2714,N_2713);
nor U2855 (N_2855,N_2718,N_2708);
xor U2856 (N_2856,N_2766,N_2713);
nand U2857 (N_2857,N_2725,N_2786);
nor U2858 (N_2858,N_2769,N_2755);
xnor U2859 (N_2859,N_2726,N_2794);
and U2860 (N_2860,N_2764,N_2792);
xor U2861 (N_2861,N_2784,N_2792);
and U2862 (N_2862,N_2768,N_2732);
nand U2863 (N_2863,N_2731,N_2732);
and U2864 (N_2864,N_2776,N_2731);
xnor U2865 (N_2865,N_2794,N_2759);
and U2866 (N_2866,N_2756,N_2733);
nand U2867 (N_2867,N_2708,N_2701);
and U2868 (N_2868,N_2729,N_2776);
xnor U2869 (N_2869,N_2713,N_2755);
xnor U2870 (N_2870,N_2743,N_2769);
nor U2871 (N_2871,N_2763,N_2726);
and U2872 (N_2872,N_2757,N_2749);
nand U2873 (N_2873,N_2767,N_2781);
and U2874 (N_2874,N_2715,N_2786);
nor U2875 (N_2875,N_2783,N_2785);
or U2876 (N_2876,N_2723,N_2777);
or U2877 (N_2877,N_2739,N_2701);
and U2878 (N_2878,N_2789,N_2765);
nand U2879 (N_2879,N_2784,N_2714);
or U2880 (N_2880,N_2752,N_2763);
and U2881 (N_2881,N_2776,N_2726);
or U2882 (N_2882,N_2752,N_2719);
or U2883 (N_2883,N_2792,N_2772);
xnor U2884 (N_2884,N_2716,N_2755);
or U2885 (N_2885,N_2725,N_2744);
or U2886 (N_2886,N_2720,N_2700);
nand U2887 (N_2887,N_2735,N_2720);
or U2888 (N_2888,N_2718,N_2734);
nor U2889 (N_2889,N_2737,N_2725);
xnor U2890 (N_2890,N_2781,N_2748);
nor U2891 (N_2891,N_2712,N_2717);
and U2892 (N_2892,N_2727,N_2708);
xnor U2893 (N_2893,N_2787,N_2724);
nand U2894 (N_2894,N_2733,N_2725);
nand U2895 (N_2895,N_2799,N_2755);
nand U2896 (N_2896,N_2798,N_2725);
nor U2897 (N_2897,N_2747,N_2778);
nand U2898 (N_2898,N_2723,N_2757);
nand U2899 (N_2899,N_2714,N_2742);
xor U2900 (N_2900,N_2871,N_2898);
or U2901 (N_2901,N_2834,N_2884);
xor U2902 (N_2902,N_2823,N_2864);
nand U2903 (N_2903,N_2868,N_2882);
xor U2904 (N_2904,N_2873,N_2812);
xnor U2905 (N_2905,N_2804,N_2839);
xnor U2906 (N_2906,N_2822,N_2851);
xor U2907 (N_2907,N_2832,N_2805);
nor U2908 (N_2908,N_2880,N_2821);
nor U2909 (N_2909,N_2887,N_2820);
nor U2910 (N_2910,N_2856,N_2876);
and U2911 (N_2911,N_2843,N_2815);
and U2912 (N_2912,N_2866,N_2886);
and U2913 (N_2913,N_2848,N_2850);
or U2914 (N_2914,N_2826,N_2810);
nand U2915 (N_2915,N_2829,N_2867);
or U2916 (N_2916,N_2814,N_2831);
or U2917 (N_2917,N_2803,N_2806);
xnor U2918 (N_2918,N_2893,N_2807);
and U2919 (N_2919,N_2860,N_2895);
xor U2920 (N_2920,N_2837,N_2863);
and U2921 (N_2921,N_2828,N_2842);
or U2922 (N_2922,N_2801,N_2870);
nand U2923 (N_2923,N_2889,N_2872);
nor U2924 (N_2924,N_2827,N_2878);
or U2925 (N_2925,N_2855,N_2836);
nor U2926 (N_2926,N_2835,N_2859);
xor U2927 (N_2927,N_2845,N_2858);
nand U2928 (N_2928,N_2841,N_2890);
nor U2929 (N_2929,N_2809,N_2847);
xor U2930 (N_2930,N_2877,N_2857);
nand U2931 (N_2931,N_2865,N_2833);
or U2932 (N_2932,N_2830,N_2802);
and U2933 (N_2933,N_2800,N_2816);
nand U2934 (N_2934,N_2817,N_2818);
and U2935 (N_2935,N_2853,N_2896);
nor U2936 (N_2936,N_2892,N_2825);
nor U2937 (N_2937,N_2846,N_2838);
xor U2938 (N_2938,N_2844,N_2808);
xor U2939 (N_2939,N_2862,N_2861);
nand U2940 (N_2940,N_2824,N_2891);
or U2941 (N_2941,N_2894,N_2854);
xnor U2942 (N_2942,N_2813,N_2849);
and U2943 (N_2943,N_2840,N_2879);
nand U2944 (N_2944,N_2875,N_2852);
and U2945 (N_2945,N_2869,N_2811);
nand U2946 (N_2946,N_2881,N_2897);
and U2947 (N_2947,N_2888,N_2874);
nand U2948 (N_2948,N_2883,N_2885);
xor U2949 (N_2949,N_2899,N_2819);
nand U2950 (N_2950,N_2800,N_2834);
nor U2951 (N_2951,N_2816,N_2866);
xnor U2952 (N_2952,N_2871,N_2836);
nand U2953 (N_2953,N_2890,N_2842);
xnor U2954 (N_2954,N_2872,N_2881);
nor U2955 (N_2955,N_2853,N_2801);
xnor U2956 (N_2956,N_2838,N_2832);
xor U2957 (N_2957,N_2823,N_2844);
nor U2958 (N_2958,N_2876,N_2846);
nor U2959 (N_2959,N_2883,N_2884);
or U2960 (N_2960,N_2850,N_2835);
nand U2961 (N_2961,N_2813,N_2874);
xnor U2962 (N_2962,N_2807,N_2888);
xor U2963 (N_2963,N_2891,N_2808);
nand U2964 (N_2964,N_2840,N_2800);
or U2965 (N_2965,N_2835,N_2870);
or U2966 (N_2966,N_2813,N_2810);
or U2967 (N_2967,N_2805,N_2874);
nand U2968 (N_2968,N_2823,N_2880);
nand U2969 (N_2969,N_2852,N_2838);
xor U2970 (N_2970,N_2875,N_2899);
and U2971 (N_2971,N_2861,N_2827);
and U2972 (N_2972,N_2810,N_2832);
nor U2973 (N_2973,N_2852,N_2832);
xnor U2974 (N_2974,N_2811,N_2848);
xor U2975 (N_2975,N_2833,N_2888);
nor U2976 (N_2976,N_2841,N_2849);
or U2977 (N_2977,N_2811,N_2818);
nor U2978 (N_2978,N_2800,N_2849);
and U2979 (N_2979,N_2829,N_2872);
nand U2980 (N_2980,N_2865,N_2876);
and U2981 (N_2981,N_2830,N_2836);
and U2982 (N_2982,N_2855,N_2840);
or U2983 (N_2983,N_2815,N_2818);
nand U2984 (N_2984,N_2839,N_2864);
xor U2985 (N_2985,N_2854,N_2852);
and U2986 (N_2986,N_2889,N_2812);
nor U2987 (N_2987,N_2863,N_2892);
nand U2988 (N_2988,N_2838,N_2874);
nor U2989 (N_2989,N_2883,N_2889);
and U2990 (N_2990,N_2836,N_2872);
nor U2991 (N_2991,N_2856,N_2877);
nand U2992 (N_2992,N_2872,N_2833);
nand U2993 (N_2993,N_2882,N_2803);
nor U2994 (N_2994,N_2887,N_2890);
and U2995 (N_2995,N_2851,N_2887);
and U2996 (N_2996,N_2819,N_2801);
and U2997 (N_2997,N_2897,N_2804);
and U2998 (N_2998,N_2878,N_2852);
nor U2999 (N_2999,N_2841,N_2876);
nor U3000 (N_3000,N_2983,N_2971);
xor U3001 (N_3001,N_2914,N_2936);
nand U3002 (N_3002,N_2968,N_2980);
and U3003 (N_3003,N_2950,N_2935);
or U3004 (N_3004,N_2966,N_2939);
or U3005 (N_3005,N_2910,N_2996);
and U3006 (N_3006,N_2972,N_2969);
xnor U3007 (N_3007,N_2981,N_2930);
or U3008 (N_3008,N_2997,N_2940);
nor U3009 (N_3009,N_2962,N_2961);
nand U3010 (N_3010,N_2982,N_2989);
xnor U3011 (N_3011,N_2959,N_2913);
nand U3012 (N_3012,N_2988,N_2919);
xor U3013 (N_3013,N_2998,N_2922);
xnor U3014 (N_3014,N_2976,N_2958);
nor U3015 (N_3015,N_2916,N_2986);
and U3016 (N_3016,N_2975,N_2956);
nor U3017 (N_3017,N_2993,N_2990);
or U3018 (N_3018,N_2925,N_2991);
xnor U3019 (N_3019,N_2960,N_2943);
xnor U3020 (N_3020,N_2946,N_2915);
nand U3021 (N_3021,N_2955,N_2924);
or U3022 (N_3022,N_2907,N_2953);
nand U3023 (N_3023,N_2906,N_2964);
xor U3024 (N_3024,N_2949,N_2920);
nor U3025 (N_3025,N_2992,N_2909);
xnor U3026 (N_3026,N_2951,N_2932);
or U3027 (N_3027,N_2923,N_2902);
nand U3028 (N_3028,N_2933,N_2984);
nand U3029 (N_3029,N_2908,N_2900);
xnor U3030 (N_3030,N_2974,N_2965);
nand U3031 (N_3031,N_2921,N_2903);
xnor U3032 (N_3032,N_2937,N_2954);
and U3033 (N_3033,N_2947,N_2978);
nand U3034 (N_3034,N_2905,N_2917);
nand U3035 (N_3035,N_2941,N_2963);
xnor U3036 (N_3036,N_2918,N_2928);
and U3037 (N_3037,N_2979,N_2926);
and U3038 (N_3038,N_2994,N_2970);
xor U3039 (N_3039,N_2938,N_2973);
and U3040 (N_3040,N_2967,N_2952);
nor U3041 (N_3041,N_2944,N_2934);
and U3042 (N_3042,N_2977,N_2985);
or U3043 (N_3043,N_2987,N_2912);
xor U3044 (N_3044,N_2904,N_2929);
nor U3045 (N_3045,N_2927,N_2942);
or U3046 (N_3046,N_2945,N_2911);
nor U3047 (N_3047,N_2948,N_2957);
nand U3048 (N_3048,N_2995,N_2999);
nand U3049 (N_3049,N_2931,N_2901);
or U3050 (N_3050,N_2946,N_2934);
xor U3051 (N_3051,N_2985,N_2908);
xor U3052 (N_3052,N_2967,N_2997);
xor U3053 (N_3053,N_2944,N_2954);
xor U3054 (N_3054,N_2946,N_2933);
nor U3055 (N_3055,N_2956,N_2933);
nor U3056 (N_3056,N_2924,N_2986);
xor U3057 (N_3057,N_2947,N_2966);
or U3058 (N_3058,N_2934,N_2941);
nor U3059 (N_3059,N_2976,N_2907);
or U3060 (N_3060,N_2926,N_2958);
xnor U3061 (N_3061,N_2945,N_2931);
and U3062 (N_3062,N_2933,N_2925);
and U3063 (N_3063,N_2995,N_2996);
xnor U3064 (N_3064,N_2912,N_2925);
nand U3065 (N_3065,N_2993,N_2949);
xor U3066 (N_3066,N_2912,N_2970);
and U3067 (N_3067,N_2931,N_2960);
nand U3068 (N_3068,N_2918,N_2960);
nor U3069 (N_3069,N_2908,N_2941);
nand U3070 (N_3070,N_2946,N_2916);
or U3071 (N_3071,N_2914,N_2943);
nor U3072 (N_3072,N_2981,N_2902);
nor U3073 (N_3073,N_2968,N_2963);
or U3074 (N_3074,N_2964,N_2930);
or U3075 (N_3075,N_2900,N_2989);
and U3076 (N_3076,N_2905,N_2956);
nor U3077 (N_3077,N_2900,N_2944);
xnor U3078 (N_3078,N_2919,N_2910);
xnor U3079 (N_3079,N_2984,N_2956);
nor U3080 (N_3080,N_2988,N_2916);
or U3081 (N_3081,N_2907,N_2900);
and U3082 (N_3082,N_2943,N_2966);
nor U3083 (N_3083,N_2958,N_2950);
or U3084 (N_3084,N_2924,N_2937);
or U3085 (N_3085,N_2995,N_2961);
or U3086 (N_3086,N_2984,N_2904);
nand U3087 (N_3087,N_2900,N_2914);
nor U3088 (N_3088,N_2923,N_2981);
nor U3089 (N_3089,N_2917,N_2929);
nor U3090 (N_3090,N_2924,N_2916);
or U3091 (N_3091,N_2949,N_2922);
nor U3092 (N_3092,N_2970,N_2985);
and U3093 (N_3093,N_2913,N_2945);
nand U3094 (N_3094,N_2981,N_2928);
and U3095 (N_3095,N_2993,N_2946);
nand U3096 (N_3096,N_2959,N_2967);
nand U3097 (N_3097,N_2927,N_2934);
nor U3098 (N_3098,N_2985,N_2915);
nand U3099 (N_3099,N_2973,N_2949);
and U3100 (N_3100,N_3010,N_3031);
xor U3101 (N_3101,N_3060,N_3084);
nor U3102 (N_3102,N_3065,N_3059);
nand U3103 (N_3103,N_3082,N_3049);
and U3104 (N_3104,N_3090,N_3055);
xnor U3105 (N_3105,N_3088,N_3089);
xnor U3106 (N_3106,N_3042,N_3014);
and U3107 (N_3107,N_3003,N_3027);
nor U3108 (N_3108,N_3034,N_3095);
or U3109 (N_3109,N_3093,N_3069);
and U3110 (N_3110,N_3085,N_3086);
or U3111 (N_3111,N_3098,N_3036);
and U3112 (N_3112,N_3064,N_3076);
xor U3113 (N_3113,N_3009,N_3061);
nor U3114 (N_3114,N_3015,N_3067);
xor U3115 (N_3115,N_3073,N_3021);
or U3116 (N_3116,N_3025,N_3026);
xnor U3117 (N_3117,N_3006,N_3053);
xnor U3118 (N_3118,N_3081,N_3046);
or U3119 (N_3119,N_3072,N_3063);
or U3120 (N_3120,N_3097,N_3039);
xor U3121 (N_3121,N_3077,N_3017);
or U3122 (N_3122,N_3038,N_3099);
nand U3123 (N_3123,N_3005,N_3080);
xnor U3124 (N_3124,N_3051,N_3040);
and U3125 (N_3125,N_3007,N_3062);
xor U3126 (N_3126,N_3068,N_3087);
xor U3127 (N_3127,N_3008,N_3043);
or U3128 (N_3128,N_3020,N_3048);
nor U3129 (N_3129,N_3092,N_3052);
or U3130 (N_3130,N_3012,N_3058);
nor U3131 (N_3131,N_3030,N_3054);
xnor U3132 (N_3132,N_3070,N_3004);
nor U3133 (N_3133,N_3079,N_3018);
nand U3134 (N_3134,N_3047,N_3032);
xor U3135 (N_3135,N_3001,N_3044);
and U3136 (N_3136,N_3023,N_3050);
and U3137 (N_3137,N_3019,N_3074);
and U3138 (N_3138,N_3013,N_3091);
nand U3139 (N_3139,N_3083,N_3022);
nand U3140 (N_3140,N_3056,N_3066);
xnor U3141 (N_3141,N_3037,N_3029);
xnor U3142 (N_3142,N_3024,N_3041);
nor U3143 (N_3143,N_3000,N_3035);
xnor U3144 (N_3144,N_3057,N_3071);
nand U3145 (N_3145,N_3016,N_3045);
nor U3146 (N_3146,N_3028,N_3002);
nor U3147 (N_3147,N_3033,N_3011);
and U3148 (N_3148,N_3096,N_3075);
nor U3149 (N_3149,N_3094,N_3078);
or U3150 (N_3150,N_3041,N_3031);
or U3151 (N_3151,N_3026,N_3045);
or U3152 (N_3152,N_3019,N_3070);
and U3153 (N_3153,N_3040,N_3005);
xnor U3154 (N_3154,N_3002,N_3007);
nor U3155 (N_3155,N_3070,N_3038);
nand U3156 (N_3156,N_3026,N_3056);
nor U3157 (N_3157,N_3019,N_3033);
or U3158 (N_3158,N_3085,N_3028);
nand U3159 (N_3159,N_3071,N_3080);
or U3160 (N_3160,N_3028,N_3067);
xnor U3161 (N_3161,N_3070,N_3056);
or U3162 (N_3162,N_3053,N_3086);
nand U3163 (N_3163,N_3026,N_3075);
nand U3164 (N_3164,N_3067,N_3063);
and U3165 (N_3165,N_3015,N_3071);
xnor U3166 (N_3166,N_3089,N_3087);
or U3167 (N_3167,N_3045,N_3092);
nor U3168 (N_3168,N_3085,N_3071);
xor U3169 (N_3169,N_3017,N_3018);
or U3170 (N_3170,N_3065,N_3063);
nor U3171 (N_3171,N_3002,N_3067);
or U3172 (N_3172,N_3025,N_3099);
or U3173 (N_3173,N_3077,N_3082);
nand U3174 (N_3174,N_3036,N_3076);
or U3175 (N_3175,N_3057,N_3036);
and U3176 (N_3176,N_3014,N_3004);
or U3177 (N_3177,N_3033,N_3051);
or U3178 (N_3178,N_3058,N_3097);
nor U3179 (N_3179,N_3024,N_3092);
or U3180 (N_3180,N_3021,N_3051);
and U3181 (N_3181,N_3080,N_3036);
or U3182 (N_3182,N_3000,N_3006);
and U3183 (N_3183,N_3078,N_3056);
nand U3184 (N_3184,N_3085,N_3008);
xnor U3185 (N_3185,N_3030,N_3032);
or U3186 (N_3186,N_3001,N_3059);
nor U3187 (N_3187,N_3054,N_3041);
and U3188 (N_3188,N_3063,N_3025);
xor U3189 (N_3189,N_3001,N_3019);
or U3190 (N_3190,N_3048,N_3005);
nor U3191 (N_3191,N_3066,N_3032);
and U3192 (N_3192,N_3046,N_3016);
nand U3193 (N_3193,N_3098,N_3035);
and U3194 (N_3194,N_3008,N_3037);
nor U3195 (N_3195,N_3092,N_3069);
xor U3196 (N_3196,N_3084,N_3001);
xor U3197 (N_3197,N_3000,N_3085);
xor U3198 (N_3198,N_3014,N_3036);
nand U3199 (N_3199,N_3047,N_3080);
and U3200 (N_3200,N_3113,N_3128);
and U3201 (N_3201,N_3122,N_3174);
or U3202 (N_3202,N_3193,N_3183);
and U3203 (N_3203,N_3157,N_3104);
and U3204 (N_3204,N_3196,N_3194);
nor U3205 (N_3205,N_3108,N_3187);
xnor U3206 (N_3206,N_3180,N_3142);
nor U3207 (N_3207,N_3154,N_3125);
nand U3208 (N_3208,N_3135,N_3130);
and U3209 (N_3209,N_3143,N_3117);
nor U3210 (N_3210,N_3153,N_3131);
or U3211 (N_3211,N_3179,N_3163);
nand U3212 (N_3212,N_3132,N_3139);
xor U3213 (N_3213,N_3176,N_3191);
or U3214 (N_3214,N_3171,N_3101);
nor U3215 (N_3215,N_3195,N_3161);
or U3216 (N_3216,N_3146,N_3172);
nor U3217 (N_3217,N_3149,N_3100);
nand U3218 (N_3218,N_3148,N_3141);
nor U3219 (N_3219,N_3133,N_3138);
xnor U3220 (N_3220,N_3119,N_3166);
and U3221 (N_3221,N_3198,N_3160);
nor U3222 (N_3222,N_3144,N_3103);
or U3223 (N_3223,N_3181,N_3134);
nor U3224 (N_3224,N_3184,N_3136);
xor U3225 (N_3225,N_3190,N_3192);
or U3226 (N_3226,N_3121,N_3156);
xor U3227 (N_3227,N_3158,N_3167);
or U3228 (N_3228,N_3123,N_3177);
and U3229 (N_3229,N_3112,N_3169);
nand U3230 (N_3230,N_3151,N_3165);
nand U3231 (N_3231,N_3164,N_3105);
or U3232 (N_3232,N_3175,N_3116);
or U3233 (N_3233,N_3145,N_3168);
nand U3234 (N_3234,N_3162,N_3152);
nand U3235 (N_3235,N_3137,N_3107);
nor U3236 (N_3236,N_3129,N_3147);
or U3237 (N_3237,N_3188,N_3106);
nor U3238 (N_3238,N_3173,N_3185);
nand U3239 (N_3239,N_3189,N_3140);
or U3240 (N_3240,N_3127,N_3102);
xnor U3241 (N_3241,N_3197,N_3109);
xnor U3242 (N_3242,N_3186,N_3178);
and U3243 (N_3243,N_3120,N_3150);
xnor U3244 (N_3244,N_3159,N_3115);
nand U3245 (N_3245,N_3114,N_3118);
or U3246 (N_3246,N_3126,N_3110);
nand U3247 (N_3247,N_3182,N_3199);
xnor U3248 (N_3248,N_3111,N_3124);
xor U3249 (N_3249,N_3170,N_3155);
nor U3250 (N_3250,N_3174,N_3168);
xor U3251 (N_3251,N_3150,N_3184);
nor U3252 (N_3252,N_3126,N_3100);
nor U3253 (N_3253,N_3161,N_3138);
nor U3254 (N_3254,N_3166,N_3183);
nor U3255 (N_3255,N_3113,N_3106);
nor U3256 (N_3256,N_3144,N_3196);
or U3257 (N_3257,N_3196,N_3169);
nor U3258 (N_3258,N_3101,N_3154);
and U3259 (N_3259,N_3111,N_3154);
or U3260 (N_3260,N_3126,N_3144);
nand U3261 (N_3261,N_3198,N_3186);
and U3262 (N_3262,N_3144,N_3198);
nor U3263 (N_3263,N_3130,N_3122);
and U3264 (N_3264,N_3117,N_3179);
xnor U3265 (N_3265,N_3193,N_3114);
nor U3266 (N_3266,N_3110,N_3115);
and U3267 (N_3267,N_3199,N_3106);
xnor U3268 (N_3268,N_3126,N_3179);
nor U3269 (N_3269,N_3170,N_3142);
and U3270 (N_3270,N_3154,N_3107);
nand U3271 (N_3271,N_3164,N_3159);
and U3272 (N_3272,N_3128,N_3174);
xor U3273 (N_3273,N_3136,N_3145);
nor U3274 (N_3274,N_3132,N_3107);
xnor U3275 (N_3275,N_3111,N_3128);
nor U3276 (N_3276,N_3110,N_3117);
or U3277 (N_3277,N_3167,N_3104);
xor U3278 (N_3278,N_3173,N_3187);
or U3279 (N_3279,N_3190,N_3160);
xor U3280 (N_3280,N_3169,N_3176);
nand U3281 (N_3281,N_3117,N_3186);
nand U3282 (N_3282,N_3188,N_3108);
and U3283 (N_3283,N_3150,N_3199);
nor U3284 (N_3284,N_3150,N_3106);
nand U3285 (N_3285,N_3131,N_3137);
and U3286 (N_3286,N_3144,N_3117);
or U3287 (N_3287,N_3134,N_3195);
nor U3288 (N_3288,N_3145,N_3179);
and U3289 (N_3289,N_3152,N_3163);
xnor U3290 (N_3290,N_3139,N_3142);
xnor U3291 (N_3291,N_3119,N_3105);
nor U3292 (N_3292,N_3192,N_3189);
xor U3293 (N_3293,N_3193,N_3171);
and U3294 (N_3294,N_3124,N_3171);
nor U3295 (N_3295,N_3166,N_3153);
nor U3296 (N_3296,N_3103,N_3120);
nor U3297 (N_3297,N_3151,N_3191);
or U3298 (N_3298,N_3142,N_3172);
and U3299 (N_3299,N_3138,N_3153);
nand U3300 (N_3300,N_3258,N_3286);
and U3301 (N_3301,N_3208,N_3227);
nor U3302 (N_3302,N_3216,N_3214);
nor U3303 (N_3303,N_3279,N_3230);
xor U3304 (N_3304,N_3201,N_3296);
xor U3305 (N_3305,N_3231,N_3234);
nand U3306 (N_3306,N_3294,N_3295);
and U3307 (N_3307,N_3259,N_3221);
and U3308 (N_3308,N_3275,N_3285);
and U3309 (N_3309,N_3266,N_3273);
nand U3310 (N_3310,N_3244,N_3284);
and U3311 (N_3311,N_3271,N_3280);
or U3312 (N_3312,N_3270,N_3247);
xnor U3313 (N_3313,N_3240,N_3290);
nor U3314 (N_3314,N_3255,N_3202);
xnor U3315 (N_3315,N_3246,N_3248);
and U3316 (N_3316,N_3281,N_3261);
xnor U3317 (N_3317,N_3241,N_3267);
nand U3318 (N_3318,N_3293,N_3210);
or U3319 (N_3319,N_3222,N_3272);
nand U3320 (N_3320,N_3298,N_3276);
or U3321 (N_3321,N_3238,N_3200);
or U3322 (N_3322,N_3228,N_3289);
xor U3323 (N_3323,N_3209,N_3287);
and U3324 (N_3324,N_3249,N_3262);
or U3325 (N_3325,N_3288,N_3203);
xnor U3326 (N_3326,N_3205,N_3263);
and U3327 (N_3327,N_3204,N_3250);
and U3328 (N_3328,N_3237,N_3235);
or U3329 (N_3329,N_3212,N_3291);
or U3330 (N_3330,N_3233,N_3215);
nand U3331 (N_3331,N_3223,N_3282);
nand U3332 (N_3332,N_3220,N_3232);
and U3333 (N_3333,N_3211,N_3268);
nor U3334 (N_3334,N_3254,N_3219);
nand U3335 (N_3335,N_3283,N_3299);
or U3336 (N_3336,N_3207,N_3260);
and U3337 (N_3337,N_3206,N_3226);
nand U3338 (N_3338,N_3252,N_3253);
and U3339 (N_3339,N_3292,N_3242);
nand U3340 (N_3340,N_3265,N_3251);
xor U3341 (N_3341,N_3256,N_3229);
xnor U3342 (N_3342,N_3236,N_3239);
nor U3343 (N_3343,N_3264,N_3243);
nand U3344 (N_3344,N_3245,N_3218);
xor U3345 (N_3345,N_3274,N_3297);
and U3346 (N_3346,N_3213,N_3225);
and U3347 (N_3347,N_3277,N_3257);
and U3348 (N_3348,N_3224,N_3278);
or U3349 (N_3349,N_3217,N_3269);
nor U3350 (N_3350,N_3258,N_3267);
xnor U3351 (N_3351,N_3223,N_3248);
nand U3352 (N_3352,N_3251,N_3218);
and U3353 (N_3353,N_3266,N_3205);
or U3354 (N_3354,N_3278,N_3279);
nand U3355 (N_3355,N_3239,N_3247);
nor U3356 (N_3356,N_3279,N_3242);
nor U3357 (N_3357,N_3267,N_3233);
or U3358 (N_3358,N_3283,N_3262);
or U3359 (N_3359,N_3228,N_3239);
nor U3360 (N_3360,N_3243,N_3236);
nor U3361 (N_3361,N_3252,N_3237);
nand U3362 (N_3362,N_3239,N_3202);
or U3363 (N_3363,N_3230,N_3228);
nand U3364 (N_3364,N_3256,N_3232);
or U3365 (N_3365,N_3288,N_3280);
and U3366 (N_3366,N_3270,N_3264);
nor U3367 (N_3367,N_3292,N_3279);
nor U3368 (N_3368,N_3210,N_3212);
nand U3369 (N_3369,N_3299,N_3268);
xor U3370 (N_3370,N_3217,N_3249);
nor U3371 (N_3371,N_3213,N_3200);
xor U3372 (N_3372,N_3202,N_3258);
nor U3373 (N_3373,N_3280,N_3222);
nand U3374 (N_3374,N_3231,N_3249);
and U3375 (N_3375,N_3240,N_3247);
and U3376 (N_3376,N_3291,N_3247);
xnor U3377 (N_3377,N_3215,N_3220);
xor U3378 (N_3378,N_3297,N_3209);
nor U3379 (N_3379,N_3209,N_3275);
nor U3380 (N_3380,N_3299,N_3273);
xor U3381 (N_3381,N_3289,N_3233);
or U3382 (N_3382,N_3203,N_3202);
or U3383 (N_3383,N_3280,N_3202);
or U3384 (N_3384,N_3259,N_3255);
nor U3385 (N_3385,N_3263,N_3223);
xor U3386 (N_3386,N_3220,N_3268);
or U3387 (N_3387,N_3277,N_3288);
nand U3388 (N_3388,N_3288,N_3211);
nand U3389 (N_3389,N_3270,N_3210);
xnor U3390 (N_3390,N_3265,N_3222);
nand U3391 (N_3391,N_3254,N_3285);
or U3392 (N_3392,N_3262,N_3220);
nor U3393 (N_3393,N_3200,N_3252);
and U3394 (N_3394,N_3289,N_3291);
and U3395 (N_3395,N_3266,N_3293);
nor U3396 (N_3396,N_3249,N_3265);
nor U3397 (N_3397,N_3245,N_3225);
and U3398 (N_3398,N_3232,N_3251);
xor U3399 (N_3399,N_3250,N_3266);
nand U3400 (N_3400,N_3385,N_3382);
xor U3401 (N_3401,N_3336,N_3386);
nor U3402 (N_3402,N_3313,N_3387);
nand U3403 (N_3403,N_3339,N_3391);
or U3404 (N_3404,N_3384,N_3305);
or U3405 (N_3405,N_3372,N_3357);
and U3406 (N_3406,N_3358,N_3355);
or U3407 (N_3407,N_3300,N_3361);
xnor U3408 (N_3408,N_3379,N_3353);
or U3409 (N_3409,N_3394,N_3397);
nand U3410 (N_3410,N_3389,N_3331);
xnor U3411 (N_3411,N_3332,N_3367);
or U3412 (N_3412,N_3399,N_3359);
or U3413 (N_3413,N_3380,N_3330);
or U3414 (N_3414,N_3375,N_3344);
or U3415 (N_3415,N_3356,N_3388);
nor U3416 (N_3416,N_3341,N_3349);
nor U3417 (N_3417,N_3365,N_3334);
nor U3418 (N_3418,N_3368,N_3396);
nor U3419 (N_3419,N_3369,N_3376);
or U3420 (N_3420,N_3337,N_3310);
nor U3421 (N_3421,N_3304,N_3398);
and U3422 (N_3422,N_3312,N_3316);
nor U3423 (N_3423,N_3302,N_3363);
and U3424 (N_3424,N_3383,N_3350);
xnor U3425 (N_3425,N_3324,N_3333);
or U3426 (N_3426,N_3348,N_3354);
nand U3427 (N_3427,N_3393,N_3343);
nand U3428 (N_3428,N_3314,N_3323);
or U3429 (N_3429,N_3335,N_3346);
nor U3430 (N_3430,N_3390,N_3320);
and U3431 (N_3431,N_3378,N_3395);
nand U3432 (N_3432,N_3362,N_3381);
and U3433 (N_3433,N_3370,N_3328);
or U3434 (N_3434,N_3371,N_3364);
nor U3435 (N_3435,N_3360,N_3329);
nand U3436 (N_3436,N_3366,N_3317);
nand U3437 (N_3437,N_3306,N_3325);
nand U3438 (N_3438,N_3326,N_3318);
nand U3439 (N_3439,N_3347,N_3308);
or U3440 (N_3440,N_3342,N_3352);
xor U3441 (N_3441,N_3340,N_3392);
and U3442 (N_3442,N_3315,N_3377);
or U3443 (N_3443,N_3309,N_3307);
or U3444 (N_3444,N_3345,N_3311);
xor U3445 (N_3445,N_3301,N_3322);
nand U3446 (N_3446,N_3351,N_3303);
or U3447 (N_3447,N_3373,N_3338);
nor U3448 (N_3448,N_3374,N_3319);
or U3449 (N_3449,N_3321,N_3327);
and U3450 (N_3450,N_3319,N_3353);
nand U3451 (N_3451,N_3338,N_3380);
and U3452 (N_3452,N_3315,N_3367);
and U3453 (N_3453,N_3370,N_3312);
or U3454 (N_3454,N_3331,N_3363);
nand U3455 (N_3455,N_3356,N_3347);
or U3456 (N_3456,N_3399,N_3304);
and U3457 (N_3457,N_3359,N_3320);
or U3458 (N_3458,N_3356,N_3312);
xnor U3459 (N_3459,N_3357,N_3352);
or U3460 (N_3460,N_3332,N_3353);
nand U3461 (N_3461,N_3351,N_3318);
and U3462 (N_3462,N_3336,N_3308);
nor U3463 (N_3463,N_3321,N_3372);
or U3464 (N_3464,N_3327,N_3339);
xor U3465 (N_3465,N_3347,N_3351);
and U3466 (N_3466,N_3395,N_3302);
nor U3467 (N_3467,N_3312,N_3390);
nand U3468 (N_3468,N_3331,N_3321);
nor U3469 (N_3469,N_3353,N_3348);
nand U3470 (N_3470,N_3337,N_3327);
or U3471 (N_3471,N_3346,N_3313);
or U3472 (N_3472,N_3331,N_3368);
or U3473 (N_3473,N_3370,N_3302);
or U3474 (N_3474,N_3314,N_3380);
nor U3475 (N_3475,N_3365,N_3364);
nor U3476 (N_3476,N_3303,N_3396);
nand U3477 (N_3477,N_3342,N_3375);
and U3478 (N_3478,N_3327,N_3331);
nor U3479 (N_3479,N_3329,N_3311);
and U3480 (N_3480,N_3314,N_3307);
nand U3481 (N_3481,N_3347,N_3379);
and U3482 (N_3482,N_3380,N_3358);
nand U3483 (N_3483,N_3346,N_3399);
nor U3484 (N_3484,N_3362,N_3349);
nand U3485 (N_3485,N_3318,N_3387);
and U3486 (N_3486,N_3314,N_3303);
or U3487 (N_3487,N_3329,N_3356);
nand U3488 (N_3488,N_3359,N_3364);
or U3489 (N_3489,N_3363,N_3343);
xnor U3490 (N_3490,N_3345,N_3326);
nor U3491 (N_3491,N_3324,N_3322);
nand U3492 (N_3492,N_3379,N_3382);
and U3493 (N_3493,N_3353,N_3306);
and U3494 (N_3494,N_3378,N_3346);
or U3495 (N_3495,N_3342,N_3308);
nor U3496 (N_3496,N_3313,N_3306);
nor U3497 (N_3497,N_3309,N_3339);
or U3498 (N_3498,N_3318,N_3347);
nand U3499 (N_3499,N_3369,N_3360);
nand U3500 (N_3500,N_3465,N_3448);
or U3501 (N_3501,N_3497,N_3443);
nor U3502 (N_3502,N_3469,N_3417);
nand U3503 (N_3503,N_3483,N_3479);
or U3504 (N_3504,N_3423,N_3488);
or U3505 (N_3505,N_3413,N_3401);
and U3506 (N_3506,N_3429,N_3486);
nand U3507 (N_3507,N_3482,N_3480);
nand U3508 (N_3508,N_3415,N_3414);
xor U3509 (N_3509,N_3406,N_3453);
or U3510 (N_3510,N_3476,N_3427);
nor U3511 (N_3511,N_3438,N_3475);
xnor U3512 (N_3512,N_3439,N_3430);
nor U3513 (N_3513,N_3462,N_3421);
xnor U3514 (N_3514,N_3418,N_3425);
nand U3515 (N_3515,N_3447,N_3440);
nand U3516 (N_3516,N_3409,N_3410);
xnor U3517 (N_3517,N_3412,N_3446);
nor U3518 (N_3518,N_3435,N_3422);
and U3519 (N_3519,N_3464,N_3411);
and U3520 (N_3520,N_3481,N_3470);
nor U3521 (N_3521,N_3485,N_3477);
and U3522 (N_3522,N_3437,N_3451);
or U3523 (N_3523,N_3463,N_3472);
xor U3524 (N_3524,N_3441,N_3433);
and U3525 (N_3525,N_3499,N_3407);
nor U3526 (N_3526,N_3408,N_3400);
and U3527 (N_3527,N_3402,N_3420);
nand U3528 (N_3528,N_3404,N_3426);
nor U3529 (N_3529,N_3436,N_3491);
nor U3530 (N_3530,N_3494,N_3484);
or U3531 (N_3531,N_3444,N_3496);
xor U3532 (N_3532,N_3474,N_3489);
or U3533 (N_3533,N_3450,N_3466);
nand U3534 (N_3534,N_3492,N_3468);
and U3535 (N_3535,N_3460,N_3432);
xor U3536 (N_3536,N_3452,N_3487);
nand U3537 (N_3537,N_3473,N_3458);
xnor U3538 (N_3538,N_3416,N_3498);
xnor U3539 (N_3539,N_3459,N_3457);
xnor U3540 (N_3540,N_3467,N_3419);
nor U3541 (N_3541,N_3431,N_3495);
or U3542 (N_3542,N_3442,N_3403);
nand U3543 (N_3543,N_3461,N_3490);
nand U3544 (N_3544,N_3478,N_3454);
xnor U3545 (N_3545,N_3471,N_3428);
xnor U3546 (N_3546,N_3405,N_3449);
or U3547 (N_3547,N_3456,N_3493);
or U3548 (N_3548,N_3455,N_3434);
nor U3549 (N_3549,N_3445,N_3424);
or U3550 (N_3550,N_3496,N_3427);
nor U3551 (N_3551,N_3410,N_3416);
nand U3552 (N_3552,N_3407,N_3404);
nor U3553 (N_3553,N_3466,N_3433);
xor U3554 (N_3554,N_3493,N_3498);
nor U3555 (N_3555,N_3425,N_3402);
or U3556 (N_3556,N_3447,N_3435);
nand U3557 (N_3557,N_3485,N_3430);
xor U3558 (N_3558,N_3475,N_3430);
and U3559 (N_3559,N_3440,N_3412);
nor U3560 (N_3560,N_3469,N_3419);
or U3561 (N_3561,N_3457,N_3429);
and U3562 (N_3562,N_3479,N_3458);
nand U3563 (N_3563,N_3490,N_3452);
xor U3564 (N_3564,N_3489,N_3439);
and U3565 (N_3565,N_3486,N_3468);
nand U3566 (N_3566,N_3412,N_3410);
or U3567 (N_3567,N_3498,N_3488);
nor U3568 (N_3568,N_3474,N_3400);
nor U3569 (N_3569,N_3482,N_3412);
xnor U3570 (N_3570,N_3400,N_3463);
xor U3571 (N_3571,N_3422,N_3467);
xor U3572 (N_3572,N_3463,N_3438);
or U3573 (N_3573,N_3495,N_3467);
xor U3574 (N_3574,N_3472,N_3441);
nand U3575 (N_3575,N_3445,N_3468);
nand U3576 (N_3576,N_3420,N_3437);
nand U3577 (N_3577,N_3480,N_3478);
nand U3578 (N_3578,N_3496,N_3429);
or U3579 (N_3579,N_3438,N_3442);
and U3580 (N_3580,N_3425,N_3445);
nand U3581 (N_3581,N_3408,N_3410);
and U3582 (N_3582,N_3492,N_3498);
or U3583 (N_3583,N_3461,N_3492);
nor U3584 (N_3584,N_3458,N_3446);
nand U3585 (N_3585,N_3425,N_3446);
xor U3586 (N_3586,N_3452,N_3460);
and U3587 (N_3587,N_3423,N_3402);
or U3588 (N_3588,N_3451,N_3413);
nor U3589 (N_3589,N_3423,N_3421);
or U3590 (N_3590,N_3440,N_3463);
nand U3591 (N_3591,N_3425,N_3466);
and U3592 (N_3592,N_3494,N_3479);
and U3593 (N_3593,N_3471,N_3473);
or U3594 (N_3594,N_3442,N_3473);
nor U3595 (N_3595,N_3476,N_3434);
nand U3596 (N_3596,N_3404,N_3457);
or U3597 (N_3597,N_3452,N_3432);
nor U3598 (N_3598,N_3402,N_3484);
or U3599 (N_3599,N_3406,N_3417);
or U3600 (N_3600,N_3578,N_3531);
nor U3601 (N_3601,N_3551,N_3550);
nand U3602 (N_3602,N_3585,N_3504);
nor U3603 (N_3603,N_3517,N_3577);
nand U3604 (N_3604,N_3536,N_3575);
nand U3605 (N_3605,N_3555,N_3553);
or U3606 (N_3606,N_3518,N_3522);
nand U3607 (N_3607,N_3594,N_3540);
or U3608 (N_3608,N_3502,N_3547);
xnor U3609 (N_3609,N_3588,N_3533);
nor U3610 (N_3610,N_3520,N_3511);
and U3611 (N_3611,N_3507,N_3526);
xnor U3612 (N_3612,N_3599,N_3557);
xor U3613 (N_3613,N_3552,N_3560);
nand U3614 (N_3614,N_3589,N_3505);
nor U3615 (N_3615,N_3597,N_3506);
and U3616 (N_3616,N_3568,N_3556);
and U3617 (N_3617,N_3580,N_3545);
nand U3618 (N_3618,N_3570,N_3583);
or U3619 (N_3619,N_3581,N_3530);
nand U3620 (N_3620,N_3500,N_3527);
and U3621 (N_3621,N_3532,N_3584);
nor U3622 (N_3622,N_3528,N_3567);
nor U3623 (N_3623,N_3537,N_3513);
or U3624 (N_3624,N_3563,N_3579);
or U3625 (N_3625,N_3587,N_3590);
nand U3626 (N_3626,N_3571,N_3591);
and U3627 (N_3627,N_3566,N_3501);
or U3628 (N_3628,N_3573,N_3525);
nand U3629 (N_3629,N_3539,N_3582);
nor U3630 (N_3630,N_3598,N_3512);
xnor U3631 (N_3631,N_3574,N_3503);
or U3632 (N_3632,N_3538,N_3509);
xnor U3633 (N_3633,N_3562,N_3595);
nand U3634 (N_3634,N_3554,N_3543);
or U3635 (N_3635,N_3576,N_3546);
and U3636 (N_3636,N_3558,N_3549);
nand U3637 (N_3637,N_3559,N_3593);
nor U3638 (N_3638,N_3510,N_3524);
and U3639 (N_3639,N_3586,N_3515);
nor U3640 (N_3640,N_3544,N_3592);
xnor U3641 (N_3641,N_3561,N_3519);
or U3642 (N_3642,N_3565,N_3569);
or U3643 (N_3643,N_3572,N_3514);
and U3644 (N_3644,N_3535,N_3542);
or U3645 (N_3645,N_3541,N_3548);
nand U3646 (N_3646,N_3523,N_3564);
or U3647 (N_3647,N_3596,N_3534);
nor U3648 (N_3648,N_3521,N_3508);
nand U3649 (N_3649,N_3529,N_3516);
xor U3650 (N_3650,N_3578,N_3581);
nand U3651 (N_3651,N_3522,N_3527);
nor U3652 (N_3652,N_3559,N_3539);
nand U3653 (N_3653,N_3508,N_3514);
or U3654 (N_3654,N_3536,N_3559);
and U3655 (N_3655,N_3584,N_3536);
xor U3656 (N_3656,N_3554,N_3503);
nand U3657 (N_3657,N_3593,N_3541);
nor U3658 (N_3658,N_3572,N_3533);
xor U3659 (N_3659,N_3578,N_3566);
nand U3660 (N_3660,N_3547,N_3503);
and U3661 (N_3661,N_3581,N_3528);
or U3662 (N_3662,N_3537,N_3505);
xnor U3663 (N_3663,N_3509,N_3504);
nor U3664 (N_3664,N_3562,N_3556);
xnor U3665 (N_3665,N_3562,N_3508);
or U3666 (N_3666,N_3555,N_3503);
nand U3667 (N_3667,N_3563,N_3505);
nor U3668 (N_3668,N_3530,N_3573);
and U3669 (N_3669,N_3551,N_3573);
nor U3670 (N_3670,N_3590,N_3517);
nand U3671 (N_3671,N_3538,N_3527);
nor U3672 (N_3672,N_3551,N_3510);
nand U3673 (N_3673,N_3577,N_3506);
and U3674 (N_3674,N_3506,N_3545);
nor U3675 (N_3675,N_3560,N_3595);
nor U3676 (N_3676,N_3532,N_3519);
nor U3677 (N_3677,N_3504,N_3529);
xnor U3678 (N_3678,N_3527,N_3595);
xor U3679 (N_3679,N_3575,N_3530);
or U3680 (N_3680,N_3533,N_3593);
nand U3681 (N_3681,N_3556,N_3565);
nand U3682 (N_3682,N_3518,N_3553);
nor U3683 (N_3683,N_3556,N_3560);
nor U3684 (N_3684,N_3583,N_3511);
nand U3685 (N_3685,N_3507,N_3534);
or U3686 (N_3686,N_3557,N_3521);
xor U3687 (N_3687,N_3594,N_3573);
xnor U3688 (N_3688,N_3589,N_3598);
or U3689 (N_3689,N_3556,N_3511);
or U3690 (N_3690,N_3563,N_3541);
and U3691 (N_3691,N_3527,N_3543);
nand U3692 (N_3692,N_3514,N_3599);
nand U3693 (N_3693,N_3541,N_3557);
or U3694 (N_3694,N_3575,N_3539);
and U3695 (N_3695,N_3509,N_3584);
xor U3696 (N_3696,N_3589,N_3522);
nor U3697 (N_3697,N_3561,N_3516);
and U3698 (N_3698,N_3556,N_3514);
xnor U3699 (N_3699,N_3512,N_3510);
nor U3700 (N_3700,N_3625,N_3642);
and U3701 (N_3701,N_3677,N_3612);
and U3702 (N_3702,N_3694,N_3683);
or U3703 (N_3703,N_3688,N_3641);
nand U3704 (N_3704,N_3660,N_3614);
nor U3705 (N_3705,N_3600,N_3621);
and U3706 (N_3706,N_3629,N_3664);
and U3707 (N_3707,N_3671,N_3645);
nor U3708 (N_3708,N_3681,N_3636);
nand U3709 (N_3709,N_3673,N_3655);
and U3710 (N_3710,N_3663,N_3689);
or U3711 (N_3711,N_3640,N_3691);
nor U3712 (N_3712,N_3674,N_3675);
and U3713 (N_3713,N_3633,N_3653);
xor U3714 (N_3714,N_3661,N_3658);
xnor U3715 (N_3715,N_3698,N_3650);
nand U3716 (N_3716,N_3638,N_3649);
nand U3717 (N_3717,N_3682,N_3632);
xor U3718 (N_3718,N_3695,N_3631);
xnor U3719 (N_3719,N_3666,N_3685);
nand U3720 (N_3720,N_3680,N_3659);
nor U3721 (N_3721,N_3607,N_3654);
and U3722 (N_3722,N_3647,N_3684);
and U3723 (N_3723,N_3616,N_3678);
nand U3724 (N_3724,N_3622,N_3696);
and U3725 (N_3725,N_3686,N_3652);
xnor U3726 (N_3726,N_3603,N_3609);
or U3727 (N_3727,N_3630,N_3639);
and U3728 (N_3728,N_3608,N_3667);
or U3729 (N_3729,N_3613,N_3615);
or U3730 (N_3730,N_3693,N_3610);
nand U3731 (N_3731,N_3692,N_3637);
and U3732 (N_3732,N_3602,N_3651);
nand U3733 (N_3733,N_3670,N_3676);
or U3734 (N_3734,N_3699,N_3604);
xnor U3735 (N_3735,N_3620,N_3665);
and U3736 (N_3736,N_3605,N_3634);
nand U3737 (N_3737,N_3624,N_3617);
nor U3738 (N_3738,N_3635,N_3626);
nor U3739 (N_3739,N_3687,N_3669);
xnor U3740 (N_3740,N_3627,N_3643);
nand U3741 (N_3741,N_3668,N_3672);
or U3742 (N_3742,N_3628,N_3662);
or U3743 (N_3743,N_3648,N_3656);
and U3744 (N_3744,N_3618,N_3679);
or U3745 (N_3745,N_3611,N_3619);
xor U3746 (N_3746,N_3646,N_3690);
xnor U3747 (N_3747,N_3657,N_3644);
nor U3748 (N_3748,N_3623,N_3697);
or U3749 (N_3749,N_3606,N_3601);
and U3750 (N_3750,N_3653,N_3691);
nor U3751 (N_3751,N_3633,N_3676);
nand U3752 (N_3752,N_3681,N_3648);
and U3753 (N_3753,N_3606,N_3695);
nand U3754 (N_3754,N_3659,N_3650);
nand U3755 (N_3755,N_3612,N_3692);
xor U3756 (N_3756,N_3691,N_3607);
or U3757 (N_3757,N_3689,N_3642);
and U3758 (N_3758,N_3664,N_3619);
nor U3759 (N_3759,N_3636,N_3663);
nor U3760 (N_3760,N_3683,N_3613);
and U3761 (N_3761,N_3644,N_3604);
nand U3762 (N_3762,N_3684,N_3611);
and U3763 (N_3763,N_3685,N_3623);
nand U3764 (N_3764,N_3610,N_3601);
nor U3765 (N_3765,N_3688,N_3623);
or U3766 (N_3766,N_3616,N_3625);
nand U3767 (N_3767,N_3685,N_3634);
nor U3768 (N_3768,N_3608,N_3677);
nor U3769 (N_3769,N_3683,N_3646);
nand U3770 (N_3770,N_3646,N_3688);
nand U3771 (N_3771,N_3602,N_3650);
or U3772 (N_3772,N_3618,N_3672);
xor U3773 (N_3773,N_3611,N_3637);
or U3774 (N_3774,N_3661,N_3688);
and U3775 (N_3775,N_3617,N_3686);
or U3776 (N_3776,N_3656,N_3693);
and U3777 (N_3777,N_3622,N_3642);
xor U3778 (N_3778,N_3685,N_3640);
xor U3779 (N_3779,N_3683,N_3635);
nand U3780 (N_3780,N_3684,N_3627);
xor U3781 (N_3781,N_3697,N_3625);
xor U3782 (N_3782,N_3606,N_3635);
or U3783 (N_3783,N_3675,N_3656);
or U3784 (N_3784,N_3665,N_3674);
and U3785 (N_3785,N_3658,N_3691);
or U3786 (N_3786,N_3654,N_3614);
or U3787 (N_3787,N_3679,N_3666);
and U3788 (N_3788,N_3661,N_3643);
or U3789 (N_3789,N_3628,N_3679);
nand U3790 (N_3790,N_3682,N_3620);
nor U3791 (N_3791,N_3655,N_3660);
and U3792 (N_3792,N_3656,N_3671);
and U3793 (N_3793,N_3610,N_3631);
nand U3794 (N_3794,N_3629,N_3660);
and U3795 (N_3795,N_3644,N_3621);
and U3796 (N_3796,N_3687,N_3690);
xnor U3797 (N_3797,N_3643,N_3639);
xor U3798 (N_3798,N_3691,N_3635);
or U3799 (N_3799,N_3670,N_3674);
xnor U3800 (N_3800,N_3750,N_3732);
nor U3801 (N_3801,N_3752,N_3780);
or U3802 (N_3802,N_3799,N_3766);
xor U3803 (N_3803,N_3737,N_3747);
nand U3804 (N_3804,N_3704,N_3702);
or U3805 (N_3805,N_3713,N_3764);
and U3806 (N_3806,N_3746,N_3719);
and U3807 (N_3807,N_3794,N_3792);
nor U3808 (N_3808,N_3768,N_3724);
and U3809 (N_3809,N_3729,N_3701);
xnor U3810 (N_3810,N_3756,N_3765);
nand U3811 (N_3811,N_3797,N_3711);
xor U3812 (N_3812,N_3790,N_3735);
or U3813 (N_3813,N_3744,N_3774);
or U3814 (N_3814,N_3721,N_3789);
nor U3815 (N_3815,N_3771,N_3754);
and U3816 (N_3816,N_3725,N_3762);
xnor U3817 (N_3817,N_3784,N_3796);
or U3818 (N_3818,N_3733,N_3753);
and U3819 (N_3819,N_3782,N_3761);
xnor U3820 (N_3820,N_3738,N_3775);
nand U3821 (N_3821,N_3706,N_3730);
or U3822 (N_3822,N_3748,N_3755);
nand U3823 (N_3823,N_3749,N_3708);
nand U3824 (N_3824,N_3716,N_3714);
xor U3825 (N_3825,N_3722,N_3791);
and U3826 (N_3826,N_3778,N_3787);
nor U3827 (N_3827,N_3763,N_3788);
xnor U3828 (N_3828,N_3795,N_3743);
nor U3829 (N_3829,N_3734,N_3741);
and U3830 (N_3830,N_3703,N_3793);
nor U3831 (N_3831,N_3717,N_3783);
xor U3832 (N_3832,N_3723,N_3777);
nor U3833 (N_3833,N_3707,N_3731);
nor U3834 (N_3834,N_3710,N_3776);
and U3835 (N_3835,N_3705,N_3798);
xnor U3836 (N_3836,N_3785,N_3712);
nor U3837 (N_3837,N_3700,N_3727);
and U3838 (N_3838,N_3751,N_3767);
and U3839 (N_3839,N_3779,N_3757);
nand U3840 (N_3840,N_3786,N_3770);
and U3841 (N_3841,N_3760,N_3758);
nor U3842 (N_3842,N_3781,N_3709);
nand U3843 (N_3843,N_3728,N_3759);
and U3844 (N_3844,N_3739,N_3740);
or U3845 (N_3845,N_3769,N_3773);
xor U3846 (N_3846,N_3720,N_3745);
nand U3847 (N_3847,N_3715,N_3742);
and U3848 (N_3848,N_3772,N_3736);
or U3849 (N_3849,N_3726,N_3718);
nor U3850 (N_3850,N_3747,N_3719);
or U3851 (N_3851,N_3704,N_3787);
xor U3852 (N_3852,N_3773,N_3789);
and U3853 (N_3853,N_3752,N_3717);
and U3854 (N_3854,N_3739,N_3726);
nor U3855 (N_3855,N_3732,N_3786);
nor U3856 (N_3856,N_3746,N_3736);
and U3857 (N_3857,N_3761,N_3701);
nor U3858 (N_3858,N_3778,N_3755);
or U3859 (N_3859,N_3780,N_3766);
xor U3860 (N_3860,N_3791,N_3748);
or U3861 (N_3861,N_3729,N_3753);
and U3862 (N_3862,N_3727,N_3750);
and U3863 (N_3863,N_3754,N_3724);
and U3864 (N_3864,N_3713,N_3779);
xnor U3865 (N_3865,N_3739,N_3748);
xnor U3866 (N_3866,N_3737,N_3773);
and U3867 (N_3867,N_3734,N_3780);
xor U3868 (N_3868,N_3701,N_3730);
nor U3869 (N_3869,N_3709,N_3740);
nand U3870 (N_3870,N_3762,N_3716);
nor U3871 (N_3871,N_3715,N_3759);
xnor U3872 (N_3872,N_3742,N_3718);
xor U3873 (N_3873,N_3743,N_3770);
and U3874 (N_3874,N_3722,N_3772);
nor U3875 (N_3875,N_3793,N_3751);
nand U3876 (N_3876,N_3751,N_3710);
nor U3877 (N_3877,N_3701,N_3779);
nand U3878 (N_3878,N_3799,N_3710);
nor U3879 (N_3879,N_3764,N_3709);
or U3880 (N_3880,N_3730,N_3797);
and U3881 (N_3881,N_3768,N_3776);
and U3882 (N_3882,N_3759,N_3751);
nor U3883 (N_3883,N_3732,N_3773);
and U3884 (N_3884,N_3771,N_3770);
xnor U3885 (N_3885,N_3740,N_3712);
or U3886 (N_3886,N_3775,N_3776);
nor U3887 (N_3887,N_3733,N_3740);
or U3888 (N_3888,N_3767,N_3768);
or U3889 (N_3889,N_3703,N_3709);
xor U3890 (N_3890,N_3736,N_3782);
and U3891 (N_3891,N_3709,N_3776);
or U3892 (N_3892,N_3702,N_3745);
or U3893 (N_3893,N_3737,N_3782);
nor U3894 (N_3894,N_3795,N_3794);
nand U3895 (N_3895,N_3713,N_3756);
nor U3896 (N_3896,N_3724,N_3711);
and U3897 (N_3897,N_3766,N_3709);
or U3898 (N_3898,N_3759,N_3768);
nor U3899 (N_3899,N_3701,N_3728);
and U3900 (N_3900,N_3879,N_3816);
nand U3901 (N_3901,N_3860,N_3868);
nor U3902 (N_3902,N_3882,N_3835);
xnor U3903 (N_3903,N_3834,N_3845);
and U3904 (N_3904,N_3852,N_3881);
nand U3905 (N_3905,N_3854,N_3814);
nand U3906 (N_3906,N_3862,N_3877);
or U3907 (N_3907,N_3819,N_3828);
nand U3908 (N_3908,N_3846,N_3832);
xor U3909 (N_3909,N_3836,N_3840);
nor U3910 (N_3910,N_3839,N_3898);
nor U3911 (N_3911,N_3866,N_3893);
or U3912 (N_3912,N_3810,N_3821);
or U3913 (N_3913,N_3875,N_3829);
and U3914 (N_3914,N_3867,N_3831);
and U3915 (N_3915,N_3885,N_3856);
nor U3916 (N_3916,N_3892,N_3806);
or U3917 (N_3917,N_3849,N_3807);
xnor U3918 (N_3918,N_3818,N_3871);
xnor U3919 (N_3919,N_3890,N_3887);
xor U3920 (N_3920,N_3802,N_3817);
nor U3921 (N_3921,N_3891,N_3804);
nand U3922 (N_3922,N_3861,N_3894);
nand U3923 (N_3923,N_3876,N_3864);
nand U3924 (N_3924,N_3895,N_3873);
and U3925 (N_3925,N_3833,N_3803);
nand U3926 (N_3926,N_3838,N_3851);
and U3927 (N_3927,N_3886,N_3880);
nor U3928 (N_3928,N_3878,N_3865);
xnor U3929 (N_3929,N_3827,N_3824);
xnor U3930 (N_3930,N_3843,N_3857);
nor U3931 (N_3931,N_3809,N_3800);
xnor U3932 (N_3932,N_3842,N_3869);
nor U3933 (N_3933,N_3811,N_3841);
and U3934 (N_3934,N_3830,N_3844);
xnor U3935 (N_3935,N_3863,N_3801);
xnor U3936 (N_3936,N_3808,N_3897);
nor U3937 (N_3937,N_3889,N_3888);
or U3938 (N_3938,N_3859,N_3874);
nand U3939 (N_3939,N_3823,N_3815);
xor U3940 (N_3940,N_3813,N_3899);
nand U3941 (N_3941,N_3826,N_3822);
nor U3942 (N_3942,N_3850,N_3870);
xnor U3943 (N_3943,N_3872,N_3883);
nor U3944 (N_3944,N_3858,N_3847);
nor U3945 (N_3945,N_3848,N_3853);
nor U3946 (N_3946,N_3820,N_3855);
and U3947 (N_3947,N_3896,N_3825);
xor U3948 (N_3948,N_3805,N_3884);
or U3949 (N_3949,N_3812,N_3837);
and U3950 (N_3950,N_3854,N_3816);
nor U3951 (N_3951,N_3899,N_3897);
nand U3952 (N_3952,N_3850,N_3890);
xor U3953 (N_3953,N_3887,N_3832);
and U3954 (N_3954,N_3896,N_3819);
or U3955 (N_3955,N_3832,N_3820);
xnor U3956 (N_3956,N_3839,N_3837);
nand U3957 (N_3957,N_3836,N_3871);
or U3958 (N_3958,N_3861,N_3822);
xnor U3959 (N_3959,N_3862,N_3838);
and U3960 (N_3960,N_3890,N_3855);
and U3961 (N_3961,N_3840,N_3810);
or U3962 (N_3962,N_3804,N_3826);
nand U3963 (N_3963,N_3827,N_3863);
nor U3964 (N_3964,N_3836,N_3898);
and U3965 (N_3965,N_3876,N_3852);
nor U3966 (N_3966,N_3863,N_3832);
or U3967 (N_3967,N_3848,N_3801);
xnor U3968 (N_3968,N_3879,N_3813);
or U3969 (N_3969,N_3832,N_3810);
nor U3970 (N_3970,N_3881,N_3856);
nand U3971 (N_3971,N_3808,N_3807);
or U3972 (N_3972,N_3820,N_3837);
xor U3973 (N_3973,N_3836,N_3832);
nor U3974 (N_3974,N_3898,N_3874);
and U3975 (N_3975,N_3831,N_3845);
xor U3976 (N_3976,N_3831,N_3841);
and U3977 (N_3977,N_3885,N_3876);
or U3978 (N_3978,N_3885,N_3846);
or U3979 (N_3979,N_3855,N_3831);
nor U3980 (N_3980,N_3806,N_3842);
or U3981 (N_3981,N_3870,N_3844);
nand U3982 (N_3982,N_3892,N_3879);
nor U3983 (N_3983,N_3896,N_3807);
xnor U3984 (N_3984,N_3837,N_3880);
or U3985 (N_3985,N_3827,N_3855);
nor U3986 (N_3986,N_3845,N_3835);
or U3987 (N_3987,N_3804,N_3852);
xor U3988 (N_3988,N_3857,N_3853);
xor U3989 (N_3989,N_3830,N_3875);
or U3990 (N_3990,N_3821,N_3895);
or U3991 (N_3991,N_3805,N_3879);
xnor U3992 (N_3992,N_3811,N_3809);
xor U3993 (N_3993,N_3845,N_3894);
xnor U3994 (N_3994,N_3833,N_3885);
or U3995 (N_3995,N_3833,N_3825);
xor U3996 (N_3996,N_3899,N_3821);
nand U3997 (N_3997,N_3863,N_3828);
nand U3998 (N_3998,N_3845,N_3827);
and U3999 (N_3999,N_3897,N_3809);
or U4000 (N_4000,N_3931,N_3966);
nand U4001 (N_4001,N_3901,N_3954);
xor U4002 (N_4002,N_3982,N_3988);
nand U4003 (N_4003,N_3958,N_3997);
xnor U4004 (N_4004,N_3915,N_3978);
nand U4005 (N_4005,N_3920,N_3971);
and U4006 (N_4006,N_3902,N_3918);
and U4007 (N_4007,N_3979,N_3928);
xnor U4008 (N_4008,N_3994,N_3984);
nor U4009 (N_4009,N_3998,N_3973);
xnor U4010 (N_4010,N_3912,N_3919);
and U4011 (N_4011,N_3989,N_3986);
nor U4012 (N_4012,N_3951,N_3910);
nor U4013 (N_4013,N_3903,N_3906);
or U4014 (N_4014,N_3991,N_3946);
and U4015 (N_4015,N_3957,N_3938);
xnor U4016 (N_4016,N_3900,N_3956);
nand U4017 (N_4017,N_3949,N_3965);
or U4018 (N_4018,N_3926,N_3977);
or U4019 (N_4019,N_3905,N_3996);
or U4020 (N_4020,N_3999,N_3941);
or U4021 (N_4021,N_3911,N_3927);
or U4022 (N_4022,N_3980,N_3960);
or U4023 (N_4023,N_3943,N_3908);
and U4024 (N_4024,N_3972,N_3962);
nor U4025 (N_4025,N_3955,N_3907);
xnor U4026 (N_4026,N_3942,N_3934);
nand U4027 (N_4027,N_3925,N_3913);
nor U4028 (N_4028,N_3953,N_3939);
xnor U4029 (N_4029,N_3940,N_3935);
nor U4030 (N_4030,N_3964,N_3947);
nand U4031 (N_4031,N_3975,N_3904);
or U4032 (N_4032,N_3922,N_3968);
nand U4033 (N_4033,N_3961,N_3916);
and U4034 (N_4034,N_3974,N_3944);
nor U4035 (N_4035,N_3970,N_3993);
xor U4036 (N_4036,N_3976,N_3950);
xnor U4037 (N_4037,N_3967,N_3995);
and U4038 (N_4038,N_3990,N_3963);
xnor U4039 (N_4039,N_3914,N_3969);
and U4040 (N_4040,N_3924,N_3952);
nand U4041 (N_4041,N_3959,N_3937);
nand U4042 (N_4042,N_3929,N_3985);
nor U4043 (N_4043,N_3930,N_3948);
nand U4044 (N_4044,N_3936,N_3945);
or U4045 (N_4045,N_3987,N_3921);
xor U4046 (N_4046,N_3981,N_3932);
and U4047 (N_4047,N_3983,N_3909);
nor U4048 (N_4048,N_3917,N_3923);
xnor U4049 (N_4049,N_3992,N_3933);
or U4050 (N_4050,N_3978,N_3925);
nor U4051 (N_4051,N_3964,N_3967);
or U4052 (N_4052,N_3931,N_3995);
and U4053 (N_4053,N_3944,N_3902);
or U4054 (N_4054,N_3981,N_3963);
nor U4055 (N_4055,N_3939,N_3994);
nand U4056 (N_4056,N_3964,N_3953);
xnor U4057 (N_4057,N_3998,N_3913);
nand U4058 (N_4058,N_3906,N_3905);
and U4059 (N_4059,N_3937,N_3976);
nand U4060 (N_4060,N_3997,N_3919);
or U4061 (N_4061,N_3901,N_3950);
or U4062 (N_4062,N_3989,N_3935);
xnor U4063 (N_4063,N_3995,N_3947);
xor U4064 (N_4064,N_3973,N_3969);
xor U4065 (N_4065,N_3950,N_3941);
and U4066 (N_4066,N_3901,N_3965);
nand U4067 (N_4067,N_3942,N_3975);
nand U4068 (N_4068,N_3906,N_3997);
nor U4069 (N_4069,N_3950,N_3974);
nand U4070 (N_4070,N_3902,N_3965);
and U4071 (N_4071,N_3916,N_3985);
xnor U4072 (N_4072,N_3988,N_3999);
and U4073 (N_4073,N_3988,N_3983);
and U4074 (N_4074,N_3938,N_3913);
nand U4075 (N_4075,N_3914,N_3935);
xnor U4076 (N_4076,N_3967,N_3951);
or U4077 (N_4077,N_3969,N_3927);
xnor U4078 (N_4078,N_3916,N_3918);
or U4079 (N_4079,N_3996,N_3929);
nand U4080 (N_4080,N_3977,N_3943);
or U4081 (N_4081,N_3964,N_3916);
xnor U4082 (N_4082,N_3992,N_3946);
xnor U4083 (N_4083,N_3992,N_3967);
nor U4084 (N_4084,N_3959,N_3984);
xor U4085 (N_4085,N_3932,N_3952);
and U4086 (N_4086,N_3950,N_3955);
and U4087 (N_4087,N_3927,N_3965);
xor U4088 (N_4088,N_3921,N_3957);
and U4089 (N_4089,N_3984,N_3944);
and U4090 (N_4090,N_3907,N_3938);
or U4091 (N_4091,N_3924,N_3970);
nor U4092 (N_4092,N_3964,N_3900);
nand U4093 (N_4093,N_3901,N_3907);
or U4094 (N_4094,N_3997,N_3909);
or U4095 (N_4095,N_3951,N_3921);
and U4096 (N_4096,N_3925,N_3989);
or U4097 (N_4097,N_3922,N_3961);
nand U4098 (N_4098,N_3973,N_3994);
nand U4099 (N_4099,N_3905,N_3937);
nand U4100 (N_4100,N_4017,N_4006);
xnor U4101 (N_4101,N_4047,N_4065);
and U4102 (N_4102,N_4066,N_4029);
nor U4103 (N_4103,N_4002,N_4090);
and U4104 (N_4104,N_4008,N_4075);
xor U4105 (N_4105,N_4068,N_4040);
xnor U4106 (N_4106,N_4089,N_4081);
xor U4107 (N_4107,N_4013,N_4004);
xor U4108 (N_4108,N_4018,N_4059);
xor U4109 (N_4109,N_4034,N_4020);
xor U4110 (N_4110,N_4045,N_4028);
nor U4111 (N_4111,N_4055,N_4063);
nand U4112 (N_4112,N_4009,N_4019);
nand U4113 (N_4113,N_4038,N_4048);
or U4114 (N_4114,N_4007,N_4085);
or U4115 (N_4115,N_4073,N_4016);
or U4116 (N_4116,N_4051,N_4022);
or U4117 (N_4117,N_4094,N_4087);
nand U4118 (N_4118,N_4095,N_4097);
nor U4119 (N_4119,N_4082,N_4026);
and U4120 (N_4120,N_4084,N_4003);
nand U4121 (N_4121,N_4042,N_4091);
and U4122 (N_4122,N_4056,N_4024);
or U4123 (N_4123,N_4031,N_4067);
or U4124 (N_4124,N_4064,N_4032);
and U4125 (N_4125,N_4025,N_4060);
or U4126 (N_4126,N_4079,N_4076);
nor U4127 (N_4127,N_4012,N_4011);
nor U4128 (N_4128,N_4093,N_4061);
nand U4129 (N_4129,N_4099,N_4070);
or U4130 (N_4130,N_4027,N_4041);
xor U4131 (N_4131,N_4044,N_4058);
and U4132 (N_4132,N_4039,N_4033);
nor U4133 (N_4133,N_4010,N_4023);
nand U4134 (N_4134,N_4035,N_4037);
or U4135 (N_4135,N_4052,N_4021);
xor U4136 (N_4136,N_4050,N_4078);
and U4137 (N_4137,N_4005,N_4030);
or U4138 (N_4138,N_4086,N_4088);
nand U4139 (N_4139,N_4074,N_4046);
or U4140 (N_4140,N_4069,N_4054);
xor U4141 (N_4141,N_4072,N_4014);
xor U4142 (N_4142,N_4001,N_4036);
nor U4143 (N_4143,N_4080,N_4053);
or U4144 (N_4144,N_4096,N_4057);
nor U4145 (N_4145,N_4062,N_4092);
and U4146 (N_4146,N_4043,N_4049);
or U4147 (N_4147,N_4077,N_4098);
xor U4148 (N_4148,N_4071,N_4015);
or U4149 (N_4149,N_4000,N_4083);
nor U4150 (N_4150,N_4078,N_4034);
xnor U4151 (N_4151,N_4025,N_4079);
xnor U4152 (N_4152,N_4012,N_4039);
nand U4153 (N_4153,N_4081,N_4018);
xnor U4154 (N_4154,N_4012,N_4066);
nand U4155 (N_4155,N_4042,N_4053);
xnor U4156 (N_4156,N_4085,N_4078);
nor U4157 (N_4157,N_4081,N_4084);
nand U4158 (N_4158,N_4078,N_4057);
and U4159 (N_4159,N_4092,N_4039);
nor U4160 (N_4160,N_4096,N_4000);
xor U4161 (N_4161,N_4014,N_4052);
or U4162 (N_4162,N_4019,N_4070);
nand U4163 (N_4163,N_4032,N_4052);
xor U4164 (N_4164,N_4068,N_4000);
xor U4165 (N_4165,N_4002,N_4065);
or U4166 (N_4166,N_4034,N_4096);
and U4167 (N_4167,N_4030,N_4076);
nor U4168 (N_4168,N_4082,N_4055);
xor U4169 (N_4169,N_4095,N_4052);
or U4170 (N_4170,N_4085,N_4098);
and U4171 (N_4171,N_4046,N_4007);
or U4172 (N_4172,N_4095,N_4018);
xor U4173 (N_4173,N_4074,N_4063);
or U4174 (N_4174,N_4001,N_4013);
nor U4175 (N_4175,N_4037,N_4084);
nor U4176 (N_4176,N_4031,N_4051);
and U4177 (N_4177,N_4070,N_4051);
xnor U4178 (N_4178,N_4041,N_4010);
nand U4179 (N_4179,N_4039,N_4099);
nand U4180 (N_4180,N_4072,N_4096);
nand U4181 (N_4181,N_4035,N_4070);
nand U4182 (N_4182,N_4053,N_4016);
nor U4183 (N_4183,N_4049,N_4092);
and U4184 (N_4184,N_4031,N_4097);
xor U4185 (N_4185,N_4036,N_4035);
xnor U4186 (N_4186,N_4058,N_4016);
nor U4187 (N_4187,N_4056,N_4048);
xnor U4188 (N_4188,N_4026,N_4052);
and U4189 (N_4189,N_4007,N_4082);
nor U4190 (N_4190,N_4010,N_4001);
and U4191 (N_4191,N_4076,N_4092);
or U4192 (N_4192,N_4037,N_4066);
or U4193 (N_4193,N_4041,N_4090);
nand U4194 (N_4194,N_4018,N_4098);
xnor U4195 (N_4195,N_4028,N_4033);
nor U4196 (N_4196,N_4063,N_4062);
and U4197 (N_4197,N_4088,N_4091);
and U4198 (N_4198,N_4008,N_4082);
nor U4199 (N_4199,N_4027,N_4089);
or U4200 (N_4200,N_4175,N_4198);
or U4201 (N_4201,N_4174,N_4109);
and U4202 (N_4202,N_4164,N_4156);
nor U4203 (N_4203,N_4110,N_4135);
nor U4204 (N_4204,N_4183,N_4125);
nand U4205 (N_4205,N_4144,N_4193);
nand U4206 (N_4206,N_4181,N_4106);
xor U4207 (N_4207,N_4131,N_4163);
and U4208 (N_4208,N_4187,N_4158);
and U4209 (N_4209,N_4191,N_4132);
xnor U4210 (N_4210,N_4194,N_4113);
or U4211 (N_4211,N_4151,N_4153);
nor U4212 (N_4212,N_4178,N_4117);
nand U4213 (N_4213,N_4103,N_4139);
xnor U4214 (N_4214,N_4166,N_4108);
or U4215 (N_4215,N_4189,N_4124);
nor U4216 (N_4216,N_4197,N_4177);
nand U4217 (N_4217,N_4122,N_4167);
nor U4218 (N_4218,N_4185,N_4188);
nor U4219 (N_4219,N_4129,N_4172);
or U4220 (N_4220,N_4192,N_4162);
nand U4221 (N_4221,N_4196,N_4195);
or U4222 (N_4222,N_4141,N_4126);
or U4223 (N_4223,N_4115,N_4123);
or U4224 (N_4224,N_4155,N_4119);
and U4225 (N_4225,N_4143,N_4186);
xnor U4226 (N_4226,N_4147,N_4179);
and U4227 (N_4227,N_4148,N_4102);
nand U4228 (N_4228,N_4101,N_4168);
xor U4229 (N_4229,N_4142,N_4107);
xor U4230 (N_4230,N_4173,N_4138);
nand U4231 (N_4231,N_4160,N_4170);
nand U4232 (N_4232,N_4199,N_4130);
and U4233 (N_4233,N_4120,N_4159);
xor U4234 (N_4234,N_4104,N_4149);
xor U4235 (N_4235,N_4111,N_4116);
and U4236 (N_4236,N_4182,N_4150);
and U4237 (N_4237,N_4165,N_4161);
nand U4238 (N_4238,N_4154,N_4169);
nand U4239 (N_4239,N_4128,N_4136);
and U4240 (N_4240,N_4137,N_4184);
and U4241 (N_4241,N_4146,N_4134);
xor U4242 (N_4242,N_4121,N_4176);
nand U4243 (N_4243,N_4171,N_4190);
xor U4244 (N_4244,N_4157,N_4152);
nor U4245 (N_4245,N_4133,N_4118);
nor U4246 (N_4246,N_4105,N_4140);
or U4247 (N_4247,N_4127,N_4112);
nor U4248 (N_4248,N_4100,N_4114);
nand U4249 (N_4249,N_4145,N_4180);
or U4250 (N_4250,N_4154,N_4111);
nand U4251 (N_4251,N_4100,N_4151);
nand U4252 (N_4252,N_4192,N_4195);
nor U4253 (N_4253,N_4153,N_4147);
or U4254 (N_4254,N_4172,N_4184);
xnor U4255 (N_4255,N_4113,N_4184);
nor U4256 (N_4256,N_4101,N_4129);
nor U4257 (N_4257,N_4165,N_4134);
nor U4258 (N_4258,N_4157,N_4172);
nor U4259 (N_4259,N_4174,N_4177);
nor U4260 (N_4260,N_4178,N_4156);
or U4261 (N_4261,N_4193,N_4166);
xnor U4262 (N_4262,N_4174,N_4130);
nor U4263 (N_4263,N_4112,N_4193);
and U4264 (N_4264,N_4135,N_4174);
nor U4265 (N_4265,N_4151,N_4154);
and U4266 (N_4266,N_4193,N_4119);
nor U4267 (N_4267,N_4195,N_4130);
nor U4268 (N_4268,N_4146,N_4124);
nor U4269 (N_4269,N_4166,N_4197);
and U4270 (N_4270,N_4159,N_4188);
nor U4271 (N_4271,N_4191,N_4159);
nand U4272 (N_4272,N_4147,N_4123);
nand U4273 (N_4273,N_4121,N_4161);
or U4274 (N_4274,N_4190,N_4193);
nand U4275 (N_4275,N_4108,N_4133);
and U4276 (N_4276,N_4144,N_4113);
xnor U4277 (N_4277,N_4195,N_4189);
and U4278 (N_4278,N_4117,N_4104);
xor U4279 (N_4279,N_4107,N_4180);
xor U4280 (N_4280,N_4141,N_4131);
xor U4281 (N_4281,N_4145,N_4132);
nor U4282 (N_4282,N_4101,N_4155);
nor U4283 (N_4283,N_4178,N_4116);
xnor U4284 (N_4284,N_4188,N_4143);
or U4285 (N_4285,N_4106,N_4178);
nor U4286 (N_4286,N_4173,N_4133);
and U4287 (N_4287,N_4122,N_4153);
nor U4288 (N_4288,N_4162,N_4173);
or U4289 (N_4289,N_4127,N_4118);
or U4290 (N_4290,N_4112,N_4103);
xor U4291 (N_4291,N_4160,N_4187);
nor U4292 (N_4292,N_4121,N_4128);
nand U4293 (N_4293,N_4135,N_4106);
or U4294 (N_4294,N_4164,N_4139);
nand U4295 (N_4295,N_4185,N_4148);
nand U4296 (N_4296,N_4156,N_4124);
nand U4297 (N_4297,N_4168,N_4143);
nor U4298 (N_4298,N_4162,N_4127);
nor U4299 (N_4299,N_4117,N_4124);
and U4300 (N_4300,N_4278,N_4202);
nor U4301 (N_4301,N_4271,N_4269);
and U4302 (N_4302,N_4282,N_4294);
nor U4303 (N_4303,N_4215,N_4213);
nor U4304 (N_4304,N_4235,N_4273);
xnor U4305 (N_4305,N_4267,N_4258);
nor U4306 (N_4306,N_4204,N_4228);
xnor U4307 (N_4307,N_4232,N_4253);
nor U4308 (N_4308,N_4250,N_4219);
or U4309 (N_4309,N_4264,N_4262);
xor U4310 (N_4310,N_4206,N_4288);
or U4311 (N_4311,N_4257,N_4207);
or U4312 (N_4312,N_4244,N_4229);
nand U4313 (N_4313,N_4283,N_4254);
and U4314 (N_4314,N_4277,N_4281);
nor U4315 (N_4315,N_4200,N_4276);
nor U4316 (N_4316,N_4227,N_4241);
or U4317 (N_4317,N_4201,N_4266);
nor U4318 (N_4318,N_4223,N_4251);
nand U4319 (N_4319,N_4298,N_4295);
nor U4320 (N_4320,N_4230,N_4299);
nand U4321 (N_4321,N_4209,N_4239);
and U4322 (N_4322,N_4237,N_4234);
xnor U4323 (N_4323,N_4290,N_4212);
nor U4324 (N_4324,N_4225,N_4246);
nand U4325 (N_4325,N_4216,N_4256);
and U4326 (N_4326,N_4203,N_4272);
or U4327 (N_4327,N_4242,N_4211);
xor U4328 (N_4328,N_4289,N_4280);
nand U4329 (N_4329,N_4243,N_4221);
or U4330 (N_4330,N_4252,N_4296);
nand U4331 (N_4331,N_4247,N_4224);
nand U4332 (N_4332,N_4291,N_4268);
or U4333 (N_4333,N_4285,N_4210);
nor U4334 (N_4334,N_4208,N_4214);
nor U4335 (N_4335,N_4286,N_4261);
nor U4336 (N_4336,N_4292,N_4236);
and U4337 (N_4337,N_4259,N_4217);
or U4338 (N_4338,N_4260,N_4297);
xnor U4339 (N_4339,N_4293,N_4284);
and U4340 (N_4340,N_4205,N_4249);
nor U4341 (N_4341,N_4238,N_4245);
and U4342 (N_4342,N_4248,N_4275);
and U4343 (N_4343,N_4274,N_4231);
nand U4344 (N_4344,N_4222,N_4220);
nand U4345 (N_4345,N_4218,N_4263);
nor U4346 (N_4346,N_4265,N_4270);
nor U4347 (N_4347,N_4279,N_4226);
nor U4348 (N_4348,N_4233,N_4255);
xor U4349 (N_4349,N_4287,N_4240);
xor U4350 (N_4350,N_4233,N_4240);
xor U4351 (N_4351,N_4230,N_4217);
and U4352 (N_4352,N_4245,N_4287);
xor U4353 (N_4353,N_4211,N_4251);
and U4354 (N_4354,N_4295,N_4206);
nor U4355 (N_4355,N_4228,N_4272);
nand U4356 (N_4356,N_4290,N_4258);
and U4357 (N_4357,N_4266,N_4229);
nand U4358 (N_4358,N_4234,N_4264);
nor U4359 (N_4359,N_4210,N_4292);
nand U4360 (N_4360,N_4213,N_4293);
nor U4361 (N_4361,N_4253,N_4240);
and U4362 (N_4362,N_4229,N_4249);
nor U4363 (N_4363,N_4251,N_4289);
nor U4364 (N_4364,N_4242,N_4214);
or U4365 (N_4365,N_4255,N_4214);
nand U4366 (N_4366,N_4204,N_4256);
and U4367 (N_4367,N_4211,N_4221);
xor U4368 (N_4368,N_4202,N_4258);
nand U4369 (N_4369,N_4203,N_4222);
nor U4370 (N_4370,N_4230,N_4244);
xnor U4371 (N_4371,N_4295,N_4230);
xor U4372 (N_4372,N_4241,N_4232);
or U4373 (N_4373,N_4293,N_4231);
nand U4374 (N_4374,N_4274,N_4200);
nor U4375 (N_4375,N_4248,N_4237);
xor U4376 (N_4376,N_4206,N_4290);
xor U4377 (N_4377,N_4208,N_4265);
nand U4378 (N_4378,N_4209,N_4256);
and U4379 (N_4379,N_4200,N_4259);
nand U4380 (N_4380,N_4281,N_4208);
xnor U4381 (N_4381,N_4287,N_4249);
xnor U4382 (N_4382,N_4228,N_4265);
or U4383 (N_4383,N_4287,N_4248);
nand U4384 (N_4384,N_4228,N_4257);
and U4385 (N_4385,N_4275,N_4259);
nor U4386 (N_4386,N_4222,N_4279);
xor U4387 (N_4387,N_4293,N_4221);
and U4388 (N_4388,N_4248,N_4254);
and U4389 (N_4389,N_4267,N_4246);
nor U4390 (N_4390,N_4223,N_4267);
xor U4391 (N_4391,N_4205,N_4276);
or U4392 (N_4392,N_4217,N_4268);
xnor U4393 (N_4393,N_4246,N_4231);
nor U4394 (N_4394,N_4250,N_4291);
and U4395 (N_4395,N_4263,N_4214);
xnor U4396 (N_4396,N_4274,N_4222);
xor U4397 (N_4397,N_4266,N_4236);
xor U4398 (N_4398,N_4227,N_4283);
nand U4399 (N_4399,N_4246,N_4239);
nand U4400 (N_4400,N_4307,N_4393);
or U4401 (N_4401,N_4300,N_4335);
and U4402 (N_4402,N_4331,N_4398);
or U4403 (N_4403,N_4329,N_4389);
or U4404 (N_4404,N_4334,N_4348);
and U4405 (N_4405,N_4396,N_4303);
nand U4406 (N_4406,N_4302,N_4315);
xor U4407 (N_4407,N_4382,N_4336);
and U4408 (N_4408,N_4317,N_4308);
and U4409 (N_4409,N_4321,N_4352);
nand U4410 (N_4410,N_4310,N_4388);
and U4411 (N_4411,N_4373,N_4361);
and U4412 (N_4412,N_4316,N_4390);
or U4413 (N_4413,N_4319,N_4301);
or U4414 (N_4414,N_4347,N_4362);
or U4415 (N_4415,N_4392,N_4395);
nand U4416 (N_4416,N_4384,N_4351);
or U4417 (N_4417,N_4366,N_4344);
nand U4418 (N_4418,N_4354,N_4391);
nor U4419 (N_4419,N_4320,N_4376);
or U4420 (N_4420,N_4375,N_4333);
nor U4421 (N_4421,N_4364,N_4349);
nor U4422 (N_4422,N_4340,N_4324);
and U4423 (N_4423,N_4304,N_4394);
nand U4424 (N_4424,N_4318,N_4325);
nor U4425 (N_4425,N_4357,N_4353);
xor U4426 (N_4426,N_4328,N_4365);
nor U4427 (N_4427,N_4346,N_4314);
nand U4428 (N_4428,N_4332,N_4355);
xor U4429 (N_4429,N_4387,N_4327);
xnor U4430 (N_4430,N_4306,N_4305);
nand U4431 (N_4431,N_4311,N_4372);
nand U4432 (N_4432,N_4326,N_4399);
nor U4433 (N_4433,N_4379,N_4380);
xor U4434 (N_4434,N_4374,N_4323);
or U4435 (N_4435,N_4343,N_4397);
nor U4436 (N_4436,N_4339,N_4345);
nor U4437 (N_4437,N_4338,N_4342);
or U4438 (N_4438,N_4378,N_4330);
nor U4439 (N_4439,N_4322,N_4360);
xor U4440 (N_4440,N_4385,N_4359);
xor U4441 (N_4441,N_4369,N_4312);
and U4442 (N_4442,N_4356,N_4350);
xnor U4443 (N_4443,N_4309,N_4370);
and U4444 (N_4444,N_4377,N_4341);
nand U4445 (N_4445,N_4371,N_4381);
or U4446 (N_4446,N_4337,N_4368);
nor U4447 (N_4447,N_4386,N_4313);
xor U4448 (N_4448,N_4383,N_4367);
and U4449 (N_4449,N_4358,N_4363);
nand U4450 (N_4450,N_4365,N_4398);
nand U4451 (N_4451,N_4347,N_4358);
nor U4452 (N_4452,N_4395,N_4351);
and U4453 (N_4453,N_4328,N_4393);
and U4454 (N_4454,N_4373,N_4306);
nor U4455 (N_4455,N_4335,N_4334);
and U4456 (N_4456,N_4366,N_4368);
nand U4457 (N_4457,N_4312,N_4372);
nor U4458 (N_4458,N_4312,N_4379);
nand U4459 (N_4459,N_4305,N_4338);
xor U4460 (N_4460,N_4322,N_4331);
nand U4461 (N_4461,N_4399,N_4356);
nor U4462 (N_4462,N_4329,N_4363);
xnor U4463 (N_4463,N_4322,N_4361);
nor U4464 (N_4464,N_4356,N_4370);
and U4465 (N_4465,N_4382,N_4389);
nand U4466 (N_4466,N_4350,N_4391);
and U4467 (N_4467,N_4310,N_4391);
or U4468 (N_4468,N_4381,N_4370);
or U4469 (N_4469,N_4322,N_4373);
xnor U4470 (N_4470,N_4355,N_4359);
or U4471 (N_4471,N_4347,N_4313);
nand U4472 (N_4472,N_4360,N_4320);
nor U4473 (N_4473,N_4337,N_4305);
nor U4474 (N_4474,N_4366,N_4332);
nor U4475 (N_4475,N_4384,N_4366);
and U4476 (N_4476,N_4348,N_4346);
and U4477 (N_4477,N_4389,N_4312);
and U4478 (N_4478,N_4361,N_4370);
or U4479 (N_4479,N_4379,N_4391);
nand U4480 (N_4480,N_4361,N_4362);
nor U4481 (N_4481,N_4353,N_4313);
or U4482 (N_4482,N_4338,N_4388);
nand U4483 (N_4483,N_4332,N_4345);
or U4484 (N_4484,N_4392,N_4317);
xnor U4485 (N_4485,N_4349,N_4369);
or U4486 (N_4486,N_4366,N_4338);
xor U4487 (N_4487,N_4386,N_4310);
and U4488 (N_4488,N_4386,N_4342);
xor U4489 (N_4489,N_4385,N_4352);
xor U4490 (N_4490,N_4350,N_4354);
or U4491 (N_4491,N_4339,N_4321);
xnor U4492 (N_4492,N_4396,N_4335);
nor U4493 (N_4493,N_4328,N_4342);
xnor U4494 (N_4494,N_4362,N_4343);
xor U4495 (N_4495,N_4329,N_4399);
xnor U4496 (N_4496,N_4398,N_4362);
xor U4497 (N_4497,N_4311,N_4359);
or U4498 (N_4498,N_4344,N_4338);
or U4499 (N_4499,N_4374,N_4320);
nand U4500 (N_4500,N_4483,N_4479);
nand U4501 (N_4501,N_4467,N_4439);
and U4502 (N_4502,N_4469,N_4470);
xor U4503 (N_4503,N_4475,N_4468);
xnor U4504 (N_4504,N_4496,N_4466);
or U4505 (N_4505,N_4445,N_4472);
and U4506 (N_4506,N_4489,N_4486);
or U4507 (N_4507,N_4443,N_4487);
xor U4508 (N_4508,N_4485,N_4406);
and U4509 (N_4509,N_4436,N_4451);
nor U4510 (N_4510,N_4463,N_4412);
xor U4511 (N_4511,N_4429,N_4449);
and U4512 (N_4512,N_4437,N_4401);
xnor U4513 (N_4513,N_4484,N_4461);
nor U4514 (N_4514,N_4454,N_4474);
nand U4515 (N_4515,N_4411,N_4482);
nand U4516 (N_4516,N_4435,N_4413);
nand U4517 (N_4517,N_4480,N_4433);
or U4518 (N_4518,N_4432,N_4418);
nand U4519 (N_4519,N_4428,N_4491);
xnor U4520 (N_4520,N_4416,N_4490);
nand U4521 (N_4521,N_4498,N_4438);
nor U4522 (N_4522,N_4465,N_4444);
nor U4523 (N_4523,N_4419,N_4442);
or U4524 (N_4524,N_4462,N_4414);
and U4525 (N_4525,N_4441,N_4464);
and U4526 (N_4526,N_4492,N_4446);
nor U4527 (N_4527,N_4497,N_4455);
nand U4528 (N_4528,N_4434,N_4477);
nor U4529 (N_4529,N_4424,N_4481);
nand U4530 (N_4530,N_4417,N_4456);
and U4531 (N_4531,N_4457,N_4425);
and U4532 (N_4532,N_4405,N_4409);
and U4533 (N_4533,N_4427,N_4460);
or U4534 (N_4534,N_4459,N_4488);
nor U4535 (N_4535,N_4430,N_4431);
nand U4536 (N_4536,N_4403,N_4494);
nor U4537 (N_4537,N_4471,N_4415);
and U4538 (N_4538,N_4458,N_4495);
nand U4539 (N_4539,N_4422,N_4410);
or U4540 (N_4540,N_4450,N_4408);
and U4541 (N_4541,N_4453,N_4476);
xnor U4542 (N_4542,N_4404,N_4420);
nand U4543 (N_4543,N_4452,N_4499);
or U4544 (N_4544,N_4400,N_4473);
nand U4545 (N_4545,N_4426,N_4448);
xnor U4546 (N_4546,N_4440,N_4407);
nand U4547 (N_4547,N_4447,N_4478);
nand U4548 (N_4548,N_4402,N_4421);
xnor U4549 (N_4549,N_4423,N_4493);
or U4550 (N_4550,N_4472,N_4489);
nor U4551 (N_4551,N_4460,N_4408);
nor U4552 (N_4552,N_4422,N_4419);
and U4553 (N_4553,N_4483,N_4433);
and U4554 (N_4554,N_4440,N_4488);
and U4555 (N_4555,N_4434,N_4469);
or U4556 (N_4556,N_4453,N_4439);
xnor U4557 (N_4557,N_4404,N_4402);
nor U4558 (N_4558,N_4487,N_4493);
or U4559 (N_4559,N_4446,N_4410);
nor U4560 (N_4560,N_4440,N_4496);
xnor U4561 (N_4561,N_4433,N_4454);
nor U4562 (N_4562,N_4405,N_4468);
and U4563 (N_4563,N_4493,N_4471);
or U4564 (N_4564,N_4423,N_4403);
nor U4565 (N_4565,N_4441,N_4488);
or U4566 (N_4566,N_4472,N_4405);
and U4567 (N_4567,N_4444,N_4457);
nor U4568 (N_4568,N_4412,N_4467);
nor U4569 (N_4569,N_4448,N_4429);
or U4570 (N_4570,N_4450,N_4401);
or U4571 (N_4571,N_4403,N_4499);
and U4572 (N_4572,N_4403,N_4445);
xor U4573 (N_4573,N_4481,N_4484);
xnor U4574 (N_4574,N_4449,N_4476);
or U4575 (N_4575,N_4496,N_4447);
nand U4576 (N_4576,N_4428,N_4499);
and U4577 (N_4577,N_4457,N_4409);
nor U4578 (N_4578,N_4433,N_4491);
xnor U4579 (N_4579,N_4430,N_4421);
nand U4580 (N_4580,N_4461,N_4407);
nor U4581 (N_4581,N_4437,N_4462);
and U4582 (N_4582,N_4423,N_4411);
xnor U4583 (N_4583,N_4449,N_4434);
and U4584 (N_4584,N_4479,N_4490);
nor U4585 (N_4585,N_4453,N_4499);
nor U4586 (N_4586,N_4460,N_4467);
or U4587 (N_4587,N_4416,N_4451);
and U4588 (N_4588,N_4447,N_4449);
nand U4589 (N_4589,N_4413,N_4410);
xor U4590 (N_4590,N_4466,N_4479);
nand U4591 (N_4591,N_4475,N_4423);
xor U4592 (N_4592,N_4487,N_4484);
or U4593 (N_4593,N_4427,N_4441);
nand U4594 (N_4594,N_4492,N_4428);
xor U4595 (N_4595,N_4420,N_4445);
nand U4596 (N_4596,N_4444,N_4416);
and U4597 (N_4597,N_4493,N_4420);
nand U4598 (N_4598,N_4484,N_4426);
and U4599 (N_4599,N_4467,N_4426);
nand U4600 (N_4600,N_4549,N_4567);
or U4601 (N_4601,N_4518,N_4581);
nor U4602 (N_4602,N_4527,N_4520);
and U4603 (N_4603,N_4595,N_4557);
nand U4604 (N_4604,N_4589,N_4584);
nor U4605 (N_4605,N_4531,N_4524);
nand U4606 (N_4606,N_4513,N_4517);
nand U4607 (N_4607,N_4574,N_4550);
nand U4608 (N_4608,N_4534,N_4539);
or U4609 (N_4609,N_4522,N_4537);
or U4610 (N_4610,N_4500,N_4556);
or U4611 (N_4611,N_4596,N_4583);
or U4612 (N_4612,N_4558,N_4515);
or U4613 (N_4613,N_4573,N_4501);
nor U4614 (N_4614,N_4536,N_4535);
or U4615 (N_4615,N_4553,N_4597);
xnor U4616 (N_4616,N_4594,N_4504);
and U4617 (N_4617,N_4571,N_4590);
and U4618 (N_4618,N_4580,N_4554);
or U4619 (N_4619,N_4587,N_4545);
and U4620 (N_4620,N_4561,N_4514);
nand U4621 (N_4621,N_4546,N_4502);
and U4622 (N_4622,N_4541,N_4523);
nand U4623 (N_4623,N_4563,N_4598);
nor U4624 (N_4624,N_4565,N_4562);
nor U4625 (N_4625,N_4559,N_4506);
xor U4626 (N_4626,N_4525,N_4579);
nor U4627 (N_4627,N_4585,N_4582);
nor U4628 (N_4628,N_4555,N_4540);
xnor U4629 (N_4629,N_4577,N_4512);
and U4630 (N_4630,N_4551,N_4552);
nor U4631 (N_4631,N_4566,N_4521);
and U4632 (N_4632,N_4572,N_4511);
and U4633 (N_4633,N_4560,N_4528);
nand U4634 (N_4634,N_4570,N_4516);
or U4635 (N_4635,N_4586,N_4519);
xor U4636 (N_4636,N_4530,N_4591);
and U4637 (N_4637,N_4588,N_4508);
nor U4638 (N_4638,N_4533,N_4569);
or U4639 (N_4639,N_4529,N_4509);
nor U4640 (N_4640,N_4507,N_4505);
or U4641 (N_4641,N_4532,N_4578);
and U4642 (N_4642,N_4526,N_4544);
nand U4643 (N_4643,N_4576,N_4593);
xnor U4644 (N_4644,N_4599,N_4542);
or U4645 (N_4645,N_4568,N_4538);
or U4646 (N_4646,N_4575,N_4592);
xor U4647 (N_4647,N_4503,N_4510);
or U4648 (N_4648,N_4564,N_4543);
nor U4649 (N_4649,N_4548,N_4547);
nor U4650 (N_4650,N_4554,N_4589);
or U4651 (N_4651,N_4520,N_4542);
and U4652 (N_4652,N_4513,N_4582);
nand U4653 (N_4653,N_4521,N_4533);
nor U4654 (N_4654,N_4501,N_4551);
nor U4655 (N_4655,N_4530,N_4503);
nand U4656 (N_4656,N_4537,N_4515);
nand U4657 (N_4657,N_4593,N_4519);
or U4658 (N_4658,N_4550,N_4596);
nand U4659 (N_4659,N_4570,N_4545);
or U4660 (N_4660,N_4501,N_4589);
and U4661 (N_4661,N_4570,N_4576);
nand U4662 (N_4662,N_4561,N_4560);
and U4663 (N_4663,N_4545,N_4559);
nand U4664 (N_4664,N_4534,N_4533);
nand U4665 (N_4665,N_4579,N_4514);
xnor U4666 (N_4666,N_4562,N_4504);
or U4667 (N_4667,N_4523,N_4596);
nor U4668 (N_4668,N_4563,N_4577);
and U4669 (N_4669,N_4582,N_4599);
or U4670 (N_4670,N_4565,N_4588);
nand U4671 (N_4671,N_4563,N_4593);
nor U4672 (N_4672,N_4524,N_4562);
nor U4673 (N_4673,N_4542,N_4532);
xor U4674 (N_4674,N_4520,N_4583);
xor U4675 (N_4675,N_4589,N_4537);
nand U4676 (N_4676,N_4538,N_4506);
nor U4677 (N_4677,N_4535,N_4556);
nor U4678 (N_4678,N_4595,N_4544);
xor U4679 (N_4679,N_4592,N_4523);
nand U4680 (N_4680,N_4555,N_4534);
xnor U4681 (N_4681,N_4511,N_4570);
nor U4682 (N_4682,N_4554,N_4535);
xnor U4683 (N_4683,N_4598,N_4572);
nand U4684 (N_4684,N_4516,N_4529);
nand U4685 (N_4685,N_4584,N_4512);
nand U4686 (N_4686,N_4595,N_4591);
or U4687 (N_4687,N_4573,N_4558);
nor U4688 (N_4688,N_4579,N_4549);
or U4689 (N_4689,N_4527,N_4507);
or U4690 (N_4690,N_4501,N_4542);
and U4691 (N_4691,N_4531,N_4521);
and U4692 (N_4692,N_4579,N_4556);
nand U4693 (N_4693,N_4578,N_4520);
nand U4694 (N_4694,N_4579,N_4561);
xnor U4695 (N_4695,N_4515,N_4502);
xor U4696 (N_4696,N_4595,N_4543);
and U4697 (N_4697,N_4546,N_4574);
nand U4698 (N_4698,N_4599,N_4550);
and U4699 (N_4699,N_4587,N_4565);
and U4700 (N_4700,N_4691,N_4686);
or U4701 (N_4701,N_4605,N_4621);
or U4702 (N_4702,N_4600,N_4643);
xnor U4703 (N_4703,N_4601,N_4633);
or U4704 (N_4704,N_4679,N_4689);
nand U4705 (N_4705,N_4653,N_4667);
xor U4706 (N_4706,N_4680,N_4642);
and U4707 (N_4707,N_4619,N_4614);
or U4708 (N_4708,N_4675,N_4681);
or U4709 (N_4709,N_4629,N_4688);
xnor U4710 (N_4710,N_4668,N_4674);
nand U4711 (N_4711,N_4662,N_4692);
nand U4712 (N_4712,N_4671,N_4661);
nand U4713 (N_4713,N_4607,N_4659);
nor U4714 (N_4714,N_4682,N_4654);
nand U4715 (N_4715,N_4664,N_4648);
and U4716 (N_4716,N_4635,N_4641);
and U4717 (N_4717,N_4697,N_4604);
nor U4718 (N_4718,N_4602,N_4696);
nor U4719 (N_4719,N_4694,N_4656);
or U4720 (N_4720,N_4683,N_4612);
nor U4721 (N_4721,N_4631,N_4673);
nand U4722 (N_4722,N_4609,N_4672);
or U4723 (N_4723,N_4610,N_4620);
xnor U4724 (N_4724,N_4655,N_4639);
nor U4725 (N_4725,N_4634,N_4628);
nor U4726 (N_4726,N_4623,N_4644);
or U4727 (N_4727,N_4608,N_4693);
xnor U4728 (N_4728,N_4618,N_4676);
nor U4729 (N_4729,N_4622,N_4651);
xnor U4730 (N_4730,N_4665,N_4615);
xnor U4731 (N_4731,N_4632,N_4638);
or U4732 (N_4732,N_4606,N_4636);
nand U4733 (N_4733,N_4666,N_4637);
or U4734 (N_4734,N_4611,N_4616);
or U4735 (N_4735,N_4650,N_4678);
nand U4736 (N_4736,N_4663,N_4617);
and U4737 (N_4737,N_4677,N_4626);
nor U4738 (N_4738,N_4657,N_4685);
and U4739 (N_4739,N_4640,N_4645);
or U4740 (N_4740,N_4699,N_4652);
nor U4741 (N_4741,N_4669,N_4627);
nand U4742 (N_4742,N_4647,N_4684);
xor U4743 (N_4743,N_4658,N_4695);
nand U4744 (N_4744,N_4613,N_4649);
xor U4745 (N_4745,N_4698,N_4687);
and U4746 (N_4746,N_4630,N_4646);
or U4747 (N_4747,N_4625,N_4624);
nor U4748 (N_4748,N_4660,N_4690);
nor U4749 (N_4749,N_4670,N_4603);
xnor U4750 (N_4750,N_4660,N_4641);
nand U4751 (N_4751,N_4614,N_4648);
or U4752 (N_4752,N_4698,N_4606);
and U4753 (N_4753,N_4653,N_4630);
and U4754 (N_4754,N_4618,N_4680);
xor U4755 (N_4755,N_4613,N_4631);
or U4756 (N_4756,N_4671,N_4686);
or U4757 (N_4757,N_4622,N_4605);
nor U4758 (N_4758,N_4637,N_4656);
nor U4759 (N_4759,N_4665,N_4625);
and U4760 (N_4760,N_4675,N_4633);
xnor U4761 (N_4761,N_4607,N_4602);
xnor U4762 (N_4762,N_4632,N_4606);
and U4763 (N_4763,N_4606,N_4609);
nor U4764 (N_4764,N_4667,N_4652);
nor U4765 (N_4765,N_4611,N_4661);
nand U4766 (N_4766,N_4634,N_4662);
or U4767 (N_4767,N_4601,N_4665);
nand U4768 (N_4768,N_4626,N_4614);
and U4769 (N_4769,N_4695,N_4640);
nand U4770 (N_4770,N_4680,N_4600);
nor U4771 (N_4771,N_4600,N_4684);
xor U4772 (N_4772,N_4672,N_4666);
nand U4773 (N_4773,N_4624,N_4664);
nor U4774 (N_4774,N_4631,N_4647);
and U4775 (N_4775,N_4668,N_4698);
nand U4776 (N_4776,N_4679,N_4615);
and U4777 (N_4777,N_4626,N_4622);
nor U4778 (N_4778,N_4631,N_4617);
or U4779 (N_4779,N_4661,N_4616);
and U4780 (N_4780,N_4660,N_4633);
nor U4781 (N_4781,N_4664,N_4668);
or U4782 (N_4782,N_4657,N_4697);
and U4783 (N_4783,N_4628,N_4633);
nor U4784 (N_4784,N_4617,N_4657);
xnor U4785 (N_4785,N_4629,N_4658);
and U4786 (N_4786,N_4666,N_4636);
xnor U4787 (N_4787,N_4687,N_4636);
and U4788 (N_4788,N_4642,N_4628);
and U4789 (N_4789,N_4631,N_4663);
and U4790 (N_4790,N_4632,N_4611);
nand U4791 (N_4791,N_4630,N_4670);
xnor U4792 (N_4792,N_4687,N_4600);
nor U4793 (N_4793,N_4660,N_4695);
and U4794 (N_4794,N_4657,N_4695);
or U4795 (N_4795,N_4635,N_4628);
and U4796 (N_4796,N_4603,N_4614);
or U4797 (N_4797,N_4610,N_4658);
and U4798 (N_4798,N_4655,N_4696);
xor U4799 (N_4799,N_4632,N_4662);
xnor U4800 (N_4800,N_4763,N_4705);
nand U4801 (N_4801,N_4732,N_4710);
xnor U4802 (N_4802,N_4762,N_4795);
or U4803 (N_4803,N_4746,N_4715);
xor U4804 (N_4804,N_4794,N_4766);
nand U4805 (N_4805,N_4709,N_4725);
xnor U4806 (N_4806,N_4750,N_4720);
and U4807 (N_4807,N_4718,N_4755);
and U4808 (N_4808,N_4756,N_4702);
xor U4809 (N_4809,N_4784,N_4786);
and U4810 (N_4810,N_4799,N_4711);
nand U4811 (N_4811,N_4721,N_4776);
nor U4812 (N_4812,N_4708,N_4730);
or U4813 (N_4813,N_4714,N_4782);
nor U4814 (N_4814,N_4733,N_4744);
nand U4815 (N_4815,N_4764,N_4768);
or U4816 (N_4816,N_4792,N_4774);
or U4817 (N_4817,N_4728,N_4741);
and U4818 (N_4818,N_4781,N_4797);
nor U4819 (N_4819,N_4724,N_4749);
xnor U4820 (N_4820,N_4713,N_4751);
nand U4821 (N_4821,N_4701,N_4723);
and U4822 (N_4822,N_4747,N_4796);
or U4823 (N_4823,N_4735,N_4752);
or U4824 (N_4824,N_4717,N_4783);
nand U4825 (N_4825,N_4771,N_4760);
or U4826 (N_4826,N_4775,N_4780);
or U4827 (N_4827,N_4700,N_4704);
nand U4828 (N_4828,N_4719,N_4777);
and U4829 (N_4829,N_4745,N_4740);
and U4830 (N_4830,N_4790,N_4727);
nor U4831 (N_4831,N_4785,N_4742);
xnor U4832 (N_4832,N_4758,N_4753);
xnor U4833 (N_4833,N_4757,N_4729);
and U4834 (N_4834,N_4703,N_4706);
nand U4835 (N_4835,N_4789,N_4778);
or U4836 (N_4836,N_4754,N_4734);
or U4837 (N_4837,N_4739,N_4767);
nand U4838 (N_4838,N_4716,N_4793);
xor U4839 (N_4839,N_4712,N_4738);
nand U4840 (N_4840,N_4748,N_4788);
nor U4841 (N_4841,N_4787,N_4772);
and U4842 (N_4842,N_4736,N_4765);
or U4843 (N_4843,N_4761,N_4726);
nor U4844 (N_4844,N_4759,N_4773);
nand U4845 (N_4845,N_4707,N_4791);
nor U4846 (N_4846,N_4798,N_4769);
and U4847 (N_4847,N_4731,N_4770);
and U4848 (N_4848,N_4722,N_4779);
nand U4849 (N_4849,N_4743,N_4737);
or U4850 (N_4850,N_4793,N_4726);
nand U4851 (N_4851,N_4759,N_4714);
or U4852 (N_4852,N_4700,N_4799);
nand U4853 (N_4853,N_4784,N_4798);
nor U4854 (N_4854,N_4750,N_4781);
xor U4855 (N_4855,N_4796,N_4744);
and U4856 (N_4856,N_4744,N_4709);
nand U4857 (N_4857,N_4762,N_4746);
nand U4858 (N_4858,N_4734,N_4760);
nand U4859 (N_4859,N_4726,N_4732);
xor U4860 (N_4860,N_4723,N_4741);
xor U4861 (N_4861,N_4732,N_4753);
nor U4862 (N_4862,N_4791,N_4751);
nand U4863 (N_4863,N_4754,N_4726);
or U4864 (N_4864,N_4763,N_4700);
nor U4865 (N_4865,N_4752,N_4709);
xor U4866 (N_4866,N_4763,N_4754);
nand U4867 (N_4867,N_4729,N_4769);
xnor U4868 (N_4868,N_4781,N_4774);
nand U4869 (N_4869,N_4734,N_4777);
nor U4870 (N_4870,N_4740,N_4755);
or U4871 (N_4871,N_4769,N_4770);
or U4872 (N_4872,N_4781,N_4742);
xor U4873 (N_4873,N_4782,N_4734);
xor U4874 (N_4874,N_4722,N_4702);
and U4875 (N_4875,N_4746,N_4772);
and U4876 (N_4876,N_4767,N_4796);
or U4877 (N_4877,N_4745,N_4784);
nor U4878 (N_4878,N_4782,N_4768);
and U4879 (N_4879,N_4752,N_4714);
xnor U4880 (N_4880,N_4741,N_4720);
nor U4881 (N_4881,N_4713,N_4747);
or U4882 (N_4882,N_4727,N_4776);
xnor U4883 (N_4883,N_4761,N_4759);
nor U4884 (N_4884,N_4793,N_4762);
and U4885 (N_4885,N_4744,N_4753);
xor U4886 (N_4886,N_4717,N_4714);
nor U4887 (N_4887,N_4760,N_4742);
xnor U4888 (N_4888,N_4700,N_4789);
xnor U4889 (N_4889,N_4751,N_4764);
and U4890 (N_4890,N_4737,N_4764);
xor U4891 (N_4891,N_4724,N_4705);
xnor U4892 (N_4892,N_4735,N_4712);
and U4893 (N_4893,N_4704,N_4756);
or U4894 (N_4894,N_4747,N_4758);
nand U4895 (N_4895,N_4711,N_4765);
and U4896 (N_4896,N_4715,N_4758);
nor U4897 (N_4897,N_4703,N_4757);
or U4898 (N_4898,N_4799,N_4740);
xnor U4899 (N_4899,N_4751,N_4701);
nor U4900 (N_4900,N_4898,N_4829);
xnor U4901 (N_4901,N_4823,N_4882);
nor U4902 (N_4902,N_4869,N_4814);
nand U4903 (N_4903,N_4809,N_4802);
nand U4904 (N_4904,N_4819,N_4828);
nor U4905 (N_4905,N_4888,N_4889);
nor U4906 (N_4906,N_4807,N_4844);
nand U4907 (N_4907,N_4816,N_4868);
xnor U4908 (N_4908,N_4826,N_4866);
and U4909 (N_4909,N_4862,N_4840);
nand U4910 (N_4910,N_4871,N_4845);
xnor U4911 (N_4911,N_4812,N_4830);
nor U4912 (N_4912,N_4891,N_4800);
or U4913 (N_4913,N_4842,N_4880);
and U4914 (N_4914,N_4832,N_4856);
xnor U4915 (N_4915,N_4883,N_4804);
nand U4916 (N_4916,N_4808,N_4818);
nand U4917 (N_4917,N_4837,N_4876);
xor U4918 (N_4918,N_4879,N_4860);
nand U4919 (N_4919,N_4892,N_4849);
nor U4920 (N_4920,N_4850,N_4875);
and U4921 (N_4921,N_4897,N_4855);
and U4922 (N_4922,N_4824,N_4805);
or U4923 (N_4923,N_4896,N_4870);
xnor U4924 (N_4924,N_4803,N_4831);
or U4925 (N_4925,N_4827,N_4836);
or U4926 (N_4926,N_4885,N_4810);
nor U4927 (N_4927,N_4873,N_4801);
xor U4928 (N_4928,N_4874,N_4847);
nand U4929 (N_4929,N_4852,N_4887);
nand U4930 (N_4930,N_4858,N_4878);
and U4931 (N_4931,N_4863,N_4886);
and U4932 (N_4932,N_4839,N_4833);
xor U4933 (N_4933,N_4834,N_4815);
nor U4934 (N_4934,N_4854,N_4851);
or U4935 (N_4935,N_4811,N_4843);
nor U4936 (N_4936,N_4877,N_4838);
or U4937 (N_4937,N_4857,N_4820);
and U4938 (N_4938,N_4867,N_4864);
nor U4939 (N_4939,N_4872,N_4899);
nor U4940 (N_4940,N_4822,N_4861);
or U4941 (N_4941,N_4895,N_4806);
and U4942 (N_4942,N_4825,N_4813);
nor U4943 (N_4943,N_4848,N_4821);
and U4944 (N_4944,N_4853,N_4881);
nand U4945 (N_4945,N_4884,N_4865);
nand U4946 (N_4946,N_4894,N_4817);
nand U4947 (N_4947,N_4859,N_4893);
xnor U4948 (N_4948,N_4890,N_4841);
or U4949 (N_4949,N_4846,N_4835);
nor U4950 (N_4950,N_4833,N_4811);
xnor U4951 (N_4951,N_4863,N_4862);
and U4952 (N_4952,N_4865,N_4826);
nor U4953 (N_4953,N_4819,N_4804);
or U4954 (N_4954,N_4838,N_4824);
nand U4955 (N_4955,N_4872,N_4881);
or U4956 (N_4956,N_4831,N_4859);
and U4957 (N_4957,N_4816,N_4888);
xor U4958 (N_4958,N_4858,N_4839);
nor U4959 (N_4959,N_4837,N_4868);
or U4960 (N_4960,N_4897,N_4861);
nand U4961 (N_4961,N_4858,N_4834);
or U4962 (N_4962,N_4886,N_4838);
nand U4963 (N_4963,N_4836,N_4809);
nor U4964 (N_4964,N_4861,N_4800);
nand U4965 (N_4965,N_4886,N_4836);
nor U4966 (N_4966,N_4891,N_4881);
or U4967 (N_4967,N_4853,N_4820);
nand U4968 (N_4968,N_4812,N_4832);
nand U4969 (N_4969,N_4804,N_4805);
nor U4970 (N_4970,N_4812,N_4833);
xor U4971 (N_4971,N_4814,N_4891);
nand U4972 (N_4972,N_4803,N_4851);
nand U4973 (N_4973,N_4880,N_4816);
xnor U4974 (N_4974,N_4821,N_4875);
nand U4975 (N_4975,N_4828,N_4888);
or U4976 (N_4976,N_4826,N_4842);
nand U4977 (N_4977,N_4857,N_4883);
or U4978 (N_4978,N_4880,N_4853);
nor U4979 (N_4979,N_4868,N_4817);
and U4980 (N_4980,N_4898,N_4895);
or U4981 (N_4981,N_4824,N_4829);
or U4982 (N_4982,N_4820,N_4892);
or U4983 (N_4983,N_4818,N_4883);
xnor U4984 (N_4984,N_4844,N_4802);
or U4985 (N_4985,N_4840,N_4879);
or U4986 (N_4986,N_4816,N_4894);
nand U4987 (N_4987,N_4889,N_4897);
nand U4988 (N_4988,N_4833,N_4815);
xor U4989 (N_4989,N_4882,N_4810);
and U4990 (N_4990,N_4874,N_4895);
and U4991 (N_4991,N_4843,N_4897);
or U4992 (N_4992,N_4882,N_4829);
nor U4993 (N_4993,N_4800,N_4857);
nor U4994 (N_4994,N_4872,N_4871);
and U4995 (N_4995,N_4893,N_4871);
nand U4996 (N_4996,N_4857,N_4880);
nor U4997 (N_4997,N_4864,N_4895);
and U4998 (N_4998,N_4887,N_4838);
and U4999 (N_4999,N_4849,N_4833);
and U5000 (N_5000,N_4966,N_4942);
nor U5001 (N_5001,N_4980,N_4952);
xor U5002 (N_5002,N_4956,N_4964);
or U5003 (N_5003,N_4921,N_4957);
or U5004 (N_5004,N_4902,N_4955);
nand U5005 (N_5005,N_4915,N_4946);
nor U5006 (N_5006,N_4933,N_4978);
nand U5007 (N_5007,N_4989,N_4965);
and U5008 (N_5008,N_4958,N_4923);
and U5009 (N_5009,N_4941,N_4929);
and U5010 (N_5010,N_4983,N_4970);
xnor U5011 (N_5011,N_4960,N_4996);
nor U5012 (N_5012,N_4982,N_4976);
nand U5013 (N_5013,N_4934,N_4979);
xor U5014 (N_5014,N_4963,N_4943);
xnor U5015 (N_5015,N_4971,N_4917);
or U5016 (N_5016,N_4901,N_4939);
nor U5017 (N_5017,N_4999,N_4992);
nor U5018 (N_5018,N_4922,N_4977);
nand U5019 (N_5019,N_4916,N_4991);
xor U5020 (N_5020,N_4905,N_4994);
and U5021 (N_5021,N_4993,N_4973);
and U5022 (N_5022,N_4985,N_4906);
and U5023 (N_5023,N_4930,N_4926);
or U5024 (N_5024,N_4910,N_4904);
xor U5025 (N_5025,N_4932,N_4908);
nor U5026 (N_5026,N_4997,N_4953);
xor U5027 (N_5027,N_4907,N_4968);
xor U5028 (N_5028,N_4987,N_4945);
nand U5029 (N_5029,N_4924,N_4928);
and U5030 (N_5030,N_4951,N_4931);
or U5031 (N_5031,N_4974,N_4938);
nand U5032 (N_5032,N_4919,N_4984);
nand U5033 (N_5033,N_4936,N_4947);
nor U5034 (N_5034,N_4975,N_4914);
nor U5035 (N_5035,N_4986,N_4937);
nor U5036 (N_5036,N_4961,N_4940);
nor U5037 (N_5037,N_4912,N_4969);
nor U5038 (N_5038,N_4981,N_4988);
nor U5039 (N_5039,N_4935,N_4962);
xor U5040 (N_5040,N_4995,N_4972);
and U5041 (N_5041,N_4998,N_4954);
or U5042 (N_5042,N_4918,N_4948);
nand U5043 (N_5043,N_4950,N_4913);
nand U5044 (N_5044,N_4925,N_4949);
xnor U5045 (N_5045,N_4959,N_4967);
xnor U5046 (N_5046,N_4911,N_4903);
and U5047 (N_5047,N_4990,N_4900);
and U5048 (N_5048,N_4920,N_4944);
nand U5049 (N_5049,N_4909,N_4927);
xor U5050 (N_5050,N_4913,N_4976);
nor U5051 (N_5051,N_4983,N_4992);
and U5052 (N_5052,N_4998,N_4956);
or U5053 (N_5053,N_4981,N_4999);
nand U5054 (N_5054,N_4934,N_4976);
nor U5055 (N_5055,N_4939,N_4919);
and U5056 (N_5056,N_4930,N_4965);
nand U5057 (N_5057,N_4937,N_4904);
xor U5058 (N_5058,N_4956,N_4927);
nor U5059 (N_5059,N_4949,N_4961);
and U5060 (N_5060,N_4915,N_4925);
and U5061 (N_5061,N_4916,N_4922);
nand U5062 (N_5062,N_4916,N_4955);
xor U5063 (N_5063,N_4908,N_4976);
nand U5064 (N_5064,N_4930,N_4906);
nor U5065 (N_5065,N_4921,N_4932);
xnor U5066 (N_5066,N_4949,N_4919);
nand U5067 (N_5067,N_4987,N_4968);
xor U5068 (N_5068,N_4900,N_4939);
nor U5069 (N_5069,N_4954,N_4979);
nor U5070 (N_5070,N_4925,N_4928);
and U5071 (N_5071,N_4938,N_4901);
or U5072 (N_5072,N_4905,N_4940);
and U5073 (N_5073,N_4968,N_4986);
nand U5074 (N_5074,N_4941,N_4978);
nor U5075 (N_5075,N_4948,N_4925);
nor U5076 (N_5076,N_4920,N_4935);
nor U5077 (N_5077,N_4959,N_4915);
nor U5078 (N_5078,N_4949,N_4944);
nor U5079 (N_5079,N_4963,N_4964);
nor U5080 (N_5080,N_4965,N_4946);
xnor U5081 (N_5081,N_4970,N_4988);
nor U5082 (N_5082,N_4943,N_4929);
nor U5083 (N_5083,N_4973,N_4986);
nor U5084 (N_5084,N_4955,N_4901);
nand U5085 (N_5085,N_4913,N_4937);
and U5086 (N_5086,N_4997,N_4952);
or U5087 (N_5087,N_4946,N_4972);
and U5088 (N_5088,N_4900,N_4917);
and U5089 (N_5089,N_4910,N_4971);
or U5090 (N_5090,N_4927,N_4954);
and U5091 (N_5091,N_4967,N_4920);
xor U5092 (N_5092,N_4911,N_4910);
nand U5093 (N_5093,N_4945,N_4927);
nand U5094 (N_5094,N_4916,N_4928);
or U5095 (N_5095,N_4901,N_4953);
nor U5096 (N_5096,N_4998,N_4975);
xnor U5097 (N_5097,N_4952,N_4939);
or U5098 (N_5098,N_4906,N_4987);
nand U5099 (N_5099,N_4936,N_4994);
nand U5100 (N_5100,N_5031,N_5035);
xor U5101 (N_5101,N_5080,N_5017);
nor U5102 (N_5102,N_5028,N_5085);
or U5103 (N_5103,N_5030,N_5020);
or U5104 (N_5104,N_5060,N_5027);
xor U5105 (N_5105,N_5075,N_5001);
xor U5106 (N_5106,N_5018,N_5029);
or U5107 (N_5107,N_5051,N_5022);
nor U5108 (N_5108,N_5041,N_5052);
nand U5109 (N_5109,N_5086,N_5070);
nor U5110 (N_5110,N_5038,N_5087);
xnor U5111 (N_5111,N_5061,N_5074);
nor U5112 (N_5112,N_5068,N_5039);
nand U5113 (N_5113,N_5033,N_5096);
nor U5114 (N_5114,N_5088,N_5055);
and U5115 (N_5115,N_5092,N_5016);
xnor U5116 (N_5116,N_5079,N_5093);
nand U5117 (N_5117,N_5059,N_5047);
and U5118 (N_5118,N_5032,N_5083);
xor U5119 (N_5119,N_5019,N_5004);
nor U5120 (N_5120,N_5008,N_5062);
xor U5121 (N_5121,N_5036,N_5010);
and U5122 (N_5122,N_5044,N_5005);
nor U5123 (N_5123,N_5090,N_5026);
or U5124 (N_5124,N_5000,N_5056);
and U5125 (N_5125,N_5054,N_5012);
or U5126 (N_5126,N_5034,N_5024);
or U5127 (N_5127,N_5002,N_5037);
xor U5128 (N_5128,N_5042,N_5011);
nand U5129 (N_5129,N_5063,N_5007);
nor U5130 (N_5130,N_5006,N_5025);
and U5131 (N_5131,N_5099,N_5053);
nor U5132 (N_5132,N_5015,N_5089);
nor U5133 (N_5133,N_5014,N_5072);
nor U5134 (N_5134,N_5081,N_5066);
nand U5135 (N_5135,N_5043,N_5064);
nor U5136 (N_5136,N_5084,N_5009);
nand U5137 (N_5137,N_5098,N_5073);
or U5138 (N_5138,N_5021,N_5077);
nand U5139 (N_5139,N_5040,N_5094);
xor U5140 (N_5140,N_5048,N_5003);
and U5141 (N_5141,N_5023,N_5069);
and U5142 (N_5142,N_5095,N_5013);
and U5143 (N_5143,N_5091,N_5071);
nand U5144 (N_5144,N_5058,N_5046);
xnor U5145 (N_5145,N_5049,N_5057);
or U5146 (N_5146,N_5050,N_5067);
nor U5147 (N_5147,N_5065,N_5045);
xor U5148 (N_5148,N_5078,N_5076);
nand U5149 (N_5149,N_5082,N_5097);
xor U5150 (N_5150,N_5052,N_5031);
nor U5151 (N_5151,N_5092,N_5096);
or U5152 (N_5152,N_5056,N_5026);
nand U5153 (N_5153,N_5018,N_5051);
nor U5154 (N_5154,N_5054,N_5024);
and U5155 (N_5155,N_5065,N_5017);
or U5156 (N_5156,N_5076,N_5065);
nor U5157 (N_5157,N_5050,N_5099);
or U5158 (N_5158,N_5074,N_5068);
xnor U5159 (N_5159,N_5092,N_5070);
or U5160 (N_5160,N_5065,N_5042);
nand U5161 (N_5161,N_5052,N_5028);
and U5162 (N_5162,N_5027,N_5094);
nand U5163 (N_5163,N_5042,N_5037);
or U5164 (N_5164,N_5024,N_5090);
nor U5165 (N_5165,N_5001,N_5041);
nand U5166 (N_5166,N_5071,N_5043);
nor U5167 (N_5167,N_5064,N_5094);
xor U5168 (N_5168,N_5068,N_5098);
xor U5169 (N_5169,N_5049,N_5083);
nand U5170 (N_5170,N_5092,N_5060);
nor U5171 (N_5171,N_5075,N_5044);
nand U5172 (N_5172,N_5013,N_5075);
nor U5173 (N_5173,N_5010,N_5071);
xnor U5174 (N_5174,N_5064,N_5095);
or U5175 (N_5175,N_5040,N_5085);
nor U5176 (N_5176,N_5050,N_5010);
or U5177 (N_5177,N_5053,N_5043);
nand U5178 (N_5178,N_5055,N_5001);
and U5179 (N_5179,N_5021,N_5033);
xor U5180 (N_5180,N_5085,N_5066);
xor U5181 (N_5181,N_5042,N_5041);
and U5182 (N_5182,N_5016,N_5015);
xnor U5183 (N_5183,N_5056,N_5069);
nand U5184 (N_5184,N_5015,N_5027);
nor U5185 (N_5185,N_5071,N_5051);
or U5186 (N_5186,N_5033,N_5039);
nand U5187 (N_5187,N_5001,N_5030);
xnor U5188 (N_5188,N_5023,N_5030);
nand U5189 (N_5189,N_5023,N_5095);
and U5190 (N_5190,N_5055,N_5072);
and U5191 (N_5191,N_5082,N_5075);
xor U5192 (N_5192,N_5043,N_5083);
and U5193 (N_5193,N_5013,N_5017);
xnor U5194 (N_5194,N_5092,N_5026);
or U5195 (N_5195,N_5074,N_5040);
and U5196 (N_5196,N_5059,N_5076);
xor U5197 (N_5197,N_5093,N_5036);
xnor U5198 (N_5198,N_5026,N_5079);
or U5199 (N_5199,N_5036,N_5038);
nor U5200 (N_5200,N_5130,N_5103);
or U5201 (N_5201,N_5198,N_5156);
xor U5202 (N_5202,N_5100,N_5168);
or U5203 (N_5203,N_5163,N_5141);
nand U5204 (N_5204,N_5108,N_5137);
or U5205 (N_5205,N_5146,N_5197);
and U5206 (N_5206,N_5152,N_5110);
and U5207 (N_5207,N_5178,N_5169);
or U5208 (N_5208,N_5101,N_5188);
nor U5209 (N_5209,N_5116,N_5195);
xnor U5210 (N_5210,N_5155,N_5185);
nor U5211 (N_5211,N_5106,N_5128);
xnor U5212 (N_5212,N_5115,N_5118);
nor U5213 (N_5213,N_5111,N_5149);
and U5214 (N_5214,N_5181,N_5192);
nor U5215 (N_5215,N_5124,N_5142);
and U5216 (N_5216,N_5160,N_5186);
xnor U5217 (N_5217,N_5174,N_5113);
and U5218 (N_5218,N_5167,N_5132);
or U5219 (N_5219,N_5199,N_5157);
and U5220 (N_5220,N_5151,N_5102);
xnor U5221 (N_5221,N_5166,N_5161);
or U5222 (N_5222,N_5122,N_5171);
and U5223 (N_5223,N_5121,N_5193);
and U5224 (N_5224,N_5140,N_5190);
or U5225 (N_5225,N_5144,N_5120);
xor U5226 (N_5226,N_5127,N_5196);
nor U5227 (N_5227,N_5175,N_5117);
xnor U5228 (N_5228,N_5154,N_5125);
xnor U5229 (N_5229,N_5172,N_5147);
and U5230 (N_5230,N_5173,N_5123);
xor U5231 (N_5231,N_5126,N_5129);
or U5232 (N_5232,N_5150,N_5135);
xor U5233 (N_5233,N_5143,N_5119);
xor U5234 (N_5234,N_5134,N_5162);
nor U5235 (N_5235,N_5165,N_5145);
xnor U5236 (N_5236,N_5138,N_5109);
nand U5237 (N_5237,N_5105,N_5107);
and U5238 (N_5238,N_5189,N_5177);
nand U5239 (N_5239,N_5170,N_5180);
nor U5240 (N_5240,N_5148,N_5159);
and U5241 (N_5241,N_5133,N_5104);
nand U5242 (N_5242,N_5136,N_5112);
nor U5243 (N_5243,N_5158,N_5187);
or U5244 (N_5244,N_5131,N_5164);
nand U5245 (N_5245,N_5183,N_5191);
xor U5246 (N_5246,N_5179,N_5139);
nor U5247 (N_5247,N_5194,N_5182);
nor U5248 (N_5248,N_5114,N_5153);
or U5249 (N_5249,N_5176,N_5184);
nand U5250 (N_5250,N_5129,N_5156);
nor U5251 (N_5251,N_5182,N_5172);
nor U5252 (N_5252,N_5186,N_5150);
nand U5253 (N_5253,N_5182,N_5123);
nor U5254 (N_5254,N_5192,N_5120);
nor U5255 (N_5255,N_5151,N_5185);
nor U5256 (N_5256,N_5180,N_5137);
xor U5257 (N_5257,N_5119,N_5190);
and U5258 (N_5258,N_5122,N_5169);
xor U5259 (N_5259,N_5176,N_5160);
nor U5260 (N_5260,N_5197,N_5189);
nand U5261 (N_5261,N_5138,N_5105);
or U5262 (N_5262,N_5119,N_5185);
or U5263 (N_5263,N_5111,N_5110);
or U5264 (N_5264,N_5178,N_5109);
and U5265 (N_5265,N_5140,N_5129);
or U5266 (N_5266,N_5123,N_5153);
nand U5267 (N_5267,N_5162,N_5126);
nand U5268 (N_5268,N_5111,N_5154);
xnor U5269 (N_5269,N_5198,N_5142);
nor U5270 (N_5270,N_5122,N_5145);
xor U5271 (N_5271,N_5120,N_5111);
and U5272 (N_5272,N_5127,N_5198);
nor U5273 (N_5273,N_5124,N_5164);
nor U5274 (N_5274,N_5101,N_5159);
and U5275 (N_5275,N_5128,N_5182);
and U5276 (N_5276,N_5144,N_5157);
or U5277 (N_5277,N_5157,N_5177);
or U5278 (N_5278,N_5193,N_5166);
xor U5279 (N_5279,N_5199,N_5164);
or U5280 (N_5280,N_5196,N_5161);
nor U5281 (N_5281,N_5162,N_5194);
nand U5282 (N_5282,N_5104,N_5129);
and U5283 (N_5283,N_5195,N_5172);
nor U5284 (N_5284,N_5100,N_5163);
nand U5285 (N_5285,N_5139,N_5153);
nor U5286 (N_5286,N_5198,N_5158);
and U5287 (N_5287,N_5155,N_5102);
nor U5288 (N_5288,N_5119,N_5123);
nor U5289 (N_5289,N_5198,N_5124);
and U5290 (N_5290,N_5165,N_5183);
nand U5291 (N_5291,N_5163,N_5196);
xor U5292 (N_5292,N_5103,N_5179);
nand U5293 (N_5293,N_5142,N_5146);
xor U5294 (N_5294,N_5164,N_5184);
xnor U5295 (N_5295,N_5188,N_5142);
and U5296 (N_5296,N_5199,N_5100);
or U5297 (N_5297,N_5101,N_5191);
nand U5298 (N_5298,N_5137,N_5144);
nor U5299 (N_5299,N_5177,N_5197);
xnor U5300 (N_5300,N_5241,N_5294);
xnor U5301 (N_5301,N_5268,N_5282);
nor U5302 (N_5302,N_5217,N_5206);
nand U5303 (N_5303,N_5293,N_5233);
xor U5304 (N_5304,N_5259,N_5290);
nand U5305 (N_5305,N_5284,N_5269);
nor U5306 (N_5306,N_5248,N_5239);
nand U5307 (N_5307,N_5225,N_5208);
nand U5308 (N_5308,N_5234,N_5237);
nand U5309 (N_5309,N_5264,N_5204);
or U5310 (N_5310,N_5212,N_5275);
xor U5311 (N_5311,N_5280,N_5283);
nand U5312 (N_5312,N_5292,N_5276);
nor U5313 (N_5313,N_5267,N_5229);
nor U5314 (N_5314,N_5246,N_5270);
nor U5315 (N_5315,N_5203,N_5257);
and U5316 (N_5316,N_5281,N_5299);
xnor U5317 (N_5317,N_5228,N_5291);
nor U5318 (N_5318,N_5289,N_5297);
or U5319 (N_5319,N_5249,N_5211);
or U5320 (N_5320,N_5263,N_5236);
nor U5321 (N_5321,N_5260,N_5202);
nand U5322 (N_5322,N_5286,N_5273);
and U5323 (N_5323,N_5232,N_5254);
nand U5324 (N_5324,N_5278,N_5222);
and U5325 (N_5325,N_5209,N_5230);
or U5326 (N_5326,N_5256,N_5218);
or U5327 (N_5327,N_5287,N_5272);
nor U5328 (N_5328,N_5296,N_5295);
xnor U5329 (N_5329,N_5223,N_5244);
xor U5330 (N_5330,N_5240,N_5265);
or U5331 (N_5331,N_5235,N_5215);
nor U5332 (N_5332,N_5226,N_5262);
xor U5333 (N_5333,N_5252,N_5227);
and U5334 (N_5334,N_5205,N_5245);
and U5335 (N_5335,N_5247,N_5261);
and U5336 (N_5336,N_5219,N_5266);
and U5337 (N_5337,N_5251,N_5279);
nor U5338 (N_5338,N_5277,N_5224);
or U5339 (N_5339,N_5213,N_5214);
or U5340 (N_5340,N_5242,N_5210);
xnor U5341 (N_5341,N_5271,N_5221);
or U5342 (N_5342,N_5288,N_5274);
xor U5343 (N_5343,N_5285,N_5200);
xnor U5344 (N_5344,N_5250,N_5207);
or U5345 (N_5345,N_5220,N_5255);
or U5346 (N_5346,N_5231,N_5253);
nor U5347 (N_5347,N_5238,N_5216);
nor U5348 (N_5348,N_5258,N_5201);
or U5349 (N_5349,N_5298,N_5243);
xnor U5350 (N_5350,N_5211,N_5214);
or U5351 (N_5351,N_5263,N_5294);
nand U5352 (N_5352,N_5266,N_5286);
nor U5353 (N_5353,N_5289,N_5215);
or U5354 (N_5354,N_5205,N_5277);
and U5355 (N_5355,N_5219,N_5292);
xor U5356 (N_5356,N_5262,N_5272);
xor U5357 (N_5357,N_5202,N_5257);
or U5358 (N_5358,N_5243,N_5281);
nor U5359 (N_5359,N_5215,N_5248);
and U5360 (N_5360,N_5297,N_5274);
or U5361 (N_5361,N_5264,N_5206);
nand U5362 (N_5362,N_5204,N_5297);
nor U5363 (N_5363,N_5230,N_5216);
nor U5364 (N_5364,N_5275,N_5250);
and U5365 (N_5365,N_5203,N_5273);
or U5366 (N_5366,N_5256,N_5203);
nor U5367 (N_5367,N_5290,N_5216);
nand U5368 (N_5368,N_5285,N_5266);
or U5369 (N_5369,N_5239,N_5256);
or U5370 (N_5370,N_5207,N_5282);
nand U5371 (N_5371,N_5200,N_5228);
nor U5372 (N_5372,N_5251,N_5275);
xor U5373 (N_5373,N_5201,N_5221);
and U5374 (N_5374,N_5218,N_5257);
xor U5375 (N_5375,N_5283,N_5268);
and U5376 (N_5376,N_5294,N_5227);
nand U5377 (N_5377,N_5218,N_5217);
nor U5378 (N_5378,N_5250,N_5294);
and U5379 (N_5379,N_5232,N_5264);
nor U5380 (N_5380,N_5244,N_5229);
nand U5381 (N_5381,N_5283,N_5264);
xnor U5382 (N_5382,N_5280,N_5213);
xor U5383 (N_5383,N_5201,N_5288);
nand U5384 (N_5384,N_5246,N_5299);
nand U5385 (N_5385,N_5225,N_5257);
nor U5386 (N_5386,N_5209,N_5292);
or U5387 (N_5387,N_5226,N_5261);
xnor U5388 (N_5388,N_5291,N_5213);
xnor U5389 (N_5389,N_5289,N_5283);
or U5390 (N_5390,N_5277,N_5270);
xnor U5391 (N_5391,N_5287,N_5280);
or U5392 (N_5392,N_5210,N_5283);
xnor U5393 (N_5393,N_5231,N_5298);
xnor U5394 (N_5394,N_5224,N_5268);
nand U5395 (N_5395,N_5289,N_5260);
nor U5396 (N_5396,N_5267,N_5270);
nand U5397 (N_5397,N_5260,N_5238);
and U5398 (N_5398,N_5245,N_5210);
or U5399 (N_5399,N_5259,N_5204);
nor U5400 (N_5400,N_5335,N_5366);
nand U5401 (N_5401,N_5336,N_5394);
xor U5402 (N_5402,N_5332,N_5316);
nor U5403 (N_5403,N_5352,N_5387);
xnor U5404 (N_5404,N_5398,N_5307);
or U5405 (N_5405,N_5383,N_5347);
and U5406 (N_5406,N_5311,N_5369);
xor U5407 (N_5407,N_5393,N_5370);
or U5408 (N_5408,N_5381,N_5360);
or U5409 (N_5409,N_5323,N_5331);
nand U5410 (N_5410,N_5382,N_5399);
and U5411 (N_5411,N_5374,N_5353);
xnor U5412 (N_5412,N_5378,N_5300);
and U5413 (N_5413,N_5385,N_5379);
and U5414 (N_5414,N_5373,N_5319);
xor U5415 (N_5415,N_5351,N_5337);
and U5416 (N_5416,N_5339,N_5356);
and U5417 (N_5417,N_5318,N_5392);
nand U5418 (N_5418,N_5341,N_5397);
or U5419 (N_5419,N_5348,N_5340);
or U5420 (N_5420,N_5380,N_5358);
nor U5421 (N_5421,N_5312,N_5302);
and U5422 (N_5422,N_5343,N_5303);
xnor U5423 (N_5423,N_5390,N_5367);
xnor U5424 (N_5424,N_5362,N_5342);
nor U5425 (N_5425,N_5327,N_5376);
and U5426 (N_5426,N_5364,N_5355);
nor U5427 (N_5427,N_5354,N_5375);
nor U5428 (N_5428,N_5396,N_5330);
or U5429 (N_5429,N_5322,N_5344);
or U5430 (N_5430,N_5328,N_5301);
nand U5431 (N_5431,N_5377,N_5315);
nand U5432 (N_5432,N_5326,N_5384);
nand U5433 (N_5433,N_5388,N_5372);
nor U5434 (N_5434,N_5305,N_5371);
and U5435 (N_5435,N_5368,N_5314);
or U5436 (N_5436,N_5346,N_5324);
nor U5437 (N_5437,N_5321,N_5349);
and U5438 (N_5438,N_5350,N_5304);
nand U5439 (N_5439,N_5310,N_5313);
xnor U5440 (N_5440,N_5325,N_5361);
and U5441 (N_5441,N_5345,N_5317);
nand U5442 (N_5442,N_5359,N_5391);
xor U5443 (N_5443,N_5333,N_5320);
and U5444 (N_5444,N_5329,N_5308);
and U5445 (N_5445,N_5306,N_5334);
and U5446 (N_5446,N_5395,N_5386);
or U5447 (N_5447,N_5357,N_5363);
and U5448 (N_5448,N_5389,N_5309);
and U5449 (N_5449,N_5338,N_5365);
xnor U5450 (N_5450,N_5339,N_5317);
xnor U5451 (N_5451,N_5349,N_5329);
nor U5452 (N_5452,N_5356,N_5355);
nand U5453 (N_5453,N_5385,N_5317);
or U5454 (N_5454,N_5378,N_5321);
nand U5455 (N_5455,N_5321,N_5335);
nand U5456 (N_5456,N_5397,N_5366);
nand U5457 (N_5457,N_5343,N_5324);
or U5458 (N_5458,N_5312,N_5310);
nand U5459 (N_5459,N_5389,N_5320);
nor U5460 (N_5460,N_5392,N_5337);
xor U5461 (N_5461,N_5315,N_5382);
and U5462 (N_5462,N_5335,N_5374);
xnor U5463 (N_5463,N_5360,N_5394);
xor U5464 (N_5464,N_5327,N_5335);
nand U5465 (N_5465,N_5307,N_5364);
nor U5466 (N_5466,N_5308,N_5349);
and U5467 (N_5467,N_5378,N_5361);
or U5468 (N_5468,N_5386,N_5306);
nand U5469 (N_5469,N_5332,N_5327);
xnor U5470 (N_5470,N_5334,N_5347);
or U5471 (N_5471,N_5311,N_5380);
and U5472 (N_5472,N_5342,N_5344);
nand U5473 (N_5473,N_5358,N_5304);
or U5474 (N_5474,N_5362,N_5306);
and U5475 (N_5475,N_5329,N_5392);
nand U5476 (N_5476,N_5360,N_5374);
nor U5477 (N_5477,N_5303,N_5365);
nand U5478 (N_5478,N_5306,N_5367);
nor U5479 (N_5479,N_5397,N_5380);
or U5480 (N_5480,N_5342,N_5311);
xnor U5481 (N_5481,N_5341,N_5318);
and U5482 (N_5482,N_5350,N_5311);
nand U5483 (N_5483,N_5325,N_5304);
xor U5484 (N_5484,N_5374,N_5385);
or U5485 (N_5485,N_5344,N_5396);
and U5486 (N_5486,N_5348,N_5381);
nand U5487 (N_5487,N_5302,N_5327);
and U5488 (N_5488,N_5325,N_5321);
or U5489 (N_5489,N_5377,N_5317);
nand U5490 (N_5490,N_5376,N_5398);
and U5491 (N_5491,N_5350,N_5354);
or U5492 (N_5492,N_5354,N_5310);
and U5493 (N_5493,N_5396,N_5347);
nor U5494 (N_5494,N_5397,N_5314);
xnor U5495 (N_5495,N_5394,N_5390);
xnor U5496 (N_5496,N_5360,N_5393);
xor U5497 (N_5497,N_5372,N_5317);
and U5498 (N_5498,N_5365,N_5305);
or U5499 (N_5499,N_5371,N_5302);
or U5500 (N_5500,N_5442,N_5449);
nor U5501 (N_5501,N_5489,N_5448);
or U5502 (N_5502,N_5440,N_5461);
xnor U5503 (N_5503,N_5410,N_5480);
or U5504 (N_5504,N_5457,N_5486);
nor U5505 (N_5505,N_5444,N_5427);
nor U5506 (N_5506,N_5418,N_5411);
nor U5507 (N_5507,N_5426,N_5409);
xnor U5508 (N_5508,N_5490,N_5481);
nand U5509 (N_5509,N_5441,N_5416);
xor U5510 (N_5510,N_5436,N_5434);
and U5511 (N_5511,N_5472,N_5478);
nor U5512 (N_5512,N_5432,N_5484);
nand U5513 (N_5513,N_5403,N_5494);
and U5514 (N_5514,N_5487,N_5459);
or U5515 (N_5515,N_5443,N_5401);
xnor U5516 (N_5516,N_5477,N_5460);
and U5517 (N_5517,N_5473,N_5419);
or U5518 (N_5518,N_5458,N_5420);
xor U5519 (N_5519,N_5479,N_5445);
nand U5520 (N_5520,N_5452,N_5464);
and U5521 (N_5521,N_5400,N_5496);
and U5522 (N_5522,N_5470,N_5433);
nand U5523 (N_5523,N_5485,N_5468);
and U5524 (N_5524,N_5471,N_5437);
nand U5525 (N_5525,N_5431,N_5498);
xnor U5526 (N_5526,N_5404,N_5451);
xor U5527 (N_5527,N_5421,N_5466);
nand U5528 (N_5528,N_5492,N_5454);
and U5529 (N_5529,N_5497,N_5424);
nand U5530 (N_5530,N_5413,N_5462);
nor U5531 (N_5531,N_5430,N_5435);
nand U5532 (N_5532,N_5455,N_5422);
nand U5533 (N_5533,N_5488,N_5463);
nand U5534 (N_5534,N_5453,N_5475);
nor U5535 (N_5535,N_5456,N_5450);
and U5536 (N_5536,N_5438,N_5493);
xor U5537 (N_5537,N_5467,N_5482);
nand U5538 (N_5538,N_5428,N_5446);
and U5539 (N_5539,N_5447,N_5408);
nand U5540 (N_5540,N_5469,N_5407);
nand U5541 (N_5541,N_5499,N_5402);
xor U5542 (N_5542,N_5474,N_5412);
and U5543 (N_5543,N_5423,N_5405);
xor U5544 (N_5544,N_5425,N_5429);
nor U5545 (N_5545,N_5483,N_5439);
and U5546 (N_5546,N_5491,N_5417);
xor U5547 (N_5547,N_5465,N_5495);
xnor U5548 (N_5548,N_5414,N_5476);
nand U5549 (N_5549,N_5406,N_5415);
nor U5550 (N_5550,N_5445,N_5417);
nand U5551 (N_5551,N_5482,N_5418);
and U5552 (N_5552,N_5462,N_5403);
nand U5553 (N_5553,N_5452,N_5442);
nand U5554 (N_5554,N_5407,N_5462);
nand U5555 (N_5555,N_5443,N_5467);
and U5556 (N_5556,N_5467,N_5497);
or U5557 (N_5557,N_5475,N_5467);
xor U5558 (N_5558,N_5404,N_5418);
nand U5559 (N_5559,N_5499,N_5434);
or U5560 (N_5560,N_5405,N_5439);
nor U5561 (N_5561,N_5491,N_5481);
nand U5562 (N_5562,N_5414,N_5499);
or U5563 (N_5563,N_5412,N_5475);
or U5564 (N_5564,N_5491,N_5467);
nand U5565 (N_5565,N_5445,N_5433);
nand U5566 (N_5566,N_5430,N_5444);
nand U5567 (N_5567,N_5429,N_5443);
nand U5568 (N_5568,N_5489,N_5429);
nor U5569 (N_5569,N_5461,N_5421);
xor U5570 (N_5570,N_5432,N_5478);
nor U5571 (N_5571,N_5405,N_5400);
xor U5572 (N_5572,N_5494,N_5451);
and U5573 (N_5573,N_5451,N_5426);
and U5574 (N_5574,N_5499,N_5437);
nand U5575 (N_5575,N_5402,N_5455);
nor U5576 (N_5576,N_5446,N_5451);
nor U5577 (N_5577,N_5402,N_5403);
xor U5578 (N_5578,N_5422,N_5419);
nand U5579 (N_5579,N_5403,N_5486);
nand U5580 (N_5580,N_5441,N_5438);
or U5581 (N_5581,N_5431,N_5429);
and U5582 (N_5582,N_5440,N_5432);
xnor U5583 (N_5583,N_5445,N_5457);
xor U5584 (N_5584,N_5447,N_5425);
nor U5585 (N_5585,N_5470,N_5493);
nor U5586 (N_5586,N_5461,N_5480);
or U5587 (N_5587,N_5457,N_5467);
nand U5588 (N_5588,N_5448,N_5492);
nand U5589 (N_5589,N_5428,N_5499);
and U5590 (N_5590,N_5445,N_5467);
or U5591 (N_5591,N_5474,N_5407);
nor U5592 (N_5592,N_5424,N_5419);
and U5593 (N_5593,N_5419,N_5472);
and U5594 (N_5594,N_5461,N_5447);
xor U5595 (N_5595,N_5435,N_5466);
or U5596 (N_5596,N_5477,N_5456);
xnor U5597 (N_5597,N_5433,N_5432);
or U5598 (N_5598,N_5467,N_5429);
and U5599 (N_5599,N_5476,N_5498);
nor U5600 (N_5600,N_5596,N_5528);
nand U5601 (N_5601,N_5598,N_5549);
xnor U5602 (N_5602,N_5560,N_5500);
xor U5603 (N_5603,N_5512,N_5526);
nor U5604 (N_5604,N_5561,N_5573);
xnor U5605 (N_5605,N_5548,N_5590);
xor U5606 (N_5606,N_5542,N_5577);
and U5607 (N_5607,N_5505,N_5517);
nor U5608 (N_5608,N_5525,N_5541);
nor U5609 (N_5609,N_5545,N_5572);
and U5610 (N_5610,N_5556,N_5565);
xnor U5611 (N_5611,N_5588,N_5570);
and U5612 (N_5612,N_5597,N_5569);
nor U5613 (N_5613,N_5584,N_5532);
or U5614 (N_5614,N_5571,N_5510);
xnor U5615 (N_5615,N_5520,N_5537);
or U5616 (N_5616,N_5594,N_5575);
xnor U5617 (N_5617,N_5523,N_5566);
or U5618 (N_5618,N_5511,N_5557);
and U5619 (N_5619,N_5589,N_5585);
and U5620 (N_5620,N_5579,N_5568);
nand U5621 (N_5621,N_5564,N_5533);
xnor U5622 (N_5622,N_5546,N_5527);
nor U5623 (N_5623,N_5536,N_5580);
and U5624 (N_5624,N_5543,N_5501);
nand U5625 (N_5625,N_5554,N_5553);
nor U5626 (N_5626,N_5529,N_5519);
or U5627 (N_5627,N_5531,N_5583);
nand U5628 (N_5628,N_5516,N_5586);
nor U5629 (N_5629,N_5524,N_5518);
and U5630 (N_5630,N_5559,N_5555);
nor U5631 (N_5631,N_5550,N_5509);
nor U5632 (N_5632,N_5574,N_5578);
and U5633 (N_5633,N_5540,N_5558);
xnor U5634 (N_5634,N_5507,N_5581);
and U5635 (N_5635,N_5515,N_5534);
nand U5636 (N_5636,N_5593,N_5567);
or U5637 (N_5637,N_5535,N_5591);
nor U5638 (N_5638,N_5506,N_5551);
nor U5639 (N_5639,N_5552,N_5539);
nor U5640 (N_5640,N_5502,N_5503);
and U5641 (N_5641,N_5538,N_5544);
xor U5642 (N_5642,N_5521,N_5522);
or U5643 (N_5643,N_5582,N_5599);
nand U5644 (N_5644,N_5595,N_5508);
nor U5645 (N_5645,N_5587,N_5514);
nand U5646 (N_5646,N_5504,N_5592);
nand U5647 (N_5647,N_5530,N_5547);
nor U5648 (N_5648,N_5576,N_5563);
nor U5649 (N_5649,N_5513,N_5562);
nand U5650 (N_5650,N_5525,N_5524);
xor U5651 (N_5651,N_5521,N_5564);
nor U5652 (N_5652,N_5564,N_5508);
nor U5653 (N_5653,N_5569,N_5552);
nand U5654 (N_5654,N_5581,N_5597);
nand U5655 (N_5655,N_5546,N_5571);
or U5656 (N_5656,N_5555,N_5547);
and U5657 (N_5657,N_5516,N_5532);
and U5658 (N_5658,N_5533,N_5571);
or U5659 (N_5659,N_5500,N_5568);
nor U5660 (N_5660,N_5547,N_5509);
or U5661 (N_5661,N_5579,N_5599);
xnor U5662 (N_5662,N_5588,N_5526);
nand U5663 (N_5663,N_5501,N_5588);
xor U5664 (N_5664,N_5534,N_5532);
nand U5665 (N_5665,N_5513,N_5502);
and U5666 (N_5666,N_5524,N_5527);
and U5667 (N_5667,N_5582,N_5548);
or U5668 (N_5668,N_5513,N_5525);
or U5669 (N_5669,N_5571,N_5500);
nand U5670 (N_5670,N_5557,N_5544);
and U5671 (N_5671,N_5512,N_5575);
nor U5672 (N_5672,N_5571,N_5531);
nand U5673 (N_5673,N_5592,N_5516);
xor U5674 (N_5674,N_5594,N_5547);
xor U5675 (N_5675,N_5569,N_5514);
nor U5676 (N_5676,N_5514,N_5548);
xnor U5677 (N_5677,N_5531,N_5576);
and U5678 (N_5678,N_5599,N_5592);
and U5679 (N_5679,N_5577,N_5540);
or U5680 (N_5680,N_5587,N_5517);
or U5681 (N_5681,N_5570,N_5511);
or U5682 (N_5682,N_5543,N_5578);
xor U5683 (N_5683,N_5561,N_5558);
nor U5684 (N_5684,N_5505,N_5550);
nor U5685 (N_5685,N_5595,N_5552);
xnor U5686 (N_5686,N_5517,N_5531);
and U5687 (N_5687,N_5581,N_5524);
xnor U5688 (N_5688,N_5501,N_5534);
xor U5689 (N_5689,N_5566,N_5541);
or U5690 (N_5690,N_5597,N_5515);
nand U5691 (N_5691,N_5526,N_5549);
nand U5692 (N_5692,N_5564,N_5581);
nor U5693 (N_5693,N_5504,N_5546);
and U5694 (N_5694,N_5565,N_5597);
nand U5695 (N_5695,N_5598,N_5504);
nand U5696 (N_5696,N_5564,N_5544);
nand U5697 (N_5697,N_5516,N_5519);
or U5698 (N_5698,N_5581,N_5506);
nand U5699 (N_5699,N_5541,N_5542);
nand U5700 (N_5700,N_5638,N_5612);
xnor U5701 (N_5701,N_5630,N_5695);
nor U5702 (N_5702,N_5605,N_5661);
xnor U5703 (N_5703,N_5604,N_5634);
and U5704 (N_5704,N_5696,N_5650);
and U5705 (N_5705,N_5639,N_5635);
and U5706 (N_5706,N_5671,N_5640);
or U5707 (N_5707,N_5675,N_5690);
or U5708 (N_5708,N_5645,N_5656);
nand U5709 (N_5709,N_5608,N_5678);
and U5710 (N_5710,N_5633,N_5619);
nand U5711 (N_5711,N_5667,N_5603);
and U5712 (N_5712,N_5688,N_5629);
and U5713 (N_5713,N_5646,N_5669);
or U5714 (N_5714,N_5672,N_5610);
and U5715 (N_5715,N_5674,N_5680);
nor U5716 (N_5716,N_5673,N_5659);
nor U5717 (N_5717,N_5648,N_5644);
or U5718 (N_5718,N_5668,N_5681);
xor U5719 (N_5719,N_5643,N_5607);
or U5720 (N_5720,N_5621,N_5662);
nor U5721 (N_5721,N_5683,N_5677);
nand U5722 (N_5722,N_5697,N_5657);
nand U5723 (N_5723,N_5622,N_5686);
xor U5724 (N_5724,N_5637,N_5628);
xnor U5725 (N_5725,N_5664,N_5693);
xnor U5726 (N_5726,N_5620,N_5615);
nor U5727 (N_5727,N_5684,N_5609);
nand U5728 (N_5728,N_5606,N_5647);
nand U5729 (N_5729,N_5685,N_5655);
and U5730 (N_5730,N_5698,N_5676);
and U5731 (N_5731,N_5692,N_5602);
nand U5732 (N_5732,N_5649,N_5689);
or U5733 (N_5733,N_5666,N_5600);
or U5734 (N_5734,N_5663,N_5687);
or U5735 (N_5735,N_5611,N_5632);
nor U5736 (N_5736,N_5641,N_5682);
nand U5737 (N_5737,N_5651,N_5694);
and U5738 (N_5738,N_5624,N_5654);
and U5739 (N_5739,N_5617,N_5660);
nor U5740 (N_5740,N_5601,N_5665);
or U5741 (N_5741,N_5658,N_5642);
and U5742 (N_5742,N_5627,N_5691);
or U5743 (N_5743,N_5670,N_5679);
nand U5744 (N_5744,N_5623,N_5614);
and U5745 (N_5745,N_5618,N_5626);
xnor U5746 (N_5746,N_5631,N_5653);
and U5747 (N_5747,N_5613,N_5625);
or U5748 (N_5748,N_5636,N_5652);
nor U5749 (N_5749,N_5616,N_5699);
and U5750 (N_5750,N_5680,N_5658);
and U5751 (N_5751,N_5686,N_5643);
or U5752 (N_5752,N_5630,N_5655);
and U5753 (N_5753,N_5642,N_5697);
nor U5754 (N_5754,N_5698,N_5664);
xnor U5755 (N_5755,N_5623,N_5681);
and U5756 (N_5756,N_5638,N_5621);
nand U5757 (N_5757,N_5687,N_5649);
and U5758 (N_5758,N_5622,N_5608);
and U5759 (N_5759,N_5632,N_5601);
or U5760 (N_5760,N_5663,N_5639);
nand U5761 (N_5761,N_5688,N_5695);
xnor U5762 (N_5762,N_5684,N_5687);
xnor U5763 (N_5763,N_5605,N_5626);
and U5764 (N_5764,N_5666,N_5636);
and U5765 (N_5765,N_5633,N_5648);
nor U5766 (N_5766,N_5671,N_5693);
xor U5767 (N_5767,N_5656,N_5652);
and U5768 (N_5768,N_5671,N_5696);
xnor U5769 (N_5769,N_5682,N_5690);
and U5770 (N_5770,N_5615,N_5617);
nor U5771 (N_5771,N_5663,N_5697);
nand U5772 (N_5772,N_5642,N_5614);
or U5773 (N_5773,N_5687,N_5619);
and U5774 (N_5774,N_5696,N_5629);
and U5775 (N_5775,N_5603,N_5620);
nand U5776 (N_5776,N_5624,N_5619);
and U5777 (N_5777,N_5621,N_5687);
xnor U5778 (N_5778,N_5608,N_5627);
xnor U5779 (N_5779,N_5692,N_5687);
or U5780 (N_5780,N_5649,N_5620);
xor U5781 (N_5781,N_5699,N_5617);
or U5782 (N_5782,N_5676,N_5624);
and U5783 (N_5783,N_5696,N_5633);
and U5784 (N_5784,N_5677,N_5642);
or U5785 (N_5785,N_5664,N_5638);
nor U5786 (N_5786,N_5682,N_5614);
nand U5787 (N_5787,N_5671,N_5660);
nand U5788 (N_5788,N_5639,N_5696);
nand U5789 (N_5789,N_5634,N_5643);
and U5790 (N_5790,N_5664,N_5617);
or U5791 (N_5791,N_5697,N_5600);
and U5792 (N_5792,N_5645,N_5663);
or U5793 (N_5793,N_5611,N_5672);
nand U5794 (N_5794,N_5691,N_5604);
xnor U5795 (N_5795,N_5654,N_5650);
xor U5796 (N_5796,N_5651,N_5678);
and U5797 (N_5797,N_5673,N_5602);
or U5798 (N_5798,N_5655,N_5627);
xnor U5799 (N_5799,N_5648,N_5601);
nor U5800 (N_5800,N_5768,N_5720);
xnor U5801 (N_5801,N_5739,N_5722);
nand U5802 (N_5802,N_5742,N_5705);
nor U5803 (N_5803,N_5712,N_5776);
nand U5804 (N_5804,N_5732,N_5747);
or U5805 (N_5805,N_5799,N_5758);
nand U5806 (N_5806,N_5736,N_5785);
nand U5807 (N_5807,N_5789,N_5754);
and U5808 (N_5808,N_5730,N_5713);
and U5809 (N_5809,N_5709,N_5749);
or U5810 (N_5810,N_5773,N_5704);
xnor U5811 (N_5811,N_5798,N_5771);
xor U5812 (N_5812,N_5764,N_5748);
and U5813 (N_5813,N_5761,N_5703);
xor U5814 (N_5814,N_5775,N_5751);
and U5815 (N_5815,N_5746,N_5769);
xnor U5816 (N_5816,N_5738,N_5716);
and U5817 (N_5817,N_5725,N_5702);
or U5818 (N_5818,N_5735,N_5726);
and U5819 (N_5819,N_5706,N_5724);
or U5820 (N_5820,N_5772,N_5753);
nor U5821 (N_5821,N_5786,N_5734);
xor U5822 (N_5822,N_5745,N_5711);
nor U5823 (N_5823,N_5795,N_5757);
nor U5824 (N_5824,N_5794,N_5715);
and U5825 (N_5825,N_5721,N_5787);
or U5826 (N_5826,N_5727,N_5737);
nand U5827 (N_5827,N_5763,N_5760);
nor U5828 (N_5828,N_5719,N_5743);
and U5829 (N_5829,N_5752,N_5774);
or U5830 (N_5830,N_5756,N_5714);
and U5831 (N_5831,N_5779,N_5759);
nand U5832 (N_5832,N_5778,N_5781);
nand U5833 (N_5833,N_5731,N_5777);
nand U5834 (N_5834,N_5741,N_5717);
nor U5835 (N_5835,N_5770,N_5733);
or U5836 (N_5836,N_5790,N_5780);
xor U5837 (N_5837,N_5792,N_5791);
xor U5838 (N_5838,N_5765,N_5782);
and U5839 (N_5839,N_5744,N_5767);
nand U5840 (N_5840,N_5750,N_5729);
or U5841 (N_5841,N_5788,N_5797);
nand U5842 (N_5842,N_5755,N_5723);
nor U5843 (N_5843,N_5710,N_5793);
nand U5844 (N_5844,N_5783,N_5708);
and U5845 (N_5845,N_5700,N_5701);
xor U5846 (N_5846,N_5740,N_5718);
xnor U5847 (N_5847,N_5728,N_5784);
xnor U5848 (N_5848,N_5766,N_5707);
and U5849 (N_5849,N_5762,N_5796);
nand U5850 (N_5850,N_5767,N_5701);
nor U5851 (N_5851,N_5703,N_5744);
or U5852 (N_5852,N_5721,N_5730);
and U5853 (N_5853,N_5732,N_5737);
nand U5854 (N_5854,N_5726,N_5754);
and U5855 (N_5855,N_5700,N_5751);
nor U5856 (N_5856,N_5756,N_5758);
and U5857 (N_5857,N_5764,N_5743);
nor U5858 (N_5858,N_5702,N_5798);
or U5859 (N_5859,N_5789,N_5713);
nor U5860 (N_5860,N_5758,N_5785);
or U5861 (N_5861,N_5747,N_5797);
nor U5862 (N_5862,N_5734,N_5744);
nand U5863 (N_5863,N_5749,N_5743);
or U5864 (N_5864,N_5774,N_5703);
nor U5865 (N_5865,N_5797,N_5770);
nand U5866 (N_5866,N_5755,N_5711);
and U5867 (N_5867,N_5733,N_5716);
or U5868 (N_5868,N_5747,N_5702);
nor U5869 (N_5869,N_5748,N_5781);
and U5870 (N_5870,N_5797,N_5751);
or U5871 (N_5871,N_5725,N_5756);
nand U5872 (N_5872,N_5794,N_5711);
xor U5873 (N_5873,N_5710,N_5717);
xor U5874 (N_5874,N_5785,N_5746);
nand U5875 (N_5875,N_5747,N_5779);
nor U5876 (N_5876,N_5739,N_5709);
xor U5877 (N_5877,N_5742,N_5793);
nand U5878 (N_5878,N_5794,N_5787);
and U5879 (N_5879,N_5785,N_5755);
xnor U5880 (N_5880,N_5786,N_5724);
nor U5881 (N_5881,N_5743,N_5710);
or U5882 (N_5882,N_5708,N_5713);
nand U5883 (N_5883,N_5744,N_5755);
and U5884 (N_5884,N_5794,N_5784);
xor U5885 (N_5885,N_5766,N_5748);
nand U5886 (N_5886,N_5777,N_5798);
nor U5887 (N_5887,N_5723,N_5780);
nor U5888 (N_5888,N_5774,N_5791);
nand U5889 (N_5889,N_5715,N_5763);
or U5890 (N_5890,N_5772,N_5737);
nor U5891 (N_5891,N_5787,N_5763);
xor U5892 (N_5892,N_5718,N_5782);
or U5893 (N_5893,N_5757,N_5756);
and U5894 (N_5894,N_5784,N_5715);
nand U5895 (N_5895,N_5777,N_5700);
nor U5896 (N_5896,N_5742,N_5708);
nand U5897 (N_5897,N_5773,N_5729);
xnor U5898 (N_5898,N_5733,N_5741);
nor U5899 (N_5899,N_5782,N_5797);
or U5900 (N_5900,N_5831,N_5848);
or U5901 (N_5901,N_5875,N_5858);
nand U5902 (N_5902,N_5802,N_5873);
xor U5903 (N_5903,N_5828,N_5888);
xnor U5904 (N_5904,N_5850,N_5845);
or U5905 (N_5905,N_5827,N_5822);
nand U5906 (N_5906,N_5832,N_5880);
or U5907 (N_5907,N_5879,N_5814);
xor U5908 (N_5908,N_5899,N_5895);
nand U5909 (N_5909,N_5892,N_5813);
xor U5910 (N_5910,N_5864,N_5874);
and U5911 (N_5911,N_5840,N_5868);
nand U5912 (N_5912,N_5869,N_5824);
and U5913 (N_5913,N_5830,N_5857);
or U5914 (N_5914,N_5801,N_5825);
nor U5915 (N_5915,N_5893,N_5837);
xor U5916 (N_5916,N_5889,N_5843);
or U5917 (N_5917,N_5890,N_5841);
xor U5918 (N_5918,N_5867,N_5815);
nand U5919 (N_5919,N_5876,N_5829);
nor U5920 (N_5920,N_5846,N_5878);
xor U5921 (N_5921,N_5821,N_5887);
and U5922 (N_5922,N_5859,N_5810);
xnor U5923 (N_5923,N_5870,N_5807);
and U5924 (N_5924,N_5839,N_5820);
or U5925 (N_5925,N_5856,N_5866);
xnor U5926 (N_5926,N_5861,N_5849);
nand U5927 (N_5927,N_5851,N_5803);
nor U5928 (N_5928,N_5852,N_5886);
nor U5929 (N_5929,N_5808,N_5800);
and U5930 (N_5930,N_5883,N_5871);
and U5931 (N_5931,N_5834,N_5855);
or U5932 (N_5932,N_5863,N_5812);
and U5933 (N_5933,N_5836,N_5898);
and U5934 (N_5934,N_5894,N_5842);
and U5935 (N_5935,N_5844,N_5865);
or U5936 (N_5936,N_5860,N_5826);
nand U5937 (N_5937,N_5823,N_5897);
and U5938 (N_5938,N_5833,N_5877);
and U5939 (N_5939,N_5818,N_5882);
and U5940 (N_5940,N_5804,N_5805);
nor U5941 (N_5941,N_5853,N_5817);
and U5942 (N_5942,N_5838,N_5806);
xor U5943 (N_5943,N_5896,N_5884);
or U5944 (N_5944,N_5872,N_5854);
and U5945 (N_5945,N_5891,N_5862);
or U5946 (N_5946,N_5885,N_5847);
or U5947 (N_5947,N_5881,N_5835);
and U5948 (N_5948,N_5811,N_5816);
nor U5949 (N_5949,N_5819,N_5809);
or U5950 (N_5950,N_5815,N_5840);
nand U5951 (N_5951,N_5824,N_5831);
xor U5952 (N_5952,N_5828,N_5808);
or U5953 (N_5953,N_5800,N_5833);
xor U5954 (N_5954,N_5825,N_5894);
nand U5955 (N_5955,N_5888,N_5840);
nor U5956 (N_5956,N_5802,N_5864);
nand U5957 (N_5957,N_5830,N_5853);
or U5958 (N_5958,N_5885,N_5833);
or U5959 (N_5959,N_5871,N_5837);
or U5960 (N_5960,N_5839,N_5805);
nor U5961 (N_5961,N_5865,N_5833);
nor U5962 (N_5962,N_5875,N_5856);
or U5963 (N_5963,N_5812,N_5878);
xor U5964 (N_5964,N_5859,N_5840);
or U5965 (N_5965,N_5851,N_5854);
or U5966 (N_5966,N_5895,N_5827);
xor U5967 (N_5967,N_5821,N_5812);
xnor U5968 (N_5968,N_5863,N_5825);
nor U5969 (N_5969,N_5839,N_5812);
nor U5970 (N_5970,N_5847,N_5818);
or U5971 (N_5971,N_5862,N_5831);
or U5972 (N_5972,N_5827,N_5853);
nor U5973 (N_5973,N_5831,N_5894);
or U5974 (N_5974,N_5837,N_5824);
or U5975 (N_5975,N_5875,N_5848);
xnor U5976 (N_5976,N_5829,N_5806);
nor U5977 (N_5977,N_5838,N_5843);
nand U5978 (N_5978,N_5868,N_5876);
or U5979 (N_5979,N_5894,N_5851);
and U5980 (N_5980,N_5869,N_5856);
nor U5981 (N_5981,N_5893,N_5872);
xor U5982 (N_5982,N_5810,N_5882);
nand U5983 (N_5983,N_5814,N_5876);
and U5984 (N_5984,N_5852,N_5882);
and U5985 (N_5985,N_5838,N_5829);
xnor U5986 (N_5986,N_5873,N_5829);
or U5987 (N_5987,N_5872,N_5860);
or U5988 (N_5988,N_5899,N_5885);
nor U5989 (N_5989,N_5884,N_5881);
nor U5990 (N_5990,N_5890,N_5814);
nor U5991 (N_5991,N_5872,N_5824);
and U5992 (N_5992,N_5896,N_5860);
xnor U5993 (N_5993,N_5830,N_5807);
nand U5994 (N_5994,N_5874,N_5859);
xor U5995 (N_5995,N_5865,N_5809);
nor U5996 (N_5996,N_5857,N_5854);
nand U5997 (N_5997,N_5829,N_5887);
and U5998 (N_5998,N_5873,N_5816);
nor U5999 (N_5999,N_5876,N_5817);
and U6000 (N_6000,N_5900,N_5926);
nand U6001 (N_6001,N_5903,N_5902);
xor U6002 (N_6002,N_5995,N_5922);
nand U6003 (N_6003,N_5996,N_5961);
or U6004 (N_6004,N_5999,N_5913);
or U6005 (N_6005,N_5947,N_5958);
xnor U6006 (N_6006,N_5935,N_5951);
and U6007 (N_6007,N_5967,N_5960);
nand U6008 (N_6008,N_5953,N_5925);
nand U6009 (N_6009,N_5950,N_5915);
and U6010 (N_6010,N_5909,N_5956);
nor U6011 (N_6011,N_5994,N_5987);
and U6012 (N_6012,N_5973,N_5949);
xnor U6013 (N_6013,N_5986,N_5948);
nand U6014 (N_6014,N_5917,N_5969);
nor U6015 (N_6015,N_5941,N_5938);
xnor U6016 (N_6016,N_5939,N_5919);
xor U6017 (N_6017,N_5934,N_5907);
and U6018 (N_6018,N_5985,N_5988);
and U6019 (N_6019,N_5920,N_5929);
nand U6020 (N_6020,N_5980,N_5933);
xnor U6021 (N_6021,N_5944,N_5916);
and U6022 (N_6022,N_5970,N_5981);
xnor U6023 (N_6023,N_5966,N_5905);
xor U6024 (N_6024,N_5962,N_5910);
nand U6025 (N_6025,N_5965,N_5940);
xnor U6026 (N_6026,N_5971,N_5975);
and U6027 (N_6027,N_5964,N_5991);
or U6028 (N_6028,N_5911,N_5954);
or U6029 (N_6029,N_5928,N_5943);
nand U6030 (N_6030,N_5989,N_5923);
nand U6031 (N_6031,N_5979,N_5952);
nor U6032 (N_6032,N_5997,N_5959);
nor U6033 (N_6033,N_5976,N_5972);
xor U6034 (N_6034,N_5945,N_5983);
xnor U6035 (N_6035,N_5990,N_5955);
or U6036 (N_6036,N_5957,N_5918);
nand U6037 (N_6037,N_5921,N_5984);
and U6038 (N_6038,N_5901,N_5974);
or U6039 (N_6039,N_5968,N_5993);
xor U6040 (N_6040,N_5946,N_5904);
and U6041 (N_6041,N_5908,N_5927);
and U6042 (N_6042,N_5912,N_5998);
nor U6043 (N_6043,N_5906,N_5937);
nand U6044 (N_6044,N_5931,N_5930);
or U6045 (N_6045,N_5942,N_5914);
or U6046 (N_6046,N_5932,N_5924);
and U6047 (N_6047,N_5978,N_5992);
xnor U6048 (N_6048,N_5936,N_5977);
nor U6049 (N_6049,N_5982,N_5963);
or U6050 (N_6050,N_5988,N_5921);
or U6051 (N_6051,N_5905,N_5930);
nor U6052 (N_6052,N_5912,N_5988);
nor U6053 (N_6053,N_5948,N_5908);
xor U6054 (N_6054,N_5944,N_5903);
xnor U6055 (N_6055,N_5999,N_5984);
nor U6056 (N_6056,N_5993,N_5929);
and U6057 (N_6057,N_5940,N_5923);
and U6058 (N_6058,N_5921,N_5939);
nor U6059 (N_6059,N_5981,N_5916);
xnor U6060 (N_6060,N_5977,N_5985);
nor U6061 (N_6061,N_5990,N_5961);
nor U6062 (N_6062,N_5951,N_5996);
and U6063 (N_6063,N_5971,N_5911);
or U6064 (N_6064,N_5906,N_5943);
nand U6065 (N_6065,N_5965,N_5944);
xnor U6066 (N_6066,N_5982,N_5914);
and U6067 (N_6067,N_5999,N_5952);
nand U6068 (N_6068,N_5901,N_5982);
xnor U6069 (N_6069,N_5956,N_5901);
xor U6070 (N_6070,N_5914,N_5946);
nand U6071 (N_6071,N_5974,N_5927);
and U6072 (N_6072,N_5900,N_5938);
and U6073 (N_6073,N_5990,N_5989);
and U6074 (N_6074,N_5970,N_5975);
nor U6075 (N_6075,N_5996,N_5969);
nor U6076 (N_6076,N_5910,N_5946);
nand U6077 (N_6077,N_5903,N_5999);
nor U6078 (N_6078,N_5977,N_5937);
or U6079 (N_6079,N_5915,N_5922);
xor U6080 (N_6080,N_5921,N_5983);
xnor U6081 (N_6081,N_5938,N_5919);
xor U6082 (N_6082,N_5976,N_5922);
and U6083 (N_6083,N_5927,N_5992);
or U6084 (N_6084,N_5967,N_5976);
nor U6085 (N_6085,N_5947,N_5916);
nand U6086 (N_6086,N_5977,N_5976);
nand U6087 (N_6087,N_5910,N_5980);
or U6088 (N_6088,N_5914,N_5950);
and U6089 (N_6089,N_5900,N_5954);
and U6090 (N_6090,N_5988,N_5943);
or U6091 (N_6091,N_5941,N_5964);
and U6092 (N_6092,N_5935,N_5926);
xor U6093 (N_6093,N_5954,N_5989);
nor U6094 (N_6094,N_5968,N_5984);
xor U6095 (N_6095,N_5969,N_5921);
or U6096 (N_6096,N_5994,N_5977);
and U6097 (N_6097,N_5909,N_5932);
xor U6098 (N_6098,N_5917,N_5990);
or U6099 (N_6099,N_5905,N_5976);
xor U6100 (N_6100,N_6016,N_6033);
and U6101 (N_6101,N_6044,N_6045);
nand U6102 (N_6102,N_6038,N_6075);
nand U6103 (N_6103,N_6055,N_6024);
nor U6104 (N_6104,N_6068,N_6091);
xor U6105 (N_6105,N_6047,N_6071);
nand U6106 (N_6106,N_6067,N_6073);
or U6107 (N_6107,N_6007,N_6049);
nand U6108 (N_6108,N_6036,N_6026);
nand U6109 (N_6109,N_6015,N_6054);
nor U6110 (N_6110,N_6041,N_6000);
and U6111 (N_6111,N_6089,N_6051);
nand U6112 (N_6112,N_6008,N_6052);
and U6113 (N_6113,N_6012,N_6023);
nand U6114 (N_6114,N_6031,N_6097);
or U6115 (N_6115,N_6017,N_6035);
nand U6116 (N_6116,N_6099,N_6066);
or U6117 (N_6117,N_6076,N_6062);
and U6118 (N_6118,N_6098,N_6058);
or U6119 (N_6119,N_6079,N_6021);
nand U6120 (N_6120,N_6085,N_6064);
nor U6121 (N_6121,N_6029,N_6050);
and U6122 (N_6122,N_6013,N_6092);
or U6123 (N_6123,N_6082,N_6048);
and U6124 (N_6124,N_6074,N_6004);
nand U6125 (N_6125,N_6090,N_6080);
nand U6126 (N_6126,N_6084,N_6009);
nor U6127 (N_6127,N_6069,N_6053);
or U6128 (N_6128,N_6065,N_6032);
and U6129 (N_6129,N_6006,N_6001);
or U6130 (N_6130,N_6095,N_6025);
nand U6131 (N_6131,N_6088,N_6094);
and U6132 (N_6132,N_6034,N_6056);
or U6133 (N_6133,N_6057,N_6059);
or U6134 (N_6134,N_6060,N_6040);
nand U6135 (N_6135,N_6070,N_6042);
nor U6136 (N_6136,N_6005,N_6002);
xnor U6137 (N_6137,N_6020,N_6028);
nand U6138 (N_6138,N_6018,N_6078);
nand U6139 (N_6139,N_6086,N_6077);
xor U6140 (N_6140,N_6072,N_6022);
xnor U6141 (N_6141,N_6083,N_6011);
xor U6142 (N_6142,N_6087,N_6093);
and U6143 (N_6143,N_6003,N_6046);
nand U6144 (N_6144,N_6010,N_6037);
and U6145 (N_6145,N_6063,N_6027);
or U6146 (N_6146,N_6043,N_6061);
nor U6147 (N_6147,N_6081,N_6014);
xnor U6148 (N_6148,N_6096,N_6019);
xor U6149 (N_6149,N_6030,N_6039);
or U6150 (N_6150,N_6088,N_6019);
xnor U6151 (N_6151,N_6046,N_6005);
nor U6152 (N_6152,N_6014,N_6048);
nor U6153 (N_6153,N_6065,N_6029);
and U6154 (N_6154,N_6095,N_6015);
nand U6155 (N_6155,N_6080,N_6038);
or U6156 (N_6156,N_6043,N_6042);
xor U6157 (N_6157,N_6045,N_6017);
and U6158 (N_6158,N_6004,N_6036);
or U6159 (N_6159,N_6012,N_6094);
and U6160 (N_6160,N_6088,N_6079);
or U6161 (N_6161,N_6041,N_6081);
xor U6162 (N_6162,N_6027,N_6032);
nand U6163 (N_6163,N_6064,N_6097);
or U6164 (N_6164,N_6035,N_6051);
nor U6165 (N_6165,N_6027,N_6081);
nand U6166 (N_6166,N_6058,N_6020);
and U6167 (N_6167,N_6012,N_6086);
nor U6168 (N_6168,N_6086,N_6071);
nand U6169 (N_6169,N_6036,N_6025);
nand U6170 (N_6170,N_6014,N_6057);
nand U6171 (N_6171,N_6040,N_6021);
or U6172 (N_6172,N_6042,N_6039);
nor U6173 (N_6173,N_6018,N_6046);
and U6174 (N_6174,N_6047,N_6020);
and U6175 (N_6175,N_6084,N_6089);
nor U6176 (N_6176,N_6067,N_6087);
xor U6177 (N_6177,N_6038,N_6018);
xnor U6178 (N_6178,N_6094,N_6013);
nor U6179 (N_6179,N_6091,N_6007);
and U6180 (N_6180,N_6032,N_6070);
xor U6181 (N_6181,N_6090,N_6011);
xnor U6182 (N_6182,N_6044,N_6091);
or U6183 (N_6183,N_6039,N_6090);
nor U6184 (N_6184,N_6054,N_6009);
or U6185 (N_6185,N_6050,N_6073);
or U6186 (N_6186,N_6005,N_6040);
nand U6187 (N_6187,N_6017,N_6014);
nand U6188 (N_6188,N_6013,N_6030);
nand U6189 (N_6189,N_6018,N_6081);
or U6190 (N_6190,N_6069,N_6015);
and U6191 (N_6191,N_6044,N_6039);
and U6192 (N_6192,N_6098,N_6054);
xnor U6193 (N_6193,N_6045,N_6001);
or U6194 (N_6194,N_6042,N_6048);
xor U6195 (N_6195,N_6004,N_6083);
nor U6196 (N_6196,N_6028,N_6087);
nand U6197 (N_6197,N_6049,N_6032);
nor U6198 (N_6198,N_6061,N_6087);
or U6199 (N_6199,N_6066,N_6076);
nor U6200 (N_6200,N_6114,N_6171);
xnor U6201 (N_6201,N_6153,N_6122);
xor U6202 (N_6202,N_6143,N_6186);
nor U6203 (N_6203,N_6168,N_6115);
nand U6204 (N_6204,N_6136,N_6189);
xnor U6205 (N_6205,N_6184,N_6105);
and U6206 (N_6206,N_6135,N_6141);
xnor U6207 (N_6207,N_6190,N_6161);
nor U6208 (N_6208,N_6158,N_6144);
nor U6209 (N_6209,N_6197,N_6103);
nand U6210 (N_6210,N_6151,N_6146);
nand U6211 (N_6211,N_6125,N_6152);
xnor U6212 (N_6212,N_6106,N_6121);
and U6213 (N_6213,N_6162,N_6169);
nor U6214 (N_6214,N_6116,N_6155);
and U6215 (N_6215,N_6188,N_6107);
nor U6216 (N_6216,N_6101,N_6118);
and U6217 (N_6217,N_6117,N_6150);
and U6218 (N_6218,N_6134,N_6163);
nor U6219 (N_6219,N_6183,N_6164);
nor U6220 (N_6220,N_6172,N_6175);
nor U6221 (N_6221,N_6109,N_6112);
nor U6222 (N_6222,N_6167,N_6142);
and U6223 (N_6223,N_6126,N_6173);
and U6224 (N_6224,N_6154,N_6157);
and U6225 (N_6225,N_6166,N_6176);
nand U6226 (N_6226,N_6124,N_6181);
or U6227 (N_6227,N_6127,N_6123);
nand U6228 (N_6228,N_6196,N_6147);
xnor U6229 (N_6229,N_6133,N_6174);
or U6230 (N_6230,N_6130,N_6120);
nand U6231 (N_6231,N_6195,N_6113);
and U6232 (N_6232,N_6179,N_6139);
nor U6233 (N_6233,N_6119,N_6148);
nand U6234 (N_6234,N_6128,N_6156);
xor U6235 (N_6235,N_6160,N_6193);
or U6236 (N_6236,N_6100,N_6132);
and U6237 (N_6237,N_6129,N_6110);
and U6238 (N_6238,N_6170,N_6140);
and U6239 (N_6239,N_6180,N_6104);
or U6240 (N_6240,N_6199,N_6138);
or U6241 (N_6241,N_6165,N_6198);
xor U6242 (N_6242,N_6108,N_6177);
or U6243 (N_6243,N_6191,N_6159);
nor U6244 (N_6244,N_6194,N_6131);
xor U6245 (N_6245,N_6182,N_6145);
nor U6246 (N_6246,N_6137,N_6185);
nor U6247 (N_6247,N_6187,N_6111);
nand U6248 (N_6248,N_6102,N_6192);
xor U6249 (N_6249,N_6178,N_6149);
xnor U6250 (N_6250,N_6146,N_6152);
xnor U6251 (N_6251,N_6165,N_6145);
xnor U6252 (N_6252,N_6155,N_6114);
xnor U6253 (N_6253,N_6166,N_6190);
nor U6254 (N_6254,N_6191,N_6124);
and U6255 (N_6255,N_6154,N_6179);
or U6256 (N_6256,N_6107,N_6145);
or U6257 (N_6257,N_6117,N_6142);
or U6258 (N_6258,N_6163,N_6148);
nand U6259 (N_6259,N_6187,N_6168);
nor U6260 (N_6260,N_6152,N_6102);
and U6261 (N_6261,N_6195,N_6123);
xor U6262 (N_6262,N_6141,N_6145);
xor U6263 (N_6263,N_6156,N_6122);
nand U6264 (N_6264,N_6128,N_6155);
nor U6265 (N_6265,N_6197,N_6176);
nor U6266 (N_6266,N_6110,N_6186);
xnor U6267 (N_6267,N_6171,N_6119);
nor U6268 (N_6268,N_6171,N_6166);
nand U6269 (N_6269,N_6143,N_6178);
and U6270 (N_6270,N_6181,N_6126);
or U6271 (N_6271,N_6155,N_6196);
xnor U6272 (N_6272,N_6197,N_6141);
nand U6273 (N_6273,N_6175,N_6112);
or U6274 (N_6274,N_6136,N_6160);
nor U6275 (N_6275,N_6150,N_6163);
and U6276 (N_6276,N_6110,N_6182);
nand U6277 (N_6277,N_6143,N_6145);
xor U6278 (N_6278,N_6181,N_6105);
or U6279 (N_6279,N_6147,N_6125);
or U6280 (N_6280,N_6162,N_6103);
or U6281 (N_6281,N_6150,N_6128);
nand U6282 (N_6282,N_6102,N_6126);
nor U6283 (N_6283,N_6109,N_6107);
or U6284 (N_6284,N_6133,N_6115);
nand U6285 (N_6285,N_6198,N_6159);
xor U6286 (N_6286,N_6172,N_6193);
xor U6287 (N_6287,N_6116,N_6174);
xor U6288 (N_6288,N_6136,N_6100);
or U6289 (N_6289,N_6155,N_6192);
nor U6290 (N_6290,N_6133,N_6125);
nand U6291 (N_6291,N_6172,N_6192);
nand U6292 (N_6292,N_6196,N_6167);
or U6293 (N_6293,N_6130,N_6163);
or U6294 (N_6294,N_6127,N_6154);
nand U6295 (N_6295,N_6173,N_6172);
nand U6296 (N_6296,N_6154,N_6122);
and U6297 (N_6297,N_6107,N_6192);
nand U6298 (N_6298,N_6102,N_6149);
nor U6299 (N_6299,N_6186,N_6157);
or U6300 (N_6300,N_6268,N_6295);
or U6301 (N_6301,N_6208,N_6249);
nand U6302 (N_6302,N_6272,N_6259);
nand U6303 (N_6303,N_6271,N_6266);
nor U6304 (N_6304,N_6297,N_6222);
or U6305 (N_6305,N_6231,N_6292);
nor U6306 (N_6306,N_6269,N_6237);
and U6307 (N_6307,N_6273,N_6244);
xor U6308 (N_6308,N_6218,N_6252);
xnor U6309 (N_6309,N_6247,N_6219);
and U6310 (N_6310,N_6270,N_6260);
or U6311 (N_6311,N_6267,N_6261);
nor U6312 (N_6312,N_6285,N_6248);
or U6313 (N_6313,N_6225,N_6211);
and U6314 (N_6314,N_6291,N_6290);
and U6315 (N_6315,N_6284,N_6293);
nand U6316 (N_6316,N_6234,N_6255);
or U6317 (N_6317,N_6280,N_6205);
nor U6318 (N_6318,N_6277,N_6283);
nor U6319 (N_6319,N_6235,N_6243);
or U6320 (N_6320,N_6262,N_6229);
nor U6321 (N_6321,N_6216,N_6246);
nand U6322 (N_6322,N_6202,N_6276);
nand U6323 (N_6323,N_6228,N_6251);
and U6324 (N_6324,N_6224,N_6298);
nor U6325 (N_6325,N_6206,N_6286);
xnor U6326 (N_6326,N_6258,N_6288);
and U6327 (N_6327,N_6294,N_6264);
nor U6328 (N_6328,N_6299,N_6213);
nand U6329 (N_6329,N_6217,N_6236);
nor U6330 (N_6330,N_6253,N_6281);
nand U6331 (N_6331,N_6233,N_6209);
xor U6332 (N_6332,N_6226,N_6275);
nand U6333 (N_6333,N_6203,N_6296);
xor U6334 (N_6334,N_6210,N_6204);
and U6335 (N_6335,N_6282,N_6212);
or U6336 (N_6336,N_6221,N_6265);
xnor U6337 (N_6337,N_6245,N_6242);
xnor U6338 (N_6338,N_6207,N_6279);
nand U6339 (N_6339,N_6215,N_6289);
nand U6340 (N_6340,N_6274,N_6241);
or U6341 (N_6341,N_6257,N_6230);
nor U6342 (N_6342,N_6254,N_6238);
nand U6343 (N_6343,N_6240,N_6287);
and U6344 (N_6344,N_6263,N_6223);
nand U6345 (N_6345,N_6278,N_6214);
nor U6346 (N_6346,N_6201,N_6250);
and U6347 (N_6347,N_6239,N_6256);
xor U6348 (N_6348,N_6232,N_6200);
nor U6349 (N_6349,N_6220,N_6227);
nand U6350 (N_6350,N_6220,N_6254);
nand U6351 (N_6351,N_6202,N_6256);
xnor U6352 (N_6352,N_6206,N_6287);
xor U6353 (N_6353,N_6263,N_6295);
and U6354 (N_6354,N_6236,N_6299);
and U6355 (N_6355,N_6273,N_6291);
or U6356 (N_6356,N_6276,N_6269);
or U6357 (N_6357,N_6264,N_6203);
nand U6358 (N_6358,N_6266,N_6257);
nand U6359 (N_6359,N_6264,N_6265);
or U6360 (N_6360,N_6297,N_6209);
nand U6361 (N_6361,N_6258,N_6263);
xor U6362 (N_6362,N_6273,N_6290);
and U6363 (N_6363,N_6269,N_6275);
and U6364 (N_6364,N_6266,N_6239);
nor U6365 (N_6365,N_6277,N_6267);
nor U6366 (N_6366,N_6218,N_6220);
and U6367 (N_6367,N_6203,N_6297);
and U6368 (N_6368,N_6205,N_6287);
nand U6369 (N_6369,N_6274,N_6211);
nor U6370 (N_6370,N_6236,N_6253);
or U6371 (N_6371,N_6257,N_6273);
or U6372 (N_6372,N_6216,N_6241);
nor U6373 (N_6373,N_6206,N_6290);
or U6374 (N_6374,N_6263,N_6237);
or U6375 (N_6375,N_6213,N_6260);
nand U6376 (N_6376,N_6210,N_6243);
or U6377 (N_6377,N_6285,N_6257);
nand U6378 (N_6378,N_6235,N_6222);
or U6379 (N_6379,N_6270,N_6261);
nor U6380 (N_6380,N_6220,N_6230);
nor U6381 (N_6381,N_6259,N_6244);
and U6382 (N_6382,N_6200,N_6242);
xor U6383 (N_6383,N_6259,N_6299);
nand U6384 (N_6384,N_6263,N_6260);
nor U6385 (N_6385,N_6237,N_6287);
nor U6386 (N_6386,N_6298,N_6285);
xnor U6387 (N_6387,N_6221,N_6271);
xor U6388 (N_6388,N_6291,N_6267);
nand U6389 (N_6389,N_6295,N_6279);
and U6390 (N_6390,N_6241,N_6256);
and U6391 (N_6391,N_6247,N_6218);
nand U6392 (N_6392,N_6246,N_6288);
and U6393 (N_6393,N_6260,N_6251);
and U6394 (N_6394,N_6245,N_6213);
nand U6395 (N_6395,N_6287,N_6278);
or U6396 (N_6396,N_6204,N_6227);
and U6397 (N_6397,N_6281,N_6202);
nand U6398 (N_6398,N_6225,N_6240);
nor U6399 (N_6399,N_6220,N_6280);
nand U6400 (N_6400,N_6395,N_6359);
and U6401 (N_6401,N_6322,N_6316);
nand U6402 (N_6402,N_6353,N_6344);
nor U6403 (N_6403,N_6342,N_6345);
nand U6404 (N_6404,N_6373,N_6365);
or U6405 (N_6405,N_6339,N_6312);
or U6406 (N_6406,N_6309,N_6326);
xnor U6407 (N_6407,N_6333,N_6381);
nand U6408 (N_6408,N_6380,N_6323);
or U6409 (N_6409,N_6363,N_6383);
nor U6410 (N_6410,N_6388,N_6329);
nand U6411 (N_6411,N_6313,N_6389);
nor U6412 (N_6412,N_6357,N_6341);
or U6413 (N_6413,N_6325,N_6347);
nor U6414 (N_6414,N_6327,N_6304);
xnor U6415 (N_6415,N_6315,N_6314);
nand U6416 (N_6416,N_6350,N_6386);
xnor U6417 (N_6417,N_6354,N_6305);
xnor U6418 (N_6418,N_6321,N_6384);
nor U6419 (N_6419,N_6375,N_6340);
xor U6420 (N_6420,N_6330,N_6378);
nor U6421 (N_6421,N_6392,N_6355);
xnor U6422 (N_6422,N_6300,N_6393);
xnor U6423 (N_6423,N_6331,N_6379);
and U6424 (N_6424,N_6361,N_6351);
and U6425 (N_6425,N_6376,N_6377);
and U6426 (N_6426,N_6362,N_6372);
and U6427 (N_6427,N_6338,N_6387);
nor U6428 (N_6428,N_6328,N_6306);
or U6429 (N_6429,N_6334,N_6346);
xor U6430 (N_6430,N_6398,N_6301);
or U6431 (N_6431,N_6385,N_6343);
xnor U6432 (N_6432,N_6307,N_6332);
nand U6433 (N_6433,N_6358,N_6317);
nor U6434 (N_6434,N_6335,N_6324);
nor U6435 (N_6435,N_6367,N_6311);
and U6436 (N_6436,N_6369,N_6349);
and U6437 (N_6437,N_6390,N_6366);
xnor U6438 (N_6438,N_6337,N_6356);
nor U6439 (N_6439,N_6374,N_6394);
xnor U6440 (N_6440,N_6320,N_6302);
nor U6441 (N_6441,N_6370,N_6318);
nand U6442 (N_6442,N_6391,N_6310);
and U6443 (N_6443,N_6368,N_6364);
nor U6444 (N_6444,N_6352,N_6303);
nor U6445 (N_6445,N_6336,N_6319);
nor U6446 (N_6446,N_6397,N_6348);
or U6447 (N_6447,N_6360,N_6399);
and U6448 (N_6448,N_6308,N_6382);
xor U6449 (N_6449,N_6396,N_6371);
and U6450 (N_6450,N_6306,N_6373);
nor U6451 (N_6451,N_6392,N_6326);
nor U6452 (N_6452,N_6336,N_6337);
xnor U6453 (N_6453,N_6383,N_6368);
or U6454 (N_6454,N_6390,N_6339);
nor U6455 (N_6455,N_6332,N_6334);
or U6456 (N_6456,N_6376,N_6308);
xnor U6457 (N_6457,N_6355,N_6364);
xnor U6458 (N_6458,N_6384,N_6324);
and U6459 (N_6459,N_6379,N_6373);
and U6460 (N_6460,N_6301,N_6324);
or U6461 (N_6461,N_6338,N_6321);
xnor U6462 (N_6462,N_6392,N_6351);
and U6463 (N_6463,N_6362,N_6387);
and U6464 (N_6464,N_6318,N_6324);
and U6465 (N_6465,N_6366,N_6325);
or U6466 (N_6466,N_6393,N_6309);
nor U6467 (N_6467,N_6352,N_6343);
xor U6468 (N_6468,N_6304,N_6345);
and U6469 (N_6469,N_6378,N_6345);
and U6470 (N_6470,N_6350,N_6356);
xnor U6471 (N_6471,N_6324,N_6377);
and U6472 (N_6472,N_6373,N_6353);
and U6473 (N_6473,N_6392,N_6312);
nand U6474 (N_6474,N_6387,N_6342);
and U6475 (N_6475,N_6321,N_6388);
and U6476 (N_6476,N_6335,N_6322);
and U6477 (N_6477,N_6378,N_6367);
and U6478 (N_6478,N_6319,N_6345);
nor U6479 (N_6479,N_6372,N_6331);
nand U6480 (N_6480,N_6356,N_6392);
nand U6481 (N_6481,N_6373,N_6396);
nand U6482 (N_6482,N_6365,N_6387);
xor U6483 (N_6483,N_6356,N_6369);
nand U6484 (N_6484,N_6340,N_6384);
or U6485 (N_6485,N_6364,N_6304);
xnor U6486 (N_6486,N_6340,N_6317);
or U6487 (N_6487,N_6345,N_6399);
and U6488 (N_6488,N_6397,N_6319);
xor U6489 (N_6489,N_6323,N_6312);
and U6490 (N_6490,N_6393,N_6369);
xor U6491 (N_6491,N_6325,N_6380);
nand U6492 (N_6492,N_6312,N_6353);
and U6493 (N_6493,N_6348,N_6307);
or U6494 (N_6494,N_6358,N_6356);
nor U6495 (N_6495,N_6384,N_6361);
and U6496 (N_6496,N_6358,N_6345);
nor U6497 (N_6497,N_6310,N_6351);
or U6498 (N_6498,N_6349,N_6372);
and U6499 (N_6499,N_6303,N_6397);
and U6500 (N_6500,N_6483,N_6427);
nand U6501 (N_6501,N_6468,N_6443);
and U6502 (N_6502,N_6472,N_6431);
nor U6503 (N_6503,N_6417,N_6451);
nand U6504 (N_6504,N_6485,N_6475);
nor U6505 (N_6505,N_6450,N_6442);
or U6506 (N_6506,N_6419,N_6411);
or U6507 (N_6507,N_6453,N_6459);
xnor U6508 (N_6508,N_6455,N_6444);
nor U6509 (N_6509,N_6400,N_6476);
or U6510 (N_6510,N_6441,N_6434);
xor U6511 (N_6511,N_6413,N_6402);
and U6512 (N_6512,N_6469,N_6478);
or U6513 (N_6513,N_6420,N_6407);
or U6514 (N_6514,N_6426,N_6477);
nand U6515 (N_6515,N_6423,N_6414);
or U6516 (N_6516,N_6461,N_6466);
nand U6517 (N_6517,N_6465,N_6457);
or U6518 (N_6518,N_6498,N_6435);
and U6519 (N_6519,N_6496,N_6471);
and U6520 (N_6520,N_6489,N_6460);
or U6521 (N_6521,N_6482,N_6412);
xnor U6522 (N_6522,N_6458,N_6432);
nor U6523 (N_6523,N_6474,N_6490);
and U6524 (N_6524,N_6452,N_6494);
nand U6525 (N_6525,N_6481,N_6408);
nand U6526 (N_6526,N_6488,N_6422);
nor U6527 (N_6527,N_6447,N_6486);
or U6528 (N_6528,N_6415,N_6404);
nor U6529 (N_6529,N_6436,N_6418);
nand U6530 (N_6530,N_6409,N_6425);
xnor U6531 (N_6531,N_6403,N_6439);
or U6532 (N_6532,N_6416,N_6421);
or U6533 (N_6533,N_6473,N_6480);
and U6534 (N_6534,N_6467,N_6424);
xnor U6535 (N_6535,N_6448,N_6492);
and U6536 (N_6536,N_6493,N_6438);
nor U6537 (N_6537,N_6464,N_6430);
nand U6538 (N_6538,N_6462,N_6437);
nand U6539 (N_6539,N_6433,N_6449);
and U6540 (N_6540,N_6479,N_6406);
or U6541 (N_6541,N_6495,N_6454);
xnor U6542 (N_6542,N_6491,N_6445);
xor U6543 (N_6543,N_6470,N_6405);
xor U6544 (N_6544,N_6429,N_6446);
xor U6545 (N_6545,N_6487,N_6484);
nand U6546 (N_6546,N_6463,N_6428);
or U6547 (N_6547,N_6440,N_6497);
or U6548 (N_6548,N_6499,N_6401);
or U6549 (N_6549,N_6410,N_6456);
or U6550 (N_6550,N_6473,N_6460);
nor U6551 (N_6551,N_6423,N_6439);
and U6552 (N_6552,N_6461,N_6426);
nand U6553 (N_6553,N_6439,N_6402);
or U6554 (N_6554,N_6415,N_6469);
and U6555 (N_6555,N_6486,N_6491);
xor U6556 (N_6556,N_6463,N_6457);
and U6557 (N_6557,N_6415,N_6441);
and U6558 (N_6558,N_6475,N_6461);
nand U6559 (N_6559,N_6463,N_6475);
nand U6560 (N_6560,N_6414,N_6431);
and U6561 (N_6561,N_6439,N_6409);
nand U6562 (N_6562,N_6419,N_6413);
and U6563 (N_6563,N_6415,N_6488);
and U6564 (N_6564,N_6491,N_6449);
nor U6565 (N_6565,N_6403,N_6474);
nand U6566 (N_6566,N_6498,N_6491);
nor U6567 (N_6567,N_6406,N_6446);
or U6568 (N_6568,N_6451,N_6464);
or U6569 (N_6569,N_6450,N_6417);
or U6570 (N_6570,N_6427,N_6476);
or U6571 (N_6571,N_6493,N_6419);
xnor U6572 (N_6572,N_6412,N_6455);
and U6573 (N_6573,N_6434,N_6408);
or U6574 (N_6574,N_6453,N_6449);
nor U6575 (N_6575,N_6493,N_6468);
or U6576 (N_6576,N_6445,N_6404);
and U6577 (N_6577,N_6418,N_6489);
or U6578 (N_6578,N_6465,N_6489);
nor U6579 (N_6579,N_6490,N_6448);
and U6580 (N_6580,N_6401,N_6425);
xnor U6581 (N_6581,N_6473,N_6469);
and U6582 (N_6582,N_6463,N_6480);
and U6583 (N_6583,N_6402,N_6446);
or U6584 (N_6584,N_6476,N_6492);
nand U6585 (N_6585,N_6472,N_6499);
xnor U6586 (N_6586,N_6481,N_6476);
nor U6587 (N_6587,N_6404,N_6441);
xor U6588 (N_6588,N_6427,N_6418);
and U6589 (N_6589,N_6431,N_6428);
nand U6590 (N_6590,N_6440,N_6445);
nand U6591 (N_6591,N_6495,N_6428);
or U6592 (N_6592,N_6459,N_6495);
nand U6593 (N_6593,N_6438,N_6415);
and U6594 (N_6594,N_6447,N_6480);
and U6595 (N_6595,N_6427,N_6478);
nand U6596 (N_6596,N_6483,N_6452);
nand U6597 (N_6597,N_6461,N_6436);
or U6598 (N_6598,N_6447,N_6498);
or U6599 (N_6599,N_6483,N_6462);
nor U6600 (N_6600,N_6507,N_6594);
and U6601 (N_6601,N_6533,N_6527);
nand U6602 (N_6602,N_6575,N_6510);
or U6603 (N_6603,N_6523,N_6553);
xor U6604 (N_6604,N_6572,N_6590);
and U6605 (N_6605,N_6557,N_6531);
nor U6606 (N_6606,N_6559,N_6556);
nand U6607 (N_6607,N_6503,N_6501);
nor U6608 (N_6608,N_6506,N_6587);
or U6609 (N_6609,N_6565,N_6597);
xor U6610 (N_6610,N_6580,N_6534);
or U6611 (N_6611,N_6524,N_6591);
or U6612 (N_6612,N_6543,N_6549);
or U6613 (N_6613,N_6509,N_6569);
nor U6614 (N_6614,N_6576,N_6568);
nor U6615 (N_6615,N_6536,N_6530);
nor U6616 (N_6616,N_6528,N_6564);
nor U6617 (N_6617,N_6513,N_6567);
nor U6618 (N_6618,N_6552,N_6500);
xnor U6619 (N_6619,N_6525,N_6560);
nor U6620 (N_6620,N_6555,N_6599);
xnor U6621 (N_6621,N_6511,N_6541);
xnor U6622 (N_6622,N_6535,N_6554);
xnor U6623 (N_6623,N_6532,N_6544);
xnor U6624 (N_6624,N_6573,N_6545);
nand U6625 (N_6625,N_6584,N_6579);
nand U6626 (N_6626,N_6521,N_6504);
and U6627 (N_6627,N_6598,N_6515);
and U6628 (N_6628,N_6517,N_6592);
and U6629 (N_6629,N_6593,N_6583);
and U6630 (N_6630,N_6566,N_6546);
and U6631 (N_6631,N_6529,N_6581);
or U6632 (N_6632,N_6516,N_6538);
nor U6633 (N_6633,N_6595,N_6558);
nor U6634 (N_6634,N_6578,N_6586);
nor U6635 (N_6635,N_6571,N_6542);
nand U6636 (N_6636,N_6502,N_6520);
nand U6637 (N_6637,N_6518,N_6512);
or U6638 (N_6638,N_6561,N_6596);
or U6639 (N_6639,N_6519,N_6562);
and U6640 (N_6640,N_6508,N_6589);
nor U6641 (N_6641,N_6551,N_6537);
xor U6642 (N_6642,N_6563,N_6547);
and U6643 (N_6643,N_6539,N_6522);
nor U6644 (N_6644,N_6582,N_6588);
and U6645 (N_6645,N_6577,N_6570);
and U6646 (N_6646,N_6574,N_6548);
xor U6647 (N_6647,N_6514,N_6540);
nand U6648 (N_6648,N_6550,N_6585);
nor U6649 (N_6649,N_6526,N_6505);
nand U6650 (N_6650,N_6511,N_6512);
xor U6651 (N_6651,N_6536,N_6557);
xnor U6652 (N_6652,N_6531,N_6556);
xnor U6653 (N_6653,N_6575,N_6522);
nand U6654 (N_6654,N_6532,N_6566);
and U6655 (N_6655,N_6545,N_6541);
xnor U6656 (N_6656,N_6566,N_6514);
nor U6657 (N_6657,N_6540,N_6590);
and U6658 (N_6658,N_6531,N_6585);
nand U6659 (N_6659,N_6529,N_6509);
nand U6660 (N_6660,N_6571,N_6504);
xnor U6661 (N_6661,N_6510,N_6573);
nand U6662 (N_6662,N_6574,N_6500);
or U6663 (N_6663,N_6525,N_6503);
and U6664 (N_6664,N_6523,N_6529);
nand U6665 (N_6665,N_6516,N_6519);
and U6666 (N_6666,N_6534,N_6587);
and U6667 (N_6667,N_6570,N_6583);
xor U6668 (N_6668,N_6524,N_6543);
nand U6669 (N_6669,N_6545,N_6596);
nand U6670 (N_6670,N_6578,N_6510);
and U6671 (N_6671,N_6535,N_6517);
nor U6672 (N_6672,N_6595,N_6507);
xnor U6673 (N_6673,N_6582,N_6525);
xnor U6674 (N_6674,N_6552,N_6571);
nand U6675 (N_6675,N_6514,N_6538);
or U6676 (N_6676,N_6573,N_6551);
and U6677 (N_6677,N_6589,N_6542);
xor U6678 (N_6678,N_6539,N_6564);
xor U6679 (N_6679,N_6552,N_6553);
xor U6680 (N_6680,N_6584,N_6567);
and U6681 (N_6681,N_6512,N_6554);
nand U6682 (N_6682,N_6562,N_6599);
nor U6683 (N_6683,N_6507,N_6563);
nand U6684 (N_6684,N_6537,N_6529);
and U6685 (N_6685,N_6539,N_6528);
nand U6686 (N_6686,N_6580,N_6528);
and U6687 (N_6687,N_6561,N_6514);
nor U6688 (N_6688,N_6545,N_6502);
nor U6689 (N_6689,N_6503,N_6524);
and U6690 (N_6690,N_6538,N_6555);
nor U6691 (N_6691,N_6595,N_6585);
or U6692 (N_6692,N_6590,N_6506);
or U6693 (N_6693,N_6556,N_6562);
xor U6694 (N_6694,N_6595,N_6501);
nand U6695 (N_6695,N_6524,N_6573);
nand U6696 (N_6696,N_6503,N_6535);
nor U6697 (N_6697,N_6584,N_6518);
xor U6698 (N_6698,N_6540,N_6527);
or U6699 (N_6699,N_6551,N_6547);
nand U6700 (N_6700,N_6692,N_6652);
nor U6701 (N_6701,N_6660,N_6616);
and U6702 (N_6702,N_6640,N_6676);
and U6703 (N_6703,N_6653,N_6655);
nand U6704 (N_6704,N_6602,N_6609);
nor U6705 (N_6705,N_6647,N_6690);
or U6706 (N_6706,N_6693,N_6642);
xor U6707 (N_6707,N_6665,N_6645);
nor U6708 (N_6708,N_6674,N_6654);
and U6709 (N_6709,N_6648,N_6679);
and U6710 (N_6710,N_6614,N_6622);
nor U6711 (N_6711,N_6682,N_6694);
or U6712 (N_6712,N_6688,N_6662);
or U6713 (N_6713,N_6699,N_6631);
xor U6714 (N_6714,N_6658,N_6678);
nand U6715 (N_6715,N_6673,N_6683);
or U6716 (N_6716,N_6623,N_6601);
nor U6717 (N_6717,N_6638,N_6684);
nand U6718 (N_6718,N_6667,N_6636);
or U6719 (N_6719,N_6619,N_6677);
nand U6720 (N_6720,N_6620,N_6681);
nor U6721 (N_6721,N_6607,N_6628);
xnor U6722 (N_6722,N_6633,N_6613);
xnor U6723 (N_6723,N_6624,N_6625);
and U6724 (N_6724,N_6605,N_6666);
or U6725 (N_6725,N_6651,N_6695);
and U6726 (N_6726,N_6606,N_6663);
nor U6727 (N_6727,N_6618,N_6626);
xnor U6728 (N_6728,N_6696,N_6697);
or U6729 (N_6729,N_6680,N_6671);
xnor U6730 (N_6730,N_6643,N_6687);
or U6731 (N_6731,N_6670,N_6627);
or U6732 (N_6732,N_6604,N_6637);
or U6733 (N_6733,N_6639,N_6612);
and U6734 (N_6734,N_6685,N_6608);
or U6735 (N_6735,N_6600,N_6659);
nand U6736 (N_6736,N_6691,N_6646);
and U6737 (N_6737,N_6661,N_6689);
and U6738 (N_6738,N_6649,N_6644);
nand U6739 (N_6739,N_6672,N_6610);
or U6740 (N_6740,N_6656,N_6664);
or U6741 (N_6741,N_6657,N_6641);
and U6742 (N_6742,N_6686,N_6603);
nand U6743 (N_6743,N_6635,N_6611);
xor U6744 (N_6744,N_6615,N_6632);
xor U6745 (N_6745,N_6675,N_6668);
xor U6746 (N_6746,N_6621,N_6630);
xor U6747 (N_6747,N_6629,N_6634);
xnor U6748 (N_6748,N_6698,N_6669);
nor U6749 (N_6749,N_6650,N_6617);
or U6750 (N_6750,N_6612,N_6634);
and U6751 (N_6751,N_6679,N_6616);
and U6752 (N_6752,N_6631,N_6648);
nand U6753 (N_6753,N_6603,N_6682);
and U6754 (N_6754,N_6652,N_6612);
and U6755 (N_6755,N_6610,N_6641);
or U6756 (N_6756,N_6699,N_6614);
xor U6757 (N_6757,N_6673,N_6680);
and U6758 (N_6758,N_6682,N_6690);
xor U6759 (N_6759,N_6648,N_6671);
xnor U6760 (N_6760,N_6653,N_6623);
nor U6761 (N_6761,N_6616,N_6653);
and U6762 (N_6762,N_6698,N_6624);
xnor U6763 (N_6763,N_6670,N_6630);
nor U6764 (N_6764,N_6646,N_6667);
nor U6765 (N_6765,N_6660,N_6674);
nor U6766 (N_6766,N_6679,N_6670);
or U6767 (N_6767,N_6640,N_6601);
nand U6768 (N_6768,N_6628,N_6685);
or U6769 (N_6769,N_6692,N_6640);
or U6770 (N_6770,N_6687,N_6633);
nand U6771 (N_6771,N_6652,N_6661);
nor U6772 (N_6772,N_6622,N_6602);
and U6773 (N_6773,N_6620,N_6633);
nor U6774 (N_6774,N_6670,N_6671);
or U6775 (N_6775,N_6620,N_6652);
nand U6776 (N_6776,N_6656,N_6646);
xor U6777 (N_6777,N_6621,N_6693);
or U6778 (N_6778,N_6664,N_6624);
nand U6779 (N_6779,N_6654,N_6653);
nand U6780 (N_6780,N_6694,N_6667);
xnor U6781 (N_6781,N_6636,N_6674);
and U6782 (N_6782,N_6682,N_6675);
nor U6783 (N_6783,N_6600,N_6692);
nand U6784 (N_6784,N_6695,N_6666);
nand U6785 (N_6785,N_6673,N_6647);
xnor U6786 (N_6786,N_6671,N_6698);
nor U6787 (N_6787,N_6692,N_6620);
xnor U6788 (N_6788,N_6652,N_6617);
nand U6789 (N_6789,N_6641,N_6671);
or U6790 (N_6790,N_6621,N_6611);
nor U6791 (N_6791,N_6603,N_6608);
and U6792 (N_6792,N_6655,N_6695);
xnor U6793 (N_6793,N_6667,N_6635);
nor U6794 (N_6794,N_6696,N_6611);
nand U6795 (N_6795,N_6673,N_6687);
or U6796 (N_6796,N_6697,N_6695);
nand U6797 (N_6797,N_6614,N_6682);
xor U6798 (N_6798,N_6672,N_6693);
nand U6799 (N_6799,N_6621,N_6662);
and U6800 (N_6800,N_6777,N_6781);
or U6801 (N_6801,N_6721,N_6709);
nand U6802 (N_6802,N_6753,N_6778);
xor U6803 (N_6803,N_6724,N_6767);
nor U6804 (N_6804,N_6755,N_6776);
nor U6805 (N_6805,N_6723,N_6798);
nor U6806 (N_6806,N_6718,N_6751);
and U6807 (N_6807,N_6762,N_6726);
or U6808 (N_6808,N_6791,N_6748);
and U6809 (N_6809,N_6733,N_6711);
xor U6810 (N_6810,N_6713,N_6710);
nor U6811 (N_6811,N_6758,N_6764);
nor U6812 (N_6812,N_6719,N_6712);
xnor U6813 (N_6813,N_6770,N_6728);
nor U6814 (N_6814,N_6790,N_6704);
or U6815 (N_6815,N_6754,N_6717);
nand U6816 (N_6816,N_6722,N_6797);
xnor U6817 (N_6817,N_6759,N_6786);
and U6818 (N_6818,N_6732,N_6763);
and U6819 (N_6819,N_6730,N_6792);
xor U6820 (N_6820,N_6700,N_6741);
and U6821 (N_6821,N_6734,N_6775);
nor U6822 (N_6822,N_6756,N_6739);
or U6823 (N_6823,N_6746,N_6750);
nor U6824 (N_6824,N_6742,N_6774);
nand U6825 (N_6825,N_6773,N_6796);
and U6826 (N_6826,N_6771,N_6765);
xnor U6827 (N_6827,N_6725,N_6766);
and U6828 (N_6828,N_6727,N_6714);
nand U6829 (N_6829,N_6785,N_6706);
nor U6830 (N_6830,N_6716,N_6708);
nor U6831 (N_6831,N_6787,N_6743);
nor U6832 (N_6832,N_6788,N_6761);
and U6833 (N_6833,N_6740,N_6752);
and U6834 (N_6834,N_6735,N_6745);
or U6835 (N_6835,N_6782,N_6720);
nor U6836 (N_6836,N_6749,N_6789);
and U6837 (N_6837,N_6799,N_6736);
nor U6838 (N_6838,N_6731,N_6715);
or U6839 (N_6839,N_6779,N_6744);
nor U6840 (N_6840,N_6768,N_6784);
nand U6841 (N_6841,N_6793,N_6783);
nand U6842 (N_6842,N_6747,N_6701);
or U6843 (N_6843,N_6794,N_6705);
nor U6844 (N_6844,N_6780,N_6769);
or U6845 (N_6845,N_6757,N_6729);
and U6846 (N_6846,N_6772,N_6703);
nor U6847 (N_6847,N_6702,N_6760);
nand U6848 (N_6848,N_6737,N_6795);
or U6849 (N_6849,N_6738,N_6707);
and U6850 (N_6850,N_6762,N_6760);
and U6851 (N_6851,N_6747,N_6722);
nor U6852 (N_6852,N_6716,N_6700);
nor U6853 (N_6853,N_6793,N_6795);
and U6854 (N_6854,N_6734,N_6744);
or U6855 (N_6855,N_6784,N_6782);
nand U6856 (N_6856,N_6758,N_6728);
nand U6857 (N_6857,N_6743,N_6718);
xor U6858 (N_6858,N_6730,N_6771);
and U6859 (N_6859,N_6754,N_6779);
or U6860 (N_6860,N_6790,N_6776);
nand U6861 (N_6861,N_6776,N_6795);
nor U6862 (N_6862,N_6790,N_6726);
nor U6863 (N_6863,N_6727,N_6739);
nand U6864 (N_6864,N_6786,N_6772);
nand U6865 (N_6865,N_6734,N_6792);
or U6866 (N_6866,N_6778,N_6798);
or U6867 (N_6867,N_6735,N_6797);
nand U6868 (N_6868,N_6777,N_6737);
nand U6869 (N_6869,N_6782,N_6779);
nand U6870 (N_6870,N_6793,N_6773);
nor U6871 (N_6871,N_6756,N_6767);
and U6872 (N_6872,N_6700,N_6750);
nand U6873 (N_6873,N_6792,N_6797);
and U6874 (N_6874,N_6727,N_6758);
and U6875 (N_6875,N_6743,N_6727);
nand U6876 (N_6876,N_6702,N_6713);
and U6877 (N_6877,N_6714,N_6774);
or U6878 (N_6878,N_6779,N_6753);
nand U6879 (N_6879,N_6783,N_6761);
nand U6880 (N_6880,N_6782,N_6748);
and U6881 (N_6881,N_6748,N_6742);
nor U6882 (N_6882,N_6747,N_6727);
xnor U6883 (N_6883,N_6762,N_6770);
xnor U6884 (N_6884,N_6727,N_6713);
or U6885 (N_6885,N_6769,N_6775);
xnor U6886 (N_6886,N_6780,N_6725);
xor U6887 (N_6887,N_6775,N_6709);
xnor U6888 (N_6888,N_6791,N_6777);
nand U6889 (N_6889,N_6745,N_6747);
nor U6890 (N_6890,N_6792,N_6723);
and U6891 (N_6891,N_6795,N_6775);
and U6892 (N_6892,N_6750,N_6705);
or U6893 (N_6893,N_6773,N_6794);
nand U6894 (N_6894,N_6735,N_6789);
nor U6895 (N_6895,N_6773,N_6797);
and U6896 (N_6896,N_6785,N_6786);
xnor U6897 (N_6897,N_6791,N_6795);
xnor U6898 (N_6898,N_6709,N_6788);
nand U6899 (N_6899,N_6757,N_6792);
xor U6900 (N_6900,N_6824,N_6818);
or U6901 (N_6901,N_6899,N_6887);
nor U6902 (N_6902,N_6800,N_6884);
xor U6903 (N_6903,N_6817,N_6888);
and U6904 (N_6904,N_6809,N_6838);
and U6905 (N_6905,N_6839,N_6866);
nor U6906 (N_6906,N_6806,N_6804);
or U6907 (N_6907,N_6844,N_6815);
nor U6908 (N_6908,N_6871,N_6843);
nor U6909 (N_6909,N_6835,N_6827);
xor U6910 (N_6910,N_6857,N_6811);
nand U6911 (N_6911,N_6807,N_6851);
or U6912 (N_6912,N_6848,N_6833);
nor U6913 (N_6913,N_6813,N_6823);
and U6914 (N_6914,N_6802,N_6822);
xnor U6915 (N_6915,N_6841,N_6803);
or U6916 (N_6916,N_6886,N_6831);
nor U6917 (N_6917,N_6821,N_6840);
and U6918 (N_6918,N_6826,N_6830);
nor U6919 (N_6919,N_6863,N_6867);
xor U6920 (N_6920,N_6875,N_6868);
or U6921 (N_6921,N_6892,N_6864);
nand U6922 (N_6922,N_6889,N_6846);
and U6923 (N_6923,N_6865,N_6805);
and U6924 (N_6924,N_6891,N_6853);
nand U6925 (N_6925,N_6825,N_6856);
xor U6926 (N_6926,N_6885,N_6852);
or U6927 (N_6927,N_6810,N_6855);
xnor U6928 (N_6928,N_6819,N_6873);
or U6929 (N_6929,N_6862,N_6828);
or U6930 (N_6930,N_6820,N_6881);
nand U6931 (N_6931,N_6860,N_6869);
xor U6932 (N_6932,N_6883,N_6816);
nor U6933 (N_6933,N_6842,N_6898);
and U6934 (N_6934,N_6882,N_6834);
xor U6935 (N_6935,N_6854,N_6801);
nor U6936 (N_6936,N_6837,N_6876);
nor U6937 (N_6937,N_6858,N_6808);
xor U6938 (N_6938,N_6814,N_6894);
or U6939 (N_6939,N_6829,N_6877);
nor U6940 (N_6940,N_6845,N_6859);
xnor U6941 (N_6941,N_6861,N_6832);
xor U6942 (N_6942,N_6872,N_6890);
nor U6943 (N_6943,N_6847,N_6896);
nand U6944 (N_6944,N_6878,N_6880);
and U6945 (N_6945,N_6874,N_6849);
and U6946 (N_6946,N_6895,N_6893);
nand U6947 (N_6947,N_6850,N_6897);
xor U6948 (N_6948,N_6836,N_6879);
or U6949 (N_6949,N_6812,N_6870);
nor U6950 (N_6950,N_6831,N_6892);
xor U6951 (N_6951,N_6859,N_6806);
nor U6952 (N_6952,N_6806,N_6849);
nor U6953 (N_6953,N_6800,N_6843);
and U6954 (N_6954,N_6834,N_6856);
xor U6955 (N_6955,N_6850,N_6810);
xor U6956 (N_6956,N_6886,N_6869);
nor U6957 (N_6957,N_6861,N_6824);
or U6958 (N_6958,N_6871,N_6894);
nand U6959 (N_6959,N_6877,N_6880);
nand U6960 (N_6960,N_6880,N_6833);
nand U6961 (N_6961,N_6820,N_6884);
and U6962 (N_6962,N_6831,N_6851);
xnor U6963 (N_6963,N_6831,N_6860);
or U6964 (N_6964,N_6872,N_6814);
and U6965 (N_6965,N_6813,N_6815);
or U6966 (N_6966,N_6873,N_6860);
and U6967 (N_6967,N_6825,N_6869);
nand U6968 (N_6968,N_6832,N_6897);
nand U6969 (N_6969,N_6836,N_6883);
and U6970 (N_6970,N_6858,N_6813);
and U6971 (N_6971,N_6875,N_6891);
xor U6972 (N_6972,N_6835,N_6845);
xnor U6973 (N_6973,N_6837,N_6805);
nand U6974 (N_6974,N_6895,N_6823);
or U6975 (N_6975,N_6876,N_6842);
and U6976 (N_6976,N_6892,N_6805);
xor U6977 (N_6977,N_6855,N_6877);
and U6978 (N_6978,N_6819,N_6882);
or U6979 (N_6979,N_6849,N_6888);
and U6980 (N_6980,N_6810,N_6864);
and U6981 (N_6981,N_6855,N_6816);
and U6982 (N_6982,N_6809,N_6808);
nand U6983 (N_6983,N_6819,N_6831);
and U6984 (N_6984,N_6816,N_6838);
or U6985 (N_6985,N_6828,N_6876);
nor U6986 (N_6986,N_6810,N_6887);
and U6987 (N_6987,N_6831,N_6857);
or U6988 (N_6988,N_6800,N_6836);
xor U6989 (N_6989,N_6864,N_6808);
nand U6990 (N_6990,N_6835,N_6805);
xnor U6991 (N_6991,N_6804,N_6865);
and U6992 (N_6992,N_6821,N_6867);
nor U6993 (N_6993,N_6801,N_6897);
and U6994 (N_6994,N_6881,N_6899);
xnor U6995 (N_6995,N_6826,N_6800);
nand U6996 (N_6996,N_6887,N_6897);
or U6997 (N_6997,N_6855,N_6878);
xor U6998 (N_6998,N_6869,N_6839);
nor U6999 (N_6999,N_6826,N_6880);
nand U7000 (N_7000,N_6960,N_6925);
xnor U7001 (N_7001,N_6956,N_6947);
xnor U7002 (N_7002,N_6917,N_6904);
nor U7003 (N_7003,N_6971,N_6998);
nand U7004 (N_7004,N_6991,N_6906);
and U7005 (N_7005,N_6993,N_6930);
nor U7006 (N_7006,N_6989,N_6962);
nand U7007 (N_7007,N_6928,N_6986);
xnor U7008 (N_7008,N_6938,N_6963);
nand U7009 (N_7009,N_6927,N_6934);
or U7010 (N_7010,N_6935,N_6936);
xor U7011 (N_7011,N_6977,N_6918);
and U7012 (N_7012,N_6983,N_6913);
or U7013 (N_7013,N_6999,N_6952);
xnor U7014 (N_7014,N_6939,N_6900);
and U7015 (N_7015,N_6987,N_6980);
or U7016 (N_7016,N_6961,N_6955);
nor U7017 (N_7017,N_6968,N_6969);
nand U7018 (N_7018,N_6995,N_6910);
xor U7019 (N_7019,N_6972,N_6954);
xnor U7020 (N_7020,N_6981,N_6903);
and U7021 (N_7021,N_6951,N_6957);
nor U7022 (N_7022,N_6933,N_6997);
nor U7023 (N_7023,N_6929,N_6944);
and U7024 (N_7024,N_6905,N_6901);
or U7025 (N_7025,N_6978,N_6908);
or U7026 (N_7026,N_6911,N_6984);
or U7027 (N_7027,N_6996,N_6931);
nor U7028 (N_7028,N_6958,N_6920);
xor U7029 (N_7029,N_6945,N_6974);
nor U7030 (N_7030,N_6982,N_6975);
xnor U7031 (N_7031,N_6924,N_6902);
or U7032 (N_7032,N_6949,N_6976);
or U7033 (N_7033,N_6909,N_6959);
nand U7034 (N_7034,N_6946,N_6915);
nand U7035 (N_7035,N_6907,N_6914);
and U7036 (N_7036,N_6990,N_6966);
and U7037 (N_7037,N_6985,N_6994);
and U7038 (N_7038,N_6950,N_6923);
and U7039 (N_7039,N_6940,N_6992);
nor U7040 (N_7040,N_6937,N_6943);
or U7041 (N_7041,N_6967,N_6921);
or U7042 (N_7042,N_6988,N_6964);
xnor U7043 (N_7043,N_6916,N_6965);
nor U7044 (N_7044,N_6948,N_6970);
nand U7045 (N_7045,N_6922,N_6941);
nand U7046 (N_7046,N_6919,N_6953);
nor U7047 (N_7047,N_6973,N_6912);
nor U7048 (N_7048,N_6942,N_6932);
xnor U7049 (N_7049,N_6926,N_6979);
nand U7050 (N_7050,N_6947,N_6969);
or U7051 (N_7051,N_6939,N_6914);
or U7052 (N_7052,N_6931,N_6947);
xnor U7053 (N_7053,N_6949,N_6905);
xnor U7054 (N_7054,N_6944,N_6961);
and U7055 (N_7055,N_6955,N_6924);
or U7056 (N_7056,N_6917,N_6957);
and U7057 (N_7057,N_6929,N_6961);
nand U7058 (N_7058,N_6918,N_6964);
nor U7059 (N_7059,N_6998,N_6962);
and U7060 (N_7060,N_6914,N_6908);
nor U7061 (N_7061,N_6944,N_6927);
and U7062 (N_7062,N_6916,N_6903);
nor U7063 (N_7063,N_6914,N_6916);
nor U7064 (N_7064,N_6956,N_6908);
and U7065 (N_7065,N_6972,N_6905);
xor U7066 (N_7066,N_6940,N_6976);
or U7067 (N_7067,N_6973,N_6904);
nand U7068 (N_7068,N_6925,N_6964);
nand U7069 (N_7069,N_6982,N_6903);
nand U7070 (N_7070,N_6933,N_6959);
nor U7071 (N_7071,N_6944,N_6962);
and U7072 (N_7072,N_6936,N_6957);
and U7073 (N_7073,N_6970,N_6935);
xnor U7074 (N_7074,N_6950,N_6996);
nor U7075 (N_7075,N_6986,N_6945);
nor U7076 (N_7076,N_6948,N_6910);
and U7077 (N_7077,N_6979,N_6910);
nor U7078 (N_7078,N_6997,N_6911);
or U7079 (N_7079,N_6935,N_6963);
nand U7080 (N_7080,N_6923,N_6979);
nand U7081 (N_7081,N_6910,N_6951);
xnor U7082 (N_7082,N_6967,N_6969);
and U7083 (N_7083,N_6915,N_6974);
nor U7084 (N_7084,N_6954,N_6921);
nor U7085 (N_7085,N_6952,N_6991);
nand U7086 (N_7086,N_6924,N_6913);
xnor U7087 (N_7087,N_6971,N_6969);
nor U7088 (N_7088,N_6909,N_6944);
nand U7089 (N_7089,N_6999,N_6958);
and U7090 (N_7090,N_6978,N_6950);
nand U7091 (N_7091,N_6929,N_6922);
and U7092 (N_7092,N_6945,N_6938);
xor U7093 (N_7093,N_6958,N_6923);
or U7094 (N_7094,N_6901,N_6911);
or U7095 (N_7095,N_6907,N_6909);
nor U7096 (N_7096,N_6943,N_6956);
xor U7097 (N_7097,N_6909,N_6954);
or U7098 (N_7098,N_6914,N_6977);
and U7099 (N_7099,N_6992,N_6976);
xnor U7100 (N_7100,N_7033,N_7048);
nand U7101 (N_7101,N_7039,N_7088);
nor U7102 (N_7102,N_7031,N_7093);
or U7103 (N_7103,N_7069,N_7057);
nor U7104 (N_7104,N_7018,N_7014);
xor U7105 (N_7105,N_7073,N_7078);
and U7106 (N_7106,N_7094,N_7000);
or U7107 (N_7107,N_7012,N_7030);
or U7108 (N_7108,N_7004,N_7064);
xor U7109 (N_7109,N_7035,N_7063);
or U7110 (N_7110,N_7036,N_7008);
xor U7111 (N_7111,N_7041,N_7089);
xnor U7112 (N_7112,N_7087,N_7086);
and U7113 (N_7113,N_7074,N_7002);
xor U7114 (N_7114,N_7022,N_7023);
nor U7115 (N_7115,N_7019,N_7083);
and U7116 (N_7116,N_7043,N_7015);
nor U7117 (N_7117,N_7021,N_7052);
nor U7118 (N_7118,N_7013,N_7020);
and U7119 (N_7119,N_7034,N_7058);
or U7120 (N_7120,N_7075,N_7076);
xnor U7121 (N_7121,N_7079,N_7005);
and U7122 (N_7122,N_7090,N_7042);
and U7123 (N_7123,N_7062,N_7085);
and U7124 (N_7124,N_7028,N_7080);
nor U7125 (N_7125,N_7055,N_7016);
nand U7126 (N_7126,N_7096,N_7065);
xor U7127 (N_7127,N_7061,N_7007);
or U7128 (N_7128,N_7095,N_7092);
nor U7129 (N_7129,N_7040,N_7053);
or U7130 (N_7130,N_7091,N_7038);
and U7131 (N_7131,N_7060,N_7024);
or U7132 (N_7132,N_7082,N_7006);
or U7133 (N_7133,N_7081,N_7097);
nand U7134 (N_7134,N_7049,N_7017);
or U7135 (N_7135,N_7077,N_7027);
xor U7136 (N_7136,N_7011,N_7046);
and U7137 (N_7137,N_7068,N_7009);
nor U7138 (N_7138,N_7066,N_7054);
xor U7139 (N_7139,N_7056,N_7029);
or U7140 (N_7140,N_7072,N_7003);
nand U7141 (N_7141,N_7001,N_7098);
or U7142 (N_7142,N_7037,N_7084);
or U7143 (N_7143,N_7099,N_7032);
or U7144 (N_7144,N_7051,N_7025);
and U7145 (N_7145,N_7071,N_7050);
xnor U7146 (N_7146,N_7047,N_7026);
xnor U7147 (N_7147,N_7070,N_7010);
xor U7148 (N_7148,N_7044,N_7059);
nand U7149 (N_7149,N_7067,N_7045);
nor U7150 (N_7150,N_7057,N_7014);
and U7151 (N_7151,N_7098,N_7013);
or U7152 (N_7152,N_7089,N_7004);
xor U7153 (N_7153,N_7080,N_7099);
xnor U7154 (N_7154,N_7021,N_7088);
or U7155 (N_7155,N_7080,N_7020);
and U7156 (N_7156,N_7016,N_7022);
nand U7157 (N_7157,N_7021,N_7022);
nand U7158 (N_7158,N_7040,N_7004);
nor U7159 (N_7159,N_7070,N_7037);
and U7160 (N_7160,N_7061,N_7089);
nor U7161 (N_7161,N_7008,N_7050);
and U7162 (N_7162,N_7045,N_7042);
xor U7163 (N_7163,N_7057,N_7005);
or U7164 (N_7164,N_7063,N_7084);
xor U7165 (N_7165,N_7054,N_7020);
nor U7166 (N_7166,N_7093,N_7036);
or U7167 (N_7167,N_7048,N_7016);
nor U7168 (N_7168,N_7081,N_7099);
and U7169 (N_7169,N_7022,N_7059);
and U7170 (N_7170,N_7086,N_7028);
nor U7171 (N_7171,N_7070,N_7030);
nand U7172 (N_7172,N_7091,N_7004);
nor U7173 (N_7173,N_7056,N_7011);
nand U7174 (N_7174,N_7065,N_7007);
xnor U7175 (N_7175,N_7083,N_7079);
and U7176 (N_7176,N_7076,N_7009);
nor U7177 (N_7177,N_7035,N_7009);
or U7178 (N_7178,N_7054,N_7063);
or U7179 (N_7179,N_7040,N_7030);
or U7180 (N_7180,N_7074,N_7096);
xnor U7181 (N_7181,N_7095,N_7062);
nand U7182 (N_7182,N_7044,N_7063);
nand U7183 (N_7183,N_7069,N_7007);
and U7184 (N_7184,N_7046,N_7087);
nand U7185 (N_7185,N_7007,N_7084);
or U7186 (N_7186,N_7015,N_7002);
nor U7187 (N_7187,N_7073,N_7019);
and U7188 (N_7188,N_7013,N_7012);
nand U7189 (N_7189,N_7093,N_7038);
and U7190 (N_7190,N_7096,N_7039);
or U7191 (N_7191,N_7073,N_7027);
nand U7192 (N_7192,N_7076,N_7095);
and U7193 (N_7193,N_7051,N_7011);
xor U7194 (N_7194,N_7079,N_7036);
or U7195 (N_7195,N_7079,N_7010);
or U7196 (N_7196,N_7092,N_7015);
nand U7197 (N_7197,N_7075,N_7070);
xor U7198 (N_7198,N_7053,N_7051);
xnor U7199 (N_7199,N_7043,N_7033);
and U7200 (N_7200,N_7108,N_7195);
or U7201 (N_7201,N_7199,N_7184);
xnor U7202 (N_7202,N_7144,N_7192);
and U7203 (N_7203,N_7148,N_7131);
or U7204 (N_7204,N_7162,N_7155);
and U7205 (N_7205,N_7109,N_7194);
or U7206 (N_7206,N_7128,N_7169);
nand U7207 (N_7207,N_7165,N_7119);
xnor U7208 (N_7208,N_7193,N_7159);
and U7209 (N_7209,N_7117,N_7100);
nor U7210 (N_7210,N_7125,N_7187);
and U7211 (N_7211,N_7126,N_7175);
nor U7212 (N_7212,N_7145,N_7178);
nor U7213 (N_7213,N_7158,N_7181);
or U7214 (N_7214,N_7110,N_7141);
and U7215 (N_7215,N_7129,N_7133);
and U7216 (N_7216,N_7142,N_7152);
xor U7217 (N_7217,N_7147,N_7112);
nand U7218 (N_7218,N_7134,N_7157);
nor U7219 (N_7219,N_7156,N_7179);
nand U7220 (N_7220,N_7124,N_7171);
nand U7221 (N_7221,N_7137,N_7153);
nand U7222 (N_7222,N_7186,N_7170);
nor U7223 (N_7223,N_7174,N_7123);
nor U7224 (N_7224,N_7172,N_7149);
nand U7225 (N_7225,N_7166,N_7140);
or U7226 (N_7226,N_7150,N_7198);
nor U7227 (N_7227,N_7102,N_7146);
and U7228 (N_7228,N_7154,N_7116);
and U7229 (N_7229,N_7136,N_7167);
and U7230 (N_7230,N_7164,N_7130);
nand U7231 (N_7231,N_7188,N_7173);
or U7232 (N_7232,N_7160,N_7106);
nand U7233 (N_7233,N_7183,N_7127);
and U7234 (N_7234,N_7107,N_7118);
nor U7235 (N_7235,N_7139,N_7168);
and U7236 (N_7236,N_7115,N_7104);
or U7237 (N_7237,N_7182,N_7122);
nor U7238 (N_7238,N_7111,N_7143);
xnor U7239 (N_7239,N_7176,N_7103);
nor U7240 (N_7240,N_7113,N_7135);
or U7241 (N_7241,N_7191,N_7101);
or U7242 (N_7242,N_7161,N_7138);
xnor U7243 (N_7243,N_7196,N_7114);
or U7244 (N_7244,N_7185,N_7189);
xnor U7245 (N_7245,N_7120,N_7105);
xor U7246 (N_7246,N_7197,N_7132);
nand U7247 (N_7247,N_7177,N_7180);
and U7248 (N_7248,N_7163,N_7190);
xor U7249 (N_7249,N_7121,N_7151);
or U7250 (N_7250,N_7145,N_7140);
nand U7251 (N_7251,N_7130,N_7166);
nand U7252 (N_7252,N_7132,N_7166);
and U7253 (N_7253,N_7159,N_7120);
or U7254 (N_7254,N_7143,N_7199);
xor U7255 (N_7255,N_7181,N_7122);
nor U7256 (N_7256,N_7139,N_7122);
xor U7257 (N_7257,N_7134,N_7170);
nor U7258 (N_7258,N_7159,N_7107);
xnor U7259 (N_7259,N_7127,N_7100);
and U7260 (N_7260,N_7160,N_7166);
and U7261 (N_7261,N_7126,N_7181);
and U7262 (N_7262,N_7121,N_7147);
nor U7263 (N_7263,N_7172,N_7158);
nand U7264 (N_7264,N_7160,N_7116);
and U7265 (N_7265,N_7189,N_7153);
nor U7266 (N_7266,N_7194,N_7136);
xnor U7267 (N_7267,N_7152,N_7159);
or U7268 (N_7268,N_7131,N_7101);
and U7269 (N_7269,N_7194,N_7198);
nor U7270 (N_7270,N_7179,N_7152);
nand U7271 (N_7271,N_7169,N_7197);
xnor U7272 (N_7272,N_7137,N_7147);
and U7273 (N_7273,N_7139,N_7184);
xor U7274 (N_7274,N_7177,N_7102);
or U7275 (N_7275,N_7125,N_7130);
xnor U7276 (N_7276,N_7175,N_7100);
xnor U7277 (N_7277,N_7159,N_7123);
nor U7278 (N_7278,N_7160,N_7175);
or U7279 (N_7279,N_7169,N_7133);
or U7280 (N_7280,N_7188,N_7157);
nor U7281 (N_7281,N_7143,N_7151);
nor U7282 (N_7282,N_7162,N_7121);
or U7283 (N_7283,N_7188,N_7101);
or U7284 (N_7284,N_7161,N_7192);
or U7285 (N_7285,N_7171,N_7174);
xor U7286 (N_7286,N_7175,N_7153);
nand U7287 (N_7287,N_7158,N_7178);
or U7288 (N_7288,N_7109,N_7148);
xnor U7289 (N_7289,N_7117,N_7131);
nand U7290 (N_7290,N_7169,N_7136);
or U7291 (N_7291,N_7176,N_7113);
nor U7292 (N_7292,N_7187,N_7161);
xor U7293 (N_7293,N_7155,N_7165);
xor U7294 (N_7294,N_7154,N_7185);
xor U7295 (N_7295,N_7168,N_7192);
nand U7296 (N_7296,N_7134,N_7187);
nor U7297 (N_7297,N_7159,N_7157);
nand U7298 (N_7298,N_7124,N_7154);
or U7299 (N_7299,N_7106,N_7191);
nor U7300 (N_7300,N_7272,N_7281);
nand U7301 (N_7301,N_7261,N_7219);
xor U7302 (N_7302,N_7260,N_7273);
nand U7303 (N_7303,N_7295,N_7264);
or U7304 (N_7304,N_7287,N_7220);
and U7305 (N_7305,N_7248,N_7232);
nand U7306 (N_7306,N_7253,N_7278);
nor U7307 (N_7307,N_7262,N_7292);
nor U7308 (N_7308,N_7284,N_7231);
or U7309 (N_7309,N_7259,N_7211);
xor U7310 (N_7310,N_7228,N_7237);
nor U7311 (N_7311,N_7227,N_7297);
nand U7312 (N_7312,N_7214,N_7216);
or U7313 (N_7313,N_7263,N_7240);
nor U7314 (N_7314,N_7243,N_7271);
nand U7315 (N_7315,N_7223,N_7293);
or U7316 (N_7316,N_7277,N_7249);
and U7317 (N_7317,N_7267,N_7268);
nand U7318 (N_7318,N_7269,N_7285);
and U7319 (N_7319,N_7254,N_7200);
nor U7320 (N_7320,N_7244,N_7289);
nor U7321 (N_7321,N_7201,N_7245);
nand U7322 (N_7322,N_7270,N_7296);
and U7323 (N_7323,N_7283,N_7229);
xnor U7324 (N_7324,N_7218,N_7221);
nor U7325 (N_7325,N_7256,N_7239);
and U7326 (N_7326,N_7266,N_7246);
nor U7327 (N_7327,N_7291,N_7212);
xnor U7328 (N_7328,N_7265,N_7257);
or U7329 (N_7329,N_7238,N_7230);
and U7330 (N_7330,N_7217,N_7294);
and U7331 (N_7331,N_7242,N_7298);
xor U7332 (N_7332,N_7226,N_7209);
nand U7333 (N_7333,N_7222,N_7280);
and U7334 (N_7334,N_7250,N_7224);
or U7335 (N_7335,N_7235,N_7203);
xor U7336 (N_7336,N_7241,N_7275);
or U7337 (N_7337,N_7213,N_7252);
xor U7338 (N_7338,N_7233,N_7282);
and U7339 (N_7339,N_7207,N_7204);
nand U7340 (N_7340,N_7234,N_7258);
and U7341 (N_7341,N_7299,N_7290);
nor U7342 (N_7342,N_7255,N_7236);
nand U7343 (N_7343,N_7205,N_7286);
or U7344 (N_7344,N_7202,N_7276);
xor U7345 (N_7345,N_7208,N_7288);
nor U7346 (N_7346,N_7215,N_7225);
and U7347 (N_7347,N_7247,N_7274);
nor U7348 (N_7348,N_7206,N_7251);
xnor U7349 (N_7349,N_7279,N_7210);
xor U7350 (N_7350,N_7288,N_7253);
xor U7351 (N_7351,N_7274,N_7256);
xnor U7352 (N_7352,N_7283,N_7224);
nor U7353 (N_7353,N_7290,N_7214);
or U7354 (N_7354,N_7208,N_7206);
and U7355 (N_7355,N_7207,N_7210);
nor U7356 (N_7356,N_7212,N_7211);
nand U7357 (N_7357,N_7245,N_7255);
nor U7358 (N_7358,N_7203,N_7229);
or U7359 (N_7359,N_7251,N_7240);
nor U7360 (N_7360,N_7230,N_7214);
nor U7361 (N_7361,N_7240,N_7247);
nand U7362 (N_7362,N_7232,N_7217);
xnor U7363 (N_7363,N_7208,N_7260);
nor U7364 (N_7364,N_7284,N_7267);
or U7365 (N_7365,N_7221,N_7259);
or U7366 (N_7366,N_7254,N_7202);
xnor U7367 (N_7367,N_7275,N_7248);
nand U7368 (N_7368,N_7210,N_7227);
or U7369 (N_7369,N_7257,N_7247);
nand U7370 (N_7370,N_7200,N_7273);
and U7371 (N_7371,N_7212,N_7210);
nand U7372 (N_7372,N_7263,N_7231);
or U7373 (N_7373,N_7231,N_7259);
nor U7374 (N_7374,N_7241,N_7216);
and U7375 (N_7375,N_7295,N_7273);
or U7376 (N_7376,N_7239,N_7222);
nand U7377 (N_7377,N_7265,N_7295);
nor U7378 (N_7378,N_7215,N_7272);
and U7379 (N_7379,N_7241,N_7239);
xnor U7380 (N_7380,N_7220,N_7269);
nand U7381 (N_7381,N_7288,N_7217);
or U7382 (N_7382,N_7298,N_7218);
nor U7383 (N_7383,N_7287,N_7270);
nor U7384 (N_7384,N_7228,N_7265);
nor U7385 (N_7385,N_7214,N_7244);
xnor U7386 (N_7386,N_7296,N_7258);
xor U7387 (N_7387,N_7213,N_7204);
xor U7388 (N_7388,N_7235,N_7225);
nand U7389 (N_7389,N_7209,N_7289);
xor U7390 (N_7390,N_7255,N_7271);
nor U7391 (N_7391,N_7241,N_7298);
nor U7392 (N_7392,N_7240,N_7202);
or U7393 (N_7393,N_7272,N_7226);
nand U7394 (N_7394,N_7241,N_7279);
nor U7395 (N_7395,N_7221,N_7215);
or U7396 (N_7396,N_7266,N_7208);
and U7397 (N_7397,N_7216,N_7221);
nor U7398 (N_7398,N_7230,N_7283);
nor U7399 (N_7399,N_7247,N_7222);
nand U7400 (N_7400,N_7327,N_7369);
xor U7401 (N_7401,N_7348,N_7309);
xnor U7402 (N_7402,N_7347,N_7362);
xor U7403 (N_7403,N_7300,N_7301);
and U7404 (N_7404,N_7390,N_7345);
and U7405 (N_7405,N_7358,N_7383);
nand U7406 (N_7406,N_7312,N_7333);
or U7407 (N_7407,N_7357,N_7343);
or U7408 (N_7408,N_7307,N_7337);
nand U7409 (N_7409,N_7320,N_7316);
and U7410 (N_7410,N_7384,N_7395);
and U7411 (N_7411,N_7354,N_7322);
nand U7412 (N_7412,N_7341,N_7380);
and U7413 (N_7413,N_7356,N_7321);
nor U7414 (N_7414,N_7328,N_7325);
or U7415 (N_7415,N_7394,N_7391);
xor U7416 (N_7416,N_7388,N_7398);
nor U7417 (N_7417,N_7366,N_7386);
nor U7418 (N_7418,N_7304,N_7346);
nand U7419 (N_7419,N_7365,N_7389);
nand U7420 (N_7420,N_7311,N_7385);
nor U7421 (N_7421,N_7326,N_7360);
nand U7422 (N_7422,N_7373,N_7368);
nand U7423 (N_7423,N_7352,N_7315);
nand U7424 (N_7424,N_7313,N_7332);
nand U7425 (N_7425,N_7396,N_7397);
and U7426 (N_7426,N_7350,N_7367);
xor U7427 (N_7427,N_7355,N_7314);
xor U7428 (N_7428,N_7378,N_7305);
nor U7429 (N_7429,N_7364,N_7331);
and U7430 (N_7430,N_7340,N_7303);
xnor U7431 (N_7431,N_7387,N_7338);
and U7432 (N_7432,N_7336,N_7381);
nor U7433 (N_7433,N_7306,N_7324);
or U7434 (N_7434,N_7339,N_7330);
or U7435 (N_7435,N_7308,N_7363);
xor U7436 (N_7436,N_7329,N_7317);
nor U7437 (N_7437,N_7376,N_7323);
xnor U7438 (N_7438,N_7351,N_7370);
nand U7439 (N_7439,N_7335,N_7319);
nand U7440 (N_7440,N_7349,N_7371);
and U7441 (N_7441,N_7393,N_7359);
nand U7442 (N_7442,N_7344,N_7372);
and U7443 (N_7443,N_7375,N_7399);
or U7444 (N_7444,N_7392,N_7302);
or U7445 (N_7445,N_7342,N_7361);
nor U7446 (N_7446,N_7377,N_7353);
xor U7447 (N_7447,N_7334,N_7382);
xnor U7448 (N_7448,N_7374,N_7318);
nor U7449 (N_7449,N_7310,N_7379);
or U7450 (N_7450,N_7369,N_7351);
and U7451 (N_7451,N_7348,N_7359);
or U7452 (N_7452,N_7340,N_7317);
xor U7453 (N_7453,N_7350,N_7338);
and U7454 (N_7454,N_7393,N_7386);
xnor U7455 (N_7455,N_7379,N_7383);
and U7456 (N_7456,N_7348,N_7317);
nor U7457 (N_7457,N_7353,N_7349);
nor U7458 (N_7458,N_7328,N_7398);
xor U7459 (N_7459,N_7311,N_7339);
xnor U7460 (N_7460,N_7384,N_7381);
and U7461 (N_7461,N_7319,N_7365);
nor U7462 (N_7462,N_7358,N_7307);
nor U7463 (N_7463,N_7393,N_7310);
nand U7464 (N_7464,N_7323,N_7393);
nor U7465 (N_7465,N_7387,N_7325);
and U7466 (N_7466,N_7343,N_7310);
nor U7467 (N_7467,N_7388,N_7399);
or U7468 (N_7468,N_7366,N_7384);
nor U7469 (N_7469,N_7347,N_7360);
and U7470 (N_7470,N_7396,N_7390);
and U7471 (N_7471,N_7327,N_7380);
nor U7472 (N_7472,N_7361,N_7317);
and U7473 (N_7473,N_7370,N_7397);
nand U7474 (N_7474,N_7380,N_7379);
nand U7475 (N_7475,N_7326,N_7319);
xor U7476 (N_7476,N_7362,N_7315);
and U7477 (N_7477,N_7366,N_7362);
or U7478 (N_7478,N_7388,N_7397);
or U7479 (N_7479,N_7376,N_7339);
xnor U7480 (N_7480,N_7302,N_7347);
or U7481 (N_7481,N_7356,N_7394);
nand U7482 (N_7482,N_7344,N_7375);
xnor U7483 (N_7483,N_7324,N_7338);
or U7484 (N_7484,N_7326,N_7327);
and U7485 (N_7485,N_7355,N_7311);
or U7486 (N_7486,N_7328,N_7387);
or U7487 (N_7487,N_7312,N_7392);
or U7488 (N_7488,N_7320,N_7384);
nand U7489 (N_7489,N_7340,N_7323);
xor U7490 (N_7490,N_7311,N_7395);
nor U7491 (N_7491,N_7363,N_7328);
nand U7492 (N_7492,N_7344,N_7397);
xnor U7493 (N_7493,N_7365,N_7369);
and U7494 (N_7494,N_7377,N_7388);
xor U7495 (N_7495,N_7394,N_7319);
xnor U7496 (N_7496,N_7305,N_7319);
nor U7497 (N_7497,N_7385,N_7351);
nand U7498 (N_7498,N_7360,N_7381);
nor U7499 (N_7499,N_7398,N_7367);
or U7500 (N_7500,N_7445,N_7417);
xor U7501 (N_7501,N_7475,N_7453);
xnor U7502 (N_7502,N_7483,N_7401);
and U7503 (N_7503,N_7462,N_7406);
nand U7504 (N_7504,N_7457,N_7485);
nand U7505 (N_7505,N_7443,N_7431);
nand U7506 (N_7506,N_7478,N_7403);
nand U7507 (N_7507,N_7410,N_7470);
nor U7508 (N_7508,N_7471,N_7494);
or U7509 (N_7509,N_7492,N_7463);
nand U7510 (N_7510,N_7432,N_7455);
nand U7511 (N_7511,N_7473,N_7466);
nand U7512 (N_7512,N_7414,N_7450);
nand U7513 (N_7513,N_7416,N_7480);
and U7514 (N_7514,N_7418,N_7499);
nor U7515 (N_7515,N_7415,N_7440);
nand U7516 (N_7516,N_7451,N_7481);
and U7517 (N_7517,N_7434,N_7436);
xor U7518 (N_7518,N_7497,N_7468);
nor U7519 (N_7519,N_7422,N_7487);
xor U7520 (N_7520,N_7458,N_7449);
and U7521 (N_7521,N_7452,N_7444);
and U7522 (N_7522,N_7407,N_7459);
nor U7523 (N_7523,N_7430,N_7437);
and U7524 (N_7524,N_7493,N_7476);
or U7525 (N_7525,N_7454,N_7488);
xor U7526 (N_7526,N_7472,N_7448);
nor U7527 (N_7527,N_7429,N_7490);
and U7528 (N_7528,N_7439,N_7482);
nor U7529 (N_7529,N_7412,N_7477);
or U7530 (N_7530,N_7498,N_7424);
nand U7531 (N_7531,N_7479,N_7467);
and U7532 (N_7532,N_7427,N_7469);
nand U7533 (N_7533,N_7400,N_7404);
xor U7534 (N_7534,N_7408,N_7405);
xor U7535 (N_7535,N_7456,N_7433);
or U7536 (N_7536,N_7438,N_7495);
and U7537 (N_7537,N_7486,N_7496);
and U7538 (N_7538,N_7419,N_7489);
nor U7539 (N_7539,N_7465,N_7464);
and U7540 (N_7540,N_7409,N_7484);
and U7541 (N_7541,N_7474,N_7402);
and U7542 (N_7542,N_7426,N_7423);
nor U7543 (N_7543,N_7442,N_7435);
and U7544 (N_7544,N_7491,N_7460);
or U7545 (N_7545,N_7461,N_7411);
nand U7546 (N_7546,N_7447,N_7425);
nand U7547 (N_7547,N_7428,N_7441);
nor U7548 (N_7548,N_7446,N_7413);
or U7549 (N_7549,N_7421,N_7420);
nor U7550 (N_7550,N_7428,N_7445);
nand U7551 (N_7551,N_7454,N_7476);
nor U7552 (N_7552,N_7484,N_7457);
or U7553 (N_7553,N_7438,N_7463);
nand U7554 (N_7554,N_7468,N_7443);
xnor U7555 (N_7555,N_7497,N_7491);
nor U7556 (N_7556,N_7484,N_7430);
nand U7557 (N_7557,N_7436,N_7453);
nor U7558 (N_7558,N_7495,N_7466);
nor U7559 (N_7559,N_7404,N_7452);
nand U7560 (N_7560,N_7499,N_7434);
nand U7561 (N_7561,N_7433,N_7475);
nor U7562 (N_7562,N_7419,N_7420);
or U7563 (N_7563,N_7467,N_7451);
nor U7564 (N_7564,N_7460,N_7440);
nand U7565 (N_7565,N_7487,N_7454);
nand U7566 (N_7566,N_7412,N_7430);
xor U7567 (N_7567,N_7485,N_7492);
or U7568 (N_7568,N_7448,N_7443);
nand U7569 (N_7569,N_7469,N_7440);
nor U7570 (N_7570,N_7468,N_7440);
nor U7571 (N_7571,N_7403,N_7453);
nor U7572 (N_7572,N_7442,N_7433);
or U7573 (N_7573,N_7467,N_7404);
or U7574 (N_7574,N_7419,N_7427);
or U7575 (N_7575,N_7448,N_7439);
xor U7576 (N_7576,N_7437,N_7459);
nor U7577 (N_7577,N_7413,N_7417);
or U7578 (N_7578,N_7411,N_7430);
xor U7579 (N_7579,N_7436,N_7460);
xnor U7580 (N_7580,N_7448,N_7471);
and U7581 (N_7581,N_7436,N_7489);
xnor U7582 (N_7582,N_7420,N_7496);
nand U7583 (N_7583,N_7424,N_7490);
and U7584 (N_7584,N_7499,N_7487);
nand U7585 (N_7585,N_7448,N_7424);
and U7586 (N_7586,N_7474,N_7418);
xnor U7587 (N_7587,N_7447,N_7444);
xor U7588 (N_7588,N_7419,N_7495);
nand U7589 (N_7589,N_7470,N_7401);
xor U7590 (N_7590,N_7411,N_7468);
and U7591 (N_7591,N_7456,N_7430);
nand U7592 (N_7592,N_7479,N_7403);
xnor U7593 (N_7593,N_7497,N_7448);
xor U7594 (N_7594,N_7435,N_7448);
nand U7595 (N_7595,N_7421,N_7442);
and U7596 (N_7596,N_7472,N_7435);
and U7597 (N_7597,N_7423,N_7453);
xor U7598 (N_7598,N_7445,N_7427);
xor U7599 (N_7599,N_7401,N_7406);
nor U7600 (N_7600,N_7581,N_7580);
or U7601 (N_7601,N_7548,N_7554);
or U7602 (N_7602,N_7523,N_7525);
xor U7603 (N_7603,N_7555,N_7579);
or U7604 (N_7604,N_7589,N_7567);
and U7605 (N_7605,N_7512,N_7573);
xor U7606 (N_7606,N_7577,N_7516);
nor U7607 (N_7607,N_7500,N_7513);
or U7608 (N_7608,N_7578,N_7522);
xor U7609 (N_7609,N_7531,N_7596);
or U7610 (N_7610,N_7562,N_7545);
xor U7611 (N_7611,N_7569,N_7550);
nor U7612 (N_7612,N_7505,N_7535);
or U7613 (N_7613,N_7518,N_7566);
nand U7614 (N_7614,N_7585,N_7506);
nor U7615 (N_7615,N_7586,N_7540);
xnor U7616 (N_7616,N_7587,N_7539);
or U7617 (N_7617,N_7574,N_7519);
nand U7618 (N_7618,N_7538,N_7546);
xor U7619 (N_7619,N_7537,N_7572);
and U7620 (N_7620,N_7552,N_7597);
nand U7621 (N_7621,N_7558,N_7511);
and U7622 (N_7622,N_7590,N_7563);
and U7623 (N_7623,N_7588,N_7568);
and U7624 (N_7624,N_7593,N_7556);
nand U7625 (N_7625,N_7598,N_7583);
xnor U7626 (N_7626,N_7532,N_7526);
nand U7627 (N_7627,N_7507,N_7536);
nor U7628 (N_7628,N_7528,N_7527);
or U7629 (N_7629,N_7530,N_7551);
nor U7630 (N_7630,N_7515,N_7534);
and U7631 (N_7631,N_7520,N_7571);
or U7632 (N_7632,N_7521,N_7517);
nor U7633 (N_7633,N_7529,N_7564);
and U7634 (N_7634,N_7510,N_7504);
xnor U7635 (N_7635,N_7501,N_7584);
or U7636 (N_7636,N_7592,N_7541);
nor U7637 (N_7637,N_7576,N_7591);
nand U7638 (N_7638,N_7524,N_7594);
or U7639 (N_7639,N_7595,N_7582);
nand U7640 (N_7640,N_7502,N_7565);
xnor U7641 (N_7641,N_7599,N_7544);
nor U7642 (N_7642,N_7547,N_7503);
nor U7643 (N_7643,N_7543,N_7559);
nand U7644 (N_7644,N_7575,N_7508);
nand U7645 (N_7645,N_7549,N_7560);
and U7646 (N_7646,N_7570,N_7553);
nand U7647 (N_7647,N_7557,N_7533);
xnor U7648 (N_7648,N_7514,N_7542);
xor U7649 (N_7649,N_7509,N_7561);
nand U7650 (N_7650,N_7590,N_7597);
xnor U7651 (N_7651,N_7581,N_7508);
xnor U7652 (N_7652,N_7513,N_7523);
xnor U7653 (N_7653,N_7515,N_7594);
xnor U7654 (N_7654,N_7578,N_7513);
or U7655 (N_7655,N_7558,N_7553);
nor U7656 (N_7656,N_7567,N_7533);
or U7657 (N_7657,N_7540,N_7593);
nand U7658 (N_7658,N_7536,N_7510);
xnor U7659 (N_7659,N_7516,N_7568);
xnor U7660 (N_7660,N_7551,N_7556);
and U7661 (N_7661,N_7508,N_7523);
nor U7662 (N_7662,N_7534,N_7575);
nand U7663 (N_7663,N_7599,N_7583);
nor U7664 (N_7664,N_7540,N_7562);
or U7665 (N_7665,N_7589,N_7557);
nor U7666 (N_7666,N_7572,N_7564);
or U7667 (N_7667,N_7517,N_7550);
xor U7668 (N_7668,N_7573,N_7595);
and U7669 (N_7669,N_7562,N_7526);
or U7670 (N_7670,N_7550,N_7535);
xor U7671 (N_7671,N_7510,N_7513);
nor U7672 (N_7672,N_7509,N_7557);
nand U7673 (N_7673,N_7507,N_7561);
nand U7674 (N_7674,N_7510,N_7566);
nand U7675 (N_7675,N_7573,N_7557);
xnor U7676 (N_7676,N_7595,N_7566);
or U7677 (N_7677,N_7547,N_7557);
or U7678 (N_7678,N_7513,N_7518);
xor U7679 (N_7679,N_7581,N_7543);
nor U7680 (N_7680,N_7538,N_7557);
nand U7681 (N_7681,N_7500,N_7582);
nand U7682 (N_7682,N_7529,N_7541);
or U7683 (N_7683,N_7575,N_7528);
nor U7684 (N_7684,N_7587,N_7521);
and U7685 (N_7685,N_7535,N_7598);
nand U7686 (N_7686,N_7583,N_7522);
nor U7687 (N_7687,N_7519,N_7571);
or U7688 (N_7688,N_7552,N_7509);
or U7689 (N_7689,N_7577,N_7580);
nand U7690 (N_7690,N_7544,N_7507);
and U7691 (N_7691,N_7515,N_7578);
and U7692 (N_7692,N_7547,N_7539);
nor U7693 (N_7693,N_7560,N_7574);
or U7694 (N_7694,N_7509,N_7560);
or U7695 (N_7695,N_7568,N_7558);
nand U7696 (N_7696,N_7571,N_7532);
nor U7697 (N_7697,N_7512,N_7524);
and U7698 (N_7698,N_7597,N_7535);
nand U7699 (N_7699,N_7551,N_7553);
nor U7700 (N_7700,N_7682,N_7673);
xor U7701 (N_7701,N_7634,N_7695);
xnor U7702 (N_7702,N_7613,N_7606);
and U7703 (N_7703,N_7647,N_7637);
nor U7704 (N_7704,N_7697,N_7610);
nor U7705 (N_7705,N_7639,N_7638);
nor U7706 (N_7706,N_7633,N_7630);
xor U7707 (N_7707,N_7640,N_7650);
nor U7708 (N_7708,N_7642,N_7604);
or U7709 (N_7709,N_7632,N_7600);
and U7710 (N_7710,N_7698,N_7660);
xor U7711 (N_7711,N_7607,N_7693);
nor U7712 (N_7712,N_7685,N_7669);
and U7713 (N_7713,N_7629,N_7671);
nor U7714 (N_7714,N_7691,N_7676);
or U7715 (N_7715,N_7621,N_7663);
xor U7716 (N_7716,N_7684,N_7618);
nor U7717 (N_7717,N_7672,N_7615);
nor U7718 (N_7718,N_7611,N_7653);
xnor U7719 (N_7719,N_7661,N_7659);
xnor U7720 (N_7720,N_7623,N_7654);
nor U7721 (N_7721,N_7689,N_7687);
and U7722 (N_7722,N_7628,N_7631);
xnor U7723 (N_7723,N_7605,N_7688);
and U7724 (N_7724,N_7646,N_7614);
and U7725 (N_7725,N_7699,N_7649);
nor U7726 (N_7726,N_7664,N_7608);
nor U7727 (N_7727,N_7601,N_7690);
nor U7728 (N_7728,N_7619,N_7636);
xor U7729 (N_7729,N_7683,N_7666);
nor U7730 (N_7730,N_7680,N_7612);
or U7731 (N_7731,N_7617,N_7679);
nand U7732 (N_7732,N_7651,N_7674);
or U7733 (N_7733,N_7662,N_7655);
nor U7734 (N_7734,N_7622,N_7667);
nand U7735 (N_7735,N_7626,N_7668);
nand U7736 (N_7736,N_7620,N_7645);
nor U7737 (N_7737,N_7602,N_7624);
or U7738 (N_7738,N_7658,N_7652);
nand U7739 (N_7739,N_7616,N_7678);
nor U7740 (N_7740,N_7681,N_7670);
and U7741 (N_7741,N_7677,N_7603);
xnor U7742 (N_7742,N_7686,N_7692);
xor U7743 (N_7743,N_7644,N_7635);
and U7744 (N_7744,N_7694,N_7641);
xnor U7745 (N_7745,N_7656,N_7696);
and U7746 (N_7746,N_7657,N_7648);
or U7747 (N_7747,N_7627,N_7609);
xor U7748 (N_7748,N_7675,N_7625);
and U7749 (N_7749,N_7665,N_7643);
or U7750 (N_7750,N_7641,N_7643);
xor U7751 (N_7751,N_7616,N_7673);
and U7752 (N_7752,N_7642,N_7624);
nand U7753 (N_7753,N_7671,N_7681);
or U7754 (N_7754,N_7620,N_7684);
nor U7755 (N_7755,N_7657,N_7609);
xnor U7756 (N_7756,N_7624,N_7678);
nor U7757 (N_7757,N_7653,N_7607);
xnor U7758 (N_7758,N_7692,N_7604);
nand U7759 (N_7759,N_7632,N_7654);
nand U7760 (N_7760,N_7697,N_7659);
and U7761 (N_7761,N_7654,N_7645);
and U7762 (N_7762,N_7677,N_7635);
xnor U7763 (N_7763,N_7671,N_7649);
and U7764 (N_7764,N_7622,N_7669);
xor U7765 (N_7765,N_7673,N_7660);
or U7766 (N_7766,N_7628,N_7692);
nor U7767 (N_7767,N_7665,N_7687);
nor U7768 (N_7768,N_7663,N_7668);
nor U7769 (N_7769,N_7696,N_7664);
nor U7770 (N_7770,N_7648,N_7688);
and U7771 (N_7771,N_7692,N_7658);
or U7772 (N_7772,N_7627,N_7623);
nand U7773 (N_7773,N_7696,N_7669);
and U7774 (N_7774,N_7643,N_7681);
xnor U7775 (N_7775,N_7681,N_7625);
and U7776 (N_7776,N_7637,N_7627);
or U7777 (N_7777,N_7647,N_7690);
nand U7778 (N_7778,N_7681,N_7669);
nand U7779 (N_7779,N_7647,N_7629);
nor U7780 (N_7780,N_7667,N_7679);
nand U7781 (N_7781,N_7626,N_7612);
nand U7782 (N_7782,N_7660,N_7637);
nor U7783 (N_7783,N_7621,N_7688);
nor U7784 (N_7784,N_7622,N_7641);
xor U7785 (N_7785,N_7644,N_7628);
xor U7786 (N_7786,N_7618,N_7645);
and U7787 (N_7787,N_7609,N_7621);
nand U7788 (N_7788,N_7636,N_7671);
nor U7789 (N_7789,N_7611,N_7685);
nor U7790 (N_7790,N_7625,N_7661);
nand U7791 (N_7791,N_7625,N_7672);
and U7792 (N_7792,N_7634,N_7664);
and U7793 (N_7793,N_7657,N_7666);
nand U7794 (N_7794,N_7620,N_7644);
nor U7795 (N_7795,N_7672,N_7646);
and U7796 (N_7796,N_7607,N_7641);
nor U7797 (N_7797,N_7699,N_7625);
xnor U7798 (N_7798,N_7681,N_7619);
nor U7799 (N_7799,N_7604,N_7662);
and U7800 (N_7800,N_7729,N_7772);
nor U7801 (N_7801,N_7776,N_7794);
xor U7802 (N_7802,N_7744,N_7725);
nor U7803 (N_7803,N_7730,N_7710);
xor U7804 (N_7804,N_7752,N_7719);
nand U7805 (N_7805,N_7713,N_7749);
and U7806 (N_7806,N_7793,N_7784);
nand U7807 (N_7807,N_7785,N_7778);
nand U7808 (N_7808,N_7705,N_7704);
xnor U7809 (N_7809,N_7783,N_7773);
and U7810 (N_7810,N_7799,N_7766);
nand U7811 (N_7811,N_7709,N_7728);
and U7812 (N_7812,N_7796,N_7762);
xnor U7813 (N_7813,N_7781,N_7751);
nand U7814 (N_7814,N_7733,N_7764);
and U7815 (N_7815,N_7754,N_7715);
nand U7816 (N_7816,N_7753,N_7788);
nor U7817 (N_7817,N_7742,N_7708);
nand U7818 (N_7818,N_7774,N_7787);
nor U7819 (N_7819,N_7779,N_7792);
and U7820 (N_7820,N_7759,N_7797);
nand U7821 (N_7821,N_7747,N_7734);
and U7822 (N_7822,N_7724,N_7760);
nor U7823 (N_7823,N_7736,N_7743);
nor U7824 (N_7824,N_7727,N_7737);
nor U7825 (N_7825,N_7735,N_7732);
or U7826 (N_7826,N_7740,N_7791);
xor U7827 (N_7827,N_7789,N_7750);
nor U7828 (N_7828,N_7765,N_7720);
or U7829 (N_7829,N_7712,N_7717);
xor U7830 (N_7830,N_7738,N_7711);
nand U7831 (N_7831,N_7786,N_7771);
nand U7832 (N_7832,N_7706,N_7716);
and U7833 (N_7833,N_7777,N_7739);
and U7834 (N_7834,N_7767,N_7769);
and U7835 (N_7835,N_7722,N_7702);
and U7836 (N_7836,N_7726,N_7780);
xnor U7837 (N_7837,N_7761,N_7703);
nor U7838 (N_7838,N_7746,N_7756);
xor U7839 (N_7839,N_7748,N_7768);
xor U7840 (N_7840,N_7790,N_7718);
nor U7841 (N_7841,N_7798,N_7782);
xnor U7842 (N_7842,N_7755,N_7763);
nand U7843 (N_7843,N_7775,N_7741);
xnor U7844 (N_7844,N_7758,N_7700);
nor U7845 (N_7845,N_7795,N_7770);
nand U7846 (N_7846,N_7701,N_7721);
xnor U7847 (N_7847,N_7723,N_7707);
nor U7848 (N_7848,N_7714,N_7757);
and U7849 (N_7849,N_7731,N_7745);
nor U7850 (N_7850,N_7721,N_7799);
xnor U7851 (N_7851,N_7731,N_7753);
nor U7852 (N_7852,N_7732,N_7747);
and U7853 (N_7853,N_7748,N_7701);
or U7854 (N_7854,N_7741,N_7753);
nor U7855 (N_7855,N_7766,N_7790);
or U7856 (N_7856,N_7740,N_7750);
nand U7857 (N_7857,N_7789,N_7705);
or U7858 (N_7858,N_7755,N_7772);
nand U7859 (N_7859,N_7778,N_7775);
nand U7860 (N_7860,N_7752,N_7703);
nor U7861 (N_7861,N_7744,N_7745);
nand U7862 (N_7862,N_7752,N_7702);
nor U7863 (N_7863,N_7781,N_7748);
nand U7864 (N_7864,N_7725,N_7755);
or U7865 (N_7865,N_7739,N_7771);
nor U7866 (N_7866,N_7710,N_7793);
nand U7867 (N_7867,N_7799,N_7723);
nand U7868 (N_7868,N_7737,N_7790);
or U7869 (N_7869,N_7763,N_7740);
nand U7870 (N_7870,N_7719,N_7767);
nor U7871 (N_7871,N_7738,N_7772);
or U7872 (N_7872,N_7767,N_7765);
nand U7873 (N_7873,N_7713,N_7797);
nand U7874 (N_7874,N_7728,N_7773);
or U7875 (N_7875,N_7755,N_7708);
and U7876 (N_7876,N_7720,N_7776);
and U7877 (N_7877,N_7789,N_7758);
and U7878 (N_7878,N_7756,N_7767);
or U7879 (N_7879,N_7791,N_7778);
and U7880 (N_7880,N_7737,N_7785);
xnor U7881 (N_7881,N_7703,N_7791);
and U7882 (N_7882,N_7779,N_7798);
and U7883 (N_7883,N_7767,N_7746);
nand U7884 (N_7884,N_7750,N_7712);
nand U7885 (N_7885,N_7764,N_7736);
and U7886 (N_7886,N_7791,N_7772);
xor U7887 (N_7887,N_7729,N_7753);
or U7888 (N_7888,N_7744,N_7793);
nand U7889 (N_7889,N_7733,N_7763);
or U7890 (N_7890,N_7797,N_7702);
nor U7891 (N_7891,N_7771,N_7795);
or U7892 (N_7892,N_7728,N_7725);
nor U7893 (N_7893,N_7726,N_7736);
and U7894 (N_7894,N_7771,N_7770);
and U7895 (N_7895,N_7758,N_7770);
nor U7896 (N_7896,N_7764,N_7724);
xor U7897 (N_7897,N_7745,N_7759);
or U7898 (N_7898,N_7793,N_7747);
nand U7899 (N_7899,N_7779,N_7744);
or U7900 (N_7900,N_7815,N_7888);
xor U7901 (N_7901,N_7881,N_7858);
nand U7902 (N_7902,N_7812,N_7872);
and U7903 (N_7903,N_7877,N_7826);
xor U7904 (N_7904,N_7885,N_7871);
xor U7905 (N_7905,N_7863,N_7817);
nor U7906 (N_7906,N_7875,N_7879);
or U7907 (N_7907,N_7816,N_7894);
nand U7908 (N_7908,N_7827,N_7898);
xor U7909 (N_7909,N_7846,N_7839);
xnor U7910 (N_7910,N_7836,N_7819);
nor U7911 (N_7911,N_7849,N_7889);
nand U7912 (N_7912,N_7856,N_7837);
and U7913 (N_7913,N_7821,N_7848);
xnor U7914 (N_7914,N_7833,N_7800);
and U7915 (N_7915,N_7845,N_7825);
nor U7916 (N_7916,N_7862,N_7802);
nand U7917 (N_7917,N_7883,N_7835);
or U7918 (N_7918,N_7824,N_7810);
xnor U7919 (N_7919,N_7860,N_7880);
nand U7920 (N_7920,N_7866,N_7887);
and U7921 (N_7921,N_7808,N_7864);
xnor U7922 (N_7922,N_7809,N_7831);
nand U7923 (N_7923,N_7855,N_7818);
nor U7924 (N_7924,N_7851,N_7861);
xor U7925 (N_7925,N_7869,N_7896);
xnor U7926 (N_7926,N_7868,N_7854);
xnor U7927 (N_7927,N_7884,N_7850);
nand U7928 (N_7928,N_7857,N_7806);
xor U7929 (N_7929,N_7841,N_7899);
nand U7930 (N_7930,N_7801,N_7829);
or U7931 (N_7931,N_7867,N_7865);
or U7932 (N_7932,N_7844,N_7878);
nand U7933 (N_7933,N_7838,N_7822);
nand U7934 (N_7934,N_7840,N_7873);
and U7935 (N_7935,N_7842,N_7874);
or U7936 (N_7936,N_7853,N_7811);
or U7937 (N_7937,N_7813,N_7847);
nand U7938 (N_7938,N_7834,N_7807);
nand U7939 (N_7939,N_7886,N_7803);
nor U7940 (N_7940,N_7828,N_7859);
nor U7941 (N_7941,N_7820,N_7852);
nor U7942 (N_7942,N_7823,N_7832);
and U7943 (N_7943,N_7895,N_7893);
xnor U7944 (N_7944,N_7830,N_7876);
or U7945 (N_7945,N_7891,N_7890);
nand U7946 (N_7946,N_7897,N_7843);
nor U7947 (N_7947,N_7805,N_7870);
or U7948 (N_7948,N_7882,N_7892);
or U7949 (N_7949,N_7814,N_7804);
xor U7950 (N_7950,N_7847,N_7828);
nand U7951 (N_7951,N_7808,N_7830);
and U7952 (N_7952,N_7826,N_7802);
xor U7953 (N_7953,N_7817,N_7808);
xnor U7954 (N_7954,N_7843,N_7819);
or U7955 (N_7955,N_7825,N_7839);
xnor U7956 (N_7956,N_7837,N_7850);
xnor U7957 (N_7957,N_7813,N_7826);
nand U7958 (N_7958,N_7868,N_7866);
xor U7959 (N_7959,N_7812,N_7866);
or U7960 (N_7960,N_7897,N_7892);
and U7961 (N_7961,N_7810,N_7830);
and U7962 (N_7962,N_7832,N_7892);
and U7963 (N_7963,N_7888,N_7834);
nor U7964 (N_7964,N_7870,N_7809);
nor U7965 (N_7965,N_7891,N_7867);
xnor U7966 (N_7966,N_7854,N_7867);
or U7967 (N_7967,N_7886,N_7857);
nand U7968 (N_7968,N_7827,N_7882);
nand U7969 (N_7969,N_7889,N_7858);
xor U7970 (N_7970,N_7842,N_7852);
xnor U7971 (N_7971,N_7833,N_7891);
or U7972 (N_7972,N_7890,N_7824);
nand U7973 (N_7973,N_7838,N_7820);
nor U7974 (N_7974,N_7833,N_7874);
nand U7975 (N_7975,N_7849,N_7880);
nand U7976 (N_7976,N_7867,N_7853);
nor U7977 (N_7977,N_7822,N_7857);
and U7978 (N_7978,N_7854,N_7828);
xnor U7979 (N_7979,N_7842,N_7853);
and U7980 (N_7980,N_7820,N_7849);
or U7981 (N_7981,N_7827,N_7858);
and U7982 (N_7982,N_7809,N_7844);
and U7983 (N_7983,N_7821,N_7873);
nand U7984 (N_7984,N_7892,N_7845);
nand U7985 (N_7985,N_7865,N_7861);
or U7986 (N_7986,N_7876,N_7895);
and U7987 (N_7987,N_7829,N_7865);
nand U7988 (N_7988,N_7835,N_7809);
or U7989 (N_7989,N_7865,N_7836);
nor U7990 (N_7990,N_7811,N_7824);
xnor U7991 (N_7991,N_7839,N_7857);
nand U7992 (N_7992,N_7884,N_7897);
nand U7993 (N_7993,N_7877,N_7869);
nor U7994 (N_7994,N_7850,N_7862);
and U7995 (N_7995,N_7824,N_7866);
nor U7996 (N_7996,N_7868,N_7828);
nand U7997 (N_7997,N_7884,N_7835);
and U7998 (N_7998,N_7863,N_7832);
xnor U7999 (N_7999,N_7840,N_7819);
and U8000 (N_8000,N_7973,N_7993);
or U8001 (N_8001,N_7990,N_7984);
and U8002 (N_8002,N_7961,N_7992);
xor U8003 (N_8003,N_7935,N_7971);
and U8004 (N_8004,N_7979,N_7952);
or U8005 (N_8005,N_7912,N_7996);
xor U8006 (N_8006,N_7947,N_7983);
nor U8007 (N_8007,N_7970,N_7960);
nand U8008 (N_8008,N_7900,N_7958);
and U8009 (N_8009,N_7995,N_7927);
or U8010 (N_8010,N_7910,N_7968);
and U8011 (N_8011,N_7929,N_7928);
nand U8012 (N_8012,N_7914,N_7981);
and U8013 (N_8013,N_7966,N_7953);
nand U8014 (N_8014,N_7956,N_7909);
nand U8015 (N_8015,N_7962,N_7940);
xor U8016 (N_8016,N_7917,N_7916);
or U8017 (N_8017,N_7988,N_7902);
and U8018 (N_8018,N_7926,N_7906);
or U8019 (N_8019,N_7923,N_7938);
and U8020 (N_8020,N_7939,N_7964);
and U8021 (N_8021,N_7946,N_7904);
or U8022 (N_8022,N_7986,N_7982);
nand U8023 (N_8023,N_7974,N_7907);
nand U8024 (N_8024,N_7919,N_7959);
or U8025 (N_8025,N_7972,N_7915);
xnor U8026 (N_8026,N_7985,N_7955);
nor U8027 (N_8027,N_7976,N_7931);
and U8028 (N_8028,N_7941,N_7937);
xor U8029 (N_8029,N_7951,N_7994);
nor U8030 (N_8030,N_7965,N_7944);
nand U8031 (N_8031,N_7933,N_7921);
and U8032 (N_8032,N_7920,N_7963);
and U8033 (N_8033,N_7905,N_7945);
and U8034 (N_8034,N_7950,N_7980);
and U8035 (N_8035,N_7948,N_7975);
and U8036 (N_8036,N_7932,N_7936);
nand U8037 (N_8037,N_7911,N_7949);
nand U8038 (N_8038,N_7934,N_7977);
or U8039 (N_8039,N_7978,N_7925);
nor U8040 (N_8040,N_7991,N_7999);
or U8041 (N_8041,N_7943,N_7997);
nand U8042 (N_8042,N_7967,N_7987);
or U8043 (N_8043,N_7918,N_7989);
nand U8044 (N_8044,N_7969,N_7998);
or U8045 (N_8045,N_7903,N_7942);
nand U8046 (N_8046,N_7922,N_7924);
nand U8047 (N_8047,N_7954,N_7908);
nand U8048 (N_8048,N_7930,N_7957);
nor U8049 (N_8049,N_7901,N_7913);
nor U8050 (N_8050,N_7956,N_7930);
or U8051 (N_8051,N_7998,N_7901);
xor U8052 (N_8052,N_7910,N_7901);
or U8053 (N_8053,N_7968,N_7954);
nor U8054 (N_8054,N_7965,N_7927);
or U8055 (N_8055,N_7933,N_7956);
xor U8056 (N_8056,N_7978,N_7921);
or U8057 (N_8057,N_7988,N_7958);
nor U8058 (N_8058,N_7920,N_7933);
xnor U8059 (N_8059,N_7958,N_7970);
nor U8060 (N_8060,N_7901,N_7954);
or U8061 (N_8061,N_7961,N_7942);
or U8062 (N_8062,N_7987,N_7920);
and U8063 (N_8063,N_7925,N_7974);
or U8064 (N_8064,N_7949,N_7900);
or U8065 (N_8065,N_7903,N_7936);
xnor U8066 (N_8066,N_7978,N_7987);
or U8067 (N_8067,N_7995,N_7956);
and U8068 (N_8068,N_7968,N_7930);
xnor U8069 (N_8069,N_7935,N_7995);
and U8070 (N_8070,N_7934,N_7982);
nand U8071 (N_8071,N_7993,N_7975);
nand U8072 (N_8072,N_7983,N_7900);
nor U8073 (N_8073,N_7901,N_7932);
and U8074 (N_8074,N_7953,N_7971);
or U8075 (N_8075,N_7980,N_7997);
nand U8076 (N_8076,N_7969,N_7936);
or U8077 (N_8077,N_7920,N_7961);
nor U8078 (N_8078,N_7915,N_7976);
xor U8079 (N_8079,N_7901,N_7968);
xnor U8080 (N_8080,N_7965,N_7966);
or U8081 (N_8081,N_7910,N_7997);
and U8082 (N_8082,N_7929,N_7941);
or U8083 (N_8083,N_7950,N_7998);
or U8084 (N_8084,N_7950,N_7993);
nor U8085 (N_8085,N_7924,N_7969);
xor U8086 (N_8086,N_7969,N_7987);
xnor U8087 (N_8087,N_7921,N_7991);
nor U8088 (N_8088,N_7971,N_7982);
nor U8089 (N_8089,N_7966,N_7971);
or U8090 (N_8090,N_7913,N_7904);
xnor U8091 (N_8091,N_7901,N_7904);
nor U8092 (N_8092,N_7919,N_7985);
or U8093 (N_8093,N_7975,N_7926);
nor U8094 (N_8094,N_7977,N_7925);
xnor U8095 (N_8095,N_7908,N_7939);
nand U8096 (N_8096,N_7911,N_7973);
nor U8097 (N_8097,N_7914,N_7950);
or U8098 (N_8098,N_7983,N_7967);
and U8099 (N_8099,N_7906,N_7947);
xor U8100 (N_8100,N_8053,N_8017);
and U8101 (N_8101,N_8098,N_8087);
nand U8102 (N_8102,N_8084,N_8011);
or U8103 (N_8103,N_8035,N_8020);
nand U8104 (N_8104,N_8019,N_8080);
xnor U8105 (N_8105,N_8096,N_8081);
and U8106 (N_8106,N_8075,N_8063);
nor U8107 (N_8107,N_8003,N_8008);
and U8108 (N_8108,N_8042,N_8085);
xnor U8109 (N_8109,N_8045,N_8072);
or U8110 (N_8110,N_8016,N_8023);
xor U8111 (N_8111,N_8059,N_8010);
and U8112 (N_8112,N_8088,N_8031);
and U8113 (N_8113,N_8090,N_8050);
or U8114 (N_8114,N_8047,N_8041);
xnor U8115 (N_8115,N_8057,N_8015);
or U8116 (N_8116,N_8060,N_8044);
xor U8117 (N_8117,N_8036,N_8027);
nand U8118 (N_8118,N_8022,N_8025);
nor U8119 (N_8119,N_8056,N_8094);
xnor U8120 (N_8120,N_8055,N_8054);
xnor U8121 (N_8121,N_8069,N_8073);
or U8122 (N_8122,N_8074,N_8005);
or U8123 (N_8123,N_8043,N_8086);
nor U8124 (N_8124,N_8079,N_8061);
nor U8125 (N_8125,N_8026,N_8082);
or U8126 (N_8126,N_8030,N_8000);
nor U8127 (N_8127,N_8049,N_8032);
xor U8128 (N_8128,N_8024,N_8038);
nand U8129 (N_8129,N_8046,N_8018);
nand U8130 (N_8130,N_8012,N_8052);
xor U8131 (N_8131,N_8062,N_8070);
xor U8132 (N_8132,N_8078,N_8083);
xnor U8133 (N_8133,N_8068,N_8028);
xnor U8134 (N_8134,N_8095,N_8029);
nor U8135 (N_8135,N_8064,N_8065);
and U8136 (N_8136,N_8037,N_8009);
nor U8137 (N_8137,N_8077,N_8089);
xor U8138 (N_8138,N_8058,N_8051);
and U8139 (N_8139,N_8091,N_8066);
or U8140 (N_8140,N_8039,N_8076);
or U8141 (N_8141,N_8097,N_8007);
or U8142 (N_8142,N_8033,N_8048);
xor U8143 (N_8143,N_8034,N_8006);
nor U8144 (N_8144,N_8071,N_8067);
nand U8145 (N_8145,N_8092,N_8004);
nor U8146 (N_8146,N_8001,N_8021);
nor U8147 (N_8147,N_8040,N_8014);
or U8148 (N_8148,N_8013,N_8093);
xor U8149 (N_8149,N_8002,N_8099);
or U8150 (N_8150,N_8022,N_8010);
and U8151 (N_8151,N_8071,N_8097);
nor U8152 (N_8152,N_8007,N_8014);
or U8153 (N_8153,N_8042,N_8078);
xor U8154 (N_8154,N_8035,N_8001);
and U8155 (N_8155,N_8033,N_8014);
xnor U8156 (N_8156,N_8032,N_8083);
and U8157 (N_8157,N_8090,N_8015);
nand U8158 (N_8158,N_8007,N_8051);
or U8159 (N_8159,N_8028,N_8033);
and U8160 (N_8160,N_8019,N_8027);
and U8161 (N_8161,N_8080,N_8025);
or U8162 (N_8162,N_8001,N_8043);
and U8163 (N_8163,N_8064,N_8059);
xnor U8164 (N_8164,N_8014,N_8041);
nor U8165 (N_8165,N_8063,N_8081);
nor U8166 (N_8166,N_8014,N_8029);
or U8167 (N_8167,N_8085,N_8064);
xnor U8168 (N_8168,N_8035,N_8066);
nand U8169 (N_8169,N_8050,N_8088);
nand U8170 (N_8170,N_8010,N_8055);
nand U8171 (N_8171,N_8082,N_8036);
nor U8172 (N_8172,N_8098,N_8007);
xor U8173 (N_8173,N_8038,N_8048);
nor U8174 (N_8174,N_8058,N_8042);
nor U8175 (N_8175,N_8027,N_8032);
nor U8176 (N_8176,N_8016,N_8050);
xor U8177 (N_8177,N_8025,N_8052);
xor U8178 (N_8178,N_8024,N_8048);
and U8179 (N_8179,N_8084,N_8087);
nand U8180 (N_8180,N_8032,N_8078);
and U8181 (N_8181,N_8001,N_8097);
and U8182 (N_8182,N_8069,N_8015);
or U8183 (N_8183,N_8074,N_8055);
or U8184 (N_8184,N_8029,N_8023);
nand U8185 (N_8185,N_8035,N_8002);
nor U8186 (N_8186,N_8083,N_8092);
nand U8187 (N_8187,N_8056,N_8049);
and U8188 (N_8188,N_8018,N_8077);
or U8189 (N_8189,N_8059,N_8045);
nand U8190 (N_8190,N_8066,N_8083);
xor U8191 (N_8191,N_8050,N_8035);
or U8192 (N_8192,N_8076,N_8036);
or U8193 (N_8193,N_8034,N_8088);
and U8194 (N_8194,N_8056,N_8027);
nand U8195 (N_8195,N_8083,N_8003);
xor U8196 (N_8196,N_8077,N_8049);
or U8197 (N_8197,N_8094,N_8079);
nor U8198 (N_8198,N_8050,N_8042);
or U8199 (N_8199,N_8092,N_8010);
or U8200 (N_8200,N_8138,N_8166);
nor U8201 (N_8201,N_8145,N_8106);
xor U8202 (N_8202,N_8144,N_8126);
nand U8203 (N_8203,N_8162,N_8109);
xor U8204 (N_8204,N_8174,N_8150);
xnor U8205 (N_8205,N_8100,N_8131);
or U8206 (N_8206,N_8123,N_8197);
nand U8207 (N_8207,N_8121,N_8198);
nor U8208 (N_8208,N_8177,N_8116);
or U8209 (N_8209,N_8103,N_8194);
and U8210 (N_8210,N_8153,N_8122);
xnor U8211 (N_8211,N_8124,N_8182);
and U8212 (N_8212,N_8196,N_8112);
xnor U8213 (N_8213,N_8193,N_8108);
nand U8214 (N_8214,N_8148,N_8159);
or U8215 (N_8215,N_8120,N_8175);
xnor U8216 (N_8216,N_8139,N_8142);
nand U8217 (N_8217,N_8141,N_8164);
and U8218 (N_8218,N_8195,N_8189);
and U8219 (N_8219,N_8115,N_8155);
nor U8220 (N_8220,N_8190,N_8140);
nor U8221 (N_8221,N_8171,N_8149);
nand U8222 (N_8222,N_8188,N_8118);
or U8223 (N_8223,N_8170,N_8101);
xnor U8224 (N_8224,N_8178,N_8119);
and U8225 (N_8225,N_8161,N_8179);
xnor U8226 (N_8226,N_8152,N_8133);
nand U8227 (N_8227,N_8151,N_8176);
or U8228 (N_8228,N_8110,N_8134);
and U8229 (N_8229,N_8163,N_8117);
nor U8230 (N_8230,N_8147,N_8154);
nand U8231 (N_8231,N_8192,N_8167);
nor U8232 (N_8232,N_8185,N_8136);
xnor U8233 (N_8233,N_8113,N_8107);
nand U8234 (N_8234,N_8199,N_8184);
or U8235 (N_8235,N_8180,N_8172);
and U8236 (N_8236,N_8157,N_8130);
nand U8237 (N_8237,N_8181,N_8125);
xnor U8238 (N_8238,N_8111,N_8105);
nor U8239 (N_8239,N_8165,N_8169);
nor U8240 (N_8240,N_8135,N_8128);
or U8241 (N_8241,N_8102,N_8143);
and U8242 (N_8242,N_8160,N_8114);
and U8243 (N_8243,N_8191,N_8158);
and U8244 (N_8244,N_8168,N_8183);
and U8245 (N_8245,N_8104,N_8187);
nor U8246 (N_8246,N_8186,N_8132);
nand U8247 (N_8247,N_8146,N_8129);
nor U8248 (N_8248,N_8127,N_8156);
nand U8249 (N_8249,N_8137,N_8173);
or U8250 (N_8250,N_8170,N_8127);
nor U8251 (N_8251,N_8125,N_8195);
xor U8252 (N_8252,N_8148,N_8166);
or U8253 (N_8253,N_8156,N_8117);
xor U8254 (N_8254,N_8130,N_8149);
nand U8255 (N_8255,N_8177,N_8117);
nand U8256 (N_8256,N_8119,N_8122);
or U8257 (N_8257,N_8148,N_8111);
or U8258 (N_8258,N_8140,N_8166);
nand U8259 (N_8259,N_8133,N_8164);
nand U8260 (N_8260,N_8152,N_8198);
or U8261 (N_8261,N_8108,N_8191);
and U8262 (N_8262,N_8160,N_8153);
nand U8263 (N_8263,N_8178,N_8124);
nor U8264 (N_8264,N_8144,N_8169);
or U8265 (N_8265,N_8164,N_8123);
nor U8266 (N_8266,N_8119,N_8191);
nor U8267 (N_8267,N_8124,N_8126);
or U8268 (N_8268,N_8115,N_8134);
xor U8269 (N_8269,N_8144,N_8146);
nor U8270 (N_8270,N_8151,N_8106);
nand U8271 (N_8271,N_8108,N_8177);
and U8272 (N_8272,N_8177,N_8195);
and U8273 (N_8273,N_8125,N_8144);
or U8274 (N_8274,N_8196,N_8194);
or U8275 (N_8275,N_8150,N_8169);
xor U8276 (N_8276,N_8195,N_8134);
and U8277 (N_8277,N_8170,N_8118);
nand U8278 (N_8278,N_8144,N_8166);
nor U8279 (N_8279,N_8172,N_8113);
nor U8280 (N_8280,N_8195,N_8188);
and U8281 (N_8281,N_8172,N_8159);
or U8282 (N_8282,N_8167,N_8129);
and U8283 (N_8283,N_8139,N_8174);
and U8284 (N_8284,N_8137,N_8129);
and U8285 (N_8285,N_8170,N_8190);
xor U8286 (N_8286,N_8165,N_8166);
nor U8287 (N_8287,N_8167,N_8126);
or U8288 (N_8288,N_8183,N_8146);
nor U8289 (N_8289,N_8193,N_8129);
and U8290 (N_8290,N_8191,N_8148);
nor U8291 (N_8291,N_8133,N_8117);
and U8292 (N_8292,N_8123,N_8104);
or U8293 (N_8293,N_8163,N_8176);
or U8294 (N_8294,N_8149,N_8196);
or U8295 (N_8295,N_8193,N_8199);
xnor U8296 (N_8296,N_8183,N_8170);
nand U8297 (N_8297,N_8170,N_8191);
nand U8298 (N_8298,N_8121,N_8130);
nor U8299 (N_8299,N_8180,N_8109);
or U8300 (N_8300,N_8255,N_8213);
xor U8301 (N_8301,N_8241,N_8275);
xor U8302 (N_8302,N_8283,N_8203);
nand U8303 (N_8303,N_8209,N_8287);
and U8304 (N_8304,N_8254,N_8238);
and U8305 (N_8305,N_8274,N_8273);
or U8306 (N_8306,N_8223,N_8221);
nor U8307 (N_8307,N_8211,N_8262);
nand U8308 (N_8308,N_8281,N_8233);
and U8309 (N_8309,N_8215,N_8280);
nand U8310 (N_8310,N_8200,N_8210);
and U8311 (N_8311,N_8244,N_8252);
or U8312 (N_8312,N_8243,N_8272);
xnor U8313 (N_8313,N_8296,N_8239);
and U8314 (N_8314,N_8284,N_8253);
or U8315 (N_8315,N_8240,N_8257);
nor U8316 (N_8316,N_8218,N_8246);
nor U8317 (N_8317,N_8299,N_8286);
or U8318 (N_8318,N_8270,N_8277);
and U8319 (N_8319,N_8228,N_8290);
nor U8320 (N_8320,N_8294,N_8263);
nand U8321 (N_8321,N_8226,N_8234);
or U8322 (N_8322,N_8245,N_8242);
nor U8323 (N_8323,N_8267,N_8265);
or U8324 (N_8324,N_8248,N_8251);
or U8325 (N_8325,N_8224,N_8208);
or U8326 (N_8326,N_8297,N_8269);
and U8327 (N_8327,N_8202,N_8235);
nor U8328 (N_8328,N_8207,N_8229);
and U8329 (N_8329,N_8285,N_8279);
nand U8330 (N_8330,N_8266,N_8205);
xnor U8331 (N_8331,N_8217,N_8288);
or U8332 (N_8332,N_8249,N_8291);
and U8333 (N_8333,N_8292,N_8259);
nand U8334 (N_8334,N_8227,N_8220);
nor U8335 (N_8335,N_8236,N_8264);
or U8336 (N_8336,N_8271,N_8225);
nor U8337 (N_8337,N_8261,N_8230);
and U8338 (N_8338,N_8214,N_8216);
xor U8339 (N_8339,N_8276,N_8258);
and U8340 (N_8340,N_8278,N_8222);
or U8341 (N_8341,N_8295,N_8204);
or U8342 (N_8342,N_8231,N_8237);
or U8343 (N_8343,N_8250,N_8232);
and U8344 (N_8344,N_8260,N_8298);
nand U8345 (N_8345,N_8289,N_8206);
nor U8346 (N_8346,N_8282,N_8268);
nor U8347 (N_8347,N_8256,N_8219);
xor U8348 (N_8348,N_8201,N_8212);
or U8349 (N_8349,N_8293,N_8247);
nand U8350 (N_8350,N_8200,N_8297);
and U8351 (N_8351,N_8258,N_8213);
or U8352 (N_8352,N_8207,N_8271);
nand U8353 (N_8353,N_8299,N_8288);
nor U8354 (N_8354,N_8291,N_8218);
xor U8355 (N_8355,N_8222,N_8254);
or U8356 (N_8356,N_8208,N_8268);
xnor U8357 (N_8357,N_8212,N_8287);
or U8358 (N_8358,N_8216,N_8260);
and U8359 (N_8359,N_8285,N_8292);
and U8360 (N_8360,N_8282,N_8273);
xnor U8361 (N_8361,N_8239,N_8286);
or U8362 (N_8362,N_8281,N_8219);
or U8363 (N_8363,N_8213,N_8284);
nand U8364 (N_8364,N_8204,N_8255);
nor U8365 (N_8365,N_8283,N_8244);
nand U8366 (N_8366,N_8281,N_8208);
nand U8367 (N_8367,N_8223,N_8263);
and U8368 (N_8368,N_8242,N_8285);
and U8369 (N_8369,N_8226,N_8213);
xor U8370 (N_8370,N_8242,N_8255);
or U8371 (N_8371,N_8263,N_8260);
and U8372 (N_8372,N_8208,N_8295);
or U8373 (N_8373,N_8203,N_8256);
and U8374 (N_8374,N_8246,N_8210);
or U8375 (N_8375,N_8255,N_8264);
and U8376 (N_8376,N_8244,N_8248);
nand U8377 (N_8377,N_8210,N_8203);
or U8378 (N_8378,N_8224,N_8281);
nor U8379 (N_8379,N_8298,N_8228);
nand U8380 (N_8380,N_8286,N_8276);
nor U8381 (N_8381,N_8265,N_8208);
xor U8382 (N_8382,N_8264,N_8287);
or U8383 (N_8383,N_8259,N_8253);
or U8384 (N_8384,N_8201,N_8250);
xnor U8385 (N_8385,N_8222,N_8244);
nor U8386 (N_8386,N_8291,N_8254);
or U8387 (N_8387,N_8295,N_8218);
xnor U8388 (N_8388,N_8222,N_8242);
and U8389 (N_8389,N_8216,N_8296);
and U8390 (N_8390,N_8204,N_8294);
or U8391 (N_8391,N_8205,N_8234);
and U8392 (N_8392,N_8214,N_8263);
xor U8393 (N_8393,N_8265,N_8202);
nor U8394 (N_8394,N_8215,N_8220);
or U8395 (N_8395,N_8233,N_8226);
nand U8396 (N_8396,N_8237,N_8254);
nor U8397 (N_8397,N_8239,N_8285);
nor U8398 (N_8398,N_8273,N_8216);
or U8399 (N_8399,N_8253,N_8222);
nand U8400 (N_8400,N_8354,N_8379);
nor U8401 (N_8401,N_8327,N_8326);
nand U8402 (N_8402,N_8399,N_8374);
and U8403 (N_8403,N_8306,N_8325);
or U8404 (N_8404,N_8303,N_8360);
or U8405 (N_8405,N_8378,N_8345);
nor U8406 (N_8406,N_8311,N_8355);
and U8407 (N_8407,N_8371,N_8336);
nor U8408 (N_8408,N_8319,N_8361);
nand U8409 (N_8409,N_8353,N_8337);
nor U8410 (N_8410,N_8349,N_8352);
or U8411 (N_8411,N_8383,N_8387);
and U8412 (N_8412,N_8365,N_8362);
nor U8413 (N_8413,N_8318,N_8348);
and U8414 (N_8414,N_8305,N_8376);
nand U8415 (N_8415,N_8312,N_8330);
xnor U8416 (N_8416,N_8366,N_8307);
xor U8417 (N_8417,N_8363,N_8394);
and U8418 (N_8418,N_8390,N_8388);
and U8419 (N_8419,N_8364,N_8396);
and U8420 (N_8420,N_8304,N_8301);
or U8421 (N_8421,N_8351,N_8315);
and U8422 (N_8422,N_8358,N_8323);
nor U8423 (N_8423,N_8367,N_8313);
nand U8424 (N_8424,N_8309,N_8391);
nand U8425 (N_8425,N_8393,N_8386);
or U8426 (N_8426,N_8370,N_8316);
xnor U8427 (N_8427,N_8310,N_8369);
xor U8428 (N_8428,N_8302,N_8317);
xnor U8429 (N_8429,N_8324,N_8356);
xnor U8430 (N_8430,N_8368,N_8389);
and U8431 (N_8431,N_8333,N_8342);
nand U8432 (N_8432,N_8321,N_8340);
nor U8433 (N_8433,N_8346,N_8377);
or U8434 (N_8434,N_8357,N_8344);
or U8435 (N_8435,N_8384,N_8343);
and U8436 (N_8436,N_8300,N_8339);
and U8437 (N_8437,N_8380,N_8398);
and U8438 (N_8438,N_8373,N_8372);
xor U8439 (N_8439,N_8341,N_8335);
nor U8440 (N_8440,N_8338,N_8329);
and U8441 (N_8441,N_8308,N_8359);
nand U8442 (N_8442,N_8332,N_8375);
xnor U8443 (N_8443,N_8350,N_8392);
and U8444 (N_8444,N_8331,N_8385);
nand U8445 (N_8445,N_8397,N_8382);
and U8446 (N_8446,N_8334,N_8328);
and U8447 (N_8447,N_8320,N_8322);
nor U8448 (N_8448,N_8347,N_8381);
or U8449 (N_8449,N_8395,N_8314);
nor U8450 (N_8450,N_8367,N_8388);
and U8451 (N_8451,N_8393,N_8353);
nor U8452 (N_8452,N_8322,N_8338);
and U8453 (N_8453,N_8334,N_8327);
and U8454 (N_8454,N_8392,N_8301);
or U8455 (N_8455,N_8332,N_8328);
nor U8456 (N_8456,N_8320,N_8316);
nand U8457 (N_8457,N_8355,N_8320);
nor U8458 (N_8458,N_8339,N_8395);
or U8459 (N_8459,N_8311,N_8342);
nand U8460 (N_8460,N_8348,N_8309);
nand U8461 (N_8461,N_8381,N_8353);
and U8462 (N_8462,N_8364,N_8311);
nor U8463 (N_8463,N_8328,N_8303);
nand U8464 (N_8464,N_8367,N_8344);
or U8465 (N_8465,N_8319,N_8311);
nand U8466 (N_8466,N_8345,N_8344);
xor U8467 (N_8467,N_8362,N_8382);
xnor U8468 (N_8468,N_8390,N_8371);
nand U8469 (N_8469,N_8338,N_8390);
and U8470 (N_8470,N_8390,N_8352);
nor U8471 (N_8471,N_8371,N_8320);
xnor U8472 (N_8472,N_8358,N_8322);
and U8473 (N_8473,N_8318,N_8367);
xor U8474 (N_8474,N_8373,N_8389);
and U8475 (N_8475,N_8387,N_8377);
xor U8476 (N_8476,N_8393,N_8359);
and U8477 (N_8477,N_8384,N_8317);
xor U8478 (N_8478,N_8329,N_8333);
nand U8479 (N_8479,N_8345,N_8339);
xnor U8480 (N_8480,N_8342,N_8382);
and U8481 (N_8481,N_8334,N_8368);
nand U8482 (N_8482,N_8368,N_8364);
or U8483 (N_8483,N_8309,N_8389);
xor U8484 (N_8484,N_8340,N_8380);
nor U8485 (N_8485,N_8327,N_8331);
nor U8486 (N_8486,N_8367,N_8349);
xnor U8487 (N_8487,N_8348,N_8384);
nand U8488 (N_8488,N_8326,N_8310);
or U8489 (N_8489,N_8340,N_8398);
nor U8490 (N_8490,N_8336,N_8368);
or U8491 (N_8491,N_8328,N_8300);
xnor U8492 (N_8492,N_8347,N_8342);
or U8493 (N_8493,N_8314,N_8304);
nor U8494 (N_8494,N_8373,N_8301);
and U8495 (N_8495,N_8349,N_8385);
xnor U8496 (N_8496,N_8348,N_8308);
and U8497 (N_8497,N_8361,N_8369);
or U8498 (N_8498,N_8328,N_8383);
nand U8499 (N_8499,N_8335,N_8353);
xor U8500 (N_8500,N_8470,N_8458);
or U8501 (N_8501,N_8479,N_8437);
or U8502 (N_8502,N_8457,N_8469);
nor U8503 (N_8503,N_8438,N_8455);
or U8504 (N_8504,N_8495,N_8445);
nand U8505 (N_8505,N_8490,N_8420);
nand U8506 (N_8506,N_8484,N_8453);
nor U8507 (N_8507,N_8425,N_8407);
nor U8508 (N_8508,N_8492,N_8465);
or U8509 (N_8509,N_8491,N_8423);
or U8510 (N_8510,N_8478,N_8485);
nand U8511 (N_8511,N_8439,N_8463);
or U8512 (N_8512,N_8405,N_8427);
nand U8513 (N_8513,N_8499,N_8411);
nor U8514 (N_8514,N_8414,N_8400);
and U8515 (N_8515,N_8450,N_8417);
nor U8516 (N_8516,N_8422,N_8496);
xnor U8517 (N_8517,N_8472,N_8431);
or U8518 (N_8518,N_8424,N_8434);
nor U8519 (N_8519,N_8440,N_8403);
nor U8520 (N_8520,N_8482,N_8446);
nor U8521 (N_8521,N_8421,N_8471);
and U8522 (N_8522,N_8408,N_8473);
nor U8523 (N_8523,N_8435,N_8454);
or U8524 (N_8524,N_8404,N_8444);
xor U8525 (N_8525,N_8452,N_8430);
nand U8526 (N_8526,N_8409,N_8415);
xor U8527 (N_8527,N_8441,N_8461);
nor U8528 (N_8528,N_8456,N_8474);
nor U8529 (N_8529,N_8402,N_8416);
and U8530 (N_8530,N_8413,N_8447);
or U8531 (N_8531,N_8448,N_8493);
xor U8532 (N_8532,N_8487,N_8467);
or U8533 (N_8533,N_8483,N_8443);
nor U8534 (N_8534,N_8480,N_8426);
or U8535 (N_8535,N_8481,N_8462);
and U8536 (N_8536,N_8477,N_8433);
nand U8537 (N_8537,N_8464,N_8419);
nand U8538 (N_8538,N_8436,N_8418);
xnor U8539 (N_8539,N_8476,N_8475);
or U8540 (N_8540,N_8410,N_8459);
or U8541 (N_8541,N_8489,N_8428);
nand U8542 (N_8542,N_8498,N_8497);
and U8543 (N_8543,N_8451,N_8406);
or U8544 (N_8544,N_8486,N_8449);
xor U8545 (N_8545,N_8432,N_8429);
or U8546 (N_8546,N_8412,N_8442);
nand U8547 (N_8547,N_8488,N_8460);
nand U8548 (N_8548,N_8494,N_8466);
xor U8549 (N_8549,N_8468,N_8401);
nor U8550 (N_8550,N_8498,N_8436);
nor U8551 (N_8551,N_8431,N_8419);
or U8552 (N_8552,N_8436,N_8496);
and U8553 (N_8553,N_8441,N_8466);
and U8554 (N_8554,N_8491,N_8413);
and U8555 (N_8555,N_8459,N_8469);
xor U8556 (N_8556,N_8412,N_8430);
or U8557 (N_8557,N_8459,N_8439);
xor U8558 (N_8558,N_8403,N_8448);
nand U8559 (N_8559,N_8422,N_8474);
and U8560 (N_8560,N_8454,N_8478);
or U8561 (N_8561,N_8445,N_8464);
and U8562 (N_8562,N_8403,N_8422);
nor U8563 (N_8563,N_8436,N_8423);
or U8564 (N_8564,N_8411,N_8406);
and U8565 (N_8565,N_8426,N_8464);
xor U8566 (N_8566,N_8400,N_8487);
nand U8567 (N_8567,N_8444,N_8473);
or U8568 (N_8568,N_8493,N_8441);
or U8569 (N_8569,N_8405,N_8434);
nand U8570 (N_8570,N_8406,N_8407);
nor U8571 (N_8571,N_8468,N_8423);
nor U8572 (N_8572,N_8462,N_8479);
and U8573 (N_8573,N_8472,N_8465);
nand U8574 (N_8574,N_8419,N_8437);
and U8575 (N_8575,N_8429,N_8461);
nand U8576 (N_8576,N_8461,N_8445);
xor U8577 (N_8577,N_8454,N_8416);
nor U8578 (N_8578,N_8460,N_8430);
xnor U8579 (N_8579,N_8484,N_8437);
and U8580 (N_8580,N_8450,N_8407);
xor U8581 (N_8581,N_8443,N_8413);
nor U8582 (N_8582,N_8437,N_8436);
xor U8583 (N_8583,N_8475,N_8481);
or U8584 (N_8584,N_8406,N_8428);
and U8585 (N_8585,N_8430,N_8496);
or U8586 (N_8586,N_8480,N_8416);
and U8587 (N_8587,N_8436,N_8441);
nor U8588 (N_8588,N_8408,N_8451);
nand U8589 (N_8589,N_8432,N_8420);
xnor U8590 (N_8590,N_8432,N_8439);
xnor U8591 (N_8591,N_8420,N_8433);
and U8592 (N_8592,N_8441,N_8453);
or U8593 (N_8593,N_8499,N_8471);
nor U8594 (N_8594,N_8499,N_8403);
nand U8595 (N_8595,N_8475,N_8462);
xor U8596 (N_8596,N_8460,N_8492);
nor U8597 (N_8597,N_8407,N_8472);
xor U8598 (N_8598,N_8439,N_8412);
nand U8599 (N_8599,N_8492,N_8462);
nor U8600 (N_8600,N_8583,N_8587);
or U8601 (N_8601,N_8578,N_8564);
nor U8602 (N_8602,N_8540,N_8572);
xor U8603 (N_8603,N_8592,N_8531);
nand U8604 (N_8604,N_8551,N_8599);
nor U8605 (N_8605,N_8503,N_8508);
nand U8606 (N_8606,N_8566,N_8500);
or U8607 (N_8607,N_8553,N_8588);
xor U8608 (N_8608,N_8548,N_8597);
and U8609 (N_8609,N_8525,N_8567);
nor U8610 (N_8610,N_8533,N_8506);
and U8611 (N_8611,N_8546,N_8589);
and U8612 (N_8612,N_8552,N_8507);
or U8613 (N_8613,N_8520,N_8547);
and U8614 (N_8614,N_8509,N_8544);
and U8615 (N_8615,N_8542,N_8517);
or U8616 (N_8616,N_8574,N_8535);
or U8617 (N_8617,N_8561,N_8523);
or U8618 (N_8618,N_8591,N_8534);
and U8619 (N_8619,N_8569,N_8570);
nor U8620 (N_8620,N_8596,N_8585);
nand U8621 (N_8621,N_8521,N_8524);
nor U8622 (N_8622,N_8532,N_8558);
nand U8623 (N_8623,N_8590,N_8539);
nand U8624 (N_8624,N_8582,N_8526);
nand U8625 (N_8625,N_8527,N_8579);
and U8626 (N_8626,N_8573,N_8543);
or U8627 (N_8627,N_8537,N_8554);
nand U8628 (N_8628,N_8515,N_8584);
and U8629 (N_8629,N_8580,N_8536);
nor U8630 (N_8630,N_8576,N_8556);
and U8631 (N_8631,N_8593,N_8519);
nand U8632 (N_8632,N_8528,N_8516);
nor U8633 (N_8633,N_8560,N_8502);
nand U8634 (N_8634,N_8598,N_8549);
nor U8635 (N_8635,N_8504,N_8541);
nor U8636 (N_8636,N_8577,N_8568);
and U8637 (N_8637,N_8555,N_8512);
xnor U8638 (N_8638,N_8505,N_8550);
xnor U8639 (N_8639,N_8565,N_8594);
or U8640 (N_8640,N_8545,N_8514);
xnor U8641 (N_8641,N_8529,N_8557);
and U8642 (N_8642,N_8513,N_8595);
xnor U8643 (N_8643,N_8518,N_8522);
and U8644 (N_8644,N_8563,N_8501);
or U8645 (N_8645,N_8538,N_8571);
nor U8646 (N_8646,N_8586,N_8511);
xor U8647 (N_8647,N_8562,N_8559);
nor U8648 (N_8648,N_8575,N_8510);
xnor U8649 (N_8649,N_8581,N_8530);
and U8650 (N_8650,N_8553,N_8525);
xnor U8651 (N_8651,N_8589,N_8564);
and U8652 (N_8652,N_8521,N_8588);
or U8653 (N_8653,N_8530,N_8508);
nand U8654 (N_8654,N_8528,N_8559);
nor U8655 (N_8655,N_8595,N_8537);
nand U8656 (N_8656,N_8539,N_8537);
nand U8657 (N_8657,N_8514,N_8526);
xor U8658 (N_8658,N_8554,N_8583);
nor U8659 (N_8659,N_8524,N_8571);
and U8660 (N_8660,N_8550,N_8551);
and U8661 (N_8661,N_8540,N_8533);
nand U8662 (N_8662,N_8575,N_8568);
or U8663 (N_8663,N_8568,N_8522);
and U8664 (N_8664,N_8557,N_8515);
and U8665 (N_8665,N_8575,N_8549);
xor U8666 (N_8666,N_8543,N_8516);
or U8667 (N_8667,N_8539,N_8579);
or U8668 (N_8668,N_8532,N_8516);
and U8669 (N_8669,N_8585,N_8508);
xnor U8670 (N_8670,N_8527,N_8568);
xor U8671 (N_8671,N_8531,N_8565);
nor U8672 (N_8672,N_8544,N_8591);
or U8673 (N_8673,N_8562,N_8589);
nor U8674 (N_8674,N_8599,N_8508);
nand U8675 (N_8675,N_8595,N_8517);
nor U8676 (N_8676,N_8576,N_8551);
xnor U8677 (N_8677,N_8590,N_8529);
and U8678 (N_8678,N_8522,N_8546);
nand U8679 (N_8679,N_8561,N_8512);
nand U8680 (N_8680,N_8513,N_8544);
xnor U8681 (N_8681,N_8576,N_8501);
xor U8682 (N_8682,N_8586,N_8534);
and U8683 (N_8683,N_8562,N_8513);
xnor U8684 (N_8684,N_8510,N_8525);
and U8685 (N_8685,N_8582,N_8583);
and U8686 (N_8686,N_8514,N_8595);
nand U8687 (N_8687,N_8560,N_8535);
xnor U8688 (N_8688,N_8588,N_8548);
xor U8689 (N_8689,N_8583,N_8591);
xor U8690 (N_8690,N_8555,N_8573);
xnor U8691 (N_8691,N_8592,N_8586);
or U8692 (N_8692,N_8506,N_8596);
nor U8693 (N_8693,N_8560,N_8585);
nand U8694 (N_8694,N_8550,N_8569);
nor U8695 (N_8695,N_8591,N_8510);
xnor U8696 (N_8696,N_8503,N_8561);
nor U8697 (N_8697,N_8593,N_8543);
nor U8698 (N_8698,N_8567,N_8581);
nand U8699 (N_8699,N_8530,N_8503);
xor U8700 (N_8700,N_8626,N_8610);
or U8701 (N_8701,N_8678,N_8691);
or U8702 (N_8702,N_8631,N_8646);
nand U8703 (N_8703,N_8687,N_8621);
or U8704 (N_8704,N_8697,N_8683);
and U8705 (N_8705,N_8698,N_8616);
and U8706 (N_8706,N_8686,N_8649);
and U8707 (N_8707,N_8624,N_8604);
xnor U8708 (N_8708,N_8670,N_8679);
and U8709 (N_8709,N_8630,N_8607);
nor U8710 (N_8710,N_8611,N_8693);
nor U8711 (N_8711,N_8688,N_8656);
nand U8712 (N_8712,N_8644,N_8677);
nand U8713 (N_8713,N_8608,N_8619);
and U8714 (N_8714,N_8650,N_8613);
nand U8715 (N_8715,N_8675,N_8676);
nor U8716 (N_8716,N_8625,N_8640);
or U8717 (N_8717,N_8685,N_8667);
nor U8718 (N_8718,N_8643,N_8668);
nand U8719 (N_8719,N_8689,N_8618);
and U8720 (N_8720,N_8682,N_8692);
and U8721 (N_8721,N_8662,N_8681);
and U8722 (N_8722,N_8654,N_8633);
or U8723 (N_8723,N_8632,N_8699);
xnor U8724 (N_8724,N_8660,N_8659);
nand U8725 (N_8725,N_8620,N_8627);
xnor U8726 (N_8726,N_8638,N_8673);
xnor U8727 (N_8727,N_8680,N_8628);
xor U8728 (N_8728,N_8652,N_8622);
nand U8729 (N_8729,N_8690,N_8623);
or U8730 (N_8730,N_8661,N_8674);
and U8731 (N_8731,N_8696,N_8601);
nand U8732 (N_8732,N_8647,N_8669);
or U8733 (N_8733,N_8602,N_8664);
and U8734 (N_8734,N_8671,N_8603);
nand U8735 (N_8735,N_8606,N_8653);
nand U8736 (N_8736,N_8615,N_8695);
or U8737 (N_8737,N_8612,N_8642);
nand U8738 (N_8738,N_8617,N_8684);
and U8739 (N_8739,N_8629,N_8636);
nand U8740 (N_8740,N_8663,N_8655);
nand U8741 (N_8741,N_8658,N_8641);
xor U8742 (N_8742,N_8645,N_8635);
xnor U8743 (N_8743,N_8651,N_8637);
xor U8744 (N_8744,N_8600,N_8648);
and U8745 (N_8745,N_8639,N_8657);
xnor U8746 (N_8746,N_8666,N_8694);
and U8747 (N_8747,N_8605,N_8672);
xor U8748 (N_8748,N_8609,N_8614);
and U8749 (N_8749,N_8634,N_8665);
nor U8750 (N_8750,N_8644,N_8640);
nor U8751 (N_8751,N_8676,N_8620);
xnor U8752 (N_8752,N_8686,N_8603);
xor U8753 (N_8753,N_8676,N_8614);
xor U8754 (N_8754,N_8642,N_8683);
or U8755 (N_8755,N_8613,N_8653);
nor U8756 (N_8756,N_8622,N_8634);
nor U8757 (N_8757,N_8673,N_8652);
nor U8758 (N_8758,N_8667,N_8616);
nand U8759 (N_8759,N_8608,N_8650);
and U8760 (N_8760,N_8651,N_8682);
nor U8761 (N_8761,N_8694,N_8682);
and U8762 (N_8762,N_8645,N_8671);
nand U8763 (N_8763,N_8686,N_8604);
xor U8764 (N_8764,N_8641,N_8695);
nand U8765 (N_8765,N_8665,N_8659);
or U8766 (N_8766,N_8673,N_8640);
or U8767 (N_8767,N_8698,N_8646);
and U8768 (N_8768,N_8651,N_8644);
nand U8769 (N_8769,N_8638,N_8611);
or U8770 (N_8770,N_8619,N_8647);
nor U8771 (N_8771,N_8632,N_8611);
or U8772 (N_8772,N_8690,N_8643);
and U8773 (N_8773,N_8646,N_8678);
xnor U8774 (N_8774,N_8678,N_8653);
and U8775 (N_8775,N_8695,N_8670);
nand U8776 (N_8776,N_8658,N_8638);
nand U8777 (N_8777,N_8693,N_8625);
nor U8778 (N_8778,N_8679,N_8662);
nor U8779 (N_8779,N_8607,N_8639);
and U8780 (N_8780,N_8691,N_8675);
nand U8781 (N_8781,N_8642,N_8661);
nor U8782 (N_8782,N_8669,N_8690);
xnor U8783 (N_8783,N_8620,N_8619);
nor U8784 (N_8784,N_8628,N_8685);
xnor U8785 (N_8785,N_8644,N_8658);
nand U8786 (N_8786,N_8610,N_8644);
or U8787 (N_8787,N_8667,N_8648);
nand U8788 (N_8788,N_8654,N_8660);
nand U8789 (N_8789,N_8620,N_8665);
nand U8790 (N_8790,N_8620,N_8653);
or U8791 (N_8791,N_8665,N_8668);
or U8792 (N_8792,N_8646,N_8656);
xnor U8793 (N_8793,N_8631,N_8623);
nor U8794 (N_8794,N_8665,N_8636);
or U8795 (N_8795,N_8682,N_8629);
and U8796 (N_8796,N_8611,N_8627);
and U8797 (N_8797,N_8627,N_8633);
xor U8798 (N_8798,N_8642,N_8674);
or U8799 (N_8799,N_8655,N_8636);
nand U8800 (N_8800,N_8719,N_8784);
or U8801 (N_8801,N_8769,N_8767);
nand U8802 (N_8802,N_8773,N_8742);
xor U8803 (N_8803,N_8702,N_8739);
and U8804 (N_8804,N_8772,N_8718);
nand U8805 (N_8805,N_8722,N_8762);
and U8806 (N_8806,N_8793,N_8755);
nor U8807 (N_8807,N_8752,N_8789);
nand U8808 (N_8808,N_8779,N_8732);
or U8809 (N_8809,N_8709,N_8712);
nor U8810 (N_8810,N_8766,N_8735);
nor U8811 (N_8811,N_8795,N_8751);
nor U8812 (N_8812,N_8775,N_8798);
and U8813 (N_8813,N_8711,N_8743);
or U8814 (N_8814,N_8726,N_8791);
xnor U8815 (N_8815,N_8760,N_8745);
nor U8816 (N_8816,N_8746,N_8749);
xnor U8817 (N_8817,N_8776,N_8753);
or U8818 (N_8818,N_8721,N_8786);
xnor U8819 (N_8819,N_8778,N_8705);
nor U8820 (N_8820,N_8731,N_8780);
xor U8821 (N_8821,N_8733,N_8761);
nor U8822 (N_8822,N_8737,N_8736);
nor U8823 (N_8823,N_8750,N_8790);
and U8824 (N_8824,N_8715,N_8796);
or U8825 (N_8825,N_8707,N_8782);
xor U8826 (N_8826,N_8730,N_8748);
nand U8827 (N_8827,N_8774,N_8700);
xor U8828 (N_8828,N_8701,N_8787);
xor U8829 (N_8829,N_8708,N_8728);
and U8830 (N_8830,N_8765,N_8741);
nor U8831 (N_8831,N_8727,N_8714);
xnor U8832 (N_8832,N_8729,N_8781);
and U8833 (N_8833,N_8724,N_8754);
nor U8834 (N_8834,N_8785,N_8720);
and U8835 (N_8835,N_8740,N_8768);
nand U8836 (N_8836,N_8716,N_8757);
and U8837 (N_8837,N_8799,N_8771);
nor U8838 (N_8838,N_8717,N_8788);
nor U8839 (N_8839,N_8770,N_8783);
nor U8840 (N_8840,N_8764,N_8797);
xnor U8841 (N_8841,N_8704,N_8747);
and U8842 (N_8842,N_8792,N_8758);
or U8843 (N_8843,N_8777,N_8710);
xnor U8844 (N_8844,N_8794,N_8738);
and U8845 (N_8845,N_8703,N_8713);
and U8846 (N_8846,N_8759,N_8723);
or U8847 (N_8847,N_8734,N_8744);
nand U8848 (N_8848,N_8725,N_8706);
or U8849 (N_8849,N_8763,N_8756);
or U8850 (N_8850,N_8752,N_8746);
xnor U8851 (N_8851,N_8771,N_8735);
nand U8852 (N_8852,N_8777,N_8771);
or U8853 (N_8853,N_8764,N_8760);
nor U8854 (N_8854,N_8752,N_8718);
and U8855 (N_8855,N_8792,N_8761);
xor U8856 (N_8856,N_8781,N_8756);
xor U8857 (N_8857,N_8712,N_8708);
nor U8858 (N_8858,N_8777,N_8709);
xor U8859 (N_8859,N_8796,N_8752);
or U8860 (N_8860,N_8709,N_8787);
or U8861 (N_8861,N_8772,N_8798);
xnor U8862 (N_8862,N_8792,N_8744);
nand U8863 (N_8863,N_8712,N_8778);
nand U8864 (N_8864,N_8736,N_8735);
and U8865 (N_8865,N_8772,N_8766);
nor U8866 (N_8866,N_8785,N_8767);
or U8867 (N_8867,N_8752,N_8736);
nand U8868 (N_8868,N_8761,N_8734);
nor U8869 (N_8869,N_8784,N_8724);
xnor U8870 (N_8870,N_8785,N_8774);
or U8871 (N_8871,N_8714,N_8715);
xor U8872 (N_8872,N_8791,N_8767);
and U8873 (N_8873,N_8790,N_8747);
and U8874 (N_8874,N_8737,N_8759);
or U8875 (N_8875,N_8797,N_8740);
and U8876 (N_8876,N_8760,N_8743);
nor U8877 (N_8877,N_8702,N_8701);
or U8878 (N_8878,N_8722,N_8732);
nand U8879 (N_8879,N_8772,N_8738);
and U8880 (N_8880,N_8788,N_8731);
nor U8881 (N_8881,N_8726,N_8781);
nor U8882 (N_8882,N_8790,N_8720);
and U8883 (N_8883,N_8713,N_8726);
and U8884 (N_8884,N_8792,N_8782);
nand U8885 (N_8885,N_8718,N_8729);
nor U8886 (N_8886,N_8707,N_8711);
nor U8887 (N_8887,N_8741,N_8700);
or U8888 (N_8888,N_8721,N_8739);
or U8889 (N_8889,N_8738,N_8741);
nor U8890 (N_8890,N_8789,N_8796);
nand U8891 (N_8891,N_8707,N_8731);
nor U8892 (N_8892,N_8770,N_8756);
xor U8893 (N_8893,N_8713,N_8720);
and U8894 (N_8894,N_8714,N_8759);
nor U8895 (N_8895,N_8740,N_8718);
nor U8896 (N_8896,N_8763,N_8745);
xnor U8897 (N_8897,N_8799,N_8760);
or U8898 (N_8898,N_8765,N_8722);
nor U8899 (N_8899,N_8799,N_8798);
and U8900 (N_8900,N_8844,N_8807);
and U8901 (N_8901,N_8856,N_8897);
or U8902 (N_8902,N_8860,N_8865);
nand U8903 (N_8903,N_8810,N_8843);
nor U8904 (N_8904,N_8876,N_8861);
nor U8905 (N_8905,N_8830,N_8854);
and U8906 (N_8906,N_8874,N_8841);
and U8907 (N_8907,N_8840,N_8824);
nor U8908 (N_8908,N_8850,N_8836);
xor U8909 (N_8909,N_8883,N_8852);
nand U8910 (N_8910,N_8878,N_8834);
or U8911 (N_8911,N_8821,N_8838);
or U8912 (N_8912,N_8858,N_8822);
xnor U8913 (N_8913,N_8851,N_8812);
and U8914 (N_8914,N_8832,N_8847);
nand U8915 (N_8915,N_8866,N_8864);
xnor U8916 (N_8916,N_8862,N_8896);
or U8917 (N_8917,N_8881,N_8871);
nand U8918 (N_8918,N_8875,N_8857);
or U8919 (N_8919,N_8873,N_8828);
or U8920 (N_8920,N_8880,N_8898);
nor U8921 (N_8921,N_8815,N_8888);
and U8922 (N_8922,N_8820,N_8891);
or U8923 (N_8923,N_8823,N_8894);
or U8924 (N_8924,N_8887,N_8890);
or U8925 (N_8925,N_8831,N_8826);
and U8926 (N_8926,N_8893,N_8884);
nand U8927 (N_8927,N_8879,N_8877);
nand U8928 (N_8928,N_8829,N_8859);
nor U8929 (N_8929,N_8818,N_8804);
and U8930 (N_8930,N_8809,N_8867);
nand U8931 (N_8931,N_8846,N_8870);
xnor U8932 (N_8932,N_8817,N_8805);
or U8933 (N_8933,N_8801,N_8863);
and U8934 (N_8934,N_8839,N_8803);
or U8935 (N_8935,N_8816,N_8814);
or U8936 (N_8936,N_8837,N_8849);
xor U8937 (N_8937,N_8889,N_8892);
nand U8938 (N_8938,N_8885,N_8842);
or U8939 (N_8939,N_8848,N_8869);
and U8940 (N_8940,N_8845,N_8802);
or U8941 (N_8941,N_8813,N_8895);
and U8942 (N_8942,N_8899,N_8827);
or U8943 (N_8943,N_8835,N_8872);
xnor U8944 (N_8944,N_8819,N_8868);
nand U8945 (N_8945,N_8800,N_8808);
nor U8946 (N_8946,N_8811,N_8806);
or U8947 (N_8947,N_8853,N_8825);
xor U8948 (N_8948,N_8833,N_8855);
nor U8949 (N_8949,N_8886,N_8882);
or U8950 (N_8950,N_8800,N_8838);
or U8951 (N_8951,N_8848,N_8851);
or U8952 (N_8952,N_8846,N_8838);
xnor U8953 (N_8953,N_8883,N_8804);
and U8954 (N_8954,N_8831,N_8880);
nand U8955 (N_8955,N_8816,N_8855);
xor U8956 (N_8956,N_8837,N_8876);
and U8957 (N_8957,N_8847,N_8841);
nand U8958 (N_8958,N_8804,N_8888);
nor U8959 (N_8959,N_8819,N_8878);
and U8960 (N_8960,N_8867,N_8823);
xor U8961 (N_8961,N_8860,N_8897);
and U8962 (N_8962,N_8804,N_8872);
nand U8963 (N_8963,N_8820,N_8874);
and U8964 (N_8964,N_8883,N_8807);
xnor U8965 (N_8965,N_8844,N_8811);
xor U8966 (N_8966,N_8882,N_8843);
or U8967 (N_8967,N_8813,N_8871);
or U8968 (N_8968,N_8891,N_8804);
and U8969 (N_8969,N_8898,N_8863);
nor U8970 (N_8970,N_8819,N_8882);
or U8971 (N_8971,N_8879,N_8866);
nor U8972 (N_8972,N_8808,N_8802);
nand U8973 (N_8973,N_8803,N_8801);
and U8974 (N_8974,N_8874,N_8895);
nand U8975 (N_8975,N_8827,N_8872);
nand U8976 (N_8976,N_8855,N_8835);
nor U8977 (N_8977,N_8861,N_8807);
nor U8978 (N_8978,N_8850,N_8896);
nor U8979 (N_8979,N_8898,N_8830);
and U8980 (N_8980,N_8865,N_8809);
nand U8981 (N_8981,N_8881,N_8887);
xor U8982 (N_8982,N_8819,N_8881);
or U8983 (N_8983,N_8813,N_8845);
xnor U8984 (N_8984,N_8826,N_8879);
and U8985 (N_8985,N_8811,N_8863);
nand U8986 (N_8986,N_8843,N_8813);
and U8987 (N_8987,N_8874,N_8834);
or U8988 (N_8988,N_8834,N_8838);
nor U8989 (N_8989,N_8836,N_8826);
xnor U8990 (N_8990,N_8840,N_8858);
and U8991 (N_8991,N_8800,N_8883);
and U8992 (N_8992,N_8878,N_8861);
xnor U8993 (N_8993,N_8806,N_8814);
nor U8994 (N_8994,N_8840,N_8878);
nor U8995 (N_8995,N_8831,N_8894);
or U8996 (N_8996,N_8888,N_8882);
nor U8997 (N_8997,N_8825,N_8847);
nand U8998 (N_8998,N_8836,N_8867);
nand U8999 (N_8999,N_8879,N_8815);
or U9000 (N_9000,N_8902,N_8906);
and U9001 (N_9001,N_8914,N_8945);
or U9002 (N_9002,N_8940,N_8989);
nand U9003 (N_9003,N_8944,N_8987);
or U9004 (N_9004,N_8928,N_8970);
nor U9005 (N_9005,N_8979,N_8998);
nor U9006 (N_9006,N_8921,N_8964);
and U9007 (N_9007,N_8962,N_8963);
nor U9008 (N_9008,N_8984,N_8923);
nor U9009 (N_9009,N_8997,N_8992);
or U9010 (N_9010,N_8934,N_8935);
xor U9011 (N_9011,N_8937,N_8941);
nor U9012 (N_9012,N_8932,N_8960);
nor U9013 (N_9013,N_8975,N_8931);
nand U9014 (N_9014,N_8994,N_8965);
or U9015 (N_9015,N_8952,N_8949);
or U9016 (N_9016,N_8911,N_8917);
nand U9017 (N_9017,N_8948,N_8978);
xor U9018 (N_9018,N_8910,N_8972);
nand U9019 (N_9019,N_8985,N_8920);
xor U9020 (N_9020,N_8991,N_8986);
nor U9021 (N_9021,N_8909,N_8956);
or U9022 (N_9022,N_8976,N_8967);
nand U9023 (N_9023,N_8988,N_8900);
xnor U9024 (N_9024,N_8939,N_8959);
nand U9025 (N_9025,N_8971,N_8946);
and U9026 (N_9026,N_8990,N_8926);
nand U9027 (N_9027,N_8982,N_8968);
or U9028 (N_9028,N_8977,N_8999);
and U9029 (N_9029,N_8912,N_8916);
xor U9030 (N_9030,N_8966,N_8927);
and U9031 (N_9031,N_8915,N_8995);
xor U9032 (N_9032,N_8942,N_8980);
xor U9033 (N_9033,N_8969,N_8904);
or U9034 (N_9034,N_8922,N_8993);
or U9035 (N_9035,N_8981,N_8919);
nand U9036 (N_9036,N_8908,N_8955);
nand U9037 (N_9037,N_8947,N_8974);
xnor U9038 (N_9038,N_8961,N_8924);
and U9039 (N_9039,N_8958,N_8943);
or U9040 (N_9040,N_8907,N_8938);
nand U9041 (N_9041,N_8933,N_8954);
xnor U9042 (N_9042,N_8930,N_8905);
or U9043 (N_9043,N_8925,N_8996);
xnor U9044 (N_9044,N_8929,N_8973);
nand U9045 (N_9045,N_8983,N_8913);
nand U9046 (N_9046,N_8901,N_8957);
nand U9047 (N_9047,N_8918,N_8951);
nand U9048 (N_9048,N_8953,N_8936);
nor U9049 (N_9049,N_8950,N_8903);
nor U9050 (N_9050,N_8911,N_8934);
xnor U9051 (N_9051,N_8924,N_8973);
xor U9052 (N_9052,N_8917,N_8910);
nor U9053 (N_9053,N_8905,N_8925);
or U9054 (N_9054,N_8929,N_8982);
nand U9055 (N_9055,N_8944,N_8943);
nor U9056 (N_9056,N_8901,N_8904);
nor U9057 (N_9057,N_8934,N_8918);
nand U9058 (N_9058,N_8900,N_8928);
nand U9059 (N_9059,N_8902,N_8910);
nand U9060 (N_9060,N_8916,N_8997);
nand U9061 (N_9061,N_8913,N_8946);
xnor U9062 (N_9062,N_8965,N_8952);
xor U9063 (N_9063,N_8972,N_8915);
nor U9064 (N_9064,N_8924,N_8912);
or U9065 (N_9065,N_8970,N_8912);
and U9066 (N_9066,N_8943,N_8986);
xnor U9067 (N_9067,N_8928,N_8967);
or U9068 (N_9068,N_8998,N_8917);
and U9069 (N_9069,N_8929,N_8922);
nand U9070 (N_9070,N_8996,N_8919);
nor U9071 (N_9071,N_8983,N_8987);
and U9072 (N_9072,N_8960,N_8987);
nand U9073 (N_9073,N_8917,N_8947);
nor U9074 (N_9074,N_8942,N_8971);
xnor U9075 (N_9075,N_8996,N_8973);
or U9076 (N_9076,N_8939,N_8941);
nand U9077 (N_9077,N_8911,N_8962);
nor U9078 (N_9078,N_8985,N_8987);
or U9079 (N_9079,N_8922,N_8917);
nor U9080 (N_9080,N_8905,N_8932);
xnor U9081 (N_9081,N_8993,N_8905);
xor U9082 (N_9082,N_8994,N_8985);
and U9083 (N_9083,N_8947,N_8998);
and U9084 (N_9084,N_8963,N_8958);
nor U9085 (N_9085,N_8940,N_8991);
nand U9086 (N_9086,N_8928,N_8948);
and U9087 (N_9087,N_8936,N_8909);
or U9088 (N_9088,N_8916,N_8925);
and U9089 (N_9089,N_8962,N_8939);
xnor U9090 (N_9090,N_8987,N_8967);
or U9091 (N_9091,N_8933,N_8983);
nor U9092 (N_9092,N_8941,N_8912);
nor U9093 (N_9093,N_8940,N_8949);
nand U9094 (N_9094,N_8929,N_8986);
and U9095 (N_9095,N_8976,N_8929);
nor U9096 (N_9096,N_8920,N_8922);
nor U9097 (N_9097,N_8908,N_8983);
or U9098 (N_9098,N_8991,N_8907);
nor U9099 (N_9099,N_8913,N_8974);
and U9100 (N_9100,N_9032,N_9027);
nor U9101 (N_9101,N_9081,N_9039);
nand U9102 (N_9102,N_9086,N_9034);
xnor U9103 (N_9103,N_9042,N_9084);
nand U9104 (N_9104,N_9093,N_9014);
nand U9105 (N_9105,N_9026,N_9036);
nand U9106 (N_9106,N_9013,N_9012);
nor U9107 (N_9107,N_9030,N_9001);
nand U9108 (N_9108,N_9079,N_9009);
nand U9109 (N_9109,N_9041,N_9046);
nor U9110 (N_9110,N_9054,N_9015);
or U9111 (N_9111,N_9033,N_9095);
or U9112 (N_9112,N_9066,N_9067);
and U9113 (N_9113,N_9083,N_9068);
or U9114 (N_9114,N_9003,N_9055);
or U9115 (N_9115,N_9076,N_9016);
nor U9116 (N_9116,N_9060,N_9087);
xor U9117 (N_9117,N_9091,N_9048);
xnor U9118 (N_9118,N_9005,N_9062);
nor U9119 (N_9119,N_9065,N_9097);
xor U9120 (N_9120,N_9058,N_9080);
or U9121 (N_9121,N_9073,N_9052);
nand U9122 (N_9122,N_9098,N_9018);
or U9123 (N_9123,N_9035,N_9092);
or U9124 (N_9124,N_9011,N_9070);
or U9125 (N_9125,N_9008,N_9043);
nand U9126 (N_9126,N_9002,N_9006);
or U9127 (N_9127,N_9096,N_9063);
and U9128 (N_9128,N_9010,N_9044);
nor U9129 (N_9129,N_9029,N_9025);
nor U9130 (N_9130,N_9089,N_9047);
xor U9131 (N_9131,N_9099,N_9085);
or U9132 (N_9132,N_9007,N_9088);
nand U9133 (N_9133,N_9072,N_9064);
xnor U9134 (N_9134,N_9031,N_9051);
nor U9135 (N_9135,N_9069,N_9078);
nor U9136 (N_9136,N_9094,N_9040);
nand U9137 (N_9137,N_9074,N_9021);
xnor U9138 (N_9138,N_9038,N_9082);
nand U9139 (N_9139,N_9061,N_9000);
nor U9140 (N_9140,N_9024,N_9049);
xnor U9141 (N_9141,N_9023,N_9022);
nand U9142 (N_9142,N_9037,N_9004);
nor U9143 (N_9143,N_9056,N_9028);
nor U9144 (N_9144,N_9019,N_9077);
xnor U9145 (N_9145,N_9071,N_9050);
nand U9146 (N_9146,N_9075,N_9059);
nand U9147 (N_9147,N_9045,N_9017);
and U9148 (N_9148,N_9053,N_9090);
nor U9149 (N_9149,N_9057,N_9020);
nand U9150 (N_9150,N_9079,N_9078);
nor U9151 (N_9151,N_9092,N_9018);
nor U9152 (N_9152,N_9084,N_9095);
nand U9153 (N_9153,N_9079,N_9097);
nand U9154 (N_9154,N_9018,N_9027);
and U9155 (N_9155,N_9065,N_9087);
xor U9156 (N_9156,N_9051,N_9093);
or U9157 (N_9157,N_9039,N_9005);
and U9158 (N_9158,N_9017,N_9050);
nor U9159 (N_9159,N_9015,N_9081);
and U9160 (N_9160,N_9004,N_9074);
xnor U9161 (N_9161,N_9044,N_9022);
nor U9162 (N_9162,N_9090,N_9020);
nand U9163 (N_9163,N_9053,N_9083);
xor U9164 (N_9164,N_9008,N_9063);
or U9165 (N_9165,N_9041,N_9096);
nand U9166 (N_9166,N_9046,N_9013);
and U9167 (N_9167,N_9080,N_9091);
nand U9168 (N_9168,N_9045,N_9035);
nand U9169 (N_9169,N_9084,N_9032);
nor U9170 (N_9170,N_9079,N_9046);
nand U9171 (N_9171,N_9019,N_9032);
or U9172 (N_9172,N_9038,N_9051);
or U9173 (N_9173,N_9070,N_9078);
xor U9174 (N_9174,N_9037,N_9010);
xnor U9175 (N_9175,N_9060,N_9025);
or U9176 (N_9176,N_9041,N_9039);
and U9177 (N_9177,N_9077,N_9092);
or U9178 (N_9178,N_9051,N_9064);
nand U9179 (N_9179,N_9004,N_9088);
and U9180 (N_9180,N_9073,N_9009);
and U9181 (N_9181,N_9057,N_9028);
xor U9182 (N_9182,N_9006,N_9011);
xnor U9183 (N_9183,N_9076,N_9078);
or U9184 (N_9184,N_9085,N_9093);
xor U9185 (N_9185,N_9095,N_9097);
and U9186 (N_9186,N_9096,N_9067);
nand U9187 (N_9187,N_9077,N_9027);
xor U9188 (N_9188,N_9026,N_9030);
nand U9189 (N_9189,N_9002,N_9015);
or U9190 (N_9190,N_9006,N_9082);
and U9191 (N_9191,N_9094,N_9044);
nand U9192 (N_9192,N_9043,N_9031);
or U9193 (N_9193,N_9045,N_9097);
or U9194 (N_9194,N_9015,N_9093);
xor U9195 (N_9195,N_9048,N_9059);
nand U9196 (N_9196,N_9075,N_9055);
or U9197 (N_9197,N_9012,N_9002);
xor U9198 (N_9198,N_9096,N_9085);
nand U9199 (N_9199,N_9052,N_9021);
xnor U9200 (N_9200,N_9130,N_9161);
or U9201 (N_9201,N_9117,N_9120);
and U9202 (N_9202,N_9105,N_9153);
xnor U9203 (N_9203,N_9113,N_9115);
nor U9204 (N_9204,N_9134,N_9118);
nor U9205 (N_9205,N_9146,N_9114);
xor U9206 (N_9206,N_9108,N_9137);
and U9207 (N_9207,N_9181,N_9189);
xnor U9208 (N_9208,N_9185,N_9183);
and U9209 (N_9209,N_9122,N_9175);
and U9210 (N_9210,N_9159,N_9155);
or U9211 (N_9211,N_9164,N_9193);
xor U9212 (N_9212,N_9144,N_9194);
and U9213 (N_9213,N_9179,N_9199);
nor U9214 (N_9214,N_9192,N_9111);
nand U9215 (N_9215,N_9178,N_9167);
xor U9216 (N_9216,N_9186,N_9169);
nor U9217 (N_9217,N_9184,N_9107);
nor U9218 (N_9218,N_9132,N_9182);
nand U9219 (N_9219,N_9198,N_9124);
xor U9220 (N_9220,N_9150,N_9142);
or U9221 (N_9221,N_9116,N_9133);
xor U9222 (N_9222,N_9191,N_9187);
and U9223 (N_9223,N_9140,N_9176);
or U9224 (N_9224,N_9157,N_9103);
xor U9225 (N_9225,N_9196,N_9154);
nand U9226 (N_9226,N_9172,N_9145);
and U9227 (N_9227,N_9166,N_9141);
xnor U9228 (N_9228,N_9101,N_9123);
xnor U9229 (N_9229,N_9112,N_9136);
nor U9230 (N_9230,N_9156,N_9125);
and U9231 (N_9231,N_9168,N_9131);
or U9232 (N_9232,N_9121,N_9163);
nor U9233 (N_9233,N_9128,N_9148);
nand U9234 (N_9234,N_9143,N_9139);
xor U9235 (N_9235,N_9160,N_9152);
nor U9236 (N_9236,N_9180,N_9109);
and U9237 (N_9237,N_9162,N_9138);
xor U9238 (N_9238,N_9151,N_9158);
nand U9239 (N_9239,N_9102,N_9190);
nand U9240 (N_9240,N_9173,N_9106);
and U9241 (N_9241,N_9127,N_9135);
and U9242 (N_9242,N_9170,N_9110);
or U9243 (N_9243,N_9149,N_9197);
xor U9244 (N_9244,N_9171,N_9147);
and U9245 (N_9245,N_9126,N_9129);
nor U9246 (N_9246,N_9195,N_9177);
nand U9247 (N_9247,N_9100,N_9165);
xor U9248 (N_9248,N_9174,N_9104);
nor U9249 (N_9249,N_9188,N_9119);
xnor U9250 (N_9250,N_9185,N_9123);
or U9251 (N_9251,N_9199,N_9160);
xnor U9252 (N_9252,N_9184,N_9144);
or U9253 (N_9253,N_9130,N_9119);
xnor U9254 (N_9254,N_9133,N_9122);
nand U9255 (N_9255,N_9198,N_9166);
xor U9256 (N_9256,N_9199,N_9121);
or U9257 (N_9257,N_9134,N_9173);
nor U9258 (N_9258,N_9121,N_9189);
xnor U9259 (N_9259,N_9142,N_9190);
or U9260 (N_9260,N_9154,N_9184);
nor U9261 (N_9261,N_9179,N_9159);
and U9262 (N_9262,N_9114,N_9175);
or U9263 (N_9263,N_9167,N_9158);
and U9264 (N_9264,N_9139,N_9185);
or U9265 (N_9265,N_9128,N_9138);
and U9266 (N_9266,N_9188,N_9105);
or U9267 (N_9267,N_9124,N_9152);
and U9268 (N_9268,N_9100,N_9151);
and U9269 (N_9269,N_9126,N_9108);
or U9270 (N_9270,N_9166,N_9122);
or U9271 (N_9271,N_9161,N_9176);
xor U9272 (N_9272,N_9140,N_9177);
nor U9273 (N_9273,N_9140,N_9198);
or U9274 (N_9274,N_9136,N_9124);
xnor U9275 (N_9275,N_9136,N_9121);
nand U9276 (N_9276,N_9124,N_9158);
or U9277 (N_9277,N_9113,N_9187);
nor U9278 (N_9278,N_9183,N_9181);
xnor U9279 (N_9279,N_9135,N_9150);
xor U9280 (N_9280,N_9170,N_9131);
nor U9281 (N_9281,N_9100,N_9166);
or U9282 (N_9282,N_9173,N_9199);
nand U9283 (N_9283,N_9147,N_9194);
xor U9284 (N_9284,N_9146,N_9105);
xnor U9285 (N_9285,N_9100,N_9125);
nand U9286 (N_9286,N_9104,N_9181);
and U9287 (N_9287,N_9165,N_9173);
nand U9288 (N_9288,N_9122,N_9192);
nor U9289 (N_9289,N_9104,N_9125);
nand U9290 (N_9290,N_9100,N_9191);
nand U9291 (N_9291,N_9111,N_9143);
and U9292 (N_9292,N_9144,N_9102);
xnor U9293 (N_9293,N_9176,N_9195);
xnor U9294 (N_9294,N_9134,N_9160);
and U9295 (N_9295,N_9175,N_9111);
xnor U9296 (N_9296,N_9185,N_9199);
or U9297 (N_9297,N_9127,N_9185);
nor U9298 (N_9298,N_9170,N_9114);
xor U9299 (N_9299,N_9187,N_9183);
xor U9300 (N_9300,N_9287,N_9294);
nand U9301 (N_9301,N_9208,N_9283);
and U9302 (N_9302,N_9227,N_9219);
nand U9303 (N_9303,N_9286,N_9293);
and U9304 (N_9304,N_9223,N_9217);
nor U9305 (N_9305,N_9258,N_9226);
xor U9306 (N_9306,N_9210,N_9222);
and U9307 (N_9307,N_9279,N_9296);
and U9308 (N_9308,N_9228,N_9257);
or U9309 (N_9309,N_9242,N_9235);
xnor U9310 (N_9310,N_9206,N_9244);
and U9311 (N_9311,N_9285,N_9280);
xnor U9312 (N_9312,N_9209,N_9271);
or U9313 (N_9313,N_9238,N_9236);
and U9314 (N_9314,N_9270,N_9290);
nand U9315 (N_9315,N_9284,N_9274);
or U9316 (N_9316,N_9213,N_9201);
or U9317 (N_9317,N_9299,N_9266);
or U9318 (N_9318,N_9230,N_9218);
or U9319 (N_9319,N_9239,N_9237);
or U9320 (N_9320,N_9215,N_9297);
xnor U9321 (N_9321,N_9216,N_9224);
or U9322 (N_9322,N_9273,N_9241);
xor U9323 (N_9323,N_9259,N_9272);
xnor U9324 (N_9324,N_9214,N_9278);
nor U9325 (N_9325,N_9263,N_9276);
xnor U9326 (N_9326,N_9229,N_9289);
nor U9327 (N_9327,N_9200,N_9248);
xor U9328 (N_9328,N_9250,N_9205);
nand U9329 (N_9329,N_9234,N_9240);
nand U9330 (N_9330,N_9262,N_9243);
nor U9331 (N_9331,N_9249,N_9211);
nand U9332 (N_9332,N_9264,N_9277);
nor U9333 (N_9333,N_9232,N_9269);
nand U9334 (N_9334,N_9252,N_9261);
and U9335 (N_9335,N_9220,N_9202);
nand U9336 (N_9336,N_9275,N_9245);
nand U9337 (N_9337,N_9207,N_9288);
or U9338 (N_9338,N_9267,N_9225);
or U9339 (N_9339,N_9251,N_9253);
or U9340 (N_9340,N_9260,N_9281);
xnor U9341 (N_9341,N_9247,N_9292);
xnor U9342 (N_9342,N_9282,N_9203);
and U9343 (N_9343,N_9246,N_9233);
nor U9344 (N_9344,N_9256,N_9255);
nor U9345 (N_9345,N_9204,N_9265);
nor U9346 (N_9346,N_9254,N_9212);
or U9347 (N_9347,N_9221,N_9268);
xnor U9348 (N_9348,N_9295,N_9298);
nor U9349 (N_9349,N_9291,N_9231);
xor U9350 (N_9350,N_9256,N_9273);
nand U9351 (N_9351,N_9201,N_9237);
xnor U9352 (N_9352,N_9278,N_9297);
and U9353 (N_9353,N_9239,N_9293);
and U9354 (N_9354,N_9218,N_9272);
nand U9355 (N_9355,N_9213,N_9266);
nand U9356 (N_9356,N_9281,N_9267);
nand U9357 (N_9357,N_9228,N_9224);
nand U9358 (N_9358,N_9282,N_9238);
xnor U9359 (N_9359,N_9236,N_9218);
or U9360 (N_9360,N_9289,N_9211);
or U9361 (N_9361,N_9235,N_9252);
nand U9362 (N_9362,N_9213,N_9284);
xor U9363 (N_9363,N_9207,N_9263);
nand U9364 (N_9364,N_9211,N_9221);
and U9365 (N_9365,N_9204,N_9259);
and U9366 (N_9366,N_9229,N_9201);
nor U9367 (N_9367,N_9247,N_9286);
xnor U9368 (N_9368,N_9296,N_9267);
xnor U9369 (N_9369,N_9242,N_9210);
and U9370 (N_9370,N_9208,N_9220);
or U9371 (N_9371,N_9241,N_9251);
nand U9372 (N_9372,N_9285,N_9274);
nand U9373 (N_9373,N_9288,N_9273);
or U9374 (N_9374,N_9273,N_9201);
or U9375 (N_9375,N_9211,N_9234);
and U9376 (N_9376,N_9220,N_9292);
nand U9377 (N_9377,N_9252,N_9244);
xnor U9378 (N_9378,N_9246,N_9235);
nand U9379 (N_9379,N_9270,N_9260);
xnor U9380 (N_9380,N_9211,N_9246);
nor U9381 (N_9381,N_9266,N_9209);
xnor U9382 (N_9382,N_9296,N_9264);
and U9383 (N_9383,N_9219,N_9225);
and U9384 (N_9384,N_9263,N_9225);
and U9385 (N_9385,N_9291,N_9263);
nand U9386 (N_9386,N_9204,N_9225);
nor U9387 (N_9387,N_9281,N_9297);
nor U9388 (N_9388,N_9218,N_9223);
xnor U9389 (N_9389,N_9261,N_9234);
or U9390 (N_9390,N_9295,N_9272);
or U9391 (N_9391,N_9203,N_9234);
xor U9392 (N_9392,N_9242,N_9200);
or U9393 (N_9393,N_9284,N_9261);
or U9394 (N_9394,N_9249,N_9257);
or U9395 (N_9395,N_9217,N_9203);
and U9396 (N_9396,N_9254,N_9289);
or U9397 (N_9397,N_9210,N_9216);
nor U9398 (N_9398,N_9256,N_9286);
xnor U9399 (N_9399,N_9217,N_9225);
xor U9400 (N_9400,N_9341,N_9380);
and U9401 (N_9401,N_9363,N_9320);
or U9402 (N_9402,N_9331,N_9399);
and U9403 (N_9403,N_9311,N_9338);
or U9404 (N_9404,N_9378,N_9394);
and U9405 (N_9405,N_9340,N_9374);
nand U9406 (N_9406,N_9334,N_9355);
nand U9407 (N_9407,N_9318,N_9351);
nor U9408 (N_9408,N_9335,N_9322);
xor U9409 (N_9409,N_9303,N_9346);
or U9410 (N_9410,N_9316,N_9314);
or U9411 (N_9411,N_9313,N_9317);
nand U9412 (N_9412,N_9389,N_9309);
or U9413 (N_9413,N_9386,N_9326);
xnor U9414 (N_9414,N_9353,N_9366);
or U9415 (N_9415,N_9332,N_9306);
nor U9416 (N_9416,N_9310,N_9336);
nand U9417 (N_9417,N_9301,N_9312);
nor U9418 (N_9418,N_9364,N_9398);
nand U9419 (N_9419,N_9377,N_9349);
xnor U9420 (N_9420,N_9381,N_9369);
and U9421 (N_9421,N_9354,N_9391);
nor U9422 (N_9422,N_9368,N_9375);
xor U9423 (N_9423,N_9356,N_9384);
nor U9424 (N_9424,N_9344,N_9304);
and U9425 (N_9425,N_9327,N_9387);
nor U9426 (N_9426,N_9324,N_9370);
xnor U9427 (N_9427,N_9373,N_9342);
xnor U9428 (N_9428,N_9307,N_9395);
and U9429 (N_9429,N_9350,N_9323);
or U9430 (N_9430,N_9397,N_9371);
xor U9431 (N_9431,N_9308,N_9359);
and U9432 (N_9432,N_9319,N_9367);
nor U9433 (N_9433,N_9361,N_9352);
nand U9434 (N_9434,N_9328,N_9393);
xor U9435 (N_9435,N_9305,N_9372);
xnor U9436 (N_9436,N_9343,N_9321);
nand U9437 (N_9437,N_9339,N_9329);
nor U9438 (N_9438,N_9337,N_9302);
nand U9439 (N_9439,N_9392,N_9357);
and U9440 (N_9440,N_9347,N_9396);
and U9441 (N_9441,N_9300,N_9348);
xor U9442 (N_9442,N_9385,N_9325);
or U9443 (N_9443,N_9358,N_9345);
and U9444 (N_9444,N_9360,N_9365);
nor U9445 (N_9445,N_9376,N_9379);
or U9446 (N_9446,N_9390,N_9382);
or U9447 (N_9447,N_9333,N_9388);
or U9448 (N_9448,N_9330,N_9362);
nor U9449 (N_9449,N_9315,N_9383);
or U9450 (N_9450,N_9325,N_9316);
and U9451 (N_9451,N_9368,N_9328);
nor U9452 (N_9452,N_9353,N_9376);
xnor U9453 (N_9453,N_9308,N_9334);
nand U9454 (N_9454,N_9364,N_9341);
and U9455 (N_9455,N_9347,N_9331);
xnor U9456 (N_9456,N_9335,N_9359);
xnor U9457 (N_9457,N_9380,N_9328);
or U9458 (N_9458,N_9323,N_9326);
nand U9459 (N_9459,N_9318,N_9339);
or U9460 (N_9460,N_9328,N_9390);
nor U9461 (N_9461,N_9337,N_9381);
nand U9462 (N_9462,N_9305,N_9327);
and U9463 (N_9463,N_9326,N_9311);
nor U9464 (N_9464,N_9387,N_9380);
nand U9465 (N_9465,N_9333,N_9340);
or U9466 (N_9466,N_9353,N_9320);
or U9467 (N_9467,N_9309,N_9359);
nor U9468 (N_9468,N_9320,N_9308);
xnor U9469 (N_9469,N_9311,N_9310);
and U9470 (N_9470,N_9358,N_9391);
or U9471 (N_9471,N_9359,N_9386);
or U9472 (N_9472,N_9371,N_9358);
or U9473 (N_9473,N_9315,N_9316);
nor U9474 (N_9474,N_9328,N_9316);
and U9475 (N_9475,N_9386,N_9362);
nor U9476 (N_9476,N_9345,N_9352);
or U9477 (N_9477,N_9345,N_9309);
and U9478 (N_9478,N_9358,N_9396);
nor U9479 (N_9479,N_9387,N_9358);
and U9480 (N_9480,N_9357,N_9340);
or U9481 (N_9481,N_9364,N_9387);
or U9482 (N_9482,N_9320,N_9356);
and U9483 (N_9483,N_9378,N_9306);
nand U9484 (N_9484,N_9371,N_9332);
nor U9485 (N_9485,N_9321,N_9381);
or U9486 (N_9486,N_9349,N_9375);
or U9487 (N_9487,N_9301,N_9346);
nand U9488 (N_9488,N_9308,N_9301);
xnor U9489 (N_9489,N_9335,N_9314);
nor U9490 (N_9490,N_9348,N_9319);
or U9491 (N_9491,N_9333,N_9359);
nand U9492 (N_9492,N_9389,N_9366);
nand U9493 (N_9493,N_9338,N_9348);
nor U9494 (N_9494,N_9359,N_9391);
or U9495 (N_9495,N_9391,N_9344);
and U9496 (N_9496,N_9324,N_9354);
or U9497 (N_9497,N_9307,N_9325);
nand U9498 (N_9498,N_9348,N_9317);
and U9499 (N_9499,N_9359,N_9390);
or U9500 (N_9500,N_9446,N_9416);
nand U9501 (N_9501,N_9415,N_9494);
and U9502 (N_9502,N_9432,N_9441);
and U9503 (N_9503,N_9461,N_9485);
and U9504 (N_9504,N_9451,N_9498);
nand U9505 (N_9505,N_9422,N_9457);
nand U9506 (N_9506,N_9420,N_9476);
and U9507 (N_9507,N_9411,N_9433);
or U9508 (N_9508,N_9481,N_9499);
or U9509 (N_9509,N_9427,N_9444);
or U9510 (N_9510,N_9408,N_9463);
or U9511 (N_9511,N_9480,N_9426);
nor U9512 (N_9512,N_9442,N_9484);
nand U9513 (N_9513,N_9495,N_9448);
xor U9514 (N_9514,N_9456,N_9472);
or U9515 (N_9515,N_9445,N_9403);
nand U9516 (N_9516,N_9400,N_9402);
and U9517 (N_9517,N_9405,N_9412);
nand U9518 (N_9518,N_9497,N_9401);
xor U9519 (N_9519,N_9443,N_9493);
and U9520 (N_9520,N_9459,N_9449);
nand U9521 (N_9521,N_9429,N_9475);
nand U9522 (N_9522,N_9490,N_9409);
and U9523 (N_9523,N_9487,N_9423);
xor U9524 (N_9524,N_9468,N_9425);
and U9525 (N_9525,N_9462,N_9413);
xor U9526 (N_9526,N_9478,N_9473);
nor U9527 (N_9527,N_9486,N_9479);
nand U9528 (N_9528,N_9466,N_9440);
xor U9529 (N_9529,N_9491,N_9410);
and U9530 (N_9530,N_9471,N_9483);
nor U9531 (N_9531,N_9450,N_9469);
xnor U9532 (N_9532,N_9465,N_9467);
and U9533 (N_9533,N_9439,N_9430);
and U9534 (N_9534,N_9488,N_9435);
or U9535 (N_9535,N_9431,N_9474);
nand U9536 (N_9536,N_9424,N_9452);
or U9537 (N_9537,N_9464,N_9458);
nor U9538 (N_9538,N_9417,N_9455);
xnor U9539 (N_9539,N_9414,N_9470);
xor U9540 (N_9540,N_9437,N_9438);
and U9541 (N_9541,N_9434,N_9428);
or U9542 (N_9542,N_9421,N_9460);
or U9543 (N_9543,N_9404,N_9447);
nand U9544 (N_9544,N_9418,N_9492);
nor U9545 (N_9545,N_9406,N_9436);
xor U9546 (N_9546,N_9482,N_9419);
nand U9547 (N_9547,N_9496,N_9489);
or U9548 (N_9548,N_9453,N_9407);
and U9549 (N_9549,N_9454,N_9477);
nand U9550 (N_9550,N_9406,N_9403);
xor U9551 (N_9551,N_9442,N_9477);
nand U9552 (N_9552,N_9440,N_9476);
or U9553 (N_9553,N_9455,N_9467);
nor U9554 (N_9554,N_9455,N_9488);
xor U9555 (N_9555,N_9438,N_9493);
or U9556 (N_9556,N_9433,N_9488);
nor U9557 (N_9557,N_9468,N_9438);
or U9558 (N_9558,N_9426,N_9427);
xor U9559 (N_9559,N_9433,N_9401);
or U9560 (N_9560,N_9480,N_9467);
nand U9561 (N_9561,N_9465,N_9464);
or U9562 (N_9562,N_9422,N_9467);
or U9563 (N_9563,N_9466,N_9433);
or U9564 (N_9564,N_9486,N_9466);
and U9565 (N_9565,N_9416,N_9433);
nor U9566 (N_9566,N_9486,N_9400);
nand U9567 (N_9567,N_9433,N_9415);
and U9568 (N_9568,N_9473,N_9474);
nor U9569 (N_9569,N_9425,N_9493);
xor U9570 (N_9570,N_9464,N_9494);
nor U9571 (N_9571,N_9434,N_9445);
nor U9572 (N_9572,N_9425,N_9482);
and U9573 (N_9573,N_9410,N_9451);
or U9574 (N_9574,N_9444,N_9414);
and U9575 (N_9575,N_9487,N_9494);
nor U9576 (N_9576,N_9463,N_9431);
and U9577 (N_9577,N_9497,N_9416);
nor U9578 (N_9578,N_9451,N_9494);
nand U9579 (N_9579,N_9428,N_9468);
or U9580 (N_9580,N_9406,N_9472);
nor U9581 (N_9581,N_9496,N_9403);
or U9582 (N_9582,N_9442,N_9444);
nand U9583 (N_9583,N_9459,N_9443);
and U9584 (N_9584,N_9422,N_9483);
and U9585 (N_9585,N_9465,N_9494);
nand U9586 (N_9586,N_9487,N_9484);
and U9587 (N_9587,N_9486,N_9480);
nor U9588 (N_9588,N_9479,N_9492);
or U9589 (N_9589,N_9497,N_9409);
xor U9590 (N_9590,N_9449,N_9440);
xor U9591 (N_9591,N_9441,N_9499);
or U9592 (N_9592,N_9420,N_9460);
or U9593 (N_9593,N_9469,N_9466);
nor U9594 (N_9594,N_9418,N_9408);
nor U9595 (N_9595,N_9473,N_9442);
nand U9596 (N_9596,N_9422,N_9469);
and U9597 (N_9597,N_9459,N_9480);
or U9598 (N_9598,N_9485,N_9482);
nand U9599 (N_9599,N_9419,N_9466);
and U9600 (N_9600,N_9511,N_9598);
and U9601 (N_9601,N_9514,N_9556);
nand U9602 (N_9602,N_9545,N_9515);
or U9603 (N_9603,N_9535,N_9531);
nor U9604 (N_9604,N_9576,N_9574);
nor U9605 (N_9605,N_9591,N_9552);
and U9606 (N_9606,N_9590,N_9549);
nor U9607 (N_9607,N_9569,N_9560);
nand U9608 (N_9608,N_9584,N_9520);
nand U9609 (N_9609,N_9586,N_9540);
nand U9610 (N_9610,N_9543,N_9581);
xnor U9611 (N_9611,N_9597,N_9506);
nand U9612 (N_9612,N_9594,N_9582);
nand U9613 (N_9613,N_9538,N_9551);
nor U9614 (N_9614,N_9573,N_9599);
or U9615 (N_9615,N_9527,N_9561);
nor U9616 (N_9616,N_9503,N_9575);
nand U9617 (N_9617,N_9588,N_9505);
nor U9618 (N_9618,N_9517,N_9518);
xnor U9619 (N_9619,N_9593,N_9596);
xor U9620 (N_9620,N_9583,N_9544);
and U9621 (N_9621,N_9570,N_9567);
or U9622 (N_9622,N_9562,N_9523);
nand U9623 (N_9623,N_9534,N_9507);
xor U9624 (N_9624,N_9530,N_9592);
nor U9625 (N_9625,N_9513,N_9502);
nor U9626 (N_9626,N_9566,N_9529);
nand U9627 (N_9627,N_9572,N_9537);
nand U9628 (N_9628,N_9522,N_9536);
and U9629 (N_9629,N_9557,N_9516);
nand U9630 (N_9630,N_9528,N_9564);
or U9631 (N_9631,N_9547,N_9546);
nor U9632 (N_9632,N_9555,N_9554);
or U9633 (N_9633,N_9521,N_9504);
xnor U9634 (N_9634,N_9559,N_9595);
nand U9635 (N_9635,N_9577,N_9525);
nand U9636 (N_9636,N_9508,N_9541);
nand U9637 (N_9637,N_9579,N_9533);
nand U9638 (N_9638,N_9532,N_9542);
nor U9639 (N_9639,N_9500,N_9558);
nor U9640 (N_9640,N_9539,N_9578);
nand U9641 (N_9641,N_9565,N_9519);
nor U9642 (N_9642,N_9509,N_9512);
nand U9643 (N_9643,N_9553,N_9580);
nand U9644 (N_9644,N_9571,N_9526);
nor U9645 (N_9645,N_9501,N_9510);
nand U9646 (N_9646,N_9563,N_9589);
xnor U9647 (N_9647,N_9587,N_9568);
xnor U9648 (N_9648,N_9524,N_9585);
nand U9649 (N_9649,N_9550,N_9548);
or U9650 (N_9650,N_9587,N_9522);
and U9651 (N_9651,N_9541,N_9561);
or U9652 (N_9652,N_9578,N_9528);
and U9653 (N_9653,N_9590,N_9542);
xor U9654 (N_9654,N_9593,N_9531);
xor U9655 (N_9655,N_9530,N_9581);
or U9656 (N_9656,N_9554,N_9553);
nor U9657 (N_9657,N_9587,N_9569);
or U9658 (N_9658,N_9564,N_9540);
and U9659 (N_9659,N_9586,N_9560);
xor U9660 (N_9660,N_9574,N_9523);
nand U9661 (N_9661,N_9537,N_9536);
xor U9662 (N_9662,N_9532,N_9531);
or U9663 (N_9663,N_9529,N_9547);
or U9664 (N_9664,N_9518,N_9509);
xor U9665 (N_9665,N_9522,N_9566);
nor U9666 (N_9666,N_9559,N_9508);
and U9667 (N_9667,N_9517,N_9529);
or U9668 (N_9668,N_9561,N_9504);
or U9669 (N_9669,N_9586,N_9563);
and U9670 (N_9670,N_9563,N_9537);
nand U9671 (N_9671,N_9574,N_9548);
xnor U9672 (N_9672,N_9558,N_9573);
nand U9673 (N_9673,N_9593,N_9517);
nor U9674 (N_9674,N_9530,N_9550);
nand U9675 (N_9675,N_9592,N_9557);
nand U9676 (N_9676,N_9536,N_9581);
xor U9677 (N_9677,N_9555,N_9589);
nor U9678 (N_9678,N_9528,N_9512);
xor U9679 (N_9679,N_9593,N_9584);
xor U9680 (N_9680,N_9588,N_9529);
xnor U9681 (N_9681,N_9579,N_9582);
or U9682 (N_9682,N_9576,N_9585);
nor U9683 (N_9683,N_9526,N_9530);
and U9684 (N_9684,N_9580,N_9568);
and U9685 (N_9685,N_9541,N_9516);
and U9686 (N_9686,N_9597,N_9564);
xor U9687 (N_9687,N_9597,N_9517);
and U9688 (N_9688,N_9570,N_9513);
nor U9689 (N_9689,N_9537,N_9567);
and U9690 (N_9690,N_9576,N_9533);
nor U9691 (N_9691,N_9570,N_9510);
xor U9692 (N_9692,N_9559,N_9515);
or U9693 (N_9693,N_9518,N_9523);
nand U9694 (N_9694,N_9543,N_9542);
or U9695 (N_9695,N_9577,N_9597);
or U9696 (N_9696,N_9574,N_9571);
nand U9697 (N_9697,N_9590,N_9551);
xnor U9698 (N_9698,N_9501,N_9599);
xnor U9699 (N_9699,N_9564,N_9582);
or U9700 (N_9700,N_9603,N_9665);
nand U9701 (N_9701,N_9680,N_9663);
nand U9702 (N_9702,N_9619,N_9695);
xor U9703 (N_9703,N_9601,N_9678);
nor U9704 (N_9704,N_9651,N_9644);
nor U9705 (N_9705,N_9650,N_9681);
xor U9706 (N_9706,N_9643,N_9669);
nor U9707 (N_9707,N_9685,N_9639);
and U9708 (N_9708,N_9667,N_9628);
and U9709 (N_9709,N_9602,N_9674);
nor U9710 (N_9710,N_9609,N_9687);
nand U9711 (N_9711,N_9615,N_9621);
nand U9712 (N_9712,N_9620,N_9618);
nand U9713 (N_9713,N_9691,N_9630);
or U9714 (N_9714,N_9653,N_9629);
xor U9715 (N_9715,N_9637,N_9677);
nor U9716 (N_9716,N_9623,N_9657);
or U9717 (N_9717,N_9627,N_9694);
and U9718 (N_9718,N_9633,N_9625);
and U9719 (N_9719,N_9655,N_9668);
nor U9720 (N_9720,N_9689,N_9690);
nor U9721 (N_9721,N_9696,N_9675);
nor U9722 (N_9722,N_9626,N_9612);
and U9723 (N_9723,N_9610,N_9671);
nand U9724 (N_9724,N_9616,N_9632);
or U9725 (N_9725,N_9613,N_9676);
nor U9726 (N_9726,N_9614,N_9638);
or U9727 (N_9727,N_9649,N_9611);
xnor U9728 (N_9728,N_9617,N_9604);
or U9729 (N_9729,N_9608,N_9606);
nand U9730 (N_9730,N_9660,N_9673);
xor U9731 (N_9731,N_9645,N_9679);
nand U9732 (N_9732,N_9658,N_9693);
nand U9733 (N_9733,N_9662,N_9670);
xnor U9734 (N_9734,N_9664,N_9631);
nor U9735 (N_9735,N_9688,N_9642);
nand U9736 (N_9736,N_9607,N_9647);
or U9737 (N_9737,N_9624,N_9659);
xnor U9738 (N_9738,N_9635,N_9648);
nor U9739 (N_9739,N_9683,N_9661);
nand U9740 (N_9740,N_9672,N_9646);
nor U9741 (N_9741,N_9641,N_9600);
and U9742 (N_9742,N_9605,N_9636);
nor U9743 (N_9743,N_9698,N_9684);
xor U9744 (N_9744,N_9686,N_9640);
nor U9745 (N_9745,N_9654,N_9699);
nor U9746 (N_9746,N_9682,N_9697);
nand U9747 (N_9747,N_9634,N_9656);
xor U9748 (N_9748,N_9692,N_9666);
and U9749 (N_9749,N_9652,N_9622);
or U9750 (N_9750,N_9611,N_9664);
nand U9751 (N_9751,N_9634,N_9659);
nand U9752 (N_9752,N_9696,N_9656);
nand U9753 (N_9753,N_9626,N_9664);
or U9754 (N_9754,N_9629,N_9669);
nand U9755 (N_9755,N_9613,N_9660);
nand U9756 (N_9756,N_9656,N_9681);
nor U9757 (N_9757,N_9690,N_9673);
and U9758 (N_9758,N_9646,N_9615);
nand U9759 (N_9759,N_9687,N_9675);
nand U9760 (N_9760,N_9608,N_9676);
xor U9761 (N_9761,N_9644,N_9602);
or U9762 (N_9762,N_9674,N_9617);
xor U9763 (N_9763,N_9673,N_9677);
and U9764 (N_9764,N_9668,N_9609);
or U9765 (N_9765,N_9636,N_9644);
xnor U9766 (N_9766,N_9668,N_9678);
nor U9767 (N_9767,N_9620,N_9689);
or U9768 (N_9768,N_9659,N_9685);
nand U9769 (N_9769,N_9627,N_9629);
or U9770 (N_9770,N_9693,N_9673);
or U9771 (N_9771,N_9694,N_9602);
nor U9772 (N_9772,N_9640,N_9656);
and U9773 (N_9773,N_9614,N_9670);
or U9774 (N_9774,N_9678,N_9624);
or U9775 (N_9775,N_9676,N_9645);
and U9776 (N_9776,N_9625,N_9667);
xnor U9777 (N_9777,N_9691,N_9699);
xor U9778 (N_9778,N_9654,N_9614);
nor U9779 (N_9779,N_9680,N_9657);
or U9780 (N_9780,N_9669,N_9633);
nor U9781 (N_9781,N_9623,N_9677);
and U9782 (N_9782,N_9664,N_9624);
nand U9783 (N_9783,N_9668,N_9667);
nand U9784 (N_9784,N_9614,N_9659);
xor U9785 (N_9785,N_9638,N_9689);
and U9786 (N_9786,N_9646,N_9653);
or U9787 (N_9787,N_9612,N_9699);
nand U9788 (N_9788,N_9633,N_9639);
nand U9789 (N_9789,N_9679,N_9647);
or U9790 (N_9790,N_9685,N_9627);
or U9791 (N_9791,N_9668,N_9674);
xnor U9792 (N_9792,N_9634,N_9654);
and U9793 (N_9793,N_9609,N_9662);
nand U9794 (N_9794,N_9675,N_9604);
nand U9795 (N_9795,N_9652,N_9655);
and U9796 (N_9796,N_9616,N_9695);
nor U9797 (N_9797,N_9605,N_9650);
nand U9798 (N_9798,N_9669,N_9690);
or U9799 (N_9799,N_9627,N_9677);
xor U9800 (N_9800,N_9788,N_9752);
nand U9801 (N_9801,N_9711,N_9773);
and U9802 (N_9802,N_9745,N_9768);
nand U9803 (N_9803,N_9775,N_9780);
and U9804 (N_9804,N_9767,N_9721);
nor U9805 (N_9805,N_9785,N_9795);
and U9806 (N_9806,N_9717,N_9730);
nand U9807 (N_9807,N_9772,N_9759);
or U9808 (N_9808,N_9797,N_9705);
xor U9809 (N_9809,N_9700,N_9729);
and U9810 (N_9810,N_9708,N_9762);
nand U9811 (N_9811,N_9741,N_9727);
nor U9812 (N_9812,N_9756,N_9726);
and U9813 (N_9813,N_9779,N_9789);
nor U9814 (N_9814,N_9751,N_9704);
nor U9815 (N_9815,N_9723,N_9706);
nand U9816 (N_9816,N_9743,N_9781);
and U9817 (N_9817,N_9766,N_9747);
nor U9818 (N_9818,N_9764,N_9718);
nand U9819 (N_9819,N_9784,N_9794);
or U9820 (N_9820,N_9739,N_9733);
or U9821 (N_9821,N_9707,N_9750);
nand U9822 (N_9822,N_9791,N_9736);
nand U9823 (N_9823,N_9755,N_9731);
or U9824 (N_9824,N_9715,N_9719);
xor U9825 (N_9825,N_9738,N_9734);
and U9826 (N_9826,N_9761,N_9703);
nand U9827 (N_9827,N_9798,N_9782);
nor U9828 (N_9828,N_9744,N_9735);
nand U9829 (N_9829,N_9793,N_9713);
nor U9830 (N_9830,N_9760,N_9799);
nor U9831 (N_9831,N_9758,N_9728);
xor U9832 (N_9832,N_9740,N_9746);
or U9833 (N_9833,N_9774,N_9712);
and U9834 (N_9834,N_9757,N_9777);
nand U9835 (N_9835,N_9754,N_9722);
nand U9836 (N_9836,N_9783,N_9786);
nand U9837 (N_9837,N_9778,N_9714);
nand U9838 (N_9838,N_9710,N_9753);
and U9839 (N_9839,N_9724,N_9701);
nor U9840 (N_9840,N_9787,N_9709);
nand U9841 (N_9841,N_9771,N_9702);
xnor U9842 (N_9842,N_9716,N_9790);
xnor U9843 (N_9843,N_9765,N_9749);
nand U9844 (N_9844,N_9742,N_9732);
xnor U9845 (N_9845,N_9776,N_9737);
and U9846 (N_9846,N_9792,N_9763);
nor U9847 (N_9847,N_9748,N_9769);
xnor U9848 (N_9848,N_9770,N_9720);
or U9849 (N_9849,N_9796,N_9725);
nor U9850 (N_9850,N_9741,N_9784);
nand U9851 (N_9851,N_9785,N_9758);
nor U9852 (N_9852,N_9786,N_9722);
and U9853 (N_9853,N_9795,N_9774);
or U9854 (N_9854,N_9765,N_9754);
or U9855 (N_9855,N_9733,N_9730);
nand U9856 (N_9856,N_9703,N_9772);
nor U9857 (N_9857,N_9797,N_9757);
nor U9858 (N_9858,N_9764,N_9774);
or U9859 (N_9859,N_9703,N_9728);
xnor U9860 (N_9860,N_9700,N_9727);
and U9861 (N_9861,N_9740,N_9703);
nor U9862 (N_9862,N_9747,N_9749);
xnor U9863 (N_9863,N_9737,N_9725);
nand U9864 (N_9864,N_9797,N_9701);
xor U9865 (N_9865,N_9751,N_9798);
xnor U9866 (N_9866,N_9797,N_9787);
and U9867 (N_9867,N_9712,N_9794);
or U9868 (N_9868,N_9714,N_9785);
or U9869 (N_9869,N_9749,N_9720);
or U9870 (N_9870,N_9727,N_9756);
or U9871 (N_9871,N_9718,N_9740);
xnor U9872 (N_9872,N_9738,N_9728);
nor U9873 (N_9873,N_9781,N_9742);
and U9874 (N_9874,N_9784,N_9735);
and U9875 (N_9875,N_9794,N_9700);
xor U9876 (N_9876,N_9756,N_9797);
or U9877 (N_9877,N_9770,N_9752);
and U9878 (N_9878,N_9781,N_9792);
xnor U9879 (N_9879,N_9780,N_9742);
nand U9880 (N_9880,N_9791,N_9709);
nand U9881 (N_9881,N_9707,N_9753);
or U9882 (N_9882,N_9762,N_9789);
and U9883 (N_9883,N_9765,N_9774);
and U9884 (N_9884,N_9717,N_9757);
nor U9885 (N_9885,N_9773,N_9710);
nand U9886 (N_9886,N_9731,N_9733);
nand U9887 (N_9887,N_9703,N_9789);
and U9888 (N_9888,N_9799,N_9740);
or U9889 (N_9889,N_9702,N_9714);
or U9890 (N_9890,N_9737,N_9775);
or U9891 (N_9891,N_9733,N_9727);
nand U9892 (N_9892,N_9754,N_9703);
nand U9893 (N_9893,N_9787,N_9724);
and U9894 (N_9894,N_9753,N_9772);
nor U9895 (N_9895,N_9798,N_9701);
xnor U9896 (N_9896,N_9718,N_9797);
or U9897 (N_9897,N_9703,N_9727);
nand U9898 (N_9898,N_9726,N_9794);
nor U9899 (N_9899,N_9751,N_9711);
nand U9900 (N_9900,N_9870,N_9871);
and U9901 (N_9901,N_9802,N_9854);
and U9902 (N_9902,N_9817,N_9823);
nor U9903 (N_9903,N_9864,N_9840);
and U9904 (N_9904,N_9844,N_9835);
or U9905 (N_9905,N_9891,N_9833);
nor U9906 (N_9906,N_9812,N_9842);
or U9907 (N_9907,N_9892,N_9847);
or U9908 (N_9908,N_9811,N_9839);
and U9909 (N_9909,N_9845,N_9814);
nor U9910 (N_9910,N_9849,N_9857);
and U9911 (N_9911,N_9824,N_9809);
or U9912 (N_9912,N_9856,N_9825);
xnor U9913 (N_9913,N_9893,N_9882);
xnor U9914 (N_9914,N_9881,N_9841);
xor U9915 (N_9915,N_9821,N_9829);
xor U9916 (N_9916,N_9818,N_9853);
and U9917 (N_9917,N_9890,N_9828);
nor U9918 (N_9918,N_9898,N_9815);
and U9919 (N_9919,N_9800,N_9863);
or U9920 (N_9920,N_9837,N_9861);
nand U9921 (N_9921,N_9869,N_9808);
nand U9922 (N_9922,N_9826,N_9873);
xor U9923 (N_9923,N_9830,N_9836);
xor U9924 (N_9924,N_9852,N_9896);
nand U9925 (N_9925,N_9813,N_9804);
nor U9926 (N_9926,N_9875,N_9820);
nand U9927 (N_9927,N_9899,N_9860);
nor U9928 (N_9928,N_9855,N_9868);
or U9929 (N_9929,N_9832,N_9827);
xor U9930 (N_9930,N_9807,N_9838);
or U9931 (N_9931,N_9801,N_9866);
nand U9932 (N_9932,N_9806,N_9843);
xnor U9933 (N_9933,N_9858,N_9874);
and U9934 (N_9934,N_9884,N_9889);
and U9935 (N_9935,N_9810,N_9877);
xor U9936 (N_9936,N_9848,N_9805);
or U9937 (N_9937,N_9897,N_9803);
nand U9938 (N_9938,N_9822,N_9879);
or U9939 (N_9939,N_9862,N_9886);
and U9940 (N_9940,N_9885,N_9880);
xnor U9941 (N_9941,N_9816,N_9819);
nor U9942 (N_9942,N_9878,N_9876);
and U9943 (N_9943,N_9850,N_9859);
xor U9944 (N_9944,N_9895,N_9831);
nand U9945 (N_9945,N_9834,N_9888);
or U9946 (N_9946,N_9887,N_9894);
nand U9947 (N_9947,N_9865,N_9851);
nor U9948 (N_9948,N_9883,N_9872);
xnor U9949 (N_9949,N_9846,N_9867);
or U9950 (N_9950,N_9801,N_9834);
or U9951 (N_9951,N_9828,N_9843);
or U9952 (N_9952,N_9890,N_9810);
nor U9953 (N_9953,N_9871,N_9862);
and U9954 (N_9954,N_9841,N_9897);
and U9955 (N_9955,N_9892,N_9826);
and U9956 (N_9956,N_9896,N_9880);
nand U9957 (N_9957,N_9822,N_9835);
xnor U9958 (N_9958,N_9826,N_9849);
nor U9959 (N_9959,N_9833,N_9819);
or U9960 (N_9960,N_9884,N_9835);
xor U9961 (N_9961,N_9869,N_9861);
xnor U9962 (N_9962,N_9875,N_9879);
and U9963 (N_9963,N_9889,N_9882);
xor U9964 (N_9964,N_9844,N_9801);
or U9965 (N_9965,N_9894,N_9838);
or U9966 (N_9966,N_9817,N_9822);
nand U9967 (N_9967,N_9870,N_9811);
nor U9968 (N_9968,N_9863,N_9899);
or U9969 (N_9969,N_9895,N_9806);
xnor U9970 (N_9970,N_9855,N_9866);
nor U9971 (N_9971,N_9848,N_9804);
or U9972 (N_9972,N_9837,N_9887);
or U9973 (N_9973,N_9810,N_9880);
nor U9974 (N_9974,N_9809,N_9834);
nor U9975 (N_9975,N_9854,N_9856);
or U9976 (N_9976,N_9853,N_9865);
nand U9977 (N_9977,N_9898,N_9809);
nand U9978 (N_9978,N_9817,N_9814);
and U9979 (N_9979,N_9859,N_9843);
nand U9980 (N_9980,N_9870,N_9894);
nor U9981 (N_9981,N_9880,N_9835);
and U9982 (N_9982,N_9816,N_9821);
or U9983 (N_9983,N_9822,N_9854);
nor U9984 (N_9984,N_9854,N_9827);
nand U9985 (N_9985,N_9885,N_9859);
nand U9986 (N_9986,N_9893,N_9877);
nor U9987 (N_9987,N_9849,N_9897);
nand U9988 (N_9988,N_9825,N_9895);
xnor U9989 (N_9989,N_9859,N_9879);
and U9990 (N_9990,N_9804,N_9878);
nor U9991 (N_9991,N_9813,N_9803);
xor U9992 (N_9992,N_9884,N_9828);
nand U9993 (N_9993,N_9895,N_9880);
xor U9994 (N_9994,N_9844,N_9811);
or U9995 (N_9995,N_9854,N_9880);
nor U9996 (N_9996,N_9890,N_9876);
xor U9997 (N_9997,N_9832,N_9800);
and U9998 (N_9998,N_9848,N_9854);
nand U9999 (N_9999,N_9874,N_9879);
nor UO_0 (O_0,N_9923,N_9919);
xor UO_1 (O_1,N_9987,N_9984);
nand UO_2 (O_2,N_9933,N_9991);
and UO_3 (O_3,N_9947,N_9995);
and UO_4 (O_4,N_9937,N_9926);
or UO_5 (O_5,N_9992,N_9955);
nor UO_6 (O_6,N_9969,N_9924);
or UO_7 (O_7,N_9998,N_9925);
or UO_8 (O_8,N_9986,N_9972);
and UO_9 (O_9,N_9968,N_9975);
and UO_10 (O_10,N_9999,N_9951);
and UO_11 (O_11,N_9963,N_9948);
or UO_12 (O_12,N_9982,N_9942);
nand UO_13 (O_13,N_9994,N_9940);
or UO_14 (O_14,N_9959,N_9900);
xor UO_15 (O_15,N_9904,N_9962);
or UO_16 (O_16,N_9989,N_9916);
and UO_17 (O_17,N_9914,N_9954);
or UO_18 (O_18,N_9931,N_9985);
xor UO_19 (O_19,N_9901,N_9967);
xnor UO_20 (O_20,N_9910,N_9960);
and UO_21 (O_21,N_9977,N_9905);
xor UO_22 (O_22,N_9907,N_9909);
nand UO_23 (O_23,N_9929,N_9917);
or UO_24 (O_24,N_9941,N_9953);
or UO_25 (O_25,N_9974,N_9932);
and UO_26 (O_26,N_9927,N_9971);
nand UO_27 (O_27,N_9946,N_9988);
and UO_28 (O_28,N_9938,N_9966);
xor UO_29 (O_29,N_9920,N_9957);
and UO_30 (O_30,N_9915,N_9935);
nor UO_31 (O_31,N_9921,N_9936);
and UO_32 (O_32,N_9902,N_9983);
and UO_33 (O_33,N_9928,N_9976);
or UO_34 (O_34,N_9950,N_9913);
and UO_35 (O_35,N_9979,N_9908);
nand UO_36 (O_36,N_9997,N_9956);
xor UO_37 (O_37,N_9939,N_9906);
nor UO_38 (O_38,N_9964,N_9911);
and UO_39 (O_39,N_9952,N_9978);
xnor UO_40 (O_40,N_9970,N_9943);
xnor UO_41 (O_41,N_9934,N_9996);
xor UO_42 (O_42,N_9944,N_9965);
xnor UO_43 (O_43,N_9918,N_9958);
and UO_44 (O_44,N_9993,N_9990);
nor UO_45 (O_45,N_9980,N_9949);
xor UO_46 (O_46,N_9922,N_9981);
and UO_47 (O_47,N_9961,N_9973);
nor UO_48 (O_48,N_9903,N_9930);
nand UO_49 (O_49,N_9912,N_9945);
nand UO_50 (O_50,N_9919,N_9990);
xor UO_51 (O_51,N_9967,N_9951);
or UO_52 (O_52,N_9904,N_9955);
nand UO_53 (O_53,N_9993,N_9927);
and UO_54 (O_54,N_9933,N_9940);
xor UO_55 (O_55,N_9994,N_9990);
and UO_56 (O_56,N_9907,N_9980);
nor UO_57 (O_57,N_9936,N_9994);
xor UO_58 (O_58,N_9909,N_9902);
xor UO_59 (O_59,N_9920,N_9963);
or UO_60 (O_60,N_9966,N_9986);
or UO_61 (O_61,N_9923,N_9976);
xor UO_62 (O_62,N_9966,N_9955);
xnor UO_63 (O_63,N_9934,N_9963);
xnor UO_64 (O_64,N_9989,N_9967);
nor UO_65 (O_65,N_9944,N_9980);
and UO_66 (O_66,N_9965,N_9924);
nor UO_67 (O_67,N_9938,N_9991);
or UO_68 (O_68,N_9942,N_9910);
and UO_69 (O_69,N_9915,N_9967);
and UO_70 (O_70,N_9950,N_9943);
or UO_71 (O_71,N_9903,N_9971);
xnor UO_72 (O_72,N_9987,N_9992);
xor UO_73 (O_73,N_9936,N_9924);
xor UO_74 (O_74,N_9925,N_9990);
and UO_75 (O_75,N_9901,N_9989);
and UO_76 (O_76,N_9963,N_9978);
and UO_77 (O_77,N_9965,N_9902);
or UO_78 (O_78,N_9973,N_9955);
nor UO_79 (O_79,N_9972,N_9999);
nand UO_80 (O_80,N_9925,N_9930);
or UO_81 (O_81,N_9974,N_9962);
xnor UO_82 (O_82,N_9949,N_9971);
and UO_83 (O_83,N_9982,N_9933);
nand UO_84 (O_84,N_9917,N_9999);
or UO_85 (O_85,N_9986,N_9945);
nor UO_86 (O_86,N_9944,N_9962);
xor UO_87 (O_87,N_9976,N_9932);
or UO_88 (O_88,N_9937,N_9917);
and UO_89 (O_89,N_9927,N_9998);
or UO_90 (O_90,N_9926,N_9959);
or UO_91 (O_91,N_9906,N_9994);
nor UO_92 (O_92,N_9934,N_9932);
or UO_93 (O_93,N_9959,N_9924);
xnor UO_94 (O_94,N_9990,N_9968);
nor UO_95 (O_95,N_9915,N_9914);
or UO_96 (O_96,N_9979,N_9987);
or UO_97 (O_97,N_9955,N_9996);
or UO_98 (O_98,N_9912,N_9965);
and UO_99 (O_99,N_9915,N_9973);
xnor UO_100 (O_100,N_9982,N_9937);
and UO_101 (O_101,N_9927,N_9908);
or UO_102 (O_102,N_9993,N_9946);
nand UO_103 (O_103,N_9905,N_9936);
nand UO_104 (O_104,N_9962,N_9923);
or UO_105 (O_105,N_9992,N_9933);
or UO_106 (O_106,N_9946,N_9986);
xnor UO_107 (O_107,N_9923,N_9975);
nand UO_108 (O_108,N_9906,N_9970);
nand UO_109 (O_109,N_9947,N_9975);
nor UO_110 (O_110,N_9943,N_9997);
nor UO_111 (O_111,N_9998,N_9965);
nand UO_112 (O_112,N_9912,N_9900);
xor UO_113 (O_113,N_9910,N_9900);
xnor UO_114 (O_114,N_9972,N_9961);
xor UO_115 (O_115,N_9935,N_9972);
nor UO_116 (O_116,N_9984,N_9976);
xnor UO_117 (O_117,N_9976,N_9992);
nor UO_118 (O_118,N_9994,N_9961);
nor UO_119 (O_119,N_9904,N_9916);
and UO_120 (O_120,N_9908,N_9986);
xnor UO_121 (O_121,N_9900,N_9947);
or UO_122 (O_122,N_9906,N_9947);
nor UO_123 (O_123,N_9930,N_9951);
nor UO_124 (O_124,N_9928,N_9935);
xor UO_125 (O_125,N_9946,N_9958);
nor UO_126 (O_126,N_9976,N_9934);
nor UO_127 (O_127,N_9951,N_9939);
or UO_128 (O_128,N_9943,N_9908);
xnor UO_129 (O_129,N_9986,N_9983);
nand UO_130 (O_130,N_9985,N_9928);
nand UO_131 (O_131,N_9907,N_9908);
xnor UO_132 (O_132,N_9990,N_9999);
nor UO_133 (O_133,N_9930,N_9959);
xnor UO_134 (O_134,N_9960,N_9914);
nand UO_135 (O_135,N_9968,N_9979);
xor UO_136 (O_136,N_9905,N_9926);
xnor UO_137 (O_137,N_9962,N_9950);
nor UO_138 (O_138,N_9996,N_9978);
nand UO_139 (O_139,N_9940,N_9967);
and UO_140 (O_140,N_9962,N_9926);
nand UO_141 (O_141,N_9955,N_9925);
xor UO_142 (O_142,N_9910,N_9979);
xnor UO_143 (O_143,N_9972,N_9906);
or UO_144 (O_144,N_9925,N_9983);
nor UO_145 (O_145,N_9908,N_9904);
and UO_146 (O_146,N_9958,N_9960);
or UO_147 (O_147,N_9999,N_9943);
and UO_148 (O_148,N_9985,N_9911);
or UO_149 (O_149,N_9969,N_9986);
xor UO_150 (O_150,N_9972,N_9971);
nor UO_151 (O_151,N_9929,N_9968);
xor UO_152 (O_152,N_9901,N_9957);
and UO_153 (O_153,N_9925,N_9928);
nand UO_154 (O_154,N_9972,N_9925);
xor UO_155 (O_155,N_9934,N_9920);
or UO_156 (O_156,N_9928,N_9945);
xor UO_157 (O_157,N_9931,N_9963);
or UO_158 (O_158,N_9975,N_9918);
nor UO_159 (O_159,N_9916,N_9962);
nor UO_160 (O_160,N_9938,N_9982);
xnor UO_161 (O_161,N_9944,N_9957);
nand UO_162 (O_162,N_9903,N_9906);
xor UO_163 (O_163,N_9948,N_9953);
nand UO_164 (O_164,N_9930,N_9956);
or UO_165 (O_165,N_9954,N_9978);
and UO_166 (O_166,N_9960,N_9989);
or UO_167 (O_167,N_9937,N_9912);
xor UO_168 (O_168,N_9955,N_9914);
or UO_169 (O_169,N_9932,N_9948);
nor UO_170 (O_170,N_9958,N_9996);
and UO_171 (O_171,N_9982,N_9915);
nor UO_172 (O_172,N_9915,N_9904);
nand UO_173 (O_173,N_9979,N_9989);
nand UO_174 (O_174,N_9936,N_9929);
nor UO_175 (O_175,N_9980,N_9933);
xor UO_176 (O_176,N_9925,N_9917);
and UO_177 (O_177,N_9988,N_9999);
nor UO_178 (O_178,N_9995,N_9922);
xnor UO_179 (O_179,N_9933,N_9976);
nor UO_180 (O_180,N_9942,N_9948);
and UO_181 (O_181,N_9909,N_9911);
and UO_182 (O_182,N_9924,N_9909);
nand UO_183 (O_183,N_9937,N_9994);
xnor UO_184 (O_184,N_9954,N_9907);
nor UO_185 (O_185,N_9900,N_9942);
nor UO_186 (O_186,N_9921,N_9950);
and UO_187 (O_187,N_9915,N_9929);
nand UO_188 (O_188,N_9993,N_9913);
xnor UO_189 (O_189,N_9960,N_9991);
nand UO_190 (O_190,N_9929,N_9931);
xnor UO_191 (O_191,N_9931,N_9947);
xor UO_192 (O_192,N_9902,N_9984);
and UO_193 (O_193,N_9927,N_9916);
and UO_194 (O_194,N_9907,N_9915);
and UO_195 (O_195,N_9916,N_9949);
or UO_196 (O_196,N_9986,N_9902);
nand UO_197 (O_197,N_9905,N_9939);
nand UO_198 (O_198,N_9930,N_9904);
nor UO_199 (O_199,N_9965,N_9977);
and UO_200 (O_200,N_9977,N_9964);
or UO_201 (O_201,N_9967,N_9994);
xor UO_202 (O_202,N_9992,N_9928);
nand UO_203 (O_203,N_9911,N_9983);
and UO_204 (O_204,N_9913,N_9927);
or UO_205 (O_205,N_9926,N_9931);
nor UO_206 (O_206,N_9922,N_9948);
nand UO_207 (O_207,N_9901,N_9969);
nor UO_208 (O_208,N_9961,N_9988);
and UO_209 (O_209,N_9908,N_9981);
nand UO_210 (O_210,N_9927,N_9943);
nand UO_211 (O_211,N_9938,N_9955);
and UO_212 (O_212,N_9981,N_9935);
xor UO_213 (O_213,N_9984,N_9947);
or UO_214 (O_214,N_9971,N_9940);
xor UO_215 (O_215,N_9945,N_9905);
nand UO_216 (O_216,N_9958,N_9972);
xor UO_217 (O_217,N_9982,N_9978);
nor UO_218 (O_218,N_9956,N_9963);
nor UO_219 (O_219,N_9913,N_9991);
nand UO_220 (O_220,N_9981,N_9941);
nand UO_221 (O_221,N_9937,N_9976);
nand UO_222 (O_222,N_9950,N_9982);
nand UO_223 (O_223,N_9941,N_9931);
xnor UO_224 (O_224,N_9900,N_9955);
and UO_225 (O_225,N_9932,N_9999);
or UO_226 (O_226,N_9983,N_9922);
or UO_227 (O_227,N_9910,N_9982);
or UO_228 (O_228,N_9997,N_9985);
nand UO_229 (O_229,N_9929,N_9962);
nor UO_230 (O_230,N_9922,N_9936);
nand UO_231 (O_231,N_9977,N_9929);
or UO_232 (O_232,N_9928,N_9949);
nand UO_233 (O_233,N_9907,N_9964);
xor UO_234 (O_234,N_9941,N_9966);
nand UO_235 (O_235,N_9908,N_9994);
nand UO_236 (O_236,N_9974,N_9903);
xor UO_237 (O_237,N_9960,N_9967);
or UO_238 (O_238,N_9963,N_9929);
or UO_239 (O_239,N_9987,N_9965);
or UO_240 (O_240,N_9906,N_9954);
nand UO_241 (O_241,N_9911,N_9937);
nand UO_242 (O_242,N_9919,N_9922);
nand UO_243 (O_243,N_9903,N_9908);
xor UO_244 (O_244,N_9988,N_9918);
and UO_245 (O_245,N_9946,N_9904);
nand UO_246 (O_246,N_9969,N_9923);
xor UO_247 (O_247,N_9998,N_9995);
and UO_248 (O_248,N_9985,N_9902);
nor UO_249 (O_249,N_9958,N_9991);
or UO_250 (O_250,N_9959,N_9957);
nor UO_251 (O_251,N_9998,N_9990);
nor UO_252 (O_252,N_9910,N_9930);
nand UO_253 (O_253,N_9943,N_9973);
nor UO_254 (O_254,N_9953,N_9907);
nor UO_255 (O_255,N_9906,N_9962);
nand UO_256 (O_256,N_9984,N_9990);
and UO_257 (O_257,N_9947,N_9964);
nand UO_258 (O_258,N_9982,N_9902);
xnor UO_259 (O_259,N_9907,N_9916);
and UO_260 (O_260,N_9971,N_9974);
or UO_261 (O_261,N_9995,N_9929);
xnor UO_262 (O_262,N_9958,N_9995);
nor UO_263 (O_263,N_9933,N_9941);
or UO_264 (O_264,N_9934,N_9977);
xor UO_265 (O_265,N_9942,N_9913);
or UO_266 (O_266,N_9974,N_9982);
nand UO_267 (O_267,N_9924,N_9983);
nand UO_268 (O_268,N_9964,N_9969);
xor UO_269 (O_269,N_9951,N_9915);
nor UO_270 (O_270,N_9915,N_9955);
or UO_271 (O_271,N_9996,N_9900);
nor UO_272 (O_272,N_9942,N_9909);
xor UO_273 (O_273,N_9918,N_9944);
nand UO_274 (O_274,N_9960,N_9954);
xnor UO_275 (O_275,N_9985,N_9998);
nor UO_276 (O_276,N_9925,N_9909);
or UO_277 (O_277,N_9902,N_9963);
nand UO_278 (O_278,N_9970,N_9915);
nor UO_279 (O_279,N_9972,N_9978);
or UO_280 (O_280,N_9997,N_9917);
nand UO_281 (O_281,N_9933,N_9985);
xor UO_282 (O_282,N_9990,N_9956);
xor UO_283 (O_283,N_9921,N_9912);
xor UO_284 (O_284,N_9936,N_9914);
and UO_285 (O_285,N_9990,N_9910);
xnor UO_286 (O_286,N_9950,N_9979);
nand UO_287 (O_287,N_9990,N_9989);
xor UO_288 (O_288,N_9959,N_9967);
or UO_289 (O_289,N_9909,N_9981);
and UO_290 (O_290,N_9900,N_9971);
or UO_291 (O_291,N_9971,N_9928);
xnor UO_292 (O_292,N_9925,N_9911);
xor UO_293 (O_293,N_9931,N_9970);
nor UO_294 (O_294,N_9994,N_9958);
and UO_295 (O_295,N_9934,N_9904);
or UO_296 (O_296,N_9905,N_9969);
nor UO_297 (O_297,N_9962,N_9964);
nand UO_298 (O_298,N_9974,N_9956);
nand UO_299 (O_299,N_9912,N_9992);
and UO_300 (O_300,N_9949,N_9931);
nand UO_301 (O_301,N_9945,N_9975);
nand UO_302 (O_302,N_9952,N_9948);
nor UO_303 (O_303,N_9944,N_9938);
or UO_304 (O_304,N_9947,N_9941);
xnor UO_305 (O_305,N_9945,N_9937);
xnor UO_306 (O_306,N_9944,N_9988);
nand UO_307 (O_307,N_9975,N_9951);
nor UO_308 (O_308,N_9981,N_9939);
and UO_309 (O_309,N_9969,N_9948);
xor UO_310 (O_310,N_9933,N_9977);
and UO_311 (O_311,N_9984,N_9900);
nor UO_312 (O_312,N_9926,N_9979);
nor UO_313 (O_313,N_9984,N_9926);
xor UO_314 (O_314,N_9972,N_9942);
nand UO_315 (O_315,N_9926,N_9949);
and UO_316 (O_316,N_9997,N_9900);
nor UO_317 (O_317,N_9967,N_9962);
nand UO_318 (O_318,N_9980,N_9982);
nor UO_319 (O_319,N_9982,N_9998);
nand UO_320 (O_320,N_9941,N_9921);
or UO_321 (O_321,N_9917,N_9983);
nand UO_322 (O_322,N_9933,N_9912);
nor UO_323 (O_323,N_9912,N_9987);
and UO_324 (O_324,N_9977,N_9931);
or UO_325 (O_325,N_9936,N_9960);
nor UO_326 (O_326,N_9904,N_9978);
and UO_327 (O_327,N_9979,N_9935);
nor UO_328 (O_328,N_9944,N_9919);
nor UO_329 (O_329,N_9970,N_9913);
or UO_330 (O_330,N_9966,N_9900);
nand UO_331 (O_331,N_9970,N_9911);
xor UO_332 (O_332,N_9958,N_9927);
nand UO_333 (O_333,N_9922,N_9913);
or UO_334 (O_334,N_9909,N_9974);
or UO_335 (O_335,N_9991,N_9932);
nand UO_336 (O_336,N_9992,N_9939);
nor UO_337 (O_337,N_9991,N_9982);
nor UO_338 (O_338,N_9981,N_9900);
and UO_339 (O_339,N_9919,N_9955);
nor UO_340 (O_340,N_9909,N_9936);
and UO_341 (O_341,N_9931,N_9964);
nor UO_342 (O_342,N_9969,N_9921);
nand UO_343 (O_343,N_9986,N_9998);
nand UO_344 (O_344,N_9902,N_9903);
nor UO_345 (O_345,N_9938,N_9950);
and UO_346 (O_346,N_9903,N_9917);
or UO_347 (O_347,N_9915,N_9968);
xor UO_348 (O_348,N_9951,N_9956);
nand UO_349 (O_349,N_9931,N_9913);
nand UO_350 (O_350,N_9905,N_9943);
nand UO_351 (O_351,N_9966,N_9929);
nand UO_352 (O_352,N_9927,N_9975);
or UO_353 (O_353,N_9994,N_9982);
and UO_354 (O_354,N_9902,N_9912);
or UO_355 (O_355,N_9923,N_9938);
nand UO_356 (O_356,N_9952,N_9928);
or UO_357 (O_357,N_9979,N_9952);
and UO_358 (O_358,N_9984,N_9991);
nand UO_359 (O_359,N_9958,N_9982);
nand UO_360 (O_360,N_9980,N_9997);
and UO_361 (O_361,N_9967,N_9942);
nor UO_362 (O_362,N_9908,N_9916);
xor UO_363 (O_363,N_9964,N_9938);
or UO_364 (O_364,N_9993,N_9998);
nor UO_365 (O_365,N_9907,N_9956);
nor UO_366 (O_366,N_9977,N_9923);
or UO_367 (O_367,N_9902,N_9948);
xnor UO_368 (O_368,N_9933,N_9986);
nor UO_369 (O_369,N_9902,N_9979);
nor UO_370 (O_370,N_9925,N_9994);
or UO_371 (O_371,N_9900,N_9943);
nand UO_372 (O_372,N_9967,N_9922);
xor UO_373 (O_373,N_9916,N_9994);
nor UO_374 (O_374,N_9964,N_9901);
and UO_375 (O_375,N_9907,N_9944);
or UO_376 (O_376,N_9961,N_9928);
and UO_377 (O_377,N_9913,N_9985);
or UO_378 (O_378,N_9922,N_9945);
nor UO_379 (O_379,N_9919,N_9915);
and UO_380 (O_380,N_9964,N_9930);
xor UO_381 (O_381,N_9986,N_9906);
nand UO_382 (O_382,N_9915,N_9986);
nand UO_383 (O_383,N_9921,N_9976);
nand UO_384 (O_384,N_9988,N_9935);
nor UO_385 (O_385,N_9928,N_9926);
nor UO_386 (O_386,N_9920,N_9936);
or UO_387 (O_387,N_9934,N_9946);
xor UO_388 (O_388,N_9932,N_9940);
nor UO_389 (O_389,N_9974,N_9921);
and UO_390 (O_390,N_9953,N_9949);
nor UO_391 (O_391,N_9956,N_9959);
and UO_392 (O_392,N_9994,N_9921);
nand UO_393 (O_393,N_9981,N_9946);
and UO_394 (O_394,N_9948,N_9980);
xor UO_395 (O_395,N_9908,N_9947);
nand UO_396 (O_396,N_9937,N_9927);
or UO_397 (O_397,N_9956,N_9934);
or UO_398 (O_398,N_9917,N_9984);
nand UO_399 (O_399,N_9997,N_9962);
or UO_400 (O_400,N_9907,N_9925);
xnor UO_401 (O_401,N_9980,N_9964);
and UO_402 (O_402,N_9919,N_9942);
or UO_403 (O_403,N_9985,N_9936);
and UO_404 (O_404,N_9920,N_9981);
nand UO_405 (O_405,N_9922,N_9930);
or UO_406 (O_406,N_9909,N_9971);
or UO_407 (O_407,N_9954,N_9930);
nand UO_408 (O_408,N_9946,N_9970);
xor UO_409 (O_409,N_9991,N_9921);
nor UO_410 (O_410,N_9983,N_9949);
or UO_411 (O_411,N_9969,N_9935);
or UO_412 (O_412,N_9970,N_9997);
nand UO_413 (O_413,N_9911,N_9930);
or UO_414 (O_414,N_9965,N_9957);
xor UO_415 (O_415,N_9965,N_9968);
and UO_416 (O_416,N_9964,N_9906);
nor UO_417 (O_417,N_9904,N_9912);
and UO_418 (O_418,N_9913,N_9940);
xnor UO_419 (O_419,N_9979,N_9961);
and UO_420 (O_420,N_9913,N_9976);
nand UO_421 (O_421,N_9989,N_9933);
nand UO_422 (O_422,N_9923,N_9958);
xnor UO_423 (O_423,N_9987,N_9978);
or UO_424 (O_424,N_9939,N_9908);
and UO_425 (O_425,N_9925,N_9974);
or UO_426 (O_426,N_9909,N_9922);
and UO_427 (O_427,N_9918,N_9917);
nor UO_428 (O_428,N_9923,N_9974);
xnor UO_429 (O_429,N_9948,N_9915);
nor UO_430 (O_430,N_9986,N_9982);
xnor UO_431 (O_431,N_9966,N_9908);
or UO_432 (O_432,N_9994,N_9973);
and UO_433 (O_433,N_9962,N_9930);
and UO_434 (O_434,N_9907,N_9972);
or UO_435 (O_435,N_9916,N_9933);
and UO_436 (O_436,N_9920,N_9922);
xor UO_437 (O_437,N_9967,N_9956);
nand UO_438 (O_438,N_9936,N_9939);
nand UO_439 (O_439,N_9959,N_9984);
nand UO_440 (O_440,N_9987,N_9949);
nor UO_441 (O_441,N_9913,N_9966);
nand UO_442 (O_442,N_9978,N_9977);
or UO_443 (O_443,N_9981,N_9904);
nor UO_444 (O_444,N_9974,N_9979);
nand UO_445 (O_445,N_9941,N_9928);
nand UO_446 (O_446,N_9962,N_9903);
xnor UO_447 (O_447,N_9996,N_9942);
and UO_448 (O_448,N_9928,N_9939);
and UO_449 (O_449,N_9960,N_9920);
nand UO_450 (O_450,N_9978,N_9902);
nor UO_451 (O_451,N_9990,N_9927);
nand UO_452 (O_452,N_9928,N_9907);
or UO_453 (O_453,N_9912,N_9975);
nand UO_454 (O_454,N_9930,N_9929);
xor UO_455 (O_455,N_9903,N_9954);
nor UO_456 (O_456,N_9956,N_9992);
or UO_457 (O_457,N_9970,N_9957);
nand UO_458 (O_458,N_9974,N_9911);
nand UO_459 (O_459,N_9974,N_9913);
or UO_460 (O_460,N_9901,N_9970);
or UO_461 (O_461,N_9999,N_9997);
nand UO_462 (O_462,N_9997,N_9945);
xnor UO_463 (O_463,N_9931,N_9946);
xnor UO_464 (O_464,N_9996,N_9989);
nor UO_465 (O_465,N_9940,N_9960);
nor UO_466 (O_466,N_9977,N_9971);
or UO_467 (O_467,N_9992,N_9994);
xnor UO_468 (O_468,N_9931,N_9928);
nor UO_469 (O_469,N_9979,N_9931);
and UO_470 (O_470,N_9979,N_9994);
nand UO_471 (O_471,N_9930,N_9965);
xnor UO_472 (O_472,N_9954,N_9917);
or UO_473 (O_473,N_9985,N_9949);
nand UO_474 (O_474,N_9989,N_9949);
or UO_475 (O_475,N_9931,N_9942);
nand UO_476 (O_476,N_9988,N_9974);
or UO_477 (O_477,N_9924,N_9946);
xnor UO_478 (O_478,N_9929,N_9987);
or UO_479 (O_479,N_9921,N_9924);
or UO_480 (O_480,N_9989,N_9966);
and UO_481 (O_481,N_9946,N_9999);
nor UO_482 (O_482,N_9903,N_9969);
nor UO_483 (O_483,N_9973,N_9919);
or UO_484 (O_484,N_9976,N_9974);
nor UO_485 (O_485,N_9950,N_9995);
xnor UO_486 (O_486,N_9943,N_9992);
or UO_487 (O_487,N_9986,N_9952);
and UO_488 (O_488,N_9925,N_9966);
xor UO_489 (O_489,N_9977,N_9936);
nand UO_490 (O_490,N_9934,N_9938);
or UO_491 (O_491,N_9974,N_9980);
xnor UO_492 (O_492,N_9982,N_9948);
or UO_493 (O_493,N_9907,N_9990);
and UO_494 (O_494,N_9939,N_9960);
and UO_495 (O_495,N_9967,N_9983);
nor UO_496 (O_496,N_9968,N_9999);
or UO_497 (O_497,N_9922,N_9973);
and UO_498 (O_498,N_9966,N_9995);
nor UO_499 (O_499,N_9937,N_9925);
and UO_500 (O_500,N_9945,N_9972);
nand UO_501 (O_501,N_9976,N_9907);
nand UO_502 (O_502,N_9918,N_9928);
nand UO_503 (O_503,N_9977,N_9973);
xnor UO_504 (O_504,N_9926,N_9916);
nand UO_505 (O_505,N_9983,N_9964);
nand UO_506 (O_506,N_9943,N_9974);
or UO_507 (O_507,N_9916,N_9932);
xor UO_508 (O_508,N_9967,N_9908);
and UO_509 (O_509,N_9976,N_9919);
and UO_510 (O_510,N_9972,N_9903);
nand UO_511 (O_511,N_9937,N_9961);
xnor UO_512 (O_512,N_9937,N_9952);
and UO_513 (O_513,N_9978,N_9975);
xnor UO_514 (O_514,N_9908,N_9931);
or UO_515 (O_515,N_9946,N_9957);
nor UO_516 (O_516,N_9916,N_9958);
and UO_517 (O_517,N_9984,N_9930);
nor UO_518 (O_518,N_9979,N_9925);
and UO_519 (O_519,N_9957,N_9994);
nand UO_520 (O_520,N_9963,N_9995);
nor UO_521 (O_521,N_9983,N_9961);
and UO_522 (O_522,N_9995,N_9945);
and UO_523 (O_523,N_9948,N_9954);
nand UO_524 (O_524,N_9934,N_9971);
nand UO_525 (O_525,N_9955,N_9949);
xnor UO_526 (O_526,N_9941,N_9942);
xnor UO_527 (O_527,N_9916,N_9966);
xor UO_528 (O_528,N_9990,N_9911);
xor UO_529 (O_529,N_9946,N_9962);
or UO_530 (O_530,N_9939,N_9994);
nand UO_531 (O_531,N_9976,N_9922);
and UO_532 (O_532,N_9949,N_9991);
or UO_533 (O_533,N_9985,N_9954);
and UO_534 (O_534,N_9927,N_9939);
and UO_535 (O_535,N_9913,N_9996);
and UO_536 (O_536,N_9973,N_9985);
xnor UO_537 (O_537,N_9931,N_9981);
nand UO_538 (O_538,N_9981,N_9910);
or UO_539 (O_539,N_9908,N_9963);
xor UO_540 (O_540,N_9979,N_9933);
nor UO_541 (O_541,N_9904,N_9920);
nor UO_542 (O_542,N_9968,N_9924);
nand UO_543 (O_543,N_9953,N_9932);
xnor UO_544 (O_544,N_9974,N_9942);
and UO_545 (O_545,N_9964,N_9939);
nor UO_546 (O_546,N_9938,N_9935);
nor UO_547 (O_547,N_9945,N_9921);
nor UO_548 (O_548,N_9906,N_9961);
or UO_549 (O_549,N_9956,N_9975);
or UO_550 (O_550,N_9945,N_9990);
or UO_551 (O_551,N_9905,N_9967);
xor UO_552 (O_552,N_9927,N_9926);
or UO_553 (O_553,N_9915,N_9912);
and UO_554 (O_554,N_9979,N_9975);
and UO_555 (O_555,N_9900,N_9913);
and UO_556 (O_556,N_9971,N_9931);
xnor UO_557 (O_557,N_9925,N_9964);
or UO_558 (O_558,N_9929,N_9908);
nor UO_559 (O_559,N_9947,N_9978);
and UO_560 (O_560,N_9957,N_9943);
nor UO_561 (O_561,N_9924,N_9987);
or UO_562 (O_562,N_9996,N_9927);
or UO_563 (O_563,N_9968,N_9957);
nand UO_564 (O_564,N_9993,N_9952);
xor UO_565 (O_565,N_9902,N_9992);
xor UO_566 (O_566,N_9970,N_9921);
nand UO_567 (O_567,N_9939,N_9967);
nand UO_568 (O_568,N_9972,N_9941);
or UO_569 (O_569,N_9929,N_9909);
nand UO_570 (O_570,N_9915,N_9941);
nor UO_571 (O_571,N_9963,N_9940);
nand UO_572 (O_572,N_9982,N_9983);
xor UO_573 (O_573,N_9931,N_9994);
and UO_574 (O_574,N_9905,N_9919);
nor UO_575 (O_575,N_9957,N_9992);
and UO_576 (O_576,N_9995,N_9931);
or UO_577 (O_577,N_9913,N_9964);
or UO_578 (O_578,N_9946,N_9928);
xnor UO_579 (O_579,N_9930,N_9940);
nor UO_580 (O_580,N_9996,N_9907);
nand UO_581 (O_581,N_9956,N_9949);
or UO_582 (O_582,N_9987,N_9901);
and UO_583 (O_583,N_9961,N_9949);
xnor UO_584 (O_584,N_9966,N_9904);
nand UO_585 (O_585,N_9947,N_9922);
nor UO_586 (O_586,N_9935,N_9961);
nand UO_587 (O_587,N_9942,N_9923);
or UO_588 (O_588,N_9912,N_9901);
nor UO_589 (O_589,N_9915,N_9908);
nand UO_590 (O_590,N_9954,N_9996);
xnor UO_591 (O_591,N_9926,N_9912);
or UO_592 (O_592,N_9999,N_9978);
xor UO_593 (O_593,N_9932,N_9913);
nor UO_594 (O_594,N_9987,N_9975);
xor UO_595 (O_595,N_9955,N_9931);
nor UO_596 (O_596,N_9932,N_9905);
and UO_597 (O_597,N_9974,N_9939);
or UO_598 (O_598,N_9937,N_9979);
xnor UO_599 (O_599,N_9918,N_9938);
xnor UO_600 (O_600,N_9914,N_9923);
xor UO_601 (O_601,N_9908,N_9961);
or UO_602 (O_602,N_9924,N_9970);
xnor UO_603 (O_603,N_9976,N_9920);
xnor UO_604 (O_604,N_9904,N_9903);
xor UO_605 (O_605,N_9961,N_9986);
and UO_606 (O_606,N_9958,N_9979);
nor UO_607 (O_607,N_9959,N_9908);
nor UO_608 (O_608,N_9948,N_9998);
xor UO_609 (O_609,N_9992,N_9989);
nor UO_610 (O_610,N_9976,N_9936);
nor UO_611 (O_611,N_9953,N_9959);
or UO_612 (O_612,N_9971,N_9935);
xor UO_613 (O_613,N_9939,N_9950);
xor UO_614 (O_614,N_9905,N_9923);
nor UO_615 (O_615,N_9951,N_9996);
and UO_616 (O_616,N_9940,N_9989);
and UO_617 (O_617,N_9982,N_9945);
nand UO_618 (O_618,N_9974,N_9936);
nor UO_619 (O_619,N_9918,N_9954);
or UO_620 (O_620,N_9978,N_9923);
and UO_621 (O_621,N_9938,N_9929);
nor UO_622 (O_622,N_9947,N_9920);
nand UO_623 (O_623,N_9940,N_9929);
nand UO_624 (O_624,N_9954,N_9908);
nor UO_625 (O_625,N_9984,N_9915);
or UO_626 (O_626,N_9996,N_9938);
nor UO_627 (O_627,N_9946,N_9911);
xnor UO_628 (O_628,N_9932,N_9936);
nand UO_629 (O_629,N_9954,N_9935);
nor UO_630 (O_630,N_9927,N_9951);
nor UO_631 (O_631,N_9960,N_9941);
nand UO_632 (O_632,N_9924,N_9945);
nand UO_633 (O_633,N_9994,N_9951);
nor UO_634 (O_634,N_9985,N_9958);
xor UO_635 (O_635,N_9951,N_9938);
nand UO_636 (O_636,N_9996,N_9950);
nand UO_637 (O_637,N_9972,N_9951);
nor UO_638 (O_638,N_9953,N_9944);
xor UO_639 (O_639,N_9943,N_9977);
nand UO_640 (O_640,N_9980,N_9916);
xnor UO_641 (O_641,N_9942,N_9966);
or UO_642 (O_642,N_9977,N_9939);
nand UO_643 (O_643,N_9909,N_9914);
or UO_644 (O_644,N_9957,N_9933);
xnor UO_645 (O_645,N_9908,N_9974);
or UO_646 (O_646,N_9929,N_9907);
xor UO_647 (O_647,N_9939,N_9991);
nor UO_648 (O_648,N_9947,N_9938);
nor UO_649 (O_649,N_9913,N_9943);
xor UO_650 (O_650,N_9942,N_9953);
nor UO_651 (O_651,N_9942,N_9977);
nand UO_652 (O_652,N_9998,N_9978);
xnor UO_653 (O_653,N_9961,N_9910);
nand UO_654 (O_654,N_9994,N_9927);
nor UO_655 (O_655,N_9929,N_9956);
xnor UO_656 (O_656,N_9991,N_9992);
and UO_657 (O_657,N_9971,N_9916);
and UO_658 (O_658,N_9929,N_9924);
nor UO_659 (O_659,N_9989,N_9925);
xnor UO_660 (O_660,N_9954,N_9955);
xor UO_661 (O_661,N_9914,N_9902);
or UO_662 (O_662,N_9930,N_9943);
nor UO_663 (O_663,N_9964,N_9921);
nand UO_664 (O_664,N_9970,N_9958);
nor UO_665 (O_665,N_9971,N_9969);
or UO_666 (O_666,N_9943,N_9934);
xnor UO_667 (O_667,N_9970,N_9948);
or UO_668 (O_668,N_9988,N_9965);
nor UO_669 (O_669,N_9977,N_9909);
nor UO_670 (O_670,N_9946,N_9948);
xor UO_671 (O_671,N_9912,N_9991);
or UO_672 (O_672,N_9914,N_9966);
and UO_673 (O_673,N_9900,N_9952);
nor UO_674 (O_674,N_9995,N_9970);
or UO_675 (O_675,N_9929,N_9979);
nand UO_676 (O_676,N_9987,N_9964);
nand UO_677 (O_677,N_9985,N_9983);
and UO_678 (O_678,N_9901,N_9951);
xor UO_679 (O_679,N_9928,N_9953);
nand UO_680 (O_680,N_9936,N_9933);
and UO_681 (O_681,N_9991,N_9957);
xor UO_682 (O_682,N_9936,N_9916);
nor UO_683 (O_683,N_9910,N_9901);
nand UO_684 (O_684,N_9974,N_9992);
nand UO_685 (O_685,N_9917,N_9907);
nand UO_686 (O_686,N_9937,N_9977);
or UO_687 (O_687,N_9922,N_9958);
nand UO_688 (O_688,N_9956,N_9940);
and UO_689 (O_689,N_9901,N_9930);
or UO_690 (O_690,N_9927,N_9988);
nor UO_691 (O_691,N_9906,N_9932);
and UO_692 (O_692,N_9920,N_9932);
or UO_693 (O_693,N_9913,N_9973);
nor UO_694 (O_694,N_9975,N_9935);
nand UO_695 (O_695,N_9982,N_9920);
xnor UO_696 (O_696,N_9958,N_9919);
nand UO_697 (O_697,N_9979,N_9924);
and UO_698 (O_698,N_9943,N_9928);
or UO_699 (O_699,N_9999,N_9983);
xor UO_700 (O_700,N_9915,N_9916);
nand UO_701 (O_701,N_9905,N_9947);
xnor UO_702 (O_702,N_9954,N_9939);
or UO_703 (O_703,N_9951,N_9904);
and UO_704 (O_704,N_9925,N_9976);
nand UO_705 (O_705,N_9975,N_9905);
or UO_706 (O_706,N_9962,N_9931);
or UO_707 (O_707,N_9989,N_9974);
nor UO_708 (O_708,N_9956,N_9913);
and UO_709 (O_709,N_9972,N_9975);
nand UO_710 (O_710,N_9969,N_9958);
nand UO_711 (O_711,N_9935,N_9941);
xor UO_712 (O_712,N_9993,N_9941);
or UO_713 (O_713,N_9997,N_9983);
nor UO_714 (O_714,N_9933,N_9910);
and UO_715 (O_715,N_9937,N_9949);
xnor UO_716 (O_716,N_9928,N_9908);
xor UO_717 (O_717,N_9985,N_9953);
nand UO_718 (O_718,N_9973,N_9939);
nand UO_719 (O_719,N_9919,N_9982);
nor UO_720 (O_720,N_9973,N_9996);
nor UO_721 (O_721,N_9914,N_9992);
or UO_722 (O_722,N_9911,N_9981);
or UO_723 (O_723,N_9990,N_9918);
and UO_724 (O_724,N_9930,N_9976);
xor UO_725 (O_725,N_9951,N_9921);
and UO_726 (O_726,N_9997,N_9992);
xnor UO_727 (O_727,N_9988,N_9993);
nand UO_728 (O_728,N_9940,N_9985);
nand UO_729 (O_729,N_9900,N_9934);
nor UO_730 (O_730,N_9954,N_9926);
nand UO_731 (O_731,N_9975,N_9998);
xor UO_732 (O_732,N_9903,N_9901);
nor UO_733 (O_733,N_9971,N_9946);
nand UO_734 (O_734,N_9909,N_9980);
or UO_735 (O_735,N_9998,N_9920);
nand UO_736 (O_736,N_9953,N_9971);
xnor UO_737 (O_737,N_9993,N_9979);
or UO_738 (O_738,N_9947,N_9990);
or UO_739 (O_739,N_9985,N_9947);
nor UO_740 (O_740,N_9992,N_9922);
nand UO_741 (O_741,N_9917,N_9986);
xor UO_742 (O_742,N_9960,N_9994);
nor UO_743 (O_743,N_9930,N_9907);
nand UO_744 (O_744,N_9927,N_9919);
or UO_745 (O_745,N_9980,N_9921);
nor UO_746 (O_746,N_9921,N_9933);
nor UO_747 (O_747,N_9942,N_9950);
or UO_748 (O_748,N_9981,N_9987);
and UO_749 (O_749,N_9991,N_9993);
or UO_750 (O_750,N_9973,N_9965);
nor UO_751 (O_751,N_9974,N_9919);
and UO_752 (O_752,N_9928,N_9975);
nand UO_753 (O_753,N_9932,N_9957);
or UO_754 (O_754,N_9982,N_9911);
and UO_755 (O_755,N_9954,N_9932);
nor UO_756 (O_756,N_9964,N_9979);
nand UO_757 (O_757,N_9998,N_9940);
xor UO_758 (O_758,N_9907,N_9995);
or UO_759 (O_759,N_9951,N_9931);
and UO_760 (O_760,N_9992,N_9926);
nand UO_761 (O_761,N_9950,N_9992);
xor UO_762 (O_762,N_9910,N_9911);
nand UO_763 (O_763,N_9956,N_9905);
xnor UO_764 (O_764,N_9945,N_9910);
or UO_765 (O_765,N_9906,N_9921);
nor UO_766 (O_766,N_9915,N_9954);
or UO_767 (O_767,N_9960,N_9998);
xor UO_768 (O_768,N_9946,N_9919);
nand UO_769 (O_769,N_9914,N_9926);
or UO_770 (O_770,N_9963,N_9958);
nor UO_771 (O_771,N_9967,N_9948);
and UO_772 (O_772,N_9920,N_9940);
nand UO_773 (O_773,N_9980,N_9987);
or UO_774 (O_774,N_9993,N_9930);
and UO_775 (O_775,N_9966,N_9903);
nor UO_776 (O_776,N_9952,N_9980);
and UO_777 (O_777,N_9950,N_9975);
and UO_778 (O_778,N_9977,N_9906);
nand UO_779 (O_779,N_9964,N_9966);
nand UO_780 (O_780,N_9997,N_9990);
nor UO_781 (O_781,N_9913,N_9901);
nand UO_782 (O_782,N_9905,N_9917);
and UO_783 (O_783,N_9981,N_9990);
nand UO_784 (O_784,N_9981,N_9917);
nor UO_785 (O_785,N_9938,N_9921);
nand UO_786 (O_786,N_9941,N_9965);
nor UO_787 (O_787,N_9971,N_9993);
nand UO_788 (O_788,N_9924,N_9950);
or UO_789 (O_789,N_9990,N_9942);
nand UO_790 (O_790,N_9937,N_9915);
xor UO_791 (O_791,N_9977,N_9913);
xnor UO_792 (O_792,N_9998,N_9932);
nor UO_793 (O_793,N_9979,N_9934);
nand UO_794 (O_794,N_9907,N_9926);
or UO_795 (O_795,N_9959,N_9975);
xor UO_796 (O_796,N_9922,N_9977);
and UO_797 (O_797,N_9978,N_9983);
and UO_798 (O_798,N_9929,N_9947);
or UO_799 (O_799,N_9958,N_9954);
xnor UO_800 (O_800,N_9976,N_9910);
xor UO_801 (O_801,N_9972,N_9956);
and UO_802 (O_802,N_9918,N_9977);
and UO_803 (O_803,N_9946,N_9967);
nand UO_804 (O_804,N_9923,N_9924);
and UO_805 (O_805,N_9934,N_9991);
or UO_806 (O_806,N_9999,N_9931);
and UO_807 (O_807,N_9943,N_9980);
or UO_808 (O_808,N_9921,N_9900);
and UO_809 (O_809,N_9937,N_9985);
nor UO_810 (O_810,N_9910,N_9969);
xor UO_811 (O_811,N_9988,N_9994);
xnor UO_812 (O_812,N_9980,N_9972);
or UO_813 (O_813,N_9925,N_9926);
nor UO_814 (O_814,N_9943,N_9989);
or UO_815 (O_815,N_9998,N_9979);
or UO_816 (O_816,N_9985,N_9930);
nor UO_817 (O_817,N_9984,N_9994);
and UO_818 (O_818,N_9967,N_9984);
and UO_819 (O_819,N_9988,N_9958);
nand UO_820 (O_820,N_9960,N_9983);
nor UO_821 (O_821,N_9918,N_9952);
and UO_822 (O_822,N_9928,N_9981);
nand UO_823 (O_823,N_9936,N_9983);
and UO_824 (O_824,N_9920,N_9905);
nor UO_825 (O_825,N_9900,N_9990);
nand UO_826 (O_826,N_9917,N_9970);
or UO_827 (O_827,N_9948,N_9976);
nor UO_828 (O_828,N_9953,N_9969);
and UO_829 (O_829,N_9901,N_9933);
nor UO_830 (O_830,N_9944,N_9922);
nand UO_831 (O_831,N_9989,N_9995);
nor UO_832 (O_832,N_9974,N_9928);
xnor UO_833 (O_833,N_9930,N_9939);
nor UO_834 (O_834,N_9996,N_9980);
xor UO_835 (O_835,N_9996,N_9926);
nand UO_836 (O_836,N_9991,N_9947);
or UO_837 (O_837,N_9941,N_9934);
nand UO_838 (O_838,N_9974,N_9901);
and UO_839 (O_839,N_9991,N_9942);
and UO_840 (O_840,N_9919,N_9953);
or UO_841 (O_841,N_9947,N_9933);
nand UO_842 (O_842,N_9959,N_9903);
xnor UO_843 (O_843,N_9951,N_9919);
xor UO_844 (O_844,N_9970,N_9918);
nor UO_845 (O_845,N_9981,N_9996);
nor UO_846 (O_846,N_9957,N_9914);
nand UO_847 (O_847,N_9990,N_9985);
and UO_848 (O_848,N_9906,N_9990);
xor UO_849 (O_849,N_9987,N_9947);
and UO_850 (O_850,N_9994,N_9934);
xnor UO_851 (O_851,N_9941,N_9974);
nor UO_852 (O_852,N_9954,N_9929);
nand UO_853 (O_853,N_9983,N_9900);
and UO_854 (O_854,N_9908,N_9910);
nand UO_855 (O_855,N_9996,N_9957);
nor UO_856 (O_856,N_9983,N_9955);
nor UO_857 (O_857,N_9957,N_9986);
or UO_858 (O_858,N_9938,N_9984);
and UO_859 (O_859,N_9918,N_9987);
and UO_860 (O_860,N_9993,N_9996);
or UO_861 (O_861,N_9957,N_9979);
nor UO_862 (O_862,N_9917,N_9911);
nand UO_863 (O_863,N_9934,N_9903);
xnor UO_864 (O_864,N_9953,N_9996);
and UO_865 (O_865,N_9996,N_9937);
and UO_866 (O_866,N_9913,N_9967);
nor UO_867 (O_867,N_9996,N_9967);
or UO_868 (O_868,N_9919,N_9979);
and UO_869 (O_869,N_9955,N_9974);
or UO_870 (O_870,N_9908,N_9972);
nor UO_871 (O_871,N_9909,N_9973);
xnor UO_872 (O_872,N_9937,N_9905);
nor UO_873 (O_873,N_9956,N_9925);
xor UO_874 (O_874,N_9979,N_9920);
nor UO_875 (O_875,N_9901,N_9982);
or UO_876 (O_876,N_9927,N_9961);
nor UO_877 (O_877,N_9935,N_9991);
nor UO_878 (O_878,N_9939,N_9931);
or UO_879 (O_879,N_9910,N_9938);
and UO_880 (O_880,N_9951,N_9908);
and UO_881 (O_881,N_9945,N_9935);
and UO_882 (O_882,N_9966,N_9948);
nor UO_883 (O_883,N_9953,N_9902);
or UO_884 (O_884,N_9982,N_9993);
xor UO_885 (O_885,N_9941,N_9988);
or UO_886 (O_886,N_9932,N_9996);
nand UO_887 (O_887,N_9922,N_9953);
nor UO_888 (O_888,N_9964,N_9952);
or UO_889 (O_889,N_9915,N_9952);
nor UO_890 (O_890,N_9959,N_9951);
and UO_891 (O_891,N_9970,N_9934);
xnor UO_892 (O_892,N_9989,N_9935);
and UO_893 (O_893,N_9981,N_9968);
nor UO_894 (O_894,N_9932,N_9926);
xnor UO_895 (O_895,N_9917,N_9931);
or UO_896 (O_896,N_9941,N_9923);
nand UO_897 (O_897,N_9935,N_9985);
nand UO_898 (O_898,N_9937,N_9986);
nand UO_899 (O_899,N_9990,N_9914);
and UO_900 (O_900,N_9938,N_9900);
nand UO_901 (O_901,N_9906,N_9951);
nor UO_902 (O_902,N_9931,N_9935);
nor UO_903 (O_903,N_9919,N_9929);
xor UO_904 (O_904,N_9970,N_9916);
and UO_905 (O_905,N_9910,N_9954);
or UO_906 (O_906,N_9968,N_9944);
or UO_907 (O_907,N_9965,N_9943);
nand UO_908 (O_908,N_9965,N_9908);
or UO_909 (O_909,N_9957,N_9942);
or UO_910 (O_910,N_9984,N_9906);
nand UO_911 (O_911,N_9981,N_9977);
or UO_912 (O_912,N_9947,N_9914);
nor UO_913 (O_913,N_9933,N_9971);
and UO_914 (O_914,N_9993,N_9926);
nand UO_915 (O_915,N_9932,N_9942);
nand UO_916 (O_916,N_9948,N_9972);
and UO_917 (O_917,N_9956,N_9920);
nand UO_918 (O_918,N_9935,N_9967);
and UO_919 (O_919,N_9962,N_9987);
or UO_920 (O_920,N_9946,N_9937);
xnor UO_921 (O_921,N_9985,N_9987);
xnor UO_922 (O_922,N_9989,N_9970);
xor UO_923 (O_923,N_9903,N_9907);
and UO_924 (O_924,N_9939,N_9989);
nand UO_925 (O_925,N_9951,N_9987);
nand UO_926 (O_926,N_9925,N_9960);
nor UO_927 (O_927,N_9905,N_9998);
nor UO_928 (O_928,N_9995,N_9918);
and UO_929 (O_929,N_9992,N_9944);
and UO_930 (O_930,N_9912,N_9983);
or UO_931 (O_931,N_9970,N_9908);
xnor UO_932 (O_932,N_9925,N_9987);
or UO_933 (O_933,N_9905,N_9941);
nor UO_934 (O_934,N_9915,N_9931);
or UO_935 (O_935,N_9902,N_9943);
nor UO_936 (O_936,N_9929,N_9941);
nor UO_937 (O_937,N_9907,N_9914);
xnor UO_938 (O_938,N_9971,N_9952);
or UO_939 (O_939,N_9909,N_9966);
or UO_940 (O_940,N_9971,N_9912);
xor UO_941 (O_941,N_9922,N_9910);
or UO_942 (O_942,N_9973,N_9966);
nand UO_943 (O_943,N_9924,N_9971);
and UO_944 (O_944,N_9914,N_9917);
nor UO_945 (O_945,N_9950,N_9944);
nand UO_946 (O_946,N_9937,N_9920);
or UO_947 (O_947,N_9989,N_9938);
nand UO_948 (O_948,N_9959,N_9963);
and UO_949 (O_949,N_9902,N_9937);
xnor UO_950 (O_950,N_9955,N_9910);
xor UO_951 (O_951,N_9963,N_9903);
xor UO_952 (O_952,N_9969,N_9988);
and UO_953 (O_953,N_9953,N_9955);
nand UO_954 (O_954,N_9952,N_9921);
and UO_955 (O_955,N_9969,N_9908);
and UO_956 (O_956,N_9931,N_9980);
or UO_957 (O_957,N_9993,N_9961);
xor UO_958 (O_958,N_9965,N_9942);
or UO_959 (O_959,N_9947,N_9953);
nand UO_960 (O_960,N_9994,N_9978);
nand UO_961 (O_961,N_9999,N_9930);
and UO_962 (O_962,N_9912,N_9918);
and UO_963 (O_963,N_9923,N_9931);
and UO_964 (O_964,N_9914,N_9945);
nand UO_965 (O_965,N_9938,N_9968);
xnor UO_966 (O_966,N_9970,N_9935);
and UO_967 (O_967,N_9956,N_9910);
nand UO_968 (O_968,N_9904,N_9941);
or UO_969 (O_969,N_9986,N_9914);
and UO_970 (O_970,N_9967,N_9920);
or UO_971 (O_971,N_9939,N_9949);
or UO_972 (O_972,N_9958,N_9999);
and UO_973 (O_973,N_9932,N_9901);
and UO_974 (O_974,N_9981,N_9992);
nand UO_975 (O_975,N_9922,N_9934);
nor UO_976 (O_976,N_9995,N_9999);
nor UO_977 (O_977,N_9902,N_9956);
xor UO_978 (O_978,N_9937,N_9918);
nand UO_979 (O_979,N_9942,N_9943);
nand UO_980 (O_980,N_9963,N_9901);
and UO_981 (O_981,N_9970,N_9974);
or UO_982 (O_982,N_9912,N_9969);
and UO_983 (O_983,N_9909,N_9987);
and UO_984 (O_984,N_9966,N_9922);
nor UO_985 (O_985,N_9997,N_9926);
nor UO_986 (O_986,N_9986,N_9958);
or UO_987 (O_987,N_9925,N_9959);
and UO_988 (O_988,N_9947,N_9940);
xnor UO_989 (O_989,N_9906,N_9997);
or UO_990 (O_990,N_9915,N_9956);
nand UO_991 (O_991,N_9966,N_9967);
nand UO_992 (O_992,N_9964,N_9951);
nand UO_993 (O_993,N_9957,N_9954);
nand UO_994 (O_994,N_9979,N_9971);
xor UO_995 (O_995,N_9986,N_9988);
xor UO_996 (O_996,N_9921,N_9916);
and UO_997 (O_997,N_9977,N_9999);
nand UO_998 (O_998,N_9970,N_9982);
xnor UO_999 (O_999,N_9975,N_9936);
and UO_1000 (O_1000,N_9903,N_9924);
or UO_1001 (O_1001,N_9909,N_9979);
and UO_1002 (O_1002,N_9975,N_9976);
nor UO_1003 (O_1003,N_9983,N_9937);
and UO_1004 (O_1004,N_9972,N_9909);
nor UO_1005 (O_1005,N_9962,N_9959);
nand UO_1006 (O_1006,N_9976,N_9988);
xor UO_1007 (O_1007,N_9991,N_9976);
or UO_1008 (O_1008,N_9929,N_9989);
and UO_1009 (O_1009,N_9970,N_9986);
nor UO_1010 (O_1010,N_9999,N_9903);
nor UO_1011 (O_1011,N_9972,N_9955);
nor UO_1012 (O_1012,N_9952,N_9909);
and UO_1013 (O_1013,N_9916,N_9968);
or UO_1014 (O_1014,N_9939,N_9920);
and UO_1015 (O_1015,N_9949,N_9914);
or UO_1016 (O_1016,N_9928,N_9998);
and UO_1017 (O_1017,N_9908,N_9942);
or UO_1018 (O_1018,N_9980,N_9973);
xnor UO_1019 (O_1019,N_9951,N_9970);
nand UO_1020 (O_1020,N_9909,N_9951);
or UO_1021 (O_1021,N_9903,N_9943);
and UO_1022 (O_1022,N_9903,N_9998);
nor UO_1023 (O_1023,N_9924,N_9949);
nand UO_1024 (O_1024,N_9908,N_9909);
and UO_1025 (O_1025,N_9931,N_9905);
nor UO_1026 (O_1026,N_9907,N_9957);
nor UO_1027 (O_1027,N_9915,N_9945);
nand UO_1028 (O_1028,N_9995,N_9933);
nor UO_1029 (O_1029,N_9959,N_9902);
and UO_1030 (O_1030,N_9924,N_9997);
and UO_1031 (O_1031,N_9928,N_9933);
xnor UO_1032 (O_1032,N_9902,N_9910);
or UO_1033 (O_1033,N_9927,N_9917);
xnor UO_1034 (O_1034,N_9967,N_9934);
nand UO_1035 (O_1035,N_9920,N_9987);
nor UO_1036 (O_1036,N_9931,N_9933);
or UO_1037 (O_1037,N_9901,N_9941);
nand UO_1038 (O_1038,N_9949,N_9905);
or UO_1039 (O_1039,N_9978,N_9922);
xor UO_1040 (O_1040,N_9939,N_9921);
and UO_1041 (O_1041,N_9915,N_9930);
and UO_1042 (O_1042,N_9974,N_9944);
xnor UO_1043 (O_1043,N_9912,N_9956);
nand UO_1044 (O_1044,N_9917,N_9996);
xor UO_1045 (O_1045,N_9984,N_9971);
nand UO_1046 (O_1046,N_9922,N_9968);
xnor UO_1047 (O_1047,N_9974,N_9977);
nor UO_1048 (O_1048,N_9968,N_9983);
nor UO_1049 (O_1049,N_9934,N_9957);
or UO_1050 (O_1050,N_9952,N_9955);
nand UO_1051 (O_1051,N_9991,N_9969);
and UO_1052 (O_1052,N_9900,N_9960);
nand UO_1053 (O_1053,N_9915,N_9960);
and UO_1054 (O_1054,N_9906,N_9919);
nand UO_1055 (O_1055,N_9964,N_9953);
or UO_1056 (O_1056,N_9969,N_9997);
nor UO_1057 (O_1057,N_9957,N_9922);
or UO_1058 (O_1058,N_9972,N_9949);
or UO_1059 (O_1059,N_9963,N_9999);
nand UO_1060 (O_1060,N_9946,N_9940);
or UO_1061 (O_1061,N_9923,N_9934);
or UO_1062 (O_1062,N_9942,N_9901);
or UO_1063 (O_1063,N_9930,N_9912);
or UO_1064 (O_1064,N_9919,N_9909);
xor UO_1065 (O_1065,N_9965,N_9910);
nor UO_1066 (O_1066,N_9963,N_9996);
or UO_1067 (O_1067,N_9956,N_9989);
and UO_1068 (O_1068,N_9902,N_9994);
or UO_1069 (O_1069,N_9993,N_9937);
xnor UO_1070 (O_1070,N_9973,N_9927);
nor UO_1071 (O_1071,N_9988,N_9928);
nor UO_1072 (O_1072,N_9919,N_9901);
xor UO_1073 (O_1073,N_9960,N_9988);
xor UO_1074 (O_1074,N_9954,N_9920);
and UO_1075 (O_1075,N_9967,N_9952);
or UO_1076 (O_1076,N_9998,N_9984);
or UO_1077 (O_1077,N_9959,N_9976);
nor UO_1078 (O_1078,N_9909,N_9931);
or UO_1079 (O_1079,N_9956,N_9968);
nand UO_1080 (O_1080,N_9985,N_9927);
or UO_1081 (O_1081,N_9976,N_9905);
and UO_1082 (O_1082,N_9968,N_9912);
xnor UO_1083 (O_1083,N_9920,N_9946);
and UO_1084 (O_1084,N_9978,N_9919);
xor UO_1085 (O_1085,N_9949,N_9933);
and UO_1086 (O_1086,N_9995,N_9930);
nor UO_1087 (O_1087,N_9951,N_9963);
and UO_1088 (O_1088,N_9992,N_9907);
xnor UO_1089 (O_1089,N_9962,N_9991);
nand UO_1090 (O_1090,N_9939,N_9912);
nand UO_1091 (O_1091,N_9982,N_9995);
and UO_1092 (O_1092,N_9999,N_9912);
or UO_1093 (O_1093,N_9922,N_9941);
xnor UO_1094 (O_1094,N_9912,N_9960);
nand UO_1095 (O_1095,N_9962,N_9902);
nand UO_1096 (O_1096,N_9965,N_9999);
nand UO_1097 (O_1097,N_9956,N_9983);
and UO_1098 (O_1098,N_9948,N_9905);
xnor UO_1099 (O_1099,N_9948,N_9918);
and UO_1100 (O_1100,N_9992,N_9953);
nor UO_1101 (O_1101,N_9917,N_9921);
nand UO_1102 (O_1102,N_9933,N_9942);
nand UO_1103 (O_1103,N_9942,N_9925);
nor UO_1104 (O_1104,N_9957,N_9935);
and UO_1105 (O_1105,N_9932,N_9923);
and UO_1106 (O_1106,N_9930,N_9967);
nand UO_1107 (O_1107,N_9955,N_9935);
nor UO_1108 (O_1108,N_9977,N_9958);
and UO_1109 (O_1109,N_9954,N_9924);
nor UO_1110 (O_1110,N_9967,N_9938);
or UO_1111 (O_1111,N_9913,N_9946);
and UO_1112 (O_1112,N_9978,N_9933);
nand UO_1113 (O_1113,N_9946,N_9987);
nor UO_1114 (O_1114,N_9931,N_9907);
nor UO_1115 (O_1115,N_9991,N_9994);
and UO_1116 (O_1116,N_9915,N_9980);
nor UO_1117 (O_1117,N_9910,N_9974);
xnor UO_1118 (O_1118,N_9957,N_9924);
xnor UO_1119 (O_1119,N_9963,N_9923);
and UO_1120 (O_1120,N_9933,N_9964);
xnor UO_1121 (O_1121,N_9938,N_9997);
nor UO_1122 (O_1122,N_9908,N_9968);
xor UO_1123 (O_1123,N_9912,N_9910);
xnor UO_1124 (O_1124,N_9912,N_9911);
or UO_1125 (O_1125,N_9932,N_9908);
or UO_1126 (O_1126,N_9908,N_9936);
nand UO_1127 (O_1127,N_9991,N_9955);
xor UO_1128 (O_1128,N_9976,N_9965);
and UO_1129 (O_1129,N_9997,N_9984);
and UO_1130 (O_1130,N_9937,N_9955);
nand UO_1131 (O_1131,N_9955,N_9978);
or UO_1132 (O_1132,N_9930,N_9935);
or UO_1133 (O_1133,N_9943,N_9955);
nor UO_1134 (O_1134,N_9947,N_9946);
and UO_1135 (O_1135,N_9950,N_9972);
nor UO_1136 (O_1136,N_9938,N_9990);
and UO_1137 (O_1137,N_9903,N_9946);
nand UO_1138 (O_1138,N_9944,N_9975);
nor UO_1139 (O_1139,N_9937,N_9964);
or UO_1140 (O_1140,N_9942,N_9961);
or UO_1141 (O_1141,N_9970,N_9933);
and UO_1142 (O_1142,N_9974,N_9983);
xor UO_1143 (O_1143,N_9976,N_9945);
and UO_1144 (O_1144,N_9927,N_9967);
nor UO_1145 (O_1145,N_9914,N_9998);
and UO_1146 (O_1146,N_9937,N_9942);
or UO_1147 (O_1147,N_9927,N_9954);
or UO_1148 (O_1148,N_9909,N_9937);
and UO_1149 (O_1149,N_9978,N_9918);
nor UO_1150 (O_1150,N_9935,N_9943);
or UO_1151 (O_1151,N_9982,N_9956);
or UO_1152 (O_1152,N_9960,N_9986);
nor UO_1153 (O_1153,N_9980,N_9993);
and UO_1154 (O_1154,N_9984,N_9949);
nor UO_1155 (O_1155,N_9924,N_9911);
xor UO_1156 (O_1156,N_9912,N_9955);
or UO_1157 (O_1157,N_9922,N_9926);
and UO_1158 (O_1158,N_9962,N_9934);
or UO_1159 (O_1159,N_9928,N_9929);
nand UO_1160 (O_1160,N_9926,N_9952);
xnor UO_1161 (O_1161,N_9966,N_9905);
or UO_1162 (O_1162,N_9967,N_9945);
nor UO_1163 (O_1163,N_9921,N_9922);
or UO_1164 (O_1164,N_9936,N_9907);
nor UO_1165 (O_1165,N_9946,N_9943);
xnor UO_1166 (O_1166,N_9977,N_9925);
or UO_1167 (O_1167,N_9944,N_9951);
nand UO_1168 (O_1168,N_9981,N_9905);
and UO_1169 (O_1169,N_9934,N_9961);
nor UO_1170 (O_1170,N_9982,N_9955);
or UO_1171 (O_1171,N_9907,N_9999);
or UO_1172 (O_1172,N_9902,N_9900);
nand UO_1173 (O_1173,N_9946,N_9907);
nor UO_1174 (O_1174,N_9974,N_9904);
or UO_1175 (O_1175,N_9994,N_9995);
xnor UO_1176 (O_1176,N_9914,N_9950);
and UO_1177 (O_1177,N_9908,N_9914);
and UO_1178 (O_1178,N_9959,N_9972);
nand UO_1179 (O_1179,N_9936,N_9952);
nand UO_1180 (O_1180,N_9913,N_9917);
nand UO_1181 (O_1181,N_9952,N_9991);
or UO_1182 (O_1182,N_9939,N_9918);
xor UO_1183 (O_1183,N_9906,N_9946);
nor UO_1184 (O_1184,N_9958,N_9944);
or UO_1185 (O_1185,N_9980,N_9975);
or UO_1186 (O_1186,N_9984,N_9907);
nor UO_1187 (O_1187,N_9934,N_9948);
nand UO_1188 (O_1188,N_9929,N_9952);
or UO_1189 (O_1189,N_9956,N_9971);
or UO_1190 (O_1190,N_9902,N_9951);
xor UO_1191 (O_1191,N_9919,N_9998);
nand UO_1192 (O_1192,N_9999,N_9909);
xor UO_1193 (O_1193,N_9933,N_9958);
or UO_1194 (O_1194,N_9970,N_9968);
nor UO_1195 (O_1195,N_9914,N_9904);
and UO_1196 (O_1196,N_9917,N_9964);
or UO_1197 (O_1197,N_9983,N_9971);
nor UO_1198 (O_1198,N_9965,N_9958);
or UO_1199 (O_1199,N_9940,N_9923);
and UO_1200 (O_1200,N_9925,N_9945);
nor UO_1201 (O_1201,N_9967,N_9911);
or UO_1202 (O_1202,N_9901,N_9984);
or UO_1203 (O_1203,N_9937,N_9932);
and UO_1204 (O_1204,N_9935,N_9987);
and UO_1205 (O_1205,N_9966,N_9946);
nor UO_1206 (O_1206,N_9971,N_9926);
nand UO_1207 (O_1207,N_9910,N_9937);
and UO_1208 (O_1208,N_9902,N_9941);
nand UO_1209 (O_1209,N_9977,N_9932);
or UO_1210 (O_1210,N_9993,N_9965);
xnor UO_1211 (O_1211,N_9970,N_9919);
nand UO_1212 (O_1212,N_9974,N_9950);
nor UO_1213 (O_1213,N_9973,N_9953);
and UO_1214 (O_1214,N_9942,N_9968);
or UO_1215 (O_1215,N_9970,N_9959);
xor UO_1216 (O_1216,N_9986,N_9922);
or UO_1217 (O_1217,N_9976,N_9993);
nand UO_1218 (O_1218,N_9911,N_9906);
xnor UO_1219 (O_1219,N_9929,N_9901);
and UO_1220 (O_1220,N_9909,N_9968);
xor UO_1221 (O_1221,N_9946,N_9952);
nor UO_1222 (O_1222,N_9992,N_9934);
or UO_1223 (O_1223,N_9926,N_9967);
and UO_1224 (O_1224,N_9938,N_9919);
nand UO_1225 (O_1225,N_9954,N_9984);
xnor UO_1226 (O_1226,N_9999,N_9902);
nand UO_1227 (O_1227,N_9909,N_9958);
nand UO_1228 (O_1228,N_9972,N_9932);
nand UO_1229 (O_1229,N_9962,N_9953);
xnor UO_1230 (O_1230,N_9924,N_9916);
nand UO_1231 (O_1231,N_9908,N_9901);
nor UO_1232 (O_1232,N_9970,N_9912);
nand UO_1233 (O_1233,N_9911,N_9958);
nand UO_1234 (O_1234,N_9948,N_9990);
nand UO_1235 (O_1235,N_9985,N_9956);
xor UO_1236 (O_1236,N_9915,N_9959);
nor UO_1237 (O_1237,N_9981,N_9989);
and UO_1238 (O_1238,N_9991,N_9999);
or UO_1239 (O_1239,N_9948,N_9940);
nor UO_1240 (O_1240,N_9989,N_9971);
and UO_1241 (O_1241,N_9994,N_9904);
nor UO_1242 (O_1242,N_9923,N_9994);
or UO_1243 (O_1243,N_9912,N_9990);
xor UO_1244 (O_1244,N_9921,N_9925);
or UO_1245 (O_1245,N_9985,N_9961);
xnor UO_1246 (O_1246,N_9975,N_9910);
xnor UO_1247 (O_1247,N_9970,N_9975);
xor UO_1248 (O_1248,N_9927,N_9910);
xnor UO_1249 (O_1249,N_9979,N_9992);
or UO_1250 (O_1250,N_9980,N_9998);
nor UO_1251 (O_1251,N_9980,N_9945);
nand UO_1252 (O_1252,N_9931,N_9987);
or UO_1253 (O_1253,N_9933,N_9996);
nand UO_1254 (O_1254,N_9995,N_9993);
or UO_1255 (O_1255,N_9995,N_9977);
nand UO_1256 (O_1256,N_9950,N_9931);
nor UO_1257 (O_1257,N_9984,N_9957);
nor UO_1258 (O_1258,N_9900,N_9901);
nand UO_1259 (O_1259,N_9922,N_9982);
nor UO_1260 (O_1260,N_9936,N_9970);
and UO_1261 (O_1261,N_9996,N_9984);
nand UO_1262 (O_1262,N_9985,N_9944);
nor UO_1263 (O_1263,N_9937,N_9960);
and UO_1264 (O_1264,N_9919,N_9948);
nand UO_1265 (O_1265,N_9989,N_9998);
nor UO_1266 (O_1266,N_9904,N_9989);
and UO_1267 (O_1267,N_9963,N_9966);
or UO_1268 (O_1268,N_9963,N_9914);
or UO_1269 (O_1269,N_9956,N_9938);
xor UO_1270 (O_1270,N_9965,N_9946);
or UO_1271 (O_1271,N_9940,N_9938);
nor UO_1272 (O_1272,N_9934,N_9935);
and UO_1273 (O_1273,N_9942,N_9955);
nand UO_1274 (O_1274,N_9935,N_9952);
and UO_1275 (O_1275,N_9948,N_9916);
nor UO_1276 (O_1276,N_9968,N_9936);
and UO_1277 (O_1277,N_9980,N_9939);
nand UO_1278 (O_1278,N_9913,N_9998);
xnor UO_1279 (O_1279,N_9910,N_9986);
xnor UO_1280 (O_1280,N_9961,N_9955);
or UO_1281 (O_1281,N_9961,N_9984);
nor UO_1282 (O_1282,N_9925,N_9947);
or UO_1283 (O_1283,N_9949,N_9932);
xor UO_1284 (O_1284,N_9908,N_9919);
nand UO_1285 (O_1285,N_9963,N_9911);
nand UO_1286 (O_1286,N_9956,N_9966);
and UO_1287 (O_1287,N_9981,N_9912);
nand UO_1288 (O_1288,N_9977,N_9930);
xnor UO_1289 (O_1289,N_9939,N_9995);
nor UO_1290 (O_1290,N_9955,N_9916);
nand UO_1291 (O_1291,N_9942,N_9998);
or UO_1292 (O_1292,N_9926,N_9909);
and UO_1293 (O_1293,N_9900,N_9985);
nor UO_1294 (O_1294,N_9945,N_9933);
nand UO_1295 (O_1295,N_9916,N_9954);
nand UO_1296 (O_1296,N_9961,N_9950);
nor UO_1297 (O_1297,N_9928,N_9993);
nand UO_1298 (O_1298,N_9914,N_9972);
nand UO_1299 (O_1299,N_9975,N_9952);
xnor UO_1300 (O_1300,N_9964,N_9916);
and UO_1301 (O_1301,N_9991,N_9917);
nor UO_1302 (O_1302,N_9932,N_9909);
or UO_1303 (O_1303,N_9960,N_9919);
nand UO_1304 (O_1304,N_9940,N_9966);
xnor UO_1305 (O_1305,N_9909,N_9969);
xor UO_1306 (O_1306,N_9952,N_9958);
nand UO_1307 (O_1307,N_9922,N_9925);
xor UO_1308 (O_1308,N_9953,N_9983);
xnor UO_1309 (O_1309,N_9901,N_9909);
xor UO_1310 (O_1310,N_9943,N_9995);
or UO_1311 (O_1311,N_9939,N_9913);
nor UO_1312 (O_1312,N_9975,N_9941);
xor UO_1313 (O_1313,N_9992,N_9978);
and UO_1314 (O_1314,N_9915,N_9964);
nand UO_1315 (O_1315,N_9987,N_9977);
nor UO_1316 (O_1316,N_9983,N_9908);
nand UO_1317 (O_1317,N_9916,N_9902);
xor UO_1318 (O_1318,N_9960,N_9955);
nor UO_1319 (O_1319,N_9992,N_9966);
nor UO_1320 (O_1320,N_9962,N_9912);
xor UO_1321 (O_1321,N_9990,N_9988);
and UO_1322 (O_1322,N_9905,N_9970);
nand UO_1323 (O_1323,N_9975,N_9924);
and UO_1324 (O_1324,N_9948,N_9909);
nand UO_1325 (O_1325,N_9916,N_9925);
xnor UO_1326 (O_1326,N_9923,N_9900);
and UO_1327 (O_1327,N_9932,N_9915);
and UO_1328 (O_1328,N_9900,N_9999);
xnor UO_1329 (O_1329,N_9940,N_9939);
nand UO_1330 (O_1330,N_9959,N_9914);
xor UO_1331 (O_1331,N_9903,N_9978);
xnor UO_1332 (O_1332,N_9985,N_9929);
nand UO_1333 (O_1333,N_9928,N_9917);
and UO_1334 (O_1334,N_9912,N_9925);
nor UO_1335 (O_1335,N_9927,N_9932);
nor UO_1336 (O_1336,N_9975,N_9948);
nand UO_1337 (O_1337,N_9962,N_9921);
nand UO_1338 (O_1338,N_9941,N_9908);
xor UO_1339 (O_1339,N_9942,N_9995);
nor UO_1340 (O_1340,N_9911,N_9980);
nor UO_1341 (O_1341,N_9997,N_9995);
nand UO_1342 (O_1342,N_9953,N_9929);
and UO_1343 (O_1343,N_9905,N_9915);
or UO_1344 (O_1344,N_9912,N_9927);
nor UO_1345 (O_1345,N_9981,N_9976);
nand UO_1346 (O_1346,N_9916,N_9960);
nand UO_1347 (O_1347,N_9931,N_9959);
nor UO_1348 (O_1348,N_9912,N_9998);
or UO_1349 (O_1349,N_9975,N_9966);
and UO_1350 (O_1350,N_9937,N_9929);
or UO_1351 (O_1351,N_9948,N_9913);
xnor UO_1352 (O_1352,N_9924,N_9973);
xnor UO_1353 (O_1353,N_9966,N_9912);
nand UO_1354 (O_1354,N_9998,N_9943);
or UO_1355 (O_1355,N_9936,N_9971);
and UO_1356 (O_1356,N_9930,N_9933);
and UO_1357 (O_1357,N_9984,N_9941);
xnor UO_1358 (O_1358,N_9986,N_9955);
nor UO_1359 (O_1359,N_9928,N_9940);
or UO_1360 (O_1360,N_9997,N_9922);
xor UO_1361 (O_1361,N_9961,N_9956);
nor UO_1362 (O_1362,N_9957,N_9998);
nor UO_1363 (O_1363,N_9913,N_9979);
xor UO_1364 (O_1364,N_9998,N_9956);
or UO_1365 (O_1365,N_9962,N_9992);
and UO_1366 (O_1366,N_9950,N_9963);
nor UO_1367 (O_1367,N_9975,N_9955);
and UO_1368 (O_1368,N_9988,N_9936);
nor UO_1369 (O_1369,N_9955,N_9958);
nand UO_1370 (O_1370,N_9952,N_9905);
or UO_1371 (O_1371,N_9950,N_9999);
nor UO_1372 (O_1372,N_9961,N_9900);
nor UO_1373 (O_1373,N_9982,N_9921);
nor UO_1374 (O_1374,N_9922,N_9975);
and UO_1375 (O_1375,N_9960,N_9976);
nor UO_1376 (O_1376,N_9908,N_9996);
nand UO_1377 (O_1377,N_9938,N_9994);
xnor UO_1378 (O_1378,N_9992,N_9905);
xor UO_1379 (O_1379,N_9947,N_9982);
and UO_1380 (O_1380,N_9945,N_9932);
or UO_1381 (O_1381,N_9921,N_9966);
xnor UO_1382 (O_1382,N_9968,N_9976);
and UO_1383 (O_1383,N_9945,N_9963);
or UO_1384 (O_1384,N_9926,N_9960);
and UO_1385 (O_1385,N_9939,N_9937);
xnor UO_1386 (O_1386,N_9923,N_9901);
and UO_1387 (O_1387,N_9917,N_9940);
nor UO_1388 (O_1388,N_9922,N_9908);
or UO_1389 (O_1389,N_9925,N_9904);
xnor UO_1390 (O_1390,N_9925,N_9932);
nor UO_1391 (O_1391,N_9965,N_9966);
nand UO_1392 (O_1392,N_9919,N_9954);
and UO_1393 (O_1393,N_9963,N_9933);
or UO_1394 (O_1394,N_9957,N_9960);
and UO_1395 (O_1395,N_9933,N_9935);
xnor UO_1396 (O_1396,N_9952,N_9982);
nor UO_1397 (O_1397,N_9947,N_9939);
xor UO_1398 (O_1398,N_9930,N_9975);
xnor UO_1399 (O_1399,N_9928,N_9903);
xnor UO_1400 (O_1400,N_9935,N_9942);
or UO_1401 (O_1401,N_9981,N_9972);
or UO_1402 (O_1402,N_9956,N_9976);
xnor UO_1403 (O_1403,N_9966,N_9954);
or UO_1404 (O_1404,N_9968,N_9940);
nand UO_1405 (O_1405,N_9965,N_9950);
nand UO_1406 (O_1406,N_9919,N_9981);
nor UO_1407 (O_1407,N_9987,N_9916);
xnor UO_1408 (O_1408,N_9976,N_9924);
xor UO_1409 (O_1409,N_9964,N_9954);
or UO_1410 (O_1410,N_9914,N_9987);
nor UO_1411 (O_1411,N_9988,N_9981);
nand UO_1412 (O_1412,N_9983,N_9910);
xnor UO_1413 (O_1413,N_9910,N_9996);
or UO_1414 (O_1414,N_9913,N_9909);
xnor UO_1415 (O_1415,N_9936,N_9999);
or UO_1416 (O_1416,N_9990,N_9979);
nand UO_1417 (O_1417,N_9957,N_9952);
nand UO_1418 (O_1418,N_9982,N_9900);
and UO_1419 (O_1419,N_9976,N_9939);
nor UO_1420 (O_1420,N_9992,N_9919);
nor UO_1421 (O_1421,N_9978,N_9926);
or UO_1422 (O_1422,N_9941,N_9913);
xor UO_1423 (O_1423,N_9917,N_9960);
nor UO_1424 (O_1424,N_9989,N_9921);
and UO_1425 (O_1425,N_9904,N_9957);
or UO_1426 (O_1426,N_9999,N_9940);
and UO_1427 (O_1427,N_9959,N_9968);
and UO_1428 (O_1428,N_9918,N_9945);
xnor UO_1429 (O_1429,N_9938,N_9992);
xor UO_1430 (O_1430,N_9903,N_9922);
and UO_1431 (O_1431,N_9945,N_9948);
nor UO_1432 (O_1432,N_9968,N_9994);
and UO_1433 (O_1433,N_9900,N_9931);
and UO_1434 (O_1434,N_9940,N_9976);
nor UO_1435 (O_1435,N_9987,N_9941);
xnor UO_1436 (O_1436,N_9935,N_9944);
or UO_1437 (O_1437,N_9999,N_9993);
or UO_1438 (O_1438,N_9932,N_9965);
or UO_1439 (O_1439,N_9953,N_9958);
nand UO_1440 (O_1440,N_9995,N_9954);
nor UO_1441 (O_1441,N_9907,N_9941);
xor UO_1442 (O_1442,N_9946,N_9902);
xor UO_1443 (O_1443,N_9971,N_9937);
or UO_1444 (O_1444,N_9966,N_9978);
and UO_1445 (O_1445,N_9956,N_9931);
or UO_1446 (O_1446,N_9934,N_9984);
xor UO_1447 (O_1447,N_9939,N_9955);
nor UO_1448 (O_1448,N_9975,N_9901);
or UO_1449 (O_1449,N_9913,N_9995);
nor UO_1450 (O_1450,N_9991,N_9925);
and UO_1451 (O_1451,N_9916,N_9923);
xor UO_1452 (O_1452,N_9974,N_9994);
nand UO_1453 (O_1453,N_9951,N_9942);
and UO_1454 (O_1454,N_9983,N_9946);
or UO_1455 (O_1455,N_9982,N_9987);
and UO_1456 (O_1456,N_9935,N_9993);
xor UO_1457 (O_1457,N_9932,N_9903);
nand UO_1458 (O_1458,N_9990,N_9953);
and UO_1459 (O_1459,N_9954,N_9988);
nand UO_1460 (O_1460,N_9964,N_9959);
xor UO_1461 (O_1461,N_9955,N_9985);
nand UO_1462 (O_1462,N_9927,N_9921);
xnor UO_1463 (O_1463,N_9992,N_9904);
nand UO_1464 (O_1464,N_9954,N_9959);
nand UO_1465 (O_1465,N_9975,N_9997);
xor UO_1466 (O_1466,N_9933,N_9987);
xnor UO_1467 (O_1467,N_9947,N_9996);
xor UO_1468 (O_1468,N_9940,N_9918);
and UO_1469 (O_1469,N_9968,N_9963);
or UO_1470 (O_1470,N_9905,N_9964);
and UO_1471 (O_1471,N_9946,N_9991);
or UO_1472 (O_1472,N_9910,N_9939);
xor UO_1473 (O_1473,N_9988,N_9989);
and UO_1474 (O_1474,N_9928,N_9955);
nand UO_1475 (O_1475,N_9918,N_9961);
and UO_1476 (O_1476,N_9964,N_9935);
nand UO_1477 (O_1477,N_9992,N_9921);
nand UO_1478 (O_1478,N_9990,N_9972);
or UO_1479 (O_1479,N_9912,N_9958);
and UO_1480 (O_1480,N_9966,N_9906);
xnor UO_1481 (O_1481,N_9968,N_9950);
nand UO_1482 (O_1482,N_9935,N_9919);
xnor UO_1483 (O_1483,N_9994,N_9944);
xnor UO_1484 (O_1484,N_9992,N_9941);
and UO_1485 (O_1485,N_9923,N_9985);
and UO_1486 (O_1486,N_9944,N_9997);
or UO_1487 (O_1487,N_9928,N_9982);
and UO_1488 (O_1488,N_9907,N_9955);
nand UO_1489 (O_1489,N_9935,N_9973);
or UO_1490 (O_1490,N_9960,N_9931);
xnor UO_1491 (O_1491,N_9972,N_9928);
and UO_1492 (O_1492,N_9926,N_9903);
nor UO_1493 (O_1493,N_9904,N_9948);
or UO_1494 (O_1494,N_9956,N_9916);
or UO_1495 (O_1495,N_9952,N_9998);
nand UO_1496 (O_1496,N_9925,N_9973);
nand UO_1497 (O_1497,N_9986,N_9994);
nand UO_1498 (O_1498,N_9973,N_9956);
nor UO_1499 (O_1499,N_9966,N_9919);
endmodule