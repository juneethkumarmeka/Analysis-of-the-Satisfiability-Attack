module basic_750_5000_1000_2_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2505,N_2507,N_2509,N_2510,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2520,N_2521,N_2522,N_2523,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2562,N_2563,N_2564,N_2565,N_2567,N_2568,N_2569,N_2570,N_2572,N_2573,N_2575,N_2576,N_2579,N_2580,N_2581,N_2583,N_2584,N_2585,N_2586,N_2587,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2624,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2639,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2658,N_2659,N_2660,N_2661,N_2663,N_2664,N_2665,N_2666,N_2667,N_2670,N_2671,N_2674,N_2675,N_2678,N_2680,N_2682,N_2684,N_2685,N_2686,N_2687,N_2690,N_2691,N_2693,N_2694,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2734,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2751,N_2752,N_2753,N_2754,N_2755,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2767,N_2768,N_2770,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2783,N_2784,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2827,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2849,N_2850,N_2852,N_2853,N_2855,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2870,N_2871,N_2872,N_2873,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2889,N_2892,N_2893,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2906,N_2907,N_2909,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2951,N_2952,N_2953,N_2954,N_2956,N_2957,N_2958,N_2960,N_2961,N_2964,N_2966,N_2968,N_2969,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2980,N_2981,N_2982,N_2983,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3009,N_3010,N_3011,N_3012,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3021,N_3022,N_3023,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3044,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3058,N_3059,N_3060,N_3064,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3075,N_3076,N_3077,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3103,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3116,N_3117,N_3118,N_3119,N_3120,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3138,N_3140,N_3141,N_3142,N_3144,N_3146,N_3147,N_3148,N_3151,N_3152,N_3153,N_3155,N_3156,N_3157,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3170,N_3171,N_3172,N_3173,N_3174,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3196,N_3197,N_3198,N_3199,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3208,N_3209,N_3210,N_3214,N_3215,N_3216,N_3218,N_3219,N_3220,N_3221,N_3222,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3232,N_3234,N_3235,N_3236,N_3237,N_3239,N_3241,N_3242,N_3243,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3259,N_3260,N_3263,N_3264,N_3265,N_3268,N_3269,N_3270,N_3272,N_3273,N_3274,N_3275,N_3276,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3288,N_3289,N_3290,N_3291,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3314,N_3315,N_3316,N_3317,N_3318,N_3321,N_3322,N_3323,N_3324,N_3325,N_3327,N_3328,N_3329,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3339,N_3340,N_3342,N_3344,N_3346,N_3348,N_3349,N_3351,N_3352,N_3353,N_3355,N_3357,N_3358,N_3359,N_3361,N_3363,N_3365,N_3366,N_3367,N_3368,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3410,N_3413,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3423,N_3424,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3455,N_3456,N_3458,N_3460,N_3461,N_3462,N_3463,N_3464,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3474,N_3477,N_3478,N_3480,N_3481,N_3483,N_3484,N_3485,N_3486,N_3488,N_3489,N_3490,N_3491,N_3493,N_3494,N_3495,N_3496,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3509,N_3510,N_3512,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3543,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3562,N_3564,N_3565,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3601,N_3602,N_3603,N_3606,N_3608,N_3609,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3632,N_3633,N_3634,N_3635,N_3636,N_3638,N_3639,N_3640,N_3642,N_3643,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3690,N_3691,N_3692,N_3693,N_3695,N_3696,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3742,N_3743,N_3744,N_3745,N_3747,N_3748,N_3750,N_3751,N_3753,N_3754,N_3755,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3765,N_3766,N_3768,N_3769,N_3770,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3781,N_3782,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3792,N_3793,N_3794,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3808,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3823,N_3824,N_3827,N_3828,N_3829,N_3831,N_3832,N_3833,N_3834,N_3838,N_3839,N_3840,N_3841,N_3842,N_3845,N_3846,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3865,N_3866,N_3867,N_3868,N_3870,N_3871,N_3872,N_3873,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3897,N_3898,N_3899,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3919,N_3920,N_3922,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3944,N_3945,N_3946,N_3947,N_3948,N_3950,N_3951,N_3952,N_3954,N_3955,N_3956,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3969,N_3973,N_3974,N_3975,N_3977,N_3978,N_3979,N_3980,N_3982,N_3984,N_3985,N_3986,N_3988,N_3989,N_3990,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4010,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4050,N_4051,N_4052,N_4054,N_4055,N_4056,N_4058,N_4061,N_4064,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4077,N_4079,N_4080,N_4081,N_4082,N_4083,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4095,N_4096,N_4097,N_4099,N_4100,N_4101,N_4103,N_4104,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4122,N_4124,N_4125,N_4128,N_4130,N_4131,N_4133,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4149,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4168,N_4169,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4181,N_4182,N_4183,N_4184,N_4187,N_4188,N_4189,N_4192,N_4193,N_4195,N_4196,N_4197,N_4198,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4249,N_4250,N_4252,N_4254,N_4256,N_4259,N_4261,N_4263,N_4264,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4274,N_4276,N_4277,N_4278,N_4279,N_4281,N_4283,N_4284,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4294,N_4295,N_4297,N_4298,N_4299,N_4301,N_4302,N_4303,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4313,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4322,N_4323,N_4324,N_4326,N_4327,N_4329,N_4330,N_4332,N_4333,N_4334,N_4336,N_4338,N_4339,N_4340,N_4342,N_4343,N_4344,N_4347,N_4348,N_4349,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4361,N_4362,N_4364,N_4365,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4388,N_4390,N_4391,N_4392,N_4393,N_4394,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4419,N_4420,N_4421,N_4422,N_4423,N_4425,N_4426,N_4428,N_4429,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4451,N_4452,N_4453,N_4454,N_4455,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4468,N_4470,N_4471,N_4472,N_4473,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4491,N_4492,N_4493,N_4497,N_4498,N_4499,N_4500,N_4501,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4534,N_4535,N_4537,N_4538,N_4539,N_4540,N_4543,N_4544,N_4545,N_4547,N_4548,N_4549,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4562,N_4564,N_4565,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4654,N_4655,N_4658,N_4659,N_4662,N_4663,N_4664,N_4667,N_4668,N_4669,N_4671,N_4672,N_4673,N_4675,N_4677,N_4680,N_4681,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4700,N_4703,N_4704,N_4705,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4761,N_4762,N_4763,N_4765,N_4766,N_4767,N_4769,N_4771,N_4772,N_4773,N_4774,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4794,N_4795,N_4796,N_4797,N_4799,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4817,N_4818,N_4819,N_4820,N_4821,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4831,N_4832,N_4833,N_4834,N_4835,N_4837,N_4838,N_4839,N_4840,N_4842,N_4843,N_4844,N_4845,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4856,N_4857,N_4858,N_4859,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4882,N_4883,N_4884,N_4886,N_4887,N_4888,N_4890,N_4893,N_4895,N_4896,N_4898,N_4899,N_4900,N_4902,N_4903,N_4904,N_4905,N_4907,N_4908,N_4909,N_4912,N_4913,N_4916,N_4917,N_4919,N_4921,N_4924,N_4925,N_4926,N_4928,N_4929,N_4930,N_4931,N_4932,N_4935,N_4937,N_4938,N_4939,N_4941,N_4944,N_4945,N_4946,N_4947,N_4948,N_4950,N_4951,N_4952,N_4954,N_4955,N_4956,N_4957,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4993,N_4994,N_4995,N_4996,N_4997,N_4999;
and U0 (N_0,In_538,In_410);
and U1 (N_1,In_274,In_404);
nor U2 (N_2,In_110,In_509);
and U3 (N_3,In_123,In_216);
nand U4 (N_4,In_500,In_311);
nand U5 (N_5,In_493,In_263);
nand U6 (N_6,In_654,In_589);
or U7 (N_7,In_413,In_208);
nor U8 (N_8,In_597,In_47);
and U9 (N_9,In_370,In_52);
nor U10 (N_10,In_341,In_77);
or U11 (N_11,In_702,In_728);
or U12 (N_12,In_695,In_548);
nand U13 (N_13,In_667,In_448);
and U14 (N_14,In_11,In_4);
nor U15 (N_15,In_429,In_373);
or U16 (N_16,In_380,In_610);
nor U17 (N_17,In_250,In_499);
or U18 (N_18,In_22,In_359);
and U19 (N_19,In_417,In_122);
and U20 (N_20,In_89,In_419);
or U21 (N_21,In_726,In_169);
nor U22 (N_22,In_599,In_465);
xor U23 (N_23,In_662,In_506);
and U24 (N_24,In_304,In_479);
xnor U25 (N_25,In_487,In_444);
or U26 (N_26,In_649,In_660);
nand U27 (N_27,In_739,In_577);
and U28 (N_28,In_23,In_226);
and U29 (N_29,In_253,In_205);
nor U30 (N_30,In_147,In_408);
nand U31 (N_31,In_378,In_368);
nor U32 (N_32,In_194,In_232);
or U33 (N_33,In_113,In_111);
and U34 (N_34,In_320,In_102);
or U35 (N_35,In_161,In_462);
nor U36 (N_36,In_525,In_683);
nand U37 (N_37,In_257,In_530);
and U38 (N_38,In_221,In_619);
nor U39 (N_39,In_570,In_151);
and U40 (N_40,In_474,In_747);
or U41 (N_41,In_162,In_129);
or U42 (N_42,In_738,In_647);
xor U43 (N_43,In_411,In_473);
nor U44 (N_44,In_691,In_635);
xor U45 (N_45,In_547,In_222);
and U46 (N_46,In_483,In_581);
or U47 (N_47,In_273,In_246);
nand U48 (N_48,In_748,In_165);
and U49 (N_49,In_397,In_240);
or U50 (N_50,In_336,In_546);
nand U51 (N_51,In_357,In_518);
nor U52 (N_52,In_282,In_449);
nor U53 (N_53,In_426,In_14);
nor U54 (N_54,In_189,In_468);
or U55 (N_55,In_590,In_564);
and U56 (N_56,In_70,In_301);
nor U57 (N_57,In_255,In_596);
or U58 (N_58,In_171,In_729);
or U59 (N_59,In_601,In_433);
nand U60 (N_60,In_478,In_621);
nor U61 (N_61,In_134,In_634);
or U62 (N_62,In_653,In_612);
and U63 (N_63,In_219,In_394);
and U64 (N_64,In_709,In_385);
or U65 (N_65,In_158,In_715);
nand U66 (N_66,In_172,In_671);
and U67 (N_67,In_497,In_181);
nor U68 (N_68,In_107,In_54);
and U69 (N_69,In_656,In_642);
and U70 (N_70,In_507,In_455);
and U71 (N_71,In_38,In_396);
nor U72 (N_72,In_749,In_197);
and U73 (N_73,In_572,In_29);
nor U74 (N_74,In_575,In_595);
nand U75 (N_75,In_296,In_708);
or U76 (N_76,In_651,In_706);
or U77 (N_77,In_733,In_228);
nand U78 (N_78,In_167,In_399);
nand U79 (N_79,In_139,In_120);
nor U80 (N_80,In_696,In_363);
and U81 (N_81,In_223,In_18);
nand U82 (N_82,In_348,In_287);
and U83 (N_83,In_543,In_632);
nor U84 (N_84,In_157,In_115);
nand U85 (N_85,In_711,In_732);
or U86 (N_86,In_101,In_160);
nor U87 (N_87,In_20,In_608);
nor U88 (N_88,In_678,In_318);
and U89 (N_89,In_0,In_594);
or U90 (N_90,In_626,In_574);
nand U91 (N_91,In_517,In_153);
and U92 (N_92,In_637,In_367);
and U93 (N_93,In_45,In_190);
or U94 (N_94,In_482,In_213);
nor U95 (N_95,In_535,In_618);
nand U96 (N_96,In_414,In_344);
nor U97 (N_97,In_442,In_329);
nand U98 (N_98,In_150,In_5);
and U99 (N_99,In_381,In_704);
nor U100 (N_100,In_204,In_103);
and U101 (N_101,In_19,In_434);
nand U102 (N_102,In_58,In_588);
nor U103 (N_103,In_536,In_379);
xnor U104 (N_104,In_511,In_592);
nand U105 (N_105,In_37,In_403);
nor U106 (N_106,In_437,In_603);
nor U107 (N_107,In_342,In_297);
nor U108 (N_108,In_633,In_125);
nor U109 (N_109,In_523,In_571);
or U110 (N_110,In_464,In_655);
nand U111 (N_111,In_95,In_176);
nor U112 (N_112,In_461,In_544);
nor U113 (N_113,In_457,In_723);
nor U114 (N_114,In_261,In_180);
xor U115 (N_115,In_384,In_576);
xor U116 (N_116,In_217,In_259);
and U117 (N_117,In_488,In_390);
nor U118 (N_118,In_645,In_358);
or U119 (N_119,In_50,In_2);
nor U120 (N_120,In_389,In_227);
and U121 (N_121,In_431,In_604);
nand U122 (N_122,In_268,In_406);
nor U123 (N_123,In_475,In_352);
or U124 (N_124,In_405,In_314);
and U125 (N_125,In_489,In_270);
nand U126 (N_126,In_108,In_224);
or U127 (N_127,In_423,In_557);
nand U128 (N_128,In_212,In_133);
and U129 (N_129,In_556,In_96);
or U130 (N_130,In_420,In_100);
nor U131 (N_131,In_361,In_606);
and U132 (N_132,In_16,In_13);
and U133 (N_133,In_476,In_229);
nand U134 (N_134,In_104,In_365);
and U135 (N_135,In_39,In_681);
or U136 (N_136,In_531,In_552);
and U137 (N_137,In_400,In_459);
nor U138 (N_138,In_533,In_332);
nand U139 (N_139,In_707,In_279);
nor U140 (N_140,In_193,In_562);
nor U141 (N_141,In_99,In_545);
or U142 (N_142,In_131,In_540);
or U143 (N_143,In_485,In_141);
or U144 (N_144,In_266,In_542);
nor U145 (N_145,In_364,In_687);
nor U146 (N_146,In_249,In_744);
and U147 (N_147,In_6,In_712);
and U148 (N_148,In_92,In_623);
nor U149 (N_149,In_166,In_10);
and U150 (N_150,In_554,In_407);
nand U151 (N_151,In_532,In_549);
nor U152 (N_152,In_196,In_666);
or U153 (N_153,In_34,In_272);
and U154 (N_154,In_665,In_105);
or U155 (N_155,In_456,In_472);
nor U156 (N_156,In_9,In_74);
nand U157 (N_157,In_701,In_534);
nor U158 (N_158,In_191,In_652);
nand U159 (N_159,In_55,In_425);
or U160 (N_160,In_236,In_602);
nor U161 (N_161,In_119,In_522);
nor U162 (N_162,In_724,In_395);
nor U163 (N_163,In_199,In_607);
nor U164 (N_164,In_614,In_322);
nor U165 (N_165,In_63,In_309);
or U166 (N_166,In_290,In_27);
nor U167 (N_167,In_112,In_713);
nor U168 (N_168,In_558,In_251);
and U169 (N_169,In_583,In_211);
and U170 (N_170,In_369,In_585);
or U171 (N_171,In_669,In_516);
nor U172 (N_172,In_690,In_638);
nor U173 (N_173,In_351,In_502);
nor U174 (N_174,In_62,In_137);
nand U175 (N_175,In_559,In_186);
or U176 (N_176,In_742,In_675);
nor U177 (N_177,In_294,In_391);
and U178 (N_178,In_560,In_680);
or U179 (N_179,In_7,In_121);
or U180 (N_180,In_512,In_452);
or U181 (N_181,In_699,In_285);
xor U182 (N_182,In_267,In_555);
nand U183 (N_183,In_625,In_349);
nand U184 (N_184,In_505,In_31);
and U185 (N_185,In_491,In_75);
nand U186 (N_186,In_68,In_321);
or U187 (N_187,In_584,In_106);
and U188 (N_188,In_245,In_41);
and U189 (N_189,In_254,In_644);
or U190 (N_190,In_288,In_537);
nand U191 (N_191,In_484,In_46);
or U192 (N_192,In_234,In_731);
and U193 (N_193,In_173,In_382);
nand U194 (N_194,In_163,In_356);
and U195 (N_195,In_82,In_53);
or U196 (N_196,In_582,In_83);
nand U197 (N_197,In_412,In_243);
and U198 (N_198,In_611,In_114);
nand U199 (N_199,In_568,In_1);
and U200 (N_200,In_90,In_278);
nor U201 (N_201,In_354,In_539);
or U202 (N_202,In_143,In_477);
and U203 (N_203,In_438,In_646);
xnor U204 (N_204,In_244,In_424);
or U205 (N_205,In_622,In_237);
and U206 (N_206,In_231,In_230);
or U207 (N_207,In_620,In_480);
or U208 (N_208,In_374,In_627);
nor U209 (N_209,In_686,In_605);
and U210 (N_210,In_60,In_293);
and U211 (N_211,In_175,In_284);
and U212 (N_212,In_513,In_44);
nand U213 (N_213,In_496,In_659);
or U214 (N_214,In_203,In_387);
and U215 (N_215,In_519,In_269);
nor U216 (N_216,In_503,In_684);
or U217 (N_217,In_201,In_362);
nand U218 (N_218,In_93,In_586);
nor U219 (N_219,In_94,In_78);
or U220 (N_220,In_127,In_640);
and U221 (N_221,In_692,In_206);
nor U222 (N_222,In_734,In_30);
nor U223 (N_223,In_520,In_312);
and U224 (N_224,In_366,In_703);
or U225 (N_225,In_593,In_214);
and U226 (N_226,In_639,In_565);
nand U227 (N_227,In_719,In_737);
nor U228 (N_228,In_315,In_298);
or U229 (N_229,In_116,In_215);
or U230 (N_230,In_170,In_3);
and U231 (N_231,In_25,In_275);
xor U232 (N_232,In_51,In_73);
or U233 (N_233,In_705,In_722);
or U234 (N_234,In_392,In_636);
nand U235 (N_235,In_710,In_310);
and U236 (N_236,In_136,In_436);
and U237 (N_237,In_154,In_745);
nand U238 (N_238,In_688,In_567);
nand U239 (N_239,In_24,In_587);
and U240 (N_240,In_643,In_156);
nand U241 (N_241,In_432,In_741);
or U242 (N_242,In_551,In_714);
nand U243 (N_243,In_42,In_353);
and U244 (N_244,In_561,In_679);
nor U245 (N_245,In_118,In_550);
and U246 (N_246,In_616,In_727);
and U247 (N_247,In_325,In_628);
or U248 (N_248,In_360,In_730);
and U249 (N_249,In_591,In_168);
nor U250 (N_250,In_388,In_164);
nand U251 (N_251,In_721,In_71);
and U252 (N_252,In_326,In_345);
nor U253 (N_253,In_441,In_598);
and U254 (N_254,In_260,In_661);
nor U255 (N_255,In_689,In_323);
nand U256 (N_256,In_280,In_508);
or U257 (N_257,In_641,In_182);
or U258 (N_258,In_339,In_693);
or U259 (N_259,In_184,In_80);
nor U260 (N_260,In_615,In_674);
and U261 (N_261,In_447,In_126);
and U262 (N_262,In_685,In_198);
or U263 (N_263,In_736,In_343);
and U264 (N_264,In_117,In_265);
or U265 (N_265,In_481,In_415);
nand U266 (N_266,In_553,In_81);
nand U267 (N_267,In_347,In_264);
nand U268 (N_268,In_295,In_490);
nand U269 (N_269,In_498,In_277);
or U270 (N_270,In_657,In_676);
nor U271 (N_271,In_28,In_252);
nand U272 (N_272,In_200,In_694);
xnor U273 (N_273,In_372,In_393);
and U274 (N_274,In_218,In_91);
nor U275 (N_275,In_578,In_398);
or U276 (N_276,In_409,In_242);
nor U277 (N_277,In_317,In_299);
and U278 (N_278,In_664,In_48);
nand U279 (N_279,In_256,In_526);
nand U280 (N_280,In_207,In_210);
or U281 (N_281,In_276,In_40);
and U282 (N_282,In_743,In_631);
nand U283 (N_283,In_155,In_109);
nand U284 (N_284,In_566,In_375);
nand U285 (N_285,In_289,In_446);
or U286 (N_286,In_527,In_12);
nor U287 (N_287,In_454,In_677);
and U288 (N_288,In_430,In_673);
nand U289 (N_289,In_418,In_271);
nor U290 (N_290,In_128,In_460);
nor U291 (N_291,In_350,In_510);
nor U292 (N_292,In_187,In_178);
or U293 (N_293,In_371,In_306);
and U294 (N_294,In_87,In_152);
and U295 (N_295,In_140,In_672);
nor U296 (N_296,In_401,In_466);
and U297 (N_297,In_233,In_428);
and U298 (N_298,In_579,In_629);
nand U299 (N_299,In_146,In_541);
or U300 (N_300,In_248,In_346);
nor U301 (N_301,In_239,In_15);
nor U302 (N_302,In_177,In_700);
nor U303 (N_303,In_624,In_528);
nor U304 (N_304,In_17,In_377);
nand U305 (N_305,In_658,In_88);
and U306 (N_306,In_331,In_86);
nor U307 (N_307,In_529,In_340);
nor U308 (N_308,In_35,In_670);
and U309 (N_309,In_79,In_65);
or U310 (N_310,In_439,In_327);
nor U311 (N_311,In_85,In_26);
nand U312 (N_312,In_292,In_179);
nand U313 (N_313,In_192,In_716);
or U314 (N_314,In_355,In_600);
or U315 (N_315,In_450,In_64);
nor U316 (N_316,In_258,In_334);
nand U317 (N_317,In_142,In_569);
nor U318 (N_318,In_328,In_613);
xnor U319 (N_319,In_335,In_67);
nand U320 (N_320,In_453,In_471);
or U321 (N_321,In_698,In_43);
or U322 (N_322,In_427,In_458);
nor U323 (N_323,In_445,In_36);
and U324 (N_324,In_72,In_663);
nand U325 (N_325,In_573,In_32);
and U326 (N_326,In_202,In_33);
and U327 (N_327,In_61,In_98);
or U328 (N_328,In_386,In_300);
nand U329 (N_329,In_333,In_337);
and U330 (N_330,In_338,In_286);
nor U331 (N_331,In_746,In_144);
and U332 (N_332,In_241,In_183);
or U333 (N_333,In_124,In_49);
and U334 (N_334,In_735,In_185);
xnor U335 (N_335,In_308,In_580);
nand U336 (N_336,In_281,In_76);
or U337 (N_337,In_402,In_247);
nor U338 (N_338,In_435,In_291);
and U339 (N_339,In_718,In_563);
nor U340 (N_340,In_303,In_97);
nor U341 (N_341,In_59,In_443);
or U342 (N_342,In_469,In_69);
or U343 (N_343,In_467,In_21);
nor U344 (N_344,In_188,In_725);
nand U345 (N_345,In_514,In_305);
xnor U346 (N_346,In_440,In_138);
xor U347 (N_347,In_422,In_494);
nor U348 (N_348,In_682,In_316);
and U349 (N_349,In_225,In_524);
or U350 (N_350,In_463,In_149);
or U351 (N_351,In_145,In_501);
nor U352 (N_352,In_8,In_330);
or U353 (N_353,In_130,In_668);
nand U354 (N_354,In_421,In_720);
or U355 (N_355,In_504,In_235);
and U356 (N_356,In_84,In_238);
nor U357 (N_357,In_220,In_630);
nor U358 (N_358,In_495,In_650);
nor U359 (N_359,In_283,In_648);
nor U360 (N_360,In_319,In_521);
nor U361 (N_361,In_302,In_66);
or U362 (N_362,In_609,In_451);
nor U363 (N_363,In_492,In_313);
nor U364 (N_364,In_376,In_515);
or U365 (N_365,In_56,In_383);
and U366 (N_366,In_324,In_135);
nor U367 (N_367,In_307,In_195);
xor U368 (N_368,In_617,In_262);
nor U369 (N_369,In_486,In_57);
or U370 (N_370,In_159,In_470);
or U371 (N_371,In_697,In_174);
and U372 (N_372,In_416,In_148);
and U373 (N_373,In_740,In_132);
or U374 (N_374,In_717,In_209);
nand U375 (N_375,In_539,In_95);
nand U376 (N_376,In_158,In_599);
or U377 (N_377,In_616,In_436);
nor U378 (N_378,In_76,In_166);
nor U379 (N_379,In_729,In_569);
nor U380 (N_380,In_368,In_41);
nor U381 (N_381,In_35,In_205);
and U382 (N_382,In_575,In_551);
or U383 (N_383,In_459,In_512);
or U384 (N_384,In_368,In_141);
nor U385 (N_385,In_12,In_225);
or U386 (N_386,In_224,In_205);
or U387 (N_387,In_264,In_312);
and U388 (N_388,In_612,In_72);
nor U389 (N_389,In_82,In_326);
or U390 (N_390,In_604,In_740);
nor U391 (N_391,In_37,In_29);
or U392 (N_392,In_710,In_411);
nor U393 (N_393,In_432,In_341);
or U394 (N_394,In_213,In_317);
or U395 (N_395,In_725,In_582);
and U396 (N_396,In_312,In_53);
or U397 (N_397,In_571,In_529);
nor U398 (N_398,In_523,In_52);
nand U399 (N_399,In_548,In_197);
or U400 (N_400,In_7,In_322);
nand U401 (N_401,In_566,In_690);
and U402 (N_402,In_237,In_167);
nand U403 (N_403,In_54,In_159);
nand U404 (N_404,In_267,In_226);
and U405 (N_405,In_650,In_331);
and U406 (N_406,In_596,In_576);
and U407 (N_407,In_38,In_319);
nand U408 (N_408,In_590,In_445);
nand U409 (N_409,In_738,In_95);
nor U410 (N_410,In_81,In_378);
nor U411 (N_411,In_611,In_358);
xnor U412 (N_412,In_54,In_99);
nand U413 (N_413,In_196,In_125);
nor U414 (N_414,In_373,In_181);
nor U415 (N_415,In_684,In_340);
nor U416 (N_416,In_319,In_281);
xor U417 (N_417,In_530,In_210);
or U418 (N_418,In_647,In_281);
and U419 (N_419,In_603,In_120);
and U420 (N_420,In_150,In_540);
nor U421 (N_421,In_551,In_421);
and U422 (N_422,In_357,In_132);
nor U423 (N_423,In_639,In_26);
and U424 (N_424,In_182,In_577);
nand U425 (N_425,In_720,In_237);
nand U426 (N_426,In_652,In_432);
and U427 (N_427,In_221,In_502);
nor U428 (N_428,In_119,In_270);
or U429 (N_429,In_260,In_558);
or U430 (N_430,In_321,In_263);
and U431 (N_431,In_636,In_178);
nor U432 (N_432,In_283,In_133);
nand U433 (N_433,In_474,In_91);
nor U434 (N_434,In_554,In_393);
nor U435 (N_435,In_222,In_439);
nor U436 (N_436,In_427,In_1);
or U437 (N_437,In_60,In_744);
nor U438 (N_438,In_670,In_195);
nor U439 (N_439,In_61,In_153);
or U440 (N_440,In_228,In_518);
or U441 (N_441,In_117,In_216);
nand U442 (N_442,In_446,In_604);
and U443 (N_443,In_392,In_409);
and U444 (N_444,In_182,In_312);
and U445 (N_445,In_482,In_130);
and U446 (N_446,In_503,In_156);
nor U447 (N_447,In_640,In_528);
and U448 (N_448,In_159,In_693);
nand U449 (N_449,In_391,In_617);
or U450 (N_450,In_118,In_364);
and U451 (N_451,In_314,In_396);
or U452 (N_452,In_525,In_466);
or U453 (N_453,In_565,In_107);
and U454 (N_454,In_551,In_628);
nor U455 (N_455,In_208,In_570);
or U456 (N_456,In_335,In_599);
nor U457 (N_457,In_258,In_160);
nand U458 (N_458,In_4,In_223);
nand U459 (N_459,In_447,In_277);
nand U460 (N_460,In_207,In_627);
and U461 (N_461,In_399,In_284);
and U462 (N_462,In_77,In_157);
and U463 (N_463,In_276,In_743);
nor U464 (N_464,In_580,In_273);
and U465 (N_465,In_129,In_138);
nor U466 (N_466,In_319,In_181);
or U467 (N_467,In_267,In_426);
or U468 (N_468,In_618,In_651);
xor U469 (N_469,In_526,In_614);
or U470 (N_470,In_265,In_56);
or U471 (N_471,In_745,In_599);
nand U472 (N_472,In_106,In_350);
nand U473 (N_473,In_23,In_725);
and U474 (N_474,In_64,In_524);
and U475 (N_475,In_424,In_8);
nand U476 (N_476,In_649,In_453);
and U477 (N_477,In_505,In_731);
and U478 (N_478,In_562,In_204);
and U479 (N_479,In_699,In_96);
nor U480 (N_480,In_329,In_393);
nor U481 (N_481,In_416,In_453);
or U482 (N_482,In_497,In_417);
and U483 (N_483,In_83,In_589);
nor U484 (N_484,In_352,In_71);
and U485 (N_485,In_459,In_726);
nand U486 (N_486,In_607,In_580);
nand U487 (N_487,In_290,In_78);
nand U488 (N_488,In_606,In_32);
nor U489 (N_489,In_195,In_122);
or U490 (N_490,In_705,In_16);
or U491 (N_491,In_309,In_107);
nand U492 (N_492,In_179,In_31);
and U493 (N_493,In_563,In_674);
nor U494 (N_494,In_349,In_486);
or U495 (N_495,In_260,In_98);
nand U496 (N_496,In_157,In_430);
nand U497 (N_497,In_464,In_95);
nor U498 (N_498,In_728,In_425);
nand U499 (N_499,In_141,In_364);
nor U500 (N_500,In_222,In_462);
or U501 (N_501,In_205,In_113);
nand U502 (N_502,In_693,In_464);
and U503 (N_503,In_309,In_450);
and U504 (N_504,In_104,In_748);
nand U505 (N_505,In_390,In_184);
and U506 (N_506,In_608,In_733);
and U507 (N_507,In_307,In_682);
nand U508 (N_508,In_684,In_565);
nor U509 (N_509,In_293,In_243);
and U510 (N_510,In_503,In_557);
nor U511 (N_511,In_7,In_87);
or U512 (N_512,In_619,In_235);
or U513 (N_513,In_702,In_220);
nand U514 (N_514,In_595,In_601);
nor U515 (N_515,In_449,In_724);
nor U516 (N_516,In_370,In_576);
nor U517 (N_517,In_105,In_504);
and U518 (N_518,In_41,In_10);
nand U519 (N_519,In_116,In_109);
and U520 (N_520,In_79,In_666);
nand U521 (N_521,In_45,In_131);
or U522 (N_522,In_576,In_121);
nand U523 (N_523,In_316,In_597);
nor U524 (N_524,In_275,In_3);
and U525 (N_525,In_705,In_236);
and U526 (N_526,In_193,In_154);
nand U527 (N_527,In_143,In_749);
nand U528 (N_528,In_386,In_646);
nand U529 (N_529,In_333,In_587);
nor U530 (N_530,In_645,In_476);
or U531 (N_531,In_549,In_40);
or U532 (N_532,In_584,In_627);
nand U533 (N_533,In_692,In_191);
nor U534 (N_534,In_84,In_208);
nand U535 (N_535,In_724,In_544);
or U536 (N_536,In_31,In_53);
and U537 (N_537,In_501,In_296);
or U538 (N_538,In_182,In_648);
and U539 (N_539,In_421,In_57);
or U540 (N_540,In_590,In_725);
or U541 (N_541,In_581,In_455);
nand U542 (N_542,In_607,In_519);
nand U543 (N_543,In_578,In_46);
or U544 (N_544,In_322,In_741);
nand U545 (N_545,In_532,In_350);
or U546 (N_546,In_269,In_233);
nand U547 (N_547,In_180,In_547);
or U548 (N_548,In_710,In_716);
nand U549 (N_549,In_645,In_341);
nor U550 (N_550,In_719,In_509);
nor U551 (N_551,In_175,In_626);
nor U552 (N_552,In_460,In_296);
nand U553 (N_553,In_235,In_80);
or U554 (N_554,In_368,In_66);
nor U555 (N_555,In_632,In_484);
nand U556 (N_556,In_598,In_649);
nor U557 (N_557,In_473,In_413);
nor U558 (N_558,In_93,In_390);
nor U559 (N_559,In_2,In_711);
nor U560 (N_560,In_719,In_144);
or U561 (N_561,In_489,In_725);
nand U562 (N_562,In_657,In_61);
nor U563 (N_563,In_447,In_169);
or U564 (N_564,In_241,In_573);
nand U565 (N_565,In_188,In_569);
xor U566 (N_566,In_367,In_198);
and U567 (N_567,In_47,In_375);
nor U568 (N_568,In_318,In_168);
nor U569 (N_569,In_322,In_77);
nand U570 (N_570,In_323,In_59);
nor U571 (N_571,In_544,In_181);
or U572 (N_572,In_254,In_745);
or U573 (N_573,In_154,In_209);
nor U574 (N_574,In_544,In_74);
and U575 (N_575,In_621,In_346);
nor U576 (N_576,In_137,In_322);
or U577 (N_577,In_148,In_208);
nor U578 (N_578,In_508,In_575);
or U579 (N_579,In_726,In_202);
nor U580 (N_580,In_541,In_479);
or U581 (N_581,In_306,In_312);
or U582 (N_582,In_204,In_640);
or U583 (N_583,In_505,In_432);
or U584 (N_584,In_451,In_618);
and U585 (N_585,In_117,In_676);
and U586 (N_586,In_144,In_717);
nand U587 (N_587,In_80,In_401);
nor U588 (N_588,In_470,In_15);
and U589 (N_589,In_228,In_545);
xnor U590 (N_590,In_711,In_686);
nand U591 (N_591,In_297,In_300);
nand U592 (N_592,In_404,In_678);
and U593 (N_593,In_131,In_95);
nor U594 (N_594,In_387,In_162);
xor U595 (N_595,In_137,In_518);
nand U596 (N_596,In_275,In_652);
xnor U597 (N_597,In_462,In_620);
nand U598 (N_598,In_623,In_355);
nor U599 (N_599,In_445,In_580);
nand U600 (N_600,In_703,In_448);
and U601 (N_601,In_651,In_539);
or U602 (N_602,In_40,In_718);
and U603 (N_603,In_680,In_134);
nor U604 (N_604,In_178,In_590);
and U605 (N_605,In_693,In_597);
and U606 (N_606,In_448,In_520);
or U607 (N_607,In_333,In_360);
nand U608 (N_608,In_508,In_36);
and U609 (N_609,In_23,In_6);
nand U610 (N_610,In_496,In_331);
nor U611 (N_611,In_556,In_329);
nand U612 (N_612,In_3,In_98);
or U613 (N_613,In_679,In_532);
or U614 (N_614,In_633,In_732);
nand U615 (N_615,In_67,In_41);
and U616 (N_616,In_266,In_575);
and U617 (N_617,In_302,In_480);
or U618 (N_618,In_225,In_13);
or U619 (N_619,In_680,In_194);
nor U620 (N_620,In_429,In_569);
or U621 (N_621,In_527,In_324);
or U622 (N_622,In_646,In_624);
nor U623 (N_623,In_348,In_102);
or U624 (N_624,In_95,In_582);
or U625 (N_625,In_461,In_712);
xnor U626 (N_626,In_129,In_558);
nor U627 (N_627,In_627,In_356);
nand U628 (N_628,In_720,In_561);
or U629 (N_629,In_67,In_455);
nor U630 (N_630,In_620,In_572);
and U631 (N_631,In_62,In_443);
and U632 (N_632,In_128,In_538);
nor U633 (N_633,In_53,In_49);
nor U634 (N_634,In_29,In_106);
xnor U635 (N_635,In_447,In_511);
xor U636 (N_636,In_428,In_114);
and U637 (N_637,In_291,In_391);
nand U638 (N_638,In_285,In_298);
nor U639 (N_639,In_107,In_683);
nand U640 (N_640,In_191,In_108);
or U641 (N_641,In_178,In_567);
xnor U642 (N_642,In_706,In_562);
nor U643 (N_643,In_591,In_469);
nor U644 (N_644,In_245,In_107);
nor U645 (N_645,In_662,In_422);
nor U646 (N_646,In_536,In_608);
nand U647 (N_647,In_56,In_328);
and U648 (N_648,In_508,In_181);
or U649 (N_649,In_249,In_358);
and U650 (N_650,In_479,In_600);
or U651 (N_651,In_395,In_462);
nor U652 (N_652,In_408,In_392);
or U653 (N_653,In_123,In_204);
or U654 (N_654,In_550,In_155);
nor U655 (N_655,In_508,In_501);
and U656 (N_656,In_496,In_247);
and U657 (N_657,In_142,In_91);
nor U658 (N_658,In_676,In_265);
or U659 (N_659,In_665,In_318);
nor U660 (N_660,In_406,In_738);
or U661 (N_661,In_59,In_148);
and U662 (N_662,In_536,In_442);
nor U663 (N_663,In_10,In_709);
or U664 (N_664,In_389,In_200);
nor U665 (N_665,In_328,In_366);
or U666 (N_666,In_229,In_689);
and U667 (N_667,In_292,In_337);
xnor U668 (N_668,In_231,In_497);
nor U669 (N_669,In_637,In_68);
nor U670 (N_670,In_575,In_686);
or U671 (N_671,In_209,In_648);
nand U672 (N_672,In_576,In_253);
nand U673 (N_673,In_330,In_236);
nor U674 (N_674,In_373,In_645);
nor U675 (N_675,In_439,In_355);
xnor U676 (N_676,In_684,In_118);
nor U677 (N_677,In_334,In_76);
nor U678 (N_678,In_743,In_424);
and U679 (N_679,In_207,In_28);
nor U680 (N_680,In_13,In_25);
xnor U681 (N_681,In_261,In_656);
or U682 (N_682,In_363,In_278);
or U683 (N_683,In_473,In_188);
nor U684 (N_684,In_544,In_253);
and U685 (N_685,In_698,In_567);
or U686 (N_686,In_543,In_688);
and U687 (N_687,In_116,In_262);
or U688 (N_688,In_572,In_426);
xnor U689 (N_689,In_455,In_659);
xor U690 (N_690,In_138,In_409);
or U691 (N_691,In_164,In_168);
or U692 (N_692,In_34,In_452);
xor U693 (N_693,In_433,In_521);
nor U694 (N_694,In_401,In_500);
nor U695 (N_695,In_281,In_589);
or U696 (N_696,In_610,In_180);
or U697 (N_697,In_206,In_150);
nor U698 (N_698,In_257,In_343);
nand U699 (N_699,In_408,In_575);
or U700 (N_700,In_149,In_84);
and U701 (N_701,In_618,In_88);
and U702 (N_702,In_315,In_694);
and U703 (N_703,In_306,In_120);
and U704 (N_704,In_705,In_544);
nor U705 (N_705,In_374,In_196);
and U706 (N_706,In_735,In_314);
or U707 (N_707,In_9,In_230);
nand U708 (N_708,In_461,In_226);
nand U709 (N_709,In_475,In_617);
and U710 (N_710,In_510,In_413);
nand U711 (N_711,In_6,In_135);
nand U712 (N_712,In_343,In_648);
or U713 (N_713,In_81,In_463);
nand U714 (N_714,In_499,In_180);
and U715 (N_715,In_396,In_101);
nand U716 (N_716,In_110,In_127);
or U717 (N_717,In_91,In_196);
nand U718 (N_718,In_604,In_544);
nor U719 (N_719,In_301,In_387);
or U720 (N_720,In_106,In_277);
nor U721 (N_721,In_272,In_377);
nand U722 (N_722,In_344,In_127);
nor U723 (N_723,In_444,In_157);
nor U724 (N_724,In_558,In_504);
and U725 (N_725,In_19,In_324);
or U726 (N_726,In_103,In_23);
nand U727 (N_727,In_315,In_80);
nor U728 (N_728,In_422,In_373);
and U729 (N_729,In_592,In_573);
nor U730 (N_730,In_714,In_487);
nor U731 (N_731,In_219,In_731);
nand U732 (N_732,In_43,In_55);
xnor U733 (N_733,In_420,In_21);
nor U734 (N_734,In_346,In_635);
xor U735 (N_735,In_364,In_608);
nand U736 (N_736,In_658,In_681);
or U737 (N_737,In_555,In_432);
nand U738 (N_738,In_735,In_639);
or U739 (N_739,In_296,In_307);
nor U740 (N_740,In_263,In_192);
or U741 (N_741,In_558,In_388);
or U742 (N_742,In_156,In_175);
nand U743 (N_743,In_720,In_230);
nor U744 (N_744,In_300,In_575);
nand U745 (N_745,In_311,In_655);
nand U746 (N_746,In_297,In_466);
and U747 (N_747,In_708,In_66);
nand U748 (N_748,In_519,In_587);
and U749 (N_749,In_73,In_36);
and U750 (N_750,In_305,In_689);
or U751 (N_751,In_696,In_142);
nor U752 (N_752,In_70,In_396);
or U753 (N_753,In_365,In_552);
nand U754 (N_754,In_497,In_107);
nand U755 (N_755,In_173,In_422);
or U756 (N_756,In_603,In_472);
and U757 (N_757,In_420,In_604);
and U758 (N_758,In_192,In_1);
or U759 (N_759,In_658,In_443);
or U760 (N_760,In_132,In_469);
nand U761 (N_761,In_279,In_141);
or U762 (N_762,In_723,In_220);
nand U763 (N_763,In_305,In_605);
nor U764 (N_764,In_532,In_554);
nand U765 (N_765,In_261,In_674);
nand U766 (N_766,In_410,In_358);
nand U767 (N_767,In_142,In_73);
or U768 (N_768,In_186,In_175);
nor U769 (N_769,In_310,In_683);
and U770 (N_770,In_708,In_749);
and U771 (N_771,In_544,In_487);
and U772 (N_772,In_261,In_659);
nor U773 (N_773,In_253,In_327);
nor U774 (N_774,In_621,In_503);
nor U775 (N_775,In_169,In_595);
nor U776 (N_776,In_108,In_741);
and U777 (N_777,In_653,In_658);
nand U778 (N_778,In_283,In_471);
or U779 (N_779,In_680,In_149);
nand U780 (N_780,In_640,In_186);
nor U781 (N_781,In_358,In_72);
nand U782 (N_782,In_305,In_604);
nand U783 (N_783,In_660,In_91);
nand U784 (N_784,In_374,In_336);
nand U785 (N_785,In_234,In_161);
nor U786 (N_786,In_296,In_685);
nor U787 (N_787,In_521,In_501);
nand U788 (N_788,In_267,In_674);
nor U789 (N_789,In_373,In_652);
and U790 (N_790,In_458,In_20);
nand U791 (N_791,In_212,In_512);
and U792 (N_792,In_39,In_223);
and U793 (N_793,In_649,In_426);
nand U794 (N_794,In_400,In_724);
xnor U795 (N_795,In_316,In_81);
and U796 (N_796,In_185,In_263);
nand U797 (N_797,In_702,In_556);
and U798 (N_798,In_575,In_217);
and U799 (N_799,In_180,In_143);
nor U800 (N_800,In_124,In_375);
nor U801 (N_801,In_324,In_168);
nor U802 (N_802,In_360,In_516);
nor U803 (N_803,In_213,In_659);
and U804 (N_804,In_44,In_362);
and U805 (N_805,In_133,In_104);
nor U806 (N_806,In_405,In_71);
and U807 (N_807,In_466,In_143);
nor U808 (N_808,In_524,In_183);
nand U809 (N_809,In_14,In_442);
nand U810 (N_810,In_638,In_53);
and U811 (N_811,In_24,In_109);
nand U812 (N_812,In_487,In_606);
nand U813 (N_813,In_361,In_340);
and U814 (N_814,In_183,In_91);
or U815 (N_815,In_160,In_612);
and U816 (N_816,In_695,In_536);
and U817 (N_817,In_10,In_161);
nor U818 (N_818,In_242,In_92);
or U819 (N_819,In_102,In_214);
nor U820 (N_820,In_120,In_492);
nor U821 (N_821,In_642,In_71);
or U822 (N_822,In_63,In_103);
and U823 (N_823,In_320,In_387);
nand U824 (N_824,In_510,In_255);
and U825 (N_825,In_534,In_277);
nor U826 (N_826,In_177,In_223);
and U827 (N_827,In_719,In_82);
nand U828 (N_828,In_87,In_399);
nor U829 (N_829,In_282,In_62);
nand U830 (N_830,In_18,In_316);
nor U831 (N_831,In_305,In_323);
nand U832 (N_832,In_639,In_75);
and U833 (N_833,In_511,In_526);
or U834 (N_834,In_689,In_488);
nor U835 (N_835,In_338,In_649);
nand U836 (N_836,In_597,In_268);
nor U837 (N_837,In_169,In_332);
nor U838 (N_838,In_705,In_515);
nor U839 (N_839,In_563,In_258);
nand U840 (N_840,In_473,In_38);
and U841 (N_841,In_462,In_584);
xnor U842 (N_842,In_317,In_14);
and U843 (N_843,In_63,In_209);
nor U844 (N_844,In_702,In_565);
and U845 (N_845,In_189,In_488);
nor U846 (N_846,In_504,In_167);
xnor U847 (N_847,In_24,In_67);
nand U848 (N_848,In_579,In_237);
and U849 (N_849,In_515,In_629);
or U850 (N_850,In_85,In_39);
and U851 (N_851,In_178,In_258);
and U852 (N_852,In_127,In_285);
or U853 (N_853,In_665,In_532);
or U854 (N_854,In_643,In_453);
or U855 (N_855,In_85,In_709);
nand U856 (N_856,In_71,In_250);
or U857 (N_857,In_330,In_700);
and U858 (N_858,In_235,In_165);
nand U859 (N_859,In_445,In_573);
or U860 (N_860,In_738,In_657);
or U861 (N_861,In_506,In_629);
and U862 (N_862,In_386,In_52);
and U863 (N_863,In_137,In_36);
nand U864 (N_864,In_48,In_183);
nand U865 (N_865,In_446,In_66);
nand U866 (N_866,In_589,In_738);
or U867 (N_867,In_403,In_247);
xnor U868 (N_868,In_394,In_591);
and U869 (N_869,In_338,In_178);
or U870 (N_870,In_666,In_690);
or U871 (N_871,In_244,In_566);
nand U872 (N_872,In_592,In_525);
nor U873 (N_873,In_210,In_259);
nand U874 (N_874,In_739,In_310);
or U875 (N_875,In_35,In_407);
and U876 (N_876,In_512,In_660);
nand U877 (N_877,In_682,In_585);
nand U878 (N_878,In_94,In_460);
or U879 (N_879,In_311,In_258);
nor U880 (N_880,In_652,In_154);
or U881 (N_881,In_127,In_390);
nor U882 (N_882,In_271,In_100);
and U883 (N_883,In_410,In_519);
nand U884 (N_884,In_449,In_244);
and U885 (N_885,In_121,In_245);
and U886 (N_886,In_478,In_548);
nor U887 (N_887,In_74,In_30);
or U888 (N_888,In_134,In_276);
nor U889 (N_889,In_284,In_517);
or U890 (N_890,In_513,In_50);
nor U891 (N_891,In_690,In_44);
nor U892 (N_892,In_399,In_290);
and U893 (N_893,In_10,In_269);
nand U894 (N_894,In_326,In_50);
or U895 (N_895,In_616,In_81);
and U896 (N_896,In_331,In_728);
or U897 (N_897,In_167,In_289);
and U898 (N_898,In_351,In_627);
and U899 (N_899,In_67,In_119);
nand U900 (N_900,In_425,In_683);
or U901 (N_901,In_365,In_443);
nand U902 (N_902,In_315,In_452);
nand U903 (N_903,In_88,In_676);
and U904 (N_904,In_430,In_134);
nand U905 (N_905,In_59,In_83);
or U906 (N_906,In_240,In_742);
nor U907 (N_907,In_645,In_629);
nor U908 (N_908,In_124,In_212);
and U909 (N_909,In_640,In_343);
and U910 (N_910,In_489,In_682);
or U911 (N_911,In_108,In_132);
nor U912 (N_912,In_323,In_395);
nor U913 (N_913,In_315,In_344);
nand U914 (N_914,In_216,In_550);
or U915 (N_915,In_194,In_154);
or U916 (N_916,In_21,In_348);
and U917 (N_917,In_353,In_145);
and U918 (N_918,In_119,In_510);
nor U919 (N_919,In_29,In_58);
and U920 (N_920,In_611,In_130);
or U921 (N_921,In_254,In_747);
and U922 (N_922,In_493,In_698);
nor U923 (N_923,In_405,In_584);
nor U924 (N_924,In_323,In_345);
nand U925 (N_925,In_576,In_339);
nand U926 (N_926,In_740,In_524);
nand U927 (N_927,In_579,In_729);
and U928 (N_928,In_347,In_624);
nand U929 (N_929,In_394,In_614);
nand U930 (N_930,In_583,In_380);
nand U931 (N_931,In_85,In_332);
nand U932 (N_932,In_502,In_577);
xnor U933 (N_933,In_373,In_417);
and U934 (N_934,In_692,In_243);
nor U935 (N_935,In_625,In_610);
nor U936 (N_936,In_443,In_427);
nand U937 (N_937,In_703,In_67);
nand U938 (N_938,In_534,In_155);
nor U939 (N_939,In_588,In_554);
nand U940 (N_940,In_725,In_292);
or U941 (N_941,In_98,In_32);
or U942 (N_942,In_734,In_31);
and U943 (N_943,In_9,In_189);
nand U944 (N_944,In_721,In_661);
nor U945 (N_945,In_285,In_708);
nor U946 (N_946,In_191,In_37);
nand U947 (N_947,In_12,In_526);
nor U948 (N_948,In_283,In_64);
nor U949 (N_949,In_67,In_422);
nand U950 (N_950,In_693,In_2);
and U951 (N_951,In_676,In_139);
and U952 (N_952,In_135,In_203);
nor U953 (N_953,In_246,In_615);
nor U954 (N_954,In_27,In_630);
and U955 (N_955,In_488,In_224);
nand U956 (N_956,In_622,In_464);
nand U957 (N_957,In_126,In_553);
or U958 (N_958,In_87,In_397);
xnor U959 (N_959,In_747,In_201);
nor U960 (N_960,In_570,In_606);
nor U961 (N_961,In_115,In_148);
or U962 (N_962,In_240,In_305);
nor U963 (N_963,In_394,In_313);
nand U964 (N_964,In_96,In_34);
or U965 (N_965,In_206,In_651);
or U966 (N_966,In_82,In_255);
nand U967 (N_967,In_481,In_251);
nor U968 (N_968,In_656,In_160);
nor U969 (N_969,In_336,In_738);
or U970 (N_970,In_671,In_355);
xor U971 (N_971,In_59,In_666);
or U972 (N_972,In_471,In_105);
and U973 (N_973,In_132,In_706);
nor U974 (N_974,In_385,In_148);
and U975 (N_975,In_564,In_575);
nor U976 (N_976,In_225,In_33);
nor U977 (N_977,In_531,In_25);
nor U978 (N_978,In_108,In_560);
and U979 (N_979,In_509,In_448);
or U980 (N_980,In_206,In_638);
and U981 (N_981,In_550,In_393);
or U982 (N_982,In_720,In_173);
xnor U983 (N_983,In_541,In_290);
and U984 (N_984,In_490,In_335);
nor U985 (N_985,In_419,In_245);
or U986 (N_986,In_543,In_187);
nor U987 (N_987,In_393,In_482);
nand U988 (N_988,In_619,In_49);
nand U989 (N_989,In_60,In_236);
nand U990 (N_990,In_524,In_118);
and U991 (N_991,In_145,In_477);
nand U992 (N_992,In_221,In_552);
nand U993 (N_993,In_423,In_256);
nor U994 (N_994,In_552,In_649);
nand U995 (N_995,In_410,In_384);
and U996 (N_996,In_428,In_417);
nor U997 (N_997,In_514,In_192);
nor U998 (N_998,In_4,In_59);
and U999 (N_999,In_653,In_149);
nand U1000 (N_1000,In_113,In_691);
and U1001 (N_1001,In_136,In_452);
nor U1002 (N_1002,In_288,In_446);
nand U1003 (N_1003,In_181,In_304);
or U1004 (N_1004,In_118,In_132);
or U1005 (N_1005,In_461,In_160);
and U1006 (N_1006,In_408,In_597);
nand U1007 (N_1007,In_498,In_220);
nand U1008 (N_1008,In_270,In_379);
and U1009 (N_1009,In_17,In_355);
nor U1010 (N_1010,In_256,In_533);
nor U1011 (N_1011,In_743,In_110);
and U1012 (N_1012,In_429,In_102);
and U1013 (N_1013,In_394,In_384);
or U1014 (N_1014,In_379,In_127);
nand U1015 (N_1015,In_546,In_205);
nand U1016 (N_1016,In_684,In_58);
or U1017 (N_1017,In_527,In_172);
or U1018 (N_1018,In_119,In_734);
or U1019 (N_1019,In_74,In_670);
nor U1020 (N_1020,In_324,In_106);
nand U1021 (N_1021,In_488,In_289);
nand U1022 (N_1022,In_75,In_620);
and U1023 (N_1023,In_652,In_47);
and U1024 (N_1024,In_278,In_490);
or U1025 (N_1025,In_267,In_186);
nand U1026 (N_1026,In_391,In_420);
nand U1027 (N_1027,In_64,In_603);
and U1028 (N_1028,In_601,In_717);
nand U1029 (N_1029,In_681,In_707);
and U1030 (N_1030,In_528,In_69);
or U1031 (N_1031,In_389,In_412);
and U1032 (N_1032,In_493,In_672);
or U1033 (N_1033,In_211,In_297);
nor U1034 (N_1034,In_32,In_79);
and U1035 (N_1035,In_237,In_747);
nor U1036 (N_1036,In_411,In_305);
nand U1037 (N_1037,In_413,In_608);
nand U1038 (N_1038,In_472,In_42);
nand U1039 (N_1039,In_160,In_333);
nor U1040 (N_1040,In_267,In_637);
or U1041 (N_1041,In_119,In_498);
and U1042 (N_1042,In_82,In_420);
nand U1043 (N_1043,In_608,In_460);
nand U1044 (N_1044,In_540,In_545);
nand U1045 (N_1045,In_218,In_719);
xor U1046 (N_1046,In_430,In_364);
or U1047 (N_1047,In_659,In_670);
and U1048 (N_1048,In_556,In_703);
and U1049 (N_1049,In_639,In_643);
or U1050 (N_1050,In_292,In_662);
or U1051 (N_1051,In_13,In_388);
and U1052 (N_1052,In_52,In_428);
nand U1053 (N_1053,In_587,In_98);
nor U1054 (N_1054,In_710,In_124);
or U1055 (N_1055,In_657,In_693);
nand U1056 (N_1056,In_368,In_684);
nand U1057 (N_1057,In_274,In_240);
nand U1058 (N_1058,In_598,In_674);
and U1059 (N_1059,In_348,In_449);
or U1060 (N_1060,In_293,In_660);
and U1061 (N_1061,In_211,In_488);
nand U1062 (N_1062,In_87,In_143);
and U1063 (N_1063,In_63,In_323);
nor U1064 (N_1064,In_644,In_369);
nand U1065 (N_1065,In_570,In_509);
nor U1066 (N_1066,In_240,In_585);
and U1067 (N_1067,In_276,In_207);
nand U1068 (N_1068,In_289,In_466);
nand U1069 (N_1069,In_310,In_562);
and U1070 (N_1070,In_78,In_662);
nand U1071 (N_1071,In_77,In_721);
and U1072 (N_1072,In_242,In_372);
nor U1073 (N_1073,In_486,In_341);
xnor U1074 (N_1074,In_453,In_170);
and U1075 (N_1075,In_552,In_228);
nor U1076 (N_1076,In_443,In_346);
nand U1077 (N_1077,In_421,In_374);
or U1078 (N_1078,In_550,In_524);
and U1079 (N_1079,In_522,In_102);
and U1080 (N_1080,In_5,In_485);
and U1081 (N_1081,In_424,In_666);
and U1082 (N_1082,In_129,In_137);
nand U1083 (N_1083,In_580,In_213);
nor U1084 (N_1084,In_532,In_473);
or U1085 (N_1085,In_258,In_189);
or U1086 (N_1086,In_696,In_157);
and U1087 (N_1087,In_575,In_382);
or U1088 (N_1088,In_223,In_151);
nand U1089 (N_1089,In_640,In_546);
and U1090 (N_1090,In_540,In_214);
nor U1091 (N_1091,In_307,In_461);
nand U1092 (N_1092,In_197,In_195);
and U1093 (N_1093,In_698,In_403);
and U1094 (N_1094,In_305,In_591);
and U1095 (N_1095,In_228,In_331);
and U1096 (N_1096,In_660,In_659);
nor U1097 (N_1097,In_416,In_418);
or U1098 (N_1098,In_494,In_275);
nor U1099 (N_1099,In_385,In_642);
nand U1100 (N_1100,In_258,In_618);
nor U1101 (N_1101,In_191,In_129);
and U1102 (N_1102,In_332,In_561);
and U1103 (N_1103,In_308,In_155);
or U1104 (N_1104,In_718,In_285);
nand U1105 (N_1105,In_149,In_340);
and U1106 (N_1106,In_257,In_166);
xor U1107 (N_1107,In_23,In_242);
or U1108 (N_1108,In_742,In_173);
nand U1109 (N_1109,In_389,In_365);
nand U1110 (N_1110,In_71,In_332);
nand U1111 (N_1111,In_540,In_93);
or U1112 (N_1112,In_220,In_570);
or U1113 (N_1113,In_309,In_682);
or U1114 (N_1114,In_713,In_492);
nor U1115 (N_1115,In_636,In_733);
or U1116 (N_1116,In_45,In_11);
nor U1117 (N_1117,In_101,In_337);
nor U1118 (N_1118,In_539,In_204);
or U1119 (N_1119,In_370,In_270);
or U1120 (N_1120,In_342,In_544);
or U1121 (N_1121,In_404,In_731);
nand U1122 (N_1122,In_501,In_481);
nor U1123 (N_1123,In_659,In_212);
nor U1124 (N_1124,In_495,In_470);
nand U1125 (N_1125,In_242,In_531);
nor U1126 (N_1126,In_701,In_214);
and U1127 (N_1127,In_634,In_683);
and U1128 (N_1128,In_149,In_133);
or U1129 (N_1129,In_660,In_465);
and U1130 (N_1130,In_244,In_480);
nor U1131 (N_1131,In_366,In_528);
nand U1132 (N_1132,In_214,In_452);
nand U1133 (N_1133,In_65,In_742);
nor U1134 (N_1134,In_740,In_463);
or U1135 (N_1135,In_238,In_489);
or U1136 (N_1136,In_267,In_608);
and U1137 (N_1137,In_638,In_370);
and U1138 (N_1138,In_444,In_652);
and U1139 (N_1139,In_465,In_236);
nor U1140 (N_1140,In_230,In_548);
nor U1141 (N_1141,In_247,In_684);
and U1142 (N_1142,In_220,In_675);
nand U1143 (N_1143,In_209,In_357);
nand U1144 (N_1144,In_660,In_349);
xnor U1145 (N_1145,In_609,In_399);
nand U1146 (N_1146,In_249,In_368);
or U1147 (N_1147,In_510,In_652);
nand U1148 (N_1148,In_314,In_744);
and U1149 (N_1149,In_623,In_721);
and U1150 (N_1150,In_112,In_247);
nor U1151 (N_1151,In_90,In_672);
nor U1152 (N_1152,In_129,In_699);
nand U1153 (N_1153,In_733,In_132);
and U1154 (N_1154,In_645,In_116);
nand U1155 (N_1155,In_716,In_627);
and U1156 (N_1156,In_325,In_463);
nand U1157 (N_1157,In_320,In_516);
and U1158 (N_1158,In_18,In_390);
or U1159 (N_1159,In_639,In_133);
nor U1160 (N_1160,In_549,In_525);
nand U1161 (N_1161,In_29,In_554);
or U1162 (N_1162,In_414,In_652);
nor U1163 (N_1163,In_415,In_293);
and U1164 (N_1164,In_712,In_484);
or U1165 (N_1165,In_279,In_129);
nor U1166 (N_1166,In_707,In_400);
nor U1167 (N_1167,In_502,In_328);
nor U1168 (N_1168,In_585,In_48);
and U1169 (N_1169,In_123,In_577);
nor U1170 (N_1170,In_287,In_557);
nand U1171 (N_1171,In_274,In_290);
and U1172 (N_1172,In_415,In_67);
nand U1173 (N_1173,In_479,In_403);
nor U1174 (N_1174,In_511,In_0);
and U1175 (N_1175,In_236,In_205);
or U1176 (N_1176,In_566,In_731);
nor U1177 (N_1177,In_745,In_89);
nand U1178 (N_1178,In_661,In_390);
or U1179 (N_1179,In_475,In_511);
nor U1180 (N_1180,In_500,In_600);
nor U1181 (N_1181,In_351,In_691);
or U1182 (N_1182,In_86,In_204);
and U1183 (N_1183,In_623,In_350);
nor U1184 (N_1184,In_655,In_16);
nor U1185 (N_1185,In_179,In_682);
nand U1186 (N_1186,In_581,In_52);
nand U1187 (N_1187,In_19,In_667);
nor U1188 (N_1188,In_333,In_372);
and U1189 (N_1189,In_108,In_424);
nand U1190 (N_1190,In_463,In_681);
and U1191 (N_1191,In_154,In_553);
nand U1192 (N_1192,In_324,In_420);
nor U1193 (N_1193,In_539,In_118);
nand U1194 (N_1194,In_637,In_581);
nand U1195 (N_1195,In_625,In_156);
and U1196 (N_1196,In_196,In_435);
nand U1197 (N_1197,In_470,In_90);
or U1198 (N_1198,In_396,In_113);
or U1199 (N_1199,In_120,In_554);
nand U1200 (N_1200,In_129,In_617);
and U1201 (N_1201,In_527,In_272);
nor U1202 (N_1202,In_356,In_278);
nor U1203 (N_1203,In_562,In_663);
nand U1204 (N_1204,In_126,In_595);
or U1205 (N_1205,In_120,In_586);
nor U1206 (N_1206,In_24,In_375);
or U1207 (N_1207,In_717,In_339);
and U1208 (N_1208,In_402,In_532);
nand U1209 (N_1209,In_727,In_381);
nor U1210 (N_1210,In_310,In_163);
or U1211 (N_1211,In_58,In_540);
nand U1212 (N_1212,In_681,In_573);
xor U1213 (N_1213,In_663,In_719);
nand U1214 (N_1214,In_116,In_140);
or U1215 (N_1215,In_302,In_149);
or U1216 (N_1216,In_25,In_261);
nand U1217 (N_1217,In_281,In_187);
and U1218 (N_1218,In_631,In_713);
nor U1219 (N_1219,In_435,In_489);
nor U1220 (N_1220,In_644,In_405);
or U1221 (N_1221,In_344,In_115);
nor U1222 (N_1222,In_466,In_379);
nor U1223 (N_1223,In_250,In_712);
nand U1224 (N_1224,In_620,In_321);
nor U1225 (N_1225,In_37,In_46);
nor U1226 (N_1226,In_326,In_472);
and U1227 (N_1227,In_62,In_335);
or U1228 (N_1228,In_704,In_546);
nor U1229 (N_1229,In_603,In_659);
nand U1230 (N_1230,In_9,In_254);
nand U1231 (N_1231,In_132,In_310);
nor U1232 (N_1232,In_194,In_369);
nand U1233 (N_1233,In_726,In_157);
nor U1234 (N_1234,In_144,In_316);
nand U1235 (N_1235,In_377,In_525);
nand U1236 (N_1236,In_321,In_730);
nand U1237 (N_1237,In_91,In_156);
nor U1238 (N_1238,In_115,In_159);
nor U1239 (N_1239,In_598,In_491);
and U1240 (N_1240,In_326,In_624);
and U1241 (N_1241,In_167,In_442);
or U1242 (N_1242,In_52,In_448);
nand U1243 (N_1243,In_717,In_221);
nand U1244 (N_1244,In_277,In_659);
and U1245 (N_1245,In_186,In_366);
and U1246 (N_1246,In_472,In_236);
and U1247 (N_1247,In_681,In_715);
nor U1248 (N_1248,In_716,In_745);
or U1249 (N_1249,In_267,In_202);
nor U1250 (N_1250,In_299,In_557);
nor U1251 (N_1251,In_476,In_263);
nand U1252 (N_1252,In_291,In_156);
nand U1253 (N_1253,In_731,In_708);
nor U1254 (N_1254,In_282,In_137);
nor U1255 (N_1255,In_502,In_446);
nor U1256 (N_1256,In_73,In_422);
nand U1257 (N_1257,In_64,In_400);
or U1258 (N_1258,In_601,In_113);
and U1259 (N_1259,In_201,In_118);
or U1260 (N_1260,In_341,In_38);
or U1261 (N_1261,In_257,In_707);
and U1262 (N_1262,In_128,In_203);
nand U1263 (N_1263,In_692,In_738);
or U1264 (N_1264,In_372,In_49);
and U1265 (N_1265,In_77,In_302);
or U1266 (N_1266,In_643,In_467);
xnor U1267 (N_1267,In_667,In_141);
or U1268 (N_1268,In_341,In_406);
xor U1269 (N_1269,In_574,In_537);
nand U1270 (N_1270,In_298,In_391);
nand U1271 (N_1271,In_487,In_252);
nor U1272 (N_1272,In_400,In_112);
nand U1273 (N_1273,In_329,In_181);
or U1274 (N_1274,In_350,In_608);
nor U1275 (N_1275,In_77,In_666);
nand U1276 (N_1276,In_627,In_203);
or U1277 (N_1277,In_445,In_636);
and U1278 (N_1278,In_510,In_333);
or U1279 (N_1279,In_180,In_171);
xnor U1280 (N_1280,In_733,In_393);
or U1281 (N_1281,In_470,In_131);
xnor U1282 (N_1282,In_720,In_2);
nand U1283 (N_1283,In_652,In_561);
xor U1284 (N_1284,In_625,In_246);
and U1285 (N_1285,In_511,In_142);
and U1286 (N_1286,In_621,In_213);
and U1287 (N_1287,In_42,In_545);
xor U1288 (N_1288,In_47,In_327);
nand U1289 (N_1289,In_565,In_524);
or U1290 (N_1290,In_561,In_87);
or U1291 (N_1291,In_284,In_368);
nor U1292 (N_1292,In_112,In_138);
and U1293 (N_1293,In_732,In_82);
nand U1294 (N_1294,In_331,In_285);
or U1295 (N_1295,In_743,In_543);
and U1296 (N_1296,In_117,In_156);
and U1297 (N_1297,In_622,In_678);
nand U1298 (N_1298,In_284,In_559);
nor U1299 (N_1299,In_36,In_701);
or U1300 (N_1300,In_200,In_666);
nor U1301 (N_1301,In_84,In_391);
and U1302 (N_1302,In_471,In_167);
and U1303 (N_1303,In_413,In_211);
and U1304 (N_1304,In_509,In_138);
and U1305 (N_1305,In_292,In_510);
nor U1306 (N_1306,In_680,In_744);
and U1307 (N_1307,In_427,In_294);
and U1308 (N_1308,In_223,In_410);
and U1309 (N_1309,In_314,In_578);
nor U1310 (N_1310,In_485,In_61);
or U1311 (N_1311,In_481,In_240);
nand U1312 (N_1312,In_396,In_636);
nand U1313 (N_1313,In_333,In_173);
nor U1314 (N_1314,In_165,In_140);
nor U1315 (N_1315,In_12,In_427);
nand U1316 (N_1316,In_278,In_5);
nand U1317 (N_1317,In_333,In_503);
or U1318 (N_1318,In_197,In_339);
nand U1319 (N_1319,In_494,In_370);
nand U1320 (N_1320,In_247,In_55);
and U1321 (N_1321,In_56,In_278);
nor U1322 (N_1322,In_304,In_50);
nor U1323 (N_1323,In_242,In_379);
nand U1324 (N_1324,In_12,In_196);
or U1325 (N_1325,In_351,In_102);
or U1326 (N_1326,In_461,In_77);
or U1327 (N_1327,In_463,In_495);
nand U1328 (N_1328,In_104,In_140);
nor U1329 (N_1329,In_420,In_343);
nor U1330 (N_1330,In_242,In_533);
nor U1331 (N_1331,In_691,In_354);
or U1332 (N_1332,In_538,In_392);
nand U1333 (N_1333,In_634,In_661);
and U1334 (N_1334,In_48,In_371);
nand U1335 (N_1335,In_590,In_591);
nand U1336 (N_1336,In_511,In_636);
nand U1337 (N_1337,In_107,In_67);
and U1338 (N_1338,In_221,In_326);
and U1339 (N_1339,In_167,In_4);
or U1340 (N_1340,In_16,In_208);
or U1341 (N_1341,In_668,In_418);
or U1342 (N_1342,In_103,In_247);
or U1343 (N_1343,In_113,In_156);
and U1344 (N_1344,In_686,In_296);
and U1345 (N_1345,In_19,In_680);
nand U1346 (N_1346,In_43,In_668);
or U1347 (N_1347,In_60,In_196);
nand U1348 (N_1348,In_440,In_746);
or U1349 (N_1349,In_743,In_319);
and U1350 (N_1350,In_731,In_341);
and U1351 (N_1351,In_584,In_661);
nand U1352 (N_1352,In_604,In_26);
nor U1353 (N_1353,In_68,In_435);
nor U1354 (N_1354,In_568,In_150);
nand U1355 (N_1355,In_469,In_383);
and U1356 (N_1356,In_578,In_100);
and U1357 (N_1357,In_79,In_551);
nor U1358 (N_1358,In_460,In_36);
nand U1359 (N_1359,In_590,In_657);
and U1360 (N_1360,In_533,In_743);
or U1361 (N_1361,In_498,In_461);
nand U1362 (N_1362,In_454,In_518);
and U1363 (N_1363,In_333,In_537);
or U1364 (N_1364,In_310,In_113);
or U1365 (N_1365,In_432,In_252);
nor U1366 (N_1366,In_366,In_76);
nor U1367 (N_1367,In_350,In_194);
nand U1368 (N_1368,In_532,In_7);
nor U1369 (N_1369,In_696,In_636);
nor U1370 (N_1370,In_617,In_412);
nand U1371 (N_1371,In_625,In_385);
or U1372 (N_1372,In_89,In_522);
or U1373 (N_1373,In_285,In_320);
or U1374 (N_1374,In_140,In_540);
or U1375 (N_1375,In_577,In_145);
nand U1376 (N_1376,In_405,In_556);
or U1377 (N_1377,In_102,In_118);
or U1378 (N_1378,In_548,In_545);
and U1379 (N_1379,In_55,In_123);
or U1380 (N_1380,In_427,In_272);
and U1381 (N_1381,In_494,In_130);
nor U1382 (N_1382,In_212,In_191);
and U1383 (N_1383,In_194,In_635);
nor U1384 (N_1384,In_297,In_572);
and U1385 (N_1385,In_420,In_666);
nor U1386 (N_1386,In_422,In_563);
nand U1387 (N_1387,In_386,In_317);
nor U1388 (N_1388,In_7,In_443);
and U1389 (N_1389,In_730,In_141);
and U1390 (N_1390,In_14,In_547);
nor U1391 (N_1391,In_167,In_259);
and U1392 (N_1392,In_93,In_257);
nand U1393 (N_1393,In_485,In_104);
nor U1394 (N_1394,In_118,In_473);
and U1395 (N_1395,In_382,In_238);
nand U1396 (N_1396,In_728,In_711);
and U1397 (N_1397,In_93,In_414);
nor U1398 (N_1398,In_583,In_16);
nand U1399 (N_1399,In_125,In_440);
and U1400 (N_1400,In_140,In_185);
nor U1401 (N_1401,In_72,In_166);
and U1402 (N_1402,In_606,In_236);
nand U1403 (N_1403,In_376,In_175);
nand U1404 (N_1404,In_198,In_0);
and U1405 (N_1405,In_623,In_29);
and U1406 (N_1406,In_184,In_90);
nand U1407 (N_1407,In_139,In_357);
and U1408 (N_1408,In_430,In_629);
or U1409 (N_1409,In_135,In_298);
nand U1410 (N_1410,In_540,In_698);
or U1411 (N_1411,In_600,In_378);
nor U1412 (N_1412,In_63,In_314);
and U1413 (N_1413,In_471,In_198);
and U1414 (N_1414,In_283,In_639);
nand U1415 (N_1415,In_594,In_210);
nor U1416 (N_1416,In_617,In_61);
nor U1417 (N_1417,In_77,In_560);
nor U1418 (N_1418,In_301,In_123);
and U1419 (N_1419,In_713,In_107);
nor U1420 (N_1420,In_438,In_514);
xor U1421 (N_1421,In_407,In_280);
or U1422 (N_1422,In_686,In_238);
or U1423 (N_1423,In_743,In_174);
and U1424 (N_1424,In_260,In_391);
or U1425 (N_1425,In_704,In_134);
or U1426 (N_1426,In_382,In_475);
or U1427 (N_1427,In_45,In_503);
and U1428 (N_1428,In_582,In_17);
and U1429 (N_1429,In_454,In_242);
nand U1430 (N_1430,In_310,In_491);
and U1431 (N_1431,In_354,In_524);
xnor U1432 (N_1432,In_122,In_663);
or U1433 (N_1433,In_496,In_745);
and U1434 (N_1434,In_705,In_73);
and U1435 (N_1435,In_256,In_570);
nand U1436 (N_1436,In_575,In_482);
nor U1437 (N_1437,In_640,In_75);
and U1438 (N_1438,In_435,In_256);
nor U1439 (N_1439,In_115,In_243);
and U1440 (N_1440,In_10,In_434);
and U1441 (N_1441,In_346,In_272);
nor U1442 (N_1442,In_4,In_600);
and U1443 (N_1443,In_673,In_191);
nand U1444 (N_1444,In_726,In_96);
nor U1445 (N_1445,In_337,In_197);
nor U1446 (N_1446,In_737,In_334);
nand U1447 (N_1447,In_641,In_175);
nor U1448 (N_1448,In_407,In_356);
or U1449 (N_1449,In_660,In_217);
and U1450 (N_1450,In_321,In_268);
nand U1451 (N_1451,In_195,In_567);
nor U1452 (N_1452,In_14,In_192);
nand U1453 (N_1453,In_27,In_540);
nor U1454 (N_1454,In_567,In_149);
and U1455 (N_1455,In_657,In_37);
or U1456 (N_1456,In_391,In_445);
nor U1457 (N_1457,In_205,In_508);
and U1458 (N_1458,In_579,In_131);
nor U1459 (N_1459,In_296,In_279);
and U1460 (N_1460,In_306,In_488);
or U1461 (N_1461,In_749,In_314);
or U1462 (N_1462,In_738,In_24);
or U1463 (N_1463,In_310,In_342);
or U1464 (N_1464,In_487,In_341);
or U1465 (N_1465,In_312,In_718);
and U1466 (N_1466,In_241,In_466);
or U1467 (N_1467,In_291,In_96);
nor U1468 (N_1468,In_36,In_226);
and U1469 (N_1469,In_626,In_352);
nand U1470 (N_1470,In_164,In_272);
nor U1471 (N_1471,In_723,In_389);
and U1472 (N_1472,In_452,In_425);
nor U1473 (N_1473,In_639,In_74);
nor U1474 (N_1474,In_523,In_462);
or U1475 (N_1475,In_496,In_463);
or U1476 (N_1476,In_441,In_13);
or U1477 (N_1477,In_25,In_585);
nor U1478 (N_1478,In_647,In_129);
nand U1479 (N_1479,In_732,In_402);
or U1480 (N_1480,In_177,In_102);
nand U1481 (N_1481,In_715,In_353);
or U1482 (N_1482,In_695,In_313);
nand U1483 (N_1483,In_567,In_694);
nand U1484 (N_1484,In_700,In_476);
nand U1485 (N_1485,In_624,In_697);
nor U1486 (N_1486,In_475,In_150);
and U1487 (N_1487,In_379,In_677);
nor U1488 (N_1488,In_189,In_422);
and U1489 (N_1489,In_170,In_21);
nand U1490 (N_1490,In_51,In_691);
nand U1491 (N_1491,In_553,In_614);
and U1492 (N_1492,In_242,In_695);
or U1493 (N_1493,In_159,In_107);
or U1494 (N_1494,In_163,In_253);
and U1495 (N_1495,In_112,In_615);
or U1496 (N_1496,In_467,In_346);
or U1497 (N_1497,In_519,In_584);
nand U1498 (N_1498,In_429,In_311);
or U1499 (N_1499,In_596,In_119);
or U1500 (N_1500,In_679,In_554);
or U1501 (N_1501,In_277,In_570);
nor U1502 (N_1502,In_575,In_39);
and U1503 (N_1503,In_143,In_579);
nand U1504 (N_1504,In_704,In_54);
and U1505 (N_1505,In_23,In_428);
nor U1506 (N_1506,In_537,In_655);
and U1507 (N_1507,In_218,In_321);
and U1508 (N_1508,In_703,In_682);
nand U1509 (N_1509,In_230,In_418);
and U1510 (N_1510,In_222,In_26);
and U1511 (N_1511,In_262,In_112);
or U1512 (N_1512,In_209,In_313);
nor U1513 (N_1513,In_333,In_433);
and U1514 (N_1514,In_631,In_88);
or U1515 (N_1515,In_12,In_304);
xnor U1516 (N_1516,In_429,In_196);
xnor U1517 (N_1517,In_408,In_395);
or U1518 (N_1518,In_246,In_255);
nand U1519 (N_1519,In_708,In_380);
or U1520 (N_1520,In_145,In_31);
or U1521 (N_1521,In_355,In_54);
and U1522 (N_1522,In_727,In_658);
or U1523 (N_1523,In_435,In_156);
and U1524 (N_1524,In_467,In_321);
nor U1525 (N_1525,In_36,In_428);
or U1526 (N_1526,In_506,In_94);
or U1527 (N_1527,In_626,In_230);
nor U1528 (N_1528,In_377,In_207);
or U1529 (N_1529,In_159,In_79);
nor U1530 (N_1530,In_39,In_377);
or U1531 (N_1531,In_265,In_748);
nand U1532 (N_1532,In_178,In_635);
nor U1533 (N_1533,In_112,In_527);
and U1534 (N_1534,In_7,In_304);
nand U1535 (N_1535,In_692,In_482);
nand U1536 (N_1536,In_398,In_184);
nor U1537 (N_1537,In_707,In_560);
nand U1538 (N_1538,In_150,In_218);
and U1539 (N_1539,In_26,In_404);
or U1540 (N_1540,In_354,In_579);
or U1541 (N_1541,In_273,In_509);
and U1542 (N_1542,In_564,In_164);
nand U1543 (N_1543,In_642,In_140);
or U1544 (N_1544,In_505,In_389);
xnor U1545 (N_1545,In_258,In_333);
nor U1546 (N_1546,In_168,In_665);
and U1547 (N_1547,In_467,In_687);
and U1548 (N_1548,In_282,In_458);
or U1549 (N_1549,In_466,In_1);
nor U1550 (N_1550,In_587,In_120);
and U1551 (N_1551,In_484,In_10);
and U1552 (N_1552,In_189,In_465);
nand U1553 (N_1553,In_606,In_539);
and U1554 (N_1554,In_314,In_576);
and U1555 (N_1555,In_249,In_430);
nand U1556 (N_1556,In_452,In_523);
or U1557 (N_1557,In_264,In_15);
or U1558 (N_1558,In_684,In_388);
nand U1559 (N_1559,In_624,In_553);
xor U1560 (N_1560,In_519,In_671);
and U1561 (N_1561,In_424,In_61);
nor U1562 (N_1562,In_223,In_499);
nor U1563 (N_1563,In_477,In_673);
and U1564 (N_1564,In_383,In_741);
xnor U1565 (N_1565,In_102,In_658);
or U1566 (N_1566,In_108,In_111);
nand U1567 (N_1567,In_428,In_478);
and U1568 (N_1568,In_600,In_323);
or U1569 (N_1569,In_53,In_38);
and U1570 (N_1570,In_57,In_174);
or U1571 (N_1571,In_292,In_227);
nand U1572 (N_1572,In_530,In_99);
or U1573 (N_1573,In_366,In_493);
and U1574 (N_1574,In_574,In_690);
nand U1575 (N_1575,In_434,In_210);
or U1576 (N_1576,In_219,In_399);
xnor U1577 (N_1577,In_72,In_335);
xnor U1578 (N_1578,In_397,In_540);
and U1579 (N_1579,In_354,In_526);
and U1580 (N_1580,In_523,In_266);
nand U1581 (N_1581,In_653,In_742);
and U1582 (N_1582,In_397,In_251);
or U1583 (N_1583,In_270,In_675);
or U1584 (N_1584,In_295,In_223);
xnor U1585 (N_1585,In_704,In_655);
xnor U1586 (N_1586,In_331,In_486);
nand U1587 (N_1587,In_238,In_172);
nor U1588 (N_1588,In_192,In_308);
and U1589 (N_1589,In_472,In_556);
nor U1590 (N_1590,In_188,In_356);
and U1591 (N_1591,In_392,In_501);
or U1592 (N_1592,In_404,In_613);
and U1593 (N_1593,In_245,In_628);
and U1594 (N_1594,In_631,In_421);
or U1595 (N_1595,In_424,In_390);
nor U1596 (N_1596,In_672,In_288);
nand U1597 (N_1597,In_382,In_144);
nand U1598 (N_1598,In_91,In_367);
or U1599 (N_1599,In_337,In_90);
and U1600 (N_1600,In_293,In_641);
and U1601 (N_1601,In_622,In_653);
nor U1602 (N_1602,In_717,In_566);
xnor U1603 (N_1603,In_684,In_298);
xor U1604 (N_1604,In_202,In_57);
nand U1605 (N_1605,In_249,In_620);
and U1606 (N_1606,In_9,In_404);
nor U1607 (N_1607,In_739,In_682);
or U1608 (N_1608,In_489,In_161);
nand U1609 (N_1609,In_580,In_151);
nor U1610 (N_1610,In_298,In_81);
nand U1611 (N_1611,In_38,In_32);
nor U1612 (N_1612,In_521,In_571);
and U1613 (N_1613,In_691,In_736);
nand U1614 (N_1614,In_194,In_405);
nor U1615 (N_1615,In_426,In_340);
nand U1616 (N_1616,In_625,In_465);
and U1617 (N_1617,In_312,In_85);
xnor U1618 (N_1618,In_412,In_294);
nor U1619 (N_1619,In_33,In_129);
and U1620 (N_1620,In_47,In_373);
nand U1621 (N_1621,In_244,In_53);
nand U1622 (N_1622,In_338,In_18);
nand U1623 (N_1623,In_735,In_149);
xor U1624 (N_1624,In_32,In_679);
nor U1625 (N_1625,In_486,In_386);
or U1626 (N_1626,In_183,In_289);
and U1627 (N_1627,In_213,In_601);
nor U1628 (N_1628,In_577,In_85);
or U1629 (N_1629,In_27,In_244);
or U1630 (N_1630,In_400,In_63);
and U1631 (N_1631,In_317,In_740);
nor U1632 (N_1632,In_314,In_79);
or U1633 (N_1633,In_244,In_747);
nor U1634 (N_1634,In_608,In_380);
or U1635 (N_1635,In_558,In_335);
nor U1636 (N_1636,In_122,In_372);
nor U1637 (N_1637,In_459,In_273);
nor U1638 (N_1638,In_741,In_372);
or U1639 (N_1639,In_662,In_590);
and U1640 (N_1640,In_611,In_680);
nand U1641 (N_1641,In_501,In_146);
nor U1642 (N_1642,In_545,In_393);
or U1643 (N_1643,In_506,In_652);
or U1644 (N_1644,In_196,In_590);
nand U1645 (N_1645,In_543,In_325);
and U1646 (N_1646,In_4,In_345);
and U1647 (N_1647,In_509,In_276);
nand U1648 (N_1648,In_237,In_146);
nor U1649 (N_1649,In_54,In_475);
or U1650 (N_1650,In_202,In_622);
or U1651 (N_1651,In_301,In_408);
nand U1652 (N_1652,In_113,In_465);
and U1653 (N_1653,In_690,In_673);
and U1654 (N_1654,In_650,In_642);
or U1655 (N_1655,In_640,In_340);
or U1656 (N_1656,In_464,In_391);
or U1657 (N_1657,In_472,In_158);
nor U1658 (N_1658,In_582,In_396);
or U1659 (N_1659,In_25,In_499);
or U1660 (N_1660,In_613,In_122);
and U1661 (N_1661,In_121,In_552);
or U1662 (N_1662,In_78,In_225);
and U1663 (N_1663,In_166,In_366);
or U1664 (N_1664,In_187,In_362);
nand U1665 (N_1665,In_554,In_380);
nand U1666 (N_1666,In_488,In_347);
nand U1667 (N_1667,In_446,In_465);
nor U1668 (N_1668,In_711,In_693);
nor U1669 (N_1669,In_488,In_428);
and U1670 (N_1670,In_547,In_215);
nand U1671 (N_1671,In_196,In_179);
or U1672 (N_1672,In_712,In_573);
and U1673 (N_1673,In_236,In_723);
nand U1674 (N_1674,In_414,In_51);
xor U1675 (N_1675,In_645,In_467);
or U1676 (N_1676,In_136,In_412);
nor U1677 (N_1677,In_525,In_414);
and U1678 (N_1678,In_430,In_0);
and U1679 (N_1679,In_351,In_118);
nand U1680 (N_1680,In_377,In_575);
and U1681 (N_1681,In_342,In_285);
nand U1682 (N_1682,In_428,In_249);
nand U1683 (N_1683,In_748,In_634);
and U1684 (N_1684,In_318,In_484);
nor U1685 (N_1685,In_309,In_546);
nor U1686 (N_1686,In_294,In_118);
xor U1687 (N_1687,In_397,In_560);
nor U1688 (N_1688,In_36,In_746);
and U1689 (N_1689,In_301,In_599);
nor U1690 (N_1690,In_688,In_18);
nor U1691 (N_1691,In_556,In_522);
nand U1692 (N_1692,In_250,In_561);
and U1693 (N_1693,In_354,In_307);
and U1694 (N_1694,In_401,In_738);
nand U1695 (N_1695,In_281,In_483);
nor U1696 (N_1696,In_548,In_415);
nor U1697 (N_1697,In_648,In_309);
nor U1698 (N_1698,In_431,In_747);
and U1699 (N_1699,In_530,In_243);
and U1700 (N_1700,In_122,In_179);
nor U1701 (N_1701,In_321,In_483);
xnor U1702 (N_1702,In_607,In_304);
nor U1703 (N_1703,In_691,In_155);
nand U1704 (N_1704,In_56,In_166);
nand U1705 (N_1705,In_590,In_745);
or U1706 (N_1706,In_320,In_31);
nand U1707 (N_1707,In_270,In_491);
and U1708 (N_1708,In_509,In_381);
or U1709 (N_1709,In_340,In_543);
nand U1710 (N_1710,In_111,In_9);
or U1711 (N_1711,In_677,In_748);
nand U1712 (N_1712,In_624,In_221);
and U1713 (N_1713,In_649,In_479);
nor U1714 (N_1714,In_736,In_638);
or U1715 (N_1715,In_22,In_56);
nor U1716 (N_1716,In_617,In_237);
nand U1717 (N_1717,In_553,In_524);
or U1718 (N_1718,In_675,In_138);
and U1719 (N_1719,In_472,In_71);
or U1720 (N_1720,In_172,In_4);
and U1721 (N_1721,In_79,In_30);
nor U1722 (N_1722,In_382,In_316);
nor U1723 (N_1723,In_152,In_651);
nor U1724 (N_1724,In_277,In_725);
or U1725 (N_1725,In_174,In_553);
xor U1726 (N_1726,In_399,In_618);
nand U1727 (N_1727,In_141,In_354);
and U1728 (N_1728,In_37,In_274);
and U1729 (N_1729,In_289,In_177);
and U1730 (N_1730,In_542,In_3);
or U1731 (N_1731,In_342,In_353);
nor U1732 (N_1732,In_660,In_377);
nor U1733 (N_1733,In_210,In_589);
nand U1734 (N_1734,In_140,In_42);
nor U1735 (N_1735,In_418,In_550);
nand U1736 (N_1736,In_665,In_346);
nor U1737 (N_1737,In_372,In_600);
nand U1738 (N_1738,In_436,In_321);
nand U1739 (N_1739,In_167,In_72);
or U1740 (N_1740,In_52,In_22);
nor U1741 (N_1741,In_267,In_623);
or U1742 (N_1742,In_630,In_467);
or U1743 (N_1743,In_514,In_575);
xnor U1744 (N_1744,In_680,In_369);
xor U1745 (N_1745,In_31,In_341);
or U1746 (N_1746,In_94,In_678);
nand U1747 (N_1747,In_720,In_607);
nor U1748 (N_1748,In_98,In_127);
or U1749 (N_1749,In_600,In_47);
and U1750 (N_1750,In_506,In_132);
or U1751 (N_1751,In_557,In_9);
or U1752 (N_1752,In_380,In_242);
or U1753 (N_1753,In_476,In_169);
and U1754 (N_1754,In_701,In_700);
or U1755 (N_1755,In_251,In_503);
and U1756 (N_1756,In_680,In_208);
nand U1757 (N_1757,In_272,In_10);
nor U1758 (N_1758,In_87,In_353);
nand U1759 (N_1759,In_50,In_592);
nor U1760 (N_1760,In_493,In_741);
nand U1761 (N_1761,In_397,In_46);
nor U1762 (N_1762,In_420,In_102);
nor U1763 (N_1763,In_501,In_78);
and U1764 (N_1764,In_231,In_38);
or U1765 (N_1765,In_677,In_107);
or U1766 (N_1766,In_697,In_484);
nand U1767 (N_1767,In_547,In_466);
and U1768 (N_1768,In_717,In_451);
and U1769 (N_1769,In_62,In_508);
nand U1770 (N_1770,In_240,In_296);
and U1771 (N_1771,In_468,In_611);
or U1772 (N_1772,In_572,In_226);
or U1773 (N_1773,In_413,In_748);
and U1774 (N_1774,In_173,In_485);
nand U1775 (N_1775,In_271,In_498);
xor U1776 (N_1776,In_309,In_579);
nand U1777 (N_1777,In_473,In_524);
nand U1778 (N_1778,In_230,In_710);
and U1779 (N_1779,In_105,In_238);
and U1780 (N_1780,In_484,In_356);
nand U1781 (N_1781,In_439,In_387);
and U1782 (N_1782,In_476,In_434);
nand U1783 (N_1783,In_91,In_672);
nor U1784 (N_1784,In_527,In_635);
nand U1785 (N_1785,In_306,In_662);
or U1786 (N_1786,In_157,In_52);
nand U1787 (N_1787,In_133,In_181);
and U1788 (N_1788,In_69,In_13);
nand U1789 (N_1789,In_587,In_406);
or U1790 (N_1790,In_106,In_418);
nor U1791 (N_1791,In_373,In_22);
or U1792 (N_1792,In_451,In_368);
nand U1793 (N_1793,In_135,In_747);
and U1794 (N_1794,In_264,In_682);
and U1795 (N_1795,In_224,In_101);
nand U1796 (N_1796,In_287,In_383);
nand U1797 (N_1797,In_422,In_181);
and U1798 (N_1798,In_684,In_236);
nand U1799 (N_1799,In_416,In_12);
or U1800 (N_1800,In_473,In_474);
nand U1801 (N_1801,In_438,In_569);
and U1802 (N_1802,In_302,In_86);
nand U1803 (N_1803,In_622,In_674);
or U1804 (N_1804,In_606,In_4);
and U1805 (N_1805,In_449,In_53);
nand U1806 (N_1806,In_202,In_593);
nor U1807 (N_1807,In_318,In_617);
or U1808 (N_1808,In_588,In_375);
nand U1809 (N_1809,In_475,In_503);
nand U1810 (N_1810,In_131,In_576);
nor U1811 (N_1811,In_619,In_658);
nor U1812 (N_1812,In_34,In_699);
nor U1813 (N_1813,In_674,In_150);
nor U1814 (N_1814,In_263,In_194);
nor U1815 (N_1815,In_650,In_201);
or U1816 (N_1816,In_485,In_694);
or U1817 (N_1817,In_717,In_681);
or U1818 (N_1818,In_104,In_103);
and U1819 (N_1819,In_497,In_699);
or U1820 (N_1820,In_495,In_363);
nand U1821 (N_1821,In_635,In_39);
nor U1822 (N_1822,In_251,In_710);
or U1823 (N_1823,In_659,In_101);
nand U1824 (N_1824,In_634,In_321);
and U1825 (N_1825,In_418,In_225);
nor U1826 (N_1826,In_150,In_212);
nand U1827 (N_1827,In_3,In_447);
xor U1828 (N_1828,In_242,In_21);
nor U1829 (N_1829,In_723,In_257);
nand U1830 (N_1830,In_215,In_250);
and U1831 (N_1831,In_273,In_114);
nor U1832 (N_1832,In_354,In_505);
and U1833 (N_1833,In_459,In_146);
or U1834 (N_1834,In_138,In_320);
or U1835 (N_1835,In_724,In_148);
and U1836 (N_1836,In_341,In_464);
or U1837 (N_1837,In_6,In_279);
nand U1838 (N_1838,In_280,In_321);
nand U1839 (N_1839,In_132,In_570);
and U1840 (N_1840,In_199,In_574);
or U1841 (N_1841,In_270,In_614);
nor U1842 (N_1842,In_282,In_634);
nand U1843 (N_1843,In_281,In_396);
nor U1844 (N_1844,In_193,In_563);
nand U1845 (N_1845,In_228,In_440);
or U1846 (N_1846,In_406,In_678);
nor U1847 (N_1847,In_188,In_223);
and U1848 (N_1848,In_10,In_403);
nor U1849 (N_1849,In_18,In_410);
nor U1850 (N_1850,In_106,In_471);
nand U1851 (N_1851,In_135,In_743);
nand U1852 (N_1852,In_293,In_342);
nor U1853 (N_1853,In_511,In_516);
and U1854 (N_1854,In_715,In_392);
nand U1855 (N_1855,In_396,In_493);
or U1856 (N_1856,In_599,In_672);
or U1857 (N_1857,In_573,In_390);
or U1858 (N_1858,In_205,In_660);
xor U1859 (N_1859,In_354,In_125);
or U1860 (N_1860,In_7,In_63);
and U1861 (N_1861,In_35,In_620);
nand U1862 (N_1862,In_421,In_376);
or U1863 (N_1863,In_629,In_449);
or U1864 (N_1864,In_381,In_474);
nand U1865 (N_1865,In_295,In_570);
nand U1866 (N_1866,In_608,In_232);
or U1867 (N_1867,In_396,In_357);
nor U1868 (N_1868,In_380,In_14);
nand U1869 (N_1869,In_477,In_341);
or U1870 (N_1870,In_582,In_111);
and U1871 (N_1871,In_606,In_70);
nand U1872 (N_1872,In_150,In_600);
nand U1873 (N_1873,In_637,In_85);
nor U1874 (N_1874,In_734,In_587);
nand U1875 (N_1875,In_551,In_663);
nor U1876 (N_1876,In_695,In_178);
or U1877 (N_1877,In_260,In_543);
nor U1878 (N_1878,In_410,In_714);
or U1879 (N_1879,In_297,In_544);
and U1880 (N_1880,In_22,In_449);
and U1881 (N_1881,In_90,In_419);
nand U1882 (N_1882,In_602,In_202);
nor U1883 (N_1883,In_275,In_644);
and U1884 (N_1884,In_597,In_644);
nor U1885 (N_1885,In_494,In_383);
nor U1886 (N_1886,In_252,In_715);
nand U1887 (N_1887,In_136,In_597);
or U1888 (N_1888,In_699,In_729);
and U1889 (N_1889,In_471,In_306);
or U1890 (N_1890,In_483,In_248);
nor U1891 (N_1891,In_471,In_110);
and U1892 (N_1892,In_683,In_283);
or U1893 (N_1893,In_145,In_557);
or U1894 (N_1894,In_35,In_286);
nor U1895 (N_1895,In_599,In_256);
and U1896 (N_1896,In_363,In_467);
or U1897 (N_1897,In_499,In_566);
or U1898 (N_1898,In_660,In_521);
and U1899 (N_1899,In_559,In_48);
or U1900 (N_1900,In_193,In_410);
and U1901 (N_1901,In_500,In_364);
nand U1902 (N_1902,In_77,In_156);
and U1903 (N_1903,In_618,In_423);
nand U1904 (N_1904,In_441,In_362);
nor U1905 (N_1905,In_211,In_10);
nor U1906 (N_1906,In_635,In_549);
or U1907 (N_1907,In_77,In_531);
or U1908 (N_1908,In_737,In_443);
or U1909 (N_1909,In_505,In_555);
or U1910 (N_1910,In_25,In_620);
nor U1911 (N_1911,In_324,In_704);
nor U1912 (N_1912,In_495,In_339);
or U1913 (N_1913,In_48,In_31);
nand U1914 (N_1914,In_276,In_49);
or U1915 (N_1915,In_466,In_615);
or U1916 (N_1916,In_106,In_352);
nor U1917 (N_1917,In_659,In_539);
nand U1918 (N_1918,In_175,In_705);
or U1919 (N_1919,In_185,In_721);
and U1920 (N_1920,In_203,In_456);
and U1921 (N_1921,In_275,In_582);
and U1922 (N_1922,In_185,In_531);
nor U1923 (N_1923,In_747,In_503);
nand U1924 (N_1924,In_193,In_47);
or U1925 (N_1925,In_715,In_561);
or U1926 (N_1926,In_76,In_488);
or U1927 (N_1927,In_70,In_281);
nand U1928 (N_1928,In_6,In_393);
nand U1929 (N_1929,In_178,In_502);
and U1930 (N_1930,In_51,In_624);
nor U1931 (N_1931,In_365,In_250);
nand U1932 (N_1932,In_242,In_535);
or U1933 (N_1933,In_574,In_433);
nor U1934 (N_1934,In_354,In_438);
and U1935 (N_1935,In_633,In_323);
or U1936 (N_1936,In_247,In_96);
and U1937 (N_1937,In_609,In_748);
and U1938 (N_1938,In_550,In_313);
and U1939 (N_1939,In_354,In_660);
or U1940 (N_1940,In_59,In_596);
or U1941 (N_1941,In_458,In_370);
or U1942 (N_1942,In_264,In_278);
and U1943 (N_1943,In_261,In_284);
or U1944 (N_1944,In_171,In_413);
nor U1945 (N_1945,In_560,In_235);
and U1946 (N_1946,In_286,In_417);
nor U1947 (N_1947,In_295,In_427);
and U1948 (N_1948,In_464,In_586);
and U1949 (N_1949,In_136,In_555);
nand U1950 (N_1950,In_373,In_45);
and U1951 (N_1951,In_621,In_655);
nor U1952 (N_1952,In_409,In_30);
nand U1953 (N_1953,In_101,In_591);
nand U1954 (N_1954,In_503,In_705);
and U1955 (N_1955,In_396,In_446);
nand U1956 (N_1956,In_278,In_323);
or U1957 (N_1957,In_102,In_311);
and U1958 (N_1958,In_186,In_556);
nand U1959 (N_1959,In_541,In_634);
or U1960 (N_1960,In_666,In_332);
or U1961 (N_1961,In_185,In_19);
and U1962 (N_1962,In_638,In_393);
or U1963 (N_1963,In_560,In_485);
and U1964 (N_1964,In_159,In_166);
or U1965 (N_1965,In_425,In_201);
nand U1966 (N_1966,In_290,In_669);
or U1967 (N_1967,In_333,In_193);
nor U1968 (N_1968,In_636,In_244);
and U1969 (N_1969,In_562,In_296);
nor U1970 (N_1970,In_331,In_697);
nand U1971 (N_1971,In_440,In_11);
nor U1972 (N_1972,In_381,In_670);
and U1973 (N_1973,In_444,In_510);
nand U1974 (N_1974,In_94,In_720);
and U1975 (N_1975,In_300,In_736);
or U1976 (N_1976,In_86,In_693);
or U1977 (N_1977,In_238,In_699);
or U1978 (N_1978,In_473,In_74);
or U1979 (N_1979,In_430,In_485);
or U1980 (N_1980,In_43,In_640);
or U1981 (N_1981,In_538,In_420);
and U1982 (N_1982,In_245,In_647);
or U1983 (N_1983,In_121,In_364);
or U1984 (N_1984,In_278,In_74);
or U1985 (N_1985,In_278,In_665);
and U1986 (N_1986,In_68,In_178);
nand U1987 (N_1987,In_704,In_481);
and U1988 (N_1988,In_545,In_263);
or U1989 (N_1989,In_148,In_53);
nand U1990 (N_1990,In_215,In_360);
nor U1991 (N_1991,In_544,In_291);
nor U1992 (N_1992,In_565,In_344);
nand U1993 (N_1993,In_425,In_535);
nand U1994 (N_1994,In_507,In_258);
nand U1995 (N_1995,In_104,In_287);
or U1996 (N_1996,In_273,In_231);
or U1997 (N_1997,In_692,In_444);
or U1998 (N_1998,In_444,In_723);
nor U1999 (N_1999,In_436,In_341);
and U2000 (N_2000,In_743,In_461);
and U2001 (N_2001,In_516,In_723);
nand U2002 (N_2002,In_498,In_237);
and U2003 (N_2003,In_656,In_379);
or U2004 (N_2004,In_559,In_652);
and U2005 (N_2005,In_619,In_252);
nor U2006 (N_2006,In_493,In_373);
and U2007 (N_2007,In_628,In_236);
or U2008 (N_2008,In_344,In_669);
and U2009 (N_2009,In_509,In_333);
and U2010 (N_2010,In_522,In_500);
nor U2011 (N_2011,In_571,In_528);
nor U2012 (N_2012,In_270,In_28);
xnor U2013 (N_2013,In_180,In_671);
or U2014 (N_2014,In_400,In_52);
nand U2015 (N_2015,In_470,In_735);
nand U2016 (N_2016,In_12,In_206);
and U2017 (N_2017,In_740,In_586);
and U2018 (N_2018,In_553,In_356);
xor U2019 (N_2019,In_410,In_690);
or U2020 (N_2020,In_508,In_628);
or U2021 (N_2021,In_309,In_541);
nand U2022 (N_2022,In_283,In_123);
and U2023 (N_2023,In_423,In_394);
nor U2024 (N_2024,In_568,In_556);
or U2025 (N_2025,In_314,In_198);
nand U2026 (N_2026,In_234,In_16);
nor U2027 (N_2027,In_437,In_164);
and U2028 (N_2028,In_531,In_248);
nor U2029 (N_2029,In_626,In_57);
nand U2030 (N_2030,In_55,In_655);
or U2031 (N_2031,In_721,In_370);
and U2032 (N_2032,In_282,In_369);
or U2033 (N_2033,In_257,In_727);
nor U2034 (N_2034,In_362,In_483);
nor U2035 (N_2035,In_22,In_741);
nor U2036 (N_2036,In_118,In_385);
nand U2037 (N_2037,In_184,In_668);
or U2038 (N_2038,In_476,In_89);
nand U2039 (N_2039,In_177,In_524);
or U2040 (N_2040,In_476,In_11);
nand U2041 (N_2041,In_700,In_570);
and U2042 (N_2042,In_472,In_708);
nand U2043 (N_2043,In_450,In_354);
nor U2044 (N_2044,In_461,In_727);
or U2045 (N_2045,In_321,In_593);
or U2046 (N_2046,In_666,In_511);
nor U2047 (N_2047,In_361,In_523);
or U2048 (N_2048,In_576,In_519);
nor U2049 (N_2049,In_75,In_98);
nand U2050 (N_2050,In_124,In_538);
or U2051 (N_2051,In_275,In_420);
nor U2052 (N_2052,In_235,In_588);
nor U2053 (N_2053,In_298,In_727);
and U2054 (N_2054,In_561,In_233);
and U2055 (N_2055,In_737,In_228);
or U2056 (N_2056,In_402,In_523);
nand U2057 (N_2057,In_338,In_302);
or U2058 (N_2058,In_449,In_161);
or U2059 (N_2059,In_198,In_733);
or U2060 (N_2060,In_258,In_255);
or U2061 (N_2061,In_172,In_703);
or U2062 (N_2062,In_681,In_120);
nand U2063 (N_2063,In_582,In_628);
and U2064 (N_2064,In_462,In_386);
and U2065 (N_2065,In_361,In_254);
nor U2066 (N_2066,In_227,In_196);
or U2067 (N_2067,In_646,In_208);
nor U2068 (N_2068,In_20,In_139);
or U2069 (N_2069,In_431,In_563);
and U2070 (N_2070,In_565,In_231);
and U2071 (N_2071,In_611,In_264);
nor U2072 (N_2072,In_430,In_178);
or U2073 (N_2073,In_740,In_477);
xnor U2074 (N_2074,In_716,In_130);
and U2075 (N_2075,In_448,In_46);
or U2076 (N_2076,In_371,In_436);
nor U2077 (N_2077,In_282,In_580);
or U2078 (N_2078,In_32,In_114);
and U2079 (N_2079,In_65,In_137);
and U2080 (N_2080,In_165,In_590);
nor U2081 (N_2081,In_576,In_548);
and U2082 (N_2082,In_131,In_93);
or U2083 (N_2083,In_432,In_672);
and U2084 (N_2084,In_682,In_543);
and U2085 (N_2085,In_110,In_489);
nand U2086 (N_2086,In_366,In_492);
and U2087 (N_2087,In_647,In_731);
nor U2088 (N_2088,In_163,In_666);
or U2089 (N_2089,In_374,In_253);
and U2090 (N_2090,In_467,In_748);
nand U2091 (N_2091,In_246,In_89);
nand U2092 (N_2092,In_330,In_599);
or U2093 (N_2093,In_317,In_661);
and U2094 (N_2094,In_250,In_97);
and U2095 (N_2095,In_43,In_666);
nor U2096 (N_2096,In_671,In_271);
nand U2097 (N_2097,In_327,In_346);
nand U2098 (N_2098,In_359,In_218);
or U2099 (N_2099,In_548,In_594);
and U2100 (N_2100,In_5,In_448);
or U2101 (N_2101,In_506,In_481);
or U2102 (N_2102,In_137,In_420);
and U2103 (N_2103,In_733,In_234);
xor U2104 (N_2104,In_604,In_223);
xnor U2105 (N_2105,In_482,In_389);
or U2106 (N_2106,In_703,In_635);
nand U2107 (N_2107,In_244,In_41);
xnor U2108 (N_2108,In_532,In_542);
or U2109 (N_2109,In_227,In_203);
nor U2110 (N_2110,In_568,In_469);
nor U2111 (N_2111,In_179,In_290);
and U2112 (N_2112,In_520,In_291);
or U2113 (N_2113,In_343,In_25);
nor U2114 (N_2114,In_626,In_346);
or U2115 (N_2115,In_715,In_731);
nand U2116 (N_2116,In_425,In_691);
nand U2117 (N_2117,In_287,In_546);
and U2118 (N_2118,In_80,In_635);
nor U2119 (N_2119,In_426,In_457);
and U2120 (N_2120,In_28,In_269);
nand U2121 (N_2121,In_48,In_418);
nand U2122 (N_2122,In_623,In_505);
and U2123 (N_2123,In_195,In_474);
and U2124 (N_2124,In_270,In_171);
nand U2125 (N_2125,In_614,In_68);
and U2126 (N_2126,In_400,In_126);
xnor U2127 (N_2127,In_709,In_247);
nor U2128 (N_2128,In_723,In_640);
or U2129 (N_2129,In_438,In_568);
or U2130 (N_2130,In_155,In_398);
xor U2131 (N_2131,In_519,In_656);
or U2132 (N_2132,In_592,In_695);
or U2133 (N_2133,In_566,In_300);
or U2134 (N_2134,In_138,In_685);
or U2135 (N_2135,In_413,In_75);
nand U2136 (N_2136,In_612,In_322);
nor U2137 (N_2137,In_714,In_718);
or U2138 (N_2138,In_738,In_462);
nor U2139 (N_2139,In_570,In_360);
nor U2140 (N_2140,In_244,In_303);
and U2141 (N_2141,In_55,In_511);
and U2142 (N_2142,In_499,In_638);
and U2143 (N_2143,In_48,In_259);
nor U2144 (N_2144,In_587,In_89);
or U2145 (N_2145,In_389,In_677);
and U2146 (N_2146,In_305,In_332);
and U2147 (N_2147,In_686,In_190);
and U2148 (N_2148,In_581,In_309);
or U2149 (N_2149,In_313,In_635);
nand U2150 (N_2150,In_559,In_672);
nor U2151 (N_2151,In_425,In_87);
nand U2152 (N_2152,In_585,In_508);
and U2153 (N_2153,In_391,In_467);
xor U2154 (N_2154,In_25,In_236);
and U2155 (N_2155,In_58,In_403);
nor U2156 (N_2156,In_488,In_545);
and U2157 (N_2157,In_342,In_708);
and U2158 (N_2158,In_189,In_182);
nand U2159 (N_2159,In_303,In_563);
or U2160 (N_2160,In_698,In_727);
or U2161 (N_2161,In_471,In_131);
and U2162 (N_2162,In_526,In_589);
nand U2163 (N_2163,In_286,In_575);
nand U2164 (N_2164,In_346,In_349);
or U2165 (N_2165,In_3,In_579);
nand U2166 (N_2166,In_588,In_318);
and U2167 (N_2167,In_50,In_174);
nor U2168 (N_2168,In_532,In_202);
and U2169 (N_2169,In_152,In_740);
or U2170 (N_2170,In_474,In_61);
or U2171 (N_2171,In_7,In_726);
and U2172 (N_2172,In_565,In_717);
or U2173 (N_2173,In_342,In_642);
and U2174 (N_2174,In_434,In_97);
and U2175 (N_2175,In_401,In_419);
and U2176 (N_2176,In_698,In_630);
nor U2177 (N_2177,In_539,In_510);
and U2178 (N_2178,In_211,In_246);
and U2179 (N_2179,In_166,In_617);
and U2180 (N_2180,In_322,In_231);
nor U2181 (N_2181,In_36,In_11);
nand U2182 (N_2182,In_34,In_53);
nor U2183 (N_2183,In_605,In_588);
or U2184 (N_2184,In_552,In_730);
or U2185 (N_2185,In_486,In_350);
or U2186 (N_2186,In_180,In_61);
nand U2187 (N_2187,In_469,In_636);
nor U2188 (N_2188,In_515,In_56);
and U2189 (N_2189,In_84,In_30);
nor U2190 (N_2190,In_358,In_87);
or U2191 (N_2191,In_343,In_511);
and U2192 (N_2192,In_655,In_227);
nor U2193 (N_2193,In_30,In_570);
nand U2194 (N_2194,In_713,In_658);
and U2195 (N_2195,In_597,In_249);
nand U2196 (N_2196,In_739,In_199);
nor U2197 (N_2197,In_616,In_732);
or U2198 (N_2198,In_654,In_674);
nor U2199 (N_2199,In_523,In_31);
nand U2200 (N_2200,In_361,In_349);
nand U2201 (N_2201,In_445,In_567);
nor U2202 (N_2202,In_695,In_476);
and U2203 (N_2203,In_378,In_695);
and U2204 (N_2204,In_669,In_719);
nor U2205 (N_2205,In_427,In_737);
nor U2206 (N_2206,In_227,In_540);
nand U2207 (N_2207,In_481,In_366);
nor U2208 (N_2208,In_679,In_451);
or U2209 (N_2209,In_594,In_247);
nor U2210 (N_2210,In_482,In_229);
or U2211 (N_2211,In_689,In_87);
or U2212 (N_2212,In_654,In_537);
nor U2213 (N_2213,In_359,In_115);
or U2214 (N_2214,In_267,In_620);
nand U2215 (N_2215,In_187,In_449);
nor U2216 (N_2216,In_388,In_79);
nor U2217 (N_2217,In_475,In_372);
or U2218 (N_2218,In_180,In_654);
nor U2219 (N_2219,In_406,In_453);
and U2220 (N_2220,In_551,In_725);
nor U2221 (N_2221,In_292,In_525);
or U2222 (N_2222,In_450,In_169);
and U2223 (N_2223,In_391,In_75);
nor U2224 (N_2224,In_651,In_204);
nor U2225 (N_2225,In_192,In_58);
nor U2226 (N_2226,In_718,In_470);
and U2227 (N_2227,In_163,In_334);
or U2228 (N_2228,In_309,In_624);
nand U2229 (N_2229,In_66,In_717);
or U2230 (N_2230,In_482,In_240);
and U2231 (N_2231,In_165,In_452);
xor U2232 (N_2232,In_5,In_193);
nor U2233 (N_2233,In_639,In_303);
nand U2234 (N_2234,In_617,In_483);
and U2235 (N_2235,In_721,In_704);
nor U2236 (N_2236,In_569,In_663);
nand U2237 (N_2237,In_244,In_163);
or U2238 (N_2238,In_384,In_213);
and U2239 (N_2239,In_305,In_614);
nand U2240 (N_2240,In_747,In_572);
and U2241 (N_2241,In_624,In_665);
nand U2242 (N_2242,In_254,In_226);
nor U2243 (N_2243,In_26,In_681);
nor U2244 (N_2244,In_346,In_523);
nor U2245 (N_2245,In_537,In_679);
or U2246 (N_2246,In_390,In_633);
nand U2247 (N_2247,In_262,In_107);
and U2248 (N_2248,In_639,In_110);
nand U2249 (N_2249,In_497,In_427);
nand U2250 (N_2250,In_614,In_364);
or U2251 (N_2251,In_297,In_661);
and U2252 (N_2252,In_127,In_531);
and U2253 (N_2253,In_683,In_161);
or U2254 (N_2254,In_569,In_466);
or U2255 (N_2255,In_274,In_187);
nor U2256 (N_2256,In_15,In_101);
nand U2257 (N_2257,In_697,In_594);
nor U2258 (N_2258,In_367,In_384);
nand U2259 (N_2259,In_123,In_617);
nand U2260 (N_2260,In_58,In_622);
or U2261 (N_2261,In_59,In_421);
and U2262 (N_2262,In_706,In_448);
nor U2263 (N_2263,In_59,In_8);
or U2264 (N_2264,In_592,In_191);
nor U2265 (N_2265,In_243,In_698);
nor U2266 (N_2266,In_282,In_570);
nor U2267 (N_2267,In_590,In_373);
xor U2268 (N_2268,In_621,In_541);
xor U2269 (N_2269,In_164,In_603);
and U2270 (N_2270,In_363,In_283);
nand U2271 (N_2271,In_80,In_393);
and U2272 (N_2272,In_613,In_631);
nand U2273 (N_2273,In_242,In_258);
and U2274 (N_2274,In_171,In_486);
nand U2275 (N_2275,In_686,In_512);
nand U2276 (N_2276,In_19,In_534);
nand U2277 (N_2277,In_566,In_633);
or U2278 (N_2278,In_242,In_286);
nand U2279 (N_2279,In_88,In_167);
and U2280 (N_2280,In_24,In_399);
or U2281 (N_2281,In_304,In_73);
or U2282 (N_2282,In_574,In_539);
and U2283 (N_2283,In_360,In_275);
nor U2284 (N_2284,In_736,In_101);
nand U2285 (N_2285,In_509,In_339);
nor U2286 (N_2286,In_189,In_592);
or U2287 (N_2287,In_130,In_445);
and U2288 (N_2288,In_158,In_253);
and U2289 (N_2289,In_747,In_84);
nor U2290 (N_2290,In_413,In_186);
nand U2291 (N_2291,In_649,In_56);
nor U2292 (N_2292,In_624,In_671);
and U2293 (N_2293,In_98,In_601);
nor U2294 (N_2294,In_536,In_12);
or U2295 (N_2295,In_88,In_260);
or U2296 (N_2296,In_458,In_671);
and U2297 (N_2297,In_35,In_55);
and U2298 (N_2298,In_639,In_266);
xnor U2299 (N_2299,In_554,In_346);
nand U2300 (N_2300,In_698,In_296);
nand U2301 (N_2301,In_707,In_415);
and U2302 (N_2302,In_575,In_225);
or U2303 (N_2303,In_498,In_373);
nand U2304 (N_2304,In_349,In_534);
nand U2305 (N_2305,In_74,In_11);
and U2306 (N_2306,In_561,In_168);
nor U2307 (N_2307,In_365,In_371);
nor U2308 (N_2308,In_281,In_52);
nand U2309 (N_2309,In_400,In_141);
or U2310 (N_2310,In_332,In_20);
nand U2311 (N_2311,In_728,In_458);
and U2312 (N_2312,In_698,In_142);
nor U2313 (N_2313,In_131,In_526);
and U2314 (N_2314,In_403,In_749);
nand U2315 (N_2315,In_203,In_613);
or U2316 (N_2316,In_584,In_326);
nand U2317 (N_2317,In_717,In_347);
nand U2318 (N_2318,In_22,In_55);
nand U2319 (N_2319,In_426,In_305);
nor U2320 (N_2320,In_325,In_420);
nor U2321 (N_2321,In_649,In_464);
nor U2322 (N_2322,In_530,In_346);
nor U2323 (N_2323,In_172,In_41);
nand U2324 (N_2324,In_489,In_194);
nand U2325 (N_2325,In_101,In_194);
nand U2326 (N_2326,In_84,In_400);
or U2327 (N_2327,In_653,In_382);
nor U2328 (N_2328,In_444,In_733);
and U2329 (N_2329,In_114,In_44);
nand U2330 (N_2330,In_219,In_426);
and U2331 (N_2331,In_744,In_424);
and U2332 (N_2332,In_113,In_469);
and U2333 (N_2333,In_690,In_55);
or U2334 (N_2334,In_86,In_222);
or U2335 (N_2335,In_534,In_101);
or U2336 (N_2336,In_152,In_360);
or U2337 (N_2337,In_310,In_293);
and U2338 (N_2338,In_234,In_320);
nand U2339 (N_2339,In_222,In_19);
or U2340 (N_2340,In_496,In_524);
nand U2341 (N_2341,In_455,In_662);
or U2342 (N_2342,In_86,In_745);
nand U2343 (N_2343,In_258,In_375);
or U2344 (N_2344,In_621,In_255);
nand U2345 (N_2345,In_569,In_299);
or U2346 (N_2346,In_434,In_286);
and U2347 (N_2347,In_580,In_555);
or U2348 (N_2348,In_393,In_167);
nor U2349 (N_2349,In_561,In_281);
and U2350 (N_2350,In_549,In_191);
and U2351 (N_2351,In_60,In_332);
nor U2352 (N_2352,In_510,In_220);
nand U2353 (N_2353,In_278,In_623);
nand U2354 (N_2354,In_320,In_160);
nor U2355 (N_2355,In_213,In_241);
nor U2356 (N_2356,In_440,In_292);
nor U2357 (N_2357,In_374,In_562);
nand U2358 (N_2358,In_509,In_190);
and U2359 (N_2359,In_239,In_690);
or U2360 (N_2360,In_11,In_496);
or U2361 (N_2361,In_675,In_74);
nor U2362 (N_2362,In_534,In_583);
or U2363 (N_2363,In_420,In_436);
or U2364 (N_2364,In_106,In_92);
or U2365 (N_2365,In_646,In_49);
or U2366 (N_2366,In_129,In_438);
nand U2367 (N_2367,In_152,In_440);
and U2368 (N_2368,In_353,In_282);
and U2369 (N_2369,In_478,In_26);
nand U2370 (N_2370,In_160,In_334);
and U2371 (N_2371,In_564,In_650);
nand U2372 (N_2372,In_410,In_198);
or U2373 (N_2373,In_185,In_728);
or U2374 (N_2374,In_706,In_413);
xnor U2375 (N_2375,In_591,In_143);
nor U2376 (N_2376,In_717,In_521);
and U2377 (N_2377,In_97,In_571);
and U2378 (N_2378,In_521,In_394);
or U2379 (N_2379,In_105,In_536);
or U2380 (N_2380,In_279,In_13);
or U2381 (N_2381,In_80,In_574);
or U2382 (N_2382,In_542,In_470);
and U2383 (N_2383,In_567,In_21);
and U2384 (N_2384,In_626,In_598);
nand U2385 (N_2385,In_255,In_406);
and U2386 (N_2386,In_99,In_110);
nand U2387 (N_2387,In_427,In_525);
or U2388 (N_2388,In_167,In_473);
and U2389 (N_2389,In_92,In_222);
nand U2390 (N_2390,In_358,In_551);
or U2391 (N_2391,In_671,In_220);
or U2392 (N_2392,In_392,In_484);
and U2393 (N_2393,In_258,In_672);
nor U2394 (N_2394,In_740,In_101);
and U2395 (N_2395,In_222,In_591);
and U2396 (N_2396,In_572,In_187);
nor U2397 (N_2397,In_301,In_23);
or U2398 (N_2398,In_625,In_714);
xor U2399 (N_2399,In_324,In_187);
and U2400 (N_2400,In_411,In_132);
nor U2401 (N_2401,In_579,In_205);
and U2402 (N_2402,In_700,In_601);
and U2403 (N_2403,In_378,In_205);
nand U2404 (N_2404,In_459,In_203);
and U2405 (N_2405,In_676,In_565);
or U2406 (N_2406,In_612,In_680);
xnor U2407 (N_2407,In_272,In_38);
xor U2408 (N_2408,In_21,In_263);
nor U2409 (N_2409,In_500,In_96);
or U2410 (N_2410,In_677,In_728);
nand U2411 (N_2411,In_158,In_316);
and U2412 (N_2412,In_532,In_331);
nand U2413 (N_2413,In_143,In_401);
nand U2414 (N_2414,In_430,In_557);
and U2415 (N_2415,In_607,In_712);
and U2416 (N_2416,In_663,In_731);
or U2417 (N_2417,In_220,In_633);
or U2418 (N_2418,In_714,In_512);
or U2419 (N_2419,In_654,In_586);
nand U2420 (N_2420,In_257,In_149);
or U2421 (N_2421,In_189,In_404);
and U2422 (N_2422,In_528,In_480);
nand U2423 (N_2423,In_143,In_155);
and U2424 (N_2424,In_393,In_238);
and U2425 (N_2425,In_257,In_341);
nor U2426 (N_2426,In_106,In_441);
and U2427 (N_2427,In_125,In_279);
and U2428 (N_2428,In_219,In_462);
nor U2429 (N_2429,In_230,In_277);
nor U2430 (N_2430,In_633,In_383);
nand U2431 (N_2431,In_82,In_296);
nand U2432 (N_2432,In_237,In_100);
or U2433 (N_2433,In_319,In_303);
nand U2434 (N_2434,In_541,In_547);
or U2435 (N_2435,In_649,In_608);
nor U2436 (N_2436,In_270,In_670);
and U2437 (N_2437,In_404,In_609);
nand U2438 (N_2438,In_84,In_467);
and U2439 (N_2439,In_291,In_607);
nor U2440 (N_2440,In_450,In_26);
nor U2441 (N_2441,In_438,In_436);
nand U2442 (N_2442,In_629,In_276);
nor U2443 (N_2443,In_374,In_380);
nor U2444 (N_2444,In_599,In_5);
or U2445 (N_2445,In_100,In_734);
nand U2446 (N_2446,In_232,In_622);
or U2447 (N_2447,In_743,In_338);
xnor U2448 (N_2448,In_400,In_648);
and U2449 (N_2449,In_328,In_133);
and U2450 (N_2450,In_86,In_631);
nor U2451 (N_2451,In_558,In_678);
nand U2452 (N_2452,In_573,In_385);
nand U2453 (N_2453,In_579,In_639);
nor U2454 (N_2454,In_249,In_417);
and U2455 (N_2455,In_289,In_613);
and U2456 (N_2456,In_22,In_11);
nor U2457 (N_2457,In_200,In_92);
nand U2458 (N_2458,In_322,In_202);
or U2459 (N_2459,In_8,In_153);
nand U2460 (N_2460,In_612,In_333);
and U2461 (N_2461,In_107,In_571);
or U2462 (N_2462,In_172,In_195);
nand U2463 (N_2463,In_343,In_268);
nand U2464 (N_2464,In_509,In_702);
nand U2465 (N_2465,In_460,In_563);
nand U2466 (N_2466,In_361,In_316);
or U2467 (N_2467,In_727,In_529);
or U2468 (N_2468,In_77,In_52);
or U2469 (N_2469,In_316,In_529);
and U2470 (N_2470,In_302,In_669);
and U2471 (N_2471,In_360,In_697);
or U2472 (N_2472,In_76,In_598);
and U2473 (N_2473,In_548,In_267);
nand U2474 (N_2474,In_510,In_572);
or U2475 (N_2475,In_396,In_267);
and U2476 (N_2476,In_505,In_534);
and U2477 (N_2477,In_277,In_22);
or U2478 (N_2478,In_28,In_145);
or U2479 (N_2479,In_60,In_398);
and U2480 (N_2480,In_208,In_275);
nor U2481 (N_2481,In_259,In_64);
and U2482 (N_2482,In_591,In_301);
nand U2483 (N_2483,In_593,In_234);
nor U2484 (N_2484,In_35,In_712);
nand U2485 (N_2485,In_260,In_647);
or U2486 (N_2486,In_700,In_273);
nor U2487 (N_2487,In_633,In_303);
or U2488 (N_2488,In_707,In_213);
nor U2489 (N_2489,In_256,In_63);
nand U2490 (N_2490,In_582,In_145);
nand U2491 (N_2491,In_360,In_424);
nand U2492 (N_2492,In_318,In_428);
and U2493 (N_2493,In_626,In_405);
nor U2494 (N_2494,In_254,In_432);
nor U2495 (N_2495,In_736,In_622);
and U2496 (N_2496,In_343,In_708);
nor U2497 (N_2497,In_286,In_657);
and U2498 (N_2498,In_702,In_536);
nor U2499 (N_2499,In_640,In_301);
and U2500 (N_2500,N_487,N_1413);
or U2501 (N_2501,N_538,N_1354);
or U2502 (N_2502,N_2372,N_714);
nand U2503 (N_2503,N_1744,N_1871);
and U2504 (N_2504,N_1016,N_2124);
nor U2505 (N_2505,N_1041,N_1527);
and U2506 (N_2506,N_56,N_2097);
or U2507 (N_2507,N_2192,N_1003);
nor U2508 (N_2508,N_535,N_500);
and U2509 (N_2509,N_799,N_876);
nand U2510 (N_2510,N_750,N_790);
nand U2511 (N_2511,N_2035,N_2450);
nor U2512 (N_2512,N_1106,N_968);
nand U2513 (N_2513,N_383,N_1532);
and U2514 (N_2514,N_2171,N_331);
or U2515 (N_2515,N_1244,N_1704);
or U2516 (N_2516,N_1913,N_1553);
nor U2517 (N_2517,N_1454,N_443);
nand U2518 (N_2518,N_164,N_1612);
nor U2519 (N_2519,N_1241,N_1531);
nor U2520 (N_2520,N_2066,N_1536);
nand U2521 (N_2521,N_1408,N_603);
nand U2522 (N_2522,N_1473,N_567);
nor U2523 (N_2523,N_2222,N_2319);
and U2524 (N_2524,N_1535,N_1654);
and U2525 (N_2525,N_226,N_1051);
and U2526 (N_2526,N_2076,N_1824);
nand U2527 (N_2527,N_721,N_1503);
or U2528 (N_2528,N_1683,N_2281);
nand U2529 (N_2529,N_398,N_2037);
nor U2530 (N_2530,N_1034,N_2277);
and U2531 (N_2531,N_969,N_1272);
and U2532 (N_2532,N_1125,N_1036);
nand U2533 (N_2533,N_1079,N_674);
and U2534 (N_2534,N_1758,N_1848);
and U2535 (N_2535,N_1463,N_23);
or U2536 (N_2536,N_1234,N_2238);
or U2537 (N_2537,N_179,N_530);
nor U2538 (N_2538,N_1167,N_1073);
or U2539 (N_2539,N_1031,N_1649);
nor U2540 (N_2540,N_82,N_1653);
and U2541 (N_2541,N_34,N_687);
or U2542 (N_2542,N_1826,N_782);
nand U2543 (N_2543,N_76,N_411);
or U2544 (N_2544,N_1950,N_2459);
nand U2545 (N_2545,N_823,N_549);
or U2546 (N_2546,N_573,N_1193);
nand U2547 (N_2547,N_427,N_280);
or U2548 (N_2548,N_1081,N_1539);
nand U2549 (N_2549,N_1435,N_414);
nor U2550 (N_2550,N_645,N_1233);
and U2551 (N_2551,N_2114,N_1169);
and U2552 (N_2552,N_38,N_2472);
nor U2553 (N_2553,N_2479,N_2149);
or U2554 (N_2554,N_16,N_1357);
nor U2555 (N_2555,N_1652,N_9);
nor U2556 (N_2556,N_1059,N_517);
nor U2557 (N_2557,N_889,N_133);
or U2558 (N_2558,N_675,N_294);
nor U2559 (N_2559,N_2389,N_1483);
and U2560 (N_2560,N_551,N_2331);
nand U2561 (N_2561,N_1297,N_1542);
nand U2562 (N_2562,N_146,N_514);
or U2563 (N_2563,N_110,N_2273);
nor U2564 (N_2564,N_1734,N_1510);
and U2565 (N_2565,N_930,N_1586);
nor U2566 (N_2566,N_639,N_1486);
nor U2567 (N_2567,N_1991,N_1462);
nor U2568 (N_2568,N_712,N_1170);
or U2569 (N_2569,N_1964,N_169);
nor U2570 (N_2570,N_2410,N_1604);
xor U2571 (N_2571,N_915,N_2174);
and U2572 (N_2572,N_2407,N_116);
or U2573 (N_2573,N_887,N_800);
nor U2574 (N_2574,N_1330,N_583);
nand U2575 (N_2575,N_2460,N_1338);
or U2576 (N_2576,N_1847,N_1960);
nor U2577 (N_2577,N_2354,N_2451);
xor U2578 (N_2578,N_749,N_352);
and U2579 (N_2579,N_222,N_1597);
or U2580 (N_2580,N_1075,N_1537);
or U2581 (N_2581,N_694,N_385);
or U2582 (N_2582,N_1718,N_334);
or U2583 (N_2583,N_1690,N_1959);
or U2584 (N_2584,N_2255,N_1452);
nor U2585 (N_2585,N_1928,N_2417);
and U2586 (N_2586,N_929,N_27);
nor U2587 (N_2587,N_1884,N_1691);
nor U2588 (N_2588,N_631,N_1563);
or U2589 (N_2589,N_453,N_817);
and U2590 (N_2590,N_2313,N_586);
or U2591 (N_2591,N_2233,N_572);
and U2592 (N_2592,N_1095,N_1580);
and U2593 (N_2593,N_1213,N_1726);
or U2594 (N_2594,N_1516,N_1460);
or U2595 (N_2595,N_1828,N_1506);
nand U2596 (N_2596,N_1398,N_1485);
or U2597 (N_2597,N_1348,N_1882);
and U2598 (N_2598,N_2143,N_78);
nor U2599 (N_2599,N_1832,N_1720);
or U2600 (N_2600,N_2006,N_2396);
or U2601 (N_2601,N_1572,N_1663);
and U2602 (N_2602,N_1534,N_311);
nor U2603 (N_2603,N_2370,N_149);
or U2604 (N_2604,N_1515,N_123);
and U2605 (N_2605,N_346,N_1850);
nor U2606 (N_2606,N_776,N_2106);
nand U2607 (N_2607,N_1468,N_426);
or U2608 (N_2608,N_600,N_1443);
nor U2609 (N_2609,N_1956,N_1390);
or U2610 (N_2610,N_475,N_2317);
and U2611 (N_2611,N_508,N_771);
nand U2612 (N_2612,N_2302,N_1194);
nor U2613 (N_2613,N_175,N_136);
nand U2614 (N_2614,N_518,N_2007);
or U2615 (N_2615,N_1189,N_990);
and U2616 (N_2616,N_495,N_958);
nor U2617 (N_2617,N_2019,N_1638);
nor U2618 (N_2618,N_858,N_2258);
nand U2619 (N_2619,N_2327,N_1795);
or U2620 (N_2620,N_1214,N_1525);
or U2621 (N_2621,N_2293,N_594);
or U2622 (N_2622,N_2467,N_2286);
nand U2623 (N_2623,N_2146,N_1749);
nand U2624 (N_2624,N_1807,N_2115);
nand U2625 (N_2625,N_1102,N_1181);
and U2626 (N_2626,N_957,N_343);
nand U2627 (N_2627,N_1936,N_1076);
and U2628 (N_2628,N_230,N_2432);
nand U2629 (N_2629,N_1456,N_1695);
or U2630 (N_2630,N_1225,N_284);
and U2631 (N_2631,N_806,N_2185);
nor U2632 (N_2632,N_2247,N_2270);
nand U2633 (N_2633,N_2107,N_2080);
nor U2634 (N_2634,N_252,N_822);
or U2635 (N_2635,N_1256,N_2126);
and U2636 (N_2636,N_860,N_1881);
or U2637 (N_2637,N_2421,N_1627);
or U2638 (N_2638,N_2147,N_1090);
nand U2639 (N_2639,N_2200,N_2343);
or U2640 (N_2640,N_345,N_1687);
nand U2641 (N_2641,N_1714,N_1210);
nand U2642 (N_2642,N_834,N_509);
nor U2643 (N_2643,N_388,N_829);
or U2644 (N_2644,N_1015,N_643);
nor U2645 (N_2645,N_1990,N_202);
xnor U2646 (N_2646,N_42,N_141);
nand U2647 (N_2647,N_2390,N_1851);
or U2648 (N_2648,N_2043,N_576);
nor U2649 (N_2649,N_135,N_646);
and U2650 (N_2650,N_491,N_323);
nand U2651 (N_2651,N_2274,N_979);
and U2652 (N_2652,N_1126,N_644);
and U2653 (N_2653,N_168,N_2340);
and U2654 (N_2654,N_429,N_2379);
nand U2655 (N_2655,N_2353,N_1074);
and U2656 (N_2656,N_1717,N_2430);
and U2657 (N_2657,N_1440,N_1405);
and U2658 (N_2658,N_558,N_75);
or U2659 (N_2659,N_1885,N_1442);
nor U2660 (N_2660,N_2294,N_1138);
and U2661 (N_2661,N_1715,N_2401);
nor U2662 (N_2662,N_1127,N_1094);
or U2663 (N_2663,N_1495,N_2388);
nand U2664 (N_2664,N_1320,N_15);
or U2665 (N_2665,N_2119,N_1711);
nand U2666 (N_2666,N_1601,N_1505);
nor U2667 (N_2667,N_1781,N_708);
or U2668 (N_2668,N_1842,N_1300);
or U2669 (N_2669,N_1009,N_238);
or U2670 (N_2670,N_599,N_940);
nor U2671 (N_2671,N_895,N_139);
xnor U2672 (N_2672,N_1900,N_1310);
nand U2673 (N_2673,N_557,N_2234);
and U2674 (N_2674,N_1737,N_1615);
or U2675 (N_2675,N_2419,N_195);
or U2676 (N_2676,N_1467,N_1569);
nand U2677 (N_2677,N_321,N_709);
and U2678 (N_2678,N_1641,N_1886);
nand U2679 (N_2679,N_45,N_1038);
or U2680 (N_2680,N_105,N_550);
or U2681 (N_2681,N_531,N_1177);
or U2682 (N_2682,N_2018,N_1312);
or U2683 (N_2683,N_614,N_1710);
and U2684 (N_2684,N_2278,N_1668);
nor U2685 (N_2685,N_2497,N_949);
nand U2686 (N_2686,N_224,N_389);
or U2687 (N_2687,N_326,N_309);
xor U2688 (N_2688,N_544,N_2257);
nor U2689 (N_2689,N_366,N_2298);
nor U2690 (N_2690,N_2264,N_2304);
and U2691 (N_2691,N_547,N_1685);
and U2692 (N_2692,N_2160,N_2225);
and U2693 (N_2693,N_2486,N_265);
and U2694 (N_2694,N_754,N_1295);
nor U2695 (N_2695,N_1666,N_1629);
or U2696 (N_2696,N_401,N_359);
nor U2697 (N_2697,N_271,N_865);
and U2698 (N_2698,N_1,N_2178);
or U2699 (N_2699,N_2142,N_1943);
nand U2700 (N_2700,N_718,N_1644);
or U2701 (N_2701,N_1411,N_2055);
or U2702 (N_2702,N_702,N_962);
nand U2703 (N_2703,N_2334,N_312);
nor U2704 (N_2704,N_1289,N_2397);
nor U2705 (N_2705,N_1517,N_1209);
nor U2706 (N_2706,N_499,N_1776);
and U2707 (N_2707,N_2060,N_376);
nand U2708 (N_2708,N_1671,N_633);
or U2709 (N_2709,N_296,N_1684);
or U2710 (N_2710,N_1618,N_1918);
and U2711 (N_2711,N_1044,N_1277);
nor U2712 (N_2712,N_1757,N_484);
or U2713 (N_2713,N_605,N_2197);
nor U2714 (N_2714,N_1812,N_1201);
nand U2715 (N_2715,N_881,N_629);
or U2716 (N_2716,N_286,N_2038);
or U2717 (N_2717,N_2168,N_766);
nor U2718 (N_2718,N_19,N_2175);
nor U2719 (N_2719,N_1874,N_292);
xor U2720 (N_2720,N_1412,N_2437);
nand U2721 (N_2721,N_512,N_148);
nand U2722 (N_2722,N_457,N_2224);
xor U2723 (N_2723,N_216,N_2475);
xnor U2724 (N_2724,N_2189,N_1377);
or U2725 (N_2725,N_1820,N_540);
nor U2726 (N_2726,N_1645,N_696);
nand U2727 (N_2727,N_465,N_201);
or U2728 (N_2728,N_763,N_2116);
and U2729 (N_2729,N_268,N_1033);
nor U2730 (N_2730,N_1393,N_1249);
nand U2731 (N_2731,N_43,N_973);
nand U2732 (N_2732,N_2001,N_1856);
or U2733 (N_2733,N_2411,N_767);
or U2734 (N_2734,N_144,N_783);
and U2735 (N_2735,N_1342,N_282);
and U2736 (N_2736,N_618,N_789);
xnor U2737 (N_2737,N_1172,N_877);
and U2738 (N_2738,N_1676,N_1313);
nor U2739 (N_2739,N_1173,N_1797);
nor U2740 (N_2740,N_1543,N_1609);
or U2741 (N_2741,N_2363,N_1195);
and U2742 (N_2742,N_938,N_1366);
nand U2743 (N_2743,N_1843,N_2047);
nor U2744 (N_2744,N_920,N_2042);
and U2745 (N_2745,N_93,N_249);
and U2746 (N_2746,N_1765,N_681);
nor U2747 (N_2747,N_1533,N_1328);
nand U2748 (N_2748,N_2034,N_1566);
or U2749 (N_2749,N_2240,N_244);
and U2750 (N_2750,N_1864,N_1010);
or U2751 (N_2751,N_1325,N_1047);
xnor U2752 (N_2752,N_2265,N_1793);
nand U2753 (N_2753,N_337,N_1899);
and U2754 (N_2754,N_794,N_1931);
or U2755 (N_2755,N_701,N_1314);
xor U2756 (N_2756,N_2373,N_113);
nand U2757 (N_2757,N_37,N_951);
and U2758 (N_2758,N_220,N_306);
and U2759 (N_2759,N_2046,N_455);
nor U2760 (N_2760,N_1385,N_1846);
or U2761 (N_2761,N_1471,N_2470);
or U2762 (N_2762,N_1407,N_575);
or U2763 (N_2763,N_597,N_32);
and U2764 (N_2764,N_1046,N_1930);
or U2765 (N_2765,N_274,N_1021);
nand U2766 (N_2766,N_1528,N_68);
nand U2767 (N_2767,N_44,N_965);
or U2768 (N_2768,N_275,N_288);
nand U2769 (N_2769,N_368,N_406);
nand U2770 (N_2770,N_1925,N_662);
nand U2771 (N_2771,N_2408,N_1679);
nor U2772 (N_2772,N_1223,N_1363);
or U2773 (N_2773,N_2485,N_104);
nand U2774 (N_2774,N_2180,N_997);
or U2775 (N_2775,N_1431,N_170);
or U2776 (N_2776,N_1524,N_641);
and U2777 (N_2777,N_2182,N_581);
xor U2778 (N_2778,N_307,N_905);
nor U2779 (N_2779,N_1133,N_1317);
or U2780 (N_2780,N_843,N_2030);
nor U2781 (N_2781,N_1457,N_317);
nor U2782 (N_2782,N_519,N_742);
nand U2783 (N_2783,N_1947,N_793);
and U2784 (N_2784,N_983,N_992);
or U2785 (N_2785,N_1049,N_497);
and U2786 (N_2786,N_774,N_1067);
nor U2787 (N_2787,N_248,N_1453);
nand U2788 (N_2788,N_1660,N_647);
and U2789 (N_2789,N_1267,N_590);
and U2790 (N_2790,N_854,N_111);
and U2791 (N_2791,N_2112,N_1981);
or U2792 (N_2792,N_2099,N_1632);
nand U2793 (N_2793,N_1865,N_1809);
nand U2794 (N_2794,N_1592,N_811);
nand U2795 (N_2795,N_1492,N_290);
or U2796 (N_2796,N_1437,N_627);
nand U2797 (N_2797,N_1810,N_541);
nor U2798 (N_2798,N_2242,N_1334);
or U2799 (N_2799,N_2318,N_2414);
nand U2800 (N_2800,N_1712,N_243);
nor U2801 (N_2801,N_2431,N_2033);
or U2802 (N_2802,N_1029,N_47);
and U2803 (N_2803,N_1188,N_2089);
nand U2804 (N_2804,N_2365,N_2263);
or U2805 (N_2805,N_842,N_277);
or U2806 (N_2806,N_1155,N_1727);
or U2807 (N_2807,N_2138,N_2436);
or U2808 (N_2808,N_1083,N_959);
or U2809 (N_2809,N_2384,N_1551);
nand U2810 (N_2810,N_926,N_1845);
or U2811 (N_2811,N_577,N_1263);
nor U2812 (N_2812,N_1299,N_1661);
xnor U2813 (N_2813,N_1203,N_1337);
and U2814 (N_2814,N_1178,N_862);
or U2815 (N_2815,N_866,N_1305);
and U2816 (N_2816,N_1613,N_2315);
and U2817 (N_2817,N_893,N_784);
or U2818 (N_2818,N_1276,N_448);
and U2819 (N_2819,N_1974,N_1284);
nor U2820 (N_2820,N_879,N_2295);
and U2821 (N_2821,N_848,N_1153);
nand U2822 (N_2822,N_1139,N_370);
nand U2823 (N_2823,N_1441,N_10);
nand U2824 (N_2824,N_293,N_803);
and U2825 (N_2825,N_2194,N_121);
and U2826 (N_2826,N_438,N_261);
nor U2827 (N_2827,N_2013,N_917);
nand U2828 (N_2828,N_66,N_1103);
or U2829 (N_2829,N_2348,N_1622);
and U2830 (N_2830,N_2422,N_1101);
or U2831 (N_2831,N_1773,N_1731);
and U2832 (N_2832,N_1910,N_1970);
nor U2833 (N_2833,N_1351,N_344);
or U2834 (N_2834,N_871,N_863);
xnor U2835 (N_2835,N_1915,N_31);
nor U2836 (N_2836,N_122,N_2312);
or U2837 (N_2837,N_1388,N_838);
nor U2838 (N_2838,N_327,N_805);
and U2839 (N_2839,N_1800,N_1549);
and U2840 (N_2840,N_1257,N_2087);
nand U2841 (N_2841,N_301,N_2271);
and U2842 (N_2842,N_394,N_67);
nor U2843 (N_2843,N_205,N_1556);
nor U2844 (N_2844,N_1647,N_2064);
nor U2845 (N_2845,N_1617,N_1221);
nor U2846 (N_2846,N_489,N_1621);
or U2847 (N_2847,N_1493,N_1331);
or U2848 (N_2848,N_304,N_2166);
and U2849 (N_2849,N_2325,N_1252);
xor U2850 (N_2850,N_1771,N_1906);
or U2851 (N_2851,N_419,N_1590);
or U2852 (N_2852,N_3,N_1365);
xnor U2853 (N_2853,N_1476,N_788);
nor U2854 (N_2854,N_8,N_1821);
or U2855 (N_2855,N_1423,N_2049);
or U2856 (N_2856,N_827,N_186);
and U2857 (N_2857,N_2387,N_1326);
nand U2858 (N_2858,N_81,N_2151);
and U2859 (N_2859,N_387,N_977);
nand U2860 (N_2860,N_381,N_830);
nor U2861 (N_2861,N_1237,N_2031);
nor U2862 (N_2862,N_1369,N_658);
nand U2863 (N_2863,N_1939,N_1735);
nand U2864 (N_2864,N_1519,N_1013);
nand U2865 (N_2865,N_1039,N_209);
nor U2866 (N_2866,N_1513,N_2382);
and U2867 (N_2867,N_166,N_477);
or U2868 (N_2868,N_548,N_2050);
and U2869 (N_2869,N_1146,N_625);
nor U2870 (N_2870,N_1166,N_2056);
nor U2871 (N_2871,N_1219,N_1914);
and U2872 (N_2872,N_972,N_1762);
nor U2873 (N_2873,N_2405,N_1078);
and U2874 (N_2874,N_797,N_1466);
and U2875 (N_2875,N_2217,N_98);
xor U2876 (N_2876,N_1065,N_441);
nor U2877 (N_2877,N_1381,N_2193);
and U2878 (N_2878,N_761,N_1406);
and U2879 (N_2879,N_143,N_892);
nand U2880 (N_2880,N_552,N_682);
and U2881 (N_2881,N_2181,N_2254);
or U2882 (N_2882,N_437,N_1787);
nor U2883 (N_2883,N_1954,N_691);
or U2884 (N_2884,N_2288,N_2195);
or U2885 (N_2885,N_1581,N_1118);
xor U2886 (N_2886,N_2113,N_1056);
or U2887 (N_2887,N_4,N_713);
nand U2888 (N_2888,N_1656,N_154);
and U2889 (N_2889,N_1250,N_2393);
nand U2890 (N_2890,N_1107,N_260);
or U2891 (N_2891,N_2177,N_1161);
and U2892 (N_2892,N_1035,N_1967);
or U2893 (N_2893,N_1963,N_686);
nand U2894 (N_2894,N_2366,N_934);
nor U2895 (N_2895,N_1403,N_1246);
and U2896 (N_2896,N_172,N_924);
nor U2897 (N_2897,N_72,N_156);
nor U2898 (N_2898,N_1258,N_2184);
and U2899 (N_2899,N_1480,N_194);
and U2900 (N_2900,N_2469,N_1841);
and U2901 (N_2901,N_1979,N_1648);
and U2902 (N_2902,N_1268,N_996);
and U2903 (N_2903,N_1054,N_2108);
and U2904 (N_2904,N_1309,N_458);
and U2905 (N_2905,N_1937,N_1251);
or U2906 (N_2906,N_360,N_1595);
nor U2907 (N_2907,N_432,N_1285);
nand U2908 (N_2908,N_833,N_462);
nand U2909 (N_2909,N_693,N_55);
or U2910 (N_2910,N_1350,N_906);
and U2911 (N_2911,N_960,N_1426);
or U2912 (N_2912,N_1084,N_1111);
nand U2913 (N_2913,N_814,N_7);
nor U2914 (N_2914,N_1834,N_1414);
nand U2915 (N_2915,N_103,N_2332);
and U2916 (N_2916,N_1565,N_65);
nor U2917 (N_2917,N_1109,N_2008);
and U2918 (N_2918,N_1344,N_479);
or U2919 (N_2919,N_1057,N_595);
nor U2920 (N_2920,N_1477,N_1750);
and U2921 (N_2921,N_2232,N_1949);
nor U2922 (N_2922,N_351,N_719);
or U2923 (N_2923,N_2139,N_835);
nand U2924 (N_2924,N_246,N_1006);
or U2925 (N_2925,N_528,N_167);
nor U2926 (N_2926,N_467,N_1500);
nor U2927 (N_2927,N_199,N_231);
nand U2928 (N_2928,N_692,N_435);
or U2929 (N_2929,N_1863,N_142);
and U2930 (N_2930,N_2476,N_2322);
nand U2931 (N_2931,N_724,N_937);
or U2932 (N_2932,N_1026,N_613);
or U2933 (N_2933,N_971,N_506);
nand U2934 (N_2934,N_859,N_483);
nor U2935 (N_2935,N_1135,N_1708);
xor U2936 (N_2936,N_2446,N_95);
and U2937 (N_2937,N_1659,N_578);
and U2938 (N_2938,N_1790,N_2069);
nand U2939 (N_2939,N_2134,N_2214);
nand U2940 (N_2940,N_241,N_828);
and U2941 (N_2941,N_1802,N_1085);
and U2942 (N_2942,N_723,N_898);
and U2943 (N_2943,N_447,N_5);
and U2944 (N_2944,N_975,N_2094);
and U2945 (N_2945,N_1722,N_537);
nor U2946 (N_2946,N_191,N_1150);
nand U2947 (N_2947,N_24,N_1672);
or U2948 (N_2948,N_1953,N_2364);
or U2949 (N_2949,N_925,N_1394);
nand U2950 (N_2950,N_680,N_235);
nor U2951 (N_2951,N_634,N_1633);
or U2952 (N_2952,N_955,N_132);
nand U2953 (N_2953,N_472,N_1425);
and U2954 (N_2954,N_2082,N_1982);
and U2955 (N_2955,N_1419,N_1582);
nand U2956 (N_2956,N_1147,N_1825);
nand U2957 (N_2957,N_2117,N_1216);
or U2958 (N_2958,N_2091,N_1894);
or U2959 (N_2959,N_1152,N_2223);
nor U2960 (N_2960,N_1747,N_1245);
xnor U2961 (N_2961,N_1760,N_124);
or U2962 (N_2962,N_1444,N_2311);
nor U2963 (N_2963,N_2280,N_1099);
or U2964 (N_2964,N_1600,N_2127);
or U2965 (N_2965,N_1196,N_2416);
nand U2966 (N_2966,N_607,N_2499);
or U2967 (N_2967,N_33,N_386);
or U2968 (N_2968,N_2003,N_1635);
and U2969 (N_2969,N_916,N_1322);
nor U2970 (N_2970,N_1705,N_1164);
and U2971 (N_2971,N_2148,N_1860);
or U2972 (N_2972,N_521,N_885);
nor U2973 (N_2973,N_2457,N_2027);
or U2974 (N_2974,N_270,N_2346);
and U2975 (N_2975,N_2473,N_2358);
nand U2976 (N_2976,N_974,N_2110);
and U2977 (N_2977,N_2227,N_1677);
nor U2978 (N_2978,N_1301,N_772);
nor U2979 (N_2979,N_661,N_1417);
nor U2980 (N_2980,N_735,N_233);
and U2981 (N_2981,N_1128,N_2399);
xnor U2982 (N_2982,N_1025,N_1876);
and U2983 (N_2983,N_1465,N_470);
nand U2984 (N_2984,N_1883,N_2424);
nand U2985 (N_2985,N_1410,N_2095);
and U2986 (N_2986,N_2204,N_532);
nor U2987 (N_2987,N_942,N_856);
or U2988 (N_2988,N_1567,N_320);
nor U2989 (N_2989,N_812,N_555);
and U2990 (N_2990,N_2219,N_1968);
nand U2991 (N_2991,N_2483,N_267);
nand U2992 (N_2992,N_602,N_1852);
and U2993 (N_2993,N_1835,N_1742);
and U2994 (N_2994,N_1724,N_1593);
nor U2995 (N_2995,N_1288,N_886);
nand U2996 (N_2996,N_2386,N_1911);
and U2997 (N_2997,N_58,N_678);
nand U2998 (N_2998,N_2418,N_1611);
nand U2999 (N_2999,N_272,N_1253);
nand U3000 (N_3000,N_1857,N_109);
nor U3001 (N_3001,N_1973,N_1228);
nor U3002 (N_3002,N_2427,N_1694);
and U3003 (N_3003,N_740,N_2162);
nor U3004 (N_3004,N_26,N_1160);
and U3005 (N_3005,N_1307,N_1340);
or U3006 (N_3006,N_71,N_837);
nor U3007 (N_3007,N_283,N_931);
or U3008 (N_3008,N_2350,N_527);
nor U3009 (N_3009,N_1018,N_1247);
or U3010 (N_3010,N_1686,N_522);
nor U3011 (N_3011,N_1464,N_2191);
nor U3012 (N_3012,N_2282,N_77);
nor U3013 (N_3013,N_1319,N_1608);
and U3014 (N_3014,N_1907,N_593);
or U3015 (N_3015,N_444,N_372);
nor U3016 (N_3016,N_984,N_659);
nand U3017 (N_3017,N_1215,N_494);
xnor U3018 (N_3018,N_635,N_114);
and U3019 (N_3019,N_1670,N_2104);
or U3020 (N_3020,N_176,N_203);
nor U3021 (N_3021,N_2228,N_445);
nand U3022 (N_3022,N_878,N_433);
nand U3023 (N_3023,N_620,N_2447);
or U3024 (N_3024,N_1799,N_2471);
or U3025 (N_3025,N_193,N_513);
or U3026 (N_3026,N_1514,N_1576);
nor U3027 (N_3027,N_852,N_2010);
nor U3028 (N_3028,N_2017,N_1159);
or U3029 (N_3029,N_780,N_913);
or U3030 (N_3030,N_49,N_163);
nor U3031 (N_3031,N_371,N_1014);
and U3032 (N_3032,N_736,N_171);
and U3033 (N_3033,N_2190,N_650);
and U3034 (N_3034,N_2402,N_1372);
nand U3035 (N_3035,N_1439,N_1753);
nand U3036 (N_3036,N_945,N_785);
nand U3037 (N_3037,N_1623,N_824);
or U3038 (N_3038,N_1124,N_2310);
nand U3039 (N_3039,N_1662,N_1957);
nand U3040 (N_3040,N_1640,N_562);
nand U3041 (N_3041,N_449,N_2452);
or U3042 (N_3042,N_341,N_1148);
xnor U3043 (N_3043,N_2067,N_1889);
or U3044 (N_3044,N_970,N_382);
or U3045 (N_3045,N_2442,N_616);
and U3046 (N_3046,N_348,N_1027);
nand U3047 (N_3047,N_741,N_628);
or U3048 (N_3048,N_2212,N_744);
nor U3049 (N_3049,N_99,N_565);
nor U3050 (N_3050,N_332,N_727);
or U3051 (N_3051,N_430,N_731);
nand U3052 (N_3052,N_315,N_1198);
and U3053 (N_3053,N_1292,N_1206);
nor U3054 (N_3054,N_18,N_1625);
xor U3055 (N_3055,N_21,N_1869);
nor U3056 (N_3056,N_1725,N_1997);
or U3057 (N_3057,N_2020,N_468);
nand U3058 (N_3058,N_83,N_1012);
nor U3059 (N_3059,N_493,N_2023);
nor U3060 (N_3060,N_2005,N_1598);
nor U3061 (N_3061,N_2229,N_1007);
and U3062 (N_3062,N_966,N_2216);
and U3063 (N_3063,N_1341,N_2179);
and U3064 (N_3064,N_2203,N_2333);
nor U3065 (N_3065,N_2137,N_902);
and U3066 (N_3066,N_39,N_1512);
or U3067 (N_3067,N_1817,N_1266);
nand U3068 (N_3068,N_1236,N_1361);
nand U3069 (N_3069,N_621,N_1669);
or U3070 (N_3070,N_2368,N_1389);
or U3071 (N_3071,N_2285,N_87);
nand U3072 (N_3072,N_137,N_2157);
or U3073 (N_3073,N_2276,N_1782);
nand U3074 (N_3074,N_1643,N_297);
nand U3075 (N_3075,N_2128,N_2044);
and U3076 (N_3076,N_1294,N_2135);
or U3077 (N_3077,N_481,N_956);
and U3078 (N_3078,N_880,N_1375);
nor U3079 (N_3079,N_2239,N_107);
nand U3080 (N_3080,N_314,N_1329);
nand U3081 (N_3081,N_2132,N_994);
or U3082 (N_3082,N_2039,N_1978);
nand U3083 (N_3083,N_1738,N_2267);
or U3084 (N_3084,N_1501,N_1995);
and U3085 (N_3085,N_798,N_197);
and U3086 (N_3086,N_964,N_1430);
nor U3087 (N_3087,N_486,N_1129);
and U3088 (N_3088,N_2231,N_751);
and U3089 (N_3089,N_2156,N_1000);
nand U3090 (N_3090,N_2351,N_919);
nand U3091 (N_3091,N_900,N_642);
and U3092 (N_3092,N_303,N_753);
and U3093 (N_3093,N_276,N_1262);
nand U3094 (N_3094,N_706,N_349);
or U3095 (N_3095,N_2291,N_2339);
nor U3096 (N_3096,N_428,N_1827);
or U3097 (N_3097,N_2260,N_70);
and U3098 (N_3098,N_402,N_120);
xor U3099 (N_3099,N_1509,N_1154);
and U3100 (N_3100,N_374,N_350);
nand U3101 (N_3101,N_2026,N_1511);
nand U3102 (N_3102,N_851,N_1942);
nand U3103 (N_3103,N_764,N_2468);
nand U3104 (N_3104,N_1628,N_2283);
and U3105 (N_3105,N_57,N_273);
or U3106 (N_3106,N_1082,N_424);
nor U3107 (N_3107,N_289,N_730);
and U3108 (N_3108,N_606,N_463);
nand U3109 (N_3109,N_1089,N_725);
and U3110 (N_3110,N_2085,N_1119);
and U3111 (N_3111,N_2323,N_1469);
nand U3112 (N_3112,N_660,N_1575);
or U3113 (N_3113,N_1992,N_601);
and U3114 (N_3114,N_247,N_1192);
and U3115 (N_3115,N_1053,N_2439);
and U3116 (N_3116,N_988,N_2109);
nor U3117 (N_3117,N_2208,N_187);
and U3118 (N_3118,N_2187,N_2256);
and U3119 (N_3119,N_2070,N_897);
nor U3120 (N_3120,N_357,N_225);
or U3121 (N_3121,N_1678,N_1490);
and U3122 (N_3122,N_1571,N_1080);
or U3123 (N_3123,N_795,N_1657);
nor U3124 (N_3124,N_421,N_126);
or U3125 (N_3125,N_183,N_1449);
nand U3126 (N_3126,N_1055,N_325);
or U3127 (N_3127,N_2377,N_1190);
or U3128 (N_3128,N_1837,N_2303);
and U3129 (N_3129,N_1502,N_1696);
nand U3130 (N_3130,N_2335,N_2261);
and U3131 (N_3131,N_138,N_2464);
nand U3132 (N_3132,N_927,N_335);
nand U3133 (N_3133,N_2435,N_1822);
nor U3134 (N_3134,N_748,N_152);
nor U3135 (N_3135,N_1401,N_2266);
or U3136 (N_3136,N_459,N_669);
or U3137 (N_3137,N_1971,N_319);
nand U3138 (N_3138,N_568,N_1803);
or U3139 (N_3139,N_1767,N_1387);
and U3140 (N_3140,N_1713,N_476);
nor U3141 (N_3141,N_1522,N_1298);
nand U3142 (N_3142,N_1208,N_2367);
or U3143 (N_3143,N_1955,N_69);
nand U3144 (N_3144,N_1287,N_218);
or U3145 (N_3145,N_1355,N_354);
or U3146 (N_3146,N_36,N_1134);
or U3147 (N_3147,N_1175,N_2308);
nor U3148 (N_3148,N_115,N_1560);
nand U3149 (N_3149,N_2198,N_1370);
nor U3150 (N_3150,N_2048,N_2392);
nand U3151 (N_3151,N_2301,N_129);
nand U3152 (N_3152,N_416,N_1579);
or U3153 (N_3153,N_640,N_869);
or U3154 (N_3154,N_1853,N_2164);
nor U3155 (N_3155,N_251,N_1728);
xnor U3156 (N_3156,N_1784,N_192);
nand U3157 (N_3157,N_1286,N_1098);
nor U3158 (N_3158,N_752,N_546);
and U3159 (N_3159,N_2458,N_781);
or U3160 (N_3160,N_229,N_1792);
and U3161 (N_3161,N_511,N_2349);
or U3162 (N_3162,N_923,N_844);
nor U3163 (N_3163,N_1062,N_716);
nand U3164 (N_3164,N_579,N_1855);
nand U3165 (N_3165,N_2209,N_993);
or U3166 (N_3166,N_342,N_2300);
nand U3167 (N_3167,N_998,N_2131);
nand U3168 (N_3168,N_1770,N_2145);
or U3169 (N_3169,N_1174,N_2425);
or U3170 (N_3170,N_391,N_1472);
nand U3171 (N_3171,N_1667,N_1844);
nand U3172 (N_3172,N_1788,N_655);
and U3173 (N_3173,N_240,N_746);
and U3174 (N_3174,N_840,N_637);
xor U3175 (N_3175,N_777,N_850);
nor U3176 (N_3176,N_569,N_434);
and U3177 (N_3177,N_1069,N_40);
nand U3178 (N_3178,N_2016,N_291);
and U3179 (N_3179,N_456,N_2360);
and U3180 (N_3180,N_574,N_460);
nor U3181 (N_3181,N_816,N_1182);
nand U3182 (N_3182,N_1665,N_2100);
and U3183 (N_3183,N_2141,N_1752);
nor U3184 (N_3184,N_1642,N_1791);
nand U3185 (N_3185,N_1587,N_1227);
nor U3186 (N_3186,N_1120,N_873);
nor U3187 (N_3187,N_1922,N_198);
nand U3188 (N_3188,N_54,N_1819);
or U3189 (N_3189,N_1605,N_417);
nor U3190 (N_3190,N_415,N_399);
nor U3191 (N_3191,N_1554,N_2466);
and U3192 (N_3192,N_697,N_779);
nor U3193 (N_3193,N_1291,N_295);
or U3194 (N_3194,N_2461,N_1043);
nand U3195 (N_3195,N_1450,N_405);
nor U3196 (N_3196,N_1183,N_200);
nor U3197 (N_3197,N_1226,N_1114);
xor U3198 (N_3198,N_2245,N_807);
or U3199 (N_3199,N_664,N_670);
and U3200 (N_3200,N_80,N_1965);
nand U3201 (N_3201,N_1614,N_796);
or U3202 (N_3202,N_1934,N_1168);
or U3203 (N_3203,N_1550,N_932);
nor U3204 (N_3204,N_134,N_466);
nor U3205 (N_3205,N_755,N_2433);
nand U3206 (N_3206,N_2272,N_2040);
or U3207 (N_3207,N_1526,N_259);
nand U3208 (N_3208,N_2130,N_1022);
nor U3209 (N_3209,N_2292,N_2014);
nor U3210 (N_3210,N_2290,N_1574);
nand U3211 (N_3211,N_1323,N_396);
and U3212 (N_3212,N_79,N_1707);
nand U3213 (N_3213,N_269,N_308);
nor U3214 (N_3214,N_1151,N_74);
or U3215 (N_3215,N_1145,N_2326);
or U3216 (N_3216,N_1386,N_1895);
or U3217 (N_3217,N_2133,N_632);
nand U3218 (N_3218,N_1149,N_63);
or U3219 (N_3219,N_882,N_1261);
and U3220 (N_3220,N_804,N_2329);
or U3221 (N_3221,N_624,N_729);
nand U3222 (N_3222,N_1446,N_1558);
or U3223 (N_3223,N_991,N_1904);
nor U3224 (N_3224,N_1868,N_1830);
or U3225 (N_3225,N_2381,N_523);
nand U3226 (N_3226,N_1421,N_1786);
nand U3227 (N_3227,N_2230,N_53);
and U3228 (N_3228,N_1280,N_609);
or U3229 (N_3229,N_2449,N_84);
and U3230 (N_3230,N_219,N_1420);
nor U3231 (N_3231,N_663,N_1548);
and U3232 (N_3232,N_685,N_2120);
or U3233 (N_3233,N_849,N_2103);
or U3234 (N_3234,N_1023,N_1144);
xnor U3235 (N_3235,N_604,N_367);
nor U3236 (N_3236,N_864,N_162);
and U3237 (N_3237,N_60,N_648);
or U3238 (N_3238,N_305,N_2374);
or U3239 (N_3239,N_2355,N_813);
and U3240 (N_3240,N_263,N_1721);
and U3241 (N_3241,N_2098,N_1998);
nand U3242 (N_3242,N_2441,N_826);
nor U3243 (N_3243,N_1805,N_2380);
nor U3244 (N_3244,N_896,N_1602);
nor U3245 (N_3245,N_256,N_1115);
and U3246 (N_3246,N_1588,N_1137);
or U3247 (N_3247,N_1409,N_1362);
nor U3248 (N_3248,N_810,N_1887);
or U3249 (N_3249,N_158,N_2153);
or U3250 (N_3250,N_1603,N_1243);
and U3251 (N_3251,N_1254,N_1719);
or U3252 (N_3252,N_2202,N_801);
or U3253 (N_3253,N_841,N_1840);
and U3254 (N_3254,N_948,N_2395);
nand U3255 (N_3255,N_2086,N_2);
nor U3256 (N_3256,N_510,N_355);
nand U3257 (N_3257,N_839,N_196);
or U3258 (N_3258,N_1862,N_1242);
and U3259 (N_3259,N_952,N_1384);
nor U3260 (N_3260,N_596,N_228);
or U3261 (N_3261,N_2489,N_46);
or U3262 (N_3262,N_874,N_2385);
or U3263 (N_3263,N_953,N_1274);
and U3264 (N_3264,N_496,N_492);
or U3265 (N_3265,N_2188,N_1358);
nor U3266 (N_3266,N_180,N_1858);
nor U3267 (N_3267,N_1282,N_1958);
and U3268 (N_3268,N_707,N_328);
or U3269 (N_3269,N_1072,N_1585);
or U3270 (N_3270,N_2498,N_1064);
nor U3271 (N_3271,N_336,N_820);
and U3272 (N_3272,N_436,N_2218);
nand U3273 (N_3273,N_985,N_756);
and U3274 (N_3274,N_28,N_1920);
nor U3275 (N_3275,N_908,N_329);
or U3276 (N_3276,N_1202,N_1985);
and U3277 (N_3277,N_1966,N_2065);
nand U3278 (N_3278,N_1011,N_1296);
nand U3279 (N_3279,N_526,N_743);
nor U3280 (N_3280,N_2336,N_2000);
nor U3281 (N_3281,N_2361,N_1197);
nand U3282 (N_3282,N_1400,N_185);
and U3283 (N_3283,N_619,N_1917);
nand U3284 (N_3284,N_1230,N_1933);
or U3285 (N_3285,N_378,N_358);
nor U3286 (N_3286,N_1700,N_1379);
nand U3287 (N_3287,N_1356,N_980);
or U3288 (N_3288,N_704,N_1716);
and U3289 (N_3289,N_1759,N_2482);
nor U3290 (N_3290,N_1699,N_237);
or U3291 (N_3291,N_208,N_1199);
or U3292 (N_3292,N_90,N_1451);
nand U3293 (N_3293,N_97,N_883);
nor U3294 (N_3294,N_1231,N_206);
and U3295 (N_3295,N_1497,N_227);
and U3296 (N_3296,N_14,N_507);
nand U3297 (N_3297,N_2284,N_1271);
and U3298 (N_3298,N_440,N_770);
nor U3299 (N_3299,N_1415,N_1594);
and U3300 (N_3300,N_651,N_2015);
or U3301 (N_3301,N_933,N_130);
nand U3302 (N_3302,N_1655,N_2077);
and U3303 (N_3303,N_715,N_482);
xor U3304 (N_3304,N_1279,N_1599);
nand U3305 (N_3305,N_2211,N_2011);
and U3306 (N_3306,N_2118,N_1248);
nor U3307 (N_3307,N_2462,N_299);
xor U3308 (N_3308,N_1658,N_1304);
or U3309 (N_3309,N_2092,N_1042);
and U3310 (N_3310,N_987,N_1763);
nor U3311 (N_3311,N_1755,N_1674);
and U3312 (N_3312,N_316,N_989);
or U3313 (N_3313,N_1761,N_2096);
nand U3314 (N_3314,N_422,N_1769);
nand U3315 (N_3315,N_1577,N_1302);
nand U3316 (N_3316,N_2237,N_773);
nor U3317 (N_3317,N_1110,N_904);
nor U3318 (N_3318,N_454,N_1880);
and U3319 (N_3319,N_22,N_1264);
nor U3320 (N_3320,N_232,N_1583);
or U3321 (N_3321,N_1070,N_695);
nor U3322 (N_3322,N_1798,N_1890);
or U3323 (N_3323,N_947,N_395);
and U3324 (N_3324,N_2169,N_408);
nor U3325 (N_3325,N_1839,N_2152);
or U3326 (N_3326,N_1929,N_1702);
or U3327 (N_3327,N_1327,N_739);
and U3328 (N_3328,N_242,N_452);
nand U3329 (N_3329,N_1530,N_1673);
and U3330 (N_3330,N_73,N_1945);
and U3331 (N_3331,N_1220,N_2296);
and U3332 (N_3332,N_1545,N_559);
nand U3333 (N_3333,N_1481,N_1200);
and U3334 (N_3334,N_1801,N_1218);
and U3335 (N_3335,N_872,N_250);
or U3336 (N_3336,N_1131,N_2307);
nor U3337 (N_3337,N_1088,N_1924);
nor U3338 (N_3338,N_380,N_2477);
or U3339 (N_3339,N_1068,N_2199);
or U3340 (N_3340,N_119,N_722);
and U3341 (N_3341,N_2316,N_410);
nand U3342 (N_3342,N_1962,N_1240);
nor U3343 (N_3343,N_1459,N_791);
nand U3344 (N_3344,N_1416,N_1434);
and U3345 (N_3345,N_1020,N_2413);
nor U3346 (N_3346,N_50,N_1186);
or U3347 (N_3347,N_918,N_870);
nor U3348 (N_3348,N_1383,N_1772);
nor U3349 (N_3349,N_654,N_2009);
and U3350 (N_3350,N_671,N_1972);
and U3351 (N_3351,N_29,N_688);
nand U3352 (N_3352,N_266,N_2415);
and U3353 (N_3353,N_125,N_1060);
or U3354 (N_3354,N_653,N_553);
or U3355 (N_3355,N_2073,N_1112);
or U3356 (N_3356,N_59,N_978);
nor U3357 (N_3357,N_1736,N_2403);
or U3358 (N_3358,N_1610,N_2246);
or U3359 (N_3359,N_287,N_1392);
xnor U3360 (N_3360,N_836,N_1838);
and U3361 (N_3361,N_1999,N_720);
and U3362 (N_3362,N_1378,N_2165);
nand U3363 (N_3363,N_1651,N_1570);
nor U3364 (N_3364,N_418,N_1650);
nand U3365 (N_3365,N_1391,N_1898);
or U3366 (N_3366,N_2341,N_1816);
or U3367 (N_3367,N_2320,N_2481);
or U3368 (N_3368,N_1359,N_2352);
nor U3369 (N_3369,N_2321,N_2356);
and U3370 (N_3370,N_999,N_471);
and U3371 (N_3371,N_907,N_1902);
or U3372 (N_3372,N_390,N_899);
nor U3373 (N_3373,N_909,N_2478);
nand U3374 (N_3374,N_488,N_747);
xnor U3375 (N_3375,N_738,N_536);
and U3376 (N_3376,N_298,N_101);
or U3377 (N_3377,N_1001,N_1158);
nor U3378 (N_3378,N_1275,N_982);
nand U3379 (N_3379,N_818,N_262);
nand U3380 (N_3380,N_775,N_1071);
or U3381 (N_3381,N_1993,N_214);
nor U3382 (N_3382,N_41,N_20);
or U3383 (N_3383,N_1589,N_425);
and U3384 (N_3384,N_1897,N_1723);
nand U3385 (N_3385,N_285,N_1368);
and U3386 (N_3386,N_1052,N_1458);
and U3387 (N_3387,N_1424,N_2102);
and U3388 (N_3388,N_1232,N_324);
nand U3389 (N_3389,N_912,N_1607);
nor U3390 (N_3390,N_1489,N_25);
and U3391 (N_3391,N_2306,N_1831);
nor U3392 (N_3392,N_1521,N_1562);
nor U3393 (N_3393,N_369,N_1681);
and U3394 (N_3394,N_1373,N_48);
and U3395 (N_3395,N_534,N_2154);
nand U3396 (N_3396,N_177,N_1422);
xnor U3397 (N_3397,N_1775,N_2111);
nand U3398 (N_3398,N_554,N_1318);
nand U3399 (N_3399,N_524,N_365);
nor U3400 (N_3400,N_1353,N_1849);
and U3401 (N_3401,N_189,N_1335);
and U3402 (N_3402,N_1428,N_533);
or U3403 (N_3403,N_1396,N_153);
nand U3404 (N_3404,N_1634,N_1606);
and U3405 (N_3405,N_234,N_726);
or U3406 (N_3406,N_501,N_1157);
and U3407 (N_3407,N_2391,N_683);
or U3408 (N_3408,N_1584,N_703);
and U3409 (N_3409,N_62,N_1541);
or U3410 (N_3410,N_589,N_1345);
or U3411 (N_3411,N_1946,N_728);
nor U3412 (N_3412,N_1316,N_1557);
and U3413 (N_3413,N_1961,N_1156);
or U3414 (N_3414,N_1751,N_1877);
xnor U3415 (N_3415,N_2299,N_1764);
and U3416 (N_3416,N_1896,N_1892);
nor U3417 (N_3417,N_944,N_1017);
nor U3418 (N_3418,N_1281,N_51);
xor U3419 (N_3419,N_1132,N_2071);
nand U3420 (N_3420,N_2434,N_1496);
nand U3421 (N_3421,N_888,N_181);
and U3422 (N_3422,N_1980,N_1427);
nand U3423 (N_3423,N_2078,N_128);
nor U3424 (N_3424,N_264,N_626);
or U3425 (N_3425,N_157,N_1813);
or U3426 (N_3426,N_2121,N_1879);
nand U3427 (N_3427,N_1701,N_1418);
nor U3428 (N_3428,N_379,N_1058);
nor U3429 (N_3429,N_608,N_1766);
or U3430 (N_3430,N_1290,N_1171);
nor U3431 (N_3431,N_112,N_1620);
nor U3432 (N_3432,N_1494,N_1815);
and U3433 (N_3433,N_1901,N_2173);
nand U3434 (N_3434,N_2314,N_2068);
and U3435 (N_3435,N_2215,N_300);
nor U3436 (N_3436,N_2344,N_950);
nand U3437 (N_3437,N_1278,N_155);
nand U3438 (N_3438,N_480,N_1212);
nor U3439 (N_3439,N_118,N_2455);
nand U3440 (N_3440,N_1987,N_733);
or U3441 (N_3441,N_758,N_2375);
nand U3442 (N_3442,N_1923,N_1140);
nand U3443 (N_3443,N_1507,N_787);
nand U3444 (N_3444,N_1371,N_928);
xnor U3445 (N_3445,N_2081,N_1975);
nor U3446 (N_3446,N_914,N_1944);
and U3447 (N_3447,N_768,N_1349);
and U3448 (N_3448,N_212,N_502);
or U3449 (N_3449,N_498,N_140);
nor U3450 (N_3450,N_1814,N_1045);
or U3451 (N_3451,N_2123,N_2324);
or U3452 (N_3452,N_2454,N_461);
nand U3453 (N_3453,N_1487,N_1087);
nor U3454 (N_3454,N_1854,N_737);
nor U3455 (N_3455,N_2079,N_1096);
nor U3456 (N_3456,N_1180,N_2487);
nand U3457 (N_3457,N_2206,N_1740);
nand U3458 (N_3458,N_853,N_339);
and U3459 (N_3459,N_1888,N_1872);
nand U3460 (N_3460,N_1455,N_2205);
xnor U3461 (N_3461,N_313,N_1692);
nand U3462 (N_3462,N_571,N_88);
nand U3463 (N_3463,N_2371,N_1048);
and U3464 (N_3464,N_2093,N_2101);
or U3465 (N_3465,N_255,N_1664);
nor U3466 (N_3466,N_1938,N_2480);
or U3467 (N_3467,N_2438,N_1352);
and U3468 (N_3468,N_1818,N_0);
and U3469 (N_3469,N_30,N_1321);
and U3470 (N_3470,N_2369,N_147);
and U3471 (N_3471,N_1395,N_667);
nand U3472 (N_3472,N_1004,N_778);
nor U3473 (N_3473,N_745,N_1706);
nand U3474 (N_3474,N_666,N_165);
nand U3475 (N_3475,N_2012,N_2236);
nor U3476 (N_3476,N_1121,N_566);
nand U3477 (N_3477,N_503,N_1024);
nand U3478 (N_3478,N_2495,N_204);
or U3479 (N_3479,N_1732,N_847);
nor U3480 (N_3480,N_2297,N_2022);
nor U3481 (N_3481,N_1037,N_1564);
or U3482 (N_3482,N_563,N_1983);
and U3483 (N_3483,N_556,N_2426);
or U3484 (N_3484,N_1315,N_954);
or U3485 (N_3485,N_1308,N_1136);
or U3486 (N_3486,N_1927,N_1996);
nor U3487 (N_3487,N_279,N_1544);
nand U3488 (N_3488,N_855,N_322);
and U3489 (N_3489,N_2494,N_1754);
nor U3490 (N_3490,N_258,N_679);
nor U3491 (N_3491,N_543,N_1093);
or U3492 (N_3492,N_2210,N_2428);
nand U3493 (N_3493,N_2183,N_1104);
nand U3494 (N_3494,N_1682,N_1207);
or U3495 (N_3495,N_2243,N_1552);
and U3496 (N_3496,N_1921,N_2059);
nand U3497 (N_3497,N_2378,N_1829);
nand U3498 (N_3498,N_2004,N_353);
or U3499 (N_3499,N_677,N_2342);
nand U3500 (N_3500,N_281,N_588);
nor U3501 (N_3501,N_976,N_1893);
nor U3502 (N_3502,N_710,N_173);
and U3503 (N_3503,N_1229,N_2105);
and U3504 (N_3504,N_1097,N_2021);
or U3505 (N_3505,N_1867,N_89);
and U3506 (N_3506,N_1559,N_2029);
or U3507 (N_3507,N_1113,N_2176);
and U3508 (N_3508,N_375,N_1402);
or U3509 (N_3509,N_580,N_967);
nand U3510 (N_3510,N_2420,N_819);
or U3511 (N_3511,N_2088,N_1836);
nor U3512 (N_3512,N_2002,N_1478);
nand U3513 (N_3513,N_717,N_2158);
or U3514 (N_3514,N_221,N_151);
or U3515 (N_3515,N_1086,N_1919);
nand U3516 (N_3516,N_2032,N_1529);
or U3517 (N_3517,N_617,N_1336);
and U3518 (N_3518,N_431,N_404);
nand U3519 (N_3519,N_1008,N_377);
nand U3520 (N_3520,N_330,N_1555);
nor U3521 (N_3521,N_2083,N_2201);
nand U3522 (N_3522,N_1940,N_1680);
or U3523 (N_3523,N_1891,N_961);
nor U3524 (N_3524,N_1806,N_1474);
and U3525 (N_3525,N_520,N_2159);
and U3526 (N_3526,N_2062,N_2412);
and U3527 (N_3527,N_591,N_1260);
nand U3528 (N_3528,N_1165,N_1143);
nand U3529 (N_3529,N_1774,N_1698);
or U3530 (N_3530,N_1688,N_1374);
and U3531 (N_3531,N_2337,N_2136);
nor U3532 (N_3532,N_2289,N_178);
nor U3533 (N_3533,N_2057,N_1878);
and U3534 (N_3534,N_1743,N_1538);
and U3535 (N_3535,N_699,N_2404);
nand U3536 (N_3536,N_2129,N_2493);
and U3537 (N_3537,N_2150,N_318);
or U3538 (N_3538,N_560,N_1429);
nor U3539 (N_3539,N_2328,N_1399);
or U3540 (N_3540,N_1745,N_1508);
or U3541 (N_3541,N_875,N_2155);
xor U3542 (N_3542,N_1689,N_2448);
and U3543 (N_3543,N_1498,N_1448);
and U3544 (N_3544,N_2253,N_420);
nand U3545 (N_3545,N_921,N_108);
and U3546 (N_3546,N_12,N_2309);
nor U3547 (N_3547,N_1804,N_1916);
and U3548 (N_3548,N_1191,N_757);
xnor U3549 (N_3549,N_759,N_1573);
or U3550 (N_3550,N_1092,N_2305);
nor U3551 (N_3551,N_2406,N_2443);
and U3552 (N_3552,N_1491,N_1908);
or U3553 (N_3553,N_1063,N_2041);
nor U3554 (N_3554,N_159,N_1547);
or U3555 (N_3555,N_808,N_809);
nor U3556 (N_3556,N_1293,N_2140);
and U3557 (N_3557,N_1265,N_1905);
nand U3558 (N_3558,N_446,N_689);
nand U3559 (N_3559,N_894,N_1259);
nor U3560 (N_3560,N_1311,N_762);
or U3561 (N_3561,N_1100,N_2052);
and U3562 (N_3562,N_474,N_86);
nor U3563 (N_3563,N_2268,N_672);
and U3564 (N_3564,N_473,N_890);
nand U3565 (N_3565,N_1116,N_2163);
nand U3566 (N_3566,N_2440,N_384);
nand U3567 (N_3567,N_1748,N_1780);
or U3568 (N_3568,N_2244,N_711);
nor U3569 (N_3569,N_1382,N_2259);
nor U3570 (N_3570,N_1540,N_310);
and U3571 (N_3571,N_1546,N_676);
or U3572 (N_3572,N_2484,N_2063);
or U3573 (N_3573,N_734,N_1903);
nor U3574 (N_3574,N_2362,N_1941);
nand U3575 (N_3575,N_1211,N_407);
nor U3576 (N_3576,N_2488,N_127);
nand U3577 (N_3577,N_561,N_1484);
or U3578 (N_3578,N_1789,N_515);
or U3579 (N_3579,N_1630,N_769);
nand U3580 (N_3580,N_1433,N_867);
nand U3581 (N_3581,N_1238,N_2252);
and U3582 (N_3582,N_582,N_1823);
nand U3583 (N_3583,N_1032,N_1224);
nand U3584 (N_3584,N_2490,N_1204);
xnor U3585 (N_3585,N_392,N_2345);
nand U3586 (N_3586,N_1866,N_1596);
and U3587 (N_3587,N_182,N_652);
nand U3588 (N_3588,N_469,N_1028);
and U3589 (N_3589,N_1270,N_1768);
nor U3590 (N_3590,N_910,N_2269);
and U3591 (N_3591,N_393,N_615);
nand U3592 (N_3592,N_690,N_2445);
and U3593 (N_3593,N_939,N_1520);
nand U3594 (N_3594,N_1951,N_903);
nor U3595 (N_3595,N_1636,N_943);
and U3596 (N_3596,N_2125,N_884);
nand U3597 (N_3597,N_821,N_362);
and U3598 (N_3598,N_2051,N_2330);
nand U3599 (N_3599,N_2074,N_936);
or U3600 (N_3600,N_1364,N_542);
and U3601 (N_3601,N_2170,N_2429);
and U3602 (N_3602,N_215,N_91);
nor U3603 (N_3603,N_1269,N_1040);
nor U3604 (N_3604,N_610,N_657);
nand U3605 (N_3605,N_1255,N_409);
or U3606 (N_3606,N_2248,N_347);
nor U3607 (N_3607,N_2084,N_450);
and U3608 (N_3608,N_1367,N_439);
and U3609 (N_3609,N_684,N_13);
and U3610 (N_3610,N_1637,N_1729);
or U3611 (N_3611,N_1141,N_190);
nor U3612 (N_3612,N_211,N_705);
or U3613 (N_3613,N_1432,N_2262);
nand U3614 (N_3614,N_1185,N_1303);
nand U3615 (N_3615,N_2220,N_1504);
nor U3616 (N_3616,N_1163,N_2172);
and U3617 (N_3617,N_700,N_2359);
or U3618 (N_3618,N_901,N_1926);
or U3619 (N_3619,N_1808,N_612);
and U3620 (N_3620,N_2054,N_2028);
or U3621 (N_3621,N_1176,N_2036);
nor U3622 (N_3622,N_1777,N_1875);
nor U3623 (N_3623,N_174,N_529);
or U3624 (N_3624,N_340,N_1447);
or U3625 (N_3625,N_765,N_1631);
xor U3626 (N_3626,N_1977,N_1333);
or U3627 (N_3627,N_831,N_946);
xor U3628 (N_3628,N_1619,N_1693);
nand U3629 (N_3629,N_2376,N_364);
or U3630 (N_3630,N_333,N_1475);
and U3631 (N_3631,N_207,N_539);
xnor U3632 (N_3632,N_1488,N_52);
nand U3633 (N_3633,N_106,N_1184);
and U3634 (N_3634,N_423,N_846);
nor U3635 (N_3635,N_1091,N_1332);
nand U3636 (N_3636,N_2058,N_656);
or U3637 (N_3637,N_1343,N_638);
and U3638 (N_3638,N_92,N_1746);
nor U3639 (N_3639,N_1626,N_1239);
nor U3640 (N_3640,N_2275,N_598);
nor U3641 (N_3641,N_2492,N_1989);
nand U3642 (N_3642,N_911,N_1019);
and U3643 (N_3643,N_2241,N_963);
xor U3644 (N_3644,N_2221,N_1870);
nor U3645 (N_3645,N_2090,N_649);
and U3646 (N_3646,N_2075,N_1796);
nor U3647 (N_3647,N_1912,N_1785);
nand U3648 (N_3648,N_210,N_257);
xor U3649 (N_3649,N_630,N_1794);
and U3650 (N_3650,N_2453,N_117);
xnor U3651 (N_3651,N_636,N_1932);
nor U3652 (N_3652,N_464,N_504);
or U3653 (N_3653,N_505,N_825);
nor U3654 (N_3654,N_1050,N_1646);
nor U3655 (N_3655,N_935,N_995);
nand U3656 (N_3656,N_1205,N_585);
or U3657 (N_3657,N_1142,N_1988);
nand U3658 (N_3658,N_61,N_35);
nor U3659 (N_3659,N_102,N_1030);
or U3660 (N_3660,N_413,N_1741);
and U3661 (N_3661,N_1952,N_622);
nand U3662 (N_3662,N_490,N_373);
and U3663 (N_3663,N_2456,N_732);
nand U3664 (N_3664,N_665,N_400);
or U3665 (N_3665,N_1783,N_1235);
nand U3666 (N_3666,N_1123,N_1873);
and U3667 (N_3667,N_1380,N_1162);
and U3668 (N_3668,N_1179,N_1935);
or U3669 (N_3669,N_1984,N_2122);
and U3670 (N_3670,N_100,N_239);
and U3671 (N_3671,N_1778,N_1436);
or U3672 (N_3672,N_2024,N_1339);
nor U3673 (N_3673,N_442,N_1306);
or U3674 (N_3674,N_1499,N_188);
nor U3675 (N_3675,N_2249,N_2398);
nand U3676 (N_3676,N_356,N_868);
or U3677 (N_3677,N_587,N_2400);
nand U3678 (N_3678,N_2226,N_891);
or U3679 (N_3679,N_1482,N_397);
nor U3680 (N_3680,N_2251,N_1739);
nor U3681 (N_3681,N_1061,N_1187);
or U3682 (N_3682,N_1861,N_584);
and U3683 (N_3683,N_2357,N_1105);
xor U3684 (N_3684,N_2196,N_2235);
or U3685 (N_3685,N_2167,N_1518);
nor U3686 (N_3686,N_1568,N_2186);
nand U3687 (N_3687,N_1122,N_2279);
or U3688 (N_3688,N_1578,N_1324);
and U3689 (N_3689,N_2394,N_698);
nor U3690 (N_3690,N_403,N_485);
nor U3691 (N_3691,N_150,N_1346);
or U3692 (N_3692,N_1130,N_1347);
and U3693 (N_3693,N_668,N_1108);
or U3694 (N_3694,N_786,N_2496);
and U3695 (N_3695,N_802,N_2423);
or U3696 (N_3696,N_1697,N_85);
or U3697 (N_3697,N_1273,N_94);
nand U3698 (N_3698,N_2061,N_1117);
nand U3699 (N_3699,N_236,N_17);
nand U3700 (N_3700,N_1969,N_1709);
or U3701 (N_3701,N_160,N_611);
and U3702 (N_3702,N_861,N_338);
nor U3703 (N_3703,N_223,N_1639);
and U3704 (N_3704,N_2144,N_623);
and U3705 (N_3705,N_1909,N_1976);
nor U3706 (N_3706,N_2491,N_2207);
and U3707 (N_3707,N_570,N_1461);
and U3708 (N_3708,N_1077,N_1624);
and U3709 (N_3709,N_1397,N_1733);
or U3710 (N_3710,N_1222,N_986);
and U3711 (N_3711,N_184,N_1561);
nor U3712 (N_3712,N_1986,N_1675);
nor U3713 (N_3713,N_1470,N_792);
or U3714 (N_3714,N_145,N_253);
nand U3715 (N_3715,N_2161,N_1479);
and U3716 (N_3716,N_2072,N_363);
xor U3717 (N_3717,N_245,N_2444);
and U3718 (N_3718,N_1859,N_941);
xor U3719 (N_3719,N_2053,N_1066);
nand U3720 (N_3720,N_922,N_545);
and U3721 (N_3721,N_832,N_2025);
nand U3722 (N_3722,N_1833,N_760);
or U3723 (N_3723,N_673,N_2347);
and U3724 (N_3724,N_161,N_96);
or U3725 (N_3725,N_1994,N_412);
nand U3726 (N_3726,N_1730,N_857);
nor U3727 (N_3727,N_1591,N_2045);
nor U3728 (N_3728,N_516,N_2338);
and U3729 (N_3729,N_1948,N_1002);
or U3730 (N_3730,N_564,N_478);
or U3731 (N_3731,N_1376,N_2213);
and U3732 (N_3732,N_213,N_2287);
nor U3733 (N_3733,N_2474,N_525);
nand U3734 (N_3734,N_451,N_1445);
and U3735 (N_3735,N_2409,N_1404);
nand U3736 (N_3736,N_1811,N_815);
nand U3737 (N_3737,N_64,N_11);
and U3738 (N_3738,N_1438,N_6);
and U3739 (N_3739,N_845,N_1703);
and U3740 (N_3740,N_361,N_1360);
nand U3741 (N_3741,N_1616,N_1779);
nor U3742 (N_3742,N_981,N_1217);
xnor U3743 (N_3743,N_1005,N_2463);
nand U3744 (N_3744,N_1756,N_592);
and U3745 (N_3745,N_278,N_217);
nand U3746 (N_3746,N_2465,N_254);
nor U3747 (N_3747,N_131,N_1283);
and U3748 (N_3748,N_2250,N_2383);
and U3749 (N_3749,N_1523,N_302);
nor U3750 (N_3750,N_1197,N_788);
or U3751 (N_3751,N_909,N_404);
nand U3752 (N_3752,N_653,N_2467);
and U3753 (N_3753,N_1019,N_1711);
and U3754 (N_3754,N_77,N_953);
nor U3755 (N_3755,N_2177,N_50);
and U3756 (N_3756,N_108,N_976);
and U3757 (N_3757,N_1238,N_1882);
nand U3758 (N_3758,N_1047,N_1881);
and U3759 (N_3759,N_1524,N_999);
and U3760 (N_3760,N_2229,N_850);
nand U3761 (N_3761,N_145,N_647);
and U3762 (N_3762,N_911,N_2141);
and U3763 (N_3763,N_915,N_1870);
nand U3764 (N_3764,N_1191,N_2339);
and U3765 (N_3765,N_467,N_1866);
nor U3766 (N_3766,N_1019,N_916);
and U3767 (N_3767,N_2085,N_42);
xor U3768 (N_3768,N_121,N_128);
and U3769 (N_3769,N_2328,N_1218);
nor U3770 (N_3770,N_208,N_1374);
and U3771 (N_3771,N_2404,N_2155);
nor U3772 (N_3772,N_1203,N_1560);
or U3773 (N_3773,N_350,N_1801);
nand U3774 (N_3774,N_2072,N_915);
nand U3775 (N_3775,N_761,N_1315);
nand U3776 (N_3776,N_1494,N_477);
and U3777 (N_3777,N_565,N_25);
or U3778 (N_3778,N_911,N_2320);
or U3779 (N_3779,N_1885,N_859);
or U3780 (N_3780,N_2315,N_1654);
nand U3781 (N_3781,N_1974,N_629);
nand U3782 (N_3782,N_1827,N_37);
nand U3783 (N_3783,N_5,N_2131);
or U3784 (N_3784,N_10,N_86);
and U3785 (N_3785,N_1812,N_2270);
and U3786 (N_3786,N_1504,N_1231);
or U3787 (N_3787,N_423,N_458);
or U3788 (N_3788,N_892,N_27);
nand U3789 (N_3789,N_709,N_370);
nand U3790 (N_3790,N_1427,N_702);
nor U3791 (N_3791,N_1489,N_1595);
or U3792 (N_3792,N_545,N_822);
nor U3793 (N_3793,N_50,N_67);
nand U3794 (N_3794,N_1319,N_2190);
nor U3795 (N_3795,N_511,N_1580);
nand U3796 (N_3796,N_41,N_549);
nor U3797 (N_3797,N_146,N_1498);
nand U3798 (N_3798,N_828,N_2322);
and U3799 (N_3799,N_1477,N_1082);
or U3800 (N_3800,N_1089,N_408);
or U3801 (N_3801,N_1960,N_219);
xor U3802 (N_3802,N_2264,N_2400);
nand U3803 (N_3803,N_1313,N_1995);
and U3804 (N_3804,N_1777,N_1511);
or U3805 (N_3805,N_1562,N_1082);
and U3806 (N_3806,N_776,N_1330);
nor U3807 (N_3807,N_1436,N_699);
and U3808 (N_3808,N_907,N_1008);
nor U3809 (N_3809,N_239,N_2034);
nor U3810 (N_3810,N_302,N_1);
nand U3811 (N_3811,N_181,N_173);
and U3812 (N_3812,N_1310,N_1965);
and U3813 (N_3813,N_1483,N_1039);
nand U3814 (N_3814,N_504,N_1164);
nand U3815 (N_3815,N_1910,N_611);
nand U3816 (N_3816,N_1314,N_2066);
nand U3817 (N_3817,N_516,N_1183);
or U3818 (N_3818,N_1453,N_2203);
nand U3819 (N_3819,N_944,N_2462);
xor U3820 (N_3820,N_908,N_981);
nor U3821 (N_3821,N_1036,N_1821);
nor U3822 (N_3822,N_1030,N_439);
nand U3823 (N_3823,N_2445,N_1024);
nor U3824 (N_3824,N_2271,N_2151);
nand U3825 (N_3825,N_680,N_2269);
and U3826 (N_3826,N_319,N_124);
nand U3827 (N_3827,N_1488,N_2473);
nor U3828 (N_3828,N_1234,N_2231);
nor U3829 (N_3829,N_1514,N_2363);
nand U3830 (N_3830,N_2313,N_2478);
xor U3831 (N_3831,N_2110,N_1873);
or U3832 (N_3832,N_495,N_729);
nand U3833 (N_3833,N_2243,N_913);
and U3834 (N_3834,N_1248,N_383);
or U3835 (N_3835,N_2485,N_1755);
nor U3836 (N_3836,N_1899,N_1267);
nor U3837 (N_3837,N_612,N_1666);
xnor U3838 (N_3838,N_2060,N_1260);
and U3839 (N_3839,N_1304,N_1569);
and U3840 (N_3840,N_2206,N_82);
nor U3841 (N_3841,N_61,N_877);
nor U3842 (N_3842,N_1152,N_1901);
and U3843 (N_3843,N_978,N_536);
and U3844 (N_3844,N_1221,N_642);
nor U3845 (N_3845,N_1837,N_918);
and U3846 (N_3846,N_1503,N_87);
or U3847 (N_3847,N_1501,N_1216);
nor U3848 (N_3848,N_345,N_1167);
or U3849 (N_3849,N_1729,N_1024);
nor U3850 (N_3850,N_147,N_1496);
nor U3851 (N_3851,N_1304,N_742);
nand U3852 (N_3852,N_1055,N_1178);
nor U3853 (N_3853,N_695,N_1788);
nor U3854 (N_3854,N_2261,N_2015);
or U3855 (N_3855,N_1723,N_1630);
nand U3856 (N_3856,N_2202,N_2407);
xor U3857 (N_3857,N_1041,N_1415);
or U3858 (N_3858,N_2372,N_1294);
or U3859 (N_3859,N_2170,N_1911);
and U3860 (N_3860,N_1288,N_120);
nand U3861 (N_3861,N_740,N_1682);
nor U3862 (N_3862,N_1886,N_712);
nor U3863 (N_3863,N_1609,N_30);
nor U3864 (N_3864,N_229,N_431);
and U3865 (N_3865,N_490,N_765);
nand U3866 (N_3866,N_655,N_2101);
nor U3867 (N_3867,N_1065,N_1021);
and U3868 (N_3868,N_2034,N_1268);
nor U3869 (N_3869,N_1523,N_2055);
nand U3870 (N_3870,N_1338,N_243);
or U3871 (N_3871,N_2479,N_1442);
or U3872 (N_3872,N_1964,N_2225);
nor U3873 (N_3873,N_707,N_1343);
nand U3874 (N_3874,N_1844,N_565);
and U3875 (N_3875,N_442,N_2088);
nor U3876 (N_3876,N_644,N_2185);
nor U3877 (N_3877,N_1380,N_2237);
nor U3878 (N_3878,N_2197,N_2260);
or U3879 (N_3879,N_292,N_2086);
nor U3880 (N_3880,N_2021,N_2375);
nand U3881 (N_3881,N_1928,N_965);
nor U3882 (N_3882,N_1911,N_939);
nor U3883 (N_3883,N_2450,N_1980);
or U3884 (N_3884,N_836,N_1184);
or U3885 (N_3885,N_1414,N_651);
or U3886 (N_3886,N_639,N_512);
and U3887 (N_3887,N_2358,N_99);
nor U3888 (N_3888,N_834,N_1695);
nor U3889 (N_3889,N_532,N_681);
nand U3890 (N_3890,N_1744,N_642);
nor U3891 (N_3891,N_1604,N_558);
and U3892 (N_3892,N_1001,N_543);
nor U3893 (N_3893,N_2025,N_1088);
or U3894 (N_3894,N_135,N_2099);
or U3895 (N_3895,N_2313,N_611);
and U3896 (N_3896,N_1037,N_1171);
or U3897 (N_3897,N_571,N_121);
or U3898 (N_3898,N_1817,N_338);
nand U3899 (N_3899,N_924,N_1416);
nand U3900 (N_3900,N_1489,N_1668);
nand U3901 (N_3901,N_399,N_119);
and U3902 (N_3902,N_1231,N_2021);
nand U3903 (N_3903,N_2421,N_357);
and U3904 (N_3904,N_2309,N_1842);
nand U3905 (N_3905,N_234,N_794);
nor U3906 (N_3906,N_397,N_841);
nor U3907 (N_3907,N_1313,N_2337);
or U3908 (N_3908,N_784,N_1079);
nand U3909 (N_3909,N_764,N_412);
and U3910 (N_3910,N_1490,N_66);
nand U3911 (N_3911,N_2179,N_732);
and U3912 (N_3912,N_78,N_81);
nor U3913 (N_3913,N_2165,N_1734);
nand U3914 (N_3914,N_469,N_582);
and U3915 (N_3915,N_1696,N_2364);
or U3916 (N_3916,N_465,N_2139);
nand U3917 (N_3917,N_1346,N_1795);
or U3918 (N_3918,N_1357,N_1870);
or U3919 (N_3919,N_143,N_761);
and U3920 (N_3920,N_2403,N_940);
or U3921 (N_3921,N_664,N_1794);
and U3922 (N_3922,N_526,N_1957);
and U3923 (N_3923,N_2117,N_236);
nor U3924 (N_3924,N_1205,N_1401);
and U3925 (N_3925,N_1653,N_1985);
nand U3926 (N_3926,N_2133,N_1997);
or U3927 (N_3927,N_2465,N_1921);
and U3928 (N_3928,N_2415,N_1148);
or U3929 (N_3929,N_1095,N_1446);
nand U3930 (N_3930,N_62,N_280);
xnor U3931 (N_3931,N_1230,N_1704);
and U3932 (N_3932,N_2005,N_1486);
and U3933 (N_3933,N_2,N_1455);
nand U3934 (N_3934,N_1494,N_2285);
nor U3935 (N_3935,N_1384,N_2387);
and U3936 (N_3936,N_2407,N_498);
or U3937 (N_3937,N_1024,N_234);
and U3938 (N_3938,N_911,N_838);
or U3939 (N_3939,N_833,N_2173);
and U3940 (N_3940,N_2083,N_1853);
nor U3941 (N_3941,N_1602,N_1684);
or U3942 (N_3942,N_56,N_769);
or U3943 (N_3943,N_814,N_156);
or U3944 (N_3944,N_494,N_1411);
nand U3945 (N_3945,N_2139,N_1650);
or U3946 (N_3946,N_1862,N_465);
nor U3947 (N_3947,N_1234,N_154);
nand U3948 (N_3948,N_1867,N_2291);
or U3949 (N_3949,N_2477,N_309);
and U3950 (N_3950,N_558,N_1417);
nand U3951 (N_3951,N_1413,N_967);
and U3952 (N_3952,N_1677,N_1891);
nand U3953 (N_3953,N_2160,N_1753);
and U3954 (N_3954,N_2136,N_578);
and U3955 (N_3955,N_338,N_269);
nor U3956 (N_3956,N_1003,N_125);
and U3957 (N_3957,N_424,N_1181);
nand U3958 (N_3958,N_1154,N_935);
and U3959 (N_3959,N_2143,N_1779);
and U3960 (N_3960,N_806,N_650);
or U3961 (N_3961,N_580,N_64);
nor U3962 (N_3962,N_172,N_1023);
and U3963 (N_3963,N_1240,N_628);
nor U3964 (N_3964,N_1626,N_583);
nand U3965 (N_3965,N_1979,N_221);
nor U3966 (N_3966,N_1342,N_300);
and U3967 (N_3967,N_846,N_1647);
nor U3968 (N_3968,N_268,N_2467);
nor U3969 (N_3969,N_1679,N_2490);
nor U3970 (N_3970,N_2075,N_1879);
or U3971 (N_3971,N_500,N_2174);
nand U3972 (N_3972,N_1377,N_1773);
nand U3973 (N_3973,N_1836,N_100);
nor U3974 (N_3974,N_2199,N_199);
and U3975 (N_3975,N_2081,N_903);
nor U3976 (N_3976,N_318,N_423);
nor U3977 (N_3977,N_738,N_1173);
and U3978 (N_3978,N_878,N_1484);
nand U3979 (N_3979,N_1020,N_741);
and U3980 (N_3980,N_1661,N_1461);
and U3981 (N_3981,N_1581,N_1719);
nor U3982 (N_3982,N_2294,N_1918);
nor U3983 (N_3983,N_2058,N_2476);
nand U3984 (N_3984,N_2149,N_1455);
and U3985 (N_3985,N_2084,N_2032);
and U3986 (N_3986,N_243,N_185);
xnor U3987 (N_3987,N_1737,N_1849);
or U3988 (N_3988,N_621,N_908);
or U3989 (N_3989,N_1863,N_1647);
or U3990 (N_3990,N_1342,N_2082);
nand U3991 (N_3991,N_1541,N_63);
nor U3992 (N_3992,N_1583,N_2015);
or U3993 (N_3993,N_444,N_1522);
or U3994 (N_3994,N_2,N_1294);
nand U3995 (N_3995,N_2170,N_2102);
nand U3996 (N_3996,N_786,N_2084);
nand U3997 (N_3997,N_1599,N_1689);
nand U3998 (N_3998,N_769,N_783);
and U3999 (N_3999,N_276,N_906);
xnor U4000 (N_4000,N_2092,N_671);
nand U4001 (N_4001,N_2365,N_1052);
nand U4002 (N_4002,N_1783,N_2414);
nand U4003 (N_4003,N_352,N_1164);
nand U4004 (N_4004,N_1877,N_2065);
nor U4005 (N_4005,N_1136,N_650);
nand U4006 (N_4006,N_209,N_2076);
nor U4007 (N_4007,N_1461,N_882);
nand U4008 (N_4008,N_1917,N_716);
nand U4009 (N_4009,N_2091,N_1598);
nor U4010 (N_4010,N_2483,N_1473);
nand U4011 (N_4011,N_2186,N_1422);
nand U4012 (N_4012,N_1180,N_458);
and U4013 (N_4013,N_1004,N_1690);
nor U4014 (N_4014,N_804,N_680);
nor U4015 (N_4015,N_2072,N_1164);
nand U4016 (N_4016,N_1616,N_951);
or U4017 (N_4017,N_1988,N_1917);
and U4018 (N_4018,N_1723,N_11);
nand U4019 (N_4019,N_1652,N_776);
or U4020 (N_4020,N_1486,N_898);
nand U4021 (N_4021,N_1030,N_1336);
or U4022 (N_4022,N_2029,N_663);
or U4023 (N_4023,N_1256,N_1812);
nor U4024 (N_4024,N_439,N_1403);
nor U4025 (N_4025,N_1828,N_519);
and U4026 (N_4026,N_367,N_262);
or U4027 (N_4027,N_152,N_773);
nor U4028 (N_4028,N_2311,N_2415);
nand U4029 (N_4029,N_1289,N_1116);
nand U4030 (N_4030,N_259,N_357);
nand U4031 (N_4031,N_285,N_885);
or U4032 (N_4032,N_2013,N_2318);
and U4033 (N_4033,N_874,N_2183);
and U4034 (N_4034,N_810,N_804);
nor U4035 (N_4035,N_1290,N_888);
or U4036 (N_4036,N_1838,N_1747);
or U4037 (N_4037,N_7,N_1742);
and U4038 (N_4038,N_512,N_1310);
and U4039 (N_4039,N_2127,N_1190);
or U4040 (N_4040,N_1842,N_1623);
nor U4041 (N_4041,N_1408,N_923);
nor U4042 (N_4042,N_1476,N_1954);
or U4043 (N_4043,N_1172,N_573);
nor U4044 (N_4044,N_2447,N_1815);
and U4045 (N_4045,N_1933,N_595);
and U4046 (N_4046,N_993,N_755);
nor U4047 (N_4047,N_2,N_1709);
nand U4048 (N_4048,N_1788,N_52);
nor U4049 (N_4049,N_1055,N_2440);
nor U4050 (N_4050,N_4,N_644);
nor U4051 (N_4051,N_1309,N_508);
and U4052 (N_4052,N_2260,N_1402);
nand U4053 (N_4053,N_2363,N_2229);
or U4054 (N_4054,N_758,N_1408);
nand U4055 (N_4055,N_981,N_588);
xnor U4056 (N_4056,N_2045,N_1502);
or U4057 (N_4057,N_1008,N_726);
and U4058 (N_4058,N_200,N_2069);
or U4059 (N_4059,N_0,N_988);
and U4060 (N_4060,N_969,N_569);
nor U4061 (N_4061,N_832,N_1072);
nand U4062 (N_4062,N_1094,N_1926);
and U4063 (N_4063,N_1354,N_515);
nor U4064 (N_4064,N_518,N_2195);
nor U4065 (N_4065,N_294,N_1644);
and U4066 (N_4066,N_776,N_554);
and U4067 (N_4067,N_1282,N_518);
xnor U4068 (N_4068,N_368,N_1653);
or U4069 (N_4069,N_2412,N_698);
or U4070 (N_4070,N_478,N_2337);
nand U4071 (N_4071,N_2002,N_1844);
and U4072 (N_4072,N_2049,N_2092);
or U4073 (N_4073,N_1781,N_1753);
nor U4074 (N_4074,N_1217,N_2142);
nor U4075 (N_4075,N_2423,N_784);
or U4076 (N_4076,N_1072,N_2345);
nor U4077 (N_4077,N_1835,N_198);
and U4078 (N_4078,N_475,N_1856);
nand U4079 (N_4079,N_1259,N_1965);
nor U4080 (N_4080,N_204,N_2342);
or U4081 (N_4081,N_421,N_2198);
nand U4082 (N_4082,N_127,N_1134);
and U4083 (N_4083,N_1152,N_2470);
and U4084 (N_4084,N_1563,N_162);
nor U4085 (N_4085,N_2250,N_1965);
and U4086 (N_4086,N_2344,N_983);
nor U4087 (N_4087,N_2163,N_305);
and U4088 (N_4088,N_1132,N_1077);
nand U4089 (N_4089,N_2407,N_1015);
nand U4090 (N_4090,N_1017,N_1990);
nor U4091 (N_4091,N_1891,N_1436);
and U4092 (N_4092,N_919,N_793);
or U4093 (N_4093,N_2142,N_2108);
and U4094 (N_4094,N_1204,N_1693);
xor U4095 (N_4095,N_1787,N_1342);
nor U4096 (N_4096,N_833,N_2467);
nand U4097 (N_4097,N_1057,N_499);
nor U4098 (N_4098,N_1883,N_167);
and U4099 (N_4099,N_254,N_848);
xor U4100 (N_4100,N_13,N_1523);
or U4101 (N_4101,N_48,N_1041);
and U4102 (N_4102,N_1738,N_1220);
nor U4103 (N_4103,N_929,N_1869);
nand U4104 (N_4104,N_2448,N_947);
and U4105 (N_4105,N_1852,N_352);
nor U4106 (N_4106,N_385,N_579);
and U4107 (N_4107,N_487,N_58);
and U4108 (N_4108,N_887,N_1635);
nand U4109 (N_4109,N_1448,N_2296);
nor U4110 (N_4110,N_1632,N_2154);
and U4111 (N_4111,N_10,N_941);
and U4112 (N_4112,N_1407,N_2305);
or U4113 (N_4113,N_1614,N_1956);
xnor U4114 (N_4114,N_793,N_2449);
nor U4115 (N_4115,N_816,N_2356);
xor U4116 (N_4116,N_2203,N_263);
or U4117 (N_4117,N_829,N_283);
or U4118 (N_4118,N_1284,N_1175);
nor U4119 (N_4119,N_1819,N_455);
nor U4120 (N_4120,N_2442,N_1008);
and U4121 (N_4121,N_1926,N_603);
nand U4122 (N_4122,N_1539,N_496);
or U4123 (N_4123,N_2439,N_392);
and U4124 (N_4124,N_1661,N_1412);
or U4125 (N_4125,N_93,N_1286);
and U4126 (N_4126,N_1709,N_330);
and U4127 (N_4127,N_2470,N_240);
or U4128 (N_4128,N_715,N_2252);
or U4129 (N_4129,N_665,N_1162);
nand U4130 (N_4130,N_2327,N_535);
and U4131 (N_4131,N_1038,N_1663);
nand U4132 (N_4132,N_804,N_1536);
nor U4133 (N_4133,N_1116,N_10);
nand U4134 (N_4134,N_588,N_12);
nand U4135 (N_4135,N_493,N_2146);
and U4136 (N_4136,N_1082,N_2443);
and U4137 (N_4137,N_1337,N_2021);
or U4138 (N_4138,N_1191,N_1272);
nor U4139 (N_4139,N_1809,N_1851);
nand U4140 (N_4140,N_2450,N_873);
or U4141 (N_4141,N_612,N_2487);
or U4142 (N_4142,N_1136,N_2267);
and U4143 (N_4143,N_675,N_1948);
xor U4144 (N_4144,N_789,N_417);
nand U4145 (N_4145,N_2158,N_952);
xor U4146 (N_4146,N_176,N_2020);
nand U4147 (N_4147,N_130,N_34);
and U4148 (N_4148,N_1392,N_1939);
xor U4149 (N_4149,N_916,N_547);
or U4150 (N_4150,N_852,N_1401);
nand U4151 (N_4151,N_688,N_1520);
or U4152 (N_4152,N_2286,N_2256);
or U4153 (N_4153,N_1738,N_447);
and U4154 (N_4154,N_291,N_1607);
nand U4155 (N_4155,N_2154,N_1558);
nand U4156 (N_4156,N_1982,N_1585);
nand U4157 (N_4157,N_1736,N_84);
and U4158 (N_4158,N_735,N_1954);
and U4159 (N_4159,N_2211,N_1391);
nor U4160 (N_4160,N_480,N_271);
or U4161 (N_4161,N_835,N_565);
and U4162 (N_4162,N_1915,N_1741);
nor U4163 (N_4163,N_1391,N_856);
or U4164 (N_4164,N_54,N_2203);
and U4165 (N_4165,N_358,N_1904);
nand U4166 (N_4166,N_1440,N_1550);
and U4167 (N_4167,N_2489,N_121);
nand U4168 (N_4168,N_1506,N_260);
nor U4169 (N_4169,N_2485,N_799);
nand U4170 (N_4170,N_973,N_2401);
and U4171 (N_4171,N_1815,N_2263);
nand U4172 (N_4172,N_405,N_247);
and U4173 (N_4173,N_275,N_553);
nand U4174 (N_4174,N_560,N_951);
and U4175 (N_4175,N_1299,N_751);
and U4176 (N_4176,N_1424,N_846);
and U4177 (N_4177,N_212,N_342);
and U4178 (N_4178,N_1248,N_525);
nor U4179 (N_4179,N_190,N_1337);
or U4180 (N_4180,N_47,N_1550);
nand U4181 (N_4181,N_846,N_477);
or U4182 (N_4182,N_247,N_1554);
nand U4183 (N_4183,N_1849,N_335);
nand U4184 (N_4184,N_2325,N_748);
and U4185 (N_4185,N_905,N_84);
nand U4186 (N_4186,N_766,N_1557);
and U4187 (N_4187,N_1544,N_905);
nand U4188 (N_4188,N_1336,N_1179);
or U4189 (N_4189,N_2088,N_1474);
nand U4190 (N_4190,N_2133,N_1120);
and U4191 (N_4191,N_1183,N_1494);
and U4192 (N_4192,N_2491,N_1533);
nor U4193 (N_4193,N_1886,N_1172);
or U4194 (N_4194,N_774,N_811);
nor U4195 (N_4195,N_2221,N_608);
nand U4196 (N_4196,N_532,N_1302);
and U4197 (N_4197,N_2324,N_635);
nor U4198 (N_4198,N_2041,N_1926);
nand U4199 (N_4199,N_2357,N_393);
nand U4200 (N_4200,N_146,N_2296);
and U4201 (N_4201,N_725,N_2163);
and U4202 (N_4202,N_494,N_1726);
nor U4203 (N_4203,N_905,N_996);
nand U4204 (N_4204,N_1307,N_44);
or U4205 (N_4205,N_1371,N_171);
or U4206 (N_4206,N_787,N_322);
and U4207 (N_4207,N_1406,N_1317);
nand U4208 (N_4208,N_1726,N_2461);
nand U4209 (N_4209,N_1708,N_715);
or U4210 (N_4210,N_2151,N_2490);
and U4211 (N_4211,N_641,N_1116);
and U4212 (N_4212,N_150,N_2372);
nand U4213 (N_4213,N_1009,N_2007);
and U4214 (N_4214,N_1742,N_1663);
nor U4215 (N_4215,N_692,N_1267);
and U4216 (N_4216,N_2095,N_1243);
nand U4217 (N_4217,N_1511,N_1146);
and U4218 (N_4218,N_1902,N_942);
and U4219 (N_4219,N_130,N_1006);
or U4220 (N_4220,N_63,N_1814);
nand U4221 (N_4221,N_1298,N_2245);
or U4222 (N_4222,N_1244,N_1286);
xor U4223 (N_4223,N_589,N_175);
nor U4224 (N_4224,N_1242,N_731);
and U4225 (N_4225,N_2389,N_1373);
nand U4226 (N_4226,N_268,N_2062);
xnor U4227 (N_4227,N_2414,N_1541);
or U4228 (N_4228,N_2331,N_2338);
nor U4229 (N_4229,N_1188,N_1945);
nor U4230 (N_4230,N_2076,N_946);
and U4231 (N_4231,N_718,N_2046);
or U4232 (N_4232,N_2183,N_517);
nand U4233 (N_4233,N_2086,N_1929);
nand U4234 (N_4234,N_786,N_2169);
nand U4235 (N_4235,N_1971,N_1549);
nand U4236 (N_4236,N_2470,N_46);
and U4237 (N_4237,N_378,N_1713);
xor U4238 (N_4238,N_2308,N_334);
nand U4239 (N_4239,N_2174,N_223);
nand U4240 (N_4240,N_1223,N_1231);
or U4241 (N_4241,N_2200,N_991);
xnor U4242 (N_4242,N_2035,N_2008);
or U4243 (N_4243,N_1801,N_952);
or U4244 (N_4244,N_370,N_1948);
or U4245 (N_4245,N_1715,N_1387);
or U4246 (N_4246,N_1036,N_1724);
and U4247 (N_4247,N_1661,N_247);
nor U4248 (N_4248,N_2255,N_1788);
nor U4249 (N_4249,N_480,N_1677);
nor U4250 (N_4250,N_1835,N_1796);
and U4251 (N_4251,N_150,N_369);
or U4252 (N_4252,N_2467,N_1352);
or U4253 (N_4253,N_916,N_2349);
or U4254 (N_4254,N_1910,N_1210);
nand U4255 (N_4255,N_526,N_475);
or U4256 (N_4256,N_472,N_1282);
xnor U4257 (N_4257,N_1907,N_1766);
and U4258 (N_4258,N_2012,N_2439);
nor U4259 (N_4259,N_76,N_423);
nor U4260 (N_4260,N_693,N_1008);
nor U4261 (N_4261,N_2032,N_1056);
nor U4262 (N_4262,N_1721,N_2371);
and U4263 (N_4263,N_712,N_97);
or U4264 (N_4264,N_1605,N_717);
xor U4265 (N_4265,N_1034,N_1617);
nand U4266 (N_4266,N_265,N_530);
and U4267 (N_4267,N_347,N_1667);
nand U4268 (N_4268,N_916,N_1808);
and U4269 (N_4269,N_212,N_1761);
nand U4270 (N_4270,N_442,N_147);
and U4271 (N_4271,N_435,N_2187);
or U4272 (N_4272,N_451,N_1928);
and U4273 (N_4273,N_1538,N_31);
nor U4274 (N_4274,N_678,N_1499);
nand U4275 (N_4275,N_1322,N_591);
nand U4276 (N_4276,N_315,N_580);
nand U4277 (N_4277,N_453,N_426);
and U4278 (N_4278,N_1950,N_1847);
nand U4279 (N_4279,N_1762,N_1703);
and U4280 (N_4280,N_1691,N_1841);
or U4281 (N_4281,N_1373,N_2403);
or U4282 (N_4282,N_421,N_1877);
nor U4283 (N_4283,N_1458,N_2075);
and U4284 (N_4284,N_2016,N_506);
and U4285 (N_4285,N_2172,N_1987);
or U4286 (N_4286,N_500,N_923);
nor U4287 (N_4287,N_1933,N_1396);
nand U4288 (N_4288,N_2346,N_1331);
nand U4289 (N_4289,N_2232,N_1911);
and U4290 (N_4290,N_2301,N_2323);
nor U4291 (N_4291,N_1379,N_876);
xor U4292 (N_4292,N_859,N_1399);
nor U4293 (N_4293,N_322,N_1213);
nor U4294 (N_4294,N_1877,N_2046);
or U4295 (N_4295,N_212,N_537);
and U4296 (N_4296,N_2019,N_897);
or U4297 (N_4297,N_1941,N_1213);
nand U4298 (N_4298,N_1516,N_1428);
nor U4299 (N_4299,N_1592,N_2122);
xnor U4300 (N_4300,N_239,N_144);
or U4301 (N_4301,N_2244,N_825);
nor U4302 (N_4302,N_2184,N_2245);
nand U4303 (N_4303,N_730,N_2283);
nor U4304 (N_4304,N_413,N_791);
nand U4305 (N_4305,N_866,N_2151);
nor U4306 (N_4306,N_1310,N_134);
and U4307 (N_4307,N_1637,N_1109);
nor U4308 (N_4308,N_1513,N_2475);
and U4309 (N_4309,N_297,N_1807);
and U4310 (N_4310,N_1258,N_2245);
nand U4311 (N_4311,N_362,N_1945);
or U4312 (N_4312,N_1486,N_1105);
or U4313 (N_4313,N_1250,N_1570);
and U4314 (N_4314,N_1891,N_2360);
or U4315 (N_4315,N_1442,N_1548);
and U4316 (N_4316,N_440,N_2281);
and U4317 (N_4317,N_1264,N_610);
and U4318 (N_4318,N_2363,N_1511);
xnor U4319 (N_4319,N_612,N_224);
nand U4320 (N_4320,N_40,N_812);
nor U4321 (N_4321,N_1175,N_983);
and U4322 (N_4322,N_2272,N_1157);
or U4323 (N_4323,N_2373,N_1490);
nor U4324 (N_4324,N_267,N_284);
nand U4325 (N_4325,N_1667,N_2053);
nor U4326 (N_4326,N_643,N_2204);
and U4327 (N_4327,N_1771,N_2358);
or U4328 (N_4328,N_2376,N_292);
and U4329 (N_4329,N_1797,N_1919);
or U4330 (N_4330,N_1639,N_1297);
xor U4331 (N_4331,N_860,N_154);
nand U4332 (N_4332,N_1981,N_767);
xor U4333 (N_4333,N_1788,N_1563);
and U4334 (N_4334,N_2356,N_2304);
or U4335 (N_4335,N_1229,N_2490);
and U4336 (N_4336,N_684,N_606);
nand U4337 (N_4337,N_1412,N_871);
nand U4338 (N_4338,N_1195,N_2119);
nand U4339 (N_4339,N_514,N_690);
and U4340 (N_4340,N_820,N_649);
nand U4341 (N_4341,N_1755,N_2306);
and U4342 (N_4342,N_2423,N_2456);
nor U4343 (N_4343,N_372,N_1549);
and U4344 (N_4344,N_1355,N_437);
or U4345 (N_4345,N_2299,N_1694);
nand U4346 (N_4346,N_408,N_2032);
nor U4347 (N_4347,N_1339,N_955);
nor U4348 (N_4348,N_2390,N_12);
nor U4349 (N_4349,N_484,N_599);
nor U4350 (N_4350,N_1268,N_2352);
and U4351 (N_4351,N_1163,N_516);
and U4352 (N_4352,N_2447,N_124);
or U4353 (N_4353,N_1097,N_2040);
nand U4354 (N_4354,N_577,N_709);
or U4355 (N_4355,N_2031,N_334);
nor U4356 (N_4356,N_1604,N_191);
or U4357 (N_4357,N_455,N_2438);
nand U4358 (N_4358,N_1704,N_1393);
and U4359 (N_4359,N_1569,N_686);
or U4360 (N_4360,N_2381,N_1484);
nand U4361 (N_4361,N_1383,N_1651);
and U4362 (N_4362,N_1648,N_682);
or U4363 (N_4363,N_1129,N_354);
or U4364 (N_4364,N_1104,N_2372);
nand U4365 (N_4365,N_2105,N_523);
nor U4366 (N_4366,N_2016,N_1147);
and U4367 (N_4367,N_1231,N_1593);
nor U4368 (N_4368,N_1764,N_194);
and U4369 (N_4369,N_141,N_1685);
or U4370 (N_4370,N_798,N_1588);
or U4371 (N_4371,N_1769,N_1448);
and U4372 (N_4372,N_1907,N_1208);
and U4373 (N_4373,N_1483,N_1330);
nand U4374 (N_4374,N_2407,N_234);
and U4375 (N_4375,N_2102,N_551);
and U4376 (N_4376,N_1974,N_1491);
and U4377 (N_4377,N_2242,N_1848);
and U4378 (N_4378,N_1178,N_2122);
nor U4379 (N_4379,N_1357,N_1732);
and U4380 (N_4380,N_2303,N_475);
nand U4381 (N_4381,N_1681,N_1252);
or U4382 (N_4382,N_819,N_637);
nor U4383 (N_4383,N_1654,N_1594);
nor U4384 (N_4384,N_2077,N_1515);
nand U4385 (N_4385,N_2216,N_1546);
or U4386 (N_4386,N_1255,N_2277);
nand U4387 (N_4387,N_124,N_1032);
or U4388 (N_4388,N_1516,N_1062);
and U4389 (N_4389,N_130,N_2478);
or U4390 (N_4390,N_114,N_1164);
or U4391 (N_4391,N_1311,N_574);
and U4392 (N_4392,N_2184,N_1692);
nand U4393 (N_4393,N_281,N_659);
and U4394 (N_4394,N_1345,N_1219);
and U4395 (N_4395,N_218,N_1672);
and U4396 (N_4396,N_2498,N_747);
and U4397 (N_4397,N_1647,N_820);
nor U4398 (N_4398,N_1476,N_1658);
nor U4399 (N_4399,N_1593,N_1952);
nor U4400 (N_4400,N_8,N_1379);
nand U4401 (N_4401,N_2246,N_1297);
or U4402 (N_4402,N_2315,N_607);
nand U4403 (N_4403,N_15,N_1504);
and U4404 (N_4404,N_1906,N_2);
nand U4405 (N_4405,N_2410,N_920);
nor U4406 (N_4406,N_1523,N_25);
nor U4407 (N_4407,N_2406,N_1783);
nand U4408 (N_4408,N_2193,N_2408);
nor U4409 (N_4409,N_129,N_745);
or U4410 (N_4410,N_1535,N_396);
or U4411 (N_4411,N_481,N_2191);
or U4412 (N_4412,N_419,N_678);
nor U4413 (N_4413,N_226,N_903);
or U4414 (N_4414,N_1846,N_2222);
nor U4415 (N_4415,N_899,N_2357);
nand U4416 (N_4416,N_1233,N_127);
nand U4417 (N_4417,N_183,N_2335);
or U4418 (N_4418,N_2439,N_1711);
nand U4419 (N_4419,N_61,N_11);
and U4420 (N_4420,N_2386,N_701);
nand U4421 (N_4421,N_961,N_508);
or U4422 (N_4422,N_921,N_1651);
and U4423 (N_4423,N_2184,N_2378);
nand U4424 (N_4424,N_270,N_1468);
and U4425 (N_4425,N_1675,N_215);
or U4426 (N_4426,N_574,N_1565);
or U4427 (N_4427,N_1035,N_1656);
nor U4428 (N_4428,N_188,N_918);
nor U4429 (N_4429,N_1311,N_1243);
or U4430 (N_4430,N_1165,N_261);
nand U4431 (N_4431,N_290,N_2108);
or U4432 (N_4432,N_2118,N_430);
or U4433 (N_4433,N_2120,N_2287);
nor U4434 (N_4434,N_1670,N_1939);
nand U4435 (N_4435,N_812,N_1547);
nor U4436 (N_4436,N_1843,N_1649);
or U4437 (N_4437,N_1637,N_42);
nor U4438 (N_4438,N_1151,N_2049);
nand U4439 (N_4439,N_2124,N_1475);
or U4440 (N_4440,N_1711,N_1488);
or U4441 (N_4441,N_2052,N_891);
nor U4442 (N_4442,N_414,N_2154);
nor U4443 (N_4443,N_555,N_2349);
and U4444 (N_4444,N_745,N_1726);
or U4445 (N_4445,N_1170,N_477);
nand U4446 (N_4446,N_1733,N_2478);
nor U4447 (N_4447,N_1328,N_716);
nand U4448 (N_4448,N_2471,N_395);
and U4449 (N_4449,N_656,N_2441);
nand U4450 (N_4450,N_1643,N_2118);
nor U4451 (N_4451,N_1261,N_866);
or U4452 (N_4452,N_2246,N_2032);
nor U4453 (N_4453,N_1292,N_453);
nand U4454 (N_4454,N_935,N_2045);
and U4455 (N_4455,N_1638,N_1546);
nand U4456 (N_4456,N_436,N_510);
xor U4457 (N_4457,N_1821,N_2401);
or U4458 (N_4458,N_151,N_1886);
nor U4459 (N_4459,N_204,N_1135);
and U4460 (N_4460,N_940,N_695);
nor U4461 (N_4461,N_229,N_1588);
nor U4462 (N_4462,N_27,N_2219);
and U4463 (N_4463,N_1837,N_1891);
or U4464 (N_4464,N_1097,N_2486);
nor U4465 (N_4465,N_737,N_243);
nor U4466 (N_4466,N_809,N_1833);
xnor U4467 (N_4467,N_1458,N_2219);
or U4468 (N_4468,N_1800,N_2046);
or U4469 (N_4469,N_2128,N_1373);
or U4470 (N_4470,N_2068,N_1195);
and U4471 (N_4471,N_840,N_408);
nor U4472 (N_4472,N_800,N_1775);
and U4473 (N_4473,N_1172,N_1889);
and U4474 (N_4474,N_1619,N_1156);
and U4475 (N_4475,N_1399,N_153);
nand U4476 (N_4476,N_1994,N_224);
and U4477 (N_4477,N_180,N_1263);
and U4478 (N_4478,N_1729,N_1254);
nand U4479 (N_4479,N_42,N_34);
and U4480 (N_4480,N_2200,N_1104);
or U4481 (N_4481,N_293,N_1452);
or U4482 (N_4482,N_2398,N_247);
and U4483 (N_4483,N_2041,N_1715);
or U4484 (N_4484,N_413,N_1984);
and U4485 (N_4485,N_1924,N_2008);
and U4486 (N_4486,N_1524,N_590);
and U4487 (N_4487,N_596,N_1851);
nand U4488 (N_4488,N_651,N_1701);
nand U4489 (N_4489,N_756,N_1844);
nor U4490 (N_4490,N_896,N_819);
and U4491 (N_4491,N_2387,N_1229);
nor U4492 (N_4492,N_1169,N_806);
nor U4493 (N_4493,N_2061,N_1713);
nor U4494 (N_4494,N_263,N_427);
nand U4495 (N_4495,N_258,N_81);
and U4496 (N_4496,N_2225,N_21);
and U4497 (N_4497,N_2140,N_999);
and U4498 (N_4498,N_2261,N_1376);
nor U4499 (N_4499,N_1676,N_303);
nand U4500 (N_4500,N_857,N_1743);
nand U4501 (N_4501,N_764,N_1017);
nand U4502 (N_4502,N_1797,N_1393);
nand U4503 (N_4503,N_1273,N_1445);
and U4504 (N_4504,N_2447,N_296);
and U4505 (N_4505,N_167,N_2336);
nand U4506 (N_4506,N_2487,N_1651);
or U4507 (N_4507,N_1516,N_2020);
and U4508 (N_4508,N_1660,N_1640);
or U4509 (N_4509,N_2030,N_941);
and U4510 (N_4510,N_2263,N_2251);
and U4511 (N_4511,N_615,N_1759);
nor U4512 (N_4512,N_1253,N_1808);
nor U4513 (N_4513,N_2012,N_325);
nand U4514 (N_4514,N_1925,N_2095);
nand U4515 (N_4515,N_523,N_1577);
and U4516 (N_4516,N_1157,N_2136);
or U4517 (N_4517,N_964,N_239);
nor U4518 (N_4518,N_1031,N_1105);
xnor U4519 (N_4519,N_1442,N_1415);
and U4520 (N_4520,N_189,N_1171);
nand U4521 (N_4521,N_183,N_1747);
or U4522 (N_4522,N_869,N_81);
and U4523 (N_4523,N_46,N_1761);
or U4524 (N_4524,N_1613,N_223);
nor U4525 (N_4525,N_2375,N_2100);
or U4526 (N_4526,N_1050,N_1899);
nand U4527 (N_4527,N_1672,N_1770);
nand U4528 (N_4528,N_1248,N_2207);
and U4529 (N_4529,N_1622,N_727);
and U4530 (N_4530,N_526,N_1854);
or U4531 (N_4531,N_536,N_1097);
or U4532 (N_4532,N_1652,N_2034);
or U4533 (N_4533,N_1899,N_1401);
xnor U4534 (N_4534,N_1595,N_574);
nor U4535 (N_4535,N_2394,N_1487);
nand U4536 (N_4536,N_2448,N_1250);
nor U4537 (N_4537,N_2154,N_990);
nand U4538 (N_4538,N_86,N_1192);
nand U4539 (N_4539,N_2451,N_107);
and U4540 (N_4540,N_2147,N_2353);
nand U4541 (N_4541,N_860,N_1562);
and U4542 (N_4542,N_1196,N_523);
or U4543 (N_4543,N_2074,N_1717);
nor U4544 (N_4544,N_1635,N_2267);
and U4545 (N_4545,N_376,N_2406);
and U4546 (N_4546,N_570,N_1415);
nor U4547 (N_4547,N_1932,N_2432);
nor U4548 (N_4548,N_2123,N_2364);
nor U4549 (N_4549,N_1586,N_1702);
or U4550 (N_4550,N_1558,N_1895);
or U4551 (N_4551,N_1071,N_1721);
nor U4552 (N_4552,N_402,N_419);
or U4553 (N_4553,N_1916,N_467);
nor U4554 (N_4554,N_1402,N_264);
nor U4555 (N_4555,N_332,N_2385);
and U4556 (N_4556,N_662,N_279);
and U4557 (N_4557,N_863,N_1333);
and U4558 (N_4558,N_1545,N_1889);
or U4559 (N_4559,N_1367,N_2085);
xnor U4560 (N_4560,N_1830,N_1406);
nor U4561 (N_4561,N_1534,N_726);
nand U4562 (N_4562,N_846,N_1066);
or U4563 (N_4563,N_390,N_784);
nor U4564 (N_4564,N_110,N_367);
and U4565 (N_4565,N_1538,N_344);
nor U4566 (N_4566,N_2444,N_929);
nand U4567 (N_4567,N_2058,N_156);
nand U4568 (N_4568,N_1878,N_2219);
nand U4569 (N_4569,N_2065,N_794);
nand U4570 (N_4570,N_318,N_1109);
or U4571 (N_4571,N_975,N_538);
nor U4572 (N_4572,N_1674,N_50);
nand U4573 (N_4573,N_2041,N_610);
nand U4574 (N_4574,N_1639,N_2352);
xnor U4575 (N_4575,N_1865,N_1312);
and U4576 (N_4576,N_1065,N_618);
nor U4577 (N_4577,N_820,N_519);
xnor U4578 (N_4578,N_2063,N_1256);
nor U4579 (N_4579,N_2299,N_1289);
and U4580 (N_4580,N_731,N_2394);
nor U4581 (N_4581,N_2369,N_1156);
or U4582 (N_4582,N_632,N_1166);
or U4583 (N_4583,N_294,N_422);
nor U4584 (N_4584,N_310,N_1929);
and U4585 (N_4585,N_2234,N_2088);
or U4586 (N_4586,N_2194,N_1595);
or U4587 (N_4587,N_2407,N_1323);
and U4588 (N_4588,N_215,N_366);
nor U4589 (N_4589,N_1595,N_586);
or U4590 (N_4590,N_815,N_720);
or U4591 (N_4591,N_1853,N_898);
nor U4592 (N_4592,N_2414,N_478);
nand U4593 (N_4593,N_2258,N_2168);
and U4594 (N_4594,N_213,N_1701);
or U4595 (N_4595,N_718,N_73);
nor U4596 (N_4596,N_1715,N_1724);
nor U4597 (N_4597,N_2306,N_1822);
or U4598 (N_4598,N_2224,N_1392);
xor U4599 (N_4599,N_1507,N_1626);
nor U4600 (N_4600,N_1577,N_1573);
or U4601 (N_4601,N_1428,N_1241);
or U4602 (N_4602,N_2002,N_2009);
and U4603 (N_4603,N_359,N_19);
nor U4604 (N_4604,N_426,N_478);
and U4605 (N_4605,N_1766,N_1200);
nand U4606 (N_4606,N_1678,N_1847);
or U4607 (N_4607,N_2149,N_1397);
and U4608 (N_4608,N_1142,N_824);
nand U4609 (N_4609,N_754,N_934);
and U4610 (N_4610,N_156,N_382);
nor U4611 (N_4611,N_62,N_177);
and U4612 (N_4612,N_151,N_2305);
or U4613 (N_4613,N_267,N_167);
nor U4614 (N_4614,N_1275,N_1317);
nand U4615 (N_4615,N_1840,N_2176);
nor U4616 (N_4616,N_1942,N_1538);
nor U4617 (N_4617,N_1553,N_1389);
and U4618 (N_4618,N_149,N_1997);
and U4619 (N_4619,N_2153,N_1314);
or U4620 (N_4620,N_965,N_2247);
nor U4621 (N_4621,N_1259,N_2371);
nand U4622 (N_4622,N_2406,N_958);
nand U4623 (N_4623,N_2147,N_1599);
nand U4624 (N_4624,N_705,N_1307);
and U4625 (N_4625,N_806,N_392);
nor U4626 (N_4626,N_1012,N_1334);
xnor U4627 (N_4627,N_1791,N_519);
nand U4628 (N_4628,N_2222,N_2099);
and U4629 (N_4629,N_1699,N_1447);
nor U4630 (N_4630,N_1224,N_88);
nand U4631 (N_4631,N_2265,N_2124);
xor U4632 (N_4632,N_760,N_2037);
nor U4633 (N_4633,N_1642,N_424);
and U4634 (N_4634,N_1667,N_221);
nand U4635 (N_4635,N_1754,N_1449);
and U4636 (N_4636,N_538,N_256);
nand U4637 (N_4637,N_1801,N_2135);
nand U4638 (N_4638,N_1616,N_1053);
or U4639 (N_4639,N_800,N_44);
or U4640 (N_4640,N_962,N_516);
nand U4641 (N_4641,N_1832,N_1091);
nand U4642 (N_4642,N_1842,N_1695);
nand U4643 (N_4643,N_600,N_1324);
or U4644 (N_4644,N_1125,N_2053);
or U4645 (N_4645,N_2342,N_530);
nor U4646 (N_4646,N_1428,N_2055);
and U4647 (N_4647,N_28,N_1352);
or U4648 (N_4648,N_1863,N_2160);
and U4649 (N_4649,N_167,N_2254);
or U4650 (N_4650,N_354,N_544);
or U4651 (N_4651,N_1715,N_1641);
nand U4652 (N_4652,N_864,N_727);
nor U4653 (N_4653,N_789,N_2014);
nor U4654 (N_4654,N_1988,N_1322);
nand U4655 (N_4655,N_1172,N_1410);
and U4656 (N_4656,N_1139,N_1680);
and U4657 (N_4657,N_55,N_2173);
or U4658 (N_4658,N_2481,N_2252);
nor U4659 (N_4659,N_936,N_340);
nor U4660 (N_4660,N_1028,N_156);
xnor U4661 (N_4661,N_1798,N_2265);
or U4662 (N_4662,N_771,N_1101);
nand U4663 (N_4663,N_21,N_2068);
nand U4664 (N_4664,N_711,N_238);
and U4665 (N_4665,N_2253,N_1815);
nor U4666 (N_4666,N_244,N_443);
nor U4667 (N_4667,N_272,N_878);
nand U4668 (N_4668,N_2456,N_1725);
nand U4669 (N_4669,N_2090,N_1000);
nand U4670 (N_4670,N_2084,N_2357);
nor U4671 (N_4671,N_1960,N_1005);
or U4672 (N_4672,N_816,N_1548);
nor U4673 (N_4673,N_916,N_754);
nand U4674 (N_4674,N_1724,N_2016);
nor U4675 (N_4675,N_350,N_2290);
and U4676 (N_4676,N_1228,N_2119);
xnor U4677 (N_4677,N_1311,N_1863);
nor U4678 (N_4678,N_1155,N_2204);
and U4679 (N_4679,N_839,N_1657);
nand U4680 (N_4680,N_463,N_157);
nand U4681 (N_4681,N_1848,N_1047);
nand U4682 (N_4682,N_1308,N_604);
nand U4683 (N_4683,N_256,N_134);
nand U4684 (N_4684,N_313,N_1256);
nand U4685 (N_4685,N_1662,N_1212);
nand U4686 (N_4686,N_2270,N_778);
nand U4687 (N_4687,N_1734,N_1723);
nor U4688 (N_4688,N_2309,N_1888);
nor U4689 (N_4689,N_1272,N_1425);
and U4690 (N_4690,N_953,N_2286);
nor U4691 (N_4691,N_1245,N_1136);
or U4692 (N_4692,N_1661,N_1339);
nor U4693 (N_4693,N_970,N_562);
and U4694 (N_4694,N_753,N_1953);
nand U4695 (N_4695,N_1986,N_333);
xor U4696 (N_4696,N_882,N_1036);
nor U4697 (N_4697,N_38,N_2267);
and U4698 (N_4698,N_537,N_677);
and U4699 (N_4699,N_1009,N_1013);
or U4700 (N_4700,N_633,N_2072);
xnor U4701 (N_4701,N_1994,N_1052);
nor U4702 (N_4702,N_2453,N_2393);
or U4703 (N_4703,N_1578,N_2339);
or U4704 (N_4704,N_963,N_285);
nand U4705 (N_4705,N_2256,N_1361);
and U4706 (N_4706,N_217,N_2412);
or U4707 (N_4707,N_931,N_1699);
nand U4708 (N_4708,N_855,N_275);
nor U4709 (N_4709,N_409,N_778);
nand U4710 (N_4710,N_773,N_2446);
and U4711 (N_4711,N_341,N_2177);
nand U4712 (N_4712,N_306,N_1525);
or U4713 (N_4713,N_304,N_2122);
and U4714 (N_4714,N_1637,N_2331);
or U4715 (N_4715,N_1087,N_1565);
and U4716 (N_4716,N_1772,N_1647);
nor U4717 (N_4717,N_1245,N_398);
or U4718 (N_4718,N_1412,N_1498);
nand U4719 (N_4719,N_768,N_2277);
nand U4720 (N_4720,N_1860,N_2432);
nor U4721 (N_4721,N_684,N_285);
nand U4722 (N_4722,N_1604,N_1724);
nor U4723 (N_4723,N_560,N_866);
and U4724 (N_4724,N_2448,N_1841);
nor U4725 (N_4725,N_206,N_2486);
and U4726 (N_4726,N_2329,N_265);
nand U4727 (N_4727,N_2024,N_338);
nor U4728 (N_4728,N_812,N_823);
xnor U4729 (N_4729,N_2042,N_1563);
nand U4730 (N_4730,N_94,N_27);
or U4731 (N_4731,N_1895,N_1077);
xnor U4732 (N_4732,N_319,N_251);
or U4733 (N_4733,N_2112,N_1232);
or U4734 (N_4734,N_327,N_2363);
nand U4735 (N_4735,N_2450,N_998);
and U4736 (N_4736,N_125,N_1588);
and U4737 (N_4737,N_1135,N_2290);
nand U4738 (N_4738,N_1591,N_963);
nor U4739 (N_4739,N_2281,N_531);
nor U4740 (N_4740,N_758,N_1124);
or U4741 (N_4741,N_60,N_460);
nor U4742 (N_4742,N_420,N_1);
nand U4743 (N_4743,N_921,N_1567);
nor U4744 (N_4744,N_141,N_731);
nand U4745 (N_4745,N_1839,N_2376);
nor U4746 (N_4746,N_1156,N_1417);
nor U4747 (N_4747,N_1402,N_925);
and U4748 (N_4748,N_2330,N_1096);
nand U4749 (N_4749,N_2396,N_4);
or U4750 (N_4750,N_1459,N_2174);
xor U4751 (N_4751,N_1184,N_1297);
nor U4752 (N_4752,N_1483,N_1236);
and U4753 (N_4753,N_1132,N_785);
and U4754 (N_4754,N_2470,N_1366);
nand U4755 (N_4755,N_885,N_479);
or U4756 (N_4756,N_1881,N_1049);
or U4757 (N_4757,N_2232,N_2048);
nor U4758 (N_4758,N_1185,N_1928);
and U4759 (N_4759,N_282,N_1796);
and U4760 (N_4760,N_1856,N_1848);
or U4761 (N_4761,N_1385,N_300);
nor U4762 (N_4762,N_1511,N_199);
and U4763 (N_4763,N_495,N_2237);
or U4764 (N_4764,N_1526,N_2106);
nand U4765 (N_4765,N_2163,N_1653);
nor U4766 (N_4766,N_146,N_570);
or U4767 (N_4767,N_1020,N_485);
or U4768 (N_4768,N_1288,N_1466);
nor U4769 (N_4769,N_78,N_221);
and U4770 (N_4770,N_743,N_80);
nor U4771 (N_4771,N_1708,N_15);
nand U4772 (N_4772,N_2023,N_752);
nand U4773 (N_4773,N_2040,N_2322);
and U4774 (N_4774,N_1613,N_1277);
or U4775 (N_4775,N_395,N_2248);
and U4776 (N_4776,N_1160,N_1929);
and U4777 (N_4777,N_2014,N_1881);
nand U4778 (N_4778,N_1512,N_1466);
nor U4779 (N_4779,N_391,N_1550);
or U4780 (N_4780,N_863,N_966);
and U4781 (N_4781,N_983,N_859);
nor U4782 (N_4782,N_645,N_2054);
and U4783 (N_4783,N_897,N_2380);
and U4784 (N_4784,N_1267,N_858);
and U4785 (N_4785,N_1143,N_246);
or U4786 (N_4786,N_2259,N_360);
nor U4787 (N_4787,N_2108,N_606);
nand U4788 (N_4788,N_342,N_1799);
nor U4789 (N_4789,N_2253,N_416);
and U4790 (N_4790,N_1042,N_1399);
or U4791 (N_4791,N_601,N_653);
nor U4792 (N_4792,N_2336,N_42);
nor U4793 (N_4793,N_2332,N_364);
nor U4794 (N_4794,N_587,N_45);
and U4795 (N_4795,N_1330,N_239);
nand U4796 (N_4796,N_2116,N_2055);
and U4797 (N_4797,N_880,N_1872);
or U4798 (N_4798,N_1433,N_1365);
and U4799 (N_4799,N_2313,N_876);
nand U4800 (N_4800,N_935,N_814);
nor U4801 (N_4801,N_2000,N_1602);
nand U4802 (N_4802,N_2048,N_872);
nor U4803 (N_4803,N_2298,N_1681);
or U4804 (N_4804,N_476,N_330);
nor U4805 (N_4805,N_350,N_2353);
nand U4806 (N_4806,N_855,N_926);
nand U4807 (N_4807,N_2077,N_1734);
and U4808 (N_4808,N_173,N_1301);
nand U4809 (N_4809,N_1981,N_335);
nor U4810 (N_4810,N_1892,N_1072);
nand U4811 (N_4811,N_1428,N_375);
nand U4812 (N_4812,N_1855,N_832);
and U4813 (N_4813,N_2299,N_1709);
nand U4814 (N_4814,N_2314,N_2456);
and U4815 (N_4815,N_343,N_853);
or U4816 (N_4816,N_1217,N_549);
and U4817 (N_4817,N_1612,N_1727);
nor U4818 (N_4818,N_125,N_2233);
or U4819 (N_4819,N_671,N_553);
nand U4820 (N_4820,N_689,N_792);
nand U4821 (N_4821,N_1785,N_1737);
nor U4822 (N_4822,N_2157,N_1790);
and U4823 (N_4823,N_570,N_1779);
nand U4824 (N_4824,N_1742,N_1703);
nor U4825 (N_4825,N_1563,N_2382);
or U4826 (N_4826,N_657,N_2143);
nor U4827 (N_4827,N_344,N_385);
or U4828 (N_4828,N_1892,N_1465);
nand U4829 (N_4829,N_335,N_1395);
nand U4830 (N_4830,N_301,N_308);
nand U4831 (N_4831,N_527,N_854);
and U4832 (N_4832,N_2270,N_2142);
nor U4833 (N_4833,N_968,N_367);
nand U4834 (N_4834,N_2306,N_1978);
nor U4835 (N_4835,N_1865,N_1385);
nor U4836 (N_4836,N_2476,N_2371);
nand U4837 (N_4837,N_1755,N_979);
and U4838 (N_4838,N_1468,N_1411);
nor U4839 (N_4839,N_671,N_469);
and U4840 (N_4840,N_953,N_2178);
or U4841 (N_4841,N_1194,N_2250);
or U4842 (N_4842,N_2321,N_59);
or U4843 (N_4843,N_2126,N_580);
and U4844 (N_4844,N_1320,N_630);
nor U4845 (N_4845,N_1852,N_2318);
or U4846 (N_4846,N_1443,N_1730);
and U4847 (N_4847,N_113,N_582);
and U4848 (N_4848,N_1548,N_2098);
and U4849 (N_4849,N_1571,N_262);
nand U4850 (N_4850,N_987,N_2402);
and U4851 (N_4851,N_2312,N_1970);
or U4852 (N_4852,N_2294,N_36);
nor U4853 (N_4853,N_845,N_2016);
or U4854 (N_4854,N_1741,N_1560);
or U4855 (N_4855,N_101,N_421);
nand U4856 (N_4856,N_554,N_2421);
or U4857 (N_4857,N_1100,N_1659);
or U4858 (N_4858,N_1224,N_1620);
nand U4859 (N_4859,N_1178,N_903);
nand U4860 (N_4860,N_129,N_1216);
and U4861 (N_4861,N_1449,N_166);
nand U4862 (N_4862,N_2493,N_1924);
nand U4863 (N_4863,N_1371,N_1110);
nor U4864 (N_4864,N_950,N_1074);
nand U4865 (N_4865,N_688,N_1937);
and U4866 (N_4866,N_1089,N_1416);
nor U4867 (N_4867,N_759,N_236);
xor U4868 (N_4868,N_2292,N_948);
nand U4869 (N_4869,N_143,N_1208);
nand U4870 (N_4870,N_1255,N_1469);
and U4871 (N_4871,N_2146,N_775);
and U4872 (N_4872,N_1271,N_1540);
and U4873 (N_4873,N_313,N_1909);
and U4874 (N_4874,N_598,N_771);
or U4875 (N_4875,N_2028,N_1587);
nand U4876 (N_4876,N_1542,N_1568);
and U4877 (N_4877,N_894,N_1361);
or U4878 (N_4878,N_1202,N_1891);
or U4879 (N_4879,N_640,N_97);
or U4880 (N_4880,N_597,N_852);
and U4881 (N_4881,N_685,N_1537);
nand U4882 (N_4882,N_294,N_203);
xnor U4883 (N_4883,N_1353,N_1756);
or U4884 (N_4884,N_931,N_2113);
nor U4885 (N_4885,N_1773,N_1313);
nor U4886 (N_4886,N_949,N_2308);
and U4887 (N_4887,N_153,N_1169);
nand U4888 (N_4888,N_1250,N_1522);
or U4889 (N_4889,N_1257,N_625);
and U4890 (N_4890,N_2154,N_839);
nor U4891 (N_4891,N_1266,N_1289);
and U4892 (N_4892,N_2131,N_864);
nor U4893 (N_4893,N_1580,N_222);
and U4894 (N_4894,N_655,N_575);
nand U4895 (N_4895,N_1258,N_2056);
and U4896 (N_4896,N_2201,N_1427);
nand U4897 (N_4897,N_2081,N_338);
nand U4898 (N_4898,N_218,N_958);
nor U4899 (N_4899,N_95,N_1768);
nand U4900 (N_4900,N_1182,N_152);
or U4901 (N_4901,N_2298,N_552);
or U4902 (N_4902,N_81,N_43);
nand U4903 (N_4903,N_755,N_748);
nor U4904 (N_4904,N_1986,N_2080);
nand U4905 (N_4905,N_1573,N_2077);
nor U4906 (N_4906,N_1274,N_352);
and U4907 (N_4907,N_2264,N_1625);
xor U4908 (N_4908,N_269,N_418);
or U4909 (N_4909,N_848,N_1580);
nand U4910 (N_4910,N_1591,N_1270);
nand U4911 (N_4911,N_1464,N_2218);
or U4912 (N_4912,N_2075,N_1097);
and U4913 (N_4913,N_1220,N_861);
nand U4914 (N_4914,N_607,N_1142);
or U4915 (N_4915,N_737,N_596);
and U4916 (N_4916,N_1012,N_2384);
nand U4917 (N_4917,N_2332,N_1534);
nor U4918 (N_4918,N_1444,N_1561);
nand U4919 (N_4919,N_1013,N_708);
and U4920 (N_4920,N_2112,N_2318);
or U4921 (N_4921,N_900,N_1458);
nand U4922 (N_4922,N_187,N_1808);
nor U4923 (N_4923,N_1335,N_1036);
xnor U4924 (N_4924,N_1186,N_708);
nor U4925 (N_4925,N_2184,N_816);
or U4926 (N_4926,N_123,N_245);
or U4927 (N_4927,N_1457,N_1298);
and U4928 (N_4928,N_536,N_354);
and U4929 (N_4929,N_309,N_1808);
or U4930 (N_4930,N_1739,N_2120);
and U4931 (N_4931,N_2406,N_1897);
and U4932 (N_4932,N_1848,N_1285);
and U4933 (N_4933,N_735,N_1803);
or U4934 (N_4934,N_928,N_1475);
nor U4935 (N_4935,N_1886,N_2259);
nand U4936 (N_4936,N_346,N_2241);
nor U4937 (N_4937,N_1514,N_484);
and U4938 (N_4938,N_1511,N_1239);
or U4939 (N_4939,N_1531,N_2141);
xnor U4940 (N_4940,N_1968,N_1984);
or U4941 (N_4941,N_962,N_1984);
and U4942 (N_4942,N_1778,N_896);
or U4943 (N_4943,N_1970,N_1300);
nor U4944 (N_4944,N_76,N_51);
nor U4945 (N_4945,N_2380,N_853);
nor U4946 (N_4946,N_887,N_696);
nand U4947 (N_4947,N_1478,N_273);
or U4948 (N_4948,N_1441,N_1472);
nor U4949 (N_4949,N_1586,N_2074);
nor U4950 (N_4950,N_2228,N_2402);
and U4951 (N_4951,N_620,N_1846);
or U4952 (N_4952,N_957,N_1373);
and U4953 (N_4953,N_1069,N_1245);
nand U4954 (N_4954,N_2010,N_1563);
or U4955 (N_4955,N_2300,N_258);
and U4956 (N_4956,N_1636,N_328);
and U4957 (N_4957,N_227,N_584);
or U4958 (N_4958,N_2190,N_2321);
nor U4959 (N_4959,N_555,N_1770);
and U4960 (N_4960,N_1477,N_2233);
nor U4961 (N_4961,N_691,N_791);
or U4962 (N_4962,N_1408,N_2470);
and U4963 (N_4963,N_287,N_2445);
and U4964 (N_4964,N_767,N_1714);
and U4965 (N_4965,N_498,N_753);
and U4966 (N_4966,N_679,N_1206);
nand U4967 (N_4967,N_41,N_2314);
or U4968 (N_4968,N_2055,N_2269);
nor U4969 (N_4969,N_2396,N_1240);
and U4970 (N_4970,N_1913,N_2025);
nor U4971 (N_4971,N_1314,N_1800);
or U4972 (N_4972,N_154,N_1729);
and U4973 (N_4973,N_969,N_2223);
or U4974 (N_4974,N_2115,N_405);
and U4975 (N_4975,N_1690,N_1612);
or U4976 (N_4976,N_2177,N_1443);
and U4977 (N_4977,N_2361,N_2160);
nor U4978 (N_4978,N_2208,N_2313);
or U4979 (N_4979,N_2093,N_451);
or U4980 (N_4980,N_18,N_2237);
nor U4981 (N_4981,N_1117,N_2452);
nor U4982 (N_4982,N_2467,N_1354);
nand U4983 (N_4983,N_1469,N_2359);
and U4984 (N_4984,N_1471,N_1965);
or U4985 (N_4985,N_0,N_668);
nor U4986 (N_4986,N_1805,N_165);
and U4987 (N_4987,N_635,N_245);
nand U4988 (N_4988,N_247,N_1555);
and U4989 (N_4989,N_1174,N_2173);
nor U4990 (N_4990,N_1626,N_1863);
nand U4991 (N_4991,N_2051,N_493);
nor U4992 (N_4992,N_726,N_209);
and U4993 (N_4993,N_866,N_2008);
nor U4994 (N_4994,N_1771,N_2268);
nand U4995 (N_4995,N_1097,N_2380);
or U4996 (N_4996,N_2427,N_1282);
nand U4997 (N_4997,N_2335,N_2107);
xnor U4998 (N_4998,N_980,N_102);
nand U4999 (N_4999,N_2183,N_391);
and UO_0 (O_0,N_2675,N_2804);
nor UO_1 (O_1,N_3494,N_2629);
or UO_2 (O_2,N_4623,N_4654);
nor UO_3 (O_3,N_2899,N_4980);
nand UO_4 (O_4,N_4577,N_4279);
nor UO_5 (O_5,N_3599,N_4106);
nor UO_6 (O_6,N_4524,N_2586);
nand UO_7 (O_7,N_3179,N_2896);
and UO_8 (O_8,N_3680,N_3534);
or UO_9 (O_9,N_4790,N_4302);
or UO_10 (O_10,N_4645,N_3014);
or UO_11 (O_11,N_4268,N_2703);
or UO_12 (O_12,N_2822,N_3093);
nor UO_13 (O_13,N_4311,N_4935);
nor UO_14 (O_14,N_3381,N_4299);
or UO_15 (O_15,N_2817,N_2736);
nand UO_16 (O_16,N_4241,N_4875);
or UO_17 (O_17,N_3242,N_2893);
nor UO_18 (O_18,N_4591,N_4284);
and UO_19 (O_19,N_4447,N_4999);
nor UO_20 (O_20,N_4818,N_3730);
nor UO_21 (O_21,N_2989,N_4783);
or UO_22 (O_22,N_3961,N_3859);
nor UO_23 (O_23,N_4641,N_2514);
and UO_24 (O_24,N_4061,N_3023);
and UO_25 (O_25,N_3272,N_4620);
xnor UO_26 (O_26,N_2545,N_4348);
nor UO_27 (O_27,N_4810,N_3792);
nor UO_28 (O_28,N_2710,N_3729);
nand UO_29 (O_29,N_3224,N_4333);
nor UO_30 (O_30,N_3246,N_2818);
nor UO_31 (O_31,N_3276,N_3503);
nor UO_32 (O_32,N_3172,N_3674);
nor UO_33 (O_33,N_2800,N_4438);
nand UO_34 (O_34,N_4157,N_2768);
nand UO_35 (O_35,N_4408,N_4187);
nor UO_36 (O_36,N_3028,N_3871);
or UO_37 (O_37,N_3623,N_3775);
nor UO_38 (O_38,N_4557,N_3453);
nor UO_39 (O_39,N_2531,N_4288);
or UO_40 (O_40,N_2953,N_2936);
nor UO_41 (O_41,N_2977,N_2633);
or UO_42 (O_42,N_4622,N_3132);
nand UO_43 (O_43,N_4269,N_3541);
and UO_44 (O_44,N_3336,N_4668);
or UO_45 (O_45,N_3116,N_4858);
and UO_46 (O_46,N_4617,N_2644);
and UO_47 (O_47,N_3331,N_2704);
nor UO_48 (O_48,N_4426,N_3300);
xnor UO_49 (O_49,N_2552,N_3423);
and UO_50 (O_50,N_2909,N_2544);
and UO_51 (O_51,N_3736,N_4970);
or UO_52 (O_52,N_2820,N_3883);
nor UO_53 (O_53,N_2961,N_4256);
and UO_54 (O_54,N_4904,N_3654);
nor UO_55 (O_55,N_3185,N_3867);
nand UO_56 (O_56,N_3977,N_3012);
or UO_57 (O_57,N_4990,N_4488);
and UO_58 (O_58,N_3872,N_3558);
or UO_59 (O_59,N_3760,N_2527);
and UO_60 (O_60,N_3108,N_3629);
or UO_61 (O_61,N_4081,N_3406);
nor UO_62 (O_62,N_4227,N_3878);
nand UO_63 (O_63,N_2747,N_4240);
nand UO_64 (O_64,N_3789,N_4983);
and UO_65 (O_65,N_3841,N_3669);
nand UO_66 (O_66,N_3784,N_4327);
or UO_67 (O_67,N_3635,N_2942);
or UO_68 (O_68,N_4979,N_4646);
and UO_69 (O_69,N_4530,N_3781);
nand UO_70 (O_70,N_4829,N_2507);
nor UO_71 (O_71,N_4254,N_3299);
or UO_72 (O_72,N_3155,N_4811);
or UO_73 (O_73,N_3460,N_3316);
or UO_74 (O_74,N_4020,N_3811);
nor UO_75 (O_75,N_3055,N_3437);
nor UO_76 (O_76,N_3787,N_4863);
nor UO_77 (O_77,N_2607,N_4204);
or UO_78 (O_78,N_3442,N_4985);
and UO_79 (O_79,N_3112,N_3470);
and UO_80 (O_80,N_4974,N_4153);
nor UO_81 (O_81,N_2528,N_2661);
nor UO_82 (O_82,N_2976,N_2648);
and UO_83 (O_83,N_3214,N_4515);
nor UO_84 (O_84,N_4422,N_3933);
nand UO_85 (O_85,N_2513,N_2696);
and UO_86 (O_86,N_2515,N_4995);
or UO_87 (O_87,N_4819,N_3474);
or UO_88 (O_88,N_3615,N_2958);
or UO_89 (O_89,N_4582,N_4843);
and UO_90 (O_90,N_4748,N_3742);
nor UO_91 (O_91,N_4162,N_3270);
and UO_92 (O_92,N_4111,N_3888);
or UO_93 (O_93,N_3123,N_4826);
nor UO_94 (O_94,N_4677,N_4893);
or UO_95 (O_95,N_3355,N_4738);
nand UO_96 (O_96,N_4362,N_3614);
and UO_97 (O_97,N_4638,N_2780);
nand UO_98 (O_98,N_4316,N_4584);
nand UO_99 (O_99,N_4016,N_4948);
or UO_100 (O_100,N_4036,N_2740);
nand UO_101 (O_101,N_4124,N_4412);
and UO_102 (O_102,N_4267,N_2755);
and UO_103 (O_103,N_2658,N_4815);
and UO_104 (O_104,N_2911,N_4652);
and UO_105 (O_105,N_3075,N_4116);
or UO_106 (O_106,N_3994,N_3861);
nor UO_107 (O_107,N_3069,N_2752);
and UO_108 (O_108,N_2579,N_2746);
nand UO_109 (O_109,N_4222,N_3676);
nor UO_110 (O_110,N_4618,N_4570);
nor UO_111 (O_111,N_3717,N_2775);
or UO_112 (O_112,N_4266,N_3547);
and UO_113 (O_113,N_3548,N_2944);
and UO_114 (O_114,N_3800,N_3557);
and UO_115 (O_115,N_4171,N_3053);
nand UO_116 (O_116,N_4834,N_3661);
and UO_117 (O_117,N_4726,N_2522);
and UO_118 (O_118,N_4814,N_3328);
or UO_119 (O_119,N_2761,N_4499);
nand UO_120 (O_120,N_3147,N_2779);
xnor UO_121 (O_121,N_4375,N_3191);
nand UO_122 (O_122,N_4216,N_3448);
and UO_123 (O_123,N_4528,N_2753);
nand UO_124 (O_124,N_4547,N_4516);
or UO_125 (O_125,N_4868,N_4031);
or UO_126 (O_126,N_3087,N_3283);
or UO_127 (O_127,N_4601,N_2729);
and UO_128 (O_128,N_2835,N_4723);
or UO_129 (O_129,N_4573,N_2565);
nand UO_130 (O_130,N_4713,N_2951);
xor UO_131 (O_131,N_3960,N_4318);
nand UO_132 (O_132,N_2762,N_3898);
or UO_133 (O_133,N_2730,N_2542);
nor UO_134 (O_134,N_3485,N_4202);
or UO_135 (O_135,N_4381,N_4593);
or UO_136 (O_136,N_4386,N_3816);
nand UO_137 (O_137,N_4356,N_3291);
and UO_138 (O_138,N_3692,N_4614);
or UO_139 (O_139,N_3201,N_2720);
and UO_140 (O_140,N_4631,N_3148);
or UO_141 (O_141,N_3011,N_4708);
and UO_142 (O_142,N_3335,N_2885);
nor UO_143 (O_143,N_4002,N_4700);
nand UO_144 (O_144,N_3181,N_3520);
or UO_145 (O_145,N_3866,N_2606);
nand UO_146 (O_146,N_4827,N_4351);
and UO_147 (O_147,N_3576,N_4443);
nand UO_148 (O_148,N_4508,N_4369);
and UO_149 (O_149,N_4378,N_4535);
and UO_150 (O_150,N_4857,N_3512);
nor UO_151 (O_151,N_2937,N_4704);
or UO_152 (O_152,N_2934,N_4048);
nand UO_153 (O_153,N_3255,N_3468);
nand UO_154 (O_154,N_2939,N_3537);
nand UO_155 (O_155,N_3279,N_2693);
nor UO_156 (O_156,N_4213,N_2639);
and UO_157 (O_157,N_3110,N_3167);
xor UO_158 (O_158,N_3006,N_3881);
or UO_159 (O_159,N_4587,N_3955);
nand UO_160 (O_160,N_3435,N_4096);
nand UO_161 (O_161,N_3098,N_4077);
nand UO_162 (O_162,N_4491,N_3719);
nor UO_163 (O_163,N_4714,N_2569);
nor UO_164 (O_164,N_4835,N_4095);
and UO_165 (O_165,N_3851,N_4912);
nor UO_166 (O_166,N_3289,N_3815);
and UO_167 (O_167,N_4179,N_3128);
and UO_168 (O_168,N_4024,N_4576);
xor UO_169 (O_169,N_2880,N_2935);
nand UO_170 (O_170,N_3382,N_3579);
or UO_171 (O_171,N_4388,N_4554);
nand UO_172 (O_172,N_3310,N_2931);
nand UO_173 (O_173,N_4621,N_4754);
or UO_174 (O_174,N_4192,N_4876);
and UO_175 (O_175,N_3997,N_4324);
and UO_176 (O_176,N_2652,N_3543);
nor UO_177 (O_177,N_4035,N_3732);
nor UO_178 (O_178,N_4849,N_2921);
and UO_179 (O_179,N_3184,N_4161);
nor UO_180 (O_180,N_4578,N_4329);
and UO_181 (O_181,N_2655,N_4907);
or UO_182 (O_182,N_3486,N_3829);
and UO_183 (O_183,N_4032,N_4962);
or UO_184 (O_184,N_3493,N_3797);
and UO_185 (O_185,N_4926,N_3428);
xor UO_186 (O_186,N_4828,N_4552);
nor UO_187 (O_187,N_3945,N_3793);
and UO_188 (O_188,N_4751,N_4233);
and UO_189 (O_189,N_3915,N_2521);
nand UO_190 (O_190,N_4777,N_3713);
or UO_191 (O_191,N_2722,N_3810);
and UO_192 (O_192,N_3753,N_3575);
and UO_193 (O_193,N_3221,N_4851);
nand UO_194 (O_194,N_4113,N_3206);
or UO_195 (O_195,N_3858,N_3294);
nor UO_196 (O_196,N_2887,N_3666);
nand UO_197 (O_197,N_4778,N_4634);
nand UO_198 (O_198,N_2573,N_4784);
nor UO_199 (O_199,N_4379,N_3973);
or UO_200 (O_200,N_4219,N_4878);
nand UO_201 (O_201,N_3904,N_2611);
and UO_202 (O_202,N_2813,N_4996);
nand UO_203 (O_203,N_4629,N_3507);
and UO_204 (O_204,N_4997,N_3786);
and UO_205 (O_205,N_2824,N_4448);
or UO_206 (O_206,N_4138,N_3903);
nand UO_207 (O_207,N_2653,N_4928);
or UO_208 (O_208,N_3646,N_4414);
or UO_209 (O_209,N_4038,N_4459);
nor UO_210 (O_210,N_4984,N_2727);
and UO_211 (O_211,N_4698,N_3342);
nor UO_212 (O_212,N_4988,N_4797);
or UO_213 (O_213,N_4596,N_4569);
nand UO_214 (O_214,N_3293,N_4107);
nor UO_215 (O_215,N_2758,N_4142);
and UO_216 (O_216,N_3038,N_3051);
and UO_217 (O_217,N_3954,N_4026);
or UO_218 (O_218,N_4001,N_2580);
or UO_219 (O_219,N_2827,N_3444);
nand UO_220 (O_220,N_3445,N_2938);
and UO_221 (O_221,N_3348,N_3838);
nor UO_222 (O_222,N_4133,N_3086);
nor UO_223 (O_223,N_3318,N_2726);
nand UO_224 (O_224,N_3387,N_4939);
or UO_225 (O_225,N_4529,N_3026);
nor UO_226 (O_226,N_2516,N_2678);
or UO_227 (O_227,N_2778,N_4357);
and UO_228 (O_228,N_3064,N_4163);
and UO_229 (O_229,N_4368,N_4390);
xnor UO_230 (O_230,N_3080,N_3127);
nor UO_231 (O_231,N_3198,N_3603);
xor UO_232 (O_232,N_2748,N_2867);
and UO_233 (O_233,N_3450,N_4028);
or UO_234 (O_234,N_2612,N_3413);
and UO_235 (O_235,N_2789,N_4595);
or UO_236 (O_236,N_2815,N_3684);
nand UO_237 (O_237,N_3021,N_2664);
and UO_238 (O_238,N_4109,N_4239);
or UO_239 (O_239,N_3993,N_3078);
and UO_240 (O_240,N_4429,N_4973);
and UO_241 (O_241,N_4667,N_3927);
or UO_242 (O_242,N_3802,N_2994);
nand UO_243 (O_243,N_4006,N_4419);
nand UO_244 (O_244,N_2949,N_3912);
or UO_245 (O_245,N_4504,N_3999);
nand UO_246 (O_246,N_3017,N_2734);
nand UO_247 (O_247,N_4866,N_3264);
and UO_248 (O_248,N_4966,N_4913);
nand UO_249 (O_249,N_4675,N_2799);
nor UO_250 (O_250,N_2805,N_3583);
and UO_251 (O_251,N_4662,N_4789);
nand UO_252 (O_252,N_4029,N_4588);
or UO_253 (O_253,N_2883,N_3842);
nand UO_254 (O_254,N_3054,N_3481);
or UO_255 (O_255,N_4347,N_4718);
and UO_256 (O_256,N_4476,N_3979);
nor UO_257 (O_257,N_2784,N_4188);
and UO_258 (O_258,N_3770,N_4717);
nor UO_259 (O_259,N_4538,N_3588);
nand UO_260 (O_260,N_3584,N_3948);
nand UO_261 (O_261,N_4687,N_4169);
nor UO_262 (O_262,N_4669,N_4313);
or UO_263 (O_263,N_4630,N_2791);
nor UO_264 (O_264,N_4119,N_3307);
nor UO_265 (O_265,N_3321,N_4201);
and UO_266 (O_266,N_4613,N_3002);
and UO_267 (O_267,N_3314,N_3183);
nand UO_268 (O_268,N_2974,N_4534);
nor UO_269 (O_269,N_4451,N_4817);
and UO_270 (O_270,N_4394,N_3721);
and UO_271 (O_271,N_3504,N_4200);
or UO_272 (O_272,N_2584,N_2701);
nor UO_273 (O_273,N_2952,N_4155);
or UO_274 (O_274,N_4590,N_3984);
xnor UO_275 (O_275,N_3862,N_2616);
and UO_276 (O_276,N_4184,N_3562);
nor UO_277 (O_277,N_3174,N_4089);
or UO_278 (O_278,N_4151,N_4177);
or UO_279 (O_279,N_2591,N_3107);
nor UO_280 (O_280,N_4384,N_3708);
nand UO_281 (O_281,N_3855,N_2631);
nor UO_282 (O_282,N_2964,N_2860);
nor UO_283 (O_283,N_4409,N_4862);
and UO_284 (O_284,N_3394,N_4431);
or UO_285 (O_285,N_4600,N_4741);
and UO_286 (O_286,N_4067,N_4354);
and UO_287 (O_287,N_4705,N_2763);
or UO_288 (O_288,N_3620,N_3509);
and UO_289 (O_289,N_2533,N_3315);
or UO_290 (O_290,N_3642,N_2666);
nand UO_291 (O_291,N_3649,N_2691);
or UO_292 (O_292,N_3613,N_4442);
or UO_293 (O_293,N_4599,N_3372);
nand UO_294 (O_294,N_2863,N_4487);
nor UO_295 (O_295,N_4088,N_4249);
nand UO_296 (O_296,N_2587,N_3390);
or UO_297 (O_297,N_4173,N_3517);
nor UO_298 (O_298,N_3625,N_3922);
or UO_299 (O_299,N_4477,N_3375);
or UO_300 (O_300,N_4047,N_4317);
nor UO_301 (O_301,N_2694,N_4309);
nor UO_302 (O_302,N_3253,N_2877);
or UO_303 (O_303,N_4110,N_4507);
nor UO_304 (O_304,N_3130,N_2560);
nor UO_305 (O_305,N_4364,N_3893);
nand UO_306 (O_306,N_3636,N_2922);
nand UO_307 (O_307,N_3089,N_4796);
nand UO_308 (O_308,N_4845,N_4609);
xnor UO_309 (O_309,N_3259,N_2642);
and UO_310 (O_310,N_3595,N_3209);
nand UO_311 (O_311,N_2684,N_3502);
nand UO_312 (O_312,N_4146,N_2770);
and UO_313 (O_313,N_3273,N_4886);
nor UO_314 (O_314,N_2558,N_3681);
or UO_315 (O_315,N_3928,N_4140);
nand UO_316 (O_316,N_4961,N_3677);
xnor UO_317 (O_317,N_3398,N_3426);
nor UO_318 (O_318,N_2793,N_2744);
nand UO_319 (O_319,N_3832,N_3794);
and UO_320 (O_320,N_2795,N_3325);
or UO_321 (O_321,N_3956,N_2844);
and UO_322 (O_322,N_3852,N_3408);
and UO_323 (O_323,N_3709,N_2509);
and UO_324 (O_324,N_3532,N_3738);
nand UO_325 (O_325,N_2914,N_3570);
nand UO_326 (O_326,N_2614,N_3963);
or UO_327 (O_327,N_4752,N_4425);
nand UO_328 (O_328,N_2900,N_4602);
or UO_329 (O_329,N_4370,N_4383);
nand UO_330 (O_330,N_4658,N_3974);
or UO_331 (O_331,N_3156,N_2991);
nand UO_332 (O_332,N_4214,N_3530);
nor UO_333 (O_333,N_3284,N_3773);
nand UO_334 (O_334,N_3941,N_4247);
nand UO_335 (O_335,N_4837,N_3846);
or UO_336 (O_336,N_2617,N_3889);
nor UO_337 (O_337,N_3250,N_4340);
nor UO_338 (O_338,N_3429,N_2575);
and UO_339 (O_339,N_4551,N_2923);
nand UO_340 (O_340,N_4968,N_2853);
and UO_341 (O_341,N_3431,N_4971);
and UO_342 (O_342,N_4485,N_3142);
or UO_343 (O_343,N_4315,N_3686);
nor UO_344 (O_344,N_4888,N_4393);
and UO_345 (O_345,N_3601,N_3281);
nand UO_346 (O_346,N_4044,N_3785);
and UO_347 (O_347,N_2972,N_4804);
or UO_348 (O_348,N_3016,N_4149);
nor UO_349 (O_349,N_2596,N_4991);
or UO_350 (O_350,N_3092,N_4355);
and UO_351 (O_351,N_4690,N_4732);
and UO_352 (O_352,N_3990,N_4385);
and UO_353 (O_353,N_2610,N_2927);
or UO_354 (O_354,N_3177,N_4695);
xor UO_355 (O_355,N_4478,N_3505);
or UO_356 (O_356,N_3380,N_4349);
nand UO_357 (O_357,N_3670,N_4532);
or UO_358 (O_358,N_3047,N_3671);
and UO_359 (O_359,N_3393,N_4005);
nand UO_360 (O_360,N_4852,N_3714);
and UO_361 (O_361,N_4734,N_2687);
xnor UO_362 (O_362,N_4071,N_4321);
or UO_363 (O_363,N_3025,N_2881);
and UO_364 (O_364,N_2978,N_2852);
nor UO_365 (O_365,N_4286,N_3070);
nand UO_366 (O_366,N_2537,N_4884);
nor UO_367 (O_367,N_4208,N_4281);
nand UO_368 (O_368,N_3814,N_2821);
or UO_369 (O_369,N_2654,N_3594);
or UO_370 (O_370,N_3225,N_4685);
and UO_371 (O_371,N_3518,N_4359);
or UO_372 (O_372,N_4402,N_3019);
or UO_373 (O_373,N_4079,N_4159);
or UO_374 (O_374,N_2618,N_2969);
nand UO_375 (O_375,N_4471,N_3344);
nand UO_376 (O_376,N_4461,N_4870);
and UO_377 (O_377,N_4441,N_3418);
nand UO_378 (O_378,N_4715,N_2719);
nor UO_379 (O_379,N_3129,N_3488);
or UO_380 (O_380,N_3672,N_4245);
nand UO_381 (O_381,N_3880,N_4903);
nand UO_382 (O_382,N_3868,N_3357);
or UO_383 (O_383,N_4549,N_3897);
or UO_384 (O_384,N_3578,N_3275);
or UO_385 (O_385,N_4023,N_2757);
nand UO_386 (O_386,N_3650,N_4839);
or UO_387 (O_387,N_2731,N_4041);
nor UO_388 (O_388,N_2806,N_3907);
and UO_389 (O_389,N_2624,N_3391);
or UO_390 (O_390,N_2585,N_3947);
and UO_391 (O_391,N_4086,N_3812);
nand UO_392 (O_392,N_4434,N_4794);
and UO_393 (O_393,N_3533,N_4018);
and UO_394 (O_394,N_2568,N_3683);
nand UO_395 (O_395,N_3483,N_2862);
or UO_396 (O_396,N_3571,N_3740);
nor UO_397 (O_397,N_4374,N_4290);
and UO_398 (O_398,N_4051,N_4182);
or UO_399 (O_399,N_3633,N_4460);
nand UO_400 (O_400,N_4372,N_3001);
nand UO_401 (O_401,N_3141,N_2843);
and UO_402 (O_402,N_3820,N_3340);
xor UO_403 (O_403,N_4655,N_4865);
nand UO_404 (O_404,N_4099,N_3296);
and UO_405 (O_405,N_3632,N_4944);
xor UO_406 (O_406,N_3559,N_3235);
or UO_407 (O_407,N_2670,N_4468);
nand UO_408 (O_408,N_3782,N_2572);
nor UO_409 (O_409,N_2798,N_4806);
nand UO_410 (O_410,N_3010,N_2620);
or UO_411 (O_411,N_2711,N_3737);
nand UO_412 (O_412,N_4101,N_2878);
and UO_413 (O_413,N_4352,N_3440);
or UO_414 (O_414,N_3833,N_3663);
or UO_415 (O_415,N_3101,N_4567);
xnor UO_416 (O_416,N_2858,N_4392);
and UO_417 (O_417,N_4847,N_4880);
nor UO_418 (O_418,N_4575,N_4689);
or UO_419 (O_419,N_2754,N_3567);
or UO_420 (O_420,N_3555,N_4568);
and UO_421 (O_421,N_4562,N_2647);
xor UO_422 (O_422,N_2674,N_2589);
nor UO_423 (O_423,N_2870,N_4749);
or UO_424 (O_424,N_2538,N_4952);
nand UO_425 (O_425,N_4730,N_2871);
nor UO_426 (O_426,N_2739,N_3490);
nand UO_427 (O_427,N_3170,N_2534);
and UO_428 (O_428,N_4503,N_3228);
nor UO_429 (O_429,N_4975,N_4505);
nor UO_430 (O_430,N_4322,N_2619);
and UO_431 (O_431,N_3723,N_4501);
nor UO_432 (O_432,N_4663,N_3951);
nor UO_433 (O_433,N_3371,N_3402);
and UO_434 (O_434,N_3964,N_2523);
and UO_435 (O_435,N_2832,N_4167);
nand UO_436 (O_436,N_4585,N_3249);
xor UO_437 (O_437,N_4774,N_2659);
or UO_438 (O_438,N_4820,N_3403);
or UO_439 (O_439,N_4122,N_3911);
or UO_440 (O_440,N_3545,N_3205);
nor UO_441 (O_441,N_2645,N_2872);
or UO_442 (O_442,N_3159,N_4398);
nand UO_443 (O_443,N_4871,N_3404);
nor UO_444 (O_444,N_3525,N_3226);
or UO_445 (O_445,N_4525,N_4693);
or UO_446 (O_446,N_3085,N_4558);
nor UO_447 (O_447,N_4571,N_2906);
or UO_448 (O_448,N_3966,N_2567);
nand UO_449 (O_449,N_4637,N_4951);
nand UO_450 (O_450,N_4498,N_2916);
nand UO_451 (O_451,N_4625,N_3126);
nand UO_452 (O_452,N_4400,N_2713);
xor UO_453 (O_453,N_3550,N_4882);
xor UO_454 (O_454,N_2946,N_4453);
and UO_455 (O_455,N_4212,N_3122);
nand UO_456 (O_456,N_3901,N_2803);
nor UO_457 (O_457,N_2504,N_3739);
nand UO_458 (O_458,N_4276,N_2995);
nor UO_459 (O_459,N_4413,N_2708);
and UO_460 (O_460,N_3361,N_3712);
nand UO_461 (O_461,N_3914,N_3056);
and UO_462 (O_462,N_4428,N_3574);
nor UO_463 (O_463,N_3349,N_3194);
or UO_464 (O_464,N_3462,N_2971);
or UO_465 (O_465,N_4154,N_3876);
and UO_466 (O_466,N_2982,N_4873);
xnor UO_467 (O_467,N_2510,N_3608);
or UO_468 (O_468,N_4215,N_4616);
nand UO_469 (O_469,N_4671,N_4519);
nor UO_470 (O_470,N_4175,N_4492);
or UO_471 (O_471,N_4297,N_4440);
nor UO_472 (O_472,N_3117,N_4543);
and UO_473 (O_473,N_4805,N_2983);
nor UO_474 (O_474,N_3424,N_2787);
and UO_475 (O_475,N_3327,N_3285);
and UO_476 (O_476,N_3887,N_3083);
nand UO_477 (O_477,N_2628,N_3779);
and UO_478 (O_478,N_4833,N_4982);
nand UO_479 (O_479,N_4211,N_4205);
xnor UO_480 (O_480,N_4792,N_3188);
nand UO_481 (O_481,N_3059,N_3434);
or UO_482 (O_482,N_3808,N_4517);
nand UO_483 (O_483,N_4228,N_4799);
and UO_484 (O_484,N_3703,N_3251);
or UO_485 (O_485,N_3624,N_3892);
nand UO_486 (O_486,N_2621,N_2535);
or UO_487 (O_487,N_3885,N_3510);
or UO_488 (O_488,N_4040,N_2875);
or UO_489 (O_489,N_3640,N_2773);
or UO_490 (O_490,N_3190,N_4758);
nor UO_491 (O_491,N_2699,N_3171);
or UO_492 (O_492,N_3587,N_3891);
nand UO_493 (O_493,N_3109,N_2505);
or UO_494 (O_494,N_3140,N_3419);
and UO_495 (O_495,N_4755,N_4782);
nand UO_496 (O_496,N_2500,N_3005);
and UO_497 (O_497,N_4773,N_3496);
and UO_498 (O_498,N_2590,N_3873);
nand UO_499 (O_499,N_4259,N_4277);
nor UO_500 (O_500,N_3265,N_3392);
or UO_501 (O_501,N_2767,N_3439);
and UO_502 (O_502,N_4344,N_4465);
nor UO_503 (O_503,N_4307,N_3241);
or UO_504 (O_504,N_4553,N_3678);
nor UO_505 (O_505,N_3041,N_3965);
nor UO_506 (O_506,N_4221,N_4462);
xnor UO_507 (O_507,N_2841,N_4021);
nand UO_508 (O_508,N_3801,N_2520);
nor UO_509 (O_509,N_3385,N_4178);
nand UO_510 (O_510,N_4709,N_3685);
and UO_511 (O_511,N_4564,N_3164);
nor UO_512 (O_512,N_3938,N_4278);
nor UO_513 (O_513,N_3060,N_2656);
nand UO_514 (O_514,N_2968,N_3527);
nand UO_515 (O_515,N_4090,N_4064);
xor UO_516 (O_516,N_4436,N_3529);
nor UO_517 (O_517,N_3232,N_4628);
nor UO_518 (O_518,N_3682,N_3227);
nand UO_519 (O_519,N_4083,N_3352);
and UO_520 (O_520,N_3498,N_3524);
nor UO_521 (O_521,N_2595,N_3030);
and UO_522 (O_522,N_4457,N_3256);
nor UO_523 (O_523,N_3478,N_2897);
and UO_524 (O_524,N_3359,N_3652);
xor UO_525 (O_525,N_3077,N_3696);
nor UO_526 (O_526,N_3222,N_3675);
nand UO_527 (O_527,N_4583,N_2930);
nand UO_528 (O_528,N_3007,N_4114);
nand UO_529 (O_529,N_4721,N_4444);
xnor UO_530 (O_530,N_3236,N_3304);
and UO_531 (O_531,N_3909,N_4929);
and UO_532 (O_532,N_3634,N_2912);
nor UO_533 (O_533,N_2772,N_3853);
or UO_534 (O_534,N_3818,N_4526);
nor UO_535 (O_535,N_3621,N_2884);
or UO_536 (O_536,N_4831,N_4353);
and UO_537 (O_537,N_4404,N_2626);
or UO_538 (O_538,N_3495,N_4605);
and UO_539 (O_539,N_3750,N_3161);
nor UO_540 (O_540,N_4509,N_2562);
nand UO_541 (O_541,N_3096,N_4210);
or UO_542 (O_542,N_2517,N_2539);
and UO_543 (O_543,N_3274,N_3351);
and UO_544 (O_544,N_3568,N_3978);
and UO_545 (O_545,N_4013,N_2792);
or UO_546 (O_546,N_3491,N_4686);
nand UO_547 (O_547,N_4510,N_4604);
nor UO_548 (O_548,N_2686,N_3377);
or UO_549 (O_549,N_4294,N_3913);
nand UO_550 (O_550,N_2864,N_2530);
and UO_551 (O_551,N_3311,N_4164);
nand UO_552 (O_552,N_3415,N_4946);
nand UO_553 (O_553,N_3932,N_3263);
or UO_554 (O_554,N_4022,N_2603);
nand UO_555 (O_555,N_4435,N_2511);
or UO_556 (O_556,N_3317,N_4174);
nor UO_557 (O_557,N_3606,N_3193);
or UO_558 (O_558,N_3734,N_4993);
and UO_559 (O_559,N_4225,N_4054);
nor UO_560 (O_560,N_3076,N_3539);
and UO_561 (O_561,N_3239,N_3728);
nor UO_562 (O_562,N_3166,N_4475);
nand UO_563 (O_563,N_2786,N_3653);
and UO_564 (O_564,N_4074,N_3989);
and UO_565 (O_565,N_4326,N_3383);
or UO_566 (O_566,N_3119,N_3687);
nand UO_567 (O_567,N_2920,N_4731);
and UO_568 (O_568,N_4072,N_4977);
nand UO_569 (O_569,N_4437,N_3451);
or UO_570 (O_570,N_4965,N_4181);
nand UO_571 (O_571,N_2543,N_4217);
xnor UO_572 (O_572,N_4237,N_3573);
and UO_573 (O_573,N_4135,N_4198);
or UO_574 (O_574,N_2928,N_4544);
nor UO_575 (O_575,N_3996,N_3609);
and UO_576 (O_576,N_2945,N_4156);
or UO_577 (O_577,N_3202,N_4759);
nand UO_578 (O_578,N_3985,N_4786);
or UO_579 (O_579,N_4416,N_2765);
nor UO_580 (O_580,N_2632,N_2839);
or UO_581 (O_581,N_3282,N_3366);
and UO_582 (O_582,N_3037,N_4118);
or UO_583 (O_583,N_4301,N_4433);
nand UO_584 (O_584,N_3551,N_4720);
nand UO_585 (O_585,N_2895,N_3034);
nor UO_586 (O_586,N_3765,N_4779);
nor UO_587 (O_587,N_2980,N_4489);
or UO_588 (O_588,N_2796,N_4410);
or UO_589 (O_589,N_2698,N_3690);
and UO_590 (O_590,N_3582,N_3103);
or UO_591 (O_591,N_4938,N_4250);
nor UO_592 (O_592,N_3519,N_3627);
or UO_593 (O_593,N_4458,N_4445);
nor UO_594 (O_594,N_3000,N_3144);
nor UO_595 (O_595,N_4750,N_3879);
and UO_596 (O_596,N_3091,N_2855);
nand UO_597 (O_597,N_2738,N_2764);
or UO_598 (O_598,N_3735,N_3707);
nand UO_599 (O_599,N_3003,N_3757);
or UO_600 (O_600,N_4147,N_2907);
nor UO_601 (O_601,N_3698,N_3039);
xnor UO_602 (O_602,N_3029,N_3899);
and UO_603 (O_603,N_3452,N_3776);
and UO_604 (O_604,N_3528,N_3937);
or UO_605 (O_605,N_3455,N_4896);
or UO_606 (O_606,N_4521,N_3339);
or UO_607 (O_607,N_3163,N_4531);
nor UO_608 (O_608,N_2913,N_4242);
xnor UO_609 (O_609,N_4639,N_4030);
or UO_610 (O_610,N_3602,N_4694);
and UO_611 (O_611,N_4045,N_4399);
and UO_612 (O_612,N_4987,N_3208);
nor UO_613 (O_613,N_4895,N_3324);
nand UO_614 (O_614,N_3755,N_3248);
nor UO_615 (O_615,N_3596,N_3743);
nand UO_616 (O_616,N_4479,N_2814);
and UO_617 (O_617,N_4097,N_3297);
and UO_618 (O_618,N_3902,N_3724);
nor UO_619 (O_619,N_2886,N_3959);
or UO_620 (O_620,N_3295,N_3186);
nand UO_621 (O_621,N_3196,N_3700);
and UO_622 (O_622,N_4559,N_3302);
nand UO_623 (O_623,N_4480,N_3477);
nand UO_624 (O_624,N_4824,N_2725);
nor UO_625 (O_625,N_4403,N_3125);
and UO_626 (O_626,N_3701,N_3804);
nand UO_627 (O_627,N_4963,N_2807);
nor UO_628 (O_628,N_3668,N_3084);
nand UO_629 (O_629,N_3405,N_4615);
nand UO_630 (O_630,N_3118,N_4960);
or UO_631 (O_631,N_3657,N_2697);
or UO_632 (O_632,N_4607,N_4753);
nand UO_633 (O_633,N_4464,N_3286);
and UO_634 (O_634,N_3363,N_4801);
or UO_635 (O_635,N_3216,N_2954);
nand UO_636 (O_636,N_2840,N_3004);
and UO_637 (O_637,N_2861,N_2849);
and UO_638 (O_638,N_4947,N_4879);
or UO_639 (O_639,N_2712,N_4716);
nor UO_640 (O_640,N_3243,N_3647);
nand UO_641 (O_641,N_2809,N_3048);
nand UO_642 (O_642,N_3173,N_2634);
xnor UO_643 (O_643,N_4455,N_4100);
or UO_644 (O_644,N_3877,N_3944);
and UO_645 (O_645,N_3894,N_3090);
and UO_646 (O_646,N_4727,N_3617);
nor UO_647 (O_647,N_2986,N_3745);
or UO_648 (O_648,N_2650,N_3886);
or UO_649 (O_649,N_4415,N_4747);
nor UO_650 (O_650,N_2892,N_4158);
xnor UO_651 (O_651,N_3049,N_4358);
and UO_652 (O_652,N_4769,N_4224);
nor UO_653 (O_653,N_3659,N_2940);
nor UO_654 (O_654,N_3538,N_2783);
or UO_655 (O_655,N_4243,N_2745);
nand UO_656 (O_656,N_4808,N_4085);
nor UO_657 (O_657,N_3515,N_4802);
or UO_658 (O_658,N_3772,N_3124);
nor UO_659 (O_659,N_2866,N_4454);
and UO_660 (O_660,N_3015,N_3813);
nand UO_661 (O_661,N_3427,N_2564);
nor UO_662 (O_662,N_2660,N_3268);
or UO_663 (O_663,N_4761,N_4978);
nand UO_664 (O_664,N_4209,N_3073);
and UO_665 (O_665,N_4339,N_2996);
nor UO_666 (O_666,N_2941,N_3926);
nand UO_667 (O_667,N_3854,N_2592);
nor UO_668 (O_668,N_4917,N_2706);
and UO_669 (O_669,N_4080,N_3940);
and UO_670 (O_670,N_4263,N_4115);
nand UO_671 (O_671,N_3135,N_3916);
nor UO_672 (O_672,N_3638,N_3598);
or UO_673 (O_673,N_3146,N_3346);
and UO_674 (O_674,N_4844,N_2723);
or UO_675 (O_675,N_4308,N_4332);
and UO_676 (O_676,N_3597,N_4069);
nand UO_677 (O_677,N_4642,N_3298);
nand UO_678 (O_678,N_3111,N_4197);
nand UO_679 (O_679,N_4673,N_2966);
and UO_680 (O_680,N_3581,N_4382);
or UO_681 (O_681,N_4010,N_4954);
nor UO_682 (O_682,N_3210,N_3052);
xor UO_683 (O_683,N_3337,N_4137);
or UO_684 (O_684,N_4813,N_2685);
or UO_685 (O_685,N_3589,N_4672);
nand UO_686 (O_686,N_4298,N_3254);
and UO_687 (O_687,N_3133,N_2690);
or UO_688 (O_688,N_4034,N_4446);
nor UO_689 (O_689,N_2999,N_2777);
or UO_690 (O_690,N_4545,N_4027);
or UO_691 (O_691,N_3301,N_3526);
nor UO_692 (O_692,N_3593,N_4937);
nand UO_693 (O_693,N_2716,N_2667);
nand UO_694 (O_694,N_3416,N_4482);
or UO_695 (O_695,N_4740,N_3693);
and UO_696 (O_696,N_2743,N_2790);
or UO_697 (O_697,N_2859,N_4234);
nand UO_698 (O_698,N_4014,N_3946);
nor UO_699 (O_699,N_4692,N_3260);
nor UO_700 (O_700,N_4696,N_4586);
nor UO_701 (O_701,N_4305,N_3138);
nor UO_702 (O_702,N_4152,N_4306);
or UO_703 (O_703,N_4969,N_4722);
or UO_704 (O_704,N_3035,N_4401);
nand UO_705 (O_705,N_2879,N_3799);
nand UO_706 (O_706,N_3704,N_4144);
and UO_707 (O_707,N_3788,N_4056);
or UO_708 (O_708,N_3334,N_3464);
nor UO_709 (O_709,N_3215,N_4520);
nor UO_710 (O_710,N_4497,N_3778);
and UO_711 (O_711,N_3456,N_2833);
and UO_712 (O_712,N_4291,N_2760);
and UO_713 (O_713,N_3506,N_4900);
or UO_714 (O_714,N_4919,N_4744);
or UO_715 (O_715,N_3630,N_2823);
or UO_716 (O_716,N_3910,N_2960);
or UO_717 (O_717,N_4626,N_4832);
nand UO_718 (O_718,N_2808,N_3931);
and UO_719 (O_719,N_4574,N_3572);
nand UO_720 (O_720,N_4803,N_3819);
or UO_721 (O_721,N_3367,N_4772);
nand UO_722 (O_722,N_3725,N_4838);
xnor UO_723 (O_723,N_4930,N_2992);
and UO_724 (O_724,N_4017,N_4781);
nor UO_725 (O_725,N_2548,N_4295);
and UO_726 (O_726,N_3895,N_3044);
xor UO_727 (O_727,N_2641,N_2549);
xor UO_728 (O_728,N_3438,N_4659);
nand UO_729 (O_729,N_3471,N_3358);
or UO_730 (O_730,N_3046,N_2957);
or UO_731 (O_731,N_4812,N_2742);
and UO_732 (O_732,N_4743,N_3705);
nand UO_733 (O_733,N_3368,N_2635);
nand UO_734 (O_734,N_2831,N_3958);
and UO_735 (O_735,N_4821,N_4373);
or UO_736 (O_736,N_4649,N_3480);
nand UO_737 (O_737,N_3626,N_4691);
and UO_738 (O_738,N_3942,N_3980);
nor UO_739 (O_739,N_3329,N_2975);
and UO_740 (O_740,N_4909,N_4310);
nand UO_741 (O_741,N_2709,N_2947);
and UO_742 (O_742,N_4139,N_4703);
nor UO_743 (O_743,N_3050,N_4195);
and UO_744 (O_744,N_4223,N_3580);
nor UO_745 (O_745,N_4887,N_3763);
or UO_746 (O_746,N_3461,N_4068);
and UO_747 (O_747,N_3870,N_4334);
nor UO_748 (O_748,N_4015,N_3071);
and UO_749 (O_749,N_3727,N_4050);
and UO_750 (O_750,N_4283,N_4610);
and UO_751 (O_751,N_2917,N_3199);
and UO_752 (O_752,N_3305,N_4742);
nand UO_753 (O_753,N_2836,N_2721);
nor UO_754 (O_754,N_4640,N_2717);
nand UO_755 (O_755,N_3831,N_3088);
nor UO_756 (O_756,N_2594,N_4594);
or UO_757 (O_757,N_3554,N_3616);
nand UO_758 (O_758,N_4274,N_3656);
nand UO_759 (O_759,N_4365,N_3523);
nor UO_760 (O_760,N_4423,N_4598);
nor UO_761 (O_761,N_3386,N_4762);
or UO_762 (O_762,N_3569,N_4411);
nor UO_763 (O_763,N_4466,N_3308);
nand UO_764 (O_764,N_3952,N_4108);
nand UO_765 (O_765,N_4246,N_3988);
nand UO_766 (O_766,N_2915,N_4270);
nor UO_767 (O_767,N_4405,N_3817);
and UO_768 (O_768,N_3290,N_3982);
and UO_769 (O_769,N_4235,N_2593);
and UO_770 (O_770,N_4877,N_3160);
nor UO_771 (O_771,N_4004,N_3396);
nor UO_772 (O_772,N_3332,N_4924);
or UO_773 (O_773,N_4303,N_4565);
or UO_774 (O_774,N_3322,N_3384);
and UO_775 (O_775,N_4407,N_3939);
nor UO_776 (O_776,N_3722,N_2597);
nand UO_777 (O_777,N_3407,N_4955);
or UO_778 (O_778,N_3067,N_4082);
nor UO_779 (O_779,N_4916,N_3176);
and UO_780 (O_780,N_2600,N_4856);
nor UO_781 (O_781,N_4632,N_4073);
and UO_782 (O_782,N_2882,N_3716);
nand UO_783 (O_783,N_4473,N_3399);
and UO_784 (O_784,N_3417,N_2816);
nor UO_785 (O_785,N_4651,N_2643);
and UO_786 (O_786,N_3748,N_4579);
nand UO_787 (O_787,N_3744,N_2842);
or UO_788 (O_788,N_3643,N_4581);
and UO_789 (O_789,N_3157,N_3549);
or UO_790 (O_790,N_3182,N_2714);
or UO_791 (O_791,N_4898,N_3365);
nor UO_792 (O_792,N_4556,N_4143);
nor UO_793 (O_793,N_4052,N_4019);
nand UO_794 (O_794,N_3280,N_4220);
or UO_795 (O_795,N_4271,N_2576);
nor UO_796 (O_796,N_4196,N_3754);
or UO_797 (O_797,N_4712,N_3094);
nand UO_798 (O_798,N_3695,N_2943);
and UO_799 (O_799,N_2985,N_3168);
nor UO_800 (O_800,N_3234,N_3269);
nand UO_801 (O_801,N_4103,N_2605);
or UO_802 (O_802,N_4125,N_4323);
nor UO_803 (O_803,N_3472,N_3691);
and UO_804 (O_804,N_4264,N_4007);
nand UO_805 (O_805,N_2546,N_3131);
or UO_806 (O_806,N_2926,N_4330);
or UO_807 (O_807,N_3018,N_2776);
or UO_808 (O_808,N_3665,N_4252);
or UO_809 (O_809,N_2502,N_4343);
nor UO_810 (O_810,N_3489,N_2988);
nand UO_811 (O_811,N_4848,N_4710);
nor UO_812 (O_812,N_2741,N_4606);
or UO_813 (O_813,N_4765,N_3204);
and UO_814 (O_814,N_2728,N_4767);
nor UO_815 (O_815,N_2663,N_4572);
nor UO_816 (O_816,N_3761,N_4791);
and UO_817 (O_817,N_4033,N_4238);
nand UO_818 (O_818,N_4463,N_2559);
nor UO_819 (O_819,N_4941,N_4506);
nand UO_820 (O_820,N_3040,N_2598);
nor UO_821 (O_821,N_3564,N_3203);
nor UO_822 (O_822,N_4603,N_2604);
and UO_823 (O_823,N_2933,N_2902);
nand UO_824 (O_824,N_3514,N_3648);
and UO_825 (O_825,N_4994,N_3917);
nand UO_826 (O_826,N_3758,N_3552);
or UO_827 (O_827,N_2646,N_3247);
and UO_828 (O_828,N_4087,N_2555);
and UO_829 (O_829,N_3986,N_2981);
and UO_830 (O_830,N_2671,N_2627);
nand UO_831 (O_831,N_4981,N_3162);
and UO_832 (O_832,N_3718,N_3962);
nand UO_833 (O_833,N_4172,N_4850);
nand UO_834 (O_834,N_4391,N_3100);
nand UO_835 (O_835,N_3751,N_3803);
nor UO_836 (O_836,N_4421,N_4650);
nand UO_837 (O_837,N_4964,N_3857);
and UO_838 (O_838,N_3027,N_3376);
or UO_839 (O_839,N_2998,N_3469);
and UO_840 (O_840,N_4633,N_4636);
nand UO_841 (O_841,N_4070,N_2929);
and UO_842 (O_842,N_4785,N_3930);
or UO_843 (O_843,N_3651,N_3449);
nor UO_844 (O_844,N_3848,N_2889);
nand UO_845 (O_845,N_4371,N_4643);
nor UO_846 (O_846,N_3747,N_4145);
or UO_847 (O_847,N_4472,N_3192);
nor UO_848 (O_848,N_3323,N_4729);
nand UO_849 (O_849,N_3420,N_3592);
nand UO_850 (O_850,N_4807,N_2956);
nand UO_851 (O_851,N_4624,N_4872);
nand UO_852 (O_852,N_3288,N_4537);
and UO_853 (O_853,N_4707,N_3501);
or UO_854 (O_854,N_2682,N_3097);
and UO_855 (O_855,N_4711,N_4931);
or UO_856 (O_856,N_4788,N_4957);
nor UO_857 (O_857,N_4950,N_3401);
or UO_858 (O_858,N_4976,N_2724);
nand UO_859 (O_859,N_2707,N_4763);
or UO_860 (O_860,N_4420,N_2547);
nor UO_861 (O_861,N_4136,N_4664);
or UO_862 (O_862,N_2556,N_4166);
and UO_863 (O_863,N_4527,N_2868);
or UO_864 (O_864,N_4376,N_3252);
and UO_865 (O_865,N_3388,N_3153);
or UO_866 (O_866,N_3828,N_3710);
nand UO_867 (O_867,N_2990,N_3850);
nand UO_868 (O_868,N_3774,N_4580);
and UO_869 (O_869,N_4699,N_4825);
or UO_870 (O_870,N_4058,N_2865);
or UO_871 (O_871,N_3655,N_2581);
or UO_872 (O_872,N_2570,N_3715);
nor UO_873 (O_873,N_4042,N_4905);
and UO_874 (O_874,N_4989,N_2550);
nor UO_875 (O_875,N_2529,N_3706);
nand UO_876 (O_876,N_4771,N_4921);
xnor UO_877 (O_877,N_3590,N_4733);
and UO_878 (O_878,N_4128,N_4523);
or UO_879 (O_879,N_2680,N_4037);
or UO_880 (O_880,N_2583,N_3378);
or UO_881 (O_881,N_4648,N_3499);
nand UO_882 (O_882,N_3187,N_4117);
nor UO_883 (O_883,N_4548,N_3834);
xnor UO_884 (O_884,N_4439,N_2819);
or UO_885 (O_885,N_3353,N_3397);
nor UO_886 (O_886,N_3827,N_3312);
nand UO_887 (O_887,N_4131,N_3120);
or UO_888 (O_888,N_4539,N_4869);
nand UO_889 (O_889,N_3969,N_4189);
or UO_890 (O_890,N_3009,N_3667);
or UO_891 (O_891,N_2665,N_2948);
nand UO_892 (O_892,N_4986,N_3446);
nand UO_893 (O_893,N_2797,N_4232);
or UO_894 (O_894,N_4066,N_4795);
and UO_895 (O_895,N_4012,N_3379);
and UO_896 (O_896,N_3081,N_3628);
or UO_897 (O_897,N_3022,N_3373);
or UO_898 (O_898,N_4756,N_4481);
or UO_899 (O_899,N_2737,N_4823);
and UO_900 (O_900,N_4518,N_3884);
nor UO_901 (O_901,N_3106,N_2601);
or UO_902 (O_902,N_4141,N_4647);
nand UO_903 (O_903,N_2774,N_3436);
or UO_904 (O_904,N_4787,N_4840);
and UO_905 (O_905,N_2759,N_3556);
nand UO_906 (O_906,N_3467,N_3463);
nor UO_907 (O_907,N_4000,N_3082);
and UO_908 (O_908,N_4289,N_3178);
nand UO_909 (O_909,N_2751,N_2845);
or UO_910 (O_910,N_4899,N_3919);
or UO_911 (O_911,N_2846,N_4449);
and UO_912 (O_912,N_3839,N_2732);
nor UO_913 (O_913,N_2700,N_4361);
or UO_914 (O_914,N_3824,N_4055);
nand UO_915 (O_915,N_2749,N_3219);
nor UO_916 (O_916,N_3189,N_3152);
nor UO_917 (O_917,N_2834,N_3702);
and UO_918 (O_918,N_4867,N_3762);
and UO_919 (O_919,N_4342,N_4861);
nor UO_920 (O_920,N_2536,N_4945);
and UO_921 (O_921,N_3920,N_2901);
nand UO_922 (O_922,N_4130,N_4908);
or UO_923 (O_923,N_4925,N_3934);
nor UO_924 (O_924,N_4484,N_3458);
xnor UO_925 (O_925,N_3218,N_3905);
xor UO_926 (O_926,N_3410,N_4757);
nand UO_927 (O_927,N_2551,N_4319);
nor UO_928 (O_928,N_3998,N_3237);
or UO_929 (O_929,N_4680,N_4470);
nor UO_930 (O_930,N_4207,N_4500);
and UO_931 (O_931,N_3535,N_4104);
nor UO_932 (O_932,N_4967,N_2873);
or UO_933 (O_933,N_3890,N_4176);
nor UO_934 (O_934,N_3975,N_3374);
or UO_935 (O_935,N_4203,N_4043);
nor UO_936 (O_936,N_4589,N_2613);
and UO_937 (O_937,N_3849,N_3068);
nand UO_938 (O_938,N_3151,N_3733);
and UO_939 (O_939,N_4854,N_4380);
or UO_940 (O_940,N_3865,N_4193);
and UO_941 (O_941,N_3134,N_4003);
nand UO_942 (O_942,N_4608,N_2876);
nor UO_943 (O_943,N_4864,N_4766);
or UO_944 (O_944,N_4932,N_4183);
nand UO_945 (O_945,N_3443,N_3768);
or UO_946 (O_946,N_3995,N_4972);
or UO_947 (O_947,N_3664,N_4735);
nor UO_948 (O_948,N_3618,N_2987);
xnor UO_949 (O_949,N_2718,N_3229);
and UO_950 (O_950,N_3619,N_4406);
nor UO_951 (O_951,N_4719,N_2997);
nor UO_952 (O_952,N_4619,N_4483);
and UO_953 (O_953,N_2526,N_3769);
nor UO_954 (O_954,N_3036,N_3798);
nor UO_955 (O_955,N_4486,N_3929);
and UO_956 (O_956,N_2609,N_4902);
or UO_957 (O_957,N_4859,N_4956);
nor UO_958 (O_958,N_3777,N_3925);
and UO_959 (O_959,N_3906,N_4285);
nor UO_960 (O_960,N_4684,N_4244);
nor UO_961 (O_961,N_2924,N_4452);
nand UO_962 (O_962,N_3950,N_4724);
nor UO_963 (O_963,N_3165,N_4780);
nor UO_964 (O_964,N_2973,N_4776);
nand UO_965 (O_965,N_2904,N_4688);
and UO_966 (O_966,N_3180,N_4853);
or UO_967 (O_967,N_4540,N_3484);
and UO_968 (O_968,N_3031,N_3540);
nor UO_969 (O_969,N_4493,N_3639);
and UO_970 (O_970,N_2715,N_3370);
xnor UO_971 (O_971,N_4555,N_2788);
and UO_972 (O_972,N_4737,N_3136);
nor UO_973 (O_973,N_4336,N_3099);
xnor UO_974 (O_974,N_3105,N_2903);
or UO_975 (O_975,N_4522,N_4432);
or UO_976 (O_976,N_3679,N_4842);
nand UO_977 (O_977,N_2503,N_3430);
nand UO_978 (O_978,N_4560,N_3845);
nor UO_979 (O_979,N_4681,N_3536);
nor UO_980 (O_980,N_3220,N_2918);
and UO_981 (O_981,N_3058,N_2850);
nand UO_982 (O_982,N_3565,N_4728);
nor UO_983 (O_983,N_4883,N_3072);
xnor UO_984 (O_984,N_4046,N_2602);
or UO_985 (O_985,N_4338,N_3309);
xnor UO_986 (O_986,N_2847,N_3577);
and UO_987 (O_987,N_3658,N_3306);
and UO_988 (O_988,N_3823,N_4612);
nor UO_989 (O_989,N_3197,N_2563);
or UO_990 (O_990,N_3766,N_3726);
nand UO_991 (O_991,N_2838,N_3644);
nand UO_992 (O_992,N_2801,N_4890);
nor UO_993 (O_993,N_3500,N_4261);
and UO_994 (O_994,N_3860,N_4739);
and UO_995 (O_995,N_2705,N_3546);
xor UO_996 (O_996,N_4229,N_4168);
nand UO_997 (O_997,N_3113,N_3840);
nor UO_998 (O_998,N_3875,N_2557);
nor UO_999 (O_999,N_2925,N_2898);
endmodule