module basic_750_5000_1000_2_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2527,N_2528,N_2529,N_2531,N_2532,N_2533,N_2534,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2545,N_2547,N_2548,N_2550,N_2551,N_2552,N_2553,N_2554,N_2558,N_2559,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2585,N_2586,N_2587,N_2590,N_2592,N_2593,N_2594,N_2595,N_2596,N_2598,N_2599,N_2601,N_2602,N_2603,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2614,N_2615,N_2616,N_2617,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2649,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2667,N_2668,N_2669,N_2672,N_2674,N_2675,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2692,N_2693,N_2694,N_2697,N_2698,N_2699,N_2700,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2709,N_2710,N_2711,N_2713,N_2714,N_2717,N_2718,N_2719,N_2720,N_2721,N_2723,N_2724,N_2725,N_2726,N_2728,N_2729,N_2730,N_2731,N_2732,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2742,N_2744,N_2745,N_2746,N_2747,N_2748,N_2750,N_2752,N_2753,N_2755,N_2757,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2769,N_2770,N_2771,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2792,N_2794,N_2795,N_2797,N_2799,N_2800,N_2802,N_2803,N_2804,N_2805,N_2806,N_2808,N_2810,N_2812,N_2813,N_2814,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2859,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2879,N_2881,N_2882,N_2883,N_2884,N_2885,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2909,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2931,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2947,N_2948,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2973,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2985,N_2988,N_2989,N_2991,N_2992,N_2994,N_2995,N_2996,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3006,N_3007,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3041,N_3042,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3086,N_3087,N_3088,N_3089,N_3091,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3100,N_3101,N_3102,N_3104,N_3105,N_3106,N_3107,N_3109,N_3110,N_3112,N_3114,N_3116,N_3117,N_3118,N_3119,N_3120,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3136,N_3137,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3149,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3164,N_3165,N_3166,N_3168,N_3170,N_3171,N_3173,N_3174,N_3175,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3192,N_3193,N_3195,N_3196,N_3197,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3207,N_3208,N_3211,N_3212,N_3214,N_3215,N_3217,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3241,N_3242,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3281,N_3283,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3293,N_3294,N_3295,N_3296,N_3301,N_3303,N_3305,N_3306,N_3308,N_3309,N_3312,N_3313,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3326,N_3327,N_3328,N_3329,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3352,N_3353,N_3357,N_3358,N_3359,N_3360,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3369,N_3370,N_3372,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3383,N_3385,N_3386,N_3387,N_3388,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3401,N_3402,N_3403,N_3404,N_3405,N_3407,N_3408,N_3410,N_3412,N_3413,N_3414,N_3416,N_3417,N_3419,N_3420,N_3422,N_3423,N_3424,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3436,N_3437,N_3438,N_3439,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3450,N_3452,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3462,N_3463,N_3464,N_3465,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3489,N_3492,N_3493,N_3494,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3516,N_3517,N_3518,N_3520,N_3521,N_3522,N_3524,N_3525,N_3527,N_3529,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3539,N_3540,N_3541,N_3542,N_3543,N_3545,N_3546,N_3548,N_3549,N_3550,N_3551,N_3552,N_3554,N_3555,N_3556,N_3557,N_3558,N_3560,N_3561,N_3562,N_3563,N_3564,N_3566,N_3567,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3585,N_3586,N_3588,N_3589,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3601,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3611,N_3613,N_3614,N_3615,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3660,N_3661,N_3663,N_3664,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3681,N_3682,N_3683,N_3684,N_3685,N_3687,N_3688,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3717,N_3718,N_3721,N_3722,N_3723,N_3724,N_3725,N_3727,N_3729,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3743,N_3744,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3754,N_3755,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3778,N_3779,N_3780,N_3781,N_3783,N_3785,N_3786,N_3787,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3807,N_3808,N_3809,N_3810,N_3811,N_3813,N_3815,N_3816,N_3817,N_3818,N_3821,N_3822,N_3823,N_3824,N_3826,N_3828,N_3829,N_3831,N_3832,N_3833,N_3834,N_3836,N_3837,N_3842,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3857,N_3858,N_3859,N_3860,N_3861,N_3863,N_3864,N_3867,N_3868,N_3869,N_3870,N_3873,N_3874,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3888,N_3890,N_3891,N_3892,N_3893,N_3894,N_3896,N_3897,N_3899,N_3900,N_3901,N_3903,N_3905,N_3906,N_3907,N_3908,N_3909,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3920,N_3923,N_3924,N_3926,N_3927,N_3929,N_3931,N_3932,N_3933,N_3934,N_3936,N_3938,N_3939,N_3940,N_3942,N_3943,N_3944,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3994,N_3995,N_3996,N_3997,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4008,N_4009,N_4010,N_4011,N_4012,N_4014,N_4015,N_4016,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4029,N_4031,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4040,N_4041,N_4042,N_4044,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4062,N_4063,N_4064,N_4065,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4080,N_4081,N_4082,N_4083,N_4084,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4112,N_4113,N_4114,N_4116,N_4117,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4134,N_4135,N_4136,N_4138,N_4139,N_4141,N_4142,N_4143,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4152,N_4154,N_4155,N_4157,N_4158,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4173,N_4174,N_4176,N_4177,N_4178,N_4180,N_4181,N_4182,N_4183,N_4184,N_4186,N_4187,N_4188,N_4190,N_4191,N_4193,N_4194,N_4195,N_4196,N_4197,N_4200,N_4201,N_4203,N_4204,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4219,N_4220,N_4221,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4230,N_4231,N_4233,N_4234,N_4235,N_4236,N_4237,N_4239,N_4240,N_4241,N_4242,N_4244,N_4245,N_4246,N_4247,N_4249,N_4250,N_4251,N_4253,N_4254,N_4255,N_4256,N_4258,N_4259,N_4261,N_4262,N_4264,N_4265,N_4266,N_4268,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4306,N_4307,N_4308,N_4309,N_4311,N_4312,N_4314,N_4315,N_4316,N_4319,N_4321,N_4323,N_4324,N_4325,N_4326,N_4327,N_4330,N_4331,N_4333,N_4334,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4350,N_4351,N_4352,N_4353,N_4354,N_4357,N_4358,N_4359,N_4360,N_4364,N_4366,N_4367,N_4370,N_4371,N_4373,N_4374,N_4376,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4407,N_4408,N_4409,N_4410,N_4412,N_4413,N_4415,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4424,N_4425,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4435,N_4436,N_4437,N_4438,N_4440,N_4441,N_4442,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4458,N_4459,N_4460,N_4462,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4480,N_4481,N_4482,N_4484,N_4486,N_4487,N_4488,N_4489,N_4491,N_4492,N_4494,N_4495,N_4496,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4516,N_4517,N_4518,N_4519,N_4521,N_4523,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4532,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4560,N_4561,N_4562,N_4563,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4586,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4598,N_4599,N_4600,N_4601,N_4603,N_4604,N_4606,N_4607,N_4608,N_4610,N_4611,N_4613,N_4614,N_4615,N_4617,N_4618,N_4619,N_4620,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4667,N_4669,N_4670,N_4671,N_4672,N_4673,N_4675,N_4676,N_4677,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4699,N_4700,N_4701,N_4702,N_4703,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4713,N_4715,N_4718,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4731,N_4732,N_4733,N_4734,N_4736,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4766,N_4767,N_4769,N_4771,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4788,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4808,N_4809,N_4810,N_4811,N_4812,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4822,N_4823,N_4825,N_4826,N_4827,N_4828,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4840,N_4842,N_4843,N_4844,N_4845,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4859,N_4862,N_4863,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4876,N_4877,N_4878,N_4879,N_4880,N_4882,N_4883,N_4884,N_4885,N_4887,N_4888,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4918,N_4919,N_4921,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4948,N_4949,N_4950,N_4951,N_4953,N_4954,N_4955,N_4958,N_4961,N_4962,N_4963,N_4964,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4977,N_4978,N_4980,N_4982,N_4985,N_4987,N_4988,N_4989,N_4990,N_4992,N_4993,N_4994,N_4995,N_4997,N_4998,N_4999;
nor U0 (N_0,In_636,In_604);
nand U1 (N_1,In_724,In_329);
nor U2 (N_2,In_77,In_109);
and U3 (N_3,In_136,In_434);
xor U4 (N_4,In_119,In_677);
and U5 (N_5,In_696,In_590);
nand U6 (N_6,In_131,In_215);
nor U7 (N_7,In_33,In_281);
nor U8 (N_8,In_229,In_314);
nor U9 (N_9,In_436,In_377);
or U10 (N_10,In_466,In_691);
or U11 (N_11,In_482,In_528);
nand U12 (N_12,In_558,In_694);
nand U13 (N_13,In_236,In_405);
nor U14 (N_14,In_397,In_239);
or U15 (N_15,In_158,In_338);
nand U16 (N_16,In_689,In_449);
nand U17 (N_17,In_633,In_246);
or U18 (N_18,In_61,In_10);
or U19 (N_19,In_627,In_453);
or U20 (N_20,In_626,In_362);
nor U21 (N_21,In_473,In_172);
nor U22 (N_22,In_7,In_403);
nand U23 (N_23,In_617,In_524);
nor U24 (N_24,In_274,In_656);
xnor U25 (N_25,In_225,In_511);
or U26 (N_26,In_634,In_97);
nand U27 (N_27,In_704,In_731);
nand U28 (N_28,In_657,In_409);
nor U29 (N_29,In_468,In_619);
nand U30 (N_30,In_586,In_115);
nand U31 (N_31,In_463,In_170);
or U32 (N_32,In_303,In_267);
nand U33 (N_33,In_536,In_85);
nor U34 (N_34,In_418,In_676);
nand U35 (N_35,In_448,In_242);
nor U36 (N_36,In_624,In_272);
nor U37 (N_37,In_530,In_262);
and U38 (N_38,In_697,In_67);
or U39 (N_39,In_173,In_166);
nor U40 (N_40,In_271,In_486);
nand U41 (N_41,In_349,In_213);
and U42 (N_42,In_143,In_576);
nor U43 (N_43,In_606,In_335);
and U44 (N_44,In_682,In_395);
nor U45 (N_45,In_415,In_317);
nand U46 (N_46,In_160,In_59);
or U47 (N_47,In_183,In_52);
and U48 (N_48,In_654,In_333);
nand U49 (N_49,In_319,In_145);
nand U50 (N_50,In_108,In_232);
nand U51 (N_51,In_37,In_388);
or U52 (N_52,In_578,In_141);
nand U53 (N_53,In_735,In_713);
nand U54 (N_54,In_614,In_568);
nand U55 (N_55,In_457,In_48);
xor U56 (N_56,In_561,In_51);
and U57 (N_57,In_423,In_599);
nand U58 (N_58,In_112,In_197);
and U59 (N_59,In_104,In_185);
nor U60 (N_60,In_135,In_219);
nand U61 (N_61,In_413,In_653);
and U62 (N_62,In_547,In_212);
and U63 (N_63,In_254,In_16);
and U64 (N_64,In_113,In_137);
nand U65 (N_65,In_357,In_666);
nand U66 (N_66,In_323,In_261);
nor U67 (N_67,In_484,In_566);
nor U68 (N_68,In_419,In_479);
nor U69 (N_69,In_149,In_35);
nand U70 (N_70,In_609,In_483);
and U71 (N_71,In_584,In_257);
and U72 (N_72,In_430,In_380);
nor U73 (N_73,In_629,In_56);
nor U74 (N_74,In_348,In_569);
and U75 (N_75,In_649,In_80);
nor U76 (N_76,In_256,In_305);
nor U77 (N_77,In_501,In_121);
nand U78 (N_78,In_543,In_527);
xnor U79 (N_79,In_575,In_640);
or U80 (N_80,In_147,In_114);
xor U81 (N_81,In_22,In_700);
nand U82 (N_82,In_517,In_712);
and U83 (N_83,In_675,In_346);
nor U84 (N_84,In_275,In_458);
and U85 (N_85,In_407,In_310);
nand U86 (N_86,In_680,In_485);
xnor U87 (N_87,In_435,In_608);
or U88 (N_88,In_294,In_45);
and U89 (N_89,In_737,In_628);
nor U90 (N_90,In_122,In_188);
nor U91 (N_91,In_559,In_643);
nand U92 (N_92,In_467,In_710);
nand U93 (N_93,In_596,In_273);
nor U94 (N_94,In_709,In_646);
or U95 (N_95,In_350,In_445);
nor U96 (N_96,In_295,In_43);
or U97 (N_97,In_107,In_662);
nor U98 (N_98,In_76,In_652);
nor U99 (N_99,In_499,In_605);
nor U100 (N_100,In_553,In_386);
and U101 (N_101,In_444,In_417);
nor U102 (N_102,In_345,In_655);
nor U103 (N_103,In_301,In_320);
and U104 (N_104,In_723,In_86);
and U105 (N_105,In_644,In_204);
nand U106 (N_106,In_111,In_332);
or U107 (N_107,In_138,In_199);
nor U108 (N_108,In_503,In_732);
and U109 (N_109,In_456,In_99);
and U110 (N_110,In_706,In_412);
or U111 (N_111,In_537,In_193);
nor U112 (N_112,In_163,In_541);
nor U113 (N_113,In_206,In_460);
nand U114 (N_114,In_390,In_279);
or U115 (N_115,In_625,In_162);
nand U116 (N_116,In_580,In_542);
or U117 (N_117,In_523,In_440);
or U118 (N_118,In_152,In_420);
and U119 (N_119,In_546,In_304);
nor U120 (N_120,In_438,In_39);
xnor U121 (N_121,In_18,In_176);
nand U122 (N_122,In_169,In_690);
and U123 (N_123,In_668,In_105);
or U124 (N_124,In_291,In_70);
or U125 (N_125,In_9,In_360);
nor U126 (N_126,In_302,In_356);
or U127 (N_127,In_285,In_481);
and U128 (N_128,In_30,In_159);
or U129 (N_129,In_32,In_5);
and U130 (N_130,In_711,In_354);
and U131 (N_131,In_366,In_591);
and U132 (N_132,In_671,In_480);
nand U133 (N_133,In_327,In_579);
xor U134 (N_134,In_359,In_607);
nand U135 (N_135,In_286,In_422);
nand U136 (N_136,In_554,In_245);
and U137 (N_137,In_521,In_540);
nor U138 (N_138,In_638,In_526);
nor U139 (N_139,In_278,In_489);
nor U140 (N_140,In_631,In_741);
and U141 (N_141,In_707,In_630);
and U142 (N_142,In_736,In_398);
nor U143 (N_143,In_178,In_308);
and U144 (N_144,In_464,In_17);
or U145 (N_145,In_117,In_341);
or U146 (N_146,In_572,In_223);
or U147 (N_147,In_148,In_637);
nand U148 (N_148,In_134,In_340);
nor U149 (N_149,In_299,In_698);
nand U150 (N_150,In_62,In_92);
nand U151 (N_151,In_125,In_684);
nand U152 (N_152,In_534,In_41);
nor U153 (N_153,In_715,In_703);
nand U154 (N_154,In_402,In_227);
nand U155 (N_155,In_410,In_392);
and U156 (N_156,In_19,In_462);
nand U157 (N_157,In_177,In_205);
xnor U158 (N_158,In_365,In_408);
and U159 (N_159,In_98,In_4);
or U160 (N_160,In_47,In_693);
and U161 (N_161,In_451,In_25);
and U162 (N_162,In_520,In_347);
and U163 (N_163,In_667,In_632);
or U164 (N_164,In_368,In_165);
and U165 (N_165,In_505,In_202);
nand U166 (N_166,In_83,In_529);
and U167 (N_167,In_384,In_182);
or U168 (N_168,In_2,In_729);
and U169 (N_169,In_248,In_93);
and U170 (N_170,In_701,In_573);
nand U171 (N_171,In_730,In_747);
nand U172 (N_172,In_132,In_476);
nand U173 (N_173,In_322,In_492);
xor U174 (N_174,In_582,In_600);
nor U175 (N_175,In_683,In_452);
nor U176 (N_176,In_391,In_151);
or U177 (N_177,In_123,In_613);
nand U178 (N_178,In_6,In_53);
or U179 (N_179,In_54,In_400);
nor U180 (N_180,In_574,In_150);
and U181 (N_181,In_21,In_324);
and U182 (N_182,In_396,In_714);
nor U183 (N_183,In_494,In_725);
or U184 (N_184,In_387,In_316);
or U185 (N_185,In_510,In_555);
or U186 (N_186,In_156,In_352);
or U187 (N_187,In_300,In_69);
nand U188 (N_188,In_531,In_669);
nand U189 (N_189,In_404,In_174);
nor U190 (N_190,In_1,In_42);
nor U191 (N_191,In_414,In_425);
or U192 (N_192,In_321,In_563);
nor U193 (N_193,In_31,In_269);
nor U194 (N_194,In_718,In_3);
nor U195 (N_195,In_118,In_331);
and U196 (N_196,In_611,In_506);
nand U197 (N_197,In_658,In_218);
and U198 (N_198,In_88,In_597);
or U199 (N_199,In_551,In_194);
nand U200 (N_200,In_101,In_616);
and U201 (N_201,In_369,In_594);
and U202 (N_202,In_57,In_589);
nor U203 (N_203,In_749,In_234);
nand U204 (N_204,In_361,In_296);
or U205 (N_205,In_210,In_65);
or U206 (N_206,In_726,In_154);
nor U207 (N_207,In_337,In_595);
and U208 (N_208,In_251,In_90);
nor U209 (N_209,In_381,In_334);
xor U210 (N_210,In_153,In_393);
nand U211 (N_211,In_238,In_355);
nor U212 (N_212,In_249,In_13);
nor U213 (N_213,In_233,In_29);
or U214 (N_214,In_424,In_120);
xor U215 (N_215,In_161,In_328);
nand U216 (N_216,In_641,In_201);
nor U217 (N_217,In_311,In_686);
or U218 (N_218,In_344,In_96);
and U219 (N_219,In_255,In_144);
nand U220 (N_220,In_214,In_209);
nand U221 (N_221,In_127,In_237);
nor U222 (N_222,In_465,In_581);
nand U223 (N_223,In_247,In_727);
nand U224 (N_224,In_263,In_203);
nor U225 (N_225,In_661,In_73);
xor U226 (N_226,In_642,In_461);
or U227 (N_227,In_488,In_235);
nor U228 (N_228,In_376,In_487);
nor U229 (N_229,In_140,In_622);
and U230 (N_230,In_439,In_89);
and U231 (N_231,In_550,In_495);
nand U232 (N_232,In_241,In_678);
or U233 (N_233,In_720,In_189);
nand U234 (N_234,In_187,In_372);
nand U235 (N_235,In_516,In_26);
nand U236 (N_236,In_78,In_639);
and U237 (N_237,In_375,In_217);
and U238 (N_238,In_343,In_94);
nor U239 (N_239,In_116,In_363);
or U240 (N_240,In_196,In_721);
nand U241 (N_241,In_744,In_593);
or U242 (N_242,In_130,In_318);
or U243 (N_243,In_307,In_28);
or U244 (N_244,In_230,In_157);
nand U245 (N_245,In_211,In_133);
nor U246 (N_246,In_401,In_474);
or U247 (N_247,In_44,In_562);
and U248 (N_248,In_374,In_184);
or U249 (N_249,In_181,In_84);
nor U250 (N_250,In_50,In_496);
and U251 (N_251,In_383,In_441);
nand U252 (N_252,In_164,In_443);
nor U253 (N_253,In_367,In_588);
nand U254 (N_254,In_175,In_282);
or U255 (N_255,In_406,In_469);
nor U256 (N_256,In_437,In_81);
nand U257 (N_257,In_567,In_733);
nand U258 (N_258,In_674,In_645);
nand U259 (N_259,In_297,In_250);
nor U260 (N_260,In_259,In_538);
and U261 (N_261,In_128,In_8);
or U262 (N_262,In_665,In_244);
or U263 (N_263,In_618,In_60);
and U264 (N_264,In_411,In_399);
or U265 (N_265,In_385,In_167);
or U266 (N_266,In_179,In_186);
and U267 (N_267,In_270,In_472);
nand U268 (N_268,In_447,In_284);
nand U269 (N_269,In_592,In_38);
nor U270 (N_270,In_478,In_240);
nand U271 (N_271,In_601,In_429);
nor U272 (N_272,In_577,In_0);
and U273 (N_273,In_265,In_716);
nor U274 (N_274,In_717,In_312);
nand U275 (N_275,In_427,In_748);
nor U276 (N_276,In_353,In_146);
nor U277 (N_277,In_293,In_659);
or U278 (N_278,In_243,In_40);
or U279 (N_279,In_564,In_535);
or U280 (N_280,In_428,In_621);
and U281 (N_281,In_110,In_557);
nand U282 (N_282,In_740,In_378);
nor U283 (N_283,In_502,In_745);
or U284 (N_284,In_277,In_71);
and U285 (N_285,In_519,In_695);
nand U286 (N_286,In_106,In_705);
nor U287 (N_287,In_339,In_364);
nor U288 (N_288,In_738,In_224);
or U289 (N_289,In_455,In_512);
or U290 (N_290,In_34,In_252);
or U291 (N_291,In_103,In_679);
or U292 (N_292,In_195,In_260);
or U293 (N_293,In_306,In_11);
and U294 (N_294,In_507,In_287);
nand U295 (N_295,In_55,In_533);
xor U296 (N_296,In_620,In_598);
nand U297 (N_297,In_615,In_504);
nor U298 (N_298,In_23,In_216);
or U299 (N_299,In_226,In_565);
or U300 (N_300,In_647,In_685);
nand U301 (N_301,In_708,In_288);
or U302 (N_302,In_743,In_500);
or U303 (N_303,In_58,In_522);
nor U304 (N_304,In_155,In_49);
nand U305 (N_305,In_681,In_446);
nor U306 (N_306,In_266,In_471);
or U307 (N_307,In_15,In_289);
and U308 (N_308,In_228,In_63);
nand U309 (N_309,In_493,In_431);
or U310 (N_310,In_664,In_651);
nor U311 (N_311,In_687,In_450);
nor U312 (N_312,In_102,In_82);
and U313 (N_313,In_142,In_192);
xnor U314 (N_314,In_75,In_513);
or U315 (N_315,In_648,In_351);
nor U316 (N_316,In_309,In_497);
or U317 (N_317,In_280,In_198);
or U318 (N_318,In_742,In_548);
nand U319 (N_319,In_722,In_129);
nand U320 (N_320,In_36,In_525);
nand U321 (N_321,In_91,In_610);
nor U322 (N_322,In_552,In_389);
nor U323 (N_323,In_673,In_699);
nor U324 (N_324,In_514,In_24);
nor U325 (N_325,In_688,In_68);
and U326 (N_326,In_454,In_587);
xor U327 (N_327,In_623,In_475);
or U328 (N_328,In_139,In_191);
or U329 (N_329,In_746,In_180);
nand U330 (N_330,In_571,In_222);
nor U331 (N_331,In_258,In_545);
nor U332 (N_332,In_325,In_370);
nor U333 (N_333,In_79,In_544);
and U334 (N_334,In_421,In_433);
and U335 (N_335,In_394,In_602);
nand U336 (N_336,In_200,In_416);
nand U337 (N_337,In_459,In_379);
nor U338 (N_338,In_20,In_231);
or U339 (N_339,In_432,In_298);
xor U340 (N_340,In_382,In_64);
nor U341 (N_341,In_560,In_14);
and U342 (N_342,In_508,In_27);
nand U343 (N_343,In_283,In_126);
and U344 (N_344,In_491,In_692);
and U345 (N_345,In_326,In_208);
nor U346 (N_346,In_74,In_336);
or U347 (N_347,In_12,In_171);
or U348 (N_348,In_498,In_207);
and U349 (N_349,In_371,In_268);
and U350 (N_350,In_539,In_221);
nor U351 (N_351,In_672,In_168);
nor U352 (N_352,In_264,In_253);
and U353 (N_353,In_719,In_95);
and U354 (N_354,In_585,In_734);
and U355 (N_355,In_532,In_549);
and U356 (N_356,In_373,In_426);
and U357 (N_357,In_490,In_509);
nand U358 (N_358,In_290,In_518);
or U359 (N_359,In_660,In_190);
or U360 (N_360,In_650,In_477);
or U361 (N_361,In_635,In_663);
nand U362 (N_362,In_330,In_66);
or U363 (N_363,In_72,In_702);
nand U364 (N_364,In_313,In_46);
and U365 (N_365,In_276,In_124);
nor U366 (N_366,In_292,In_739);
nand U367 (N_367,In_442,In_670);
nand U368 (N_368,In_728,In_612);
nand U369 (N_369,In_87,In_220);
or U370 (N_370,In_100,In_603);
or U371 (N_371,In_470,In_570);
nor U372 (N_372,In_315,In_342);
and U373 (N_373,In_515,In_556);
or U374 (N_374,In_358,In_583);
nand U375 (N_375,In_499,In_263);
or U376 (N_376,In_362,In_158);
and U377 (N_377,In_248,In_258);
nor U378 (N_378,In_141,In_528);
or U379 (N_379,In_227,In_75);
nor U380 (N_380,In_240,In_536);
nand U381 (N_381,In_221,In_680);
nor U382 (N_382,In_607,In_218);
nand U383 (N_383,In_513,In_646);
or U384 (N_384,In_500,In_550);
and U385 (N_385,In_403,In_676);
nand U386 (N_386,In_612,In_611);
and U387 (N_387,In_526,In_462);
nand U388 (N_388,In_275,In_627);
and U389 (N_389,In_416,In_593);
nor U390 (N_390,In_570,In_366);
or U391 (N_391,In_23,In_192);
or U392 (N_392,In_294,In_248);
nor U393 (N_393,In_480,In_133);
or U394 (N_394,In_83,In_437);
nor U395 (N_395,In_611,In_158);
nor U396 (N_396,In_312,In_354);
and U397 (N_397,In_490,In_567);
and U398 (N_398,In_642,In_463);
nor U399 (N_399,In_436,In_555);
or U400 (N_400,In_137,In_575);
nand U401 (N_401,In_254,In_39);
or U402 (N_402,In_611,In_650);
and U403 (N_403,In_320,In_572);
nand U404 (N_404,In_642,In_620);
or U405 (N_405,In_322,In_200);
or U406 (N_406,In_253,In_625);
or U407 (N_407,In_726,In_693);
or U408 (N_408,In_640,In_693);
nand U409 (N_409,In_731,In_512);
and U410 (N_410,In_24,In_612);
nand U411 (N_411,In_508,In_649);
nor U412 (N_412,In_392,In_78);
and U413 (N_413,In_531,In_677);
and U414 (N_414,In_320,In_238);
and U415 (N_415,In_656,In_90);
nor U416 (N_416,In_492,In_327);
nor U417 (N_417,In_8,In_360);
or U418 (N_418,In_303,In_424);
nand U419 (N_419,In_185,In_169);
and U420 (N_420,In_93,In_129);
nor U421 (N_421,In_566,In_305);
and U422 (N_422,In_469,In_717);
or U423 (N_423,In_246,In_428);
and U424 (N_424,In_717,In_323);
nand U425 (N_425,In_727,In_166);
and U426 (N_426,In_656,In_582);
nand U427 (N_427,In_669,In_527);
nor U428 (N_428,In_66,In_573);
and U429 (N_429,In_431,In_190);
and U430 (N_430,In_600,In_411);
or U431 (N_431,In_348,In_657);
and U432 (N_432,In_36,In_77);
nor U433 (N_433,In_194,In_715);
or U434 (N_434,In_347,In_643);
nor U435 (N_435,In_307,In_222);
or U436 (N_436,In_370,In_614);
and U437 (N_437,In_159,In_522);
and U438 (N_438,In_475,In_717);
and U439 (N_439,In_278,In_363);
or U440 (N_440,In_703,In_275);
nor U441 (N_441,In_47,In_90);
or U442 (N_442,In_329,In_603);
and U443 (N_443,In_266,In_642);
nor U444 (N_444,In_440,In_227);
or U445 (N_445,In_638,In_503);
nand U446 (N_446,In_200,In_523);
nand U447 (N_447,In_188,In_562);
and U448 (N_448,In_412,In_270);
or U449 (N_449,In_353,In_101);
nor U450 (N_450,In_227,In_78);
nand U451 (N_451,In_471,In_573);
nor U452 (N_452,In_576,In_748);
nor U453 (N_453,In_558,In_444);
nor U454 (N_454,In_304,In_630);
nand U455 (N_455,In_235,In_426);
and U456 (N_456,In_86,In_469);
or U457 (N_457,In_285,In_86);
nand U458 (N_458,In_502,In_653);
or U459 (N_459,In_530,In_301);
or U460 (N_460,In_450,In_387);
and U461 (N_461,In_408,In_738);
nand U462 (N_462,In_282,In_211);
nand U463 (N_463,In_37,In_382);
nand U464 (N_464,In_732,In_117);
nand U465 (N_465,In_467,In_470);
nor U466 (N_466,In_637,In_223);
nor U467 (N_467,In_95,In_569);
and U468 (N_468,In_251,In_656);
and U469 (N_469,In_456,In_317);
nor U470 (N_470,In_223,In_556);
or U471 (N_471,In_155,In_454);
and U472 (N_472,In_321,In_219);
or U473 (N_473,In_506,In_467);
and U474 (N_474,In_568,In_208);
nor U475 (N_475,In_452,In_612);
nor U476 (N_476,In_378,In_481);
or U477 (N_477,In_313,In_414);
nand U478 (N_478,In_478,In_458);
and U479 (N_479,In_469,In_243);
nor U480 (N_480,In_385,In_703);
or U481 (N_481,In_179,In_684);
nor U482 (N_482,In_143,In_514);
nand U483 (N_483,In_529,In_665);
nor U484 (N_484,In_60,In_266);
nand U485 (N_485,In_394,In_22);
and U486 (N_486,In_1,In_625);
nand U487 (N_487,In_558,In_185);
nor U488 (N_488,In_610,In_331);
nand U489 (N_489,In_644,In_178);
and U490 (N_490,In_232,In_368);
or U491 (N_491,In_285,In_549);
or U492 (N_492,In_740,In_386);
nand U493 (N_493,In_473,In_307);
nor U494 (N_494,In_553,In_603);
nor U495 (N_495,In_286,In_415);
and U496 (N_496,In_472,In_141);
or U497 (N_497,In_745,In_131);
and U498 (N_498,In_501,In_284);
or U499 (N_499,In_409,In_593);
and U500 (N_500,In_409,In_344);
nand U501 (N_501,In_530,In_537);
and U502 (N_502,In_486,In_348);
nand U503 (N_503,In_657,In_304);
and U504 (N_504,In_318,In_153);
or U505 (N_505,In_406,In_260);
or U506 (N_506,In_516,In_267);
and U507 (N_507,In_348,In_666);
nor U508 (N_508,In_157,In_92);
and U509 (N_509,In_87,In_221);
nor U510 (N_510,In_95,In_284);
nand U511 (N_511,In_309,In_624);
nand U512 (N_512,In_736,In_83);
or U513 (N_513,In_428,In_459);
and U514 (N_514,In_4,In_325);
and U515 (N_515,In_329,In_205);
or U516 (N_516,In_108,In_415);
nand U517 (N_517,In_451,In_316);
nand U518 (N_518,In_548,In_495);
nor U519 (N_519,In_622,In_387);
or U520 (N_520,In_550,In_716);
nand U521 (N_521,In_360,In_204);
nor U522 (N_522,In_82,In_448);
nand U523 (N_523,In_272,In_125);
or U524 (N_524,In_157,In_704);
or U525 (N_525,In_27,In_380);
xor U526 (N_526,In_669,In_650);
nor U527 (N_527,In_256,In_180);
or U528 (N_528,In_744,In_476);
or U529 (N_529,In_425,In_375);
or U530 (N_530,In_683,In_607);
and U531 (N_531,In_696,In_561);
nand U532 (N_532,In_670,In_51);
and U533 (N_533,In_606,In_333);
and U534 (N_534,In_748,In_672);
nor U535 (N_535,In_249,In_329);
or U536 (N_536,In_744,In_484);
and U537 (N_537,In_644,In_371);
and U538 (N_538,In_390,In_394);
nand U539 (N_539,In_509,In_693);
nor U540 (N_540,In_62,In_6);
nor U541 (N_541,In_671,In_104);
nand U542 (N_542,In_629,In_721);
and U543 (N_543,In_512,In_663);
or U544 (N_544,In_274,In_55);
and U545 (N_545,In_672,In_150);
nand U546 (N_546,In_360,In_371);
nand U547 (N_547,In_184,In_601);
or U548 (N_548,In_53,In_459);
nor U549 (N_549,In_304,In_582);
nor U550 (N_550,In_16,In_544);
or U551 (N_551,In_577,In_17);
nor U552 (N_552,In_24,In_540);
nor U553 (N_553,In_147,In_190);
and U554 (N_554,In_438,In_449);
or U555 (N_555,In_300,In_592);
and U556 (N_556,In_544,In_76);
nand U557 (N_557,In_329,In_683);
and U558 (N_558,In_92,In_122);
or U559 (N_559,In_545,In_321);
nand U560 (N_560,In_132,In_245);
or U561 (N_561,In_252,In_645);
nor U562 (N_562,In_567,In_661);
nor U563 (N_563,In_401,In_318);
and U564 (N_564,In_730,In_43);
nand U565 (N_565,In_542,In_609);
nor U566 (N_566,In_626,In_69);
and U567 (N_567,In_123,In_279);
nor U568 (N_568,In_499,In_346);
or U569 (N_569,In_203,In_696);
nand U570 (N_570,In_174,In_323);
or U571 (N_571,In_23,In_341);
nor U572 (N_572,In_208,In_112);
or U573 (N_573,In_357,In_274);
nor U574 (N_574,In_557,In_494);
and U575 (N_575,In_89,In_77);
nor U576 (N_576,In_477,In_488);
nor U577 (N_577,In_680,In_650);
nor U578 (N_578,In_236,In_207);
and U579 (N_579,In_599,In_634);
and U580 (N_580,In_452,In_553);
nand U581 (N_581,In_158,In_702);
nor U582 (N_582,In_574,In_583);
or U583 (N_583,In_473,In_413);
and U584 (N_584,In_727,In_512);
nand U585 (N_585,In_244,In_701);
and U586 (N_586,In_373,In_439);
nor U587 (N_587,In_573,In_314);
or U588 (N_588,In_405,In_158);
xnor U589 (N_589,In_734,In_334);
nor U590 (N_590,In_16,In_155);
and U591 (N_591,In_257,In_199);
and U592 (N_592,In_693,In_4);
nor U593 (N_593,In_338,In_466);
or U594 (N_594,In_129,In_748);
or U595 (N_595,In_600,In_399);
or U596 (N_596,In_717,In_33);
or U597 (N_597,In_66,In_666);
nand U598 (N_598,In_146,In_539);
nor U599 (N_599,In_376,In_88);
or U600 (N_600,In_421,In_531);
and U601 (N_601,In_552,In_381);
nand U602 (N_602,In_267,In_121);
nand U603 (N_603,In_323,In_14);
and U604 (N_604,In_637,In_370);
nand U605 (N_605,In_313,In_61);
and U606 (N_606,In_210,In_185);
nor U607 (N_607,In_268,In_443);
and U608 (N_608,In_644,In_506);
nand U609 (N_609,In_216,In_357);
and U610 (N_610,In_158,In_324);
nor U611 (N_611,In_142,In_86);
nand U612 (N_612,In_477,In_105);
nor U613 (N_613,In_10,In_698);
and U614 (N_614,In_606,In_237);
or U615 (N_615,In_347,In_390);
nand U616 (N_616,In_592,In_215);
nor U617 (N_617,In_73,In_175);
or U618 (N_618,In_272,In_410);
or U619 (N_619,In_457,In_37);
nand U620 (N_620,In_309,In_116);
and U621 (N_621,In_325,In_292);
nand U622 (N_622,In_344,In_347);
nor U623 (N_623,In_67,In_110);
nand U624 (N_624,In_640,In_214);
or U625 (N_625,In_61,In_562);
nor U626 (N_626,In_68,In_337);
nand U627 (N_627,In_454,In_473);
or U628 (N_628,In_521,In_351);
or U629 (N_629,In_119,In_712);
nand U630 (N_630,In_154,In_226);
nand U631 (N_631,In_380,In_439);
nand U632 (N_632,In_513,In_611);
or U633 (N_633,In_198,In_12);
or U634 (N_634,In_588,In_494);
nor U635 (N_635,In_89,In_626);
nand U636 (N_636,In_397,In_726);
nor U637 (N_637,In_382,In_224);
and U638 (N_638,In_257,In_179);
or U639 (N_639,In_24,In_221);
nand U640 (N_640,In_18,In_568);
nor U641 (N_641,In_55,In_195);
nand U642 (N_642,In_26,In_10);
nand U643 (N_643,In_529,In_329);
nor U644 (N_644,In_98,In_488);
nand U645 (N_645,In_174,In_584);
nand U646 (N_646,In_14,In_293);
nor U647 (N_647,In_336,In_227);
nor U648 (N_648,In_474,In_516);
nand U649 (N_649,In_258,In_308);
nand U650 (N_650,In_488,In_552);
nand U651 (N_651,In_436,In_278);
nor U652 (N_652,In_237,In_682);
nor U653 (N_653,In_349,In_609);
nand U654 (N_654,In_409,In_427);
and U655 (N_655,In_315,In_226);
or U656 (N_656,In_153,In_296);
nor U657 (N_657,In_82,In_208);
nor U658 (N_658,In_619,In_43);
and U659 (N_659,In_598,In_21);
and U660 (N_660,In_705,In_198);
or U661 (N_661,In_296,In_390);
or U662 (N_662,In_437,In_744);
nor U663 (N_663,In_247,In_341);
and U664 (N_664,In_593,In_122);
nor U665 (N_665,In_270,In_326);
nand U666 (N_666,In_596,In_228);
and U667 (N_667,In_642,In_568);
nand U668 (N_668,In_215,In_257);
nor U669 (N_669,In_182,In_130);
nand U670 (N_670,In_741,In_234);
nor U671 (N_671,In_156,In_356);
nor U672 (N_672,In_361,In_233);
nor U673 (N_673,In_381,In_245);
nand U674 (N_674,In_135,In_644);
nor U675 (N_675,In_321,In_118);
nor U676 (N_676,In_519,In_397);
nor U677 (N_677,In_514,In_331);
or U678 (N_678,In_399,In_213);
nand U679 (N_679,In_75,In_712);
or U680 (N_680,In_321,In_90);
xnor U681 (N_681,In_345,In_674);
and U682 (N_682,In_572,In_7);
nor U683 (N_683,In_626,In_150);
or U684 (N_684,In_7,In_231);
nor U685 (N_685,In_420,In_472);
and U686 (N_686,In_447,In_172);
or U687 (N_687,In_691,In_76);
or U688 (N_688,In_423,In_476);
or U689 (N_689,In_676,In_680);
nand U690 (N_690,In_736,In_150);
nand U691 (N_691,In_296,In_364);
and U692 (N_692,In_403,In_545);
nor U693 (N_693,In_485,In_252);
or U694 (N_694,In_185,In_501);
and U695 (N_695,In_500,In_660);
nand U696 (N_696,In_286,In_145);
nand U697 (N_697,In_140,In_573);
and U698 (N_698,In_425,In_631);
and U699 (N_699,In_356,In_340);
nand U700 (N_700,In_559,In_434);
or U701 (N_701,In_131,In_565);
nand U702 (N_702,In_248,In_80);
and U703 (N_703,In_548,In_512);
nand U704 (N_704,In_389,In_51);
nand U705 (N_705,In_460,In_509);
nor U706 (N_706,In_231,In_736);
nor U707 (N_707,In_103,In_515);
nand U708 (N_708,In_689,In_195);
or U709 (N_709,In_208,In_423);
or U710 (N_710,In_180,In_183);
nand U711 (N_711,In_688,In_684);
nor U712 (N_712,In_621,In_418);
nand U713 (N_713,In_733,In_703);
nor U714 (N_714,In_543,In_512);
nand U715 (N_715,In_412,In_330);
nor U716 (N_716,In_169,In_41);
or U717 (N_717,In_320,In_210);
or U718 (N_718,In_500,In_259);
and U719 (N_719,In_146,In_225);
or U720 (N_720,In_30,In_6);
or U721 (N_721,In_12,In_495);
or U722 (N_722,In_259,In_398);
and U723 (N_723,In_736,In_740);
nand U724 (N_724,In_730,In_680);
or U725 (N_725,In_736,In_402);
nor U726 (N_726,In_527,In_468);
or U727 (N_727,In_510,In_629);
nor U728 (N_728,In_720,In_644);
and U729 (N_729,In_536,In_398);
or U730 (N_730,In_186,In_547);
nand U731 (N_731,In_627,In_133);
or U732 (N_732,In_744,In_440);
and U733 (N_733,In_401,In_110);
and U734 (N_734,In_673,In_197);
or U735 (N_735,In_146,In_642);
nand U736 (N_736,In_648,In_509);
nand U737 (N_737,In_585,In_663);
nand U738 (N_738,In_411,In_641);
or U739 (N_739,In_736,In_486);
and U740 (N_740,In_481,In_191);
and U741 (N_741,In_531,In_487);
nand U742 (N_742,In_429,In_32);
and U743 (N_743,In_298,In_217);
nor U744 (N_744,In_413,In_206);
or U745 (N_745,In_619,In_667);
nand U746 (N_746,In_523,In_8);
nor U747 (N_747,In_270,In_204);
nor U748 (N_748,In_96,In_620);
and U749 (N_749,In_464,In_22);
and U750 (N_750,In_264,In_158);
nand U751 (N_751,In_284,In_608);
nand U752 (N_752,In_221,In_582);
and U753 (N_753,In_142,In_502);
nand U754 (N_754,In_280,In_626);
or U755 (N_755,In_718,In_184);
or U756 (N_756,In_8,In_215);
nand U757 (N_757,In_327,In_257);
and U758 (N_758,In_243,In_588);
and U759 (N_759,In_507,In_720);
and U760 (N_760,In_524,In_37);
or U761 (N_761,In_407,In_524);
nand U762 (N_762,In_3,In_670);
nor U763 (N_763,In_38,In_594);
and U764 (N_764,In_251,In_328);
or U765 (N_765,In_113,In_20);
or U766 (N_766,In_392,In_82);
nor U767 (N_767,In_575,In_405);
nor U768 (N_768,In_420,In_466);
nand U769 (N_769,In_205,In_408);
and U770 (N_770,In_93,In_292);
and U771 (N_771,In_745,In_435);
nand U772 (N_772,In_327,In_266);
or U773 (N_773,In_222,In_32);
or U774 (N_774,In_723,In_99);
nor U775 (N_775,In_529,In_473);
and U776 (N_776,In_115,In_166);
nor U777 (N_777,In_261,In_604);
nor U778 (N_778,In_543,In_39);
nor U779 (N_779,In_575,In_10);
or U780 (N_780,In_63,In_214);
nor U781 (N_781,In_505,In_417);
and U782 (N_782,In_201,In_223);
nor U783 (N_783,In_172,In_304);
or U784 (N_784,In_564,In_729);
nor U785 (N_785,In_232,In_74);
and U786 (N_786,In_573,In_316);
or U787 (N_787,In_255,In_16);
or U788 (N_788,In_269,In_30);
and U789 (N_789,In_263,In_157);
and U790 (N_790,In_21,In_66);
nand U791 (N_791,In_644,In_147);
or U792 (N_792,In_398,In_293);
nand U793 (N_793,In_668,In_551);
or U794 (N_794,In_519,In_337);
nor U795 (N_795,In_490,In_349);
or U796 (N_796,In_53,In_120);
nor U797 (N_797,In_644,In_29);
and U798 (N_798,In_269,In_207);
nand U799 (N_799,In_225,In_76);
nor U800 (N_800,In_483,In_699);
nor U801 (N_801,In_56,In_667);
or U802 (N_802,In_703,In_334);
nor U803 (N_803,In_18,In_364);
and U804 (N_804,In_442,In_552);
nand U805 (N_805,In_187,In_701);
or U806 (N_806,In_119,In_165);
nand U807 (N_807,In_363,In_594);
nand U808 (N_808,In_646,In_359);
and U809 (N_809,In_137,In_652);
or U810 (N_810,In_214,In_479);
nor U811 (N_811,In_684,In_674);
nor U812 (N_812,In_220,In_309);
nor U813 (N_813,In_497,In_663);
and U814 (N_814,In_203,In_218);
or U815 (N_815,In_467,In_515);
nand U816 (N_816,In_36,In_21);
or U817 (N_817,In_384,In_341);
nor U818 (N_818,In_387,In_108);
and U819 (N_819,In_574,In_327);
or U820 (N_820,In_439,In_33);
or U821 (N_821,In_308,In_126);
nand U822 (N_822,In_508,In_66);
and U823 (N_823,In_65,In_15);
xnor U824 (N_824,In_741,In_586);
nor U825 (N_825,In_364,In_450);
nand U826 (N_826,In_571,In_78);
or U827 (N_827,In_672,In_621);
or U828 (N_828,In_453,In_707);
or U829 (N_829,In_612,In_351);
and U830 (N_830,In_409,In_235);
nor U831 (N_831,In_477,In_309);
nand U832 (N_832,In_549,In_392);
or U833 (N_833,In_270,In_56);
and U834 (N_834,In_704,In_420);
nand U835 (N_835,In_132,In_483);
nor U836 (N_836,In_414,In_375);
or U837 (N_837,In_121,In_701);
nand U838 (N_838,In_9,In_483);
and U839 (N_839,In_210,In_278);
or U840 (N_840,In_274,In_503);
nand U841 (N_841,In_672,In_102);
nand U842 (N_842,In_424,In_94);
or U843 (N_843,In_374,In_153);
nor U844 (N_844,In_647,In_141);
or U845 (N_845,In_551,In_133);
nand U846 (N_846,In_72,In_94);
nand U847 (N_847,In_152,In_266);
nand U848 (N_848,In_277,In_181);
nand U849 (N_849,In_528,In_737);
and U850 (N_850,In_438,In_382);
nor U851 (N_851,In_330,In_132);
nor U852 (N_852,In_480,In_444);
nor U853 (N_853,In_360,In_226);
nand U854 (N_854,In_238,In_447);
nand U855 (N_855,In_727,In_86);
nor U856 (N_856,In_572,In_69);
nand U857 (N_857,In_256,In_152);
or U858 (N_858,In_677,In_414);
nand U859 (N_859,In_417,In_603);
or U860 (N_860,In_364,In_680);
nand U861 (N_861,In_187,In_411);
nor U862 (N_862,In_447,In_635);
nor U863 (N_863,In_462,In_143);
or U864 (N_864,In_152,In_697);
and U865 (N_865,In_290,In_117);
nor U866 (N_866,In_535,In_511);
nor U867 (N_867,In_636,In_541);
and U868 (N_868,In_103,In_522);
and U869 (N_869,In_156,In_417);
nand U870 (N_870,In_107,In_324);
nor U871 (N_871,In_538,In_436);
nor U872 (N_872,In_550,In_661);
or U873 (N_873,In_549,In_40);
or U874 (N_874,In_733,In_212);
or U875 (N_875,In_133,In_96);
nor U876 (N_876,In_85,In_48);
and U877 (N_877,In_720,In_105);
or U878 (N_878,In_434,In_68);
nand U879 (N_879,In_36,In_512);
nand U880 (N_880,In_495,In_155);
nand U881 (N_881,In_620,In_329);
nor U882 (N_882,In_403,In_118);
nor U883 (N_883,In_451,In_424);
or U884 (N_884,In_100,In_447);
and U885 (N_885,In_8,In_373);
and U886 (N_886,In_13,In_38);
nand U887 (N_887,In_149,In_209);
nor U888 (N_888,In_254,In_435);
nand U889 (N_889,In_244,In_605);
or U890 (N_890,In_749,In_534);
nand U891 (N_891,In_116,In_624);
and U892 (N_892,In_105,In_498);
nand U893 (N_893,In_453,In_17);
or U894 (N_894,In_342,In_657);
or U895 (N_895,In_679,In_738);
nand U896 (N_896,In_317,In_573);
or U897 (N_897,In_116,In_136);
or U898 (N_898,In_149,In_132);
and U899 (N_899,In_624,In_577);
nand U900 (N_900,In_324,In_459);
and U901 (N_901,In_537,In_409);
or U902 (N_902,In_224,In_115);
or U903 (N_903,In_27,In_242);
nor U904 (N_904,In_739,In_404);
nand U905 (N_905,In_748,In_640);
nand U906 (N_906,In_593,In_20);
and U907 (N_907,In_112,In_401);
nand U908 (N_908,In_153,In_284);
and U909 (N_909,In_14,In_539);
nor U910 (N_910,In_253,In_278);
nor U911 (N_911,In_457,In_445);
or U912 (N_912,In_190,In_26);
or U913 (N_913,In_371,In_84);
nand U914 (N_914,In_600,In_152);
xnor U915 (N_915,In_323,In_321);
and U916 (N_916,In_304,In_9);
nor U917 (N_917,In_470,In_381);
or U918 (N_918,In_196,In_719);
nand U919 (N_919,In_512,In_28);
nor U920 (N_920,In_243,In_197);
xnor U921 (N_921,In_236,In_431);
and U922 (N_922,In_547,In_598);
nor U923 (N_923,In_317,In_18);
nor U924 (N_924,In_328,In_649);
nor U925 (N_925,In_204,In_679);
nor U926 (N_926,In_185,In_447);
or U927 (N_927,In_674,In_653);
or U928 (N_928,In_714,In_353);
and U929 (N_929,In_581,In_132);
nand U930 (N_930,In_140,In_221);
and U931 (N_931,In_4,In_557);
and U932 (N_932,In_242,In_572);
or U933 (N_933,In_612,In_477);
and U934 (N_934,In_13,In_367);
or U935 (N_935,In_745,In_658);
or U936 (N_936,In_151,In_597);
or U937 (N_937,In_448,In_251);
and U938 (N_938,In_553,In_607);
nor U939 (N_939,In_590,In_207);
nand U940 (N_940,In_376,In_576);
nor U941 (N_941,In_390,In_442);
or U942 (N_942,In_466,In_667);
or U943 (N_943,In_496,In_382);
nor U944 (N_944,In_514,In_628);
and U945 (N_945,In_420,In_213);
nor U946 (N_946,In_55,In_294);
or U947 (N_947,In_543,In_367);
or U948 (N_948,In_265,In_277);
and U949 (N_949,In_343,In_244);
nor U950 (N_950,In_447,In_174);
nand U951 (N_951,In_106,In_28);
nand U952 (N_952,In_303,In_368);
or U953 (N_953,In_27,In_320);
or U954 (N_954,In_668,In_20);
and U955 (N_955,In_644,In_564);
nor U956 (N_956,In_307,In_289);
or U957 (N_957,In_325,In_339);
or U958 (N_958,In_22,In_614);
and U959 (N_959,In_579,In_108);
nand U960 (N_960,In_581,In_507);
nand U961 (N_961,In_218,In_682);
nor U962 (N_962,In_630,In_523);
or U963 (N_963,In_600,In_12);
and U964 (N_964,In_578,In_430);
nor U965 (N_965,In_110,In_368);
or U966 (N_966,In_196,In_262);
nand U967 (N_967,In_629,In_291);
and U968 (N_968,In_732,In_689);
nand U969 (N_969,In_469,In_699);
nor U970 (N_970,In_384,In_583);
or U971 (N_971,In_21,In_244);
or U972 (N_972,In_631,In_302);
or U973 (N_973,In_527,In_582);
and U974 (N_974,In_567,In_731);
nand U975 (N_975,In_610,In_32);
nand U976 (N_976,In_513,In_376);
and U977 (N_977,In_638,In_554);
and U978 (N_978,In_582,In_588);
and U979 (N_979,In_467,In_634);
nand U980 (N_980,In_662,In_271);
nand U981 (N_981,In_401,In_545);
nand U982 (N_982,In_424,In_65);
nor U983 (N_983,In_75,In_275);
or U984 (N_984,In_162,In_594);
or U985 (N_985,In_323,In_413);
or U986 (N_986,In_341,In_245);
nand U987 (N_987,In_731,In_664);
or U988 (N_988,In_62,In_338);
and U989 (N_989,In_310,In_668);
nor U990 (N_990,In_348,In_608);
or U991 (N_991,In_605,In_319);
nor U992 (N_992,In_465,In_308);
and U993 (N_993,In_22,In_239);
nand U994 (N_994,In_103,In_350);
nand U995 (N_995,In_653,In_143);
or U996 (N_996,In_556,In_614);
nor U997 (N_997,In_322,In_568);
nor U998 (N_998,In_14,In_657);
nand U999 (N_999,In_382,In_39);
or U1000 (N_1000,In_287,In_397);
nand U1001 (N_1001,In_661,In_334);
or U1002 (N_1002,In_457,In_177);
or U1003 (N_1003,In_466,In_403);
and U1004 (N_1004,In_199,In_280);
xor U1005 (N_1005,In_601,In_385);
or U1006 (N_1006,In_196,In_0);
nor U1007 (N_1007,In_135,In_22);
nor U1008 (N_1008,In_303,In_105);
or U1009 (N_1009,In_214,In_304);
or U1010 (N_1010,In_379,In_588);
or U1011 (N_1011,In_397,In_257);
and U1012 (N_1012,In_124,In_732);
or U1013 (N_1013,In_609,In_368);
and U1014 (N_1014,In_249,In_241);
nand U1015 (N_1015,In_340,In_209);
or U1016 (N_1016,In_568,In_165);
or U1017 (N_1017,In_702,In_216);
nand U1018 (N_1018,In_284,In_573);
and U1019 (N_1019,In_740,In_335);
or U1020 (N_1020,In_286,In_651);
or U1021 (N_1021,In_295,In_243);
and U1022 (N_1022,In_194,In_136);
or U1023 (N_1023,In_370,In_691);
nor U1024 (N_1024,In_48,In_380);
and U1025 (N_1025,In_221,In_666);
and U1026 (N_1026,In_457,In_583);
nand U1027 (N_1027,In_290,In_113);
or U1028 (N_1028,In_419,In_132);
nand U1029 (N_1029,In_681,In_486);
or U1030 (N_1030,In_423,In_412);
and U1031 (N_1031,In_75,In_362);
and U1032 (N_1032,In_326,In_501);
and U1033 (N_1033,In_356,In_514);
nor U1034 (N_1034,In_437,In_39);
or U1035 (N_1035,In_654,In_34);
or U1036 (N_1036,In_76,In_325);
or U1037 (N_1037,In_609,In_445);
nand U1038 (N_1038,In_509,In_722);
nor U1039 (N_1039,In_141,In_225);
and U1040 (N_1040,In_244,In_383);
or U1041 (N_1041,In_376,In_296);
and U1042 (N_1042,In_125,In_151);
nand U1043 (N_1043,In_370,In_716);
nand U1044 (N_1044,In_601,In_541);
and U1045 (N_1045,In_292,In_119);
nor U1046 (N_1046,In_426,In_9);
and U1047 (N_1047,In_699,In_495);
nor U1048 (N_1048,In_219,In_366);
nand U1049 (N_1049,In_97,In_105);
and U1050 (N_1050,In_146,In_706);
nor U1051 (N_1051,In_260,In_739);
nor U1052 (N_1052,In_574,In_103);
and U1053 (N_1053,In_307,In_153);
or U1054 (N_1054,In_696,In_419);
nor U1055 (N_1055,In_511,In_715);
nand U1056 (N_1056,In_51,In_63);
or U1057 (N_1057,In_392,In_681);
and U1058 (N_1058,In_369,In_270);
nor U1059 (N_1059,In_472,In_640);
nand U1060 (N_1060,In_92,In_42);
nor U1061 (N_1061,In_507,In_444);
or U1062 (N_1062,In_88,In_258);
or U1063 (N_1063,In_118,In_702);
or U1064 (N_1064,In_190,In_304);
or U1065 (N_1065,In_6,In_257);
nor U1066 (N_1066,In_454,In_638);
or U1067 (N_1067,In_472,In_70);
nor U1068 (N_1068,In_226,In_123);
or U1069 (N_1069,In_731,In_572);
or U1070 (N_1070,In_435,In_449);
and U1071 (N_1071,In_717,In_148);
nand U1072 (N_1072,In_299,In_363);
nor U1073 (N_1073,In_476,In_505);
and U1074 (N_1074,In_539,In_688);
nand U1075 (N_1075,In_226,In_727);
or U1076 (N_1076,In_564,In_731);
and U1077 (N_1077,In_724,In_55);
nand U1078 (N_1078,In_570,In_607);
and U1079 (N_1079,In_209,In_116);
or U1080 (N_1080,In_664,In_410);
or U1081 (N_1081,In_347,In_542);
nand U1082 (N_1082,In_403,In_620);
nor U1083 (N_1083,In_251,In_77);
nor U1084 (N_1084,In_401,In_179);
nand U1085 (N_1085,In_227,In_260);
and U1086 (N_1086,In_273,In_226);
or U1087 (N_1087,In_335,In_737);
nand U1088 (N_1088,In_423,In_444);
nor U1089 (N_1089,In_370,In_565);
and U1090 (N_1090,In_522,In_30);
nand U1091 (N_1091,In_161,In_166);
or U1092 (N_1092,In_634,In_604);
nand U1093 (N_1093,In_675,In_149);
nand U1094 (N_1094,In_231,In_212);
or U1095 (N_1095,In_217,In_593);
nor U1096 (N_1096,In_500,In_47);
xor U1097 (N_1097,In_586,In_738);
and U1098 (N_1098,In_707,In_141);
nor U1099 (N_1099,In_189,In_272);
or U1100 (N_1100,In_599,In_472);
xnor U1101 (N_1101,In_164,In_533);
nor U1102 (N_1102,In_681,In_398);
or U1103 (N_1103,In_274,In_79);
nor U1104 (N_1104,In_281,In_312);
and U1105 (N_1105,In_699,In_34);
or U1106 (N_1106,In_189,In_145);
or U1107 (N_1107,In_281,In_387);
nand U1108 (N_1108,In_292,In_453);
or U1109 (N_1109,In_69,In_711);
nand U1110 (N_1110,In_610,In_650);
nor U1111 (N_1111,In_603,In_676);
nand U1112 (N_1112,In_225,In_99);
and U1113 (N_1113,In_359,In_387);
nand U1114 (N_1114,In_45,In_42);
and U1115 (N_1115,In_352,In_170);
and U1116 (N_1116,In_665,In_454);
nor U1117 (N_1117,In_241,In_33);
nand U1118 (N_1118,In_420,In_72);
or U1119 (N_1119,In_633,In_440);
nor U1120 (N_1120,In_699,In_493);
nor U1121 (N_1121,In_553,In_20);
nor U1122 (N_1122,In_251,In_432);
or U1123 (N_1123,In_102,In_244);
nand U1124 (N_1124,In_596,In_460);
nand U1125 (N_1125,In_689,In_481);
nand U1126 (N_1126,In_734,In_257);
or U1127 (N_1127,In_230,In_92);
nand U1128 (N_1128,In_467,In_571);
or U1129 (N_1129,In_71,In_555);
or U1130 (N_1130,In_525,In_537);
nand U1131 (N_1131,In_329,In_515);
nor U1132 (N_1132,In_318,In_694);
and U1133 (N_1133,In_461,In_214);
xor U1134 (N_1134,In_41,In_129);
nand U1135 (N_1135,In_112,In_388);
nor U1136 (N_1136,In_259,In_229);
nor U1137 (N_1137,In_283,In_535);
or U1138 (N_1138,In_200,In_524);
nand U1139 (N_1139,In_258,In_595);
and U1140 (N_1140,In_391,In_214);
xnor U1141 (N_1141,In_597,In_269);
nand U1142 (N_1142,In_717,In_557);
nor U1143 (N_1143,In_160,In_617);
and U1144 (N_1144,In_277,In_647);
nand U1145 (N_1145,In_618,In_214);
or U1146 (N_1146,In_654,In_359);
and U1147 (N_1147,In_89,In_239);
nand U1148 (N_1148,In_162,In_178);
nor U1149 (N_1149,In_357,In_392);
or U1150 (N_1150,In_605,In_533);
nand U1151 (N_1151,In_237,In_463);
nor U1152 (N_1152,In_716,In_590);
nand U1153 (N_1153,In_240,In_227);
and U1154 (N_1154,In_275,In_623);
nand U1155 (N_1155,In_136,In_115);
and U1156 (N_1156,In_203,In_619);
or U1157 (N_1157,In_95,In_300);
or U1158 (N_1158,In_507,In_579);
and U1159 (N_1159,In_746,In_260);
nand U1160 (N_1160,In_437,In_218);
nor U1161 (N_1161,In_526,In_233);
nand U1162 (N_1162,In_41,In_520);
and U1163 (N_1163,In_341,In_523);
and U1164 (N_1164,In_276,In_555);
nor U1165 (N_1165,In_2,In_83);
xnor U1166 (N_1166,In_527,In_706);
nand U1167 (N_1167,In_115,In_88);
or U1168 (N_1168,In_473,In_372);
and U1169 (N_1169,In_390,In_319);
nor U1170 (N_1170,In_160,In_155);
nand U1171 (N_1171,In_369,In_610);
nand U1172 (N_1172,In_317,In_207);
or U1173 (N_1173,In_299,In_450);
nand U1174 (N_1174,In_138,In_632);
and U1175 (N_1175,In_243,In_177);
or U1176 (N_1176,In_342,In_721);
nand U1177 (N_1177,In_682,In_612);
nand U1178 (N_1178,In_64,In_100);
or U1179 (N_1179,In_260,In_11);
nand U1180 (N_1180,In_29,In_561);
and U1181 (N_1181,In_271,In_671);
nand U1182 (N_1182,In_588,In_523);
nor U1183 (N_1183,In_89,In_330);
or U1184 (N_1184,In_612,In_566);
or U1185 (N_1185,In_418,In_599);
and U1186 (N_1186,In_435,In_11);
or U1187 (N_1187,In_33,In_122);
or U1188 (N_1188,In_117,In_557);
and U1189 (N_1189,In_227,In_14);
nor U1190 (N_1190,In_314,In_338);
or U1191 (N_1191,In_344,In_139);
or U1192 (N_1192,In_19,In_455);
or U1193 (N_1193,In_67,In_618);
nor U1194 (N_1194,In_532,In_525);
nand U1195 (N_1195,In_432,In_635);
nor U1196 (N_1196,In_340,In_673);
or U1197 (N_1197,In_7,In_488);
nor U1198 (N_1198,In_125,In_594);
nand U1199 (N_1199,In_590,In_33);
and U1200 (N_1200,In_346,In_153);
and U1201 (N_1201,In_291,In_572);
and U1202 (N_1202,In_557,In_408);
nand U1203 (N_1203,In_105,In_55);
or U1204 (N_1204,In_334,In_339);
nand U1205 (N_1205,In_546,In_543);
and U1206 (N_1206,In_114,In_485);
nor U1207 (N_1207,In_542,In_273);
and U1208 (N_1208,In_693,In_13);
and U1209 (N_1209,In_309,In_676);
and U1210 (N_1210,In_228,In_117);
nand U1211 (N_1211,In_670,In_690);
or U1212 (N_1212,In_231,In_209);
and U1213 (N_1213,In_27,In_715);
and U1214 (N_1214,In_699,In_693);
nand U1215 (N_1215,In_738,In_685);
nor U1216 (N_1216,In_354,In_161);
nand U1217 (N_1217,In_580,In_368);
and U1218 (N_1218,In_536,In_541);
and U1219 (N_1219,In_41,In_513);
nor U1220 (N_1220,In_387,In_552);
and U1221 (N_1221,In_700,In_517);
or U1222 (N_1222,In_349,In_544);
or U1223 (N_1223,In_665,In_110);
nand U1224 (N_1224,In_101,In_566);
nor U1225 (N_1225,In_384,In_532);
nand U1226 (N_1226,In_576,In_580);
or U1227 (N_1227,In_137,In_279);
and U1228 (N_1228,In_661,In_200);
and U1229 (N_1229,In_371,In_421);
nor U1230 (N_1230,In_481,In_295);
or U1231 (N_1231,In_265,In_488);
nor U1232 (N_1232,In_47,In_66);
or U1233 (N_1233,In_106,In_335);
nor U1234 (N_1234,In_104,In_158);
or U1235 (N_1235,In_383,In_28);
nor U1236 (N_1236,In_482,In_172);
or U1237 (N_1237,In_451,In_348);
or U1238 (N_1238,In_714,In_265);
or U1239 (N_1239,In_92,In_658);
nand U1240 (N_1240,In_144,In_95);
or U1241 (N_1241,In_337,In_248);
nor U1242 (N_1242,In_606,In_85);
nand U1243 (N_1243,In_37,In_600);
nand U1244 (N_1244,In_659,In_67);
nor U1245 (N_1245,In_52,In_675);
nor U1246 (N_1246,In_533,In_244);
or U1247 (N_1247,In_730,In_572);
nor U1248 (N_1248,In_106,In_162);
or U1249 (N_1249,In_94,In_451);
nor U1250 (N_1250,In_204,In_163);
xor U1251 (N_1251,In_380,In_247);
nand U1252 (N_1252,In_264,In_262);
nor U1253 (N_1253,In_125,In_598);
nand U1254 (N_1254,In_177,In_29);
nor U1255 (N_1255,In_470,In_63);
and U1256 (N_1256,In_195,In_408);
nand U1257 (N_1257,In_568,In_362);
nor U1258 (N_1258,In_324,In_662);
nor U1259 (N_1259,In_533,In_590);
or U1260 (N_1260,In_295,In_484);
or U1261 (N_1261,In_600,In_203);
nand U1262 (N_1262,In_333,In_349);
nor U1263 (N_1263,In_157,In_136);
nand U1264 (N_1264,In_144,In_427);
xor U1265 (N_1265,In_77,In_107);
or U1266 (N_1266,In_538,In_48);
and U1267 (N_1267,In_127,In_610);
and U1268 (N_1268,In_647,In_375);
and U1269 (N_1269,In_129,In_281);
and U1270 (N_1270,In_243,In_267);
and U1271 (N_1271,In_251,In_173);
or U1272 (N_1272,In_563,In_36);
nor U1273 (N_1273,In_526,In_701);
or U1274 (N_1274,In_17,In_581);
nand U1275 (N_1275,In_638,In_483);
nand U1276 (N_1276,In_522,In_641);
nand U1277 (N_1277,In_590,In_307);
and U1278 (N_1278,In_104,In_318);
nor U1279 (N_1279,In_396,In_127);
and U1280 (N_1280,In_439,In_132);
nor U1281 (N_1281,In_369,In_320);
and U1282 (N_1282,In_453,In_250);
nand U1283 (N_1283,In_234,In_585);
nor U1284 (N_1284,In_47,In_566);
nand U1285 (N_1285,In_18,In_149);
nor U1286 (N_1286,In_337,In_263);
nor U1287 (N_1287,In_67,In_179);
nor U1288 (N_1288,In_30,In_618);
and U1289 (N_1289,In_114,In_443);
and U1290 (N_1290,In_506,In_651);
nand U1291 (N_1291,In_330,In_605);
nor U1292 (N_1292,In_748,In_367);
nand U1293 (N_1293,In_204,In_713);
or U1294 (N_1294,In_662,In_694);
nor U1295 (N_1295,In_190,In_711);
nand U1296 (N_1296,In_145,In_203);
or U1297 (N_1297,In_59,In_475);
nor U1298 (N_1298,In_582,In_3);
or U1299 (N_1299,In_379,In_70);
and U1300 (N_1300,In_391,In_279);
nand U1301 (N_1301,In_708,In_362);
and U1302 (N_1302,In_289,In_271);
nor U1303 (N_1303,In_341,In_575);
nand U1304 (N_1304,In_262,In_464);
and U1305 (N_1305,In_359,In_139);
or U1306 (N_1306,In_643,In_374);
nand U1307 (N_1307,In_195,In_499);
nor U1308 (N_1308,In_229,In_705);
or U1309 (N_1309,In_487,In_72);
or U1310 (N_1310,In_83,In_734);
or U1311 (N_1311,In_437,In_237);
or U1312 (N_1312,In_549,In_695);
nor U1313 (N_1313,In_655,In_467);
or U1314 (N_1314,In_549,In_742);
nor U1315 (N_1315,In_119,In_54);
or U1316 (N_1316,In_633,In_716);
and U1317 (N_1317,In_475,In_732);
or U1318 (N_1318,In_661,In_462);
and U1319 (N_1319,In_282,In_673);
nand U1320 (N_1320,In_538,In_453);
nor U1321 (N_1321,In_32,In_299);
and U1322 (N_1322,In_348,In_291);
and U1323 (N_1323,In_29,In_34);
and U1324 (N_1324,In_319,In_701);
and U1325 (N_1325,In_7,In_506);
and U1326 (N_1326,In_415,In_704);
and U1327 (N_1327,In_694,In_327);
or U1328 (N_1328,In_734,In_89);
nor U1329 (N_1329,In_216,In_167);
nand U1330 (N_1330,In_634,In_446);
nand U1331 (N_1331,In_590,In_542);
and U1332 (N_1332,In_728,In_732);
nand U1333 (N_1333,In_589,In_727);
and U1334 (N_1334,In_74,In_363);
nor U1335 (N_1335,In_609,In_322);
and U1336 (N_1336,In_5,In_225);
xnor U1337 (N_1337,In_614,In_587);
nand U1338 (N_1338,In_616,In_219);
nor U1339 (N_1339,In_121,In_583);
nor U1340 (N_1340,In_749,In_516);
nand U1341 (N_1341,In_235,In_419);
or U1342 (N_1342,In_57,In_726);
nand U1343 (N_1343,In_220,In_240);
and U1344 (N_1344,In_341,In_137);
nor U1345 (N_1345,In_524,In_262);
and U1346 (N_1346,In_641,In_584);
nor U1347 (N_1347,In_155,In_168);
nor U1348 (N_1348,In_4,In_564);
nand U1349 (N_1349,In_15,In_726);
nor U1350 (N_1350,In_741,In_623);
nor U1351 (N_1351,In_110,In_501);
or U1352 (N_1352,In_150,In_428);
nand U1353 (N_1353,In_713,In_521);
nor U1354 (N_1354,In_558,In_390);
nand U1355 (N_1355,In_72,In_27);
nand U1356 (N_1356,In_511,In_672);
and U1357 (N_1357,In_472,In_154);
and U1358 (N_1358,In_661,In_87);
and U1359 (N_1359,In_470,In_706);
nand U1360 (N_1360,In_248,In_334);
nor U1361 (N_1361,In_607,In_560);
nor U1362 (N_1362,In_123,In_614);
nor U1363 (N_1363,In_398,In_128);
and U1364 (N_1364,In_470,In_473);
or U1365 (N_1365,In_502,In_150);
nor U1366 (N_1366,In_535,In_22);
nor U1367 (N_1367,In_351,In_621);
nor U1368 (N_1368,In_702,In_527);
nor U1369 (N_1369,In_686,In_67);
nor U1370 (N_1370,In_419,In_130);
or U1371 (N_1371,In_647,In_103);
or U1372 (N_1372,In_726,In_293);
nand U1373 (N_1373,In_283,In_134);
nor U1374 (N_1374,In_567,In_530);
or U1375 (N_1375,In_194,In_527);
nand U1376 (N_1376,In_652,In_585);
nand U1377 (N_1377,In_625,In_130);
or U1378 (N_1378,In_227,In_522);
nor U1379 (N_1379,In_734,In_66);
nand U1380 (N_1380,In_570,In_80);
or U1381 (N_1381,In_141,In_331);
or U1382 (N_1382,In_362,In_177);
nand U1383 (N_1383,In_639,In_686);
or U1384 (N_1384,In_594,In_698);
and U1385 (N_1385,In_562,In_49);
nand U1386 (N_1386,In_451,In_657);
and U1387 (N_1387,In_560,In_285);
or U1388 (N_1388,In_283,In_521);
or U1389 (N_1389,In_333,In_578);
and U1390 (N_1390,In_408,In_196);
nor U1391 (N_1391,In_729,In_474);
or U1392 (N_1392,In_478,In_521);
nor U1393 (N_1393,In_600,In_742);
nor U1394 (N_1394,In_330,In_589);
or U1395 (N_1395,In_548,In_486);
nor U1396 (N_1396,In_613,In_122);
nand U1397 (N_1397,In_307,In_166);
nor U1398 (N_1398,In_345,In_316);
nor U1399 (N_1399,In_268,In_613);
nor U1400 (N_1400,In_635,In_220);
nand U1401 (N_1401,In_404,In_292);
nand U1402 (N_1402,In_59,In_429);
or U1403 (N_1403,In_353,In_219);
or U1404 (N_1404,In_248,In_54);
nand U1405 (N_1405,In_723,In_304);
or U1406 (N_1406,In_51,In_646);
and U1407 (N_1407,In_107,In_125);
nor U1408 (N_1408,In_648,In_577);
and U1409 (N_1409,In_239,In_491);
nand U1410 (N_1410,In_562,In_378);
nand U1411 (N_1411,In_377,In_572);
or U1412 (N_1412,In_689,In_252);
and U1413 (N_1413,In_652,In_445);
nand U1414 (N_1414,In_123,In_749);
nor U1415 (N_1415,In_308,In_19);
and U1416 (N_1416,In_361,In_29);
nor U1417 (N_1417,In_706,In_44);
and U1418 (N_1418,In_367,In_503);
nor U1419 (N_1419,In_16,In_745);
or U1420 (N_1420,In_282,In_635);
or U1421 (N_1421,In_379,In_462);
nand U1422 (N_1422,In_416,In_328);
nand U1423 (N_1423,In_326,In_459);
or U1424 (N_1424,In_707,In_375);
nor U1425 (N_1425,In_699,In_344);
or U1426 (N_1426,In_165,In_590);
nand U1427 (N_1427,In_663,In_57);
and U1428 (N_1428,In_216,In_438);
and U1429 (N_1429,In_279,In_745);
nor U1430 (N_1430,In_328,In_584);
nor U1431 (N_1431,In_369,In_56);
and U1432 (N_1432,In_323,In_60);
and U1433 (N_1433,In_668,In_3);
or U1434 (N_1434,In_117,In_182);
nor U1435 (N_1435,In_120,In_102);
and U1436 (N_1436,In_375,In_372);
nor U1437 (N_1437,In_729,In_595);
nor U1438 (N_1438,In_536,In_269);
and U1439 (N_1439,In_490,In_669);
nor U1440 (N_1440,In_588,In_155);
or U1441 (N_1441,In_271,In_575);
nor U1442 (N_1442,In_89,In_142);
and U1443 (N_1443,In_468,In_371);
nand U1444 (N_1444,In_95,In_634);
nor U1445 (N_1445,In_710,In_453);
nand U1446 (N_1446,In_718,In_158);
and U1447 (N_1447,In_380,In_368);
or U1448 (N_1448,In_588,In_193);
and U1449 (N_1449,In_627,In_240);
or U1450 (N_1450,In_80,In_289);
or U1451 (N_1451,In_491,In_700);
and U1452 (N_1452,In_457,In_613);
nor U1453 (N_1453,In_364,In_559);
nand U1454 (N_1454,In_748,In_238);
or U1455 (N_1455,In_465,In_193);
or U1456 (N_1456,In_622,In_182);
or U1457 (N_1457,In_89,In_303);
and U1458 (N_1458,In_289,In_651);
and U1459 (N_1459,In_441,In_482);
nand U1460 (N_1460,In_534,In_705);
nor U1461 (N_1461,In_227,In_664);
and U1462 (N_1462,In_480,In_458);
nand U1463 (N_1463,In_579,In_229);
nor U1464 (N_1464,In_447,In_179);
nor U1465 (N_1465,In_450,In_437);
and U1466 (N_1466,In_540,In_305);
nand U1467 (N_1467,In_553,In_26);
nand U1468 (N_1468,In_240,In_321);
and U1469 (N_1469,In_29,In_630);
and U1470 (N_1470,In_396,In_260);
or U1471 (N_1471,In_511,In_68);
nand U1472 (N_1472,In_512,In_613);
nand U1473 (N_1473,In_87,In_269);
or U1474 (N_1474,In_436,In_83);
nor U1475 (N_1475,In_239,In_100);
or U1476 (N_1476,In_47,In_426);
nor U1477 (N_1477,In_310,In_44);
and U1478 (N_1478,In_175,In_671);
nand U1479 (N_1479,In_741,In_730);
nand U1480 (N_1480,In_253,In_72);
or U1481 (N_1481,In_339,In_379);
or U1482 (N_1482,In_293,In_94);
and U1483 (N_1483,In_429,In_572);
or U1484 (N_1484,In_458,In_730);
or U1485 (N_1485,In_594,In_637);
nor U1486 (N_1486,In_508,In_145);
or U1487 (N_1487,In_116,In_725);
nand U1488 (N_1488,In_253,In_619);
or U1489 (N_1489,In_270,In_186);
or U1490 (N_1490,In_452,In_302);
and U1491 (N_1491,In_713,In_433);
nand U1492 (N_1492,In_316,In_357);
nand U1493 (N_1493,In_505,In_59);
nand U1494 (N_1494,In_695,In_233);
nor U1495 (N_1495,In_739,In_490);
or U1496 (N_1496,In_721,In_644);
nand U1497 (N_1497,In_140,In_29);
or U1498 (N_1498,In_172,In_376);
nand U1499 (N_1499,In_35,In_143);
nand U1500 (N_1500,In_383,In_457);
or U1501 (N_1501,In_375,In_406);
nand U1502 (N_1502,In_648,In_682);
nor U1503 (N_1503,In_220,In_252);
or U1504 (N_1504,In_675,In_574);
nor U1505 (N_1505,In_101,In_392);
or U1506 (N_1506,In_464,In_503);
and U1507 (N_1507,In_494,In_649);
or U1508 (N_1508,In_497,In_540);
nand U1509 (N_1509,In_710,In_704);
nor U1510 (N_1510,In_59,In_62);
nor U1511 (N_1511,In_117,In_392);
nor U1512 (N_1512,In_29,In_192);
and U1513 (N_1513,In_102,In_78);
or U1514 (N_1514,In_124,In_399);
and U1515 (N_1515,In_378,In_574);
nand U1516 (N_1516,In_449,In_40);
or U1517 (N_1517,In_672,In_246);
or U1518 (N_1518,In_418,In_176);
nor U1519 (N_1519,In_305,In_227);
and U1520 (N_1520,In_658,In_21);
nand U1521 (N_1521,In_191,In_477);
xnor U1522 (N_1522,In_410,In_669);
and U1523 (N_1523,In_687,In_544);
or U1524 (N_1524,In_599,In_720);
or U1525 (N_1525,In_105,In_152);
or U1526 (N_1526,In_107,In_331);
nand U1527 (N_1527,In_438,In_430);
xnor U1528 (N_1528,In_534,In_380);
or U1529 (N_1529,In_677,In_148);
nand U1530 (N_1530,In_509,In_122);
and U1531 (N_1531,In_450,In_560);
nand U1532 (N_1532,In_392,In_244);
or U1533 (N_1533,In_672,In_209);
nor U1534 (N_1534,In_566,In_522);
or U1535 (N_1535,In_562,In_294);
and U1536 (N_1536,In_507,In_519);
nand U1537 (N_1537,In_744,In_66);
nand U1538 (N_1538,In_406,In_458);
nor U1539 (N_1539,In_458,In_223);
and U1540 (N_1540,In_301,In_421);
nand U1541 (N_1541,In_322,In_676);
and U1542 (N_1542,In_289,In_717);
nand U1543 (N_1543,In_129,In_383);
nand U1544 (N_1544,In_680,In_351);
or U1545 (N_1545,In_89,In_272);
or U1546 (N_1546,In_669,In_651);
or U1547 (N_1547,In_497,In_42);
nand U1548 (N_1548,In_731,In_293);
nand U1549 (N_1549,In_10,In_53);
nand U1550 (N_1550,In_294,In_222);
nor U1551 (N_1551,In_441,In_684);
nand U1552 (N_1552,In_664,In_439);
or U1553 (N_1553,In_521,In_731);
nor U1554 (N_1554,In_255,In_306);
or U1555 (N_1555,In_541,In_307);
nor U1556 (N_1556,In_616,In_239);
and U1557 (N_1557,In_690,In_187);
nand U1558 (N_1558,In_296,In_555);
and U1559 (N_1559,In_187,In_527);
nor U1560 (N_1560,In_437,In_461);
nor U1561 (N_1561,In_405,In_69);
and U1562 (N_1562,In_476,In_208);
nand U1563 (N_1563,In_325,In_291);
nand U1564 (N_1564,In_194,In_608);
nand U1565 (N_1565,In_704,In_208);
nand U1566 (N_1566,In_523,In_42);
nand U1567 (N_1567,In_409,In_429);
and U1568 (N_1568,In_555,In_2);
nor U1569 (N_1569,In_1,In_248);
or U1570 (N_1570,In_483,In_663);
or U1571 (N_1571,In_488,In_382);
nor U1572 (N_1572,In_695,In_507);
nor U1573 (N_1573,In_515,In_627);
and U1574 (N_1574,In_500,In_567);
nand U1575 (N_1575,In_182,In_364);
nor U1576 (N_1576,In_127,In_478);
nand U1577 (N_1577,In_316,In_83);
nor U1578 (N_1578,In_67,In_557);
nand U1579 (N_1579,In_482,In_560);
nand U1580 (N_1580,In_675,In_188);
nor U1581 (N_1581,In_275,In_130);
nand U1582 (N_1582,In_379,In_274);
or U1583 (N_1583,In_723,In_714);
nand U1584 (N_1584,In_314,In_426);
and U1585 (N_1585,In_122,In_322);
or U1586 (N_1586,In_601,In_338);
and U1587 (N_1587,In_522,In_636);
nand U1588 (N_1588,In_494,In_602);
nor U1589 (N_1589,In_214,In_747);
or U1590 (N_1590,In_387,In_617);
and U1591 (N_1591,In_162,In_376);
nand U1592 (N_1592,In_353,In_278);
nor U1593 (N_1593,In_575,In_635);
nand U1594 (N_1594,In_48,In_80);
nand U1595 (N_1595,In_481,In_138);
and U1596 (N_1596,In_82,In_738);
and U1597 (N_1597,In_158,In_65);
nand U1598 (N_1598,In_381,In_405);
and U1599 (N_1599,In_405,In_318);
xnor U1600 (N_1600,In_130,In_737);
or U1601 (N_1601,In_417,In_640);
nor U1602 (N_1602,In_725,In_359);
nand U1603 (N_1603,In_232,In_66);
nand U1604 (N_1604,In_617,In_20);
or U1605 (N_1605,In_170,In_86);
and U1606 (N_1606,In_590,In_425);
nand U1607 (N_1607,In_477,In_220);
or U1608 (N_1608,In_106,In_501);
xor U1609 (N_1609,In_550,In_440);
and U1610 (N_1610,In_214,In_580);
and U1611 (N_1611,In_391,In_476);
nor U1612 (N_1612,In_115,In_41);
nor U1613 (N_1613,In_481,In_35);
and U1614 (N_1614,In_574,In_697);
and U1615 (N_1615,In_71,In_207);
or U1616 (N_1616,In_541,In_67);
nand U1617 (N_1617,In_250,In_632);
or U1618 (N_1618,In_706,In_35);
xor U1619 (N_1619,In_294,In_182);
or U1620 (N_1620,In_65,In_467);
and U1621 (N_1621,In_462,In_463);
or U1622 (N_1622,In_312,In_310);
or U1623 (N_1623,In_413,In_91);
nor U1624 (N_1624,In_292,In_212);
nand U1625 (N_1625,In_46,In_302);
nand U1626 (N_1626,In_134,In_20);
or U1627 (N_1627,In_631,In_42);
nand U1628 (N_1628,In_336,In_42);
or U1629 (N_1629,In_83,In_320);
or U1630 (N_1630,In_361,In_271);
or U1631 (N_1631,In_65,In_286);
and U1632 (N_1632,In_578,In_57);
and U1633 (N_1633,In_528,In_68);
or U1634 (N_1634,In_579,In_585);
or U1635 (N_1635,In_392,In_457);
or U1636 (N_1636,In_465,In_152);
and U1637 (N_1637,In_156,In_550);
nor U1638 (N_1638,In_295,In_278);
nand U1639 (N_1639,In_76,In_355);
or U1640 (N_1640,In_291,In_398);
and U1641 (N_1641,In_596,In_136);
or U1642 (N_1642,In_678,In_447);
and U1643 (N_1643,In_626,In_351);
nand U1644 (N_1644,In_38,In_63);
nor U1645 (N_1645,In_554,In_158);
or U1646 (N_1646,In_689,In_369);
and U1647 (N_1647,In_345,In_717);
or U1648 (N_1648,In_83,In_30);
or U1649 (N_1649,In_326,In_197);
or U1650 (N_1650,In_623,In_333);
and U1651 (N_1651,In_748,In_147);
and U1652 (N_1652,In_634,In_736);
or U1653 (N_1653,In_93,In_134);
and U1654 (N_1654,In_420,In_667);
or U1655 (N_1655,In_739,In_262);
or U1656 (N_1656,In_52,In_609);
nor U1657 (N_1657,In_386,In_178);
nor U1658 (N_1658,In_704,In_679);
nand U1659 (N_1659,In_612,In_39);
nor U1660 (N_1660,In_532,In_61);
nor U1661 (N_1661,In_142,In_490);
or U1662 (N_1662,In_623,In_434);
nand U1663 (N_1663,In_290,In_596);
or U1664 (N_1664,In_354,In_357);
nand U1665 (N_1665,In_27,In_57);
nand U1666 (N_1666,In_276,In_44);
nand U1667 (N_1667,In_109,In_21);
nor U1668 (N_1668,In_481,In_506);
nor U1669 (N_1669,In_731,In_354);
or U1670 (N_1670,In_695,In_383);
and U1671 (N_1671,In_718,In_136);
or U1672 (N_1672,In_393,In_411);
nand U1673 (N_1673,In_710,In_202);
or U1674 (N_1674,In_746,In_731);
nor U1675 (N_1675,In_733,In_166);
nand U1676 (N_1676,In_156,In_346);
or U1677 (N_1677,In_569,In_549);
nand U1678 (N_1678,In_678,In_202);
nor U1679 (N_1679,In_58,In_507);
or U1680 (N_1680,In_72,In_293);
nand U1681 (N_1681,In_539,In_115);
nand U1682 (N_1682,In_77,In_315);
and U1683 (N_1683,In_683,In_10);
and U1684 (N_1684,In_367,In_167);
and U1685 (N_1685,In_196,In_324);
and U1686 (N_1686,In_234,In_580);
nand U1687 (N_1687,In_397,In_622);
nor U1688 (N_1688,In_403,In_386);
and U1689 (N_1689,In_525,In_388);
and U1690 (N_1690,In_497,In_606);
nand U1691 (N_1691,In_300,In_551);
nor U1692 (N_1692,In_536,In_3);
nand U1693 (N_1693,In_24,In_704);
and U1694 (N_1694,In_275,In_336);
nand U1695 (N_1695,In_6,In_249);
and U1696 (N_1696,In_294,In_499);
nand U1697 (N_1697,In_270,In_710);
and U1698 (N_1698,In_654,In_305);
nor U1699 (N_1699,In_50,In_565);
and U1700 (N_1700,In_3,In_127);
nand U1701 (N_1701,In_734,In_23);
nor U1702 (N_1702,In_392,In_651);
or U1703 (N_1703,In_648,In_410);
nor U1704 (N_1704,In_176,In_701);
nor U1705 (N_1705,In_477,In_730);
or U1706 (N_1706,In_308,In_10);
xnor U1707 (N_1707,In_127,In_191);
nor U1708 (N_1708,In_183,In_597);
nor U1709 (N_1709,In_257,In_228);
nor U1710 (N_1710,In_228,In_476);
and U1711 (N_1711,In_17,In_663);
nand U1712 (N_1712,In_394,In_29);
xnor U1713 (N_1713,In_488,In_660);
nand U1714 (N_1714,In_587,In_611);
nand U1715 (N_1715,In_468,In_220);
nor U1716 (N_1716,In_739,In_340);
nor U1717 (N_1717,In_94,In_417);
nand U1718 (N_1718,In_188,In_632);
and U1719 (N_1719,In_367,In_398);
and U1720 (N_1720,In_42,In_313);
nand U1721 (N_1721,In_322,In_269);
and U1722 (N_1722,In_200,In_343);
nand U1723 (N_1723,In_156,In_186);
nor U1724 (N_1724,In_423,In_60);
and U1725 (N_1725,In_325,In_557);
nand U1726 (N_1726,In_233,In_128);
nor U1727 (N_1727,In_549,In_244);
and U1728 (N_1728,In_123,In_78);
or U1729 (N_1729,In_53,In_402);
or U1730 (N_1730,In_365,In_169);
and U1731 (N_1731,In_212,In_463);
and U1732 (N_1732,In_129,In_431);
nor U1733 (N_1733,In_668,In_663);
or U1734 (N_1734,In_593,In_100);
nor U1735 (N_1735,In_287,In_198);
or U1736 (N_1736,In_73,In_296);
nand U1737 (N_1737,In_97,In_716);
or U1738 (N_1738,In_14,In_249);
and U1739 (N_1739,In_102,In_544);
or U1740 (N_1740,In_633,In_545);
nor U1741 (N_1741,In_19,In_465);
nor U1742 (N_1742,In_41,In_233);
nand U1743 (N_1743,In_299,In_357);
nor U1744 (N_1744,In_228,In_480);
nand U1745 (N_1745,In_727,In_466);
nand U1746 (N_1746,In_124,In_556);
or U1747 (N_1747,In_635,In_251);
and U1748 (N_1748,In_115,In_668);
nor U1749 (N_1749,In_736,In_129);
and U1750 (N_1750,In_330,In_6);
nor U1751 (N_1751,In_550,In_52);
or U1752 (N_1752,In_421,In_699);
and U1753 (N_1753,In_269,In_566);
and U1754 (N_1754,In_154,In_115);
nor U1755 (N_1755,In_132,In_737);
nor U1756 (N_1756,In_165,In_591);
xor U1757 (N_1757,In_153,In_84);
or U1758 (N_1758,In_305,In_166);
or U1759 (N_1759,In_504,In_571);
nor U1760 (N_1760,In_475,In_707);
and U1761 (N_1761,In_405,In_462);
or U1762 (N_1762,In_687,In_632);
or U1763 (N_1763,In_473,In_588);
nand U1764 (N_1764,In_267,In_217);
and U1765 (N_1765,In_136,In_648);
and U1766 (N_1766,In_644,In_352);
and U1767 (N_1767,In_651,In_84);
nor U1768 (N_1768,In_560,In_544);
nand U1769 (N_1769,In_460,In_445);
nor U1770 (N_1770,In_1,In_183);
nor U1771 (N_1771,In_92,In_275);
nand U1772 (N_1772,In_547,In_517);
nand U1773 (N_1773,In_108,In_72);
nand U1774 (N_1774,In_538,In_668);
and U1775 (N_1775,In_141,In_182);
or U1776 (N_1776,In_679,In_727);
nor U1777 (N_1777,In_513,In_37);
nor U1778 (N_1778,In_34,In_577);
and U1779 (N_1779,In_665,In_367);
nor U1780 (N_1780,In_229,In_186);
nor U1781 (N_1781,In_310,In_682);
nor U1782 (N_1782,In_50,In_392);
and U1783 (N_1783,In_505,In_331);
or U1784 (N_1784,In_348,In_461);
and U1785 (N_1785,In_433,In_571);
nor U1786 (N_1786,In_685,In_703);
or U1787 (N_1787,In_559,In_594);
nor U1788 (N_1788,In_576,In_364);
nand U1789 (N_1789,In_624,In_425);
nor U1790 (N_1790,In_346,In_24);
or U1791 (N_1791,In_682,In_322);
and U1792 (N_1792,In_590,In_529);
nand U1793 (N_1793,In_136,In_81);
nor U1794 (N_1794,In_455,In_693);
and U1795 (N_1795,In_589,In_165);
and U1796 (N_1796,In_279,In_548);
nand U1797 (N_1797,In_110,In_714);
or U1798 (N_1798,In_598,In_513);
nand U1799 (N_1799,In_330,In_222);
and U1800 (N_1800,In_85,In_672);
nand U1801 (N_1801,In_400,In_251);
and U1802 (N_1802,In_486,In_513);
nor U1803 (N_1803,In_515,In_16);
and U1804 (N_1804,In_414,In_124);
and U1805 (N_1805,In_498,In_454);
or U1806 (N_1806,In_170,In_252);
and U1807 (N_1807,In_408,In_228);
nand U1808 (N_1808,In_446,In_748);
and U1809 (N_1809,In_232,In_88);
nor U1810 (N_1810,In_262,In_721);
nand U1811 (N_1811,In_259,In_220);
or U1812 (N_1812,In_170,In_400);
or U1813 (N_1813,In_428,In_265);
nand U1814 (N_1814,In_216,In_28);
nor U1815 (N_1815,In_299,In_330);
or U1816 (N_1816,In_709,In_250);
nand U1817 (N_1817,In_198,In_646);
and U1818 (N_1818,In_66,In_641);
nand U1819 (N_1819,In_45,In_327);
nand U1820 (N_1820,In_35,In_216);
or U1821 (N_1821,In_682,In_710);
or U1822 (N_1822,In_620,In_313);
nand U1823 (N_1823,In_188,In_283);
or U1824 (N_1824,In_382,In_683);
or U1825 (N_1825,In_83,In_179);
or U1826 (N_1826,In_68,In_205);
nor U1827 (N_1827,In_733,In_700);
nor U1828 (N_1828,In_524,In_441);
and U1829 (N_1829,In_509,In_296);
or U1830 (N_1830,In_705,In_231);
nand U1831 (N_1831,In_94,In_344);
or U1832 (N_1832,In_527,In_685);
and U1833 (N_1833,In_6,In_439);
and U1834 (N_1834,In_199,In_174);
or U1835 (N_1835,In_275,In_164);
or U1836 (N_1836,In_26,In_611);
nand U1837 (N_1837,In_126,In_502);
or U1838 (N_1838,In_425,In_21);
nand U1839 (N_1839,In_163,In_193);
or U1840 (N_1840,In_114,In_93);
and U1841 (N_1841,In_286,In_221);
and U1842 (N_1842,In_677,In_271);
and U1843 (N_1843,In_471,In_90);
or U1844 (N_1844,In_255,In_24);
nand U1845 (N_1845,In_421,In_162);
xnor U1846 (N_1846,In_102,In_243);
or U1847 (N_1847,In_248,In_482);
and U1848 (N_1848,In_322,In_655);
and U1849 (N_1849,In_407,In_629);
or U1850 (N_1850,In_715,In_426);
nor U1851 (N_1851,In_396,In_190);
nand U1852 (N_1852,In_367,In_196);
nand U1853 (N_1853,In_743,In_523);
or U1854 (N_1854,In_565,In_225);
or U1855 (N_1855,In_78,In_243);
nand U1856 (N_1856,In_136,In_122);
nand U1857 (N_1857,In_718,In_685);
nand U1858 (N_1858,In_183,In_722);
or U1859 (N_1859,In_481,In_651);
and U1860 (N_1860,In_62,In_543);
or U1861 (N_1861,In_24,In_157);
nor U1862 (N_1862,In_230,In_591);
and U1863 (N_1863,In_106,In_355);
and U1864 (N_1864,In_27,In_566);
or U1865 (N_1865,In_125,In_638);
nor U1866 (N_1866,In_610,In_427);
nor U1867 (N_1867,In_366,In_345);
nor U1868 (N_1868,In_223,In_27);
nand U1869 (N_1869,In_595,In_56);
or U1870 (N_1870,In_18,In_86);
nor U1871 (N_1871,In_649,In_492);
xnor U1872 (N_1872,In_569,In_279);
or U1873 (N_1873,In_648,In_537);
nand U1874 (N_1874,In_400,In_202);
or U1875 (N_1875,In_594,In_386);
and U1876 (N_1876,In_217,In_137);
nand U1877 (N_1877,In_530,In_514);
nor U1878 (N_1878,In_467,In_617);
or U1879 (N_1879,In_584,In_748);
nand U1880 (N_1880,In_699,In_150);
nand U1881 (N_1881,In_178,In_283);
and U1882 (N_1882,In_562,In_497);
nor U1883 (N_1883,In_656,In_509);
nor U1884 (N_1884,In_697,In_735);
or U1885 (N_1885,In_112,In_619);
nor U1886 (N_1886,In_129,In_447);
nor U1887 (N_1887,In_538,In_10);
and U1888 (N_1888,In_385,In_648);
nor U1889 (N_1889,In_350,In_126);
or U1890 (N_1890,In_46,In_108);
nand U1891 (N_1891,In_480,In_331);
and U1892 (N_1892,In_595,In_157);
and U1893 (N_1893,In_725,In_400);
or U1894 (N_1894,In_100,In_542);
or U1895 (N_1895,In_166,In_42);
or U1896 (N_1896,In_584,In_413);
nand U1897 (N_1897,In_249,In_180);
and U1898 (N_1898,In_498,In_624);
and U1899 (N_1899,In_282,In_595);
or U1900 (N_1900,In_409,In_188);
and U1901 (N_1901,In_186,In_380);
nand U1902 (N_1902,In_587,In_597);
and U1903 (N_1903,In_7,In_600);
and U1904 (N_1904,In_195,In_21);
and U1905 (N_1905,In_245,In_76);
or U1906 (N_1906,In_673,In_679);
and U1907 (N_1907,In_177,In_423);
or U1908 (N_1908,In_125,In_235);
nand U1909 (N_1909,In_642,In_296);
nand U1910 (N_1910,In_524,In_637);
and U1911 (N_1911,In_421,In_588);
or U1912 (N_1912,In_100,In_610);
or U1913 (N_1913,In_700,In_531);
and U1914 (N_1914,In_510,In_24);
nor U1915 (N_1915,In_598,In_744);
or U1916 (N_1916,In_191,In_455);
nor U1917 (N_1917,In_605,In_726);
nand U1918 (N_1918,In_190,In_350);
nor U1919 (N_1919,In_492,In_259);
and U1920 (N_1920,In_68,In_184);
nand U1921 (N_1921,In_686,In_87);
nor U1922 (N_1922,In_42,In_172);
nor U1923 (N_1923,In_417,In_246);
nor U1924 (N_1924,In_250,In_123);
or U1925 (N_1925,In_736,In_14);
nor U1926 (N_1926,In_717,In_458);
and U1927 (N_1927,In_632,In_56);
nand U1928 (N_1928,In_322,In_216);
nor U1929 (N_1929,In_88,In_259);
nor U1930 (N_1930,In_550,In_668);
and U1931 (N_1931,In_138,In_699);
nor U1932 (N_1932,In_481,In_714);
nor U1933 (N_1933,In_423,In_277);
or U1934 (N_1934,In_654,In_643);
nand U1935 (N_1935,In_743,In_342);
nand U1936 (N_1936,In_710,In_222);
or U1937 (N_1937,In_535,In_144);
or U1938 (N_1938,In_81,In_462);
or U1939 (N_1939,In_209,In_366);
or U1940 (N_1940,In_342,In_625);
nand U1941 (N_1941,In_74,In_101);
nor U1942 (N_1942,In_713,In_451);
or U1943 (N_1943,In_617,In_268);
and U1944 (N_1944,In_569,In_1);
and U1945 (N_1945,In_336,In_205);
nor U1946 (N_1946,In_583,In_380);
or U1947 (N_1947,In_518,In_65);
or U1948 (N_1948,In_22,In_284);
and U1949 (N_1949,In_290,In_681);
nor U1950 (N_1950,In_246,In_257);
nand U1951 (N_1951,In_636,In_44);
and U1952 (N_1952,In_629,In_458);
nor U1953 (N_1953,In_180,In_181);
nor U1954 (N_1954,In_130,In_589);
nand U1955 (N_1955,In_541,In_91);
or U1956 (N_1956,In_288,In_347);
nor U1957 (N_1957,In_700,In_148);
and U1958 (N_1958,In_612,In_647);
xnor U1959 (N_1959,In_598,In_601);
and U1960 (N_1960,In_373,In_694);
nor U1961 (N_1961,In_258,In_193);
or U1962 (N_1962,In_532,In_95);
or U1963 (N_1963,In_518,In_583);
nor U1964 (N_1964,In_180,In_522);
nand U1965 (N_1965,In_324,In_592);
nor U1966 (N_1966,In_636,In_647);
or U1967 (N_1967,In_70,In_701);
or U1968 (N_1968,In_620,In_266);
or U1969 (N_1969,In_271,In_45);
and U1970 (N_1970,In_293,In_700);
and U1971 (N_1971,In_361,In_184);
and U1972 (N_1972,In_84,In_129);
nor U1973 (N_1973,In_660,In_410);
nand U1974 (N_1974,In_502,In_631);
nor U1975 (N_1975,In_155,In_280);
and U1976 (N_1976,In_200,In_163);
or U1977 (N_1977,In_342,In_748);
nor U1978 (N_1978,In_605,In_485);
and U1979 (N_1979,In_685,In_679);
or U1980 (N_1980,In_382,In_240);
nor U1981 (N_1981,In_445,In_147);
nor U1982 (N_1982,In_349,In_705);
or U1983 (N_1983,In_5,In_566);
nor U1984 (N_1984,In_562,In_494);
or U1985 (N_1985,In_603,In_230);
nand U1986 (N_1986,In_533,In_51);
and U1987 (N_1987,In_429,In_526);
and U1988 (N_1988,In_350,In_618);
or U1989 (N_1989,In_237,In_55);
and U1990 (N_1990,In_709,In_122);
nand U1991 (N_1991,In_633,In_213);
nand U1992 (N_1992,In_86,In_493);
or U1993 (N_1993,In_536,In_15);
and U1994 (N_1994,In_629,In_281);
nor U1995 (N_1995,In_106,In_390);
nor U1996 (N_1996,In_624,In_79);
or U1997 (N_1997,In_451,In_106);
nor U1998 (N_1998,In_150,In_411);
and U1999 (N_1999,In_255,In_436);
or U2000 (N_2000,In_393,In_559);
or U2001 (N_2001,In_454,In_294);
and U2002 (N_2002,In_352,In_298);
nand U2003 (N_2003,In_605,In_599);
and U2004 (N_2004,In_86,In_343);
nor U2005 (N_2005,In_610,In_160);
or U2006 (N_2006,In_725,In_146);
nor U2007 (N_2007,In_615,In_520);
and U2008 (N_2008,In_45,In_747);
and U2009 (N_2009,In_486,In_503);
or U2010 (N_2010,In_31,In_337);
nand U2011 (N_2011,In_184,In_264);
and U2012 (N_2012,In_77,In_306);
or U2013 (N_2013,In_718,In_738);
and U2014 (N_2014,In_20,In_427);
nand U2015 (N_2015,In_309,In_749);
and U2016 (N_2016,In_282,In_702);
and U2017 (N_2017,In_301,In_719);
and U2018 (N_2018,In_243,In_627);
or U2019 (N_2019,In_347,In_585);
or U2020 (N_2020,In_499,In_472);
nand U2021 (N_2021,In_516,In_102);
or U2022 (N_2022,In_71,In_414);
and U2023 (N_2023,In_199,In_23);
or U2024 (N_2024,In_185,In_153);
nand U2025 (N_2025,In_96,In_600);
nor U2026 (N_2026,In_456,In_17);
and U2027 (N_2027,In_341,In_540);
xor U2028 (N_2028,In_320,In_148);
or U2029 (N_2029,In_225,In_3);
nand U2030 (N_2030,In_178,In_170);
and U2031 (N_2031,In_386,In_167);
nand U2032 (N_2032,In_221,In_162);
nand U2033 (N_2033,In_23,In_146);
nand U2034 (N_2034,In_236,In_134);
nand U2035 (N_2035,In_44,In_148);
nand U2036 (N_2036,In_356,In_111);
or U2037 (N_2037,In_410,In_34);
or U2038 (N_2038,In_501,In_474);
nand U2039 (N_2039,In_274,In_247);
nor U2040 (N_2040,In_207,In_708);
nand U2041 (N_2041,In_678,In_483);
nand U2042 (N_2042,In_560,In_171);
nor U2043 (N_2043,In_142,In_428);
and U2044 (N_2044,In_593,In_500);
or U2045 (N_2045,In_53,In_650);
xnor U2046 (N_2046,In_342,In_687);
or U2047 (N_2047,In_230,In_402);
nand U2048 (N_2048,In_659,In_690);
nor U2049 (N_2049,In_42,In_270);
nor U2050 (N_2050,In_183,In_38);
and U2051 (N_2051,In_425,In_49);
or U2052 (N_2052,In_358,In_638);
or U2053 (N_2053,In_121,In_521);
or U2054 (N_2054,In_697,In_487);
nand U2055 (N_2055,In_535,In_222);
or U2056 (N_2056,In_465,In_2);
nand U2057 (N_2057,In_470,In_677);
or U2058 (N_2058,In_522,In_29);
nand U2059 (N_2059,In_17,In_671);
and U2060 (N_2060,In_125,In_178);
and U2061 (N_2061,In_660,In_477);
nand U2062 (N_2062,In_64,In_716);
nor U2063 (N_2063,In_378,In_457);
and U2064 (N_2064,In_190,In_422);
or U2065 (N_2065,In_157,In_286);
or U2066 (N_2066,In_217,In_36);
or U2067 (N_2067,In_560,In_330);
nand U2068 (N_2068,In_218,In_390);
nand U2069 (N_2069,In_421,In_47);
nand U2070 (N_2070,In_102,In_354);
nor U2071 (N_2071,In_543,In_64);
and U2072 (N_2072,In_30,In_57);
or U2073 (N_2073,In_303,In_107);
or U2074 (N_2074,In_521,In_344);
or U2075 (N_2075,In_336,In_571);
or U2076 (N_2076,In_489,In_211);
and U2077 (N_2077,In_611,In_200);
nand U2078 (N_2078,In_24,In_466);
or U2079 (N_2079,In_745,In_308);
nand U2080 (N_2080,In_275,In_599);
and U2081 (N_2081,In_509,In_15);
nor U2082 (N_2082,In_602,In_178);
and U2083 (N_2083,In_454,In_348);
and U2084 (N_2084,In_167,In_184);
nand U2085 (N_2085,In_157,In_234);
nand U2086 (N_2086,In_402,In_495);
and U2087 (N_2087,In_673,In_350);
and U2088 (N_2088,In_382,In_533);
nor U2089 (N_2089,In_435,In_587);
nand U2090 (N_2090,In_257,In_277);
nor U2091 (N_2091,In_425,In_165);
nor U2092 (N_2092,In_143,In_426);
nor U2093 (N_2093,In_592,In_747);
nor U2094 (N_2094,In_307,In_130);
or U2095 (N_2095,In_10,In_547);
nand U2096 (N_2096,In_216,In_14);
and U2097 (N_2097,In_100,In_504);
nand U2098 (N_2098,In_701,In_470);
and U2099 (N_2099,In_738,In_277);
nor U2100 (N_2100,In_61,In_748);
or U2101 (N_2101,In_52,In_302);
and U2102 (N_2102,In_667,In_373);
or U2103 (N_2103,In_17,In_241);
or U2104 (N_2104,In_656,In_240);
nor U2105 (N_2105,In_472,In_699);
nand U2106 (N_2106,In_254,In_431);
or U2107 (N_2107,In_291,In_132);
and U2108 (N_2108,In_107,In_528);
nor U2109 (N_2109,In_469,In_61);
nand U2110 (N_2110,In_667,In_256);
nor U2111 (N_2111,In_432,In_351);
or U2112 (N_2112,In_371,In_749);
nand U2113 (N_2113,In_256,In_588);
and U2114 (N_2114,In_527,In_262);
and U2115 (N_2115,In_476,In_74);
and U2116 (N_2116,In_685,In_159);
nand U2117 (N_2117,In_204,In_522);
or U2118 (N_2118,In_470,In_657);
nor U2119 (N_2119,In_625,In_318);
nand U2120 (N_2120,In_536,In_562);
nor U2121 (N_2121,In_206,In_172);
or U2122 (N_2122,In_27,In_449);
or U2123 (N_2123,In_456,In_360);
or U2124 (N_2124,In_272,In_132);
nor U2125 (N_2125,In_721,In_438);
or U2126 (N_2126,In_210,In_579);
and U2127 (N_2127,In_390,In_328);
or U2128 (N_2128,In_651,In_264);
and U2129 (N_2129,In_715,In_716);
nand U2130 (N_2130,In_595,In_436);
or U2131 (N_2131,In_231,In_560);
nor U2132 (N_2132,In_147,In_242);
nand U2133 (N_2133,In_429,In_189);
and U2134 (N_2134,In_694,In_184);
or U2135 (N_2135,In_369,In_54);
nor U2136 (N_2136,In_6,In_78);
nor U2137 (N_2137,In_245,In_255);
and U2138 (N_2138,In_446,In_368);
and U2139 (N_2139,In_407,In_572);
or U2140 (N_2140,In_288,In_585);
and U2141 (N_2141,In_675,In_622);
nand U2142 (N_2142,In_22,In_233);
nor U2143 (N_2143,In_275,In_528);
and U2144 (N_2144,In_665,In_267);
or U2145 (N_2145,In_584,In_146);
nand U2146 (N_2146,In_377,In_693);
or U2147 (N_2147,In_103,In_611);
nand U2148 (N_2148,In_615,In_32);
or U2149 (N_2149,In_91,In_345);
and U2150 (N_2150,In_200,In_180);
nor U2151 (N_2151,In_2,In_421);
or U2152 (N_2152,In_113,In_303);
or U2153 (N_2153,In_176,In_719);
nor U2154 (N_2154,In_717,In_15);
nor U2155 (N_2155,In_58,In_672);
nor U2156 (N_2156,In_358,In_315);
nand U2157 (N_2157,In_546,In_596);
or U2158 (N_2158,In_63,In_264);
or U2159 (N_2159,In_380,In_272);
and U2160 (N_2160,In_145,In_148);
nand U2161 (N_2161,In_166,In_679);
nand U2162 (N_2162,In_295,In_588);
and U2163 (N_2163,In_67,In_421);
and U2164 (N_2164,In_661,In_58);
nand U2165 (N_2165,In_200,In_492);
and U2166 (N_2166,In_197,In_605);
xor U2167 (N_2167,In_558,In_149);
or U2168 (N_2168,In_168,In_398);
nand U2169 (N_2169,In_588,In_461);
and U2170 (N_2170,In_269,In_686);
and U2171 (N_2171,In_226,In_450);
and U2172 (N_2172,In_465,In_264);
nand U2173 (N_2173,In_5,In_442);
or U2174 (N_2174,In_389,In_359);
and U2175 (N_2175,In_338,In_671);
and U2176 (N_2176,In_44,In_649);
nor U2177 (N_2177,In_680,In_78);
or U2178 (N_2178,In_162,In_78);
and U2179 (N_2179,In_323,In_325);
xor U2180 (N_2180,In_458,In_596);
nand U2181 (N_2181,In_489,In_228);
or U2182 (N_2182,In_386,In_651);
and U2183 (N_2183,In_526,In_248);
or U2184 (N_2184,In_14,In_421);
and U2185 (N_2185,In_386,In_507);
and U2186 (N_2186,In_653,In_312);
and U2187 (N_2187,In_690,In_436);
and U2188 (N_2188,In_454,In_600);
nand U2189 (N_2189,In_450,In_215);
nand U2190 (N_2190,In_498,In_484);
nor U2191 (N_2191,In_148,In_719);
nand U2192 (N_2192,In_416,In_299);
nand U2193 (N_2193,In_556,In_354);
nor U2194 (N_2194,In_32,In_420);
and U2195 (N_2195,In_114,In_190);
or U2196 (N_2196,In_523,In_105);
or U2197 (N_2197,In_158,In_211);
or U2198 (N_2198,In_73,In_109);
nand U2199 (N_2199,In_275,In_665);
or U2200 (N_2200,In_426,In_253);
nor U2201 (N_2201,In_209,In_54);
nor U2202 (N_2202,In_123,In_630);
nand U2203 (N_2203,In_37,In_48);
and U2204 (N_2204,In_30,In_62);
nand U2205 (N_2205,In_222,In_247);
nand U2206 (N_2206,In_183,In_610);
nor U2207 (N_2207,In_731,In_491);
and U2208 (N_2208,In_415,In_83);
and U2209 (N_2209,In_49,In_377);
nor U2210 (N_2210,In_402,In_407);
or U2211 (N_2211,In_518,In_5);
nor U2212 (N_2212,In_392,In_448);
and U2213 (N_2213,In_23,In_258);
nand U2214 (N_2214,In_633,In_266);
nor U2215 (N_2215,In_638,In_99);
and U2216 (N_2216,In_681,In_249);
nand U2217 (N_2217,In_368,In_354);
or U2218 (N_2218,In_501,In_741);
or U2219 (N_2219,In_588,In_369);
or U2220 (N_2220,In_440,In_716);
or U2221 (N_2221,In_147,In_291);
nor U2222 (N_2222,In_468,In_23);
nand U2223 (N_2223,In_509,In_455);
or U2224 (N_2224,In_580,In_547);
or U2225 (N_2225,In_116,In_202);
or U2226 (N_2226,In_460,In_48);
and U2227 (N_2227,In_376,In_378);
nor U2228 (N_2228,In_96,In_71);
and U2229 (N_2229,In_535,In_213);
and U2230 (N_2230,In_268,In_683);
nand U2231 (N_2231,In_48,In_594);
or U2232 (N_2232,In_449,In_703);
nor U2233 (N_2233,In_552,In_398);
nor U2234 (N_2234,In_675,In_723);
and U2235 (N_2235,In_591,In_349);
nand U2236 (N_2236,In_214,In_350);
and U2237 (N_2237,In_516,In_668);
or U2238 (N_2238,In_477,In_425);
and U2239 (N_2239,In_6,In_437);
nor U2240 (N_2240,In_345,In_291);
nand U2241 (N_2241,In_126,In_196);
nor U2242 (N_2242,In_63,In_346);
and U2243 (N_2243,In_591,In_652);
nand U2244 (N_2244,In_243,In_298);
and U2245 (N_2245,In_267,In_412);
nor U2246 (N_2246,In_554,In_560);
nand U2247 (N_2247,In_506,In_736);
nand U2248 (N_2248,In_304,In_654);
nand U2249 (N_2249,In_657,In_208);
and U2250 (N_2250,In_20,In_611);
and U2251 (N_2251,In_524,In_94);
nor U2252 (N_2252,In_615,In_360);
and U2253 (N_2253,In_686,In_667);
or U2254 (N_2254,In_41,In_592);
nand U2255 (N_2255,In_455,In_271);
nand U2256 (N_2256,In_533,In_476);
nand U2257 (N_2257,In_474,In_536);
and U2258 (N_2258,In_690,In_700);
or U2259 (N_2259,In_416,In_320);
and U2260 (N_2260,In_479,In_598);
nand U2261 (N_2261,In_652,In_5);
and U2262 (N_2262,In_73,In_626);
nor U2263 (N_2263,In_147,In_451);
xnor U2264 (N_2264,In_207,In_480);
and U2265 (N_2265,In_100,In_349);
nand U2266 (N_2266,In_515,In_178);
and U2267 (N_2267,In_679,In_740);
and U2268 (N_2268,In_67,In_672);
and U2269 (N_2269,In_683,In_131);
nor U2270 (N_2270,In_649,In_158);
nand U2271 (N_2271,In_409,In_59);
nand U2272 (N_2272,In_325,In_567);
nor U2273 (N_2273,In_47,In_104);
nand U2274 (N_2274,In_118,In_257);
nand U2275 (N_2275,In_2,In_345);
nand U2276 (N_2276,In_424,In_748);
nor U2277 (N_2277,In_227,In_244);
and U2278 (N_2278,In_349,In_16);
nand U2279 (N_2279,In_705,In_426);
and U2280 (N_2280,In_36,In_664);
nand U2281 (N_2281,In_698,In_352);
nand U2282 (N_2282,In_489,In_356);
nor U2283 (N_2283,In_586,In_475);
nand U2284 (N_2284,In_106,In_149);
and U2285 (N_2285,In_137,In_474);
nor U2286 (N_2286,In_707,In_182);
and U2287 (N_2287,In_323,In_545);
and U2288 (N_2288,In_547,In_251);
nand U2289 (N_2289,In_167,In_682);
and U2290 (N_2290,In_234,In_160);
or U2291 (N_2291,In_97,In_732);
nor U2292 (N_2292,In_271,In_17);
nor U2293 (N_2293,In_135,In_36);
and U2294 (N_2294,In_89,In_229);
and U2295 (N_2295,In_519,In_71);
nor U2296 (N_2296,In_81,In_290);
and U2297 (N_2297,In_353,In_626);
nand U2298 (N_2298,In_513,In_653);
or U2299 (N_2299,In_273,In_221);
or U2300 (N_2300,In_374,In_504);
and U2301 (N_2301,In_553,In_615);
or U2302 (N_2302,In_63,In_158);
and U2303 (N_2303,In_599,In_580);
nor U2304 (N_2304,In_247,In_748);
and U2305 (N_2305,In_574,In_702);
and U2306 (N_2306,In_605,In_67);
or U2307 (N_2307,In_314,In_378);
nand U2308 (N_2308,In_717,In_267);
nor U2309 (N_2309,In_94,In_17);
nor U2310 (N_2310,In_323,In_168);
or U2311 (N_2311,In_202,In_141);
nor U2312 (N_2312,In_741,In_719);
and U2313 (N_2313,In_28,In_415);
nand U2314 (N_2314,In_517,In_492);
nor U2315 (N_2315,In_5,In_267);
or U2316 (N_2316,In_106,In_470);
and U2317 (N_2317,In_608,In_477);
nand U2318 (N_2318,In_486,In_396);
or U2319 (N_2319,In_148,In_38);
or U2320 (N_2320,In_599,In_717);
nor U2321 (N_2321,In_311,In_634);
nand U2322 (N_2322,In_330,In_511);
nand U2323 (N_2323,In_13,In_443);
nor U2324 (N_2324,In_626,In_693);
nor U2325 (N_2325,In_501,In_684);
nor U2326 (N_2326,In_489,In_173);
nand U2327 (N_2327,In_176,In_275);
nand U2328 (N_2328,In_683,In_103);
and U2329 (N_2329,In_143,In_219);
nor U2330 (N_2330,In_211,In_421);
nand U2331 (N_2331,In_53,In_191);
and U2332 (N_2332,In_712,In_531);
and U2333 (N_2333,In_514,In_151);
nor U2334 (N_2334,In_222,In_306);
or U2335 (N_2335,In_248,In_161);
nand U2336 (N_2336,In_571,In_44);
or U2337 (N_2337,In_699,In_333);
or U2338 (N_2338,In_248,In_397);
nand U2339 (N_2339,In_471,In_495);
nor U2340 (N_2340,In_125,In_176);
nand U2341 (N_2341,In_161,In_645);
nand U2342 (N_2342,In_745,In_252);
and U2343 (N_2343,In_484,In_515);
and U2344 (N_2344,In_537,In_140);
nor U2345 (N_2345,In_380,In_681);
nor U2346 (N_2346,In_684,In_648);
and U2347 (N_2347,In_328,In_629);
or U2348 (N_2348,In_628,In_134);
nor U2349 (N_2349,In_161,In_698);
nand U2350 (N_2350,In_420,In_262);
nor U2351 (N_2351,In_237,In_468);
nand U2352 (N_2352,In_308,In_573);
nor U2353 (N_2353,In_579,In_425);
or U2354 (N_2354,In_627,In_692);
nor U2355 (N_2355,In_58,In_683);
or U2356 (N_2356,In_630,In_222);
nand U2357 (N_2357,In_511,In_710);
or U2358 (N_2358,In_151,In_330);
nand U2359 (N_2359,In_708,In_725);
or U2360 (N_2360,In_548,In_579);
nor U2361 (N_2361,In_103,In_605);
or U2362 (N_2362,In_225,In_206);
and U2363 (N_2363,In_74,In_432);
nor U2364 (N_2364,In_705,In_602);
nor U2365 (N_2365,In_125,In_264);
xor U2366 (N_2366,In_535,In_581);
and U2367 (N_2367,In_570,In_693);
nand U2368 (N_2368,In_428,In_714);
and U2369 (N_2369,In_190,In_140);
and U2370 (N_2370,In_187,In_2);
nand U2371 (N_2371,In_390,In_47);
and U2372 (N_2372,In_545,In_658);
and U2373 (N_2373,In_732,In_550);
or U2374 (N_2374,In_563,In_116);
or U2375 (N_2375,In_558,In_477);
or U2376 (N_2376,In_719,In_24);
or U2377 (N_2377,In_375,In_125);
and U2378 (N_2378,In_360,In_396);
and U2379 (N_2379,In_133,In_458);
nand U2380 (N_2380,In_84,In_256);
or U2381 (N_2381,In_470,In_319);
nand U2382 (N_2382,In_419,In_454);
nand U2383 (N_2383,In_468,In_429);
nor U2384 (N_2384,In_507,In_410);
nor U2385 (N_2385,In_317,In_570);
nor U2386 (N_2386,In_185,In_680);
xnor U2387 (N_2387,In_733,In_668);
and U2388 (N_2388,In_209,In_484);
nor U2389 (N_2389,In_65,In_627);
nand U2390 (N_2390,In_186,In_216);
nor U2391 (N_2391,In_678,In_263);
and U2392 (N_2392,In_675,In_523);
and U2393 (N_2393,In_425,In_120);
or U2394 (N_2394,In_675,In_355);
nand U2395 (N_2395,In_332,In_652);
and U2396 (N_2396,In_558,In_50);
and U2397 (N_2397,In_726,In_404);
and U2398 (N_2398,In_725,In_484);
or U2399 (N_2399,In_613,In_577);
nand U2400 (N_2400,In_124,In_46);
nor U2401 (N_2401,In_20,In_387);
and U2402 (N_2402,In_389,In_562);
nor U2403 (N_2403,In_154,In_55);
or U2404 (N_2404,In_19,In_190);
nor U2405 (N_2405,In_219,In_62);
nand U2406 (N_2406,In_456,In_115);
nand U2407 (N_2407,In_21,In_695);
nand U2408 (N_2408,In_733,In_608);
nand U2409 (N_2409,In_224,In_373);
or U2410 (N_2410,In_253,In_47);
nand U2411 (N_2411,In_28,In_677);
and U2412 (N_2412,In_16,In_630);
nand U2413 (N_2413,In_110,In_530);
nand U2414 (N_2414,In_562,In_335);
nor U2415 (N_2415,In_282,In_431);
nand U2416 (N_2416,In_256,In_668);
nor U2417 (N_2417,In_590,In_586);
nor U2418 (N_2418,In_529,In_282);
and U2419 (N_2419,In_661,In_672);
or U2420 (N_2420,In_705,In_143);
nor U2421 (N_2421,In_682,In_420);
nor U2422 (N_2422,In_658,In_260);
nand U2423 (N_2423,In_250,In_451);
or U2424 (N_2424,In_335,In_644);
or U2425 (N_2425,In_606,In_25);
or U2426 (N_2426,In_489,In_728);
nand U2427 (N_2427,In_98,In_356);
nand U2428 (N_2428,In_630,In_609);
or U2429 (N_2429,In_261,In_80);
nand U2430 (N_2430,In_412,In_207);
nor U2431 (N_2431,In_86,In_129);
nand U2432 (N_2432,In_343,In_698);
or U2433 (N_2433,In_135,In_66);
and U2434 (N_2434,In_453,In_222);
or U2435 (N_2435,In_302,In_388);
and U2436 (N_2436,In_444,In_368);
and U2437 (N_2437,In_97,In_45);
or U2438 (N_2438,In_176,In_159);
nand U2439 (N_2439,In_127,In_352);
or U2440 (N_2440,In_515,In_367);
or U2441 (N_2441,In_650,In_626);
or U2442 (N_2442,In_178,In_165);
nand U2443 (N_2443,In_364,In_297);
nor U2444 (N_2444,In_377,In_68);
and U2445 (N_2445,In_426,In_538);
nor U2446 (N_2446,In_713,In_227);
nor U2447 (N_2447,In_377,In_641);
and U2448 (N_2448,In_278,In_388);
nand U2449 (N_2449,In_467,In_699);
nor U2450 (N_2450,In_393,In_502);
and U2451 (N_2451,In_31,In_444);
nor U2452 (N_2452,In_75,In_617);
or U2453 (N_2453,In_242,In_646);
and U2454 (N_2454,In_214,In_313);
and U2455 (N_2455,In_662,In_628);
nor U2456 (N_2456,In_426,In_451);
and U2457 (N_2457,In_208,In_554);
nor U2458 (N_2458,In_389,In_583);
and U2459 (N_2459,In_18,In_225);
nand U2460 (N_2460,In_709,In_654);
or U2461 (N_2461,In_717,In_371);
nand U2462 (N_2462,In_232,In_380);
nand U2463 (N_2463,In_108,In_651);
or U2464 (N_2464,In_572,In_244);
and U2465 (N_2465,In_523,In_607);
nand U2466 (N_2466,In_454,In_652);
or U2467 (N_2467,In_341,In_263);
and U2468 (N_2468,In_453,In_577);
nor U2469 (N_2469,In_470,In_398);
and U2470 (N_2470,In_663,In_618);
nand U2471 (N_2471,In_370,In_303);
or U2472 (N_2472,In_546,In_660);
nor U2473 (N_2473,In_281,In_363);
nor U2474 (N_2474,In_631,In_638);
nor U2475 (N_2475,In_332,In_413);
nand U2476 (N_2476,In_641,In_374);
or U2477 (N_2477,In_171,In_112);
or U2478 (N_2478,In_135,In_211);
nand U2479 (N_2479,In_294,In_44);
and U2480 (N_2480,In_86,In_568);
nor U2481 (N_2481,In_743,In_264);
or U2482 (N_2482,In_701,In_388);
nor U2483 (N_2483,In_512,In_128);
nor U2484 (N_2484,In_585,In_442);
and U2485 (N_2485,In_454,In_162);
and U2486 (N_2486,In_202,In_439);
and U2487 (N_2487,In_317,In_307);
nor U2488 (N_2488,In_395,In_371);
and U2489 (N_2489,In_372,In_471);
or U2490 (N_2490,In_402,In_425);
nand U2491 (N_2491,In_278,In_690);
or U2492 (N_2492,In_54,In_575);
and U2493 (N_2493,In_496,In_556);
or U2494 (N_2494,In_307,In_382);
or U2495 (N_2495,In_378,In_524);
nor U2496 (N_2496,In_270,In_453);
or U2497 (N_2497,In_477,In_699);
or U2498 (N_2498,In_57,In_222);
and U2499 (N_2499,In_696,In_723);
xor U2500 (N_2500,N_664,N_131);
or U2501 (N_2501,N_1022,N_2249);
nor U2502 (N_2502,N_2171,N_1632);
nand U2503 (N_2503,N_904,N_2243);
nor U2504 (N_2504,N_1815,N_799);
and U2505 (N_2505,N_1809,N_1360);
nand U2506 (N_2506,N_2302,N_171);
or U2507 (N_2507,N_519,N_2111);
nor U2508 (N_2508,N_1492,N_462);
nand U2509 (N_2509,N_2495,N_844);
nor U2510 (N_2510,N_794,N_782);
and U2511 (N_2511,N_193,N_1451);
nor U2512 (N_2512,N_672,N_1519);
nor U2513 (N_2513,N_528,N_1377);
nor U2514 (N_2514,N_1475,N_1418);
nor U2515 (N_2515,N_839,N_414);
nor U2516 (N_2516,N_638,N_1265);
and U2517 (N_2517,N_153,N_2319);
and U2518 (N_2518,N_2188,N_1134);
and U2519 (N_2519,N_360,N_681);
and U2520 (N_2520,N_1270,N_1738);
nor U2521 (N_2521,N_450,N_89);
or U2522 (N_2522,N_2436,N_2443);
nor U2523 (N_2523,N_41,N_1088);
nand U2524 (N_2524,N_1692,N_966);
and U2525 (N_2525,N_110,N_603);
or U2526 (N_2526,N_1476,N_751);
nand U2527 (N_2527,N_1294,N_1646);
or U2528 (N_2528,N_1822,N_768);
nor U2529 (N_2529,N_539,N_515);
nand U2530 (N_2530,N_1101,N_695);
nand U2531 (N_2531,N_1302,N_2140);
xnor U2532 (N_2532,N_125,N_1041);
or U2533 (N_2533,N_925,N_1080);
xnor U2534 (N_2534,N_692,N_1096);
or U2535 (N_2535,N_597,N_1702);
nand U2536 (N_2536,N_2290,N_2445);
nor U2537 (N_2537,N_823,N_1729);
or U2538 (N_2538,N_740,N_656);
nor U2539 (N_2539,N_1131,N_533);
nand U2540 (N_2540,N_31,N_811);
nand U2541 (N_2541,N_1526,N_1971);
and U2542 (N_2542,N_847,N_407);
nor U2543 (N_2543,N_1221,N_1261);
or U2544 (N_2544,N_480,N_1207);
or U2545 (N_2545,N_1517,N_1649);
and U2546 (N_2546,N_798,N_1356);
and U2547 (N_2547,N_854,N_315);
or U2548 (N_2548,N_1660,N_2077);
nor U2549 (N_2549,N_955,N_1549);
nor U2550 (N_2550,N_1706,N_831);
or U2551 (N_2551,N_2322,N_2204);
and U2552 (N_2552,N_2080,N_772);
nand U2553 (N_2553,N_649,N_1631);
and U2554 (N_2554,N_1239,N_253);
or U2555 (N_2555,N_60,N_1774);
and U2556 (N_2556,N_1500,N_401);
or U2557 (N_2557,N_2274,N_513);
nor U2558 (N_2558,N_1629,N_1453);
or U2559 (N_2559,N_424,N_1037);
or U2560 (N_2560,N_210,N_1769);
or U2561 (N_2561,N_1384,N_706);
nand U2562 (N_2562,N_94,N_749);
or U2563 (N_2563,N_2106,N_425);
nand U2564 (N_2564,N_2058,N_977);
nor U2565 (N_2565,N_1182,N_393);
nor U2566 (N_2566,N_444,N_71);
and U2567 (N_2567,N_227,N_1299);
nand U2568 (N_2568,N_1956,N_568);
nor U2569 (N_2569,N_1454,N_541);
nor U2570 (N_2570,N_1181,N_1054);
nor U2571 (N_2571,N_1189,N_1399);
nor U2572 (N_2572,N_1922,N_2202);
nand U2573 (N_2573,N_911,N_292);
nor U2574 (N_2574,N_1947,N_2063);
nor U2575 (N_2575,N_2345,N_349);
and U2576 (N_2576,N_116,N_2263);
and U2577 (N_2577,N_1613,N_2296);
or U2578 (N_2578,N_1503,N_1485);
and U2579 (N_2579,N_1657,N_2328);
and U2580 (N_2580,N_1557,N_1495);
and U2581 (N_2581,N_1627,N_1874);
nor U2582 (N_2582,N_1714,N_2374);
nor U2583 (N_2583,N_483,N_2219);
or U2584 (N_2584,N_1014,N_720);
nor U2585 (N_2585,N_2144,N_50);
nor U2586 (N_2586,N_867,N_1885);
nand U2587 (N_2587,N_19,N_687);
nand U2588 (N_2588,N_427,N_2121);
nor U2589 (N_2589,N_591,N_908);
nor U2590 (N_2590,N_1634,N_1001);
and U2591 (N_2591,N_1522,N_1183);
and U2592 (N_2592,N_1919,N_1044);
or U2593 (N_2593,N_374,N_2360);
nor U2594 (N_2594,N_832,N_1295);
nand U2595 (N_2595,N_506,N_1925);
or U2596 (N_2596,N_1565,N_1090);
and U2597 (N_2597,N_228,N_946);
nor U2598 (N_2598,N_2254,N_454);
nor U2599 (N_2599,N_1915,N_1471);
nor U2600 (N_2600,N_1621,N_49);
nor U2601 (N_2601,N_268,N_1619);
and U2602 (N_2602,N_574,N_939);
or U2603 (N_2603,N_2371,N_181);
and U2604 (N_2604,N_2057,N_1078);
and U2605 (N_2605,N_2275,N_1029);
or U2606 (N_2606,N_1857,N_1380);
or U2607 (N_2607,N_884,N_1313);
and U2608 (N_2608,N_1846,N_113);
or U2609 (N_2609,N_792,N_2124);
nor U2610 (N_2610,N_366,N_203);
nor U2611 (N_2611,N_1970,N_93);
or U2612 (N_2612,N_284,N_775);
and U2613 (N_2613,N_367,N_2075);
nor U2614 (N_2614,N_371,N_891);
nor U2615 (N_2615,N_2220,N_916);
or U2616 (N_2616,N_129,N_452);
nor U2617 (N_2617,N_2242,N_2133);
nand U2618 (N_2618,N_1378,N_912);
or U2619 (N_2619,N_245,N_1048);
and U2620 (N_2620,N_1905,N_752);
or U2621 (N_2621,N_469,N_1833);
nand U2622 (N_2622,N_2348,N_1260);
nand U2623 (N_2623,N_2422,N_573);
nor U2624 (N_2624,N_1094,N_376);
and U2625 (N_2625,N_1154,N_1208);
nor U2626 (N_2626,N_1287,N_492);
or U2627 (N_2627,N_763,N_1891);
nor U2628 (N_2628,N_753,N_279);
nor U2629 (N_2629,N_679,N_2136);
or U2630 (N_2630,N_363,N_187);
nand U2631 (N_2631,N_1830,N_1862);
and U2632 (N_2632,N_2480,N_883);
nor U2633 (N_2633,N_1811,N_1580);
or U2634 (N_2634,N_460,N_1367);
nor U2635 (N_2635,N_1123,N_2143);
xor U2636 (N_2636,N_1750,N_886);
nor U2637 (N_2637,N_600,N_442);
or U2638 (N_2638,N_2245,N_2320);
nor U2639 (N_2639,N_1490,N_805);
and U2640 (N_2640,N_824,N_1249);
xor U2641 (N_2641,N_170,N_39);
and U2642 (N_2642,N_1608,N_1);
nor U2643 (N_2643,N_422,N_1355);
nor U2644 (N_2644,N_1494,N_1444);
nand U2645 (N_2645,N_1537,N_1117);
nor U2646 (N_2646,N_2305,N_1006);
or U2647 (N_2647,N_2358,N_431);
or U2648 (N_2648,N_310,N_777);
and U2649 (N_2649,N_2457,N_1257);
or U2650 (N_2650,N_107,N_2336);
nand U2651 (N_2651,N_261,N_846);
nand U2652 (N_2652,N_2011,N_1344);
and U2653 (N_2653,N_2064,N_953);
or U2654 (N_2654,N_249,N_2247);
nor U2655 (N_2655,N_625,N_567);
and U2656 (N_2656,N_379,N_489);
or U2657 (N_2657,N_267,N_739);
nor U2658 (N_2658,N_377,N_4);
and U2659 (N_2659,N_156,N_2496);
nand U2660 (N_2660,N_1800,N_1732);
nand U2661 (N_2661,N_1593,N_570);
nor U2662 (N_2662,N_269,N_1902);
and U2663 (N_2663,N_905,N_184);
and U2664 (N_2664,N_791,N_224);
nand U2665 (N_2665,N_2309,N_1171);
or U2666 (N_2666,N_1814,N_1097);
nor U2667 (N_2667,N_2197,N_608);
or U2668 (N_2668,N_1720,N_1013);
nor U2669 (N_2669,N_1895,N_578);
nand U2670 (N_2670,N_2375,N_1733);
nand U2671 (N_2671,N_1790,N_1338);
and U2672 (N_2672,N_12,N_1734);
nand U2673 (N_2673,N_339,N_2353);
or U2674 (N_2674,N_2180,N_1887);
nor U2675 (N_2675,N_252,N_2450);
nor U2676 (N_2676,N_1335,N_77);
nand U2677 (N_2677,N_1039,N_816);
nand U2678 (N_2678,N_2,N_481);
or U2679 (N_2679,N_1264,N_1170);
nor U2680 (N_2680,N_1327,N_1510);
nand U2681 (N_2681,N_1056,N_2205);
nand U2682 (N_2682,N_2287,N_938);
nand U2683 (N_2683,N_1528,N_1986);
or U2684 (N_2684,N_2122,N_714);
nand U2685 (N_2685,N_1047,N_1877);
nor U2686 (N_2686,N_2034,N_2303);
or U2687 (N_2687,N_1879,N_2065);
nor U2688 (N_2688,N_434,N_935);
and U2689 (N_2689,N_1076,N_343);
and U2690 (N_2690,N_877,N_1177);
nor U2691 (N_2691,N_1673,N_72);
nand U2692 (N_2692,N_1268,N_150);
nand U2693 (N_2693,N_2300,N_2473);
and U2694 (N_2694,N_974,N_1550);
and U2695 (N_2695,N_1408,N_748);
nor U2696 (N_2696,N_958,N_728);
or U2697 (N_2697,N_853,N_1553);
nor U2698 (N_2698,N_1841,N_561);
nor U2699 (N_2699,N_28,N_731);
nor U2700 (N_2700,N_2331,N_1026);
nor U2701 (N_2701,N_1278,N_1369);
nand U2702 (N_2702,N_1043,N_1897);
or U2703 (N_2703,N_2493,N_1643);
and U2704 (N_2704,N_2250,N_395);
and U2705 (N_2705,N_2039,N_810);
and U2706 (N_2706,N_1405,N_464);
or U2707 (N_2707,N_1577,N_1403);
and U2708 (N_2708,N_614,N_286);
nand U2709 (N_2709,N_1276,N_1598);
nand U2710 (N_2710,N_97,N_814);
nand U2711 (N_2711,N_2280,N_504);
and U2712 (N_2712,N_85,N_1770);
or U2713 (N_2713,N_467,N_1320);
nor U2714 (N_2714,N_2131,N_1633);
or U2715 (N_2715,N_2053,N_1513);
or U2716 (N_2716,N_1715,N_841);
or U2717 (N_2717,N_2286,N_1086);
and U2718 (N_2718,N_2424,N_120);
and U2719 (N_2719,N_248,N_423);
or U2720 (N_2720,N_1396,N_633);
nor U2721 (N_2721,N_281,N_352);
and U2722 (N_2722,N_2414,N_258);
nand U2723 (N_2723,N_2076,N_1283);
nand U2724 (N_2724,N_2052,N_1133);
or U2725 (N_2725,N_2107,N_2224);
and U2726 (N_2726,N_1920,N_1095);
or U2727 (N_2727,N_321,N_1099);
and U2728 (N_2728,N_1178,N_2038);
and U2729 (N_2729,N_301,N_635);
nor U2730 (N_2730,N_986,N_1334);
nor U2731 (N_2731,N_2432,N_961);
and U2732 (N_2732,N_1918,N_1420);
and U2733 (N_2733,N_75,N_180);
nor U2734 (N_2734,N_1772,N_2090);
or U2735 (N_2735,N_473,N_648);
or U2736 (N_2736,N_2163,N_722);
and U2737 (N_2737,N_1638,N_1309);
and U2738 (N_2738,N_2334,N_1425);
nand U2739 (N_2739,N_644,N_1591);
or U2740 (N_2740,N_959,N_2380);
or U2741 (N_2741,N_1435,N_1036);
nand U2742 (N_2742,N_1609,N_1217);
nand U2743 (N_2743,N_217,N_1602);
or U2744 (N_2744,N_887,N_1579);
and U2745 (N_2745,N_640,N_737);
nor U2746 (N_2746,N_283,N_582);
nor U2747 (N_2747,N_2168,N_1542);
nand U2748 (N_2748,N_232,N_369);
and U2749 (N_2749,N_1543,N_2475);
nor U2750 (N_2750,N_1228,N_1639);
or U2751 (N_2751,N_980,N_1703);
nand U2752 (N_2752,N_322,N_892);
or U2753 (N_2753,N_1271,N_496);
or U2754 (N_2754,N_95,N_137);
and U2755 (N_2755,N_98,N_985);
nand U2756 (N_2756,N_1780,N_22);
nand U2757 (N_2757,N_1321,N_1524);
or U2758 (N_2758,N_2354,N_1878);
nand U2759 (N_2759,N_601,N_400);
and U2760 (N_2760,N_362,N_783);
nand U2761 (N_2761,N_641,N_902);
and U2762 (N_2762,N_174,N_2024);
xnor U2763 (N_2763,N_221,N_290);
nor U2764 (N_2764,N_1427,N_599);
nand U2765 (N_2765,N_2119,N_2004);
nor U2766 (N_2766,N_356,N_2105);
nand U2767 (N_2767,N_1124,N_453);
and U2768 (N_2768,N_2373,N_825);
nand U2769 (N_2769,N_1817,N_2104);
nand U2770 (N_2770,N_970,N_318);
or U2771 (N_2771,N_1719,N_1436);
nand U2772 (N_2772,N_666,N_2023);
nor U2773 (N_2773,N_1948,N_647);
and U2774 (N_2774,N_1132,N_335);
and U2775 (N_2775,N_804,N_1910);
nand U2776 (N_2776,N_2027,N_1429);
and U2777 (N_2777,N_1128,N_677);
and U2778 (N_2778,N_2051,N_700);
nand U2779 (N_2779,N_1219,N_838);
nor U2780 (N_2780,N_1303,N_689);
or U2781 (N_2781,N_1917,N_2074);
and U2782 (N_2782,N_2466,N_61);
and U2783 (N_2783,N_390,N_2096);
and U2784 (N_2784,N_2426,N_1301);
or U2785 (N_2785,N_1470,N_9);
or U2786 (N_2786,N_2318,N_2194);
and U2787 (N_2787,N_1392,N_188);
or U2788 (N_2788,N_2304,N_1137);
nor U2789 (N_2789,N_2001,N_250);
or U2790 (N_2790,N_2033,N_2120);
nand U2791 (N_2791,N_1059,N_936);
nand U2792 (N_2792,N_212,N_1142);
nand U2793 (N_2793,N_1664,N_826);
and U2794 (N_2794,N_2013,N_2279);
nor U2795 (N_2795,N_544,N_1541);
or U2796 (N_2796,N_1546,N_2073);
and U2797 (N_2797,N_1472,N_214);
and U2798 (N_2798,N_2208,N_87);
nor U2799 (N_2799,N_458,N_923);
nand U2800 (N_2800,N_1760,N_233);
and U2801 (N_2801,N_160,N_757);
and U2802 (N_2802,N_1890,N_1694);
and U2803 (N_2803,N_646,N_1753);
nor U2804 (N_2804,N_2031,N_1489);
nand U2805 (N_2805,N_1824,N_1289);
or U2806 (N_2806,N_627,N_375);
nor U2807 (N_2807,N_2376,N_1950);
or U2808 (N_2808,N_2463,N_1379);
nand U2809 (N_2809,N_1985,N_2086);
or U2810 (N_2810,N_2297,N_915);
nand U2811 (N_2811,N_559,N_1414);
or U2812 (N_2812,N_975,N_1431);
or U2813 (N_2813,N_750,N_1826);
nor U2814 (N_2814,N_2157,N_1647);
or U2815 (N_2815,N_575,N_1316);
and U2816 (N_2816,N_1158,N_1125);
and U2817 (N_2817,N_2252,N_1477);
or U2818 (N_2818,N_2041,N_2129);
or U2819 (N_2819,N_1375,N_1866);
or U2820 (N_2820,N_385,N_429);
and U2821 (N_2821,N_304,N_2409);
nand U2822 (N_2822,N_433,N_621);
xnor U2823 (N_2823,N_795,N_779);
nor U2824 (N_2824,N_191,N_211);
and U2825 (N_2825,N_1539,N_1233);
and U2826 (N_2826,N_577,N_121);
or U2827 (N_2827,N_325,N_556);
nand U2828 (N_2828,N_10,N_1223);
nand U2829 (N_2829,N_1558,N_251);
and U2830 (N_2830,N_907,N_1701);
nand U2831 (N_2831,N_2145,N_1461);
or U2832 (N_2832,N_585,N_1349);
and U2833 (N_2833,N_1348,N_1652);
or U2834 (N_2834,N_1507,N_1411);
and U2835 (N_2835,N_1279,N_552);
nand U2836 (N_2836,N_1242,N_1084);
and U2837 (N_2837,N_1739,N_402);
or U2838 (N_2838,N_23,N_1654);
nor U2839 (N_2839,N_394,N_1661);
nand U2840 (N_2840,N_2244,N_1198);
nor U2841 (N_2841,N_1247,N_760);
nand U2842 (N_2842,N_1209,N_1081);
nor U2843 (N_2843,N_618,N_1386);
and U2844 (N_2844,N_124,N_1617);
and U2845 (N_2845,N_981,N_2311);
nand U2846 (N_2846,N_1656,N_1623);
or U2847 (N_2847,N_1590,N_852);
or U2848 (N_2848,N_2029,N_43);
and U2849 (N_2849,N_964,N_2449);
or U2850 (N_2850,N_1187,N_532);
nor U2851 (N_2851,N_2465,N_1118);
nor U2852 (N_2852,N_1987,N_688);
or U2853 (N_2853,N_2214,N_2301);
nor U2854 (N_2854,N_2170,N_2260);
nand U2855 (N_2855,N_1346,N_53);
nand U2856 (N_2856,N_1122,N_2153);
nor U2857 (N_2857,N_38,N_247);
and U2858 (N_2858,N_1576,N_1535);
nand U2859 (N_2859,N_388,N_605);
nand U2860 (N_2860,N_2370,N_514);
nand U2861 (N_2861,N_312,N_344);
nand U2862 (N_2862,N_1512,N_703);
or U2863 (N_2863,N_572,N_368);
nand U2864 (N_2864,N_1416,N_470);
or U2865 (N_2865,N_507,N_1685);
nor U2866 (N_2866,N_2471,N_1025);
nor U2867 (N_2867,N_1404,N_2226);
nand U2868 (N_2868,N_1675,N_860);
nor U2869 (N_2869,N_1515,N_921);
and U2870 (N_2870,N_167,N_494);
nand U2871 (N_2871,N_1110,N_1193);
or U2872 (N_2872,N_1191,N_196);
nand U2873 (N_2873,N_1343,N_185);
or U2874 (N_2874,N_1180,N_128);
or U2875 (N_2875,N_161,N_1997);
nor U2876 (N_2876,N_1777,N_1305);
or U2877 (N_2877,N_1468,N_2403);
and U2878 (N_2878,N_1382,N_330);
nor U2879 (N_2879,N_1234,N_1135);
nor U2880 (N_2880,N_1562,N_736);
or U2881 (N_2881,N_501,N_1445);
or U2882 (N_2882,N_1038,N_1936);
or U2883 (N_2883,N_2240,N_1401);
and U2884 (N_2884,N_1448,N_2020);
or U2885 (N_2885,N_1275,N_579);
or U2886 (N_2886,N_1916,N_337);
and U2887 (N_2887,N_2385,N_2454);
and U2888 (N_2888,N_1889,N_2390);
nand U2889 (N_2889,N_208,N_1018);
nor U2890 (N_2890,N_2216,N_55);
and U2891 (N_2891,N_1371,N_2350);
nor U2892 (N_2892,N_1563,N_576);
and U2893 (N_2893,N_1782,N_1620);
or U2894 (N_2894,N_756,N_74);
nand U2895 (N_2895,N_734,N_1138);
or U2896 (N_2896,N_1373,N_403);
or U2897 (N_2897,N_2448,N_2135);
and U2898 (N_2898,N_1793,N_178);
and U2899 (N_2899,N_2372,N_1871);
and U2900 (N_2900,N_704,N_956);
and U2901 (N_2901,N_1073,N_1676);
nand U2902 (N_2902,N_36,N_937);
and U2903 (N_2903,N_2489,N_719);
or U2904 (N_2904,N_309,N_1368);
nand U2905 (N_2905,N_1949,N_1341);
nor U2906 (N_2906,N_866,N_456);
or U2907 (N_2907,N_540,N_1258);
and U2908 (N_2908,N_620,N_718);
nor U2909 (N_2909,N_842,N_383);
and U2910 (N_2910,N_2333,N_439);
or U2911 (N_2911,N_285,N_2460);
or U2912 (N_2912,N_879,N_931);
nand U2913 (N_2913,N_698,N_1163);
or U2914 (N_2914,N_1722,N_735);
and U2915 (N_2915,N_943,N_554);
and U2916 (N_2916,N_733,N_830);
or U2917 (N_2917,N_1407,N_1554);
and U2918 (N_2918,N_1921,N_2388);
nor U2919 (N_2919,N_1152,N_1717);
or U2920 (N_2920,N_1070,N_872);
xor U2921 (N_2921,N_1575,N_2416);
and U2922 (N_2922,N_2072,N_143);
nand U2923 (N_2923,N_2397,N_969);
nand U2924 (N_2924,N_195,N_1269);
nor U2925 (N_2925,N_34,N_1398);
nand U2926 (N_2926,N_671,N_2094);
and U2927 (N_2927,N_206,N_152);
nor U2928 (N_2928,N_1236,N_1060);
or U2929 (N_2929,N_1230,N_1960);
nor U2930 (N_2930,N_1761,N_690);
nand U2931 (N_2931,N_1559,N_54);
and U2932 (N_2932,N_683,N_822);
nor U2933 (N_2933,N_1449,N_606);
nor U2934 (N_2934,N_2406,N_1779);
nor U2935 (N_2935,N_1820,N_562);
and U2936 (N_2936,N_354,N_503);
and U2937 (N_2937,N_2233,N_549);
nand U2938 (N_2938,N_331,N_1696);
and U2939 (N_2939,N_2198,N_1277);
nor U2940 (N_2940,N_993,N_968);
nand U2941 (N_2941,N_1419,N_1545);
or U2942 (N_2942,N_1465,N_1286);
nand U2943 (N_2943,N_859,N_1072);
nor U2944 (N_2944,N_1940,N_1496);
nand U2945 (N_2945,N_2339,N_2175);
and U2946 (N_2946,N_1642,N_987);
and U2947 (N_2947,N_1516,N_2060);
or U2948 (N_2948,N_829,N_347);
and U2949 (N_2949,N_2264,N_2462);
nand U2950 (N_2950,N_11,N_1644);
and U2951 (N_2951,N_865,N_1479);
xnor U2952 (N_2952,N_910,N_1778);
nor U2953 (N_2953,N_645,N_2470);
or U2954 (N_2954,N_413,N_493);
or U2955 (N_2955,N_1683,N_108);
nand U2956 (N_2956,N_164,N_1984);
nand U2957 (N_2957,N_835,N_586);
or U2958 (N_2958,N_1622,N_2025);
nor U2959 (N_2959,N_2444,N_2439);
nand U2960 (N_2960,N_1151,N_1009);
nor U2961 (N_2961,N_169,N_2126);
and U2962 (N_2962,N_2281,N_2415);
nor U2963 (N_2963,N_882,N_476);
and U2964 (N_2964,N_1204,N_2097);
nand U2965 (N_2965,N_1245,N_133);
nand U2966 (N_2966,N_1751,N_746);
or U2967 (N_2967,N_341,N_2078);
or U2968 (N_2968,N_1121,N_2442);
and U2969 (N_2969,N_2270,N_346);
nand U2970 (N_2970,N_674,N_1173);
nor U2971 (N_2971,N_2391,N_100);
nand U2972 (N_2972,N_2419,N_2166);
nor U2973 (N_2973,N_2285,N_2019);
and U2974 (N_2974,N_2014,N_1486);
and U2975 (N_2975,N_1821,N_1340);
and U2976 (N_2976,N_505,N_2177);
and U2977 (N_2977,N_1161,N_2026);
nand U2978 (N_2978,N_373,N_1238);
xor U2979 (N_2979,N_303,N_1106);
and U2980 (N_2980,N_1941,N_1827);
nand U2981 (N_2981,N_47,N_650);
nand U2982 (N_2982,N_1266,N_1016);
and U2983 (N_2983,N_2417,N_2248);
nand U2984 (N_2984,N_1801,N_2317);
and U2985 (N_2985,N_42,N_2284);
and U2986 (N_2986,N_1240,N_404);
nor U2987 (N_2987,N_1584,N_200);
or U2988 (N_2988,N_1645,N_35);
or U2989 (N_2989,N_1808,N_76);
and U2990 (N_2990,N_2282,N_954);
and U2991 (N_2991,N_2159,N_2467);
nand U2992 (N_2992,N_1533,N_1856);
nand U2993 (N_2993,N_51,N_1536);
or U2994 (N_2994,N_1058,N_386);
nand U2995 (N_2995,N_300,N_1359);
nor U2996 (N_2996,N_2330,N_1159);
nor U2997 (N_2997,N_364,N_2367);
nand U2998 (N_2998,N_617,N_2269);
and U2999 (N_2999,N_1655,N_590);
xnor U3000 (N_3000,N_1111,N_104);
nor U3001 (N_3001,N_868,N_1861);
nand U3002 (N_3002,N_2383,N_1604);
nand U3003 (N_3003,N_109,N_1030);
or U3004 (N_3004,N_1450,N_1361);
nand U3005 (N_3005,N_2127,N_2459);
nor U3006 (N_3006,N_2176,N_1254);
or U3007 (N_3007,N_765,N_781);
nor U3008 (N_3008,N_1803,N_498);
nor U3009 (N_3009,N_202,N_2200);
or U3010 (N_3010,N_971,N_2497);
or U3011 (N_3011,N_1374,N_788);
and U3012 (N_3012,N_118,N_1315);
and U3013 (N_3013,N_729,N_1928);
and U3014 (N_3014,N_435,N_2082);
nand U3015 (N_3015,N_260,N_593);
or U3016 (N_3016,N_2420,N_652);
nand U3017 (N_3017,N_1914,N_1556);
nand U3018 (N_3018,N_84,N_694);
or U3019 (N_3019,N_1805,N_2441);
nor U3020 (N_3020,N_112,N_1310);
or U3021 (N_3021,N_2392,N_1547);
nor U3022 (N_3022,N_282,N_1788);
nand U3023 (N_3023,N_670,N_3);
or U3024 (N_3024,N_992,N_2461);
or U3025 (N_3025,N_1108,N_1437);
nor U3026 (N_3026,N_440,N_5);
nor U3027 (N_3027,N_2071,N_1282);
nor U3028 (N_3028,N_2323,N_392);
and U3029 (N_3029,N_2325,N_1612);
nor U3030 (N_3030,N_630,N_266);
or U3031 (N_3031,N_918,N_676);
and U3032 (N_3032,N_1698,N_667);
and U3033 (N_3033,N_2137,N_1666);
or U3034 (N_3034,N_1210,N_333);
and U3035 (N_3035,N_622,N_1764);
and U3036 (N_3036,N_1981,N_637);
and U3037 (N_3037,N_2259,N_216);
or U3038 (N_3038,N_724,N_1735);
nand U3039 (N_3039,N_1658,N_2044);
nand U3040 (N_3040,N_495,N_2288);
or U3041 (N_3041,N_2421,N_2256);
nor U3042 (N_3042,N_2418,N_1988);
and U3043 (N_3043,N_1186,N_1443);
and U3044 (N_3044,N_767,N_1049);
or U3045 (N_3045,N_334,N_1908);
nor U3046 (N_3046,N_1713,N_1785);
xnor U3047 (N_3047,N_1179,N_903);
nor U3048 (N_3048,N_29,N_537);
or U3049 (N_3049,N_2299,N_607);
and U3050 (N_3050,N_1409,N_317);
nor U3051 (N_3051,N_1907,N_1784);
nor U3052 (N_3052,N_1679,N_996);
nor U3053 (N_3053,N_1045,N_840);
and U3054 (N_3054,N_274,N_726);
and U3055 (N_3055,N_1083,N_1263);
nand U3056 (N_3056,N_2092,N_2359);
and U3057 (N_3057,N_909,N_2116);
and U3058 (N_3058,N_994,N_2018);
nand U3059 (N_3059,N_33,N_1031);
nand U3060 (N_3060,N_148,N_1747);
nor U3061 (N_3061,N_1028,N_1410);
nand U3062 (N_3062,N_1807,N_81);
and U3063 (N_3063,N_1888,N_1749);
or U3064 (N_3064,N_1211,N_338);
nor U3065 (N_3065,N_405,N_1990);
nand U3066 (N_3066,N_2009,N_165);
and U3067 (N_3067,N_685,N_1098);
nor U3068 (N_3068,N_1605,N_833);
or U3069 (N_3069,N_1452,N_332);
nor U3070 (N_3070,N_30,N_1898);
nor U3071 (N_3071,N_1707,N_222);
nand U3072 (N_3072,N_2393,N_1300);
and U3073 (N_3073,N_901,N_1757);
and U3074 (N_3074,N_1573,N_1426);
nor U3075 (N_3075,N_2440,N_1991);
and U3076 (N_3076,N_1812,N_272);
or U3077 (N_3077,N_978,N_858);
nor U3078 (N_3078,N_721,N_631);
nand U3079 (N_3079,N_766,N_218);
and U3080 (N_3080,N_1252,N_380);
and U3081 (N_3081,N_448,N_83);
and U3082 (N_3082,N_2049,N_820);
or U3083 (N_3083,N_154,N_2488);
and U3084 (N_3084,N_1003,N_468);
nor U3085 (N_3085,N_1832,N_2369);
or U3086 (N_3086,N_1331,N_548);
or U3087 (N_3087,N_2266,N_1951);
nor U3088 (N_3088,N_948,N_461);
nor U3089 (N_3089,N_1873,N_32);
or U3090 (N_3090,N_1859,N_1206);
nor U3091 (N_3091,N_1759,N_1190);
and U3092 (N_3092,N_2059,N_1394);
nand U3093 (N_3093,N_1791,N_716);
and U3094 (N_3094,N_1653,N_96);
or U3095 (N_3095,N_1854,N_2265);
nor U3096 (N_3096,N_967,N_2185);
nor U3097 (N_3097,N_516,N_79);
and U3098 (N_3098,N_2477,N_1312);
or U3099 (N_3099,N_2261,N_1682);
xor U3100 (N_3100,N_1668,N_2196);
and U3101 (N_3101,N_2095,N_557);
or U3102 (N_3102,N_234,N_655);
or U3103 (N_3103,N_1624,N_1804);
and U3104 (N_3104,N_1322,N_511);
nand U3105 (N_3105,N_995,N_960);
or U3106 (N_3106,N_1061,N_686);
nor U3107 (N_3107,N_2000,N_1883);
or U3108 (N_3108,N_1678,N_500);
or U3109 (N_3109,N_1127,N_1288);
or U3110 (N_3110,N_488,N_2089);
nor U3111 (N_3111,N_237,N_2378);
and U3112 (N_3112,N_1446,N_1972);
nand U3113 (N_3113,N_1250,N_802);
or U3114 (N_3114,N_1466,N_2184);
or U3115 (N_3115,N_336,N_2382);
and U3116 (N_3116,N_183,N_1587);
nor U3117 (N_3117,N_1689,N_502);
or U3118 (N_3118,N_2338,N_856);
or U3119 (N_3119,N_1880,N_1298);
nand U3120 (N_3120,N_2482,N_813);
and U3121 (N_3121,N_52,N_1455);
and U3122 (N_3122,N_661,N_1930);
and U3123 (N_3123,N_2099,N_663);
or U3124 (N_3124,N_1548,N_898);
nor U3125 (N_3125,N_1996,N_546);
or U3126 (N_3126,N_2148,N_800);
nor U3127 (N_3127,N_1766,N_1202);
and U3128 (N_3128,N_668,N_1358);
nor U3129 (N_3129,N_1226,N_1899);
and U3130 (N_3130,N_6,N_982);
nand U3131 (N_3131,N_571,N_1725);
nand U3132 (N_3132,N_2469,N_1965);
nand U3133 (N_3133,N_408,N_1107);
and U3134 (N_3134,N_2101,N_2312);
nor U3135 (N_3135,N_1691,N_1756);
nand U3136 (N_3136,N_2292,N_2423);
and U3137 (N_3137,N_62,N_890);
and U3138 (N_3138,N_384,N_1284);
nor U3139 (N_3139,N_864,N_1243);
or U3140 (N_3140,N_2191,N_2431);
nor U3141 (N_3141,N_520,N_712);
nor U3142 (N_3142,N_65,N_1428);
or U3143 (N_3143,N_1197,N_1002);
nand U3144 (N_3144,N_1912,N_484);
nand U3145 (N_3145,N_1103,N_897);
nor U3146 (N_3146,N_1218,N_1686);
nand U3147 (N_3147,N_2225,N_24);
or U3148 (N_3148,N_855,N_873);
nand U3149 (N_3149,N_412,N_391);
or U3150 (N_3150,N_806,N_1964);
nor U3151 (N_3151,N_1544,N_708);
and U3152 (N_3152,N_2276,N_634);
nor U3153 (N_3153,N_1157,N_837);
and U3154 (N_3154,N_2400,N_1572);
and U3155 (N_3155,N_1063,N_2232);
nand U3156 (N_3156,N_1292,N_2239);
or U3157 (N_3157,N_497,N_1843);
or U3158 (N_3158,N_1606,N_2268);
or U3159 (N_3159,N_933,N_2165);
and U3160 (N_3160,N_1337,N_220);
nor U3161 (N_3161,N_2047,N_463);
nor U3162 (N_3162,N_2398,N_2048);
nand U3163 (N_3163,N_665,N_2012);
nand U3164 (N_3164,N_2213,N_1293);
nand U3165 (N_3165,N_365,N_2067);
and U3166 (N_3166,N_2007,N_2056);
and U3167 (N_3167,N_1352,N_466);
or U3168 (N_3168,N_1975,N_1942);
nor U3169 (N_3169,N_808,N_14);
and U3170 (N_3170,N_2410,N_238);
nand U3171 (N_3171,N_1004,N_15);
or U3172 (N_3172,N_361,N_594);
nand U3173 (N_3173,N_1958,N_482);
nand U3174 (N_3174,N_895,N_1781);
nand U3175 (N_3175,N_17,N_64);
nor U3176 (N_3176,N_1570,N_149);
and U3177 (N_3177,N_7,N_1336);
nand U3178 (N_3178,N_2472,N_2128);
nand U3179 (N_3179,N_1387,N_2139);
and U3180 (N_3180,N_1823,N_2192);
or U3181 (N_3181,N_611,N_809);
nand U3182 (N_3182,N_2042,N_596);
nor U3183 (N_3183,N_1737,N_381);
or U3184 (N_3184,N_1231,N_581);
nand U3185 (N_3185,N_973,N_68);
nor U3186 (N_3186,N_1851,N_1592);
nand U3187 (N_3187,N_2387,N_797);
nor U3188 (N_3188,N_1509,N_2227);
and U3189 (N_3189,N_1640,N_565);
and U3190 (N_3190,N_776,N_2147);
or U3191 (N_3191,N_1586,N_263);
or U3192 (N_3192,N_295,N_551);
nand U3193 (N_3193,N_755,N_1695);
nand U3194 (N_3194,N_2032,N_1705);
nand U3195 (N_3195,N_1402,N_1222);
or U3196 (N_3196,N_1852,N_273);
nor U3197 (N_3197,N_194,N_397);
and U3198 (N_3198,N_1376,N_869);
and U3199 (N_3199,N_744,N_522);
nor U3200 (N_3200,N_1201,N_1175);
nor U3201 (N_3201,N_914,N_1796);
or U3202 (N_3202,N_1797,N_1954);
or U3203 (N_3203,N_1520,N_1870);
or U3204 (N_3204,N_843,N_410);
nor U3205 (N_3205,N_754,N_1955);
and U3206 (N_3206,N_1502,N_2006);
nand U3207 (N_3207,N_1372,N_1771);
nand U3208 (N_3208,N_1119,N_934);
or U3209 (N_3209,N_430,N_906);
nor U3210 (N_3210,N_1139,N_1672);
nand U3211 (N_3211,N_236,N_134);
and U3212 (N_3212,N_0,N_1775);
or U3213 (N_3213,N_1601,N_254);
nand U3214 (N_3214,N_418,N_1798);
and U3215 (N_3215,N_771,N_1872);
and U3216 (N_3216,N_616,N_785);
nand U3217 (N_3217,N_271,N_1636);
or U3218 (N_3218,N_2115,N_1412);
or U3219 (N_3219,N_1430,N_1143);
and U3220 (N_3220,N_1493,N_2230);
and U3221 (N_3221,N_1067,N_2346);
nand U3222 (N_3222,N_475,N_86);
or U3223 (N_3223,N_223,N_949);
and U3224 (N_3224,N_1027,N_711);
and U3225 (N_3225,N_1087,N_1232);
or U3226 (N_3226,N_1064,N_1864);
nor U3227 (N_3227,N_73,N_1473);
or U3228 (N_3228,N_1763,N_1498);
and U3229 (N_3229,N_2084,N_1089);
nand U3230 (N_3230,N_2055,N_2206);
and U3231 (N_3231,N_2030,N_1799);
nor U3232 (N_3232,N_1165,N_1931);
nand U3233 (N_3233,N_1324,N_2190);
nor U3234 (N_3234,N_817,N_1711);
nand U3235 (N_3235,N_560,N_406);
nor U3236 (N_3236,N_592,N_1136);
and U3237 (N_3237,N_1116,N_1244);
nand U3238 (N_3238,N_1406,N_2054);
xnor U3239 (N_3239,N_530,N_2427);
nand U3240 (N_3240,N_215,N_917);
nor U3241 (N_3241,N_870,N_1148);
and U3242 (N_3242,N_1532,N_658);
nor U3243 (N_3243,N_566,N_1332);
nand U3244 (N_3244,N_262,N_2366);
and U3245 (N_3245,N_1935,N_2437);
nor U3246 (N_3246,N_1578,N_2207);
or U3247 (N_3247,N_930,N_1730);
or U3248 (N_3248,N_2088,N_1768);
nand U3249 (N_3249,N_1727,N_2394);
nor U3250 (N_3250,N_705,N_1943);
and U3251 (N_3251,N_2228,N_598);
or U3252 (N_3252,N_1141,N_1600);
and U3253 (N_3253,N_486,N_1306);
or U3254 (N_3254,N_1388,N_1184);
and U3255 (N_3255,N_1665,N_881);
and U3256 (N_3256,N_465,N_1953);
nand U3257 (N_3257,N_1712,N_353);
nor U3258 (N_3258,N_1196,N_16);
nor U3259 (N_3259,N_1560,N_793);
or U3260 (N_3260,N_27,N_998);
nor U3261 (N_3261,N_1933,N_1342);
nand U3262 (N_3262,N_1057,N_1460);
and U3263 (N_3263,N_2396,N_1366);
and U3264 (N_3264,N_78,N_784);
or U3265 (N_3265,N_848,N_2173);
and U3266 (N_3266,N_1172,N_88);
or U3267 (N_3267,N_358,N_201);
or U3268 (N_3268,N_529,N_1091);
nor U3269 (N_3269,N_1740,N_1052);
or U3270 (N_3270,N_1903,N_1102);
or U3271 (N_3271,N_963,N_91);
and U3272 (N_3272,N_742,N_443);
and U3273 (N_3273,N_2258,N_827);
or U3274 (N_3274,N_256,N_1583);
or U3275 (N_3275,N_1569,N_1307);
and U3276 (N_3276,N_1144,N_947);
nor U3277 (N_3277,N_1484,N_186);
or U3278 (N_3278,N_1892,N_2340);
and U3279 (N_3279,N_2008,N_2218);
nor U3280 (N_3280,N_615,N_517);
and U3281 (N_3281,N_899,N_1596);
or U3282 (N_3282,N_1463,N_265);
and U3283 (N_3283,N_983,N_2453);
nand U3284 (N_3284,N_518,N_278);
and U3285 (N_3285,N_550,N_235);
or U3286 (N_3286,N_1481,N_2085);
nor U3287 (N_3287,N_2389,N_1482);
nor U3288 (N_3288,N_2337,N_1721);
or U3289 (N_3289,N_876,N_659);
or U3290 (N_3290,N_1527,N_1626);
and U3291 (N_3291,N_1350,N_2117);
or U3292 (N_3292,N_547,N_1838);
nor U3293 (N_3293,N_138,N_155);
nand U3294 (N_3294,N_2498,N_2468);
nor U3295 (N_3295,N_1129,N_2413);
xnor U3296 (N_3296,N_639,N_764);
nor U3297 (N_3297,N_102,N_1518);
and U3298 (N_3298,N_140,N_1505);
nor U3299 (N_3299,N_1836,N_2187);
and U3300 (N_3300,N_691,N_1215);
or U3301 (N_3301,N_1304,N_610);
xor U3302 (N_3302,N_8,N_294);
nand U3303 (N_3303,N_420,N_1551);
and U3304 (N_3304,N_197,N_1741);
nand U3305 (N_3305,N_2411,N_732);
and U3306 (N_3306,N_1840,N_2203);
or U3307 (N_3307,N_1105,N_348);
and U3308 (N_3308,N_126,N_288);
or U3309 (N_3309,N_1724,N_801);
nor U3310 (N_3310,N_989,N_2081);
nand U3311 (N_3311,N_1909,N_2199);
and U3312 (N_3312,N_1610,N_1383);
nand U3313 (N_3313,N_1886,N_569);
nor U3314 (N_3314,N_1962,N_1982);
or U3315 (N_3315,N_1079,N_1235);
and U3316 (N_3316,N_2046,N_1957);
nand U3317 (N_3317,N_398,N_1628);
and U3318 (N_3318,N_432,N_1615);
or U3319 (N_3319,N_1051,N_2335);
nor U3320 (N_3320,N_1671,N_770);
nand U3321 (N_3321,N_1582,N_1203);
nor U3322 (N_3322,N_447,N_182);
and U3323 (N_3323,N_1267,N_1681);
nor U3324 (N_3324,N_747,N_46);
nor U3325 (N_3325,N_845,N_2428);
or U3326 (N_3326,N_190,N_1959);
nor U3327 (N_3327,N_1023,N_1828);
or U3328 (N_3328,N_880,N_1783);
nor U3329 (N_3329,N_1849,N_2186);
or U3330 (N_3330,N_2308,N_2150);
nor U3331 (N_3331,N_2267,N_276);
or U3332 (N_3332,N_1176,N_2352);
or U3333 (N_3333,N_157,N_1442);
and U3334 (N_3334,N_922,N_359);
and U3335 (N_3335,N_329,N_2277);
and U3336 (N_3336,N_1835,N_2102);
nand U3337 (N_3337,N_526,N_1650);
nor U3338 (N_3338,N_1728,N_2327);
and U3339 (N_3339,N_1977,N_2002);
nand U3340 (N_3340,N_1199,N_2483);
nand U3341 (N_3341,N_162,N_69);
and U3342 (N_3342,N_1794,N_243);
or U3343 (N_3343,N_1109,N_1104);
and U3344 (N_3344,N_1280,N_1397);
or U3345 (N_3345,N_2138,N_2479);
nand U3346 (N_3346,N_1938,N_199);
or U3347 (N_3347,N_834,N_1166);
or U3348 (N_3348,N_1323,N_2015);
nand U3349 (N_3349,N_1353,N_2342);
or U3350 (N_3350,N_1192,N_542);
nor U3351 (N_3351,N_417,N_421);
nor U3352 (N_3352,N_1641,N_738);
or U3353 (N_3353,N_990,N_1989);
xnor U3354 (N_3354,N_1934,N_1364);
nand U3355 (N_3355,N_1618,N_2146);
or U3356 (N_3356,N_176,N_2241);
and U3357 (N_3357,N_490,N_2154);
nor U3358 (N_3358,N_2201,N_2435);
nand U3359 (N_3359,N_1900,N_1837);
nor U3360 (N_3360,N_1625,N_1979);
or U3361 (N_3361,N_1262,N_478);
nor U3362 (N_3362,N_2246,N_114);
and U3363 (N_3363,N_105,N_2481);
nand U3364 (N_3364,N_988,N_1501);
or U3365 (N_3365,N_919,N_1748);
nand U3366 (N_3366,N_1499,N_1050);
nand U3367 (N_3367,N_136,N_1112);
nor U3368 (N_3368,N_1253,N_1174);
and U3369 (N_3369,N_1999,N_2474);
nor U3370 (N_3370,N_1214,N_240);
nand U3371 (N_3371,N_370,N_1066);
nand U3372 (N_3372,N_828,N_2399);
nor U3373 (N_3373,N_1333,N_213);
nor U3374 (N_3374,N_26,N_940);
and U3375 (N_3375,N_2412,N_2195);
or U3376 (N_3376,N_2491,N_2178);
nor U3377 (N_3377,N_2193,N_595);
nand U3378 (N_3378,N_1684,N_991);
nand U3379 (N_3379,N_1802,N_1946);
nor U3380 (N_3380,N_999,N_678);
or U3381 (N_3381,N_1568,N_1904);
and U3382 (N_3382,N_1969,N_1844);
and U3383 (N_3383,N_1395,N_1024);
or U3384 (N_3384,N_769,N_1994);
and U3385 (N_3385,N_449,N_1432);
and U3386 (N_3386,N_580,N_57);
or U3387 (N_3387,N_787,N_485);
and U3388 (N_3388,N_1514,N_296);
nand U3389 (N_3389,N_2142,N_1850);
nor U3390 (N_3390,N_1365,N_2125);
or U3391 (N_3391,N_2130,N_1867);
or U3392 (N_3392,N_762,N_2003);
nand U3393 (N_3393,N_2235,N_142);
nand U3394 (N_3394,N_812,N_715);
and U3395 (N_3395,N_145,N_2291);
and U3396 (N_3396,N_2257,N_1945);
nand U3397 (N_3397,N_2215,N_2181);
and U3398 (N_3398,N_2098,N_242);
or U3399 (N_3399,N_1581,N_1071);
and U3400 (N_3400,N_1659,N_1155);
nor U3401 (N_3401,N_555,N_1523);
nand U3402 (N_3402,N_863,N_111);
nor U3403 (N_3403,N_241,N_18);
nand U3404 (N_3404,N_1697,N_455);
nor U3405 (N_3405,N_357,N_1792);
or U3406 (N_3406,N_175,N_2293);
nand U3407 (N_3407,N_1317,N_382);
nor U3408 (N_3408,N_2404,N_2210);
or U3409 (N_3409,N_1032,N_302);
nor U3410 (N_3410,N_436,N_1865);
and U3411 (N_3411,N_1561,N_1274);
nor U3412 (N_3412,N_2341,N_972);
nor U3413 (N_3413,N_1019,N_697);
or U3414 (N_3414,N_307,N_1225);
nand U3415 (N_3415,N_2212,N_177);
nor U3416 (N_3416,N_1021,N_426);
and U3417 (N_3417,N_2010,N_1530);
nor U3418 (N_3418,N_1194,N_1281);
nor U3419 (N_3419,N_2114,N_945);
and U3420 (N_3420,N_612,N_1227);
nor U3421 (N_3421,N_1115,N_924);
nor U3422 (N_3422,N_1363,N_342);
xor U3423 (N_3423,N_127,N_1831);
nor U3424 (N_3424,N_1017,N_1216);
or U3425 (N_3425,N_2283,N_204);
nor U3426 (N_3426,N_1616,N_979);
nor U3427 (N_3427,N_1511,N_2152);
nor U3428 (N_3428,N_1046,N_1924);
nor U3429 (N_3429,N_1834,N_1525);
xor U3430 (N_3430,N_2169,N_1153);
nand U3431 (N_3431,N_1929,N_1339);
nor U3432 (N_3432,N_1205,N_1167);
and U3433 (N_3433,N_1092,N_1571);
or U3434 (N_3434,N_1896,N_2211);
and U3435 (N_3435,N_538,N_257);
or U3436 (N_3436,N_306,N_1015);
and U3437 (N_3437,N_1663,N_2377);
nor U3438 (N_3438,N_2402,N_928);
and U3439 (N_3439,N_2271,N_1731);
and U3440 (N_3440,N_299,N_2368);
and U3441 (N_3441,N_20,N_1169);
nand U3442 (N_3442,N_2433,N_1574);
or U3443 (N_3443,N_159,N_487);
nand U3444 (N_3444,N_1008,N_623);
nand U3445 (N_3445,N_298,N_944);
nor U3446 (N_3446,N_2068,N_1745);
nand U3447 (N_3447,N_1053,N_1229);
nor U3448 (N_3448,N_209,N_328);
or U3449 (N_3449,N_66,N_1926);
or U3450 (N_3450,N_1389,N_163);
or U3451 (N_3451,N_1423,N_1065);
nand U3452 (N_3452,N_173,N_378);
nand U3453 (N_3453,N_1611,N_225);
nand U3454 (N_3454,N_1040,N_45);
and U3455 (N_3455,N_2273,N_1506);
and U3456 (N_3456,N_1467,N_1007);
nor U3457 (N_3457,N_106,N_2236);
nor U3458 (N_3458,N_1433,N_2485);
and U3459 (N_3459,N_63,N_1390);
nor U3460 (N_3460,N_2161,N_1531);
nor U3461 (N_3461,N_1251,N_2021);
or U3462 (N_3462,N_1126,N_1034);
nand U3463 (N_3463,N_1391,N_2384);
nand U3464 (N_3464,N_1674,N_741);
and U3465 (N_3465,N_558,N_1010);
and U3466 (N_3466,N_636,N_786);
nor U3467 (N_3467,N_2499,N_1150);
nor U3468 (N_3468,N_1818,N_1978);
or U3469 (N_3469,N_773,N_2162);
or U3470 (N_3470,N_1259,N_1961);
and U3471 (N_3471,N_441,N_1318);
and U3472 (N_3472,N_1881,N_2093);
or U3473 (N_3473,N_355,N_56);
and U3474 (N_3474,N_1708,N_759);
nand U3475 (N_3475,N_2447,N_796);
or U3476 (N_3476,N_1752,N_1603);
nand U3477 (N_3477,N_1588,N_1422);
nor U3478 (N_3478,N_1497,N_2355);
or U3479 (N_3479,N_1966,N_1351);
nor U3480 (N_3480,N_192,N_471);
or U3481 (N_3481,N_474,N_1974);
or U3482 (N_3482,N_713,N_389);
nor U3483 (N_3483,N_1710,N_2349);
or U3484 (N_3484,N_2364,N_1848);
and U3485 (N_3485,N_1457,N_723);
or U3486 (N_3486,N_2083,N_2401);
nand U3487 (N_3487,N_1816,N_308);
or U3488 (N_3488,N_1459,N_277);
nor U3489 (N_3489,N_419,N_563);
or U3490 (N_3490,N_67,N_1795);
nand U3491 (N_3491,N_836,N_2118);
and U3492 (N_3492,N_1635,N_2316);
and U3493 (N_3493,N_231,N_727);
and U3494 (N_3494,N_1742,N_37);
nand U3495 (N_3495,N_372,N_1540);
and U3496 (N_3496,N_2361,N_1555);
or U3497 (N_3497,N_1314,N_1491);
nand U3498 (N_3498,N_2112,N_1973);
nand U3499 (N_3499,N_523,N_1521);
and U3500 (N_3500,N_512,N_1693);
or U3501 (N_3501,N_1597,N_229);
nor U3502 (N_3502,N_139,N_2141);
nor U3503 (N_3503,N_743,N_1120);
or U3504 (N_3504,N_545,N_1937);
nor U3505 (N_3505,N_553,N_1662);
nand U3506 (N_3506,N_289,N_438);
or U3507 (N_3507,N_48,N_1385);
nand U3508 (N_3508,N_1325,N_643);
nor U3509 (N_3509,N_957,N_1913);
or U3510 (N_3510,N_2478,N_2313);
nor U3511 (N_3511,N_1413,N_219);
or U3512 (N_3512,N_324,N_123);
or U3513 (N_3513,N_1670,N_1074);
nor U3514 (N_3514,N_130,N_1968);
or U3515 (N_3515,N_942,N_58);
nand U3516 (N_3516,N_1296,N_305);
xnor U3517 (N_3517,N_1168,N_350);
nand U3518 (N_3518,N_1185,N_13);
and U3519 (N_3519,N_1272,N_1754);
and U3520 (N_3520,N_1068,N_141);
nand U3521 (N_3521,N_525,N_2351);
xor U3522 (N_3522,N_2070,N_2164);
or U3523 (N_3523,N_543,N_1894);
nor U3524 (N_3524,N_2016,N_2386);
nor U3525 (N_3525,N_1700,N_2149);
or U3526 (N_3526,N_701,N_583);
nor U3527 (N_3527,N_1487,N_2061);
or U3528 (N_3528,N_396,N_2363);
or U3529 (N_3529,N_1381,N_411);
and U3530 (N_3530,N_1983,N_40);
nand U3531 (N_3531,N_323,N_2050);
and U3532 (N_3532,N_2231,N_351);
and U3533 (N_3533,N_1529,N_1447);
nand U3534 (N_3534,N_2294,N_255);
or U3535 (N_3535,N_660,N_774);
or U3536 (N_3536,N_1114,N_1417);
nor U3537 (N_3537,N_642,N_259);
and U3538 (N_3538,N_778,N_1100);
or U3539 (N_3539,N_1776,N_1875);
and U3540 (N_3540,N_1967,N_326);
nand U3541 (N_3541,N_1483,N_2160);
and U3542 (N_3542,N_1164,N_2022);
nor U3543 (N_3543,N_709,N_2229);
nor U3544 (N_3544,N_862,N_437);
nor U3545 (N_3545,N_2476,N_2234);
and U3546 (N_3546,N_239,N_1441);
or U3547 (N_3547,N_965,N_2310);
or U3548 (N_3548,N_628,N_2347);
and U3549 (N_3549,N_609,N_2155);
nand U3550 (N_3550,N_1595,N_132);
nand U3551 (N_3551,N_1882,N_270);
or U3552 (N_3552,N_2062,N_2321);
or U3553 (N_3553,N_927,N_2458);
and U3554 (N_3554,N_1723,N_1438);
nor U3555 (N_3555,N_871,N_1357);
and U3556 (N_3556,N_2043,N_2222);
nor U3557 (N_3557,N_1716,N_2151);
nor U3558 (N_3558,N_893,N_1195);
or U3559 (N_3559,N_888,N_327);
and U3560 (N_3560,N_147,N_1869);
and U3561 (N_3561,N_1773,N_1677);
and U3562 (N_3562,N_1093,N_1853);
or U3563 (N_3563,N_680,N_2295);
nand U3564 (N_3564,N_2103,N_1311);
nand U3565 (N_3565,N_2156,N_2045);
and U3566 (N_3566,N_1813,N_2017);
nor U3567 (N_3567,N_962,N_662);
nor U3568 (N_3568,N_226,N_1637);
nand U3569 (N_3569,N_684,N_1188);
or U3570 (N_3570,N_2289,N_717);
and U3571 (N_3571,N_1630,N_119);
and U3572 (N_3572,N_629,N_527);
and U3573 (N_3573,N_1687,N_1755);
and U3574 (N_3574,N_669,N_1488);
nor U3575 (N_3575,N_144,N_889);
nor U3576 (N_3576,N_1819,N_1146);
nor U3577 (N_3577,N_44,N_531);
or U3578 (N_3578,N_707,N_2091);
and U3579 (N_3579,N_1077,N_1011);
nand U3580 (N_3580,N_508,N_1055);
nor U3581 (N_3581,N_2005,N_2306);
or U3582 (N_3582,N_745,N_619);
nor U3583 (N_3583,N_1690,N_1993);
and U3584 (N_3584,N_1246,N_1069);
or U3585 (N_3585,N_524,N_230);
and U3586 (N_3586,N_1508,N_70);
nand U3587 (N_3587,N_1939,N_1354);
or U3588 (N_3588,N_1140,N_92);
or U3589 (N_3589,N_1248,N_2079);
nor U3590 (N_3590,N_1789,N_1370);
nor U3591 (N_3591,N_59,N_1995);
or U3592 (N_3592,N_2492,N_874);
xnor U3593 (N_3593,N_2451,N_1688);
and U3594 (N_3594,N_761,N_314);
nor U3595 (N_3595,N_2262,N_275);
and U3596 (N_3596,N_291,N_2446);
and U3597 (N_3597,N_1704,N_1944);
nand U3598 (N_3598,N_1594,N_122);
and U3599 (N_3599,N_1156,N_99);
and U3600 (N_3600,N_287,N_1237);
or U3601 (N_3601,N_2182,N_1825);
and U3602 (N_3602,N_819,N_1130);
nor U3603 (N_3603,N_1787,N_2278);
nor U3604 (N_3604,N_207,N_2329);
and U3605 (N_3605,N_1718,N_849);
nand U3606 (N_3606,N_1906,N_2307);
xor U3607 (N_3607,N_319,N_1669);
and U3608 (N_3608,N_1113,N_951);
or U3609 (N_3609,N_146,N_1319);
nand U3610 (N_3610,N_632,N_1504);
nor U3611 (N_3611,N_1699,N_673);
and U3612 (N_3612,N_1480,N_1651);
nor U3613 (N_3613,N_2087,N_2452);
nand U3614 (N_3614,N_1474,N_445);
and U3615 (N_3615,N_1762,N_850);
nor U3616 (N_3616,N_459,N_1149);
or U3617 (N_3617,N_913,N_1709);
nor U3618 (N_3618,N_657,N_472);
and U3619 (N_3619,N_1075,N_2362);
nor U3620 (N_3620,N_1746,N_115);
nor U3621 (N_3621,N_818,N_1743);
or U3622 (N_3622,N_1421,N_587);
nand U3623 (N_3623,N_311,N_2179);
nand U3624 (N_3624,N_2490,N_564);
or U3625 (N_3625,N_2221,N_789);
and U3626 (N_3626,N_1829,N_815);
nor U3627 (N_3627,N_1012,N_821);
nand U3628 (N_3628,N_80,N_1160);
nand U3629 (N_3629,N_205,N_2487);
nand U3630 (N_3630,N_790,N_2066);
nor U3631 (N_3631,N_1241,N_588);
or U3632 (N_3632,N_2174,N_929);
and U3633 (N_3633,N_293,N_2037);
nor U3634 (N_3634,N_316,N_1868);
nand U3635 (N_3635,N_2040,N_1085);
nor U3636 (N_3636,N_2172,N_25);
or U3637 (N_3637,N_264,N_725);
or U3638 (N_3638,N_1589,N_166);
or U3639 (N_3639,N_446,N_1434);
and U3640 (N_3640,N_2110,N_1863);
nor U3641 (N_3641,N_2209,N_1758);
or U3642 (N_3642,N_952,N_2456);
nand U3643 (N_3643,N_2434,N_415);
nand U3644 (N_3644,N_730,N_2381);
or U3645 (N_3645,N_2100,N_2255);
nor U3646 (N_3646,N_1767,N_1992);
or U3647 (N_3647,N_1786,N_1614);
or U3648 (N_3648,N_1330,N_2484);
nand U3649 (N_3649,N_2344,N_521);
and U3650 (N_3650,N_2123,N_1440);
nand U3651 (N_3651,N_1963,N_2223);
and U3652 (N_3652,N_2425,N_1806);
and U3653 (N_3653,N_1393,N_696);
and U3654 (N_3654,N_2356,N_1424);
nand U3655 (N_3655,N_1876,N_135);
or U3656 (N_3656,N_1538,N_158);
nand U3657 (N_3657,N_1212,N_2464);
nand U3658 (N_3658,N_900,N_894);
nor U3659 (N_3659,N_1200,N_1893);
or U3660 (N_3660,N_1765,N_950);
or U3661 (N_3661,N_1290,N_1607);
or U3662 (N_3662,N_857,N_399);
nand U3663 (N_3663,N_2395,N_1952);
and U3664 (N_3664,N_2455,N_479);
or U3665 (N_3665,N_1000,N_1224);
nor U3666 (N_3666,N_510,N_2343);
or U3667 (N_3667,N_1567,N_172);
and U3668 (N_3668,N_1439,N_1736);
or U3669 (N_3669,N_875,N_1255);
nand U3670 (N_3670,N_1566,N_179);
nor U3671 (N_3671,N_1291,N_491);
and U3672 (N_3672,N_807,N_758);
or U3673 (N_3673,N_1035,N_1998);
or U3674 (N_3674,N_2132,N_1285);
or U3675 (N_3675,N_2315,N_1297);
nand U3676 (N_3676,N_90,N_1020);
nor U3677 (N_3677,N_1162,N_2108);
or U3678 (N_3678,N_1033,N_653);
nor U3679 (N_3679,N_654,N_2158);
or U3680 (N_3680,N_589,N_682);
or U3681 (N_3681,N_2408,N_409);
nand U3682 (N_3682,N_693,N_624);
or U3683 (N_3683,N_2314,N_602);
nand U3684 (N_3684,N_2183,N_198);
or U3685 (N_3685,N_499,N_2405);
or U3686 (N_3686,N_584,N_2134);
and U3687 (N_3687,N_2069,N_675);
nand U3688 (N_3688,N_1599,N_535);
and U3689 (N_3689,N_1273,N_2167);
nand U3690 (N_3690,N_2332,N_2324);
nor U3691 (N_3691,N_2251,N_2365);
and U3692 (N_3692,N_1810,N_1726);
nand U3693 (N_3693,N_1884,N_2438);
nand U3694 (N_3694,N_861,N_1911);
or U3695 (N_3695,N_1308,N_2429);
nor U3696 (N_3696,N_1845,N_2298);
or U3697 (N_3697,N_984,N_878);
nand U3698 (N_3698,N_941,N_604);
or U3699 (N_3699,N_1976,N_2238);
nand U3700 (N_3700,N_1082,N_101);
nor U3701 (N_3701,N_21,N_699);
nor U3702 (N_3702,N_2253,N_82);
nand U3703 (N_3703,N_536,N_1744);
or U3704 (N_3704,N_1564,N_851);
or U3705 (N_3705,N_457,N_244);
nor U3706 (N_3706,N_534,N_1415);
nand U3707 (N_3707,N_1062,N_2486);
nor U3708 (N_3708,N_896,N_1839);
and U3709 (N_3709,N_1145,N_416);
xnor U3710 (N_3710,N_151,N_1256);
or U3711 (N_3711,N_1680,N_702);
and U3712 (N_3712,N_1042,N_1980);
nand U3713 (N_3713,N_2189,N_387);
or U3714 (N_3714,N_1362,N_2326);
or U3715 (N_3715,N_926,N_1469);
nand U3716 (N_3716,N_1855,N_2430);
and U3717 (N_3717,N_1462,N_2407);
or U3718 (N_3718,N_1213,N_1585);
nor U3719 (N_3719,N_1005,N_297);
or U3720 (N_3720,N_1842,N_803);
nor U3721 (N_3721,N_428,N_1147);
nor U3722 (N_3722,N_246,N_651);
xor U3723 (N_3723,N_710,N_1400);
nor U3724 (N_3724,N_1458,N_1478);
nor U3725 (N_3725,N_2109,N_1847);
and U3726 (N_3726,N_2035,N_477);
nand U3727 (N_3727,N_280,N_1345);
nor U3728 (N_3728,N_2028,N_451);
nor U3729 (N_3729,N_2113,N_2036);
nor U3730 (N_3730,N_1329,N_1901);
or U3731 (N_3731,N_103,N_1858);
xnor U3732 (N_3732,N_168,N_613);
or U3733 (N_3733,N_1220,N_997);
and U3734 (N_3734,N_1347,N_313);
nand U3735 (N_3735,N_2494,N_2217);
xor U3736 (N_3736,N_1927,N_1648);
nor U3737 (N_3737,N_189,N_1667);
nand U3738 (N_3738,N_920,N_932);
and U3739 (N_3739,N_2272,N_340);
nand U3740 (N_3740,N_885,N_2357);
nand U3741 (N_3741,N_1464,N_345);
or U3742 (N_3742,N_2379,N_117);
or U3743 (N_3743,N_780,N_1552);
and U3744 (N_3744,N_1456,N_2237);
nor U3745 (N_3745,N_1534,N_1326);
nand U3746 (N_3746,N_509,N_1328);
nand U3747 (N_3747,N_626,N_976);
or U3748 (N_3748,N_1860,N_1932);
nand U3749 (N_3749,N_1923,N_320);
nor U3750 (N_3750,N_448,N_2165);
or U3751 (N_3751,N_557,N_2060);
nand U3752 (N_3752,N_532,N_2321);
and U3753 (N_3753,N_238,N_2194);
nand U3754 (N_3754,N_1130,N_2109);
and U3755 (N_3755,N_61,N_1257);
nand U3756 (N_3756,N_1884,N_374);
or U3757 (N_3757,N_2300,N_347);
nand U3758 (N_3758,N_2497,N_979);
nand U3759 (N_3759,N_365,N_73);
or U3760 (N_3760,N_1742,N_464);
or U3761 (N_3761,N_2037,N_2443);
or U3762 (N_3762,N_1002,N_1352);
or U3763 (N_3763,N_669,N_2369);
nor U3764 (N_3764,N_983,N_1448);
or U3765 (N_3765,N_1493,N_2260);
or U3766 (N_3766,N_2184,N_2065);
or U3767 (N_3767,N_2273,N_1577);
or U3768 (N_3768,N_734,N_685);
or U3769 (N_3769,N_1528,N_1677);
nand U3770 (N_3770,N_2308,N_362);
or U3771 (N_3771,N_1769,N_1220);
or U3772 (N_3772,N_1812,N_2086);
nand U3773 (N_3773,N_1898,N_422);
nand U3774 (N_3774,N_789,N_1208);
nor U3775 (N_3775,N_2261,N_343);
or U3776 (N_3776,N_521,N_547);
or U3777 (N_3777,N_1077,N_1082);
nor U3778 (N_3778,N_1069,N_624);
or U3779 (N_3779,N_287,N_2309);
nor U3780 (N_3780,N_2128,N_462);
or U3781 (N_3781,N_1691,N_990);
and U3782 (N_3782,N_963,N_363);
or U3783 (N_3783,N_1403,N_1750);
or U3784 (N_3784,N_1141,N_375);
or U3785 (N_3785,N_536,N_2345);
nand U3786 (N_3786,N_745,N_369);
nand U3787 (N_3787,N_2208,N_1989);
nand U3788 (N_3788,N_1142,N_684);
or U3789 (N_3789,N_824,N_1476);
or U3790 (N_3790,N_1355,N_2365);
or U3791 (N_3791,N_2346,N_1941);
nand U3792 (N_3792,N_704,N_1204);
or U3793 (N_3793,N_133,N_2230);
nand U3794 (N_3794,N_124,N_121);
nor U3795 (N_3795,N_1907,N_2156);
and U3796 (N_3796,N_1644,N_2313);
nand U3797 (N_3797,N_1398,N_542);
nor U3798 (N_3798,N_1506,N_894);
nor U3799 (N_3799,N_6,N_1124);
nor U3800 (N_3800,N_1379,N_1696);
and U3801 (N_3801,N_1272,N_16);
and U3802 (N_3802,N_1264,N_1550);
nor U3803 (N_3803,N_882,N_904);
nand U3804 (N_3804,N_276,N_2027);
nand U3805 (N_3805,N_968,N_2479);
or U3806 (N_3806,N_967,N_499);
or U3807 (N_3807,N_284,N_851);
xor U3808 (N_3808,N_1393,N_2401);
nor U3809 (N_3809,N_1934,N_2007);
and U3810 (N_3810,N_744,N_937);
nand U3811 (N_3811,N_280,N_1671);
or U3812 (N_3812,N_2424,N_2005);
nand U3813 (N_3813,N_2221,N_8);
nor U3814 (N_3814,N_1843,N_24);
or U3815 (N_3815,N_1995,N_113);
nor U3816 (N_3816,N_548,N_2293);
nor U3817 (N_3817,N_342,N_806);
and U3818 (N_3818,N_1293,N_1042);
nor U3819 (N_3819,N_1942,N_723);
or U3820 (N_3820,N_1440,N_1389);
or U3821 (N_3821,N_805,N_619);
and U3822 (N_3822,N_401,N_1713);
nand U3823 (N_3823,N_2192,N_1255);
and U3824 (N_3824,N_2323,N_1470);
nand U3825 (N_3825,N_2014,N_2476);
and U3826 (N_3826,N_278,N_126);
or U3827 (N_3827,N_2058,N_856);
or U3828 (N_3828,N_2054,N_1611);
nand U3829 (N_3829,N_2455,N_2235);
nand U3830 (N_3830,N_613,N_2338);
and U3831 (N_3831,N_1969,N_2109);
nor U3832 (N_3832,N_1445,N_1299);
or U3833 (N_3833,N_594,N_1385);
and U3834 (N_3834,N_2275,N_1833);
nand U3835 (N_3835,N_835,N_80);
nand U3836 (N_3836,N_1829,N_2078);
nand U3837 (N_3837,N_1050,N_11);
nand U3838 (N_3838,N_271,N_888);
nor U3839 (N_3839,N_2240,N_2470);
nand U3840 (N_3840,N_1665,N_2443);
nand U3841 (N_3841,N_1343,N_1731);
nand U3842 (N_3842,N_1304,N_146);
or U3843 (N_3843,N_355,N_367);
or U3844 (N_3844,N_2135,N_1412);
nor U3845 (N_3845,N_1428,N_63);
and U3846 (N_3846,N_832,N_1826);
or U3847 (N_3847,N_74,N_399);
or U3848 (N_3848,N_2229,N_625);
nor U3849 (N_3849,N_355,N_29);
or U3850 (N_3850,N_183,N_2413);
or U3851 (N_3851,N_1119,N_2491);
nand U3852 (N_3852,N_1493,N_2134);
and U3853 (N_3853,N_2428,N_1108);
and U3854 (N_3854,N_860,N_557);
or U3855 (N_3855,N_394,N_1124);
nand U3856 (N_3856,N_177,N_1117);
nor U3857 (N_3857,N_1208,N_804);
or U3858 (N_3858,N_1228,N_2331);
nor U3859 (N_3859,N_1288,N_740);
and U3860 (N_3860,N_1982,N_785);
or U3861 (N_3861,N_497,N_2480);
nor U3862 (N_3862,N_265,N_1903);
nor U3863 (N_3863,N_1229,N_2409);
nand U3864 (N_3864,N_719,N_74);
nand U3865 (N_3865,N_2192,N_1026);
nand U3866 (N_3866,N_791,N_201);
nand U3867 (N_3867,N_2152,N_774);
and U3868 (N_3868,N_1303,N_448);
nand U3869 (N_3869,N_1880,N_1678);
nor U3870 (N_3870,N_2231,N_1111);
nor U3871 (N_3871,N_545,N_712);
nand U3872 (N_3872,N_962,N_559);
nor U3873 (N_3873,N_1575,N_646);
nor U3874 (N_3874,N_31,N_939);
nand U3875 (N_3875,N_1809,N_1759);
nand U3876 (N_3876,N_2193,N_1737);
nand U3877 (N_3877,N_1787,N_691);
and U3878 (N_3878,N_1610,N_1930);
and U3879 (N_3879,N_1877,N_2330);
and U3880 (N_3880,N_2282,N_2396);
nor U3881 (N_3881,N_2383,N_67);
nand U3882 (N_3882,N_120,N_1376);
nand U3883 (N_3883,N_498,N_2027);
and U3884 (N_3884,N_344,N_684);
and U3885 (N_3885,N_898,N_2380);
nor U3886 (N_3886,N_1852,N_2076);
nor U3887 (N_3887,N_2477,N_604);
nand U3888 (N_3888,N_1054,N_2355);
and U3889 (N_3889,N_485,N_1348);
nor U3890 (N_3890,N_475,N_947);
nor U3891 (N_3891,N_536,N_1622);
or U3892 (N_3892,N_2040,N_640);
nand U3893 (N_3893,N_1311,N_806);
or U3894 (N_3894,N_334,N_1666);
and U3895 (N_3895,N_1146,N_813);
xor U3896 (N_3896,N_225,N_2475);
nand U3897 (N_3897,N_1846,N_2424);
nand U3898 (N_3898,N_1976,N_2147);
or U3899 (N_3899,N_713,N_671);
nand U3900 (N_3900,N_866,N_581);
nor U3901 (N_3901,N_1624,N_1114);
xor U3902 (N_3902,N_1651,N_896);
nand U3903 (N_3903,N_561,N_639);
and U3904 (N_3904,N_956,N_2195);
nor U3905 (N_3905,N_22,N_1534);
or U3906 (N_3906,N_1241,N_584);
or U3907 (N_3907,N_565,N_304);
nand U3908 (N_3908,N_105,N_127);
or U3909 (N_3909,N_1318,N_101);
or U3910 (N_3910,N_1554,N_807);
nor U3911 (N_3911,N_775,N_2418);
nor U3912 (N_3912,N_1289,N_1606);
nand U3913 (N_3913,N_2038,N_271);
nand U3914 (N_3914,N_33,N_425);
xnor U3915 (N_3915,N_998,N_1547);
or U3916 (N_3916,N_1961,N_1186);
or U3917 (N_3917,N_1563,N_422);
or U3918 (N_3918,N_303,N_1462);
or U3919 (N_3919,N_1493,N_301);
and U3920 (N_3920,N_1569,N_30);
nor U3921 (N_3921,N_2474,N_270);
or U3922 (N_3922,N_1776,N_354);
nand U3923 (N_3923,N_147,N_1810);
and U3924 (N_3924,N_371,N_840);
or U3925 (N_3925,N_527,N_997);
nor U3926 (N_3926,N_1979,N_1849);
nor U3927 (N_3927,N_968,N_841);
or U3928 (N_3928,N_1276,N_2477);
and U3929 (N_3929,N_1710,N_73);
nand U3930 (N_3930,N_2168,N_1948);
nor U3931 (N_3931,N_2286,N_577);
nor U3932 (N_3932,N_854,N_950);
or U3933 (N_3933,N_1789,N_284);
nand U3934 (N_3934,N_2217,N_466);
or U3935 (N_3935,N_90,N_215);
or U3936 (N_3936,N_493,N_213);
or U3937 (N_3937,N_288,N_490);
nand U3938 (N_3938,N_1567,N_663);
or U3939 (N_3939,N_2482,N_485);
nor U3940 (N_3940,N_2086,N_2322);
nand U3941 (N_3941,N_557,N_2055);
or U3942 (N_3942,N_759,N_96);
nand U3943 (N_3943,N_2443,N_12);
or U3944 (N_3944,N_731,N_2147);
nor U3945 (N_3945,N_4,N_672);
and U3946 (N_3946,N_2029,N_865);
nand U3947 (N_3947,N_83,N_1459);
or U3948 (N_3948,N_1326,N_1828);
nand U3949 (N_3949,N_1208,N_1632);
nand U3950 (N_3950,N_832,N_1345);
and U3951 (N_3951,N_1070,N_164);
and U3952 (N_3952,N_827,N_2136);
and U3953 (N_3953,N_2434,N_1030);
and U3954 (N_3954,N_451,N_1291);
nor U3955 (N_3955,N_119,N_1712);
or U3956 (N_3956,N_21,N_1486);
nand U3957 (N_3957,N_2149,N_707);
nor U3958 (N_3958,N_1190,N_2199);
nor U3959 (N_3959,N_831,N_1288);
or U3960 (N_3960,N_2322,N_367);
and U3961 (N_3961,N_305,N_362);
nor U3962 (N_3962,N_158,N_2179);
nand U3963 (N_3963,N_966,N_2048);
nor U3964 (N_3964,N_2446,N_1894);
or U3965 (N_3965,N_2059,N_303);
or U3966 (N_3966,N_953,N_1178);
nor U3967 (N_3967,N_428,N_733);
nor U3968 (N_3968,N_2223,N_1215);
or U3969 (N_3969,N_1921,N_1133);
nor U3970 (N_3970,N_1835,N_74);
or U3971 (N_3971,N_511,N_2326);
nand U3972 (N_3972,N_1555,N_1026);
and U3973 (N_3973,N_1767,N_902);
nor U3974 (N_3974,N_1123,N_373);
and U3975 (N_3975,N_2091,N_2311);
and U3976 (N_3976,N_28,N_2389);
nand U3977 (N_3977,N_1835,N_1107);
and U3978 (N_3978,N_2472,N_1040);
and U3979 (N_3979,N_1739,N_1658);
and U3980 (N_3980,N_2069,N_1886);
and U3981 (N_3981,N_1697,N_1209);
or U3982 (N_3982,N_2367,N_2042);
xor U3983 (N_3983,N_2254,N_1878);
nand U3984 (N_3984,N_2029,N_2306);
and U3985 (N_3985,N_24,N_676);
or U3986 (N_3986,N_1448,N_1499);
and U3987 (N_3987,N_2369,N_2305);
nor U3988 (N_3988,N_1552,N_1316);
or U3989 (N_3989,N_2459,N_234);
nand U3990 (N_3990,N_211,N_1866);
and U3991 (N_3991,N_912,N_931);
or U3992 (N_3992,N_139,N_1460);
nand U3993 (N_3993,N_2073,N_26);
or U3994 (N_3994,N_181,N_1817);
nand U3995 (N_3995,N_1552,N_1450);
nand U3996 (N_3996,N_2251,N_2085);
and U3997 (N_3997,N_1978,N_1126);
nand U3998 (N_3998,N_1530,N_412);
or U3999 (N_3999,N_187,N_2151);
nor U4000 (N_4000,N_215,N_40);
and U4001 (N_4001,N_294,N_2192);
nand U4002 (N_4002,N_2148,N_1310);
or U4003 (N_4003,N_2213,N_2270);
or U4004 (N_4004,N_2471,N_1480);
or U4005 (N_4005,N_227,N_1844);
or U4006 (N_4006,N_880,N_1032);
nor U4007 (N_4007,N_1891,N_2346);
or U4008 (N_4008,N_1392,N_850);
nand U4009 (N_4009,N_1860,N_2353);
or U4010 (N_4010,N_1572,N_473);
or U4011 (N_4011,N_2207,N_834);
nor U4012 (N_4012,N_1848,N_2070);
or U4013 (N_4013,N_1227,N_1299);
or U4014 (N_4014,N_1300,N_33);
and U4015 (N_4015,N_2476,N_2274);
and U4016 (N_4016,N_2413,N_1782);
nand U4017 (N_4017,N_420,N_700);
nand U4018 (N_4018,N_1936,N_2091);
nand U4019 (N_4019,N_1119,N_119);
or U4020 (N_4020,N_152,N_736);
nand U4021 (N_4021,N_104,N_2313);
nor U4022 (N_4022,N_1583,N_655);
and U4023 (N_4023,N_189,N_2378);
nand U4024 (N_4024,N_1914,N_240);
nor U4025 (N_4025,N_1279,N_1427);
nand U4026 (N_4026,N_833,N_1451);
or U4027 (N_4027,N_2071,N_408);
or U4028 (N_4028,N_629,N_2101);
nand U4029 (N_4029,N_464,N_2041);
or U4030 (N_4030,N_229,N_362);
or U4031 (N_4031,N_2254,N_358);
and U4032 (N_4032,N_1567,N_1400);
nand U4033 (N_4033,N_219,N_1068);
or U4034 (N_4034,N_1801,N_2446);
and U4035 (N_4035,N_826,N_972);
and U4036 (N_4036,N_957,N_1501);
or U4037 (N_4037,N_502,N_903);
and U4038 (N_4038,N_2439,N_2197);
nand U4039 (N_4039,N_634,N_1559);
nor U4040 (N_4040,N_1748,N_1637);
or U4041 (N_4041,N_542,N_1187);
and U4042 (N_4042,N_2080,N_2318);
and U4043 (N_4043,N_1485,N_1708);
or U4044 (N_4044,N_1240,N_387);
nor U4045 (N_4045,N_2248,N_1353);
nor U4046 (N_4046,N_566,N_585);
nand U4047 (N_4047,N_675,N_334);
or U4048 (N_4048,N_1195,N_1951);
and U4049 (N_4049,N_709,N_1236);
nand U4050 (N_4050,N_1528,N_1458);
nor U4051 (N_4051,N_2196,N_2295);
or U4052 (N_4052,N_875,N_1840);
nand U4053 (N_4053,N_1132,N_1977);
nor U4054 (N_4054,N_2254,N_1083);
and U4055 (N_4055,N_2472,N_1295);
nor U4056 (N_4056,N_1693,N_1592);
nand U4057 (N_4057,N_1773,N_2044);
nor U4058 (N_4058,N_1663,N_1691);
nand U4059 (N_4059,N_2230,N_61);
or U4060 (N_4060,N_500,N_1971);
nor U4061 (N_4061,N_1064,N_2060);
or U4062 (N_4062,N_114,N_1467);
nor U4063 (N_4063,N_1663,N_771);
and U4064 (N_4064,N_379,N_1905);
nand U4065 (N_4065,N_652,N_1221);
nor U4066 (N_4066,N_1473,N_1472);
or U4067 (N_4067,N_70,N_2376);
or U4068 (N_4068,N_1282,N_963);
nand U4069 (N_4069,N_1024,N_1124);
or U4070 (N_4070,N_1819,N_516);
nor U4071 (N_4071,N_2482,N_875);
or U4072 (N_4072,N_348,N_2260);
nor U4073 (N_4073,N_1176,N_39);
or U4074 (N_4074,N_2300,N_786);
nand U4075 (N_4075,N_1362,N_773);
or U4076 (N_4076,N_1818,N_1035);
or U4077 (N_4077,N_2041,N_527);
or U4078 (N_4078,N_1522,N_607);
xnor U4079 (N_4079,N_537,N_479);
nand U4080 (N_4080,N_2455,N_701);
or U4081 (N_4081,N_951,N_138);
nor U4082 (N_4082,N_1392,N_995);
xor U4083 (N_4083,N_353,N_1484);
and U4084 (N_4084,N_732,N_820);
and U4085 (N_4085,N_352,N_1305);
and U4086 (N_4086,N_1993,N_1426);
or U4087 (N_4087,N_239,N_1742);
or U4088 (N_4088,N_449,N_1981);
or U4089 (N_4089,N_250,N_965);
and U4090 (N_4090,N_2491,N_2045);
nor U4091 (N_4091,N_1876,N_99);
or U4092 (N_4092,N_1419,N_2001);
nand U4093 (N_4093,N_1333,N_1927);
or U4094 (N_4094,N_996,N_367);
or U4095 (N_4095,N_68,N_1617);
and U4096 (N_4096,N_1690,N_234);
nand U4097 (N_4097,N_824,N_1606);
nor U4098 (N_4098,N_1545,N_670);
and U4099 (N_4099,N_2017,N_237);
nand U4100 (N_4100,N_2102,N_75);
nand U4101 (N_4101,N_1385,N_785);
or U4102 (N_4102,N_1227,N_757);
and U4103 (N_4103,N_1414,N_1950);
nor U4104 (N_4104,N_15,N_1696);
nor U4105 (N_4105,N_1047,N_2275);
and U4106 (N_4106,N_194,N_1769);
nor U4107 (N_4107,N_1651,N_2085);
nor U4108 (N_4108,N_1922,N_410);
nand U4109 (N_4109,N_1048,N_725);
nand U4110 (N_4110,N_714,N_1561);
or U4111 (N_4111,N_1114,N_1301);
nor U4112 (N_4112,N_232,N_687);
and U4113 (N_4113,N_1787,N_367);
or U4114 (N_4114,N_1382,N_1618);
nor U4115 (N_4115,N_1611,N_778);
nand U4116 (N_4116,N_904,N_57);
nor U4117 (N_4117,N_1451,N_2340);
and U4118 (N_4118,N_1602,N_1771);
or U4119 (N_4119,N_842,N_2125);
and U4120 (N_4120,N_731,N_495);
nor U4121 (N_4121,N_256,N_1499);
nand U4122 (N_4122,N_1736,N_2384);
nor U4123 (N_4123,N_2486,N_1319);
nand U4124 (N_4124,N_2268,N_2479);
and U4125 (N_4125,N_203,N_253);
or U4126 (N_4126,N_2268,N_380);
and U4127 (N_4127,N_2002,N_762);
nor U4128 (N_4128,N_426,N_294);
nor U4129 (N_4129,N_2358,N_1208);
and U4130 (N_4130,N_579,N_391);
nor U4131 (N_4131,N_1786,N_2367);
nand U4132 (N_4132,N_1844,N_2090);
and U4133 (N_4133,N_1464,N_804);
and U4134 (N_4134,N_1136,N_1022);
nor U4135 (N_4135,N_2346,N_162);
nand U4136 (N_4136,N_411,N_6);
and U4137 (N_4137,N_2423,N_252);
nand U4138 (N_4138,N_448,N_1720);
or U4139 (N_4139,N_568,N_2011);
nand U4140 (N_4140,N_2319,N_334);
nand U4141 (N_4141,N_1083,N_1177);
and U4142 (N_4142,N_361,N_1246);
and U4143 (N_4143,N_337,N_1252);
nor U4144 (N_4144,N_2452,N_1724);
or U4145 (N_4145,N_675,N_1433);
and U4146 (N_4146,N_1683,N_1191);
nand U4147 (N_4147,N_1320,N_80);
nand U4148 (N_4148,N_646,N_57);
and U4149 (N_4149,N_2370,N_1547);
and U4150 (N_4150,N_1079,N_1828);
nor U4151 (N_4151,N_1432,N_2458);
nor U4152 (N_4152,N_1286,N_954);
nor U4153 (N_4153,N_2452,N_2489);
and U4154 (N_4154,N_1635,N_1554);
and U4155 (N_4155,N_1116,N_1375);
and U4156 (N_4156,N_1763,N_2233);
or U4157 (N_4157,N_1377,N_378);
nand U4158 (N_4158,N_1041,N_518);
nand U4159 (N_4159,N_1700,N_1064);
and U4160 (N_4160,N_1330,N_188);
or U4161 (N_4161,N_1361,N_929);
nand U4162 (N_4162,N_1609,N_2329);
nor U4163 (N_4163,N_1980,N_1249);
or U4164 (N_4164,N_542,N_2105);
and U4165 (N_4165,N_2331,N_2283);
and U4166 (N_4166,N_2123,N_1343);
nand U4167 (N_4167,N_395,N_1958);
and U4168 (N_4168,N_1447,N_2192);
and U4169 (N_4169,N_1676,N_70);
nor U4170 (N_4170,N_1281,N_849);
and U4171 (N_4171,N_912,N_685);
nand U4172 (N_4172,N_2440,N_1196);
nor U4173 (N_4173,N_2191,N_1152);
and U4174 (N_4174,N_2094,N_844);
and U4175 (N_4175,N_1485,N_461);
nor U4176 (N_4176,N_915,N_829);
or U4177 (N_4177,N_1106,N_1152);
nand U4178 (N_4178,N_199,N_1177);
nand U4179 (N_4179,N_276,N_652);
nand U4180 (N_4180,N_1037,N_1860);
and U4181 (N_4181,N_255,N_235);
or U4182 (N_4182,N_625,N_2324);
and U4183 (N_4183,N_193,N_424);
and U4184 (N_4184,N_527,N_1788);
and U4185 (N_4185,N_764,N_785);
nor U4186 (N_4186,N_1721,N_1569);
nor U4187 (N_4187,N_466,N_1329);
nor U4188 (N_4188,N_1701,N_1611);
and U4189 (N_4189,N_1954,N_2474);
nand U4190 (N_4190,N_727,N_19);
nor U4191 (N_4191,N_2151,N_283);
nand U4192 (N_4192,N_1838,N_1587);
and U4193 (N_4193,N_1235,N_1702);
nand U4194 (N_4194,N_893,N_791);
and U4195 (N_4195,N_1741,N_941);
nor U4196 (N_4196,N_729,N_800);
nor U4197 (N_4197,N_2120,N_1925);
nor U4198 (N_4198,N_477,N_1094);
or U4199 (N_4199,N_2258,N_300);
and U4200 (N_4200,N_439,N_1602);
and U4201 (N_4201,N_322,N_789);
and U4202 (N_4202,N_1209,N_2474);
nand U4203 (N_4203,N_975,N_1486);
and U4204 (N_4204,N_877,N_2438);
and U4205 (N_4205,N_367,N_465);
nand U4206 (N_4206,N_1804,N_2430);
or U4207 (N_4207,N_949,N_1142);
and U4208 (N_4208,N_1118,N_1218);
nor U4209 (N_4209,N_1816,N_2355);
and U4210 (N_4210,N_948,N_656);
nor U4211 (N_4211,N_2371,N_2261);
or U4212 (N_4212,N_570,N_2121);
and U4213 (N_4213,N_901,N_945);
nor U4214 (N_4214,N_1123,N_1769);
xor U4215 (N_4215,N_2061,N_721);
and U4216 (N_4216,N_2032,N_582);
nand U4217 (N_4217,N_1053,N_2373);
or U4218 (N_4218,N_1314,N_2180);
nand U4219 (N_4219,N_60,N_533);
nand U4220 (N_4220,N_861,N_2398);
and U4221 (N_4221,N_1467,N_866);
nand U4222 (N_4222,N_2096,N_2412);
nand U4223 (N_4223,N_1282,N_1562);
nor U4224 (N_4224,N_2267,N_531);
or U4225 (N_4225,N_417,N_2383);
nor U4226 (N_4226,N_537,N_2123);
nor U4227 (N_4227,N_2208,N_975);
nor U4228 (N_4228,N_1234,N_703);
or U4229 (N_4229,N_1592,N_2028);
and U4230 (N_4230,N_2466,N_1910);
and U4231 (N_4231,N_2453,N_1603);
nand U4232 (N_4232,N_177,N_2091);
or U4233 (N_4233,N_2235,N_656);
nor U4234 (N_4234,N_2082,N_2364);
or U4235 (N_4235,N_329,N_1044);
and U4236 (N_4236,N_376,N_1542);
or U4237 (N_4237,N_2144,N_33);
nor U4238 (N_4238,N_1750,N_1273);
and U4239 (N_4239,N_1416,N_383);
and U4240 (N_4240,N_957,N_871);
nor U4241 (N_4241,N_889,N_308);
nor U4242 (N_4242,N_1973,N_810);
or U4243 (N_4243,N_1868,N_711);
and U4244 (N_4244,N_2156,N_1330);
or U4245 (N_4245,N_823,N_1700);
or U4246 (N_4246,N_292,N_2190);
or U4247 (N_4247,N_845,N_8);
nor U4248 (N_4248,N_2070,N_1637);
nor U4249 (N_4249,N_1863,N_362);
or U4250 (N_4250,N_585,N_468);
nor U4251 (N_4251,N_475,N_1636);
or U4252 (N_4252,N_145,N_416);
nor U4253 (N_4253,N_1055,N_752);
nand U4254 (N_4254,N_2125,N_1180);
or U4255 (N_4255,N_573,N_942);
nand U4256 (N_4256,N_2372,N_1020);
and U4257 (N_4257,N_500,N_1954);
nor U4258 (N_4258,N_27,N_1387);
or U4259 (N_4259,N_814,N_803);
or U4260 (N_4260,N_932,N_1728);
nor U4261 (N_4261,N_2293,N_2383);
or U4262 (N_4262,N_1632,N_2448);
nand U4263 (N_4263,N_400,N_2394);
nor U4264 (N_4264,N_1385,N_215);
or U4265 (N_4265,N_640,N_2176);
nor U4266 (N_4266,N_1444,N_411);
nand U4267 (N_4267,N_458,N_1704);
and U4268 (N_4268,N_327,N_73);
or U4269 (N_4269,N_2492,N_144);
nor U4270 (N_4270,N_2331,N_2207);
nor U4271 (N_4271,N_2119,N_1008);
nand U4272 (N_4272,N_1749,N_324);
nand U4273 (N_4273,N_473,N_1895);
and U4274 (N_4274,N_2426,N_708);
nor U4275 (N_4275,N_391,N_1923);
nor U4276 (N_4276,N_2391,N_43);
and U4277 (N_4277,N_407,N_934);
nand U4278 (N_4278,N_475,N_1966);
nand U4279 (N_4279,N_2241,N_1388);
and U4280 (N_4280,N_658,N_226);
xnor U4281 (N_4281,N_372,N_90);
nand U4282 (N_4282,N_1307,N_1115);
or U4283 (N_4283,N_62,N_2236);
and U4284 (N_4284,N_2401,N_1929);
or U4285 (N_4285,N_2470,N_1098);
nand U4286 (N_4286,N_2145,N_2470);
nand U4287 (N_4287,N_730,N_2286);
nor U4288 (N_4288,N_1614,N_165);
and U4289 (N_4289,N_989,N_2113);
and U4290 (N_4290,N_2047,N_525);
or U4291 (N_4291,N_1290,N_2251);
or U4292 (N_4292,N_868,N_609);
and U4293 (N_4293,N_1781,N_594);
and U4294 (N_4294,N_1891,N_1635);
and U4295 (N_4295,N_241,N_254);
nand U4296 (N_4296,N_1037,N_1290);
and U4297 (N_4297,N_1717,N_829);
or U4298 (N_4298,N_1591,N_1736);
or U4299 (N_4299,N_1918,N_1281);
nand U4300 (N_4300,N_841,N_212);
and U4301 (N_4301,N_1761,N_2352);
nand U4302 (N_4302,N_12,N_1937);
and U4303 (N_4303,N_452,N_812);
nand U4304 (N_4304,N_884,N_585);
or U4305 (N_4305,N_1685,N_535);
nand U4306 (N_4306,N_1145,N_1265);
and U4307 (N_4307,N_11,N_2077);
and U4308 (N_4308,N_2220,N_1829);
nor U4309 (N_4309,N_1356,N_609);
and U4310 (N_4310,N_135,N_731);
nand U4311 (N_4311,N_1311,N_522);
nand U4312 (N_4312,N_1382,N_1577);
nand U4313 (N_4313,N_689,N_1187);
nor U4314 (N_4314,N_2385,N_1512);
nor U4315 (N_4315,N_263,N_2450);
or U4316 (N_4316,N_1433,N_1712);
and U4317 (N_4317,N_1729,N_719);
nand U4318 (N_4318,N_1666,N_2436);
and U4319 (N_4319,N_1500,N_317);
or U4320 (N_4320,N_2020,N_128);
nand U4321 (N_4321,N_2081,N_1590);
and U4322 (N_4322,N_1363,N_2079);
or U4323 (N_4323,N_2315,N_1551);
or U4324 (N_4324,N_2388,N_2231);
nand U4325 (N_4325,N_2119,N_1617);
nor U4326 (N_4326,N_2179,N_2379);
and U4327 (N_4327,N_153,N_157);
or U4328 (N_4328,N_555,N_258);
and U4329 (N_4329,N_1597,N_287);
nor U4330 (N_4330,N_1582,N_2378);
nand U4331 (N_4331,N_2033,N_2026);
and U4332 (N_4332,N_2406,N_825);
or U4333 (N_4333,N_1253,N_2433);
or U4334 (N_4334,N_455,N_1886);
nor U4335 (N_4335,N_1314,N_266);
nor U4336 (N_4336,N_13,N_1509);
nor U4337 (N_4337,N_263,N_1964);
and U4338 (N_4338,N_655,N_1105);
nor U4339 (N_4339,N_902,N_1491);
nor U4340 (N_4340,N_827,N_1110);
nand U4341 (N_4341,N_2479,N_1149);
or U4342 (N_4342,N_1203,N_2358);
nor U4343 (N_4343,N_611,N_132);
and U4344 (N_4344,N_1185,N_1793);
nand U4345 (N_4345,N_1457,N_679);
nor U4346 (N_4346,N_291,N_830);
or U4347 (N_4347,N_394,N_1399);
or U4348 (N_4348,N_517,N_1256);
nor U4349 (N_4349,N_2340,N_1572);
or U4350 (N_4350,N_1561,N_698);
or U4351 (N_4351,N_40,N_2209);
and U4352 (N_4352,N_277,N_547);
xor U4353 (N_4353,N_2397,N_182);
nand U4354 (N_4354,N_1223,N_2291);
and U4355 (N_4355,N_2224,N_956);
or U4356 (N_4356,N_1724,N_379);
nor U4357 (N_4357,N_2324,N_919);
nand U4358 (N_4358,N_689,N_986);
and U4359 (N_4359,N_2238,N_931);
nor U4360 (N_4360,N_2101,N_899);
or U4361 (N_4361,N_1866,N_911);
nand U4362 (N_4362,N_1892,N_359);
and U4363 (N_4363,N_1729,N_437);
or U4364 (N_4364,N_745,N_189);
nand U4365 (N_4365,N_431,N_1438);
or U4366 (N_4366,N_699,N_568);
and U4367 (N_4367,N_1171,N_1767);
nand U4368 (N_4368,N_1004,N_2288);
nor U4369 (N_4369,N_499,N_175);
nor U4370 (N_4370,N_2142,N_2249);
and U4371 (N_4371,N_1037,N_2434);
or U4372 (N_4372,N_2177,N_2236);
and U4373 (N_4373,N_554,N_2296);
or U4374 (N_4374,N_2191,N_445);
nand U4375 (N_4375,N_1336,N_1144);
nand U4376 (N_4376,N_1808,N_397);
or U4377 (N_4377,N_220,N_2100);
and U4378 (N_4378,N_1409,N_1793);
or U4379 (N_4379,N_1143,N_2474);
nor U4380 (N_4380,N_1562,N_1164);
or U4381 (N_4381,N_596,N_1837);
or U4382 (N_4382,N_1617,N_1124);
or U4383 (N_4383,N_2319,N_1080);
or U4384 (N_4384,N_1745,N_2387);
and U4385 (N_4385,N_687,N_740);
and U4386 (N_4386,N_2070,N_923);
or U4387 (N_4387,N_581,N_2120);
or U4388 (N_4388,N_1048,N_42);
nand U4389 (N_4389,N_1098,N_223);
nand U4390 (N_4390,N_1382,N_2207);
or U4391 (N_4391,N_1205,N_1451);
nor U4392 (N_4392,N_1302,N_1081);
or U4393 (N_4393,N_2180,N_1773);
and U4394 (N_4394,N_1778,N_1295);
and U4395 (N_4395,N_1270,N_583);
or U4396 (N_4396,N_380,N_629);
or U4397 (N_4397,N_296,N_2112);
or U4398 (N_4398,N_2074,N_410);
nand U4399 (N_4399,N_575,N_167);
and U4400 (N_4400,N_720,N_1023);
nor U4401 (N_4401,N_2240,N_139);
nand U4402 (N_4402,N_735,N_323);
or U4403 (N_4403,N_1805,N_183);
nand U4404 (N_4404,N_1926,N_1972);
nand U4405 (N_4405,N_1483,N_723);
or U4406 (N_4406,N_759,N_2021);
nand U4407 (N_4407,N_2234,N_757);
nand U4408 (N_4408,N_149,N_1809);
and U4409 (N_4409,N_449,N_593);
nand U4410 (N_4410,N_1476,N_2453);
nand U4411 (N_4411,N_695,N_2377);
and U4412 (N_4412,N_1596,N_1404);
nand U4413 (N_4413,N_1408,N_2389);
or U4414 (N_4414,N_884,N_1766);
and U4415 (N_4415,N_1957,N_425);
nor U4416 (N_4416,N_378,N_1095);
nand U4417 (N_4417,N_176,N_936);
or U4418 (N_4418,N_2437,N_1893);
nand U4419 (N_4419,N_1244,N_696);
nand U4420 (N_4420,N_1989,N_2004);
and U4421 (N_4421,N_2223,N_2472);
nor U4422 (N_4422,N_812,N_353);
nand U4423 (N_4423,N_1241,N_1979);
nor U4424 (N_4424,N_201,N_1791);
nor U4425 (N_4425,N_2444,N_718);
or U4426 (N_4426,N_1929,N_1277);
nor U4427 (N_4427,N_383,N_447);
or U4428 (N_4428,N_169,N_1527);
nand U4429 (N_4429,N_1816,N_479);
or U4430 (N_4430,N_1026,N_2215);
nand U4431 (N_4431,N_1885,N_744);
nand U4432 (N_4432,N_2025,N_1437);
or U4433 (N_4433,N_745,N_849);
nor U4434 (N_4434,N_1081,N_737);
nand U4435 (N_4435,N_1013,N_1921);
or U4436 (N_4436,N_2422,N_117);
or U4437 (N_4437,N_1429,N_781);
and U4438 (N_4438,N_2417,N_605);
nor U4439 (N_4439,N_1067,N_622);
or U4440 (N_4440,N_1082,N_692);
nor U4441 (N_4441,N_1412,N_2128);
nand U4442 (N_4442,N_2318,N_1679);
or U4443 (N_4443,N_1789,N_2315);
and U4444 (N_4444,N_988,N_204);
or U4445 (N_4445,N_1238,N_2243);
and U4446 (N_4446,N_1281,N_1121);
nand U4447 (N_4447,N_1282,N_651);
xnor U4448 (N_4448,N_631,N_1999);
or U4449 (N_4449,N_2398,N_1789);
nor U4450 (N_4450,N_541,N_67);
nor U4451 (N_4451,N_1944,N_1856);
nor U4452 (N_4452,N_1518,N_2236);
and U4453 (N_4453,N_528,N_1080);
or U4454 (N_4454,N_1233,N_1417);
nand U4455 (N_4455,N_1232,N_518);
nor U4456 (N_4456,N_1370,N_536);
nand U4457 (N_4457,N_497,N_851);
nand U4458 (N_4458,N_2370,N_1590);
and U4459 (N_4459,N_727,N_1874);
nand U4460 (N_4460,N_1183,N_721);
or U4461 (N_4461,N_632,N_233);
nor U4462 (N_4462,N_1802,N_1327);
or U4463 (N_4463,N_2431,N_2487);
nand U4464 (N_4464,N_2464,N_901);
nand U4465 (N_4465,N_2384,N_2446);
nand U4466 (N_4466,N_2309,N_2482);
or U4467 (N_4467,N_972,N_1757);
nor U4468 (N_4468,N_1043,N_1027);
nor U4469 (N_4469,N_1559,N_2088);
or U4470 (N_4470,N_1232,N_1194);
and U4471 (N_4471,N_980,N_161);
nor U4472 (N_4472,N_2376,N_1435);
and U4473 (N_4473,N_726,N_148);
and U4474 (N_4474,N_477,N_1934);
and U4475 (N_4475,N_1517,N_1162);
and U4476 (N_4476,N_536,N_448);
nor U4477 (N_4477,N_940,N_268);
nand U4478 (N_4478,N_1773,N_1823);
and U4479 (N_4479,N_1822,N_286);
nand U4480 (N_4480,N_775,N_2347);
nor U4481 (N_4481,N_1675,N_696);
nand U4482 (N_4482,N_2157,N_1341);
nor U4483 (N_4483,N_1510,N_42);
nor U4484 (N_4484,N_2154,N_1861);
nand U4485 (N_4485,N_28,N_1392);
or U4486 (N_4486,N_1320,N_396);
and U4487 (N_4487,N_2449,N_2129);
or U4488 (N_4488,N_2287,N_175);
nand U4489 (N_4489,N_1611,N_2081);
and U4490 (N_4490,N_2104,N_429);
nand U4491 (N_4491,N_2087,N_544);
nor U4492 (N_4492,N_71,N_1756);
or U4493 (N_4493,N_225,N_1342);
and U4494 (N_4494,N_1714,N_1503);
or U4495 (N_4495,N_2044,N_968);
nand U4496 (N_4496,N_1386,N_729);
nor U4497 (N_4497,N_753,N_2274);
and U4498 (N_4498,N_110,N_1057);
xnor U4499 (N_4499,N_1814,N_398);
nand U4500 (N_4500,N_1921,N_179);
nor U4501 (N_4501,N_704,N_1382);
or U4502 (N_4502,N_1182,N_1067);
nor U4503 (N_4503,N_746,N_1015);
nand U4504 (N_4504,N_2086,N_1571);
and U4505 (N_4505,N_2271,N_2222);
nand U4506 (N_4506,N_1179,N_247);
or U4507 (N_4507,N_95,N_1188);
nor U4508 (N_4508,N_1568,N_2403);
nand U4509 (N_4509,N_1742,N_1566);
and U4510 (N_4510,N_1517,N_505);
nor U4511 (N_4511,N_291,N_588);
and U4512 (N_4512,N_816,N_1847);
nor U4513 (N_4513,N_608,N_657);
and U4514 (N_4514,N_1507,N_1111);
nand U4515 (N_4515,N_694,N_520);
nand U4516 (N_4516,N_1720,N_167);
nor U4517 (N_4517,N_1511,N_1040);
or U4518 (N_4518,N_1540,N_1504);
or U4519 (N_4519,N_2448,N_2187);
nand U4520 (N_4520,N_329,N_961);
or U4521 (N_4521,N_910,N_2161);
nand U4522 (N_4522,N_1855,N_2228);
nor U4523 (N_4523,N_111,N_1792);
nor U4524 (N_4524,N_2359,N_2426);
nor U4525 (N_4525,N_2290,N_226);
and U4526 (N_4526,N_417,N_1640);
nor U4527 (N_4527,N_902,N_360);
and U4528 (N_4528,N_273,N_521);
nor U4529 (N_4529,N_906,N_1716);
nand U4530 (N_4530,N_1284,N_640);
and U4531 (N_4531,N_1480,N_2070);
or U4532 (N_4532,N_1346,N_1953);
or U4533 (N_4533,N_142,N_1156);
or U4534 (N_4534,N_1445,N_2373);
and U4535 (N_4535,N_2010,N_2368);
xnor U4536 (N_4536,N_2277,N_1767);
nor U4537 (N_4537,N_190,N_1278);
nand U4538 (N_4538,N_2188,N_31);
or U4539 (N_4539,N_392,N_1702);
and U4540 (N_4540,N_2125,N_1400);
and U4541 (N_4541,N_1591,N_1671);
nor U4542 (N_4542,N_2101,N_865);
or U4543 (N_4543,N_1596,N_380);
and U4544 (N_4544,N_1087,N_980);
xnor U4545 (N_4545,N_226,N_1894);
nand U4546 (N_4546,N_2311,N_234);
or U4547 (N_4547,N_711,N_490);
nor U4548 (N_4548,N_1094,N_823);
and U4549 (N_4549,N_333,N_1431);
nand U4550 (N_4550,N_376,N_108);
nor U4551 (N_4551,N_416,N_1020);
nand U4552 (N_4552,N_618,N_1609);
nand U4553 (N_4553,N_76,N_326);
or U4554 (N_4554,N_1898,N_309);
and U4555 (N_4555,N_142,N_318);
and U4556 (N_4556,N_1835,N_548);
and U4557 (N_4557,N_390,N_1414);
and U4558 (N_4558,N_128,N_1506);
or U4559 (N_4559,N_1671,N_1313);
and U4560 (N_4560,N_1594,N_2139);
or U4561 (N_4561,N_1934,N_2269);
nand U4562 (N_4562,N_1559,N_881);
or U4563 (N_4563,N_921,N_1169);
nand U4564 (N_4564,N_1891,N_2349);
or U4565 (N_4565,N_451,N_648);
or U4566 (N_4566,N_882,N_2034);
or U4567 (N_4567,N_670,N_1301);
nor U4568 (N_4568,N_2385,N_2125);
and U4569 (N_4569,N_1637,N_1370);
and U4570 (N_4570,N_1449,N_1140);
nand U4571 (N_4571,N_924,N_340);
nor U4572 (N_4572,N_1719,N_322);
and U4573 (N_4573,N_305,N_1561);
and U4574 (N_4574,N_1888,N_85);
nor U4575 (N_4575,N_1702,N_114);
nand U4576 (N_4576,N_369,N_2315);
and U4577 (N_4577,N_1186,N_992);
nand U4578 (N_4578,N_1582,N_2451);
nor U4579 (N_4579,N_2135,N_787);
nor U4580 (N_4580,N_2307,N_2103);
and U4581 (N_4581,N_2477,N_2347);
or U4582 (N_4582,N_1956,N_110);
nand U4583 (N_4583,N_2219,N_1617);
and U4584 (N_4584,N_973,N_221);
and U4585 (N_4585,N_136,N_1452);
and U4586 (N_4586,N_306,N_714);
nand U4587 (N_4587,N_1126,N_1589);
and U4588 (N_4588,N_809,N_2250);
nand U4589 (N_4589,N_1740,N_305);
nor U4590 (N_4590,N_1101,N_1145);
nor U4591 (N_4591,N_1142,N_785);
and U4592 (N_4592,N_236,N_2434);
and U4593 (N_4593,N_2258,N_1480);
nor U4594 (N_4594,N_1098,N_468);
or U4595 (N_4595,N_1403,N_1996);
nor U4596 (N_4596,N_2075,N_2191);
or U4597 (N_4597,N_1885,N_2429);
and U4598 (N_4598,N_241,N_2131);
and U4599 (N_4599,N_1319,N_1349);
or U4600 (N_4600,N_1547,N_1448);
nand U4601 (N_4601,N_2256,N_761);
and U4602 (N_4602,N_672,N_535);
or U4603 (N_4603,N_191,N_662);
or U4604 (N_4604,N_391,N_996);
or U4605 (N_4605,N_1179,N_2237);
and U4606 (N_4606,N_1277,N_1750);
nor U4607 (N_4607,N_403,N_702);
nor U4608 (N_4608,N_1576,N_1355);
nor U4609 (N_4609,N_210,N_305);
nor U4610 (N_4610,N_703,N_1291);
or U4611 (N_4611,N_1001,N_2361);
nor U4612 (N_4612,N_1883,N_147);
nand U4613 (N_4613,N_509,N_749);
or U4614 (N_4614,N_1230,N_624);
nand U4615 (N_4615,N_2413,N_795);
or U4616 (N_4616,N_1950,N_395);
nor U4617 (N_4617,N_1163,N_2341);
nand U4618 (N_4618,N_2246,N_1947);
and U4619 (N_4619,N_2483,N_588);
nor U4620 (N_4620,N_541,N_2345);
and U4621 (N_4621,N_2032,N_457);
nand U4622 (N_4622,N_733,N_2142);
nand U4623 (N_4623,N_382,N_1436);
nor U4624 (N_4624,N_1757,N_1092);
or U4625 (N_4625,N_1268,N_1385);
nor U4626 (N_4626,N_563,N_2424);
nand U4627 (N_4627,N_989,N_740);
nor U4628 (N_4628,N_1417,N_868);
nand U4629 (N_4629,N_1600,N_478);
or U4630 (N_4630,N_1786,N_1116);
nand U4631 (N_4631,N_1910,N_1009);
and U4632 (N_4632,N_1087,N_1797);
or U4633 (N_4633,N_1585,N_112);
nand U4634 (N_4634,N_236,N_123);
and U4635 (N_4635,N_1766,N_1658);
and U4636 (N_4636,N_805,N_51);
or U4637 (N_4637,N_1903,N_638);
nor U4638 (N_4638,N_394,N_583);
nor U4639 (N_4639,N_1783,N_2275);
or U4640 (N_4640,N_192,N_99);
and U4641 (N_4641,N_1777,N_505);
and U4642 (N_4642,N_616,N_697);
nand U4643 (N_4643,N_982,N_613);
and U4644 (N_4644,N_396,N_918);
and U4645 (N_4645,N_245,N_434);
nand U4646 (N_4646,N_331,N_414);
nand U4647 (N_4647,N_446,N_2153);
nand U4648 (N_4648,N_167,N_2057);
nand U4649 (N_4649,N_62,N_93);
or U4650 (N_4650,N_1736,N_1599);
nand U4651 (N_4651,N_66,N_450);
nand U4652 (N_4652,N_1379,N_1760);
or U4653 (N_4653,N_2020,N_1032);
nor U4654 (N_4654,N_2332,N_1566);
or U4655 (N_4655,N_2276,N_764);
nand U4656 (N_4656,N_2053,N_816);
and U4657 (N_4657,N_575,N_2169);
and U4658 (N_4658,N_2435,N_1539);
or U4659 (N_4659,N_2384,N_570);
nor U4660 (N_4660,N_611,N_407);
or U4661 (N_4661,N_1239,N_819);
nand U4662 (N_4662,N_846,N_576);
or U4663 (N_4663,N_1324,N_144);
and U4664 (N_4664,N_357,N_582);
and U4665 (N_4665,N_405,N_1270);
nor U4666 (N_4666,N_1521,N_2143);
and U4667 (N_4667,N_2100,N_1572);
nand U4668 (N_4668,N_2197,N_62);
nor U4669 (N_4669,N_1260,N_306);
or U4670 (N_4670,N_1763,N_1053);
or U4671 (N_4671,N_277,N_66);
nor U4672 (N_4672,N_951,N_1083);
and U4673 (N_4673,N_2277,N_746);
nand U4674 (N_4674,N_103,N_778);
or U4675 (N_4675,N_2090,N_161);
or U4676 (N_4676,N_967,N_260);
and U4677 (N_4677,N_204,N_2005);
nor U4678 (N_4678,N_580,N_1879);
or U4679 (N_4679,N_412,N_122);
nand U4680 (N_4680,N_68,N_726);
and U4681 (N_4681,N_1324,N_834);
nor U4682 (N_4682,N_986,N_988);
and U4683 (N_4683,N_1341,N_500);
and U4684 (N_4684,N_403,N_248);
nand U4685 (N_4685,N_1161,N_1489);
nand U4686 (N_4686,N_820,N_2485);
or U4687 (N_4687,N_2049,N_2221);
nor U4688 (N_4688,N_2222,N_1885);
nor U4689 (N_4689,N_2254,N_1381);
nor U4690 (N_4690,N_2280,N_485);
or U4691 (N_4691,N_2208,N_2198);
nand U4692 (N_4692,N_1218,N_236);
or U4693 (N_4693,N_2169,N_390);
xnor U4694 (N_4694,N_898,N_2134);
or U4695 (N_4695,N_1655,N_1918);
or U4696 (N_4696,N_1309,N_662);
nand U4697 (N_4697,N_1106,N_449);
or U4698 (N_4698,N_725,N_1558);
or U4699 (N_4699,N_2429,N_2249);
nand U4700 (N_4700,N_2185,N_1935);
and U4701 (N_4701,N_301,N_1039);
nor U4702 (N_4702,N_1029,N_1961);
nor U4703 (N_4703,N_891,N_1435);
and U4704 (N_4704,N_265,N_2148);
and U4705 (N_4705,N_648,N_1097);
and U4706 (N_4706,N_376,N_2036);
nand U4707 (N_4707,N_911,N_2052);
nand U4708 (N_4708,N_1062,N_753);
nand U4709 (N_4709,N_317,N_1097);
nor U4710 (N_4710,N_725,N_1553);
and U4711 (N_4711,N_1618,N_154);
or U4712 (N_4712,N_955,N_1398);
and U4713 (N_4713,N_2097,N_2178);
nor U4714 (N_4714,N_2121,N_1717);
and U4715 (N_4715,N_1496,N_1611);
nand U4716 (N_4716,N_1417,N_1651);
or U4717 (N_4717,N_640,N_799);
nor U4718 (N_4718,N_1185,N_1041);
nor U4719 (N_4719,N_260,N_563);
nand U4720 (N_4720,N_1858,N_1092);
nand U4721 (N_4721,N_1872,N_247);
nor U4722 (N_4722,N_635,N_1184);
and U4723 (N_4723,N_961,N_1050);
nor U4724 (N_4724,N_800,N_2326);
or U4725 (N_4725,N_29,N_387);
nor U4726 (N_4726,N_2127,N_593);
nor U4727 (N_4727,N_1166,N_1895);
nand U4728 (N_4728,N_1640,N_2137);
or U4729 (N_4729,N_829,N_2233);
or U4730 (N_4730,N_1567,N_924);
nor U4731 (N_4731,N_2313,N_2222);
and U4732 (N_4732,N_472,N_2323);
and U4733 (N_4733,N_2337,N_1556);
and U4734 (N_4734,N_2052,N_62);
nand U4735 (N_4735,N_1676,N_1537);
nand U4736 (N_4736,N_870,N_323);
nor U4737 (N_4737,N_987,N_1121);
or U4738 (N_4738,N_450,N_583);
and U4739 (N_4739,N_413,N_216);
or U4740 (N_4740,N_1786,N_1464);
nand U4741 (N_4741,N_1936,N_1811);
nor U4742 (N_4742,N_1691,N_1067);
nor U4743 (N_4743,N_1572,N_36);
nand U4744 (N_4744,N_1664,N_850);
nand U4745 (N_4745,N_1689,N_755);
nand U4746 (N_4746,N_1754,N_761);
nand U4747 (N_4747,N_2124,N_1485);
nor U4748 (N_4748,N_2347,N_637);
or U4749 (N_4749,N_563,N_309);
and U4750 (N_4750,N_1858,N_62);
and U4751 (N_4751,N_526,N_846);
or U4752 (N_4752,N_669,N_244);
or U4753 (N_4753,N_2440,N_665);
or U4754 (N_4754,N_2092,N_859);
and U4755 (N_4755,N_1349,N_2258);
nand U4756 (N_4756,N_1430,N_933);
or U4757 (N_4757,N_465,N_523);
and U4758 (N_4758,N_154,N_1675);
nor U4759 (N_4759,N_792,N_1457);
and U4760 (N_4760,N_192,N_2442);
nor U4761 (N_4761,N_1233,N_689);
and U4762 (N_4762,N_301,N_2373);
nand U4763 (N_4763,N_2134,N_2198);
nand U4764 (N_4764,N_627,N_311);
and U4765 (N_4765,N_530,N_1065);
nand U4766 (N_4766,N_1301,N_1964);
or U4767 (N_4767,N_1723,N_1668);
and U4768 (N_4768,N_656,N_1124);
and U4769 (N_4769,N_798,N_491);
and U4770 (N_4770,N_2361,N_2276);
nand U4771 (N_4771,N_2410,N_647);
nand U4772 (N_4772,N_1974,N_625);
and U4773 (N_4773,N_1219,N_186);
and U4774 (N_4774,N_1403,N_691);
and U4775 (N_4775,N_2286,N_1602);
and U4776 (N_4776,N_2192,N_113);
nand U4777 (N_4777,N_820,N_2206);
or U4778 (N_4778,N_2239,N_429);
or U4779 (N_4779,N_644,N_1994);
nand U4780 (N_4780,N_877,N_1245);
and U4781 (N_4781,N_2192,N_626);
and U4782 (N_4782,N_1998,N_1476);
or U4783 (N_4783,N_1002,N_221);
nand U4784 (N_4784,N_2025,N_530);
or U4785 (N_4785,N_1847,N_578);
or U4786 (N_4786,N_256,N_1946);
nand U4787 (N_4787,N_805,N_645);
nand U4788 (N_4788,N_1181,N_834);
and U4789 (N_4789,N_726,N_2155);
nor U4790 (N_4790,N_362,N_731);
nor U4791 (N_4791,N_1637,N_1430);
or U4792 (N_4792,N_749,N_1932);
or U4793 (N_4793,N_1439,N_137);
and U4794 (N_4794,N_504,N_611);
and U4795 (N_4795,N_2084,N_2403);
and U4796 (N_4796,N_1073,N_1099);
nor U4797 (N_4797,N_270,N_1198);
nor U4798 (N_4798,N_67,N_582);
and U4799 (N_4799,N_1066,N_1974);
or U4800 (N_4800,N_1261,N_1089);
nand U4801 (N_4801,N_586,N_39);
nand U4802 (N_4802,N_216,N_2159);
nand U4803 (N_4803,N_373,N_973);
nor U4804 (N_4804,N_187,N_1809);
nand U4805 (N_4805,N_1600,N_2247);
and U4806 (N_4806,N_516,N_262);
and U4807 (N_4807,N_821,N_1929);
nand U4808 (N_4808,N_2248,N_1649);
or U4809 (N_4809,N_992,N_284);
xnor U4810 (N_4810,N_1539,N_1921);
nor U4811 (N_4811,N_1450,N_64);
and U4812 (N_4812,N_1041,N_2402);
nor U4813 (N_4813,N_5,N_1494);
xnor U4814 (N_4814,N_196,N_923);
and U4815 (N_4815,N_2416,N_965);
or U4816 (N_4816,N_1084,N_1728);
and U4817 (N_4817,N_1457,N_2411);
nand U4818 (N_4818,N_252,N_809);
nor U4819 (N_4819,N_955,N_843);
and U4820 (N_4820,N_1019,N_1741);
and U4821 (N_4821,N_1769,N_1594);
and U4822 (N_4822,N_158,N_442);
or U4823 (N_4823,N_316,N_815);
and U4824 (N_4824,N_364,N_953);
xor U4825 (N_4825,N_691,N_175);
or U4826 (N_4826,N_545,N_814);
nand U4827 (N_4827,N_779,N_819);
and U4828 (N_4828,N_1073,N_671);
nor U4829 (N_4829,N_1149,N_922);
and U4830 (N_4830,N_863,N_510);
nor U4831 (N_4831,N_2069,N_2096);
nand U4832 (N_4832,N_1494,N_1052);
nor U4833 (N_4833,N_1119,N_889);
and U4834 (N_4834,N_2287,N_2107);
nor U4835 (N_4835,N_873,N_1328);
or U4836 (N_4836,N_2038,N_2323);
and U4837 (N_4837,N_2431,N_242);
nor U4838 (N_4838,N_2226,N_112);
nand U4839 (N_4839,N_1093,N_1274);
nand U4840 (N_4840,N_2484,N_2490);
and U4841 (N_4841,N_1961,N_1534);
nor U4842 (N_4842,N_2390,N_793);
nand U4843 (N_4843,N_924,N_2077);
and U4844 (N_4844,N_1564,N_761);
nor U4845 (N_4845,N_1437,N_1627);
and U4846 (N_4846,N_890,N_1233);
and U4847 (N_4847,N_2183,N_449);
nand U4848 (N_4848,N_2424,N_1340);
nand U4849 (N_4849,N_628,N_1216);
and U4850 (N_4850,N_657,N_771);
or U4851 (N_4851,N_833,N_1299);
nand U4852 (N_4852,N_2332,N_1620);
nor U4853 (N_4853,N_774,N_1091);
nand U4854 (N_4854,N_836,N_21);
or U4855 (N_4855,N_114,N_1637);
nor U4856 (N_4856,N_706,N_1987);
and U4857 (N_4857,N_2314,N_684);
nand U4858 (N_4858,N_1393,N_234);
or U4859 (N_4859,N_2391,N_868);
nor U4860 (N_4860,N_1849,N_982);
nand U4861 (N_4861,N_1321,N_1600);
nor U4862 (N_4862,N_1643,N_827);
xnor U4863 (N_4863,N_1642,N_1628);
and U4864 (N_4864,N_760,N_882);
or U4865 (N_4865,N_155,N_588);
or U4866 (N_4866,N_831,N_86);
nor U4867 (N_4867,N_1135,N_916);
nand U4868 (N_4868,N_1175,N_800);
nor U4869 (N_4869,N_2416,N_1012);
nand U4870 (N_4870,N_1961,N_1366);
and U4871 (N_4871,N_871,N_2381);
and U4872 (N_4872,N_855,N_1242);
nand U4873 (N_4873,N_1702,N_837);
nand U4874 (N_4874,N_2043,N_1197);
and U4875 (N_4875,N_612,N_340);
nor U4876 (N_4876,N_1936,N_687);
nor U4877 (N_4877,N_1478,N_1110);
or U4878 (N_4878,N_778,N_1407);
nand U4879 (N_4879,N_1622,N_1211);
and U4880 (N_4880,N_1561,N_1389);
and U4881 (N_4881,N_774,N_1531);
and U4882 (N_4882,N_126,N_1917);
or U4883 (N_4883,N_41,N_1535);
nand U4884 (N_4884,N_2437,N_985);
or U4885 (N_4885,N_618,N_1223);
and U4886 (N_4886,N_1956,N_1868);
nand U4887 (N_4887,N_2040,N_529);
and U4888 (N_4888,N_678,N_319);
nor U4889 (N_4889,N_566,N_1597);
or U4890 (N_4890,N_2475,N_809);
and U4891 (N_4891,N_1185,N_2391);
or U4892 (N_4892,N_1055,N_574);
nor U4893 (N_4893,N_727,N_2452);
or U4894 (N_4894,N_1609,N_545);
nor U4895 (N_4895,N_1975,N_123);
or U4896 (N_4896,N_1495,N_1898);
nor U4897 (N_4897,N_557,N_922);
nor U4898 (N_4898,N_383,N_338);
and U4899 (N_4899,N_1169,N_1699);
or U4900 (N_4900,N_594,N_70);
or U4901 (N_4901,N_85,N_1867);
nand U4902 (N_4902,N_403,N_2111);
xor U4903 (N_4903,N_2344,N_2272);
xor U4904 (N_4904,N_1875,N_1394);
nand U4905 (N_4905,N_1845,N_824);
or U4906 (N_4906,N_2431,N_2437);
nor U4907 (N_4907,N_2442,N_1355);
nand U4908 (N_4908,N_31,N_1239);
nor U4909 (N_4909,N_421,N_1827);
nand U4910 (N_4910,N_1923,N_1506);
or U4911 (N_4911,N_1382,N_907);
and U4912 (N_4912,N_1759,N_2198);
or U4913 (N_4913,N_2446,N_1582);
or U4914 (N_4914,N_1022,N_1045);
nor U4915 (N_4915,N_1990,N_2387);
nor U4916 (N_4916,N_1679,N_753);
and U4917 (N_4917,N_1067,N_389);
nor U4918 (N_4918,N_2385,N_1657);
or U4919 (N_4919,N_2477,N_1143);
and U4920 (N_4920,N_1575,N_1665);
nor U4921 (N_4921,N_2440,N_587);
nor U4922 (N_4922,N_763,N_115);
nand U4923 (N_4923,N_1396,N_1817);
nor U4924 (N_4924,N_1270,N_105);
nor U4925 (N_4925,N_2078,N_515);
and U4926 (N_4926,N_1072,N_880);
nand U4927 (N_4927,N_2412,N_1921);
nor U4928 (N_4928,N_2334,N_1807);
nor U4929 (N_4929,N_923,N_2066);
nand U4930 (N_4930,N_2080,N_414);
or U4931 (N_4931,N_329,N_848);
nand U4932 (N_4932,N_2310,N_1684);
nor U4933 (N_4933,N_691,N_1659);
or U4934 (N_4934,N_2068,N_2144);
or U4935 (N_4935,N_2170,N_2094);
or U4936 (N_4936,N_1835,N_1690);
or U4937 (N_4937,N_2407,N_1512);
nor U4938 (N_4938,N_262,N_1919);
nor U4939 (N_4939,N_2173,N_318);
or U4940 (N_4940,N_1209,N_2150);
nor U4941 (N_4941,N_725,N_2195);
nand U4942 (N_4942,N_1848,N_1553);
nor U4943 (N_4943,N_1919,N_444);
nor U4944 (N_4944,N_1920,N_1938);
or U4945 (N_4945,N_1095,N_1489);
and U4946 (N_4946,N_1986,N_2036);
or U4947 (N_4947,N_2240,N_1786);
and U4948 (N_4948,N_1836,N_1106);
nand U4949 (N_4949,N_377,N_98);
or U4950 (N_4950,N_1962,N_855);
nand U4951 (N_4951,N_1355,N_2257);
or U4952 (N_4952,N_1467,N_1727);
or U4953 (N_4953,N_704,N_1833);
and U4954 (N_4954,N_602,N_388);
and U4955 (N_4955,N_471,N_325);
nor U4956 (N_4956,N_738,N_823);
nand U4957 (N_4957,N_1655,N_2050);
and U4958 (N_4958,N_2480,N_600);
nor U4959 (N_4959,N_273,N_837);
or U4960 (N_4960,N_437,N_1226);
nand U4961 (N_4961,N_2392,N_118);
nor U4962 (N_4962,N_69,N_297);
and U4963 (N_4963,N_1778,N_1578);
and U4964 (N_4964,N_499,N_2245);
or U4965 (N_4965,N_2236,N_1682);
or U4966 (N_4966,N_62,N_1807);
nor U4967 (N_4967,N_1127,N_1094);
or U4968 (N_4968,N_1338,N_1328);
or U4969 (N_4969,N_1515,N_761);
or U4970 (N_4970,N_1260,N_67);
nand U4971 (N_4971,N_2277,N_1238);
or U4972 (N_4972,N_62,N_2231);
nand U4973 (N_4973,N_320,N_1639);
and U4974 (N_4974,N_800,N_1680);
and U4975 (N_4975,N_2273,N_1152);
nand U4976 (N_4976,N_155,N_1182);
xor U4977 (N_4977,N_2267,N_979);
and U4978 (N_4978,N_1345,N_1672);
or U4979 (N_4979,N_1520,N_837);
and U4980 (N_4980,N_1303,N_114);
and U4981 (N_4981,N_1898,N_2438);
nor U4982 (N_4982,N_1422,N_178);
and U4983 (N_4983,N_2471,N_2380);
nor U4984 (N_4984,N_494,N_421);
and U4985 (N_4985,N_1415,N_1079);
nand U4986 (N_4986,N_99,N_1059);
nand U4987 (N_4987,N_1029,N_2141);
nor U4988 (N_4988,N_1247,N_1810);
xor U4989 (N_4989,N_2336,N_872);
nor U4990 (N_4990,N_2482,N_1941);
nor U4991 (N_4991,N_1812,N_228);
and U4992 (N_4992,N_1363,N_1202);
nand U4993 (N_4993,N_483,N_1314);
nand U4994 (N_4994,N_2426,N_899);
and U4995 (N_4995,N_1102,N_2348);
nand U4996 (N_4996,N_1381,N_1300);
nor U4997 (N_4997,N_1511,N_1541);
and U4998 (N_4998,N_199,N_675);
and U4999 (N_4999,N_1057,N_2018);
nor UO_0 (O_0,N_4690,N_3769);
nor UO_1 (O_1,N_4712,N_4928);
nand UO_2 (O_2,N_4348,N_3212);
nand UO_3 (O_3,N_4732,N_4402);
or UO_4 (O_4,N_2508,N_4340);
nand UO_5 (O_5,N_4659,N_2808);
nor UO_6 (O_6,N_3318,N_2871);
nand UO_7 (O_7,N_2844,N_2633);
nand UO_8 (O_8,N_2732,N_4370);
and UO_9 (O_9,N_4567,N_2989);
and UO_10 (O_10,N_4893,N_4691);
nor UO_11 (O_11,N_3019,N_2765);
nor UO_12 (O_12,N_3799,N_2706);
and UO_13 (O_13,N_4999,N_3966);
nor UO_14 (O_14,N_2964,N_3855);
or UO_15 (O_15,N_4098,N_2978);
nor UO_16 (O_16,N_3305,N_2850);
or UO_17 (O_17,N_2742,N_3638);
nand UO_18 (O_18,N_3824,N_4713);
and UO_19 (O_19,N_3599,N_3249);
nor UO_20 (O_20,N_4739,N_3467);
nor UO_21 (O_21,N_3494,N_4667);
and UO_22 (O_22,N_2879,N_3395);
and UO_23 (O_23,N_2501,N_3053);
or UO_24 (O_24,N_4510,N_4064);
or UO_25 (O_25,N_3846,N_3798);
nand UO_26 (O_26,N_2699,N_3487);
nor UO_27 (O_27,N_2786,N_4094);
nand UO_28 (O_28,N_4469,N_3687);
nor UO_29 (O_29,N_4794,N_3690);
nor UO_30 (O_30,N_2954,N_2719);
and UO_31 (O_31,N_4562,N_4455);
or UO_32 (O_32,N_2855,N_2817);
and UO_33 (O_33,N_2635,N_2652);
nor UO_34 (O_34,N_4109,N_4220);
and UO_35 (O_35,N_3807,N_2833);
nor UO_36 (O_36,N_4163,N_3738);
and UO_37 (O_37,N_3332,N_3059);
nand UO_38 (O_38,N_2840,N_4486);
nor UO_39 (O_39,N_4049,N_3534);
or UO_40 (O_40,N_3347,N_4188);
nor UO_41 (O_41,N_4701,N_4547);
nor UO_42 (O_42,N_4347,N_2774);
nor UO_43 (O_43,N_3772,N_3554);
and UO_44 (O_44,N_2576,N_4496);
nor UO_45 (O_45,N_4842,N_3463);
nor UO_46 (O_46,N_3673,N_2957);
or UO_47 (O_47,N_2962,N_2554);
nand UO_48 (O_48,N_4624,N_3154);
nor UO_49 (O_49,N_3958,N_3258);
or UO_50 (O_50,N_3221,N_3765);
nor UO_51 (O_51,N_4670,N_2863);
and UO_52 (O_52,N_2516,N_4377);
or UO_53 (O_53,N_2838,N_3450);
or UO_54 (O_54,N_4056,N_4020);
nor UO_55 (O_55,N_2926,N_2991);
nor UO_56 (O_56,N_3723,N_4143);
nand UO_57 (O_57,N_2794,N_4762);
nor UO_58 (O_58,N_2728,N_3119);
nand UO_59 (O_59,N_3976,N_4409);
and UO_60 (O_60,N_3269,N_4640);
and UO_61 (O_61,N_3166,N_3036);
nor UO_62 (O_62,N_3674,N_3663);
nor UO_63 (O_63,N_4040,N_4844);
and UO_64 (O_64,N_3439,N_3861);
nand UO_65 (O_65,N_4723,N_3833);
nor UO_66 (O_66,N_4108,N_2853);
nand UO_67 (O_67,N_3652,N_3618);
nor UO_68 (O_68,N_3391,N_4758);
and UO_69 (O_69,N_4751,N_4008);
and UO_70 (O_70,N_3142,N_3571);
or UO_71 (O_71,N_3804,N_4556);
or UO_72 (O_72,N_3390,N_3196);
xnor UO_73 (O_73,N_3288,N_3177);
or UO_74 (O_74,N_3522,N_3107);
nor UO_75 (O_75,N_4018,N_4502);
nand UO_76 (O_76,N_2866,N_4993);
and UO_77 (O_77,N_3883,N_3076);
nand UO_78 (O_78,N_3333,N_3864);
nor UO_79 (O_79,N_2569,N_3942);
or UO_80 (O_80,N_2650,N_3289);
and UO_81 (O_81,N_3295,N_2709);
nor UO_82 (O_82,N_3473,N_4428);
and UO_83 (O_83,N_4544,N_4116);
and UO_84 (O_84,N_3884,N_3290);
and UO_85 (O_85,N_2660,N_2686);
or UO_86 (O_86,N_4619,N_2724);
and UO_87 (O_87,N_4782,N_3831);
and UO_88 (O_88,N_3983,N_3388);
and UO_89 (O_89,N_3348,N_4838);
nor UO_90 (O_90,N_4628,N_3486);
nor UO_91 (O_91,N_3546,N_3968);
or UO_92 (O_92,N_4171,N_3014);
nand UO_93 (O_93,N_3424,N_4442);
nand UO_94 (O_94,N_4664,N_4871);
and UO_95 (O_95,N_3714,N_4197);
or UO_96 (O_96,N_2615,N_4903);
nand UO_97 (O_97,N_4776,N_4973);
nand UO_98 (O_98,N_3617,N_4090);
nand UO_99 (O_99,N_4289,N_4692);
nor UO_100 (O_100,N_2935,N_4021);
or UO_101 (O_101,N_4048,N_3823);
or UO_102 (O_102,N_3342,N_3383);
nor UO_103 (O_103,N_4650,N_2929);
nand UO_104 (O_104,N_3033,N_4990);
or UO_105 (O_105,N_3256,N_4648);
or UO_106 (O_106,N_4954,N_2718);
nand UO_107 (O_107,N_4219,N_2856);
nor UO_108 (O_108,N_3647,N_3178);
nand UO_109 (O_109,N_4523,N_4300);
nand UO_110 (O_110,N_4777,N_3443);
nand UO_111 (O_111,N_3327,N_3123);
nor UO_112 (O_112,N_4706,N_2893);
or UO_113 (O_113,N_4229,N_4119);
nor UO_114 (O_114,N_4334,N_4298);
nand UO_115 (O_115,N_4448,N_3294);
or UO_116 (O_116,N_2619,N_4870);
or UO_117 (O_117,N_4521,N_2521);
or UO_118 (O_118,N_3078,N_3842);
nand UO_119 (O_119,N_2874,N_2625);
nand UO_120 (O_120,N_4584,N_2581);
or UO_121 (O_121,N_4798,N_4078);
nand UO_122 (O_122,N_3149,N_4506);
nand UO_123 (O_123,N_4590,N_3124);
nand UO_124 (O_124,N_4508,N_4050);
or UO_125 (O_125,N_3713,N_2636);
or UO_126 (O_126,N_4390,N_3959);
nor UO_127 (O_127,N_3620,N_4528);
nor UO_128 (O_128,N_4345,N_2781);
and UO_129 (O_129,N_2892,N_3259);
xor UO_130 (O_130,N_4073,N_3488);
nor UO_131 (O_131,N_3746,N_3199);
nand UO_132 (O_132,N_3649,N_3200);
nor UO_133 (O_133,N_3152,N_4376);
nor UO_134 (O_134,N_4814,N_3146);
nor UO_135 (O_135,N_3964,N_3670);
or UO_136 (O_136,N_3574,N_4482);
nand UO_137 (O_137,N_2744,N_4208);
and UO_138 (O_138,N_4287,N_4791);
nand UO_139 (O_139,N_3129,N_3207);
nor UO_140 (O_140,N_3403,N_2750);
and UO_141 (O_141,N_4047,N_2571);
and UO_142 (O_142,N_3496,N_3161);
nand UO_143 (O_143,N_4308,N_4186);
nand UO_144 (O_144,N_2762,N_3882);
and UO_145 (O_145,N_2661,N_4961);
and UO_146 (O_146,N_4872,N_2927);
or UO_147 (O_147,N_2587,N_3410);
or UO_148 (O_148,N_2955,N_3264);
or UO_149 (O_149,N_4470,N_3678);
nor UO_150 (O_150,N_3817,N_4773);
and UO_151 (O_151,N_3876,N_3988);
or UO_152 (O_152,N_3570,N_4265);
nor UO_153 (O_153,N_4459,N_3900);
nand UO_154 (O_154,N_3860,N_4077);
or UO_155 (O_155,N_4183,N_3064);
or UO_156 (O_156,N_4212,N_4467);
or UO_157 (O_157,N_4909,N_4918);
or UO_158 (O_158,N_3009,N_4350);
and UO_159 (O_159,N_3011,N_3500);
nand UO_160 (O_160,N_3965,N_2813);
nor UO_161 (O_161,N_4446,N_3321);
and UO_162 (O_162,N_3062,N_4525);
nor UO_163 (O_163,N_2561,N_4392);
nand UO_164 (O_164,N_3858,N_3362);
nor UO_165 (O_165,N_3818,N_2537);
xor UO_166 (O_166,N_3072,N_4859);
and UO_167 (O_167,N_2784,N_3479);
and UO_168 (O_168,N_2981,N_2685);
and UO_169 (O_169,N_3979,N_3734);
and UO_170 (O_170,N_4672,N_4210);
nor UO_171 (O_171,N_2647,N_3067);
nor UO_172 (O_172,N_4614,N_2723);
or UO_173 (O_173,N_4400,N_3625);
and UO_174 (O_174,N_3668,N_3850);
xnor UO_175 (O_175,N_3733,N_3685);
nand UO_176 (O_176,N_3543,N_2766);
nor UO_177 (O_177,N_3797,N_4393);
nand UO_178 (O_178,N_3776,N_3029);
and UO_179 (O_179,N_3157,N_3913);
or UO_180 (O_180,N_4103,N_3065);
nor UO_181 (O_181,N_3524,N_4820);
nor UO_182 (O_182,N_3634,N_3632);
and UO_183 (O_183,N_4834,N_4000);
nor UO_184 (O_184,N_4427,N_3667);
or UO_185 (O_185,N_3548,N_2726);
nor UO_186 (O_186,N_2645,N_3120);
nor UO_187 (O_187,N_2529,N_3512);
or UO_188 (O_188,N_4187,N_3012);
nand UO_189 (O_189,N_3749,N_4034);
and UO_190 (O_190,N_3285,N_4126);
or UO_191 (O_191,N_4687,N_4771);
or UO_192 (O_192,N_2642,N_4721);
nand UO_193 (O_193,N_3969,N_3266);
and UO_194 (O_194,N_4071,N_2500);
nand UO_195 (O_195,N_3896,N_3729);
nor UO_196 (O_196,N_3313,N_3429);
and UO_197 (O_197,N_4611,N_3897);
nand UO_198 (O_198,N_3084,N_4967);
nor UO_199 (O_199,N_3767,N_3039);
nand UO_200 (O_200,N_2565,N_4413);
or UO_201 (O_201,N_4940,N_2835);
nand UO_202 (O_202,N_4271,N_4450);
nand UO_203 (O_203,N_2608,N_4729);
nand UO_204 (O_204,N_4759,N_2983);
and UO_205 (O_205,N_2637,N_4817);
nor UO_206 (O_206,N_4811,N_2564);
or UO_207 (O_207,N_3442,N_2914);
nand UO_208 (O_208,N_3984,N_4339);
or UO_209 (O_209,N_4695,N_4346);
or UO_210 (O_210,N_4152,N_3128);
and UO_211 (O_211,N_2511,N_3591);
and UO_212 (O_212,N_3502,N_4635);
and UO_213 (O_213,N_3633,N_2525);
or UO_214 (O_214,N_4826,N_4994);
nor UO_215 (O_215,N_3405,N_4312);
and UO_216 (O_216,N_3270,N_3914);
and UO_217 (O_217,N_4276,N_2839);
and UO_218 (O_218,N_3781,N_3379);
and UO_219 (O_219,N_4638,N_3535);
nor UO_220 (O_220,N_4288,N_4868);
or UO_221 (O_221,N_4404,N_3943);
and UO_222 (O_222,N_4319,N_2603);
or UO_223 (O_223,N_4132,N_3518);
or UO_224 (O_224,N_3560,N_3892);
nor UO_225 (O_225,N_3068,N_4138);
or UO_226 (O_226,N_2867,N_4507);
nand UO_227 (O_227,N_3455,N_3493);
and UO_228 (O_228,N_4856,N_3619);
nand UO_229 (O_229,N_4675,N_3628);
and UO_230 (O_230,N_4069,N_4795);
nor UO_231 (O_231,N_3809,N_4465);
or UO_232 (O_232,N_2522,N_3569);
or UO_233 (O_233,N_3878,N_4949);
nand UO_234 (O_234,N_2851,N_3999);
nand UO_235 (O_235,N_3049,N_4738);
or UO_236 (O_236,N_3562,N_3683);
nor UO_237 (O_237,N_3365,N_2654);
and UO_238 (O_238,N_2904,N_2736);
and UO_239 (O_239,N_4569,N_4244);
nand UO_240 (O_240,N_2711,N_3963);
or UO_241 (O_241,N_3609,N_3002);
or UO_242 (O_242,N_2953,N_3790);
xnor UO_243 (O_243,N_4818,N_3386);
or UO_244 (O_244,N_3960,N_3905);
and UO_245 (O_245,N_3932,N_3792);
and UO_246 (O_246,N_2995,N_4015);
or UO_247 (O_247,N_4245,N_3038);
nor UO_248 (O_248,N_2888,N_3066);
nand UO_249 (O_249,N_3047,N_4869);
and UO_250 (O_250,N_3179,N_2507);
and UO_251 (O_251,N_4499,N_4731);
nand UO_252 (O_252,N_4907,N_4371);
and UO_253 (O_253,N_2797,N_2969);
and UO_254 (O_254,N_4599,N_3417);
nor UO_255 (O_255,N_4429,N_3627);
nor UO_256 (O_256,N_2804,N_3694);
nor UO_257 (O_257,N_3890,N_2911);
nand UO_258 (O_258,N_4515,N_3888);
nand UO_259 (O_259,N_2976,N_3430);
nor UO_260 (O_260,N_2631,N_4657);
and UO_261 (O_261,N_4060,N_2607);
and UO_262 (O_262,N_4734,N_3567);
nand UO_263 (O_263,N_2824,N_3147);
or UO_264 (O_264,N_4728,N_4632);
or UO_265 (O_265,N_3069,N_2865);
nor UO_266 (O_266,N_4694,N_4074);
nand UO_267 (O_267,N_4044,N_4681);
nand UO_268 (O_268,N_2644,N_2942);
and UO_269 (O_269,N_3603,N_3995);
and UO_270 (O_270,N_3697,N_4549);
nand UO_271 (O_271,N_4488,N_4398);
and UO_272 (O_272,N_2541,N_3225);
nand UO_273 (O_273,N_4494,N_3324);
and UO_274 (O_274,N_3927,N_4148);
nor UO_275 (O_275,N_2923,N_3070);
or UO_276 (O_276,N_2900,N_4093);
and UO_277 (O_277,N_3394,N_3821);
nor UO_278 (O_278,N_2859,N_4606);
and UO_279 (O_279,N_3116,N_4828);
or UO_280 (O_280,N_4884,N_2966);
nor UO_281 (O_281,N_3229,N_3681);
and UO_282 (O_282,N_3810,N_4272);
or UO_283 (O_283,N_3661,N_3725);
and UO_284 (O_284,N_4931,N_2934);
or UO_285 (O_285,N_3903,N_4440);
or UO_286 (O_286,N_3051,N_3608);
nor UO_287 (O_287,N_4673,N_4665);
nor UO_288 (O_288,N_4191,N_4929);
nand UO_289 (O_289,N_4899,N_4808);
or UO_290 (O_290,N_4495,N_4292);
or UO_291 (O_291,N_4580,N_3579);
nand UO_292 (O_292,N_2901,N_3739);
and UO_293 (O_293,N_3000,N_4330);
or UO_294 (O_294,N_4424,N_3848);
and UO_295 (O_295,N_3615,N_3482);
or UO_296 (O_296,N_2623,N_3185);
or UO_297 (O_297,N_3048,N_2821);
or UO_298 (O_298,N_3510,N_3658);
and UO_299 (O_299,N_3158,N_3117);
nor UO_300 (O_300,N_4246,N_4594);
and UO_301 (O_301,N_3614,N_4203);
and UO_302 (O_302,N_3308,N_2812);
nor UO_303 (O_303,N_2593,N_3275);
nor UO_304 (O_304,N_4480,N_4610);
or UO_305 (O_305,N_3329,N_2533);
nor UO_306 (O_306,N_3236,N_4207);
and UO_307 (O_307,N_3672,N_3434);
nor UO_308 (O_308,N_2915,N_3452);
nand UO_309 (O_309,N_4102,N_4916);
nand UO_310 (O_310,N_3557,N_2918);
nor UO_311 (O_311,N_4421,N_3642);
nand UO_312 (O_312,N_2611,N_3168);
nand UO_313 (O_313,N_3561,N_4299);
nand UO_314 (O_314,N_2710,N_4978);
nor UO_315 (O_315,N_4812,N_3432);
and UO_316 (O_316,N_3013,N_2534);
nor UO_317 (O_317,N_2931,N_4661);
nor UO_318 (O_318,N_4989,N_4823);
nor UO_319 (O_319,N_4853,N_3703);
nand UO_320 (O_320,N_3173,N_3315);
nand UO_321 (O_321,N_3779,N_3370);
or UO_322 (O_322,N_4432,N_4283);
nand UO_323 (O_323,N_3626,N_3363);
nand UO_324 (O_324,N_3273,N_3955);
nor UO_325 (O_325,N_4539,N_4653);
or UO_326 (O_326,N_4693,N_3197);
or UO_327 (O_327,N_4810,N_3431);
and UO_328 (O_328,N_4699,N_2509);
and UO_329 (O_329,N_3542,N_4139);
nor UO_330 (O_330,N_3915,N_2841);
and UO_331 (O_331,N_4822,N_2545);
and UO_332 (O_332,N_3975,N_3364);
and UO_333 (O_333,N_2606,N_2885);
nor UO_334 (O_334,N_2897,N_4352);
and UO_335 (O_335,N_4962,N_3233);
or UO_336 (O_336,N_4325,N_3859);
and UO_337 (O_337,N_2789,N_4749);
and UO_338 (O_338,N_3489,N_2540);
nor UO_339 (O_339,N_4315,N_3581);
nor UO_340 (O_340,N_3754,N_2902);
nor UO_341 (O_341,N_2634,N_4651);
nand UO_342 (O_342,N_4600,N_4342);
nand UO_343 (O_343,N_3139,N_3250);
nand UO_344 (O_344,N_4052,N_4264);
or UO_345 (O_345,N_4297,N_4086);
nor UO_346 (O_346,N_4608,N_4215);
and UO_347 (O_347,N_3228,N_2767);
or UO_348 (O_348,N_2700,N_2678);
nor UO_349 (O_349,N_4302,N_3961);
or UO_350 (O_350,N_3607,N_3505);
nor UO_351 (O_351,N_4677,N_4545);
or UO_352 (O_352,N_3026,N_4380);
nand UO_353 (O_353,N_3594,N_4561);
and UO_354 (O_354,N_4689,N_3934);
and UO_355 (O_355,N_3268,N_4141);
nand UO_356 (O_356,N_4038,N_3114);
or UO_357 (O_357,N_2601,N_4051);
and UO_358 (O_358,N_3151,N_2999);
or UO_359 (O_359,N_4784,N_3972);
nor UO_360 (O_360,N_3531,N_4702);
xnor UO_361 (O_361,N_2788,N_2968);
and UO_362 (O_362,N_3001,N_4792);
and UO_363 (O_363,N_4581,N_4946);
nand UO_364 (O_364,N_4998,N_4785);
and UO_365 (O_365,N_4630,N_3917);
and UO_366 (O_366,N_3974,N_4593);
and UO_367 (O_367,N_4745,N_3709);
and UO_368 (O_368,N_2553,N_2890);
nor UO_369 (O_369,N_3444,N_2825);
and UO_370 (O_370,N_3646,N_3241);
or UO_371 (O_371,N_4529,N_3260);
and UO_372 (O_372,N_4634,N_3320);
nand UO_373 (O_373,N_3372,N_4742);
or UO_374 (O_374,N_3412,N_4671);
nand UO_375 (O_375,N_4214,N_3936);
nor UO_376 (O_376,N_4877,N_2679);
or UO_377 (O_377,N_4053,N_3028);
nand UO_378 (O_378,N_4468,N_3336);
or UO_379 (O_379,N_4089,N_2558);
nand UO_380 (O_380,N_4033,N_3226);
nand UO_381 (O_381,N_4037,N_2980);
nand UO_382 (O_382,N_4752,N_3580);
or UO_383 (O_383,N_4754,N_2937);
or UO_384 (O_384,N_2520,N_3203);
or UO_385 (O_385,N_2621,N_2814);
nor UO_386 (O_386,N_3223,N_4136);
or UO_387 (O_387,N_4857,N_4162);
and UO_388 (O_388,N_3711,N_4239);
or UO_389 (O_389,N_3700,N_4551);
and UO_390 (O_390,N_4686,N_3701);
nand UO_391 (O_391,N_3045,N_3413);
and UO_392 (O_392,N_4577,N_2580);
or UO_393 (O_393,N_4306,N_3237);
nor UO_394 (O_394,N_4970,N_3109);
nand UO_395 (O_395,N_3732,N_4992);
nor UO_396 (O_396,N_3093,N_2528);
xor UO_397 (O_397,N_4603,N_3122);
or UO_398 (O_398,N_4969,N_2646);
and UO_399 (O_399,N_3637,N_4344);
nor UO_400 (O_400,N_3868,N_4519);
or UO_401 (O_401,N_3339,N_4224);
nand UO_402 (O_402,N_3317,N_3155);
or UO_403 (O_403,N_4168,N_4843);
and UO_404 (O_404,N_3351,N_4351);
xor UO_405 (O_405,N_3533,N_3328);
or UO_406 (O_406,N_2720,N_3578);
xnor UO_407 (O_407,N_4285,N_2583);
or UO_408 (O_408,N_3695,N_3087);
nand UO_409 (O_409,N_4801,N_2763);
nor UO_410 (O_410,N_3242,N_4256);
nor UO_411 (O_411,N_3880,N_3475);
xor UO_412 (O_412,N_2566,N_2828);
nor UO_413 (O_413,N_4447,N_4157);
nand UO_414 (O_414,N_4656,N_3105);
or UO_415 (O_415,N_4487,N_3485);
and UO_416 (O_416,N_3477,N_3301);
nor UO_417 (O_417,N_4228,N_4958);
and UO_418 (O_418,N_2847,N_4902);
nor UO_419 (O_419,N_4572,N_3251);
or UO_420 (O_420,N_3385,N_4883);
nand UO_421 (O_421,N_3470,N_4755);
or UO_422 (O_422,N_3393,N_4850);
and UO_423 (O_423,N_2731,N_3468);
and UO_424 (O_424,N_4280,N_2664);
or UO_425 (O_425,N_4890,N_4504);
nand UO_426 (O_426,N_4113,N_2523);
nand UO_427 (O_427,N_3967,N_2919);
or UO_428 (O_428,N_3211,N_2829);
or UO_429 (O_429,N_4087,N_2917);
or UO_430 (O_430,N_3724,N_3133);
and UO_431 (O_431,N_4201,N_4436);
or UO_432 (O_432,N_4803,N_3926);
nand UO_433 (O_433,N_4511,N_4067);
and UO_434 (O_434,N_3267,N_4724);
nand UO_435 (O_435,N_4835,N_3254);
and UO_436 (O_436,N_3281,N_4885);
and UO_437 (O_437,N_3164,N_3089);
or UO_438 (O_438,N_2775,N_3712);
and UO_439 (O_439,N_4932,N_3773);
nor UO_440 (O_440,N_3287,N_3110);
and UO_441 (O_441,N_4799,N_2690);
and UO_442 (O_442,N_4036,N_4396);
and UO_443 (O_443,N_4968,N_2536);
or UO_444 (O_444,N_2643,N_4733);
nor UO_445 (O_445,N_3077,N_4472);
nor UO_446 (O_446,N_2837,N_4977);
or UO_447 (O_447,N_2517,N_4879);
and UO_448 (O_448,N_2539,N_4441);
or UO_449 (O_449,N_3731,N_3832);
or UO_450 (O_450,N_4796,N_3215);
or UO_451 (O_451,N_3457,N_3909);
nand UO_452 (O_452,N_3186,N_3794);
and UO_453 (O_453,N_3536,N_4080);
and UO_454 (O_454,N_3255,N_3131);
nor UO_455 (O_455,N_2669,N_4887);
nand UO_456 (O_456,N_4290,N_3655);
and UO_457 (O_457,N_3702,N_3589);
nor UO_458 (O_458,N_4786,N_4891);
or UO_459 (O_459,N_4491,N_4181);
and UO_460 (O_460,N_4326,N_3752);
or UO_461 (O_461,N_3148,N_4337);
and UO_462 (O_462,N_4065,N_4045);
nand UO_463 (O_463,N_2674,N_4259);
nand UO_464 (O_464,N_4382,N_2779);
nand UO_465 (O_465,N_4629,N_4669);
nor UO_466 (O_466,N_4397,N_3796);
xnor UO_467 (O_467,N_4307,N_4068);
nand UO_468 (O_468,N_3214,N_2656);
and UO_469 (O_469,N_3021,N_4783);
and UO_470 (O_470,N_4541,N_3973);
nor UO_471 (O_471,N_3771,N_3404);
or UO_472 (O_472,N_4540,N_2752);
or UO_473 (O_473,N_3576,N_2940);
nand UO_474 (O_474,N_3611,N_4827);
nor UO_475 (O_475,N_2559,N_4725);
nand UO_476 (O_476,N_3183,N_2745);
and UO_477 (O_477,N_4788,N_4249);
or UO_478 (O_478,N_3503,N_2806);
and UO_479 (O_479,N_3075,N_4031);
nand UO_480 (O_480,N_3017,N_3181);
nor UO_481 (O_481,N_2684,N_3556);
and UO_482 (O_482,N_3074,N_3829);
and UO_483 (O_483,N_2884,N_3879);
nand UO_484 (O_484,N_4184,N_3808);
and UO_485 (O_485,N_4722,N_4736);
and UO_486 (O_486,N_3952,N_2777);
nand UO_487 (O_487,N_2605,N_2663);
nor UO_488 (O_488,N_2582,N_2948);
nand UO_489 (O_489,N_2747,N_3506);
and UO_490 (O_490,N_4955,N_3996);
and UO_491 (O_491,N_3881,N_4646);
and UO_492 (O_492,N_3248,N_3758);
nand UO_493 (O_493,N_2641,N_2675);
nand UO_494 (O_494,N_2826,N_4433);
nand UO_495 (O_495,N_3691,N_3869);
and UO_496 (O_496,N_3768,N_3525);
or UO_497 (O_497,N_3532,N_4105);
nor UO_498 (O_498,N_4825,N_4930);
nor UO_499 (O_499,N_2883,N_3940);
nor UO_500 (O_500,N_3022,N_4926);
or UO_501 (O_501,N_4097,N_3826);
or UO_502 (O_502,N_4937,N_4084);
or UO_503 (O_503,N_4643,N_3024);
nor UO_504 (O_504,N_4401,N_3572);
and UO_505 (O_505,N_3710,N_2945);
and UO_506 (O_506,N_2568,N_2960);
and UO_507 (O_507,N_4367,N_4003);
and UO_508 (O_508,N_4591,N_3309);
or UO_509 (O_509,N_3789,N_2970);
nand UO_510 (O_510,N_4019,N_2703);
and UO_511 (O_511,N_4913,N_3894);
nor UO_512 (O_512,N_2882,N_3037);
and UO_513 (O_513,N_3735,N_2869);
or UO_514 (O_514,N_2843,N_3950);
or UO_515 (O_515,N_3303,N_4430);
or UO_516 (O_516,N_2598,N_2896);
or UO_517 (O_517,N_4321,N_3828);
and UO_518 (O_518,N_4333,N_3132);
and UO_519 (O_519,N_3136,N_4816);
xnor UO_520 (O_520,N_4797,N_4912);
nand UO_521 (O_521,N_3778,N_4418);
nand UO_522 (O_522,N_3929,N_4819);
or UO_523 (O_523,N_3737,N_4237);
and UO_524 (O_524,N_4408,N_4091);
or UO_525 (O_525,N_2551,N_2667);
or UO_526 (O_526,N_4293,N_3083);
nand UO_527 (O_527,N_3948,N_4882);
nor UO_528 (O_528,N_3787,N_2887);
nor UO_529 (O_529,N_2864,N_4613);
nand UO_530 (O_530,N_3419,N_3545);
nand UO_531 (O_531,N_3863,N_2979);
nand UO_532 (O_532,N_2513,N_3188);
nor UO_533 (O_533,N_4167,N_4550);
and UO_534 (O_534,N_4373,N_4481);
and UO_535 (O_535,N_3715,N_4832);
and UO_536 (O_536,N_4637,N_2692);
nor UO_537 (O_537,N_3459,N_2697);
or UO_538 (O_538,N_3235,N_3722);
nand UO_539 (O_539,N_2996,N_4471);
and UO_540 (O_540,N_3427,N_2862);
and UO_541 (O_541,N_4170,N_4023);
or UO_542 (O_542,N_4741,N_3095);
or UO_543 (O_543,N_3727,N_2771);
and UO_544 (O_544,N_4462,N_4062);
or UO_545 (O_545,N_2689,N_2810);
and UO_546 (O_546,N_4649,N_4010);
nand UO_547 (O_547,N_4254,N_3396);
nor UO_548 (O_548,N_3717,N_3648);
xnor UO_549 (O_549,N_3507,N_2665);
nor UO_550 (O_550,N_2543,N_2640);
nor UO_551 (O_551,N_3057,N_3238);
nand UO_552 (O_552,N_4652,N_2881);
and UO_553 (O_553,N_2688,N_4836);
nor UO_554 (O_554,N_2921,N_2906);
nand UO_555 (O_555,N_4873,N_4225);
or UO_556 (O_556,N_4647,N_3392);
nand UO_557 (O_557,N_4303,N_3376);
and UO_558 (O_558,N_4452,N_4697);
nor UO_559 (O_559,N_4291,N_4235);
nor UO_560 (O_560,N_3761,N_4761);
and UO_561 (O_561,N_3639,N_2848);
nand UO_562 (O_562,N_3101,N_2502);
nor UO_563 (O_563,N_4378,N_4534);
nand UO_564 (O_564,N_4128,N_3456);
or UO_565 (O_565,N_3165,N_4971);
and UO_566 (O_566,N_3462,N_4586);
nor UO_567 (O_567,N_4353,N_2994);
nor UO_568 (O_568,N_4764,N_4178);
nor UO_569 (O_569,N_3682,N_3901);
and UO_570 (O_570,N_3873,N_4004);
and UO_571 (O_571,N_3990,N_3202);
and UO_572 (O_572,N_3337,N_4489);
nand UO_573 (O_573,N_4598,N_4155);
nor UO_574 (O_574,N_4135,N_3408);
and UO_575 (O_575,N_4718,N_4769);
nand UO_576 (O_576,N_4582,N_2616);
nand UO_577 (O_577,N_2992,N_4934);
nand UO_578 (O_578,N_4114,N_4642);
and UO_579 (O_579,N_2965,N_2956);
and UO_580 (O_580,N_4680,N_3606);
nor UO_581 (O_581,N_4921,N_3762);
nand UO_582 (O_582,N_3997,N_4445);
or UO_583 (O_583,N_2907,N_3175);
and UO_584 (O_584,N_3748,N_2782);
nand UO_585 (O_585,N_4837,N_4063);
and UO_586 (O_586,N_4154,N_3088);
nand UO_587 (O_587,N_3931,N_3791);
nor UO_588 (O_588,N_4995,N_3271);
nor UO_589 (O_589,N_3740,N_3193);
or UO_590 (O_590,N_2818,N_3343);
nand UO_591 (O_591,N_2721,N_4182);
nor UO_592 (O_592,N_3350,N_3205);
and UO_593 (O_593,N_4101,N_3447);
or UO_594 (O_594,N_2590,N_2653);
nand UO_595 (O_595,N_2677,N_2538);
nand UO_596 (O_596,N_3933,N_4234);
and UO_597 (O_597,N_3751,N_3509);
and UO_598 (O_598,N_3184,N_4809);
nand UO_599 (O_599,N_2702,N_4700);
or UO_600 (O_600,N_4894,N_3056);
nand UO_601 (O_601,N_4016,N_3182);
or UO_602 (O_602,N_3621,N_3423);
nand UO_603 (O_603,N_3192,N_2738);
nor UO_604 (O_604,N_4104,N_3541);
nor UO_605 (O_605,N_3448,N_4746);
or UO_606 (O_606,N_3852,N_3564);
nor UO_607 (O_607,N_2610,N_4011);
nand UO_608 (O_608,N_3016,N_4951);
nor UO_609 (O_609,N_4294,N_4518);
nor UO_610 (O_610,N_2898,N_4399);
nand UO_611 (O_611,N_3437,N_4715);
nand UO_612 (O_612,N_3811,N_4120);
or UO_613 (O_613,N_3563,N_4498);
and UO_614 (O_614,N_4895,N_2985);
and UO_615 (O_615,N_4781,N_2967);
and UO_616 (O_616,N_3369,N_4057);
nand UO_617 (O_617,N_3775,N_4530);
nand UO_618 (O_618,N_3605,N_4601);
and UO_619 (O_619,N_2760,N_4526);
nor UO_620 (O_620,N_3704,N_3582);
nor UO_621 (O_621,N_4324,N_4035);
nand UO_622 (O_622,N_3224,N_3245);
and UO_623 (O_623,N_4117,N_3671);
or UO_624 (O_624,N_2795,N_3322);
nand UO_625 (O_625,N_4950,N_2925);
and UO_626 (O_626,N_2769,N_4840);
and UO_627 (O_627,N_3750,N_2913);
nor UO_628 (O_628,N_3949,N_4553);
nand UO_629 (O_629,N_3402,N_4473);
and UO_630 (O_630,N_2870,N_2903);
nor UO_631 (O_631,N_3923,N_3583);
and UO_632 (O_632,N_4005,N_3588);
nor UO_633 (O_633,N_4639,N_3231);
nand UO_634 (O_634,N_3345,N_3550);
nand UO_635 (O_635,N_2527,N_2895);
nand UO_636 (O_636,N_3801,N_2627);
nor UO_637 (O_637,N_4939,N_3664);
and UO_638 (O_638,N_2672,N_2683);
nor UO_639 (O_639,N_4662,N_4683);
or UO_640 (O_640,N_3708,N_4477);
and UO_641 (O_641,N_4941,N_4001);
nor UO_642 (O_642,N_2503,N_4615);
xnor UO_643 (O_643,N_4568,N_4273);
nand UO_644 (O_644,N_3641,N_4517);
or UO_645 (O_645,N_4919,N_4112);
nand UO_646 (O_646,N_4150,N_3159);
and UO_647 (O_647,N_3492,N_4660);
nor UO_648 (O_648,N_2563,N_4286);
or UO_649 (O_649,N_3907,N_3367);
and UO_650 (O_650,N_4997,N_2694);
nand UO_651 (O_651,N_3433,N_2713);
and UO_652 (O_652,N_3010,N_3359);
or UO_653 (O_653,N_4012,N_3558);
nand UO_654 (O_654,N_3375,N_3566);
nand UO_655 (O_655,N_3669,N_3414);
nand UO_656 (O_656,N_4142,N_3660);
and UO_657 (O_657,N_4341,N_4027);
nand UO_658 (O_658,N_4360,N_3511);
and UO_659 (O_659,N_2785,N_3344);
or UO_660 (O_660,N_4088,N_4831);
nor UO_661 (O_661,N_4546,N_3253);
nand UO_662 (O_662,N_4099,N_2515);
and UO_663 (O_663,N_4760,N_4092);
and UO_664 (O_664,N_3970,N_2746);
nand UO_665 (O_665,N_3630,N_2626);
nor UO_666 (O_666,N_2737,N_2639);
or UO_667 (O_667,N_3980,N_3645);
or UO_668 (O_668,N_2705,N_3513);
nor UO_669 (O_669,N_3144,N_3079);
nand UO_670 (O_670,N_4703,N_3263);
and UO_671 (O_671,N_4573,N_2868);
and UO_672 (O_672,N_4327,N_4158);
and UO_673 (O_673,N_4200,N_4655);
and UO_674 (O_674,N_3650,N_4800);
and UO_675 (O_675,N_4654,N_4059);
or UO_676 (O_676,N_3520,N_3693);
and UO_677 (O_677,N_4107,N_3696);
or UO_678 (O_678,N_3877,N_4964);
nor UO_679 (O_679,N_4579,N_3575);
or UO_680 (O_680,N_4658,N_3246);
nor UO_681 (O_681,N_4247,N_4055);
and UO_682 (O_682,N_3785,N_2739);
and UO_683 (O_683,N_3378,N_4460);
nand UO_684 (O_684,N_4123,N_2959);
or UO_685 (O_685,N_3458,N_3743);
nor UO_686 (O_686,N_3465,N_3744);
nor UO_687 (O_687,N_3585,N_4542);
nand UO_688 (O_688,N_4552,N_2614);
nand UO_689 (O_689,N_4258,N_3593);
nor UO_690 (O_690,N_3857,N_3891);
or UO_691 (O_691,N_4388,N_3018);
or UO_692 (O_692,N_4867,N_3081);
or UO_693 (O_693,N_4766,N_3991);
nor UO_694 (O_694,N_4121,N_4083);
and UO_695 (O_695,N_3920,N_4779);
nand UO_696 (O_696,N_3041,N_4802);
nor UO_697 (O_697,N_3265,N_3257);
nor UO_698 (O_698,N_4709,N_3027);
and UO_699 (O_699,N_2830,N_3981);
or UO_700 (O_700,N_4354,N_4331);
nand UO_701 (O_701,N_4711,N_3052);
nor UO_702 (O_702,N_3438,N_4082);
and UO_703 (O_703,N_3549,N_3622);
nor UO_704 (O_704,N_4072,N_4943);
nand UO_705 (O_705,N_3800,N_3407);
and UO_706 (O_706,N_3374,N_2854);
and UO_707 (O_707,N_3469,N_3360);
nand UO_708 (O_708,N_4888,N_3986);
nand UO_709 (O_709,N_2505,N_3006);
nor UO_710 (O_710,N_3034,N_3688);
or UO_711 (O_711,N_2852,N_3276);
and UO_712 (O_712,N_4385,N_3401);
or UO_713 (O_713,N_2547,N_2939);
or UO_714 (O_714,N_3847,N_2586);
nand UO_715 (O_715,N_2941,N_4684);
nor UO_716 (O_716,N_4589,N_3126);
nand UO_717 (O_717,N_4417,N_2668);
and UO_718 (O_718,N_4316,N_4125);
or UO_719 (O_719,N_3783,N_4740);
or UO_720 (O_720,N_4389,N_4311);
or UO_721 (O_721,N_3684,N_4966);
and UO_722 (O_722,N_3156,N_4938);
or UO_723 (O_723,N_2905,N_3874);
or UO_724 (O_724,N_4512,N_4173);
nand UO_725 (O_725,N_4425,N_2971);
xnor UO_726 (O_726,N_3640,N_3261);
nor UO_727 (O_727,N_3340,N_2773);
nor UO_728 (O_728,N_3334,N_3239);
and UO_729 (O_729,N_4833,N_3551);
and UO_730 (O_730,N_3636,N_4336);
or UO_731 (O_731,N_2800,N_3802);
nor UO_732 (O_732,N_4438,N_3899);
nor UO_733 (O_733,N_2704,N_4146);
or UO_734 (O_734,N_3143,N_2891);
nand UO_735 (O_735,N_3098,N_4774);
or UO_736 (O_736,N_3924,N_2961);
or UO_737 (O_737,N_3091,N_3086);
or UO_738 (O_738,N_3323,N_4484);
nand UO_739 (O_739,N_3654,N_4230);
and UO_740 (O_740,N_4282,N_4437);
or UO_741 (O_741,N_4852,N_2922);
or UO_742 (O_742,N_2594,N_4190);
or UO_743 (O_743,N_4458,N_3042);
and UO_744 (O_744,N_4982,N_4268);
or UO_745 (O_745,N_4466,N_3195);
nor UO_746 (O_746,N_4422,N_2827);
nand UO_747 (O_747,N_4301,N_3352);
nor UO_748 (O_748,N_4743,N_3623);
nand UO_749 (O_749,N_2504,N_2638);
nor UO_750 (O_750,N_2975,N_2916);
or UO_751 (O_751,N_3055,N_3793);
nand UO_752 (O_752,N_3604,N_3656);
nor UO_753 (O_753,N_4505,N_4213);
nand UO_754 (O_754,N_3516,N_4804);
xor UO_755 (O_755,N_4688,N_2596);
nand UO_756 (O_756,N_4274,N_4231);
and UO_757 (O_757,N_3573,N_3481);
and UO_758 (O_758,N_4636,N_4516);
nand UO_759 (O_759,N_4240,N_3174);
and UO_760 (O_760,N_4641,N_3552);
nand UO_761 (O_761,N_3283,N_4987);
nand UO_762 (O_762,N_3978,N_2842);
and UO_763 (O_763,N_4563,N_3286);
or UO_764 (O_764,N_3613,N_4555);
or UO_765 (O_765,N_2575,N_3736);
nand UO_766 (O_766,N_4122,N_4513);
and UO_767 (O_767,N_4548,N_3454);
nor UO_768 (O_768,N_3100,N_4209);
or UO_769 (O_769,N_3358,N_2849);
nand UO_770 (O_770,N_3274,N_3499);
and UO_771 (O_771,N_3208,N_4892);
nor UO_772 (O_772,N_3795,N_3555);
nand UO_773 (O_773,N_4851,N_3335);
nor UO_774 (O_774,N_3134,N_4174);
nand UO_775 (O_775,N_2757,N_3851);
nand UO_776 (O_776,N_4323,N_3849);
nand UO_777 (O_777,N_4194,N_4845);
nor UO_778 (O_778,N_2764,N_3537);
nor UO_779 (O_779,N_4129,N_3657);
nand UO_780 (O_780,N_4767,N_4407);
and UO_781 (O_781,N_4570,N_3030);
or UO_782 (O_782,N_4620,N_2803);
nand UO_783 (O_783,N_3312,N_4227);
nand UO_784 (O_784,N_4145,N_2622);
nand UO_785 (O_785,N_3677,N_3474);
nor UO_786 (O_786,N_4974,N_4474);
or UO_787 (O_787,N_4262,N_3112);
nor UO_788 (O_788,N_3420,N_2875);
or UO_789 (O_789,N_3397,N_2792);
nand UO_790 (O_790,N_4775,N_2573);
nor UO_791 (O_791,N_2735,N_2928);
or UO_792 (O_792,N_4855,N_3104);
nand UO_793 (O_793,N_3160,N_2585);
nand UO_794 (O_794,N_3471,N_2579);
or UO_795 (O_795,N_4456,N_3338);
xnor UO_796 (O_796,N_3272,N_3939);
and UO_797 (O_797,N_4682,N_4196);
and UO_798 (O_798,N_2682,N_3592);
nand UO_799 (O_799,N_4278,N_2783);
or UO_800 (O_800,N_3953,N_4726);
or UO_801 (O_801,N_3911,N_3501);
nor UO_802 (O_802,N_3601,N_3377);
or UO_803 (O_803,N_2734,N_2524);
or UO_804 (O_804,N_3597,N_4910);
nor UO_805 (O_805,N_3220,N_4753);
nor UO_806 (O_806,N_4707,N_2612);
nor UO_807 (O_807,N_4604,N_3845);
or UO_808 (O_808,N_3756,N_2680);
nor UO_809 (O_809,N_4415,N_4216);
or UO_810 (O_810,N_3217,N_3747);
nand UO_811 (O_811,N_3096,N_3755);
nor UO_812 (O_812,N_4727,N_2617);
nor UO_813 (O_813,N_4866,N_3296);
or UO_814 (O_814,N_2531,N_3938);
nand UO_815 (O_815,N_4944,N_4041);
and UO_816 (O_816,N_3854,N_4261);
nor UO_817 (O_817,N_4134,N_2506);
or UO_818 (O_818,N_3992,N_4042);
nand UO_819 (O_819,N_3956,N_3586);
nand UO_820 (O_820,N_4131,N_3514);
nor UO_821 (O_821,N_3844,N_3020);
nor UO_822 (O_822,N_3094,N_3912);
nor UO_823 (O_823,N_4535,N_4403);
or UO_824 (O_824,N_3234,N_2550);
or UO_825 (O_825,N_4166,N_4757);
and UO_826 (O_826,N_3977,N_3007);
and UO_827 (O_827,N_4748,N_4449);
and UO_828 (O_828,N_3718,N_2958);
nor UO_829 (O_829,N_4963,N_3595);
and UO_830 (O_830,N_3476,N_4451);
nor UO_831 (O_831,N_3836,N_3870);
and UO_832 (O_832,N_3346,N_3252);
or UO_833 (O_833,N_3539,N_4790);
nor UO_834 (O_834,N_3774,N_2820);
and UO_835 (O_835,N_4130,N_2519);
nand UO_836 (O_836,N_3707,N_2698);
nor UO_837 (O_837,N_3472,N_4250);
nor UO_838 (O_838,N_3416,N_3130);
nand UO_839 (O_839,N_4763,N_3822);
nor UO_840 (O_840,N_2729,N_3944);
nor UO_841 (O_841,N_3705,N_2909);
nor UO_842 (O_842,N_4195,N_2834);
or UO_843 (O_843,N_4914,N_4750);
nand UO_844 (O_844,N_3326,N_4945);
or UO_845 (O_845,N_3698,N_4696);
nand UO_846 (O_846,N_3137,N_3982);
and UO_847 (O_847,N_4394,N_3118);
nand UO_848 (O_848,N_3080,N_3635);
nand UO_849 (O_849,N_3306,N_3035);
nor UO_850 (O_850,N_3054,N_4364);
and UO_851 (O_851,N_2572,N_2624);
and UO_852 (O_852,N_2920,N_4935);
and UO_853 (O_853,N_4270,N_4236);
and UO_854 (O_854,N_2687,N_3760);
nand UO_855 (O_855,N_3527,N_3676);
or UO_856 (O_856,N_4953,N_3867);
nand UO_857 (O_857,N_3764,N_4206);
nor UO_858 (O_858,N_4927,N_2998);
or UO_859 (O_859,N_4277,N_3834);
nand UO_860 (O_860,N_3721,N_4905);
nor UO_861 (O_861,N_2753,N_3050);
nor UO_862 (O_862,N_2832,N_4571);
or UO_863 (O_863,N_4233,N_2725);
and UO_864 (O_864,N_3102,N_4435);
or UO_865 (O_865,N_3127,N_4815);
nor UO_866 (O_866,N_4501,N_2761);
nor UO_867 (O_867,N_2899,N_3441);
nand UO_868 (O_868,N_3478,N_4592);
and UO_869 (O_869,N_2570,N_4676);
nand UO_870 (O_870,N_2748,N_2823);
and UO_871 (O_871,N_2567,N_4454);
and UO_872 (O_872,N_4644,N_3073);
or UO_873 (O_873,N_4475,N_3816);
nand UO_874 (O_874,N_4295,N_3624);
nand UO_875 (O_875,N_4625,N_4988);
nor UO_876 (O_876,N_3908,N_2805);
or UO_877 (O_877,N_2873,N_4744);
or UO_878 (O_878,N_4878,N_3540);
nand UO_879 (O_879,N_4358,N_4405);
or UO_880 (O_880,N_2787,N_2562);
and UO_881 (O_881,N_3644,N_2655);
and UO_882 (O_882,N_4284,N_4025);
or UO_883 (O_883,N_3483,N_4387);
and UO_884 (O_884,N_3319,N_3140);
and UO_885 (O_885,N_2776,N_4357);
and UO_886 (O_886,N_4374,N_4177);
and UO_887 (O_887,N_2707,N_3446);
nor UO_888 (O_888,N_4176,N_2872);
nor UO_889 (O_889,N_4915,N_4900);
or UO_890 (O_890,N_4906,N_2982);
or UO_891 (O_891,N_2780,N_3596);
or UO_892 (O_892,N_3498,N_2717);
nor UO_893 (O_893,N_4410,N_4251);
nor UO_894 (O_894,N_4165,N_4204);
and UO_895 (O_895,N_2514,N_4633);
or UO_896 (O_896,N_3951,N_4985);
nor UO_897 (O_897,N_4147,N_4241);
xnor UO_898 (O_898,N_2947,N_3153);
nand UO_899 (O_899,N_2595,N_4296);
nor UO_900 (O_900,N_3436,N_3521);
and UO_901 (O_901,N_3125,N_4058);
and UO_902 (O_902,N_4193,N_3357);
nand UO_903 (O_903,N_3853,N_2924);
or UO_904 (O_904,N_4880,N_2977);
nand UO_905 (O_905,N_4936,N_4805);
nor UO_906 (O_906,N_3837,N_3222);
and UO_907 (O_907,N_3815,N_4560);
and UO_908 (O_908,N_3757,N_4617);
and UO_909 (O_909,N_4980,N_2628);
or UO_910 (O_910,N_3987,N_4874);
nand UO_911 (O_911,N_4281,N_3046);
or UO_912 (O_912,N_2548,N_3316);
nand UO_913 (O_913,N_4395,N_2816);
or UO_914 (O_914,N_4169,N_3517);
or UO_915 (O_915,N_4557,N_4211);
nor UO_916 (O_916,N_4778,N_3428);
or UO_917 (O_917,N_2938,N_4527);
nor UO_918 (O_918,N_4492,N_3227);
and UO_919 (O_919,N_2819,N_3025);
nor UO_920 (O_920,N_4149,N_4002);
xor UO_921 (O_921,N_4663,N_3445);
and UO_922 (O_922,N_4386,N_2620);
and UO_923 (O_923,N_2831,N_3631);
and UO_924 (O_924,N_4076,N_4532);
or UO_925 (O_925,N_3994,N_3679);
nand UO_926 (O_926,N_3598,N_2963);
nor UO_927 (O_927,N_4863,N_4679);
or UO_928 (O_928,N_4793,N_4223);
or UO_929 (O_929,N_3204,N_4576);
nor UO_930 (O_930,N_4338,N_3893);
nor UO_931 (O_931,N_3293,N_4304);
nand UO_932 (O_932,N_4854,N_3653);
and UO_933 (O_933,N_4106,N_4583);
or UO_934 (O_934,N_2518,N_4431);
nand UO_935 (O_935,N_3529,N_2944);
and UO_936 (O_936,N_4161,N_4578);
nor UO_937 (O_937,N_4266,N_4607);
and UO_938 (O_938,N_2936,N_4543);
nor UO_939 (O_939,N_4710,N_3763);
and UO_940 (O_940,N_2693,N_3097);
or UO_941 (O_941,N_3985,N_2730);
nand UO_942 (O_942,N_4536,N_3508);
nor UO_943 (O_943,N_4029,N_2602);
nor UO_944 (O_944,N_4381,N_3989);
nand UO_945 (O_945,N_3004,N_4009);
nand UO_946 (O_946,N_2632,N_2662);
nor UO_947 (O_947,N_3141,N_3813);
or UO_948 (O_948,N_4420,N_2681);
nor UO_949 (O_949,N_4509,N_4538);
or UO_950 (O_950,N_4503,N_2578);
and UO_951 (O_951,N_2574,N_4901);
or UO_952 (O_952,N_2943,N_2790);
nor UO_953 (O_953,N_4279,N_4022);
nor UO_954 (O_954,N_4876,N_2755);
or UO_955 (O_955,N_4309,N_4024);
or UO_956 (O_956,N_2802,N_4075);
and UO_957 (O_957,N_2799,N_3916);
nor UO_958 (O_958,N_4054,N_3063);
nor UO_959 (O_959,N_4255,N_2889);
nor UO_960 (O_960,N_2577,N_4862);
and UO_961 (O_961,N_2952,N_2770);
or UO_962 (O_962,N_3187,N_4911);
nor UO_963 (O_963,N_4500,N_4419);
nand UO_964 (O_964,N_4618,N_4627);
nand UO_965 (O_965,N_3003,N_2973);
nand UO_966 (O_966,N_4478,N_4383);
and UO_967 (O_967,N_3766,N_3780);
nand UO_968 (O_968,N_4164,N_3692);
or UO_969 (O_969,N_3464,N_3023);
and UO_970 (O_970,N_3219,N_3387);
nor UO_971 (O_971,N_3786,N_4575);
nand UO_972 (O_972,N_4081,N_3353);
nand UO_973 (O_973,N_3044,N_3957);
nand UO_974 (O_974,N_3058,N_2894);
and UO_975 (O_975,N_2552,N_4972);
nor UO_976 (O_976,N_2778,N_4948);
nor UO_977 (O_977,N_3497,N_3422);
or UO_978 (O_978,N_4275,N_2714);
or UO_979 (O_979,N_4253,N_4453);
nand UO_980 (O_980,N_4412,N_4100);
and UO_981 (O_981,N_4359,N_2609);
nand UO_982 (O_982,N_2912,N_3180);
or UO_983 (O_983,N_3232,N_4574);
or UO_984 (O_984,N_3629,N_4476);
or UO_985 (O_985,N_3082,N_4366);
or UO_986 (O_986,N_4124,N_2649);
or UO_987 (O_987,N_4070,N_3675);
and UO_988 (O_988,N_4391,N_3906);
nand UO_989 (O_989,N_4014,N_3171);
or UO_990 (O_990,N_3366,N_4942);
nand UO_991 (O_991,N_2599,N_3201);
and UO_992 (O_992,N_3106,N_2629);
or UO_993 (O_993,N_4026,N_4849);
nor UO_994 (O_994,N_4127,N_3170);
or UO_995 (O_995,N_3803,N_4221);
nand UO_996 (O_996,N_4314,N_4242);
and UO_997 (O_997,N_2592,N_4180);
nor UO_998 (O_998,N_2988,N_4904);
nor UO_999 (O_999,N_3247,N_2532);
endmodule