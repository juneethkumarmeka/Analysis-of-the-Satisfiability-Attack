module basic_2500_25000_3000_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_505,In_2428);
and U1 (N_1,In_2453,In_685);
nand U2 (N_2,In_2373,In_2334);
nand U3 (N_3,In_2017,In_2451);
or U4 (N_4,In_408,In_1754);
or U5 (N_5,In_17,In_584);
nand U6 (N_6,In_2374,In_519);
and U7 (N_7,In_1230,In_1522);
and U8 (N_8,In_2426,In_1502);
nor U9 (N_9,In_2155,In_2203);
nor U10 (N_10,In_1246,In_382);
and U11 (N_11,In_1590,In_2488);
nand U12 (N_12,In_756,In_496);
and U13 (N_13,In_867,In_1922);
and U14 (N_14,In_315,In_527);
and U15 (N_15,In_2268,In_1232);
or U16 (N_16,In_1313,In_2255);
or U17 (N_17,In_615,In_153);
or U18 (N_18,In_1802,In_2404);
nor U19 (N_19,In_281,In_1954);
nand U20 (N_20,In_1379,In_28);
or U21 (N_21,In_1739,In_2183);
and U22 (N_22,In_1799,In_1850);
xnor U23 (N_23,In_1082,In_1429);
nor U24 (N_24,In_1872,In_2001);
nor U25 (N_25,In_658,In_1224);
nand U26 (N_26,In_856,In_46);
and U27 (N_27,In_363,In_356);
xnor U28 (N_28,In_1844,In_344);
nand U29 (N_29,In_889,In_1177);
or U30 (N_30,In_1801,In_574);
nor U31 (N_31,In_249,In_455);
or U32 (N_32,In_1603,In_2012);
nor U33 (N_33,In_1772,In_438);
xnor U34 (N_34,In_1228,In_553);
or U35 (N_35,In_536,In_499);
and U36 (N_36,In_969,In_1178);
or U37 (N_37,In_2124,In_1546);
or U38 (N_38,In_482,In_1107);
and U39 (N_39,In_1867,In_732);
and U40 (N_40,In_1573,In_1255);
xnor U41 (N_41,In_504,In_2260);
and U42 (N_42,In_336,In_1800);
and U43 (N_43,In_1466,In_69);
nand U44 (N_44,In_1758,In_1181);
nand U45 (N_45,In_529,In_650);
and U46 (N_46,In_2135,In_1910);
nor U47 (N_47,In_2307,In_1747);
or U48 (N_48,In_1184,In_1681);
nor U49 (N_49,In_287,In_2091);
nor U50 (N_50,In_1698,In_88);
or U51 (N_51,In_1881,In_82);
nor U52 (N_52,In_1212,In_781);
or U53 (N_53,In_47,In_908);
and U54 (N_54,In_722,In_6);
xnor U55 (N_55,In_864,In_152);
nand U56 (N_56,In_1609,In_823);
nor U57 (N_57,In_1500,In_852);
and U58 (N_58,In_888,In_105);
xnor U59 (N_59,In_2010,In_21);
and U60 (N_60,In_592,In_510);
nor U61 (N_61,In_2213,In_237);
nor U62 (N_62,In_1266,In_1200);
xor U63 (N_63,In_760,In_911);
and U64 (N_64,In_2154,In_954);
and U65 (N_65,In_1841,In_1796);
or U66 (N_66,In_1656,In_1343);
nor U67 (N_67,In_2371,In_1786);
nand U68 (N_68,In_447,In_330);
or U69 (N_69,In_1891,In_1365);
nor U70 (N_70,In_2323,In_525);
nand U71 (N_71,In_1068,In_746);
or U72 (N_72,In_557,In_1031);
nor U73 (N_73,In_1939,In_426);
and U74 (N_74,In_668,In_2342);
nor U75 (N_75,In_1812,In_812);
nand U76 (N_76,In_1767,In_1140);
or U77 (N_77,In_342,In_484);
nand U78 (N_78,In_2184,In_1706);
or U79 (N_79,In_577,In_2309);
and U80 (N_80,In_905,In_2249);
nand U81 (N_81,In_1483,In_2463);
or U82 (N_82,In_1599,In_1871);
nand U83 (N_83,In_871,In_2347);
nor U84 (N_84,In_294,In_590);
nand U85 (N_85,In_1790,In_2176);
nor U86 (N_86,In_2494,In_646);
or U87 (N_87,In_815,In_593);
nand U88 (N_88,In_440,In_1370);
nor U89 (N_89,In_2218,In_478);
xnor U90 (N_90,In_236,In_1159);
or U91 (N_91,In_1852,In_120);
and U92 (N_92,In_853,In_1962);
and U93 (N_93,In_524,In_1320);
xnor U94 (N_94,In_1651,In_2002);
xor U95 (N_95,In_2493,In_1303);
xnor U96 (N_96,In_755,In_99);
nor U97 (N_97,In_149,In_544);
and U98 (N_98,In_422,In_2125);
nand U99 (N_99,In_1360,In_1007);
and U100 (N_100,In_807,In_246);
and U101 (N_101,In_443,In_475);
or U102 (N_102,In_1538,In_979);
and U103 (N_103,In_2299,In_345);
or U104 (N_104,In_174,In_10);
nand U105 (N_105,In_1334,In_873);
xnor U106 (N_106,In_2093,In_890);
xor U107 (N_107,In_625,In_1416);
and U108 (N_108,In_1724,In_663);
xor U109 (N_109,In_1037,In_2330);
or U110 (N_110,In_2219,In_83);
and U111 (N_111,In_456,In_2057);
nor U112 (N_112,In_1208,In_2435);
or U113 (N_113,In_224,In_1169);
and U114 (N_114,In_1444,In_1057);
and U115 (N_115,In_2384,In_697);
xnor U116 (N_116,In_1602,In_859);
and U117 (N_117,In_2272,In_1435);
nor U118 (N_118,In_328,In_1322);
or U119 (N_119,In_2465,In_1620);
or U120 (N_120,In_513,In_1991);
nor U121 (N_121,In_517,In_1482);
xnor U122 (N_122,In_2430,In_2496);
or U123 (N_123,In_2170,In_521);
or U124 (N_124,In_948,In_1015);
xor U125 (N_125,In_273,In_2225);
and U126 (N_126,In_1845,In_441);
nor U127 (N_127,In_1454,In_2150);
nor U128 (N_128,In_816,In_599);
nand U129 (N_129,In_61,In_1022);
nor U130 (N_130,In_2245,In_1137);
or U131 (N_131,In_860,In_1869);
nand U132 (N_132,In_1198,In_789);
nand U133 (N_133,In_1557,In_2321);
and U134 (N_134,In_1286,In_2437);
and U135 (N_135,In_1262,In_636);
nand U136 (N_136,In_1021,In_2224);
or U137 (N_137,In_762,In_213);
and U138 (N_138,In_2174,In_1525);
nor U139 (N_139,In_1146,In_2270);
xnor U140 (N_140,In_724,In_1478);
nand U141 (N_141,In_269,In_1851);
xnor U142 (N_142,In_768,In_1696);
or U143 (N_143,In_2181,In_2398);
nor U144 (N_144,In_2499,In_2177);
nor U145 (N_145,In_813,In_824);
and U146 (N_146,In_1979,In_1367);
or U147 (N_147,In_1016,In_1849);
xnor U148 (N_148,In_208,In_1472);
or U149 (N_149,In_2305,In_151);
and U150 (N_150,In_1654,In_1885);
or U151 (N_151,In_2208,In_148);
and U152 (N_152,In_1475,In_63);
and U153 (N_153,In_167,In_1364);
xnor U154 (N_154,In_1161,In_329);
nand U155 (N_155,In_1465,In_1927);
nor U156 (N_156,In_1858,In_1539);
xnor U157 (N_157,In_952,In_2236);
and U158 (N_158,In_474,In_1086);
nor U159 (N_159,In_512,In_2345);
or U160 (N_160,In_2361,In_1090);
and U161 (N_161,In_1211,In_1529);
and U162 (N_162,In_1895,In_218);
or U163 (N_163,In_2313,In_1026);
and U164 (N_164,In_935,In_189);
nand U165 (N_165,In_1759,In_212);
xnor U166 (N_166,In_947,In_2264);
nand U167 (N_167,In_155,In_1403);
xor U168 (N_168,In_839,In_645);
and U169 (N_169,In_40,In_1668);
nor U170 (N_170,In_1160,In_891);
or U171 (N_171,In_371,In_1480);
nor U172 (N_172,In_624,In_922);
and U173 (N_173,In_1730,In_678);
or U174 (N_174,In_1325,In_876);
nand U175 (N_175,In_534,In_316);
xor U176 (N_176,In_731,In_2073);
xnor U177 (N_177,In_1302,In_1513);
and U178 (N_178,In_1448,In_3);
or U179 (N_179,In_1804,In_1521);
nand U180 (N_180,In_940,In_292);
nor U181 (N_181,In_2257,In_2033);
xor U182 (N_182,In_2417,In_1424);
nand U183 (N_183,In_333,In_106);
or U184 (N_184,In_1616,In_1055);
and U185 (N_185,In_798,In_11);
nand U186 (N_186,In_2215,In_1578);
nor U187 (N_187,In_960,In_2084);
nand U188 (N_188,In_2030,In_690);
and U189 (N_189,In_479,In_1911);
xor U190 (N_190,In_405,In_1685);
xnor U191 (N_191,In_469,In_1652);
nor U192 (N_192,In_1614,In_1226);
nor U193 (N_193,In_1780,In_2369);
xor U194 (N_194,In_702,In_1234);
and U195 (N_195,In_1565,In_162);
and U196 (N_196,In_729,In_666);
xor U197 (N_197,In_2442,In_930);
or U198 (N_198,In_270,In_2092);
and U199 (N_199,In_1278,In_1915);
xor U200 (N_200,In_1241,In_1151);
and U201 (N_201,In_2348,In_1079);
and U202 (N_202,In_1345,In_1105);
xnor U203 (N_203,In_2405,In_700);
nand U204 (N_204,In_235,In_1680);
and U205 (N_205,In_2443,In_1704);
or U206 (N_206,In_1664,In_620);
or U207 (N_207,In_64,In_1768);
and U208 (N_208,In_29,In_1694);
or U209 (N_209,In_1422,In_1324);
or U210 (N_210,In_2069,In_1914);
and U211 (N_211,In_2271,In_2157);
and U212 (N_212,In_656,In_1217);
xor U213 (N_213,In_2175,In_2473);
nor U214 (N_214,In_1346,In_2457);
xor U215 (N_215,In_794,In_628);
nor U216 (N_216,In_412,In_2138);
xnor U217 (N_217,In_243,In_753);
xor U218 (N_218,In_95,In_1814);
and U219 (N_219,In_424,In_2188);
or U220 (N_220,In_2034,In_1762);
xor U221 (N_221,In_1705,In_288);
and U222 (N_222,In_537,In_2427);
or U223 (N_223,In_1632,In_101);
or U224 (N_224,In_214,In_1611);
or U225 (N_225,In_738,In_1818);
xor U226 (N_226,In_248,In_837);
and U227 (N_227,In_79,In_809);
nor U228 (N_228,In_141,In_1013);
nor U229 (N_229,In_1039,In_1798);
nor U230 (N_230,In_1221,In_1485);
nand U231 (N_231,In_2031,In_130);
and U232 (N_232,In_460,In_104);
or U233 (N_233,In_875,In_1456);
or U234 (N_234,In_1463,In_1156);
nor U235 (N_235,In_1714,In_2195);
nor U236 (N_236,In_406,In_1537);
and U237 (N_237,In_623,In_1366);
xnor U238 (N_238,In_1846,In_1750);
or U239 (N_239,In_1725,In_546);
and U240 (N_240,In_276,In_1859);
nand U241 (N_241,In_93,In_1967);
nor U242 (N_242,In_1552,In_1987);
xnor U243 (N_243,In_800,In_1516);
and U244 (N_244,In_486,In_1820);
nand U245 (N_245,In_579,In_819);
and U246 (N_246,In_638,In_974);
nor U247 (N_247,In_2179,In_296);
and U248 (N_248,In_1375,In_2288);
nor U249 (N_249,In_1190,In_1476);
nand U250 (N_250,In_1707,In_1534);
xor U251 (N_251,In_1604,In_785);
and U252 (N_252,In_659,In_1250);
nor U253 (N_253,In_733,In_1102);
nor U254 (N_254,In_1936,In_57);
xor U255 (N_255,In_507,In_1660);
nor U256 (N_256,In_2353,In_634);
nand U257 (N_257,In_164,In_1460);
nor U258 (N_258,In_59,In_439);
nand U259 (N_259,In_2087,In_1711);
xnor U260 (N_260,In_432,In_1765);
nor U261 (N_261,In_1506,In_2379);
or U262 (N_262,In_1623,In_1917);
and U263 (N_263,In_2376,In_2327);
nand U264 (N_264,In_1543,In_2005);
xnor U265 (N_265,In_65,In_264);
or U266 (N_266,In_1204,In_2137);
nor U267 (N_267,In_644,In_2252);
and U268 (N_268,In_274,In_1209);
or U269 (N_269,In_283,In_415);
nor U270 (N_270,In_126,In_914);
or U271 (N_271,In_1000,In_290);
and U272 (N_272,In_1880,In_1587);
and U273 (N_273,In_2067,In_467);
or U274 (N_274,In_1127,In_1023);
xor U275 (N_275,In_767,In_1598);
nor U276 (N_276,In_770,In_530);
nand U277 (N_277,In_882,In_1843);
xnor U278 (N_278,In_1953,In_1621);
nand U279 (N_279,In_848,In_887);
xor U280 (N_280,In_1828,In_1999);
or U281 (N_281,In_1912,In_2212);
and U282 (N_282,In_1884,In_1008);
xor U283 (N_283,In_540,In_221);
nor U284 (N_284,In_796,In_588);
or U285 (N_285,In_1899,In_1358);
nor U286 (N_286,In_2363,In_701);
and U287 (N_287,In_2364,In_70);
and U288 (N_288,In_991,In_2011);
nand U289 (N_289,In_1053,In_437);
and U290 (N_290,In_1029,In_2356);
xor U291 (N_291,In_254,In_1333);
nor U292 (N_292,In_1494,In_1940);
xnor U293 (N_293,In_1699,In_124);
xor U294 (N_294,In_619,In_1318);
nand U295 (N_295,In_334,In_2482);
nor U296 (N_296,In_1340,In_2394);
xor U297 (N_297,In_1701,In_1390);
or U298 (N_298,In_2253,In_2420);
or U299 (N_299,In_1183,In_399);
nand U300 (N_300,In_721,In_1256);
nor U301 (N_301,In_1982,In_715);
nor U302 (N_302,In_1094,In_1756);
or U303 (N_303,In_2332,In_727);
and U304 (N_304,In_1376,In_554);
xor U305 (N_305,In_1109,In_917);
xor U306 (N_306,In_869,In_1959);
nand U307 (N_307,In_341,In_1129);
nand U308 (N_308,In_2080,In_1964);
xor U309 (N_309,In_841,In_985);
nor U310 (N_310,In_1042,In_1838);
nor U311 (N_311,In_188,In_1687);
nor U312 (N_312,In_2226,In_2285);
or U313 (N_313,In_2397,In_718);
or U314 (N_314,In_2378,In_497);
and U315 (N_315,In_1244,In_2411);
xor U316 (N_316,In_2278,In_1051);
and U317 (N_317,In_2118,In_1847);
nand U318 (N_318,In_855,In_844);
or U319 (N_319,In_203,In_123);
nor U320 (N_320,In_1399,In_2282);
nand U321 (N_321,In_1793,In_2450);
nor U322 (N_322,In_778,In_1001);
nor U323 (N_323,In_2265,In_1888);
and U324 (N_324,In_1996,In_944);
xor U325 (N_325,In_2362,In_1056);
xor U326 (N_326,In_925,In_159);
and U327 (N_327,In_339,In_1520);
nand U328 (N_328,In_657,In_231);
nand U329 (N_329,In_490,In_388);
nor U330 (N_330,In_2359,In_118);
and U331 (N_331,In_2237,In_1957);
or U332 (N_332,In_1458,In_319);
xor U333 (N_333,In_2075,In_1717);
nand U334 (N_334,In_35,In_1906);
or U335 (N_335,In_215,In_977);
or U336 (N_336,In_639,In_1132);
xnor U337 (N_337,In_1561,In_850);
xnor U338 (N_338,In_1973,In_2015);
nor U339 (N_339,In_1378,In_1570);
or U340 (N_340,In_2455,In_1298);
and U341 (N_341,In_1736,In_1721);
nor U342 (N_342,In_711,In_495);
nand U343 (N_343,In_1175,In_987);
xnor U344 (N_344,In_2107,In_547);
nand U345 (N_345,In_2214,In_2304);
xor U346 (N_346,In_1672,In_774);
or U347 (N_347,In_373,In_862);
xor U348 (N_348,In_626,In_2419);
nor U349 (N_349,In_261,In_600);
xor U350 (N_350,In_902,In_1417);
or U351 (N_351,In_133,In_1138);
nor U352 (N_352,In_1541,In_1729);
nand U353 (N_353,In_779,In_16);
or U354 (N_354,In_522,In_1391);
nor U355 (N_355,In_383,In_278);
and U356 (N_356,In_2368,In_849);
xnor U357 (N_357,In_1653,In_631);
xor U358 (N_358,In_1369,In_128);
or U359 (N_359,In_431,In_1594);
or U360 (N_360,In_2349,In_2040);
or U361 (N_361,In_103,In_2467);
or U362 (N_362,In_1389,In_451);
nor U363 (N_363,In_2338,In_1331);
nand U364 (N_364,In_2143,In_158);
xor U365 (N_365,In_1533,In_298);
nor U366 (N_366,In_321,In_306);
xor U367 (N_367,In_532,In_2166);
xnor U368 (N_368,In_466,In_1792);
and U369 (N_369,In_48,In_1441);
or U370 (N_370,In_750,In_1060);
xor U371 (N_371,In_2227,In_1062);
and U372 (N_372,In_239,In_42);
nand U373 (N_373,In_200,In_1203);
nand U374 (N_374,In_2382,In_323);
xnor U375 (N_375,In_1174,In_1356);
xnor U376 (N_376,In_303,In_2461);
xnor U377 (N_377,In_1644,In_1030);
xnor U378 (N_378,In_1312,In_913);
xnor U379 (N_379,In_181,In_2229);
and U380 (N_380,In_2325,In_618);
xnor U381 (N_381,In_187,In_1426);
xor U382 (N_382,In_801,In_771);
xor U383 (N_383,In_1201,In_1760);
and U384 (N_384,In_1288,In_2019);
or U385 (N_385,In_1737,In_1104);
or U386 (N_386,In_2308,In_1150);
nor U387 (N_387,In_222,In_1193);
or U388 (N_388,In_607,In_2127);
or U389 (N_389,In_1924,In_1410);
nand U390 (N_390,In_1931,In_1547);
nand U391 (N_391,In_461,In_44);
xor U392 (N_392,In_327,In_166);
and U393 (N_393,In_19,In_1024);
xnor U394 (N_394,In_1716,In_780);
nand U395 (N_395,In_1438,In_1819);
nand U396 (N_396,In_1240,In_608);
and U397 (N_397,In_1111,In_2258);
or U398 (N_398,In_2395,In_2238);
and U399 (N_399,In_1134,In_1144);
nand U400 (N_400,In_1563,In_393);
xnor U401 (N_401,In_585,In_372);
xnor U402 (N_402,In_216,In_2210);
or U403 (N_403,In_705,In_1070);
nor U404 (N_404,In_1607,In_555);
nor U405 (N_405,In_468,In_1341);
or U406 (N_406,In_241,In_1344);
or U407 (N_407,In_1167,In_27);
nor U408 (N_408,In_1682,In_2475);
nor U409 (N_409,In_1690,In_660);
nand U410 (N_410,In_986,In_1427);
and U411 (N_411,In_2312,In_2331);
nand U412 (N_412,In_1077,In_1098);
xnor U413 (N_413,In_317,In_1374);
xor U414 (N_414,In_539,In_936);
xor U415 (N_415,In_352,In_2162);
and U416 (N_416,In_1164,In_835);
xor U417 (N_417,In_2491,In_442);
and U418 (N_418,In_41,In_2160);
xnor U419 (N_419,In_597,In_2410);
or U420 (N_420,In_545,In_18);
or U421 (N_421,In_1254,In_217);
xnor U422 (N_422,In_2167,In_146);
nor U423 (N_423,In_1301,In_1745);
xor U424 (N_424,In_420,In_1815);
xor U425 (N_425,In_309,In_1045);
or U426 (N_426,In_1469,In_693);
nand U427 (N_427,In_2365,In_1139);
nor U428 (N_428,In_1257,In_1723);
nor U429 (N_429,In_1452,In_1455);
and U430 (N_430,In_2099,In_1113);
xor U431 (N_431,In_635,In_15);
xor U432 (N_432,In_178,In_307);
nand U433 (N_433,In_2490,In_1227);
nand U434 (N_434,In_7,In_2063);
xor U435 (N_435,In_1304,In_1329);
nand U436 (N_436,In_260,In_2027);
nand U437 (N_437,In_1133,In_156);
nand U438 (N_438,In_1994,In_761);
xnor U439 (N_439,In_2277,In_2098);
nand U440 (N_440,In_509,In_1596);
or U441 (N_441,In_161,In_942);
and U442 (N_442,In_684,In_282);
nand U443 (N_443,In_1453,In_1805);
or U444 (N_444,In_1807,In_2100);
nand U445 (N_445,In_1213,In_804);
nor U446 (N_446,In_1586,In_2316);
or U447 (N_447,In_2440,In_1662);
and U448 (N_448,In_1507,In_5);
and U449 (N_449,In_80,In_1613);
nand U450 (N_450,In_654,In_2464);
or U451 (N_451,In_271,In_347);
nand U452 (N_452,In_1670,In_168);
or U453 (N_453,In_1330,In_528);
or U454 (N_454,In_1925,In_2128);
or U455 (N_455,In_1528,In_1011);
nand U456 (N_456,In_857,In_473);
and U457 (N_457,In_295,In_1530);
or U458 (N_458,In_1649,In_1131);
xor U459 (N_459,In_671,In_872);
xor U460 (N_460,In_783,In_1985);
nor U461 (N_461,In_1921,In_1813);
nand U462 (N_462,In_357,In_22);
and U463 (N_463,In_1856,In_683);
or U464 (N_464,In_2003,In_2014);
nand U465 (N_465,In_494,In_1806);
nand U466 (N_466,In_1323,In_829);
xnor U467 (N_467,In_833,In_953);
nor U468 (N_468,In_1674,In_210);
and U469 (N_469,In_707,In_2117);
or U470 (N_470,In_1440,In_1210);
and U471 (N_471,In_962,In_233);
and U472 (N_472,In_1617,In_1835);
and U473 (N_473,In_941,In_476);
and U474 (N_474,In_2295,In_2487);
xor U475 (N_475,In_531,In_591);
or U476 (N_476,In_2452,In_183);
or U477 (N_477,In_1752,In_831);
nand U478 (N_478,In_1997,In_1788);
or U479 (N_479,In_2201,In_2424);
xor U480 (N_480,In_1975,In_653);
nor U481 (N_481,In_958,In_1130);
and U482 (N_482,In_1406,In_772);
nand U483 (N_483,In_1143,In_1479);
or U484 (N_484,In_1218,In_1097);
xnor U485 (N_485,In_2230,In_395);
xor U486 (N_486,In_1457,In_2083);
or U487 (N_487,In_1067,In_2444);
nand U488 (N_488,In_946,In_1532);
xnor U489 (N_489,In_1497,In_113);
xnor U490 (N_490,In_376,In_1176);
xnor U491 (N_491,In_924,In_2393);
nand U492 (N_492,In_713,In_2468);
nor U493 (N_493,In_594,In_1284);
xnor U494 (N_494,In_1550,In_2243);
and U495 (N_495,In_797,In_1293);
or U496 (N_496,In_514,In_1148);
and U497 (N_497,In_179,In_1692);
and U498 (N_498,In_775,In_232);
xor U499 (N_499,In_1972,In_1551);
nand U500 (N_500,In_116,In_2110);
xor U501 (N_501,In_452,In_1797);
and U502 (N_502,In_2492,In_2311);
nand U503 (N_503,In_2498,In_13);
or U504 (N_504,In_520,In_2048);
nand U505 (N_505,In_541,In_951);
nand U506 (N_506,In_1300,In_2476);
nor U507 (N_507,In_675,In_1731);
and U508 (N_508,In_1825,In_407);
nand U509 (N_509,In_2077,In_1980);
and U510 (N_510,In_877,In_377);
nand U511 (N_511,In_1048,In_563);
or U512 (N_512,In_854,In_1703);
nor U513 (N_513,In_1968,In_2367);
and U514 (N_514,In_605,In_1166);
xor U515 (N_515,In_2097,In_1075);
xor U516 (N_516,In_2132,In_98);
nand U517 (N_517,In_2418,In_1544);
and U518 (N_518,In_2189,In_560);
xor U519 (N_519,In_633,In_2042);
nand U520 (N_520,In_1535,In_277);
xnor U521 (N_521,In_1988,In_2053);
nor U522 (N_522,In_37,In_2037);
or U523 (N_523,In_2234,In_1803);
nand U524 (N_524,In_1496,In_2262);
or U525 (N_525,In_1646,In_706);
xor U526 (N_526,In_2296,In_416);
xnor U527 (N_527,In_351,In_2025);
or U528 (N_528,In_1605,In_2263);
nor U529 (N_529,In_324,In_0);
or U530 (N_530,In_968,In_1064);
xnor U531 (N_531,In_1220,In_1307);
and U532 (N_532,In_1415,In_434);
xnor U533 (N_533,In_1781,In_1192);
nand U534 (N_534,In_1753,In_1420);
nor U535 (N_535,In_51,In_81);
or U536 (N_536,In_228,In_2337);
nand U537 (N_537,In_2228,In_1387);
and U538 (N_538,In_1258,In_787);
and U539 (N_539,In_2207,In_1488);
and U540 (N_540,In_1495,In_523);
or U541 (N_541,In_879,In_223);
or U542 (N_542,In_142,In_186);
or U543 (N_543,In_135,In_2089);
nand U544 (N_544,In_259,In_1295);
and U545 (N_545,In_1404,In_1439);
nor U546 (N_546,In_1386,In_1400);
nand U547 (N_547,In_1920,In_87);
or U548 (N_548,In_881,In_1308);
xor U549 (N_549,In_2186,In_799);
and U550 (N_550,In_206,In_1071);
and U551 (N_551,In_1046,In_565);
nor U552 (N_552,In_263,In_1155);
nor U553 (N_553,In_1950,In_2409);
nand U554 (N_554,In_2495,In_1394);
nor U555 (N_555,In_1152,In_1902);
xnor U556 (N_556,In_26,In_949);
or U557 (N_557,In_275,In_583);
nor U558 (N_558,In_1896,In_901);
and U559 (N_559,In_2381,In_2412);
xor U560 (N_560,In_1734,In_2064);
xnor U561 (N_561,In_696,In_1571);
xor U562 (N_562,In_337,In_1004);
or U563 (N_563,In_2222,In_1831);
xnor U564 (N_564,In_1584,In_2123);
or U565 (N_565,In_14,In_757);
xnor U566 (N_566,In_571,In_2047);
or U567 (N_567,In_934,In_559);
and U568 (N_568,In_970,In_988);
nand U569 (N_569,In_735,In_2415);
xor U570 (N_570,In_1898,In_2013);
or U571 (N_571,In_2406,In_2193);
xor U572 (N_572,In_1900,In_325);
nand U573 (N_573,In_2044,In_2106);
and U574 (N_574,In_744,In_516);
and U575 (N_575,In_1095,In_2241);
nor U576 (N_576,In_788,In_983);
and U577 (N_577,In_1,In_1036);
and U578 (N_578,In_1567,In_2292);
or U579 (N_579,In_664,In_1591);
and U580 (N_580,In_795,In_1065);
nor U581 (N_581,In_538,In_1149);
xnor U582 (N_582,In_1615,In_1624);
xnor U583 (N_583,In_1294,In_1984);
xnor U584 (N_584,In_2429,In_129);
nor U585 (N_585,In_1306,In_1811);
and U586 (N_586,In_1119,In_1773);
xor U587 (N_587,In_90,In_1504);
or U588 (N_588,In_137,In_1321);
nand U589 (N_589,In_2071,In_2020);
and U590 (N_590,In_699,In_1832);
and U591 (N_591,In_1271,In_1206);
or U592 (N_592,In_1471,In_280);
nor U593 (N_593,In_335,In_242);
and U594 (N_594,In_1517,In_1893);
or U595 (N_595,In_1678,In_2039);
and U596 (N_596,In_1746,In_1492);
nand U597 (N_597,In_289,In_2105);
nand U598 (N_598,In_165,In_2206);
and U599 (N_599,In_1270,In_1147);
and U600 (N_600,In_897,In_1291);
xor U601 (N_601,In_912,In_1216);
or U602 (N_602,In_1296,In_2281);
nor U603 (N_603,In_279,In_2469);
nand U604 (N_604,In_880,In_368);
nor U605 (N_605,In_1398,In_1648);
xnor U606 (N_606,In_140,In_1697);
nor U607 (N_607,In_866,In_971);
nor U608 (N_608,In_1679,In_2054);
xnor U609 (N_609,In_1782,In_810);
nor U610 (N_610,In_643,In_2016);
nand U611 (N_611,In_627,In_182);
nand U612 (N_612,In_503,In_1677);
nand U613 (N_613,In_2136,In_1938);
nand U614 (N_614,In_1816,In_2115);
xnor U615 (N_615,In_493,In_1861);
xnor U616 (N_616,In_1247,In_1742);
xnor U617 (N_617,In_950,In_1332);
nand U618 (N_618,In_2116,In_1545);
xnor U619 (N_619,In_1978,In_1225);
and U620 (N_620,In_1992,In_2052);
xor U621 (N_621,In_331,In_318);
xnor U622 (N_622,In_471,In_978);
or U623 (N_623,In_1965,In_549);
and U624 (N_624,In_60,In_2062);
nor U625 (N_625,In_1857,In_2141);
or U626 (N_626,In_1955,In_2000);
xor U627 (N_627,In_487,In_959);
nor U628 (N_628,In_1585,In_648);
and U629 (N_629,In_1583,In_691);
or U630 (N_630,In_2246,In_1135);
nand U631 (N_631,In_2108,In_498);
nor U632 (N_632,In_2172,In_1830);
or U633 (N_633,In_1158,In_52);
nor U634 (N_634,In_1741,In_267);
nand U635 (N_635,In_576,In_240);
or U636 (N_636,In_501,In_195);
and U637 (N_637,In_1348,In_2142);
nor U638 (N_638,In_1963,In_365);
nand U639 (N_639,In_2114,In_1474);
nand U640 (N_640,In_489,In_1467);
xnor U641 (N_641,In_892,In_550);
nor U642 (N_642,In_2085,In_589);
nor U643 (N_643,In_2377,In_1635);
nand U644 (N_644,In_1879,In_2462);
and U645 (N_645,In_2328,In_846);
xnor U646 (N_646,In_2438,In_928);
nand U647 (N_647,In_759,In_2144);
or U648 (N_648,In_677,In_2303);
and U649 (N_649,In_956,In_423);
and U650 (N_650,In_204,In_2088);
nor U651 (N_651,In_2149,In_995);
xnor U652 (N_652,In_190,In_817);
nand U653 (N_653,In_1328,In_1749);
xnor U654 (N_654,In_2103,In_792);
xor U655 (N_655,In_421,In_1913);
nand U656 (N_656,In_68,In_1402);
and U657 (N_657,In_196,In_1355);
xnor U658 (N_658,In_1817,In_814);
nor U659 (N_659,In_793,In_1233);
or U660 (N_660,In_1085,In_1112);
or U661 (N_661,In_1512,In_1414);
nand U662 (N_662,In_1958,In_1794);
and U663 (N_663,In_2389,In_965);
and U664 (N_664,In_1882,In_893);
and U665 (N_665,In_2387,In_209);
and U666 (N_666,In_836,In_1034);
xnor U667 (N_667,In_1054,In_2421);
or U668 (N_668,In_2036,In_2380);
and U669 (N_669,In_982,In_139);
nand U670 (N_670,In_1923,In_1359);
nand U671 (N_671,In_900,In_1117);
or U672 (N_672,In_990,In_198);
xor U673 (N_673,In_2273,In_1770);
nand U674 (N_674,In_1777,In_1855);
xor U675 (N_675,In_2161,In_2478);
xnor U676 (N_676,In_1688,In_211);
nand U677 (N_677,In_1447,In_1283);
xnor U678 (N_678,In_2202,In_205);
xnor U679 (N_679,In_397,In_575);
or U680 (N_680,In_427,In_2094);
nand U681 (N_681,In_1943,In_2022);
nand U682 (N_682,In_1165,In_251);
xor U683 (N_683,In_366,In_2153);
nand U684 (N_684,In_967,In_2314);
or U685 (N_685,In_884,In_2279);
nand U686 (N_686,In_1316,In_353);
or U687 (N_687,In_749,In_1505);
or U688 (N_688,In_392,In_567);
xnor U689 (N_689,In_157,In_1061);
nand U690 (N_690,In_2196,In_730);
xor U691 (N_691,In_1163,In_1863);
nand U692 (N_692,In_2148,In_1775);
or U693 (N_693,In_1866,In_1371);
or U694 (N_694,In_596,In_2497);
nand U695 (N_695,In_1693,In_606);
xor U696 (N_696,In_163,In_937);
nand U697 (N_697,In_1172,In_2129);
and U698 (N_698,In_883,In_2432);
nand U699 (N_699,In_1377,In_74);
or U700 (N_700,In_1574,In_2101);
xnor U701 (N_701,In_500,In_2038);
nand U702 (N_702,In_202,In_1657);
xnor U703 (N_703,In_1700,In_127);
nand U704 (N_704,In_2130,In_1173);
nor U705 (N_705,In_570,In_993);
nand U706 (N_706,In_2261,In_1981);
and U707 (N_707,In_1600,In_1909);
or U708 (N_708,In_1436,In_411);
nand U709 (N_709,In_723,In_1047);
nand U710 (N_710,In_1168,In_361);
nand U711 (N_711,In_66,In_1428);
and U712 (N_712,In_1120,In_2035);
or U713 (N_713,In_483,In_1418);
nand U714 (N_714,In_1764,In_832);
nand U715 (N_715,In_1249,In_927);
or U716 (N_716,In_199,In_1719);
or U717 (N_717,In_621,In_1050);
xnor U718 (N_718,In_1998,In_1695);
xor U719 (N_719,In_1986,In_1889);
nor U720 (N_720,In_1450,In_1442);
nor U721 (N_721,In_125,In_1995);
and U722 (N_722,In_1214,In_1887);
xnor U723 (N_723,In_2240,In_1408);
nor U724 (N_724,In_1809,In_1171);
nand U725 (N_725,In_2274,In_1827);
or U726 (N_726,In_2111,In_1518);
xor U727 (N_727,In_2358,In_1503);
nand U728 (N_728,In_535,In_998);
nor U729 (N_729,In_1645,In_285);
and U730 (N_730,In_2119,In_918);
xnor U731 (N_731,In_2139,In_1014);
nor U732 (N_732,In_1421,In_286);
nor U733 (N_733,In_821,In_2055);
and U734 (N_734,In_350,In_1059);
nor U735 (N_735,In_1412,In_1489);
xor U736 (N_736,In_2336,In_1735);
xnor U737 (N_737,In_1088,In_433);
and U738 (N_738,In_598,In_1873);
nor U739 (N_739,In_1824,In_1290);
and U740 (N_740,In_1837,In_710);
xor U741 (N_741,In_604,In_1486);
nor U742 (N_742,In_403,In_1589);
xnor U743 (N_743,In_1548,In_1951);
nand U744 (N_744,In_915,In_1751);
nand U745 (N_745,In_2306,In_1702);
xor U746 (N_746,In_1299,In_2291);
nor U747 (N_747,In_919,In_1093);
and U748 (N_748,In_518,In_1977);
nand U749 (N_749,In_1385,In_143);
nor U750 (N_750,In_2471,In_170);
xnor U751 (N_751,In_1069,In_1025);
nor U752 (N_752,In_704,In_1631);
nor U753 (N_753,In_1219,In_1562);
nand U754 (N_754,In_58,In_679);
and U755 (N_755,In_1941,In_1259);
nor U756 (N_756,In_943,In_1285);
and U757 (N_757,In_1647,In_670);
xnor U758 (N_758,In_54,In_1627);
xnor U759 (N_759,In_2109,In_1388);
nand U760 (N_760,In_1946,In_830);
and U761 (N_761,In_1971,In_2072);
nand U762 (N_762,In_2449,In_1126);
xor U763 (N_763,In_492,In_865);
and U764 (N_764,In_818,In_358);
and U765 (N_765,In_1691,In_244);
nand U766 (N_766,In_4,In_355);
or U767 (N_767,In_1121,In_1066);
and U768 (N_768,In_587,In_1686);
nand U769 (N_769,In_1462,In_655);
or U770 (N_770,In_255,In_2070);
nor U771 (N_771,In_2351,In_1243);
nor U772 (N_772,In_603,In_1187);
nor U773 (N_773,In_999,In_362);
nor U774 (N_774,In_2425,In_2319);
nand U775 (N_775,In_394,In_300);
and U776 (N_776,In_805,In_62);
or U777 (N_777,In_2209,In_1363);
xnor U778 (N_778,In_1310,In_806);
nor U779 (N_779,In_2297,In_1315);
and U780 (N_780,In_1430,In_515);
and U781 (N_781,In_238,In_533);
nand U782 (N_782,In_957,In_629);
or U783 (N_783,In_1554,In_932);
nand U784 (N_784,In_2402,In_907);
xnor U785 (N_785,In_1822,In_265);
nor U786 (N_786,In_121,In_1407);
nor U787 (N_787,In_258,In_734);
xnor U788 (N_788,In_1401,In_2346);
and U789 (N_789,In_1966,In_963);
nand U790 (N_790,In_1006,In_107);
nand U791 (N_791,In_2400,In_1035);
and U792 (N_792,In_2433,In_1223);
nand U793 (N_793,In_1012,In_1523);
nor U794 (N_794,In_472,In_71);
xor U795 (N_795,In_20,In_1434);
nor U796 (N_796,In_1833,In_36);
xor U797 (N_797,In_2446,In_2283);
xor U798 (N_798,In_1839,In_1829);
xor U799 (N_799,In_2081,In_933);
nand U800 (N_800,In_1515,In_847);
nand U801 (N_801,In_2448,In_338);
or U802 (N_802,In_558,In_1157);
or U803 (N_803,In_1397,In_2399);
nor U804 (N_804,In_1560,In_1498);
xor U805 (N_805,In_1125,In_253);
or U806 (N_806,In_1918,In_2335);
and U807 (N_807,In_1267,In_2390);
xnor U808 (N_808,In_1287,In_252);
and U809 (N_809,In_1501,In_613);
and U810 (N_810,In_1372,In_502);
xnor U811 (N_811,In_1018,In_2173);
or U812 (N_812,In_1667,In_1003);
or U813 (N_813,In_2165,In_1451);
nand U814 (N_814,In_2164,In_417);
or U815 (N_815,In_1784,In_425);
nand U816 (N_816,In_2198,In_2401);
xor U817 (N_817,In_1821,In_1392);
nand U818 (N_818,In_1526,In_2147);
xnor U819 (N_819,In_320,In_1890);
and U820 (N_820,In_2254,In_1419);
nor U821 (N_821,In_2122,In_906);
and U822 (N_822,In_410,In_100);
xnor U823 (N_823,In_1265,In_1194);
xor U824 (N_824,In_1468,In_1027);
nand U825 (N_825,In_1186,In_641);
nor U826 (N_826,In_1289,In_1840);
nor U827 (N_827,In_1063,In_1443);
xnor U828 (N_828,In_1261,In_1791);
xnor U829 (N_829,In_602,In_389);
nand U830 (N_830,In_2231,In_1010);
xor U831 (N_831,In_1976,In_736);
and U832 (N_832,In_843,In_2133);
xnor U833 (N_833,In_354,In_2204);
nand U834 (N_834,In_870,In_694);
nand U835 (N_835,In_444,In_1883);
nand U836 (N_836,In_2477,In_1948);
nor U837 (N_837,In_112,In_972);
nor U838 (N_838,In_573,In_1726);
or U839 (N_839,In_1413,In_1949);
and U840 (N_840,In_84,In_378);
and U841 (N_841,In_1353,In_1942);
nor U842 (N_842,In_1272,In_909);
and U843 (N_843,In_548,In_2185);
and U844 (N_844,In_1182,In_1595);
or U845 (N_845,In_1892,In_1625);
xor U846 (N_846,In_826,In_1597);
or U847 (N_847,In_1579,In_1432);
or U848 (N_848,In_720,In_1044);
xor U849 (N_849,In_1763,In_1718);
or U850 (N_850,In_1038,In_1073);
nor U851 (N_851,In_402,In_448);
nor U852 (N_852,In_1643,In_2483);
and U853 (N_853,In_2339,In_1626);
nor U854 (N_854,In_2280,In_740);
nand U855 (N_855,In_230,In_1043);
and U856 (N_856,In_1876,In_418);
or U857 (N_857,In_1383,In_2247);
and U858 (N_858,In_2180,In_838);
and U859 (N_859,In_1002,In_2200);
or U860 (N_860,In_86,In_1188);
and U861 (N_861,In_551,In_1755);
xnor U862 (N_862,In_1633,In_820);
nand U863 (N_863,In_1834,In_1744);
and U864 (N_864,In_1826,In_2043);
nor U865 (N_865,In_1423,In_1382);
or U866 (N_866,In_2439,In_1273);
or U867 (N_867,In_349,In_1622);
and U868 (N_868,In_680,In_895);
and U869 (N_869,In_649,In_2152);
xnor U870 (N_870,In_896,In_291);
nor U871 (N_871,In_1527,In_67);
nand U872 (N_872,In_380,In_1860);
xnor U873 (N_873,In_802,In_1339);
nor U874 (N_874,In_1235,In_739);
xor U875 (N_875,In_488,In_1612);
and U876 (N_876,In_1789,In_1245);
and U877 (N_877,In_293,In_2357);
xor U878 (N_878,In_97,In_784);
or U879 (N_879,In_55,In_175);
nand U880 (N_880,In_2060,In_1878);
xnor U881 (N_881,In_1928,In_1009);
nand U882 (N_882,In_247,In_2414);
nor U883 (N_883,In_617,In_1373);
xor U884 (N_884,In_1352,In_1536);
or U885 (N_885,In_2223,In_2235);
nand U886 (N_886,In_134,In_304);
or U887 (N_887,In_1628,In_364);
nor U888 (N_888,In_1260,In_1877);
xor U889 (N_889,In_2259,In_754);
xnor U890 (N_890,In_752,In_1549);
nand U891 (N_891,In_2056,In_404);
and U892 (N_892,In_1774,In_2082);
xnor U893 (N_893,In_2049,In_1974);
xnor U894 (N_894,In_2178,In_470);
or U895 (N_895,In_1769,In_1576);
nor U896 (N_896,In_916,In_2251);
and U897 (N_897,In_964,In_2159);
or U898 (N_898,In_1683,In_923);
or U899 (N_899,In_147,In_1380);
nand U900 (N_900,In_966,In_119);
nor U901 (N_901,In_429,In_387);
nor U902 (N_902,In_1926,In_2102);
xor U903 (N_903,In_457,In_1251);
and U904 (N_904,In_878,In_2066);
xor U905 (N_905,In_1141,In_191);
or U906 (N_906,In_2242,In_2171);
or U907 (N_907,In_1778,In_76);
nand U908 (N_908,In_1637,In_1269);
xnor U909 (N_909,In_477,In_1354);
and U910 (N_910,In_73,In_651);
nor U911 (N_911,In_2408,In_172);
nor U912 (N_912,In_1853,In_1279);
nand U913 (N_913,In_2317,In_464);
or U914 (N_914,In_1709,In_552);
and U915 (N_915,In_193,In_308);
nor U916 (N_916,In_689,In_1592);
xor U917 (N_917,In_2029,In_1490);
xnor U918 (N_918,In_1327,In_2211);
or U919 (N_919,In_822,In_227);
nor U920 (N_920,In_556,In_122);
or U921 (N_921,In_2396,In_2383);
and U922 (N_922,In_138,In_1556);
nand U923 (N_923,In_1952,In_384);
or U924 (N_924,In_1519,In_1650);
nor U925 (N_925,In_1349,In_764);
and U926 (N_926,In_1671,In_825);
nor U927 (N_927,In_1076,In_102);
and U928 (N_928,In_1618,In_1091);
nand U929 (N_929,In_1566,In_1281);
xor U930 (N_930,In_1908,In_1947);
nand U931 (N_931,In_640,In_145);
nand U932 (N_932,In_108,In_1553);
xor U933 (N_933,In_2484,In_1081);
or U934 (N_934,In_12,In_2079);
and U935 (N_935,In_1092,In_662);
nor U936 (N_936,In_2191,In_1785);
nand U937 (N_937,In_2021,In_1395);
xnor U938 (N_938,In_2050,In_2324);
nor U939 (N_939,In_1362,In_1277);
xor U940 (N_940,In_169,In_1738);
xor U941 (N_941,In_1708,In_340);
and U942 (N_942,In_2294,In_858);
or U943 (N_943,In_712,In_1106);
nor U944 (N_944,In_1901,In_921);
or U945 (N_945,In_1636,In_1669);
or U946 (N_946,In_1464,In_898);
xor U947 (N_947,In_980,In_1335);
nand U948 (N_948,In_945,In_2120);
nor U949 (N_949,In_2286,In_401);
or U950 (N_950,In_1848,In_616);
nor U951 (N_951,In_2454,In_1274);
nand U952 (N_952,In_109,In_2096);
nand U953 (N_953,In_1886,In_1836);
or U954 (N_954,In_144,In_2447);
nand U955 (N_955,In_1409,In_2008);
and U956 (N_956,In_485,In_2113);
and U957 (N_957,In_714,In_1317);
nand U958 (N_958,In_96,In_1305);
or U959 (N_959,In_50,In_1017);
xnor U960 (N_960,In_1425,In_301);
or U961 (N_961,In_1684,In_2416);
and U962 (N_962,In_1449,In_984);
nor U963 (N_963,In_2232,In_266);
nor U964 (N_964,In_379,In_2386);
xor U965 (N_965,In_1559,In_1202);
nand U966 (N_966,In_2256,In_1100);
and U967 (N_967,In_868,In_1655);
nor U968 (N_968,In_673,In_1275);
and U969 (N_969,In_1743,In_1116);
or U970 (N_970,In_332,In_1634);
and U971 (N_971,In_1153,In_2140);
or U972 (N_972,In_2481,In_1199);
or U973 (N_973,In_465,In_1593);
xor U974 (N_974,In_1569,In_481);
and U975 (N_975,In_359,In_1509);
or U976 (N_976,In_1446,In_1115);
nor U977 (N_977,In_110,In_1795);
nand U978 (N_978,In_390,In_601);
and U979 (N_979,In_661,In_2388);
and U980 (N_980,In_609,In_1189);
nor U981 (N_981,In_1710,In_790);
or U982 (N_982,In_845,In_2248);
or U983 (N_983,In_1282,In_2250);
and U984 (N_984,In_742,In_709);
or U985 (N_985,In_234,In_346);
and U986 (N_986,In_2095,In_2068);
nand U987 (N_987,In_2445,In_719);
xnor U988 (N_988,In_1905,In_1019);
nand U989 (N_989,In_2474,In_2300);
nor U990 (N_990,In_1229,In_766);
nand U991 (N_991,In_1207,In_2343);
nand U992 (N_992,In_1110,In_1337);
xor U993 (N_993,In_1231,In_2131);
nand U994 (N_994,In_1396,In_920);
xnor U995 (N_995,In_1242,In_428);
and U996 (N_996,In_1292,In_1929);
nor U997 (N_997,In_154,In_566);
xnor U998 (N_998,In_647,In_85);
xor U999 (N_999,In_386,In_1311);
xnor U1000 (N_1000,In_2320,In_8);
nor U1001 (N_1001,In_1020,In_2354);
and U1002 (N_1002,In_25,In_38);
or U1003 (N_1003,In_1897,In_542);
xnor U1004 (N_1004,In_1179,In_2301);
nand U1005 (N_1005,In_409,In_197);
or U1006 (N_1006,In_2086,In_2004);
nand U1007 (N_1007,In_996,In_136);
nor U1008 (N_1008,In_2018,In_1874);
or U1009 (N_1009,In_1639,In_808);
nand U1010 (N_1010,In_171,In_1084);
and U1011 (N_1011,In_229,In_1487);
nand U1012 (N_1012,In_2370,In_842);
xor U1013 (N_1013,In_1990,In_1582);
or U1014 (N_1014,In_374,In_2076);
or U1015 (N_1015,In_1854,In_1531);
nand U1016 (N_1016,In_1932,In_2168);
nand U1017 (N_1017,In_256,In_219);
nor U1018 (N_1018,In_568,In_313);
and U1019 (N_1019,In_430,In_53);
xnor U1020 (N_1020,In_737,In_2058);
xnor U1021 (N_1021,In_459,In_458);
and U1022 (N_1022,In_874,In_1944);
and U1023 (N_1023,In_637,In_2009);
or U1024 (N_1024,In_43,In_2391);
nor U1025 (N_1025,In_1808,In_225);
xor U1026 (N_1026,In_1215,In_1180);
xor U1027 (N_1027,In_2146,In_572);
nand U1028 (N_1028,In_1903,In_1875);
nor U1029 (N_1029,In_667,In_997);
nand U1030 (N_1030,In_773,In_78);
xor U1031 (N_1031,In_1641,In_1638);
and U1032 (N_1032,In_2413,In_2385);
nor U1033 (N_1033,In_220,In_1128);
nand U1034 (N_1034,In_1514,In_1540);
and U1035 (N_1035,In_49,In_562);
nand U1036 (N_1036,In_582,In_786);
xor U1037 (N_1037,In_717,In_1969);
nand U1038 (N_1038,In_2216,In_885);
nand U1039 (N_1039,In_1601,In_310);
nor U1040 (N_1040,In_1078,In_1197);
nor U1041 (N_1041,In_1933,In_1606);
and U1042 (N_1042,In_160,In_595);
or U1043 (N_1043,In_72,In_989);
or U1044 (N_1044,In_1766,In_1351);
and U1045 (N_1045,In_1783,In_2112);
and U1046 (N_1046,In_2217,In_2197);
nor U1047 (N_1047,In_1555,In_811);
and U1048 (N_1048,In_2431,In_201);
nand U1049 (N_1049,In_1136,In_1640);
or U1050 (N_1050,In_1350,In_981);
or U1051 (N_1051,In_23,In_385);
or U1052 (N_1052,In_1970,In_2065);
xnor U1053 (N_1053,In_56,In_2233);
or U1054 (N_1054,In_2158,In_992);
xnor U1055 (N_1055,In_2156,In_1123);
and U1056 (N_1056,In_2341,In_2221);
nand U1057 (N_1057,In_445,In_2470);
or U1058 (N_1058,In_454,In_34);
xnor U1059 (N_1059,In_686,In_1431);
and U1060 (N_1060,In_1103,In_1268);
nand U1061 (N_1061,In_192,In_2436);
xor U1062 (N_1062,In_1757,In_2267);
or U1063 (N_1063,In_2026,In_1868);
xor U1064 (N_1064,In_612,In_453);
and U1065 (N_1065,In_491,In_1689);
nor U1066 (N_1066,In_2032,In_77);
or U1067 (N_1067,In_1665,In_1326);
xnor U1068 (N_1068,In_2028,In_692);
xnor U1069 (N_1069,In_2182,In_305);
or U1070 (N_1070,In_2352,In_284);
nand U1071 (N_1071,In_1405,In_1437);
nand U1072 (N_1072,In_1493,In_1630);
xor U1073 (N_1073,In_1099,In_1114);
nand U1074 (N_1074,In_360,In_1040);
nor U1075 (N_1075,In_763,In_1074);
nor U1076 (N_1076,In_2480,In_777);
and U1077 (N_1077,In_2006,In_185);
nand U1078 (N_1078,In_1309,In_299);
and U1079 (N_1079,In_1096,In_370);
and U1080 (N_1080,In_2134,In_726);
nor U1081 (N_1081,In_580,In_910);
nand U1082 (N_1082,In_1761,In_2479);
nor U1083 (N_1083,In_2074,In_1663);
and U1084 (N_1084,In_2284,In_89);
xor U1085 (N_1085,In_1713,In_1368);
xor U1086 (N_1086,In_1087,In_2023);
and U1087 (N_1087,In_632,In_1484);
nand U1088 (N_1088,In_2310,In_929);
nor U1089 (N_1089,In_973,In_630);
nand U1090 (N_1090,In_1237,In_375);
and U1091 (N_1091,In_1041,In_695);
and U1092 (N_1092,In_1748,In_2205);
and U1093 (N_1093,In_728,In_367);
nand U1094 (N_1094,In_1510,In_398);
or U1095 (N_1095,In_1185,In_610);
or U1096 (N_1096,In_1411,In_1524);
or U1097 (N_1097,In_1661,In_2);
nor U1098 (N_1098,In_903,In_1477);
nand U1099 (N_1099,In_2329,In_1629);
nand U1100 (N_1100,In_1989,In_506);
nand U1101 (N_1101,In_262,In_30);
and U1102 (N_1102,In_2269,In_2472);
nand U1103 (N_1103,In_1732,In_2423);
nor U1104 (N_1104,In_1445,In_827);
nand U1105 (N_1105,In_975,In_2322);
nor U1106 (N_1106,In_131,In_1740);
and U1107 (N_1107,In_1961,In_462);
xor U1108 (N_1108,In_622,In_2266);
or U1109 (N_1109,In_302,In_184);
and U1110 (N_1110,In_343,In_861);
and U1111 (N_1111,In_642,In_1236);
nand U1112 (N_1112,In_1619,In_682);
and U1113 (N_1113,In_1028,In_245);
and U1114 (N_1114,In_769,In_314);
xnor U1115 (N_1115,In_31,In_1658);
and U1116 (N_1116,In_111,In_2163);
nand U1117 (N_1117,In_1577,In_976);
and U1118 (N_1118,In_1072,In_173);
nand U1119 (N_1119,In_652,In_511);
or U1120 (N_1120,In_2489,In_904);
nor U1121 (N_1121,In_955,In_1771);
nor U1122 (N_1122,In_396,In_1361);
nand U1123 (N_1123,In_115,In_2169);
nand U1124 (N_1124,In_851,In_688);
or U1125 (N_1125,In_1357,In_1473);
or U1126 (N_1126,In_1581,In_2293);
xor U1127 (N_1127,In_2422,In_1297);
xnor U1128 (N_1128,In_180,In_1779);
nor U1129 (N_1129,In_886,In_2199);
xor U1130 (N_1130,In_1239,In_2041);
nand U1131 (N_1131,In_2375,In_480);
and U1132 (N_1132,In_926,In_450);
nand U1133 (N_1133,In_1960,In_1253);
nor U1134 (N_1134,In_207,In_1568);
nor U1135 (N_1135,In_1124,In_1393);
or U1136 (N_1136,In_994,In_1870);
and U1137 (N_1137,In_747,In_1314);
and U1138 (N_1138,In_449,In_312);
nor U1139 (N_1139,In_1459,In_782);
or U1140 (N_1140,In_132,In_1564);
xor U1141 (N_1141,In_1715,In_1276);
and U1142 (N_1142,In_2061,In_322);
and U1143 (N_1143,In_39,In_1727);
or U1144 (N_1144,In_2372,In_961);
nand U1145 (N_1145,In_2104,In_508);
nand U1146 (N_1146,In_311,In_2194);
nand U1147 (N_1147,In_391,In_435);
nor U1148 (N_1148,In_413,In_1280);
nor U1149 (N_1149,In_581,In_1263);
or U1150 (N_1150,In_1642,In_765);
and U1151 (N_1151,In_2458,In_446);
xnor U1152 (N_1152,In_1934,In_1347);
nor U1153 (N_1153,In_176,In_2355);
xor U1154 (N_1154,In_2151,In_2051);
and U1155 (N_1155,In_1810,In_1993);
nand U1156 (N_1156,In_1676,In_776);
and U1157 (N_1157,In_703,In_1907);
or U1158 (N_1158,In_1052,In_1470);
nor U1159 (N_1159,In_1945,In_564);
and U1160 (N_1160,In_91,In_741);
nor U1161 (N_1161,In_1336,In_1089);
or U1162 (N_1162,In_751,In_828);
nand U1163 (N_1163,In_1319,In_2275);
nand U1164 (N_1164,In_2298,In_2407);
nor U1165 (N_1165,In_1154,In_939);
or U1166 (N_1166,In_92,In_2434);
nor U1167 (N_1167,In_681,In_1461);
or U1168 (N_1168,In_665,In_1252);
nor U1169 (N_1169,In_2459,In_9);
nand U1170 (N_1170,In_436,In_463);
nand U1171 (N_1171,In_1916,In_1580);
xor U1172 (N_1172,In_1935,In_803);
xor U1173 (N_1173,In_2046,In_748);
nand U1174 (N_1174,In_1118,In_2441);
nand U1175 (N_1175,In_1191,In_1588);
nor U1176 (N_1176,In_1558,In_2024);
xnor U1177 (N_1177,In_2289,In_561);
xnor U1178 (N_1178,In_1033,In_226);
nand U1179 (N_1179,In_743,In_716);
xnor U1180 (N_1180,In_1049,In_2187);
nand U1181 (N_1181,In_1491,In_326);
nand U1182 (N_1182,In_2220,In_2344);
xnor U1183 (N_1183,In_2244,In_1381);
nand U1184 (N_1184,In_698,In_863);
or U1185 (N_1185,In_1675,In_2007);
or U1186 (N_1186,In_1904,In_1919);
nand U1187 (N_1187,In_2239,In_1248);
nand U1188 (N_1188,In_2392,In_745);
and U1189 (N_1189,In_1722,In_2190);
and U1190 (N_1190,In_369,In_543);
or U1191 (N_1191,In_33,In_1433);
nand U1192 (N_1192,In_687,In_1862);
xnor U1193 (N_1193,In_1575,In_586);
xor U1194 (N_1194,In_2466,In_2333);
and U1195 (N_1195,In_725,In_419);
or U1196 (N_1196,In_32,In_931);
nor U1197 (N_1197,In_45,In_1776);
xor U1198 (N_1198,In_1728,In_1145);
xnor U1199 (N_1199,In_1823,In_674);
and U1200 (N_1200,In_1222,In_2302);
xor U1201 (N_1201,In_2078,In_2276);
or U1202 (N_1202,In_2126,In_1499);
or U1203 (N_1203,In_177,In_2403);
nand U1204 (N_1204,In_2045,In_1005);
nand U1205 (N_1205,In_150,In_1032);
or U1206 (N_1206,In_1342,In_1083);
and U1207 (N_1207,In_894,In_1733);
or U1208 (N_1208,In_2486,In_2360);
nand U1209 (N_1209,In_1122,In_2090);
nor U1210 (N_1210,In_708,In_669);
nor U1211 (N_1211,In_569,In_2456);
and U1212 (N_1212,In_1572,In_400);
xnor U1213 (N_1213,In_1101,In_114);
nand U1214 (N_1214,In_578,In_1264);
nand U1215 (N_1215,In_1108,In_1937);
or U1216 (N_1216,In_899,In_257);
nand U1217 (N_1217,In_1864,In_834);
nor U1218 (N_1218,In_2059,In_2121);
xor U1219 (N_1219,In_1930,In_1894);
nand U1220 (N_1220,In_1659,In_24);
xor U1221 (N_1221,In_1511,In_2315);
and U1222 (N_1222,In_2192,In_1195);
or U1223 (N_1223,In_2290,In_414);
and U1224 (N_1224,In_1712,In_1162);
nand U1225 (N_1225,In_840,In_348);
nand U1226 (N_1226,In_2366,In_1338);
nand U1227 (N_1227,In_676,In_2145);
nand U1228 (N_1228,In_1058,In_614);
nor U1229 (N_1229,In_1956,In_672);
xor U1230 (N_1230,In_1142,In_758);
or U1231 (N_1231,In_1787,In_1608);
nor U1232 (N_1232,In_1842,In_117);
and U1233 (N_1233,In_1196,In_2485);
nand U1234 (N_1234,In_2326,In_1205);
xor U1235 (N_1235,In_1542,In_1080);
xnor U1236 (N_1236,In_611,In_272);
or U1237 (N_1237,In_194,In_1238);
nand U1238 (N_1238,In_1666,In_1673);
and U1239 (N_1239,In_1720,In_526);
or U1240 (N_1240,In_791,In_2287);
nand U1241 (N_1241,In_2318,In_2340);
and U1242 (N_1242,In_75,In_268);
nand U1243 (N_1243,In_1865,In_1170);
and U1244 (N_1244,In_938,In_1610);
nand U1245 (N_1245,In_1481,In_381);
and U1246 (N_1246,In_297,In_2460);
and U1247 (N_1247,In_250,In_2350);
xnor U1248 (N_1248,In_94,In_1983);
or U1249 (N_1249,In_1508,In_1384);
xor U1250 (N_1250,In_2323,In_1589);
and U1251 (N_1251,In_1912,In_1008);
nand U1252 (N_1252,In_128,In_2046);
nand U1253 (N_1253,In_2312,In_451);
and U1254 (N_1254,In_1311,In_1158);
xnor U1255 (N_1255,In_2176,In_2047);
and U1256 (N_1256,In_588,In_1724);
nor U1257 (N_1257,In_1593,In_1533);
or U1258 (N_1258,In_1191,In_528);
and U1259 (N_1259,In_569,In_302);
xor U1260 (N_1260,In_970,In_1792);
and U1261 (N_1261,In_2123,In_183);
nor U1262 (N_1262,In_880,In_1503);
or U1263 (N_1263,In_1878,In_1187);
xor U1264 (N_1264,In_342,In_43);
xor U1265 (N_1265,In_106,In_1753);
or U1266 (N_1266,In_1639,In_209);
nor U1267 (N_1267,In_352,In_1942);
or U1268 (N_1268,In_2116,In_1277);
and U1269 (N_1269,In_1938,In_2143);
nand U1270 (N_1270,In_2293,In_922);
xor U1271 (N_1271,In_1793,In_1645);
nor U1272 (N_1272,In_1663,In_1933);
xor U1273 (N_1273,In_174,In_1113);
or U1274 (N_1274,In_2036,In_1666);
nand U1275 (N_1275,In_534,In_1362);
nand U1276 (N_1276,In_1000,In_43);
xor U1277 (N_1277,In_1719,In_1931);
nand U1278 (N_1278,In_1303,In_1767);
nor U1279 (N_1279,In_1867,In_88);
and U1280 (N_1280,In_8,In_806);
nor U1281 (N_1281,In_1045,In_2423);
and U1282 (N_1282,In_1495,In_535);
or U1283 (N_1283,In_2009,In_239);
xor U1284 (N_1284,In_1544,In_1333);
nand U1285 (N_1285,In_2159,In_1309);
xnor U1286 (N_1286,In_2425,In_2041);
xnor U1287 (N_1287,In_576,In_1632);
nand U1288 (N_1288,In_943,In_1338);
nor U1289 (N_1289,In_2078,In_844);
or U1290 (N_1290,In_248,In_1273);
xnor U1291 (N_1291,In_84,In_2019);
nor U1292 (N_1292,In_2470,In_2378);
nor U1293 (N_1293,In_2252,In_272);
and U1294 (N_1294,In_273,In_1818);
and U1295 (N_1295,In_1811,In_2299);
nor U1296 (N_1296,In_941,In_503);
nor U1297 (N_1297,In_1385,In_2073);
xor U1298 (N_1298,In_1564,In_1010);
and U1299 (N_1299,In_679,In_390);
nor U1300 (N_1300,In_625,In_131);
or U1301 (N_1301,In_1370,In_1545);
xnor U1302 (N_1302,In_376,In_1384);
xnor U1303 (N_1303,In_1720,In_1954);
nand U1304 (N_1304,In_1967,In_1390);
nor U1305 (N_1305,In_1537,In_2005);
or U1306 (N_1306,In_325,In_1781);
and U1307 (N_1307,In_1626,In_701);
nand U1308 (N_1308,In_651,In_2378);
xnor U1309 (N_1309,In_1578,In_1941);
xnor U1310 (N_1310,In_657,In_1382);
or U1311 (N_1311,In_2430,In_2494);
or U1312 (N_1312,In_801,In_504);
and U1313 (N_1313,In_458,In_2130);
or U1314 (N_1314,In_2013,In_1644);
or U1315 (N_1315,In_1796,In_1174);
nand U1316 (N_1316,In_2468,In_2084);
xor U1317 (N_1317,In_2468,In_1185);
or U1318 (N_1318,In_616,In_634);
nor U1319 (N_1319,In_2339,In_1857);
and U1320 (N_1320,In_1874,In_1955);
xnor U1321 (N_1321,In_2304,In_499);
xor U1322 (N_1322,In_1690,In_1954);
and U1323 (N_1323,In_1424,In_45);
or U1324 (N_1324,In_1365,In_2067);
nand U1325 (N_1325,In_1311,In_260);
nand U1326 (N_1326,In_476,In_1016);
nor U1327 (N_1327,In_1378,In_2408);
nor U1328 (N_1328,In_2352,In_985);
nand U1329 (N_1329,In_1973,In_406);
nand U1330 (N_1330,In_106,In_2164);
or U1331 (N_1331,In_727,In_1103);
and U1332 (N_1332,In_2356,In_991);
and U1333 (N_1333,In_331,In_1072);
and U1334 (N_1334,In_899,In_30);
xnor U1335 (N_1335,In_22,In_1606);
nor U1336 (N_1336,In_627,In_2017);
or U1337 (N_1337,In_2374,In_2402);
nor U1338 (N_1338,In_1868,In_2130);
and U1339 (N_1339,In_469,In_2219);
nand U1340 (N_1340,In_1472,In_1841);
xor U1341 (N_1341,In_909,In_2326);
or U1342 (N_1342,In_1311,In_795);
and U1343 (N_1343,In_1830,In_860);
xnor U1344 (N_1344,In_2108,In_980);
xnor U1345 (N_1345,In_321,In_1921);
or U1346 (N_1346,In_1248,In_804);
xor U1347 (N_1347,In_1025,In_1765);
nand U1348 (N_1348,In_1051,In_2184);
nand U1349 (N_1349,In_333,In_1615);
nor U1350 (N_1350,In_47,In_1723);
or U1351 (N_1351,In_2146,In_1386);
or U1352 (N_1352,In_933,In_2109);
xnor U1353 (N_1353,In_2425,In_646);
nand U1354 (N_1354,In_1685,In_719);
xor U1355 (N_1355,In_924,In_2078);
nor U1356 (N_1356,In_1281,In_1800);
or U1357 (N_1357,In_2033,In_653);
and U1358 (N_1358,In_220,In_171);
and U1359 (N_1359,In_1134,In_2453);
or U1360 (N_1360,In_2337,In_166);
or U1361 (N_1361,In_1814,In_1190);
or U1362 (N_1362,In_986,In_987);
or U1363 (N_1363,In_2363,In_1364);
xor U1364 (N_1364,In_1788,In_262);
xor U1365 (N_1365,In_2341,In_919);
xnor U1366 (N_1366,In_1765,In_2157);
or U1367 (N_1367,In_755,In_816);
or U1368 (N_1368,In_917,In_101);
nor U1369 (N_1369,In_2241,In_463);
and U1370 (N_1370,In_438,In_543);
nor U1371 (N_1371,In_1871,In_1283);
and U1372 (N_1372,In_2314,In_1495);
nor U1373 (N_1373,In_968,In_1868);
nand U1374 (N_1374,In_1899,In_1051);
nor U1375 (N_1375,In_2353,In_81);
nor U1376 (N_1376,In_1361,In_2442);
or U1377 (N_1377,In_1798,In_1023);
and U1378 (N_1378,In_2496,In_2432);
nor U1379 (N_1379,In_1742,In_1726);
and U1380 (N_1380,In_556,In_1156);
or U1381 (N_1381,In_2175,In_2370);
nor U1382 (N_1382,In_2134,In_2405);
or U1383 (N_1383,In_1290,In_68);
or U1384 (N_1384,In_476,In_713);
nor U1385 (N_1385,In_536,In_511);
xor U1386 (N_1386,In_1183,In_92);
or U1387 (N_1387,In_2141,In_1969);
nor U1388 (N_1388,In_477,In_1318);
and U1389 (N_1389,In_2253,In_377);
xnor U1390 (N_1390,In_353,In_1845);
nand U1391 (N_1391,In_571,In_2338);
nand U1392 (N_1392,In_1582,In_1790);
nor U1393 (N_1393,In_1717,In_1870);
or U1394 (N_1394,In_1605,In_752);
nor U1395 (N_1395,In_147,In_123);
xnor U1396 (N_1396,In_358,In_1422);
nor U1397 (N_1397,In_1486,In_1838);
and U1398 (N_1398,In_2362,In_2094);
nand U1399 (N_1399,In_1015,In_1329);
nand U1400 (N_1400,In_1964,In_2187);
nor U1401 (N_1401,In_1600,In_852);
xor U1402 (N_1402,In_2104,In_1398);
and U1403 (N_1403,In_1441,In_1167);
nor U1404 (N_1404,In_2022,In_2428);
xor U1405 (N_1405,In_2058,In_526);
and U1406 (N_1406,In_1888,In_1233);
nand U1407 (N_1407,In_2135,In_902);
nand U1408 (N_1408,In_1239,In_1129);
or U1409 (N_1409,In_1724,In_2488);
or U1410 (N_1410,In_88,In_184);
and U1411 (N_1411,In_483,In_1612);
and U1412 (N_1412,In_2176,In_2234);
or U1413 (N_1413,In_1261,In_1265);
xnor U1414 (N_1414,In_1851,In_456);
xor U1415 (N_1415,In_1607,In_2469);
xor U1416 (N_1416,In_1561,In_2404);
xnor U1417 (N_1417,In_1951,In_311);
or U1418 (N_1418,In_320,In_1592);
nand U1419 (N_1419,In_235,In_778);
nand U1420 (N_1420,In_467,In_1204);
nand U1421 (N_1421,In_716,In_652);
nand U1422 (N_1422,In_1155,In_876);
nor U1423 (N_1423,In_2043,In_663);
or U1424 (N_1424,In_1035,In_1827);
or U1425 (N_1425,In_511,In_1349);
and U1426 (N_1426,In_2129,In_1329);
nor U1427 (N_1427,In_481,In_2138);
xnor U1428 (N_1428,In_1389,In_2041);
nand U1429 (N_1429,In_981,In_410);
or U1430 (N_1430,In_1741,In_1214);
nand U1431 (N_1431,In_1985,In_970);
nand U1432 (N_1432,In_51,In_1183);
or U1433 (N_1433,In_230,In_2265);
and U1434 (N_1434,In_1785,In_2326);
nor U1435 (N_1435,In_1451,In_1946);
xor U1436 (N_1436,In_2470,In_2386);
xnor U1437 (N_1437,In_1155,In_211);
and U1438 (N_1438,In_2468,In_2169);
nor U1439 (N_1439,In_288,In_1019);
nor U1440 (N_1440,In_1210,In_885);
nor U1441 (N_1441,In_1017,In_1038);
nor U1442 (N_1442,In_83,In_1377);
xnor U1443 (N_1443,In_1836,In_655);
nor U1444 (N_1444,In_958,In_1122);
or U1445 (N_1445,In_619,In_396);
or U1446 (N_1446,In_2446,In_444);
and U1447 (N_1447,In_1145,In_22);
and U1448 (N_1448,In_620,In_2208);
nor U1449 (N_1449,In_1720,In_422);
nor U1450 (N_1450,In_2010,In_316);
nand U1451 (N_1451,In_29,In_350);
or U1452 (N_1452,In_711,In_23);
nand U1453 (N_1453,In_1587,In_978);
or U1454 (N_1454,In_529,In_208);
nor U1455 (N_1455,In_1736,In_1364);
nand U1456 (N_1456,In_270,In_23);
nor U1457 (N_1457,In_2186,In_501);
nand U1458 (N_1458,In_856,In_191);
xnor U1459 (N_1459,In_2325,In_993);
and U1460 (N_1460,In_1513,In_1286);
or U1461 (N_1461,In_1719,In_2386);
and U1462 (N_1462,In_939,In_403);
and U1463 (N_1463,In_1266,In_1267);
xnor U1464 (N_1464,In_2169,In_2258);
xor U1465 (N_1465,In_1731,In_1883);
nand U1466 (N_1466,In_1563,In_445);
and U1467 (N_1467,In_1553,In_272);
or U1468 (N_1468,In_2140,In_1171);
nand U1469 (N_1469,In_2099,In_130);
and U1470 (N_1470,In_1977,In_2046);
nor U1471 (N_1471,In_2327,In_877);
and U1472 (N_1472,In_1459,In_2186);
nor U1473 (N_1473,In_387,In_120);
nor U1474 (N_1474,In_1566,In_2319);
nor U1475 (N_1475,In_1608,In_2356);
and U1476 (N_1476,In_701,In_2046);
or U1477 (N_1477,In_1070,In_644);
or U1478 (N_1478,In_1487,In_520);
xor U1479 (N_1479,In_2339,In_981);
and U1480 (N_1480,In_943,In_1054);
xnor U1481 (N_1481,In_2032,In_546);
nand U1482 (N_1482,In_1133,In_1810);
and U1483 (N_1483,In_2431,In_1166);
or U1484 (N_1484,In_916,In_2408);
nand U1485 (N_1485,In_1612,In_1331);
nor U1486 (N_1486,In_1447,In_386);
nor U1487 (N_1487,In_628,In_1803);
or U1488 (N_1488,In_1233,In_582);
or U1489 (N_1489,In_2487,In_1344);
and U1490 (N_1490,In_1035,In_504);
xnor U1491 (N_1491,In_994,In_636);
and U1492 (N_1492,In_1785,In_1969);
nor U1493 (N_1493,In_712,In_619);
nor U1494 (N_1494,In_130,In_1513);
or U1495 (N_1495,In_913,In_564);
nand U1496 (N_1496,In_1408,In_1350);
xor U1497 (N_1497,In_635,In_212);
nand U1498 (N_1498,In_1547,In_291);
and U1499 (N_1499,In_1806,In_299);
nor U1500 (N_1500,In_1002,In_2461);
nand U1501 (N_1501,In_2236,In_1375);
and U1502 (N_1502,In_354,In_1598);
and U1503 (N_1503,In_374,In_1293);
xnor U1504 (N_1504,In_2122,In_844);
xor U1505 (N_1505,In_655,In_1700);
nor U1506 (N_1506,In_160,In_1367);
nor U1507 (N_1507,In_1495,In_871);
xnor U1508 (N_1508,In_181,In_2223);
and U1509 (N_1509,In_1453,In_2417);
nand U1510 (N_1510,In_2162,In_2136);
nor U1511 (N_1511,In_1086,In_644);
nor U1512 (N_1512,In_1773,In_693);
or U1513 (N_1513,In_1904,In_1824);
xnor U1514 (N_1514,In_1832,In_152);
and U1515 (N_1515,In_1657,In_2164);
nand U1516 (N_1516,In_659,In_1403);
nand U1517 (N_1517,In_2309,In_36);
nand U1518 (N_1518,In_1563,In_2053);
nand U1519 (N_1519,In_1210,In_1595);
and U1520 (N_1520,In_595,In_251);
nand U1521 (N_1521,In_328,In_1315);
xnor U1522 (N_1522,In_825,In_416);
nor U1523 (N_1523,In_1830,In_2136);
nand U1524 (N_1524,In_1743,In_514);
and U1525 (N_1525,In_1639,In_2243);
xnor U1526 (N_1526,In_1688,In_1652);
nand U1527 (N_1527,In_439,In_57);
nand U1528 (N_1528,In_1258,In_1921);
nor U1529 (N_1529,In_2294,In_2101);
xor U1530 (N_1530,In_210,In_239);
xor U1531 (N_1531,In_1565,In_179);
nor U1532 (N_1532,In_55,In_1741);
and U1533 (N_1533,In_911,In_900);
and U1534 (N_1534,In_2209,In_61);
and U1535 (N_1535,In_2092,In_1610);
or U1536 (N_1536,In_674,In_2096);
xor U1537 (N_1537,In_2232,In_1943);
nand U1538 (N_1538,In_182,In_2274);
xnor U1539 (N_1539,In_1326,In_1842);
or U1540 (N_1540,In_1778,In_2150);
nand U1541 (N_1541,In_1608,In_81);
and U1542 (N_1542,In_2387,In_1020);
and U1543 (N_1543,In_376,In_1915);
xnor U1544 (N_1544,In_735,In_1557);
or U1545 (N_1545,In_90,In_1318);
or U1546 (N_1546,In_969,In_427);
xnor U1547 (N_1547,In_1577,In_485);
nand U1548 (N_1548,In_1321,In_827);
nor U1549 (N_1549,In_955,In_2185);
nor U1550 (N_1550,In_315,In_1749);
nor U1551 (N_1551,In_2016,In_1914);
xor U1552 (N_1552,In_1160,In_213);
nand U1553 (N_1553,In_1765,In_2249);
xnor U1554 (N_1554,In_1890,In_2422);
nor U1555 (N_1555,In_2184,In_2294);
or U1556 (N_1556,In_1607,In_1458);
or U1557 (N_1557,In_58,In_388);
nand U1558 (N_1558,In_1622,In_2412);
nand U1559 (N_1559,In_1790,In_2064);
nand U1560 (N_1560,In_2102,In_329);
and U1561 (N_1561,In_2395,In_1077);
or U1562 (N_1562,In_531,In_491);
nand U1563 (N_1563,In_783,In_1811);
and U1564 (N_1564,In_399,In_301);
and U1565 (N_1565,In_2440,In_2419);
nand U1566 (N_1566,In_2364,In_803);
nor U1567 (N_1567,In_651,In_1406);
nor U1568 (N_1568,In_761,In_1176);
nor U1569 (N_1569,In_2130,In_116);
nor U1570 (N_1570,In_1144,In_1142);
xor U1571 (N_1571,In_2136,In_189);
and U1572 (N_1572,In_2115,In_690);
xnor U1573 (N_1573,In_1553,In_1746);
xnor U1574 (N_1574,In_925,In_1936);
xor U1575 (N_1575,In_849,In_1740);
nand U1576 (N_1576,In_709,In_1555);
or U1577 (N_1577,In_2274,In_955);
xor U1578 (N_1578,In_575,In_909);
nor U1579 (N_1579,In_266,In_2114);
and U1580 (N_1580,In_881,In_1534);
or U1581 (N_1581,In_341,In_2173);
xnor U1582 (N_1582,In_51,In_897);
xor U1583 (N_1583,In_2492,In_1204);
xor U1584 (N_1584,In_1833,In_1759);
or U1585 (N_1585,In_1293,In_1715);
nand U1586 (N_1586,In_541,In_2355);
xor U1587 (N_1587,In_60,In_1491);
nand U1588 (N_1588,In_1888,In_353);
and U1589 (N_1589,In_1923,In_237);
or U1590 (N_1590,In_921,In_1668);
nor U1591 (N_1591,In_2117,In_1850);
or U1592 (N_1592,In_2020,In_128);
xnor U1593 (N_1593,In_2382,In_842);
xor U1594 (N_1594,In_1444,In_1013);
and U1595 (N_1595,In_1757,In_1084);
or U1596 (N_1596,In_1639,In_1374);
and U1597 (N_1597,In_1093,In_1117);
nand U1598 (N_1598,In_2495,In_471);
nor U1599 (N_1599,In_862,In_1700);
xnor U1600 (N_1600,In_757,In_1968);
nand U1601 (N_1601,In_2224,In_1492);
and U1602 (N_1602,In_1256,In_328);
or U1603 (N_1603,In_1586,In_1985);
or U1604 (N_1604,In_1133,In_2456);
or U1605 (N_1605,In_308,In_870);
nand U1606 (N_1606,In_555,In_1719);
xnor U1607 (N_1607,In_1060,In_1616);
xor U1608 (N_1608,In_331,In_380);
or U1609 (N_1609,In_817,In_1147);
nand U1610 (N_1610,In_1778,In_1446);
or U1611 (N_1611,In_2357,In_1632);
nor U1612 (N_1612,In_2106,In_1835);
nor U1613 (N_1613,In_2088,In_1409);
nor U1614 (N_1614,In_34,In_890);
xor U1615 (N_1615,In_597,In_361);
and U1616 (N_1616,In_1846,In_1900);
xor U1617 (N_1617,In_2008,In_35);
and U1618 (N_1618,In_1860,In_845);
xnor U1619 (N_1619,In_451,In_428);
xnor U1620 (N_1620,In_1998,In_796);
and U1621 (N_1621,In_2317,In_128);
nor U1622 (N_1622,In_1919,In_1721);
and U1623 (N_1623,In_1419,In_1520);
xnor U1624 (N_1624,In_2197,In_734);
and U1625 (N_1625,In_1242,In_2221);
or U1626 (N_1626,In_1463,In_2077);
or U1627 (N_1627,In_1608,In_114);
and U1628 (N_1628,In_2265,In_288);
xnor U1629 (N_1629,In_1348,In_1318);
nor U1630 (N_1630,In_2150,In_2465);
and U1631 (N_1631,In_1853,In_187);
nand U1632 (N_1632,In_2081,In_1667);
and U1633 (N_1633,In_1669,In_1007);
nor U1634 (N_1634,In_1629,In_1473);
nor U1635 (N_1635,In_554,In_192);
xor U1636 (N_1636,In_45,In_1067);
and U1637 (N_1637,In_371,In_1446);
and U1638 (N_1638,In_2422,In_1950);
nor U1639 (N_1639,In_29,In_867);
nor U1640 (N_1640,In_1886,In_1242);
nor U1641 (N_1641,In_1840,In_562);
nand U1642 (N_1642,In_1514,In_877);
nand U1643 (N_1643,In_867,In_1286);
nand U1644 (N_1644,In_1200,In_2150);
nor U1645 (N_1645,In_2475,In_188);
and U1646 (N_1646,In_1295,In_2216);
and U1647 (N_1647,In_1574,In_936);
nand U1648 (N_1648,In_2035,In_1752);
nor U1649 (N_1649,In_1110,In_1864);
and U1650 (N_1650,In_755,In_1634);
or U1651 (N_1651,In_678,In_2303);
nor U1652 (N_1652,In_672,In_1785);
nand U1653 (N_1653,In_1615,In_1342);
nor U1654 (N_1654,In_417,In_1916);
xnor U1655 (N_1655,In_1161,In_1147);
nor U1656 (N_1656,In_1521,In_1737);
xnor U1657 (N_1657,In_750,In_530);
nand U1658 (N_1658,In_2464,In_176);
and U1659 (N_1659,In_514,In_1385);
nor U1660 (N_1660,In_633,In_2008);
and U1661 (N_1661,In_1030,In_2005);
xor U1662 (N_1662,In_575,In_1522);
nand U1663 (N_1663,In_1906,In_1855);
xnor U1664 (N_1664,In_76,In_793);
nand U1665 (N_1665,In_988,In_1599);
nand U1666 (N_1666,In_752,In_110);
and U1667 (N_1667,In_665,In_1749);
and U1668 (N_1668,In_2224,In_1947);
and U1669 (N_1669,In_1106,In_982);
and U1670 (N_1670,In_1077,In_2190);
nand U1671 (N_1671,In_1402,In_2468);
xor U1672 (N_1672,In_1127,In_1130);
or U1673 (N_1673,In_917,In_2430);
nand U1674 (N_1674,In_454,In_481);
or U1675 (N_1675,In_934,In_1689);
nand U1676 (N_1676,In_1644,In_202);
nand U1677 (N_1677,In_247,In_2311);
xor U1678 (N_1678,In_881,In_1198);
xor U1679 (N_1679,In_552,In_841);
xnor U1680 (N_1680,In_1800,In_2052);
xor U1681 (N_1681,In_1807,In_828);
nor U1682 (N_1682,In_754,In_1504);
nor U1683 (N_1683,In_983,In_312);
nor U1684 (N_1684,In_367,In_490);
and U1685 (N_1685,In_1213,In_2198);
or U1686 (N_1686,In_1599,In_787);
xnor U1687 (N_1687,In_1479,In_2464);
nor U1688 (N_1688,In_158,In_2448);
nand U1689 (N_1689,In_158,In_2378);
or U1690 (N_1690,In_1219,In_157);
xnor U1691 (N_1691,In_433,In_151);
xnor U1692 (N_1692,In_682,In_1753);
xor U1693 (N_1693,In_1461,In_233);
or U1694 (N_1694,In_1828,In_201);
xnor U1695 (N_1695,In_165,In_2365);
nand U1696 (N_1696,In_513,In_842);
nor U1697 (N_1697,In_798,In_595);
and U1698 (N_1698,In_1798,In_1071);
nor U1699 (N_1699,In_369,In_1875);
nor U1700 (N_1700,In_314,In_2346);
or U1701 (N_1701,In_1302,In_2183);
or U1702 (N_1702,In_1060,In_906);
or U1703 (N_1703,In_2052,In_2001);
or U1704 (N_1704,In_1890,In_721);
or U1705 (N_1705,In_1837,In_460);
nor U1706 (N_1706,In_1158,In_262);
or U1707 (N_1707,In_1228,In_1143);
xor U1708 (N_1708,In_1480,In_1345);
nor U1709 (N_1709,In_487,In_610);
xor U1710 (N_1710,In_1979,In_2388);
nand U1711 (N_1711,In_1524,In_826);
or U1712 (N_1712,In_32,In_2467);
or U1713 (N_1713,In_2135,In_1359);
xnor U1714 (N_1714,In_725,In_529);
or U1715 (N_1715,In_2434,In_1215);
nor U1716 (N_1716,In_339,In_1844);
nor U1717 (N_1717,In_1822,In_115);
nor U1718 (N_1718,In_1261,In_232);
nor U1719 (N_1719,In_1619,In_1032);
nand U1720 (N_1720,In_34,In_145);
nand U1721 (N_1721,In_797,In_119);
nand U1722 (N_1722,In_268,In_1260);
or U1723 (N_1723,In_1143,In_1657);
or U1724 (N_1724,In_1880,In_863);
nor U1725 (N_1725,In_505,In_2179);
or U1726 (N_1726,In_1956,In_1887);
xor U1727 (N_1727,In_1878,In_2012);
or U1728 (N_1728,In_410,In_242);
nor U1729 (N_1729,In_44,In_846);
and U1730 (N_1730,In_185,In_369);
nor U1731 (N_1731,In_1052,In_310);
or U1732 (N_1732,In_1485,In_1413);
nand U1733 (N_1733,In_961,In_2254);
nor U1734 (N_1734,In_1816,In_2095);
xor U1735 (N_1735,In_470,In_2165);
xor U1736 (N_1736,In_1380,In_13);
nor U1737 (N_1737,In_1723,In_2443);
nor U1738 (N_1738,In_1316,In_91);
nand U1739 (N_1739,In_2431,In_234);
or U1740 (N_1740,In_1410,In_1439);
or U1741 (N_1741,In_816,In_858);
nand U1742 (N_1742,In_1734,In_24);
nor U1743 (N_1743,In_73,In_618);
nor U1744 (N_1744,In_328,In_1518);
and U1745 (N_1745,In_1675,In_190);
xor U1746 (N_1746,In_1183,In_499);
nand U1747 (N_1747,In_384,In_1292);
nand U1748 (N_1748,In_2011,In_2168);
and U1749 (N_1749,In_88,In_468);
nand U1750 (N_1750,In_686,In_1094);
or U1751 (N_1751,In_1661,In_2089);
or U1752 (N_1752,In_1435,In_93);
or U1753 (N_1753,In_490,In_2141);
nor U1754 (N_1754,In_1614,In_793);
and U1755 (N_1755,In_2042,In_1633);
xnor U1756 (N_1756,In_1346,In_107);
nand U1757 (N_1757,In_707,In_1604);
and U1758 (N_1758,In_634,In_80);
nor U1759 (N_1759,In_1715,In_765);
and U1760 (N_1760,In_480,In_1752);
nor U1761 (N_1761,In_877,In_989);
and U1762 (N_1762,In_470,In_151);
xor U1763 (N_1763,In_1493,In_1801);
xnor U1764 (N_1764,In_278,In_825);
nand U1765 (N_1765,In_2085,In_1091);
xor U1766 (N_1766,In_1649,In_322);
nor U1767 (N_1767,In_474,In_2059);
and U1768 (N_1768,In_80,In_2412);
nand U1769 (N_1769,In_2415,In_2228);
nand U1770 (N_1770,In_2421,In_2245);
nor U1771 (N_1771,In_1426,In_1781);
or U1772 (N_1772,In_253,In_1457);
xor U1773 (N_1773,In_1649,In_625);
nand U1774 (N_1774,In_296,In_495);
nor U1775 (N_1775,In_614,In_1277);
xor U1776 (N_1776,In_55,In_1584);
or U1777 (N_1777,In_1375,In_163);
nand U1778 (N_1778,In_1721,In_332);
or U1779 (N_1779,In_471,In_323);
nor U1780 (N_1780,In_1729,In_1578);
xnor U1781 (N_1781,In_2417,In_83);
nor U1782 (N_1782,In_2237,In_2413);
nand U1783 (N_1783,In_904,In_2289);
xnor U1784 (N_1784,In_621,In_643);
xor U1785 (N_1785,In_53,In_1637);
nor U1786 (N_1786,In_1183,In_848);
xnor U1787 (N_1787,In_1010,In_2110);
or U1788 (N_1788,In_2010,In_1863);
or U1789 (N_1789,In_2095,In_401);
and U1790 (N_1790,In_11,In_1676);
or U1791 (N_1791,In_1508,In_989);
nor U1792 (N_1792,In_1538,In_2106);
nand U1793 (N_1793,In_227,In_2233);
xnor U1794 (N_1794,In_2278,In_222);
or U1795 (N_1795,In_49,In_539);
or U1796 (N_1796,In_1205,In_794);
nor U1797 (N_1797,In_1818,In_2018);
and U1798 (N_1798,In_495,In_1198);
nand U1799 (N_1799,In_1728,In_813);
or U1800 (N_1800,In_146,In_1304);
nand U1801 (N_1801,In_520,In_1985);
and U1802 (N_1802,In_630,In_30);
or U1803 (N_1803,In_515,In_1730);
nor U1804 (N_1804,In_890,In_1645);
nand U1805 (N_1805,In_3,In_1768);
or U1806 (N_1806,In_1977,In_1060);
nor U1807 (N_1807,In_180,In_2464);
and U1808 (N_1808,In_433,In_1773);
and U1809 (N_1809,In_1845,In_1649);
or U1810 (N_1810,In_1406,In_1845);
xnor U1811 (N_1811,In_894,In_737);
xnor U1812 (N_1812,In_126,In_456);
nor U1813 (N_1813,In_95,In_2456);
nand U1814 (N_1814,In_1747,In_696);
and U1815 (N_1815,In_1644,In_1417);
or U1816 (N_1816,In_530,In_1607);
or U1817 (N_1817,In_1351,In_1708);
nand U1818 (N_1818,In_853,In_614);
and U1819 (N_1819,In_1497,In_819);
or U1820 (N_1820,In_2469,In_2107);
and U1821 (N_1821,In_1408,In_1265);
or U1822 (N_1822,In_218,In_1791);
nand U1823 (N_1823,In_909,In_2077);
nand U1824 (N_1824,In_14,In_1006);
nand U1825 (N_1825,In_1046,In_2293);
nand U1826 (N_1826,In_2411,In_1162);
nor U1827 (N_1827,In_561,In_2208);
or U1828 (N_1828,In_902,In_2329);
xnor U1829 (N_1829,In_209,In_2017);
nor U1830 (N_1830,In_258,In_1931);
nor U1831 (N_1831,In_2343,In_1491);
and U1832 (N_1832,In_1823,In_1301);
nor U1833 (N_1833,In_271,In_1821);
nand U1834 (N_1834,In_1855,In_523);
or U1835 (N_1835,In_688,In_388);
nor U1836 (N_1836,In_1329,In_1860);
nand U1837 (N_1837,In_2318,In_1492);
nand U1838 (N_1838,In_883,In_238);
xor U1839 (N_1839,In_921,In_2261);
nand U1840 (N_1840,In_365,In_1998);
nor U1841 (N_1841,In_521,In_25);
nand U1842 (N_1842,In_1543,In_629);
xor U1843 (N_1843,In_505,In_2225);
xor U1844 (N_1844,In_1758,In_783);
xnor U1845 (N_1845,In_2286,In_2005);
or U1846 (N_1846,In_867,In_970);
or U1847 (N_1847,In_1904,In_2392);
and U1848 (N_1848,In_151,In_1527);
nand U1849 (N_1849,In_1047,In_1924);
xor U1850 (N_1850,In_139,In_1735);
and U1851 (N_1851,In_1631,In_1449);
nor U1852 (N_1852,In_1356,In_197);
nand U1853 (N_1853,In_1924,In_72);
and U1854 (N_1854,In_2161,In_493);
or U1855 (N_1855,In_227,In_265);
xnor U1856 (N_1856,In_556,In_1537);
nand U1857 (N_1857,In_1441,In_900);
xnor U1858 (N_1858,In_88,In_1142);
xor U1859 (N_1859,In_1278,In_1099);
and U1860 (N_1860,In_2379,In_2353);
nand U1861 (N_1861,In_2013,In_1529);
and U1862 (N_1862,In_30,In_888);
nand U1863 (N_1863,In_2181,In_1824);
or U1864 (N_1864,In_1183,In_562);
xnor U1865 (N_1865,In_952,In_1672);
nor U1866 (N_1866,In_2039,In_2029);
or U1867 (N_1867,In_420,In_1581);
xnor U1868 (N_1868,In_1636,In_1277);
or U1869 (N_1869,In_1680,In_1717);
nand U1870 (N_1870,In_737,In_804);
nor U1871 (N_1871,In_510,In_1430);
nand U1872 (N_1872,In_1718,In_2370);
and U1873 (N_1873,In_1826,In_960);
and U1874 (N_1874,In_2074,In_1725);
xnor U1875 (N_1875,In_819,In_1361);
nor U1876 (N_1876,In_1523,In_558);
or U1877 (N_1877,In_920,In_1978);
xnor U1878 (N_1878,In_2431,In_2384);
or U1879 (N_1879,In_197,In_49);
and U1880 (N_1880,In_1641,In_1072);
xor U1881 (N_1881,In_798,In_1469);
or U1882 (N_1882,In_1052,In_422);
or U1883 (N_1883,In_2408,In_340);
or U1884 (N_1884,In_1624,In_1154);
or U1885 (N_1885,In_391,In_750);
and U1886 (N_1886,In_2037,In_902);
nor U1887 (N_1887,In_1981,In_399);
or U1888 (N_1888,In_1528,In_1234);
or U1889 (N_1889,In_2270,In_2163);
nand U1890 (N_1890,In_1252,In_1798);
xor U1891 (N_1891,In_1710,In_750);
or U1892 (N_1892,In_888,In_1063);
or U1893 (N_1893,In_2491,In_2227);
and U1894 (N_1894,In_53,In_409);
and U1895 (N_1895,In_2197,In_2084);
xnor U1896 (N_1896,In_1801,In_2251);
and U1897 (N_1897,In_68,In_687);
and U1898 (N_1898,In_2429,In_2396);
nand U1899 (N_1899,In_228,In_1625);
and U1900 (N_1900,In_2432,In_84);
xnor U1901 (N_1901,In_310,In_2265);
xnor U1902 (N_1902,In_1703,In_1716);
nand U1903 (N_1903,In_2261,In_232);
or U1904 (N_1904,In_966,In_987);
xnor U1905 (N_1905,In_163,In_626);
or U1906 (N_1906,In_1686,In_83);
nand U1907 (N_1907,In_1536,In_2198);
nor U1908 (N_1908,In_2367,In_737);
or U1909 (N_1909,In_1422,In_1918);
or U1910 (N_1910,In_1488,In_872);
xnor U1911 (N_1911,In_2329,In_786);
nor U1912 (N_1912,In_1372,In_1079);
xnor U1913 (N_1913,In_1756,In_1887);
or U1914 (N_1914,In_1793,In_1322);
and U1915 (N_1915,In_56,In_2288);
or U1916 (N_1916,In_394,In_160);
and U1917 (N_1917,In_798,In_2248);
nor U1918 (N_1918,In_230,In_1318);
or U1919 (N_1919,In_618,In_1627);
or U1920 (N_1920,In_2152,In_1971);
and U1921 (N_1921,In_1107,In_998);
nand U1922 (N_1922,In_1709,In_1333);
xnor U1923 (N_1923,In_1416,In_2004);
nand U1924 (N_1924,In_1130,In_655);
and U1925 (N_1925,In_1143,In_1710);
xnor U1926 (N_1926,In_2067,In_1786);
nor U1927 (N_1927,In_1050,In_661);
or U1928 (N_1928,In_113,In_1968);
and U1929 (N_1929,In_2112,In_557);
and U1930 (N_1930,In_297,In_1077);
nor U1931 (N_1931,In_2169,In_2086);
xor U1932 (N_1932,In_1997,In_1811);
nand U1933 (N_1933,In_416,In_1582);
xnor U1934 (N_1934,In_1294,In_216);
xor U1935 (N_1935,In_1796,In_1879);
xnor U1936 (N_1936,In_60,In_1280);
nand U1937 (N_1937,In_1149,In_862);
nand U1938 (N_1938,In_1557,In_27);
xor U1939 (N_1939,In_2144,In_2214);
xnor U1940 (N_1940,In_2326,In_1802);
and U1941 (N_1941,In_44,In_812);
or U1942 (N_1942,In_1767,In_958);
nand U1943 (N_1943,In_2368,In_46);
xnor U1944 (N_1944,In_529,In_1918);
nor U1945 (N_1945,In_380,In_595);
and U1946 (N_1946,In_2432,In_1870);
xnor U1947 (N_1947,In_2268,In_1136);
nor U1948 (N_1948,In_1265,In_1165);
nand U1949 (N_1949,In_1193,In_920);
and U1950 (N_1950,In_1417,In_287);
xor U1951 (N_1951,In_672,In_2304);
nor U1952 (N_1952,In_2319,In_1322);
or U1953 (N_1953,In_59,In_161);
or U1954 (N_1954,In_312,In_2349);
or U1955 (N_1955,In_32,In_2179);
nand U1956 (N_1956,In_1211,In_790);
nor U1957 (N_1957,In_1145,In_446);
and U1958 (N_1958,In_986,In_1205);
nor U1959 (N_1959,In_970,In_2349);
nor U1960 (N_1960,In_1347,In_1024);
nand U1961 (N_1961,In_1984,In_701);
or U1962 (N_1962,In_1503,In_2068);
and U1963 (N_1963,In_414,In_70);
or U1964 (N_1964,In_2156,In_643);
and U1965 (N_1965,In_2492,In_1402);
xnor U1966 (N_1966,In_995,In_763);
xor U1967 (N_1967,In_685,In_1526);
and U1968 (N_1968,In_1308,In_461);
xnor U1969 (N_1969,In_2378,In_500);
nor U1970 (N_1970,In_2378,In_757);
and U1971 (N_1971,In_213,In_1614);
xnor U1972 (N_1972,In_1867,In_754);
or U1973 (N_1973,In_1778,In_1260);
nand U1974 (N_1974,In_872,In_1934);
nor U1975 (N_1975,In_765,In_724);
xor U1976 (N_1976,In_1139,In_1714);
nor U1977 (N_1977,In_1974,In_1045);
xnor U1978 (N_1978,In_1560,In_885);
and U1979 (N_1979,In_409,In_949);
nor U1980 (N_1980,In_1289,In_2293);
xnor U1981 (N_1981,In_669,In_2215);
nor U1982 (N_1982,In_2216,In_1384);
nor U1983 (N_1983,In_2135,In_162);
xor U1984 (N_1984,In_177,In_1356);
and U1985 (N_1985,In_1079,In_807);
nand U1986 (N_1986,In_700,In_2203);
or U1987 (N_1987,In_1301,In_1650);
nand U1988 (N_1988,In_559,In_755);
or U1989 (N_1989,In_43,In_347);
and U1990 (N_1990,In_1460,In_1260);
nand U1991 (N_1991,In_901,In_2421);
nand U1992 (N_1992,In_78,In_1348);
nand U1993 (N_1993,In_1099,In_1874);
nor U1994 (N_1994,In_801,In_1357);
nor U1995 (N_1995,In_2172,In_1178);
nor U1996 (N_1996,In_1643,In_177);
nor U1997 (N_1997,In_793,In_530);
nor U1998 (N_1998,In_842,In_1509);
nor U1999 (N_1999,In_49,In_710);
xor U2000 (N_2000,In_1185,In_2223);
nor U2001 (N_2001,In_1923,In_1463);
nor U2002 (N_2002,In_2195,In_1594);
or U2003 (N_2003,In_2394,In_2260);
or U2004 (N_2004,In_478,In_2037);
nand U2005 (N_2005,In_330,In_1315);
nand U2006 (N_2006,In_1487,In_1611);
and U2007 (N_2007,In_1191,In_789);
nor U2008 (N_2008,In_1272,In_505);
or U2009 (N_2009,In_1841,In_2355);
nor U2010 (N_2010,In_618,In_1850);
xor U2011 (N_2011,In_1063,In_2201);
xor U2012 (N_2012,In_1765,In_1269);
and U2013 (N_2013,In_1716,In_1106);
xnor U2014 (N_2014,In_1362,In_405);
xnor U2015 (N_2015,In_616,In_1188);
nand U2016 (N_2016,In_1433,In_2340);
nor U2017 (N_2017,In_2291,In_74);
nand U2018 (N_2018,In_2369,In_330);
and U2019 (N_2019,In_504,In_2298);
xnor U2020 (N_2020,In_2101,In_455);
or U2021 (N_2021,In_2133,In_230);
or U2022 (N_2022,In_355,In_161);
or U2023 (N_2023,In_1459,In_1583);
or U2024 (N_2024,In_1928,In_1599);
xnor U2025 (N_2025,In_1557,In_494);
nor U2026 (N_2026,In_1222,In_2046);
nor U2027 (N_2027,In_1314,In_944);
and U2028 (N_2028,In_1652,In_2479);
and U2029 (N_2029,In_2300,In_2124);
nand U2030 (N_2030,In_2007,In_423);
or U2031 (N_2031,In_1511,In_1522);
nor U2032 (N_2032,In_137,In_354);
nand U2033 (N_2033,In_1029,In_992);
nand U2034 (N_2034,In_432,In_936);
nand U2035 (N_2035,In_128,In_1904);
nand U2036 (N_2036,In_1487,In_1962);
nand U2037 (N_2037,In_2331,In_2326);
nor U2038 (N_2038,In_1082,In_85);
or U2039 (N_2039,In_589,In_66);
nand U2040 (N_2040,In_949,In_1939);
or U2041 (N_2041,In_613,In_1921);
nor U2042 (N_2042,In_326,In_2291);
nor U2043 (N_2043,In_2015,In_32);
xor U2044 (N_2044,In_1406,In_1182);
or U2045 (N_2045,In_1704,In_1537);
nand U2046 (N_2046,In_1825,In_1860);
nor U2047 (N_2047,In_630,In_1352);
nand U2048 (N_2048,In_392,In_508);
or U2049 (N_2049,In_1225,In_1109);
nor U2050 (N_2050,In_205,In_1461);
xor U2051 (N_2051,In_1412,In_95);
xor U2052 (N_2052,In_1441,In_2386);
nand U2053 (N_2053,In_1608,In_2485);
xor U2054 (N_2054,In_498,In_2119);
xnor U2055 (N_2055,In_1032,In_1753);
xnor U2056 (N_2056,In_2314,In_2046);
nor U2057 (N_2057,In_1327,In_380);
or U2058 (N_2058,In_1298,In_1292);
and U2059 (N_2059,In_444,In_822);
xor U2060 (N_2060,In_2087,In_529);
and U2061 (N_2061,In_2116,In_771);
and U2062 (N_2062,In_1393,In_1479);
or U2063 (N_2063,In_598,In_2399);
or U2064 (N_2064,In_2281,In_1635);
or U2065 (N_2065,In_857,In_2308);
xnor U2066 (N_2066,In_1148,In_87);
xnor U2067 (N_2067,In_2365,In_784);
or U2068 (N_2068,In_1503,In_1449);
nand U2069 (N_2069,In_1,In_1121);
xor U2070 (N_2070,In_1495,In_1735);
and U2071 (N_2071,In_722,In_943);
and U2072 (N_2072,In_2182,In_2038);
xnor U2073 (N_2073,In_1170,In_2473);
or U2074 (N_2074,In_289,In_1902);
or U2075 (N_2075,In_1687,In_773);
xor U2076 (N_2076,In_1353,In_885);
and U2077 (N_2077,In_447,In_45);
or U2078 (N_2078,In_2064,In_2028);
xnor U2079 (N_2079,In_85,In_9);
or U2080 (N_2080,In_1507,In_2383);
or U2081 (N_2081,In_531,In_714);
nand U2082 (N_2082,In_1964,In_1645);
and U2083 (N_2083,In_2234,In_2449);
and U2084 (N_2084,In_1894,In_2347);
xnor U2085 (N_2085,In_1299,In_365);
xnor U2086 (N_2086,In_1540,In_1496);
or U2087 (N_2087,In_1973,In_1879);
nor U2088 (N_2088,In_1520,In_1448);
and U2089 (N_2089,In_298,In_8);
xor U2090 (N_2090,In_1216,In_2231);
nand U2091 (N_2091,In_1313,In_2388);
xnor U2092 (N_2092,In_1064,In_465);
xor U2093 (N_2093,In_2109,In_676);
and U2094 (N_2094,In_335,In_1339);
and U2095 (N_2095,In_1149,In_992);
xor U2096 (N_2096,In_2362,In_415);
and U2097 (N_2097,In_998,In_2273);
nor U2098 (N_2098,In_921,In_851);
nor U2099 (N_2099,In_2290,In_573);
or U2100 (N_2100,In_240,In_2139);
nor U2101 (N_2101,In_353,In_188);
nor U2102 (N_2102,In_54,In_2004);
xor U2103 (N_2103,In_2075,In_1981);
nor U2104 (N_2104,In_1259,In_291);
nor U2105 (N_2105,In_687,In_70);
and U2106 (N_2106,In_326,In_864);
or U2107 (N_2107,In_314,In_1104);
nor U2108 (N_2108,In_1216,In_2040);
and U2109 (N_2109,In_1162,In_118);
or U2110 (N_2110,In_1244,In_1120);
nor U2111 (N_2111,In_1040,In_347);
xnor U2112 (N_2112,In_464,In_862);
and U2113 (N_2113,In_1012,In_1815);
and U2114 (N_2114,In_1285,In_1866);
or U2115 (N_2115,In_1406,In_1197);
or U2116 (N_2116,In_789,In_2180);
and U2117 (N_2117,In_514,In_50);
nand U2118 (N_2118,In_1653,In_1992);
or U2119 (N_2119,In_798,In_1081);
or U2120 (N_2120,In_1864,In_1049);
nand U2121 (N_2121,In_820,In_2068);
and U2122 (N_2122,In_1116,In_670);
and U2123 (N_2123,In_1932,In_1385);
or U2124 (N_2124,In_1655,In_2389);
and U2125 (N_2125,In_385,In_543);
xor U2126 (N_2126,In_1833,In_278);
nor U2127 (N_2127,In_1638,In_549);
xnor U2128 (N_2128,In_574,In_1283);
xnor U2129 (N_2129,In_889,In_759);
nor U2130 (N_2130,In_1624,In_77);
and U2131 (N_2131,In_134,In_2041);
xor U2132 (N_2132,In_1210,In_303);
nand U2133 (N_2133,In_65,In_1405);
or U2134 (N_2134,In_1144,In_1143);
nand U2135 (N_2135,In_17,In_1095);
xnor U2136 (N_2136,In_2497,In_2153);
and U2137 (N_2137,In_1936,In_1016);
and U2138 (N_2138,In_213,In_2389);
and U2139 (N_2139,In_1833,In_2413);
xor U2140 (N_2140,In_1607,In_1610);
xor U2141 (N_2141,In_2131,In_2109);
xor U2142 (N_2142,In_1411,In_380);
nand U2143 (N_2143,In_2210,In_1118);
xnor U2144 (N_2144,In_1874,In_2016);
or U2145 (N_2145,In_1336,In_275);
nand U2146 (N_2146,In_1795,In_1889);
or U2147 (N_2147,In_1790,In_1808);
nor U2148 (N_2148,In_970,In_2139);
nor U2149 (N_2149,In_2468,In_1378);
nor U2150 (N_2150,In_1963,In_1661);
or U2151 (N_2151,In_1019,In_17);
xor U2152 (N_2152,In_1058,In_1030);
nand U2153 (N_2153,In_177,In_763);
and U2154 (N_2154,In_1350,In_1156);
xnor U2155 (N_2155,In_947,In_2045);
nand U2156 (N_2156,In_1213,In_175);
xnor U2157 (N_2157,In_36,In_1119);
and U2158 (N_2158,In_1033,In_1819);
nor U2159 (N_2159,In_127,In_483);
xor U2160 (N_2160,In_812,In_1392);
and U2161 (N_2161,In_1829,In_84);
and U2162 (N_2162,In_1277,In_833);
xor U2163 (N_2163,In_1559,In_1881);
nor U2164 (N_2164,In_142,In_1831);
nand U2165 (N_2165,In_937,In_719);
and U2166 (N_2166,In_1383,In_2464);
nor U2167 (N_2167,In_2406,In_626);
nand U2168 (N_2168,In_1592,In_1880);
nand U2169 (N_2169,In_2184,In_1418);
xnor U2170 (N_2170,In_310,In_1440);
or U2171 (N_2171,In_1157,In_564);
or U2172 (N_2172,In_252,In_2);
and U2173 (N_2173,In_1347,In_1346);
and U2174 (N_2174,In_2408,In_1271);
nand U2175 (N_2175,In_265,In_1103);
nor U2176 (N_2176,In_47,In_2351);
nor U2177 (N_2177,In_2218,In_2330);
and U2178 (N_2178,In_543,In_328);
nor U2179 (N_2179,In_2163,In_937);
nand U2180 (N_2180,In_1093,In_272);
or U2181 (N_2181,In_507,In_1454);
or U2182 (N_2182,In_1449,In_2354);
or U2183 (N_2183,In_1666,In_1773);
nor U2184 (N_2184,In_1524,In_656);
nor U2185 (N_2185,In_335,In_285);
and U2186 (N_2186,In_802,In_132);
nand U2187 (N_2187,In_11,In_1289);
and U2188 (N_2188,In_1194,In_33);
nand U2189 (N_2189,In_2027,In_983);
nor U2190 (N_2190,In_1643,In_1902);
nor U2191 (N_2191,In_1063,In_2139);
nor U2192 (N_2192,In_2092,In_678);
nor U2193 (N_2193,In_601,In_2492);
and U2194 (N_2194,In_1834,In_1250);
nand U2195 (N_2195,In_2256,In_1365);
or U2196 (N_2196,In_830,In_1456);
and U2197 (N_2197,In_1395,In_2164);
xor U2198 (N_2198,In_85,In_1821);
nor U2199 (N_2199,In_976,In_1384);
xor U2200 (N_2200,In_1045,In_2061);
nor U2201 (N_2201,In_721,In_99);
xnor U2202 (N_2202,In_1312,In_155);
nand U2203 (N_2203,In_1935,In_823);
xor U2204 (N_2204,In_1125,In_898);
nand U2205 (N_2205,In_976,In_127);
and U2206 (N_2206,In_905,In_2383);
xnor U2207 (N_2207,In_1294,In_2132);
or U2208 (N_2208,In_293,In_2314);
nand U2209 (N_2209,In_1444,In_1609);
and U2210 (N_2210,In_0,In_2250);
and U2211 (N_2211,In_2166,In_1565);
nor U2212 (N_2212,In_2263,In_1250);
and U2213 (N_2213,In_634,In_1471);
nand U2214 (N_2214,In_334,In_1112);
nand U2215 (N_2215,In_1122,In_1130);
or U2216 (N_2216,In_1218,In_787);
or U2217 (N_2217,In_143,In_292);
nand U2218 (N_2218,In_821,In_1584);
and U2219 (N_2219,In_1894,In_1151);
xor U2220 (N_2220,In_1998,In_576);
or U2221 (N_2221,In_432,In_2468);
xnor U2222 (N_2222,In_921,In_1482);
or U2223 (N_2223,In_2080,In_2366);
and U2224 (N_2224,In_1017,In_2461);
nand U2225 (N_2225,In_1123,In_1213);
nand U2226 (N_2226,In_2176,In_706);
and U2227 (N_2227,In_14,In_252);
xor U2228 (N_2228,In_2195,In_1489);
nor U2229 (N_2229,In_1639,In_2173);
nand U2230 (N_2230,In_303,In_985);
xor U2231 (N_2231,In_750,In_837);
or U2232 (N_2232,In_383,In_256);
or U2233 (N_2233,In_855,In_2216);
nand U2234 (N_2234,In_1839,In_1213);
nand U2235 (N_2235,In_1254,In_706);
xor U2236 (N_2236,In_356,In_763);
or U2237 (N_2237,In_660,In_2422);
or U2238 (N_2238,In_17,In_194);
nand U2239 (N_2239,In_1330,In_1705);
xor U2240 (N_2240,In_250,In_1412);
and U2241 (N_2241,In_2181,In_1177);
nand U2242 (N_2242,In_2146,In_42);
nor U2243 (N_2243,In_1096,In_707);
nand U2244 (N_2244,In_1772,In_776);
nor U2245 (N_2245,In_206,In_304);
nor U2246 (N_2246,In_804,In_2121);
and U2247 (N_2247,In_1746,In_1783);
nor U2248 (N_2248,In_825,In_1984);
nand U2249 (N_2249,In_407,In_2341);
nand U2250 (N_2250,In_37,In_417);
nor U2251 (N_2251,In_2071,In_1890);
nand U2252 (N_2252,In_1060,In_360);
nor U2253 (N_2253,In_2052,In_930);
and U2254 (N_2254,In_217,In_1623);
or U2255 (N_2255,In_1392,In_1124);
nand U2256 (N_2256,In_2336,In_1109);
or U2257 (N_2257,In_1099,In_1756);
nor U2258 (N_2258,In_642,In_212);
xor U2259 (N_2259,In_1441,In_1613);
nor U2260 (N_2260,In_1427,In_992);
or U2261 (N_2261,In_1715,In_597);
nor U2262 (N_2262,In_75,In_2349);
xor U2263 (N_2263,In_1949,In_566);
or U2264 (N_2264,In_1630,In_1391);
and U2265 (N_2265,In_1621,In_1238);
or U2266 (N_2266,In_1350,In_1946);
nor U2267 (N_2267,In_2163,In_101);
and U2268 (N_2268,In_1065,In_1020);
and U2269 (N_2269,In_813,In_2263);
nand U2270 (N_2270,In_1334,In_679);
or U2271 (N_2271,In_889,In_2160);
and U2272 (N_2272,In_1137,In_2381);
nor U2273 (N_2273,In_2026,In_2191);
xor U2274 (N_2274,In_1724,In_2360);
and U2275 (N_2275,In_1919,In_369);
and U2276 (N_2276,In_1553,In_1341);
and U2277 (N_2277,In_172,In_1748);
nand U2278 (N_2278,In_1514,In_1203);
and U2279 (N_2279,In_373,In_2399);
and U2280 (N_2280,In_1711,In_190);
and U2281 (N_2281,In_834,In_1487);
or U2282 (N_2282,In_808,In_2413);
nor U2283 (N_2283,In_774,In_2390);
nor U2284 (N_2284,In_646,In_639);
nand U2285 (N_2285,In_1889,In_1924);
xnor U2286 (N_2286,In_1540,In_1289);
and U2287 (N_2287,In_2499,In_2152);
nor U2288 (N_2288,In_1537,In_1709);
nand U2289 (N_2289,In_561,In_360);
xnor U2290 (N_2290,In_640,In_249);
and U2291 (N_2291,In_1880,In_65);
or U2292 (N_2292,In_1510,In_910);
and U2293 (N_2293,In_2308,In_1954);
and U2294 (N_2294,In_338,In_1025);
or U2295 (N_2295,In_2153,In_1484);
xor U2296 (N_2296,In_1879,In_1748);
and U2297 (N_2297,In_828,In_2146);
nand U2298 (N_2298,In_2477,In_2103);
or U2299 (N_2299,In_2091,In_1370);
nor U2300 (N_2300,In_877,In_2130);
xnor U2301 (N_2301,In_2173,In_2483);
xor U2302 (N_2302,In_2061,In_243);
nand U2303 (N_2303,In_548,In_1069);
and U2304 (N_2304,In_1931,In_922);
and U2305 (N_2305,In_511,In_1639);
and U2306 (N_2306,In_2497,In_1097);
nand U2307 (N_2307,In_2378,In_399);
xnor U2308 (N_2308,In_2442,In_999);
xor U2309 (N_2309,In_2246,In_1186);
or U2310 (N_2310,In_2395,In_289);
xnor U2311 (N_2311,In_923,In_649);
or U2312 (N_2312,In_2476,In_2119);
xor U2313 (N_2313,In_441,In_1160);
or U2314 (N_2314,In_91,In_2173);
nor U2315 (N_2315,In_951,In_175);
or U2316 (N_2316,In_845,In_365);
nand U2317 (N_2317,In_2423,In_702);
nand U2318 (N_2318,In_1598,In_1997);
nand U2319 (N_2319,In_220,In_1974);
nor U2320 (N_2320,In_567,In_2391);
nor U2321 (N_2321,In_1791,In_2009);
and U2322 (N_2322,In_442,In_1710);
nor U2323 (N_2323,In_1296,In_1024);
nor U2324 (N_2324,In_1268,In_1608);
nand U2325 (N_2325,In_762,In_484);
xor U2326 (N_2326,In_1458,In_178);
and U2327 (N_2327,In_2332,In_2202);
nor U2328 (N_2328,In_1161,In_794);
or U2329 (N_2329,In_2248,In_1864);
nor U2330 (N_2330,In_1551,In_2111);
and U2331 (N_2331,In_1022,In_286);
xnor U2332 (N_2332,In_1814,In_434);
nand U2333 (N_2333,In_1472,In_2342);
or U2334 (N_2334,In_533,In_2153);
nand U2335 (N_2335,In_416,In_1292);
xnor U2336 (N_2336,In_282,In_2146);
xor U2337 (N_2337,In_1427,In_1642);
or U2338 (N_2338,In_2107,In_2416);
nand U2339 (N_2339,In_800,In_603);
nand U2340 (N_2340,In_2359,In_1952);
xor U2341 (N_2341,In_582,In_884);
xor U2342 (N_2342,In_1463,In_570);
nor U2343 (N_2343,In_1485,In_2363);
or U2344 (N_2344,In_96,In_455);
nand U2345 (N_2345,In_623,In_1923);
nor U2346 (N_2346,In_2313,In_2210);
nand U2347 (N_2347,In_1276,In_446);
nor U2348 (N_2348,In_186,In_389);
nand U2349 (N_2349,In_788,In_1022);
or U2350 (N_2350,In_933,In_364);
nor U2351 (N_2351,In_111,In_185);
xnor U2352 (N_2352,In_646,In_102);
nand U2353 (N_2353,In_260,In_90);
or U2354 (N_2354,In_2268,In_2437);
or U2355 (N_2355,In_1751,In_1655);
and U2356 (N_2356,In_321,In_2229);
xor U2357 (N_2357,In_577,In_133);
and U2358 (N_2358,In_1150,In_1259);
xor U2359 (N_2359,In_437,In_584);
or U2360 (N_2360,In_1207,In_968);
xnor U2361 (N_2361,In_546,In_1810);
nand U2362 (N_2362,In_656,In_2167);
or U2363 (N_2363,In_504,In_1434);
or U2364 (N_2364,In_2326,In_2398);
nand U2365 (N_2365,In_353,In_1000);
or U2366 (N_2366,In_2418,In_846);
or U2367 (N_2367,In_698,In_1691);
nand U2368 (N_2368,In_1119,In_482);
or U2369 (N_2369,In_791,In_1072);
nand U2370 (N_2370,In_141,In_1470);
nor U2371 (N_2371,In_1614,In_1585);
nand U2372 (N_2372,In_1264,In_1729);
or U2373 (N_2373,In_403,In_924);
nor U2374 (N_2374,In_1800,In_1111);
or U2375 (N_2375,In_630,In_3);
nand U2376 (N_2376,In_837,In_2471);
nor U2377 (N_2377,In_101,In_2178);
or U2378 (N_2378,In_48,In_2169);
and U2379 (N_2379,In_144,In_353);
xor U2380 (N_2380,In_679,In_563);
xor U2381 (N_2381,In_229,In_2472);
nor U2382 (N_2382,In_2376,In_617);
nor U2383 (N_2383,In_1782,In_864);
or U2384 (N_2384,In_221,In_328);
nand U2385 (N_2385,In_1945,In_783);
or U2386 (N_2386,In_2380,In_2322);
xnor U2387 (N_2387,In_149,In_1975);
or U2388 (N_2388,In_1505,In_242);
nor U2389 (N_2389,In_508,In_1471);
xnor U2390 (N_2390,In_428,In_1647);
or U2391 (N_2391,In_986,In_1428);
nand U2392 (N_2392,In_1752,In_1843);
and U2393 (N_2393,In_557,In_2234);
xor U2394 (N_2394,In_1333,In_487);
nand U2395 (N_2395,In_1166,In_2449);
and U2396 (N_2396,In_1899,In_596);
or U2397 (N_2397,In_2020,In_610);
xor U2398 (N_2398,In_1526,In_280);
xor U2399 (N_2399,In_1543,In_1265);
and U2400 (N_2400,In_2041,In_2289);
nand U2401 (N_2401,In_1154,In_2448);
or U2402 (N_2402,In_465,In_1579);
and U2403 (N_2403,In_1315,In_1678);
nand U2404 (N_2404,In_2297,In_475);
or U2405 (N_2405,In_1026,In_1924);
or U2406 (N_2406,In_2082,In_1254);
nand U2407 (N_2407,In_712,In_2282);
nand U2408 (N_2408,In_697,In_594);
and U2409 (N_2409,In_2269,In_2055);
nand U2410 (N_2410,In_1121,In_2299);
and U2411 (N_2411,In_1011,In_2150);
nor U2412 (N_2412,In_1555,In_490);
nand U2413 (N_2413,In_121,In_958);
xnor U2414 (N_2414,In_1175,In_1271);
or U2415 (N_2415,In_2109,In_885);
and U2416 (N_2416,In_449,In_2330);
xor U2417 (N_2417,In_116,In_118);
or U2418 (N_2418,In_1473,In_1923);
and U2419 (N_2419,In_689,In_52);
and U2420 (N_2420,In_325,In_1957);
xor U2421 (N_2421,In_1865,In_2247);
nor U2422 (N_2422,In_312,In_1317);
and U2423 (N_2423,In_1669,In_1535);
xor U2424 (N_2424,In_1359,In_2147);
nand U2425 (N_2425,In_1857,In_1620);
and U2426 (N_2426,In_1399,In_1267);
xnor U2427 (N_2427,In_2479,In_1471);
or U2428 (N_2428,In_989,In_446);
xor U2429 (N_2429,In_65,In_2051);
nand U2430 (N_2430,In_2097,In_1033);
and U2431 (N_2431,In_1230,In_267);
nor U2432 (N_2432,In_2334,In_493);
and U2433 (N_2433,In_1438,In_536);
xor U2434 (N_2434,In_1899,In_473);
xnor U2435 (N_2435,In_502,In_2400);
xor U2436 (N_2436,In_488,In_141);
and U2437 (N_2437,In_1647,In_1827);
nor U2438 (N_2438,In_753,In_1884);
nand U2439 (N_2439,In_790,In_800);
or U2440 (N_2440,In_493,In_666);
nor U2441 (N_2441,In_361,In_155);
and U2442 (N_2442,In_122,In_658);
and U2443 (N_2443,In_787,In_1835);
xnor U2444 (N_2444,In_2154,In_1991);
or U2445 (N_2445,In_207,In_1377);
and U2446 (N_2446,In_1357,In_808);
nand U2447 (N_2447,In_2066,In_1578);
and U2448 (N_2448,In_2189,In_2310);
nor U2449 (N_2449,In_1784,In_1175);
xnor U2450 (N_2450,In_829,In_1356);
and U2451 (N_2451,In_1624,In_1239);
nor U2452 (N_2452,In_204,In_1223);
nor U2453 (N_2453,In_2362,In_27);
or U2454 (N_2454,In_2337,In_484);
nand U2455 (N_2455,In_2382,In_319);
and U2456 (N_2456,In_151,In_1134);
nand U2457 (N_2457,In_2277,In_333);
or U2458 (N_2458,In_1162,In_1530);
xnor U2459 (N_2459,In_1340,In_157);
nand U2460 (N_2460,In_1632,In_901);
xnor U2461 (N_2461,In_1450,In_2417);
xor U2462 (N_2462,In_1841,In_1252);
xnor U2463 (N_2463,In_1455,In_2412);
xnor U2464 (N_2464,In_720,In_1337);
or U2465 (N_2465,In_2455,In_1136);
and U2466 (N_2466,In_1585,In_2098);
nand U2467 (N_2467,In_129,In_894);
or U2468 (N_2468,In_1125,In_491);
nand U2469 (N_2469,In_2273,In_1523);
nor U2470 (N_2470,In_2478,In_2219);
and U2471 (N_2471,In_2216,In_2392);
or U2472 (N_2472,In_1254,In_385);
nand U2473 (N_2473,In_2231,In_31);
nor U2474 (N_2474,In_2032,In_2285);
nand U2475 (N_2475,In_1791,In_987);
nor U2476 (N_2476,In_1661,In_1388);
and U2477 (N_2477,In_2485,In_1971);
nand U2478 (N_2478,In_2323,In_1753);
and U2479 (N_2479,In_954,In_601);
nand U2480 (N_2480,In_2038,In_1697);
and U2481 (N_2481,In_598,In_368);
nand U2482 (N_2482,In_2314,In_1413);
nand U2483 (N_2483,In_1775,In_533);
xor U2484 (N_2484,In_2104,In_2132);
xor U2485 (N_2485,In_2181,In_752);
or U2486 (N_2486,In_171,In_560);
nor U2487 (N_2487,In_706,In_1164);
xor U2488 (N_2488,In_1557,In_296);
and U2489 (N_2489,In_1037,In_78);
or U2490 (N_2490,In_395,In_731);
nor U2491 (N_2491,In_60,In_977);
xnor U2492 (N_2492,In_1572,In_1225);
or U2493 (N_2493,In_1328,In_2220);
xor U2494 (N_2494,In_212,In_107);
and U2495 (N_2495,In_1473,In_326);
nand U2496 (N_2496,In_2040,In_1823);
nor U2497 (N_2497,In_2311,In_2333);
xor U2498 (N_2498,In_553,In_2252);
xor U2499 (N_2499,In_2150,In_619);
xor U2500 (N_2500,In_999,In_1561);
or U2501 (N_2501,In_1562,In_13);
xor U2502 (N_2502,In_1143,In_1955);
xor U2503 (N_2503,In_2427,In_79);
or U2504 (N_2504,In_1148,In_2404);
and U2505 (N_2505,In_1047,In_1182);
and U2506 (N_2506,In_2384,In_2460);
nor U2507 (N_2507,In_429,In_1970);
xnor U2508 (N_2508,In_1822,In_1552);
xnor U2509 (N_2509,In_308,In_2188);
or U2510 (N_2510,In_1666,In_2478);
or U2511 (N_2511,In_289,In_1065);
nor U2512 (N_2512,In_549,In_2420);
nor U2513 (N_2513,In_1780,In_2375);
xnor U2514 (N_2514,In_1346,In_136);
xnor U2515 (N_2515,In_203,In_52);
or U2516 (N_2516,In_609,In_2097);
nand U2517 (N_2517,In_449,In_1631);
nor U2518 (N_2518,In_1410,In_552);
nor U2519 (N_2519,In_1378,In_1952);
nor U2520 (N_2520,In_1040,In_2058);
nand U2521 (N_2521,In_1926,In_2492);
nand U2522 (N_2522,In_1582,In_698);
and U2523 (N_2523,In_388,In_2418);
or U2524 (N_2524,In_993,In_2307);
nor U2525 (N_2525,In_1985,In_2051);
and U2526 (N_2526,In_1678,In_826);
nor U2527 (N_2527,In_778,In_1717);
xnor U2528 (N_2528,In_1519,In_1627);
xnor U2529 (N_2529,In_1151,In_138);
nand U2530 (N_2530,In_261,In_1344);
and U2531 (N_2531,In_1311,In_1404);
xor U2532 (N_2532,In_1155,In_1998);
or U2533 (N_2533,In_2184,In_1324);
nand U2534 (N_2534,In_786,In_2168);
nor U2535 (N_2535,In_1905,In_2232);
and U2536 (N_2536,In_1152,In_2398);
nor U2537 (N_2537,In_672,In_1659);
xnor U2538 (N_2538,In_417,In_1447);
nor U2539 (N_2539,In_755,In_1343);
or U2540 (N_2540,In_1444,In_1689);
and U2541 (N_2541,In_558,In_1658);
xnor U2542 (N_2542,In_1159,In_509);
nand U2543 (N_2543,In_2477,In_2248);
nand U2544 (N_2544,In_1531,In_2038);
nor U2545 (N_2545,In_215,In_325);
nand U2546 (N_2546,In_653,In_581);
nand U2547 (N_2547,In_2307,In_200);
nor U2548 (N_2548,In_1413,In_818);
nor U2549 (N_2549,In_1755,In_414);
xor U2550 (N_2550,In_2395,In_941);
and U2551 (N_2551,In_165,In_1473);
nor U2552 (N_2552,In_2431,In_1491);
and U2553 (N_2553,In_1755,In_313);
or U2554 (N_2554,In_1972,In_2214);
xnor U2555 (N_2555,In_2454,In_933);
or U2556 (N_2556,In_341,In_713);
xor U2557 (N_2557,In_233,In_1305);
xnor U2558 (N_2558,In_1622,In_994);
and U2559 (N_2559,In_812,In_34);
or U2560 (N_2560,In_874,In_2430);
nor U2561 (N_2561,In_2450,In_742);
or U2562 (N_2562,In_1035,In_1259);
or U2563 (N_2563,In_995,In_768);
and U2564 (N_2564,In_1982,In_1431);
nand U2565 (N_2565,In_629,In_911);
xnor U2566 (N_2566,In_2435,In_2010);
nand U2567 (N_2567,In_2340,In_1426);
nand U2568 (N_2568,In_397,In_494);
or U2569 (N_2569,In_381,In_1807);
nand U2570 (N_2570,In_1193,In_44);
and U2571 (N_2571,In_896,In_2063);
nor U2572 (N_2572,In_1145,In_231);
and U2573 (N_2573,In_816,In_2218);
and U2574 (N_2574,In_2210,In_1916);
or U2575 (N_2575,In_2391,In_1805);
or U2576 (N_2576,In_1513,In_2315);
nor U2577 (N_2577,In_1966,In_334);
xnor U2578 (N_2578,In_1838,In_2229);
and U2579 (N_2579,In_1929,In_2453);
xor U2580 (N_2580,In_294,In_681);
nand U2581 (N_2581,In_104,In_1956);
xnor U2582 (N_2582,In_493,In_1608);
and U2583 (N_2583,In_1431,In_1401);
nor U2584 (N_2584,In_1968,In_825);
or U2585 (N_2585,In_1837,In_210);
xor U2586 (N_2586,In_448,In_2484);
and U2587 (N_2587,In_1472,In_1780);
xor U2588 (N_2588,In_1565,In_1865);
nor U2589 (N_2589,In_310,In_2382);
xnor U2590 (N_2590,In_1548,In_1610);
nand U2591 (N_2591,In_1602,In_2408);
nand U2592 (N_2592,In_1728,In_582);
nor U2593 (N_2593,In_1250,In_1172);
nor U2594 (N_2594,In_1633,In_1122);
xor U2595 (N_2595,In_1031,In_348);
and U2596 (N_2596,In_2470,In_1168);
nor U2597 (N_2597,In_927,In_43);
or U2598 (N_2598,In_2014,In_1157);
or U2599 (N_2599,In_374,In_267);
and U2600 (N_2600,In_2498,In_454);
or U2601 (N_2601,In_1787,In_1821);
or U2602 (N_2602,In_1441,In_2092);
nor U2603 (N_2603,In_546,In_2000);
xor U2604 (N_2604,In_2422,In_2389);
and U2605 (N_2605,In_1519,In_1319);
nand U2606 (N_2606,In_887,In_1403);
nor U2607 (N_2607,In_1282,In_1437);
or U2608 (N_2608,In_1948,In_1607);
and U2609 (N_2609,In_989,In_789);
xnor U2610 (N_2610,In_1966,In_382);
xor U2611 (N_2611,In_596,In_2384);
nand U2612 (N_2612,In_878,In_1441);
nand U2613 (N_2613,In_723,In_1572);
nand U2614 (N_2614,In_121,In_2228);
nor U2615 (N_2615,In_2402,In_978);
nand U2616 (N_2616,In_939,In_1373);
or U2617 (N_2617,In_1053,In_130);
or U2618 (N_2618,In_517,In_73);
and U2619 (N_2619,In_1214,In_1680);
and U2620 (N_2620,In_1874,In_792);
or U2621 (N_2621,In_2248,In_2463);
nand U2622 (N_2622,In_1117,In_2488);
nand U2623 (N_2623,In_812,In_340);
nor U2624 (N_2624,In_1281,In_2289);
xor U2625 (N_2625,In_2395,In_979);
nand U2626 (N_2626,In_1787,In_2278);
nor U2627 (N_2627,In_1247,In_1752);
xor U2628 (N_2628,In_1251,In_1537);
or U2629 (N_2629,In_2357,In_2042);
and U2630 (N_2630,In_849,In_1469);
nand U2631 (N_2631,In_1602,In_600);
nand U2632 (N_2632,In_627,In_2332);
nor U2633 (N_2633,In_1104,In_345);
and U2634 (N_2634,In_252,In_1297);
nand U2635 (N_2635,In_946,In_877);
nand U2636 (N_2636,In_1290,In_769);
nor U2637 (N_2637,In_862,In_1385);
nand U2638 (N_2638,In_2341,In_871);
or U2639 (N_2639,In_1591,In_520);
nor U2640 (N_2640,In_353,In_2375);
or U2641 (N_2641,In_1974,In_324);
or U2642 (N_2642,In_894,In_224);
or U2643 (N_2643,In_1283,In_1575);
or U2644 (N_2644,In_435,In_189);
nand U2645 (N_2645,In_870,In_273);
or U2646 (N_2646,In_1881,In_153);
and U2647 (N_2647,In_1586,In_668);
nand U2648 (N_2648,In_236,In_865);
nand U2649 (N_2649,In_675,In_42);
xnor U2650 (N_2650,In_1735,In_1832);
and U2651 (N_2651,In_2291,In_1280);
nand U2652 (N_2652,In_2444,In_2467);
and U2653 (N_2653,In_272,In_2244);
or U2654 (N_2654,In_1668,In_2033);
nor U2655 (N_2655,In_1733,In_1969);
or U2656 (N_2656,In_1298,In_2136);
or U2657 (N_2657,In_1295,In_152);
xor U2658 (N_2658,In_1622,In_1807);
nand U2659 (N_2659,In_2111,In_33);
xnor U2660 (N_2660,In_2274,In_1503);
xnor U2661 (N_2661,In_1221,In_808);
nand U2662 (N_2662,In_1787,In_1512);
xor U2663 (N_2663,In_1497,In_2188);
or U2664 (N_2664,In_623,In_1560);
nor U2665 (N_2665,In_810,In_710);
nor U2666 (N_2666,In_1530,In_822);
nor U2667 (N_2667,In_296,In_65);
nand U2668 (N_2668,In_1920,In_1684);
nor U2669 (N_2669,In_405,In_1143);
and U2670 (N_2670,In_158,In_1130);
nor U2671 (N_2671,In_2292,In_2055);
and U2672 (N_2672,In_924,In_1165);
nor U2673 (N_2673,In_1589,In_944);
and U2674 (N_2674,In_1838,In_2432);
xnor U2675 (N_2675,In_2076,In_916);
nor U2676 (N_2676,In_2093,In_1767);
xnor U2677 (N_2677,In_307,In_2493);
and U2678 (N_2678,In_2005,In_410);
and U2679 (N_2679,In_1243,In_374);
xor U2680 (N_2680,In_2207,In_750);
or U2681 (N_2681,In_246,In_106);
or U2682 (N_2682,In_2331,In_519);
nand U2683 (N_2683,In_953,In_662);
xnor U2684 (N_2684,In_1726,In_242);
or U2685 (N_2685,In_479,In_698);
or U2686 (N_2686,In_1725,In_666);
nor U2687 (N_2687,In_1525,In_1328);
nand U2688 (N_2688,In_628,In_982);
xnor U2689 (N_2689,In_1510,In_436);
and U2690 (N_2690,In_1464,In_1364);
xor U2691 (N_2691,In_1442,In_81);
nor U2692 (N_2692,In_639,In_1221);
xnor U2693 (N_2693,In_847,In_2192);
and U2694 (N_2694,In_1795,In_2250);
nor U2695 (N_2695,In_419,In_2051);
nor U2696 (N_2696,In_2124,In_353);
and U2697 (N_2697,In_2127,In_507);
nor U2698 (N_2698,In_1720,In_1650);
nor U2699 (N_2699,In_2127,In_1633);
xor U2700 (N_2700,In_1899,In_979);
nor U2701 (N_2701,In_2000,In_1037);
or U2702 (N_2702,In_2225,In_560);
nor U2703 (N_2703,In_440,In_575);
xnor U2704 (N_2704,In_1122,In_856);
xor U2705 (N_2705,In_442,In_1920);
or U2706 (N_2706,In_1364,In_1372);
nand U2707 (N_2707,In_0,In_1853);
and U2708 (N_2708,In_774,In_1523);
and U2709 (N_2709,In_2133,In_306);
nand U2710 (N_2710,In_1105,In_1975);
or U2711 (N_2711,In_2324,In_1887);
xnor U2712 (N_2712,In_436,In_1978);
nand U2713 (N_2713,In_1451,In_1294);
xor U2714 (N_2714,In_2324,In_354);
nand U2715 (N_2715,In_1915,In_1244);
nand U2716 (N_2716,In_2029,In_2188);
nand U2717 (N_2717,In_186,In_1290);
nor U2718 (N_2718,In_2116,In_2399);
or U2719 (N_2719,In_1290,In_693);
or U2720 (N_2720,In_277,In_1208);
nand U2721 (N_2721,In_550,In_2322);
or U2722 (N_2722,In_837,In_2343);
nor U2723 (N_2723,In_698,In_1209);
nand U2724 (N_2724,In_231,In_1364);
xor U2725 (N_2725,In_590,In_1938);
and U2726 (N_2726,In_557,In_1056);
nand U2727 (N_2727,In_2301,In_1794);
or U2728 (N_2728,In_212,In_1717);
or U2729 (N_2729,In_1230,In_1077);
and U2730 (N_2730,In_340,In_2293);
nor U2731 (N_2731,In_2091,In_267);
or U2732 (N_2732,In_2359,In_1701);
or U2733 (N_2733,In_770,In_1756);
nor U2734 (N_2734,In_1011,In_927);
nor U2735 (N_2735,In_1959,In_506);
and U2736 (N_2736,In_952,In_583);
nor U2737 (N_2737,In_162,In_455);
nor U2738 (N_2738,In_840,In_859);
nor U2739 (N_2739,In_327,In_2291);
and U2740 (N_2740,In_343,In_1198);
nor U2741 (N_2741,In_1562,In_1903);
nand U2742 (N_2742,In_1928,In_966);
or U2743 (N_2743,In_261,In_1675);
nand U2744 (N_2744,In_2044,In_1525);
nor U2745 (N_2745,In_1536,In_2013);
xor U2746 (N_2746,In_381,In_487);
and U2747 (N_2747,In_1492,In_694);
xor U2748 (N_2748,In_834,In_874);
nand U2749 (N_2749,In_388,In_42);
nor U2750 (N_2750,In_2138,In_1466);
nand U2751 (N_2751,In_1729,In_1869);
or U2752 (N_2752,In_350,In_802);
nand U2753 (N_2753,In_560,In_364);
or U2754 (N_2754,In_1787,In_1400);
and U2755 (N_2755,In_170,In_138);
and U2756 (N_2756,In_1017,In_1463);
xnor U2757 (N_2757,In_1717,In_2299);
xor U2758 (N_2758,In_1847,In_1887);
xor U2759 (N_2759,In_1368,In_893);
or U2760 (N_2760,In_2058,In_2372);
xnor U2761 (N_2761,In_154,In_517);
or U2762 (N_2762,In_872,In_1652);
or U2763 (N_2763,In_2050,In_73);
xnor U2764 (N_2764,In_758,In_2344);
and U2765 (N_2765,In_753,In_943);
xor U2766 (N_2766,In_2341,In_2393);
nand U2767 (N_2767,In_1808,In_1024);
nand U2768 (N_2768,In_1792,In_579);
nor U2769 (N_2769,In_1431,In_910);
or U2770 (N_2770,In_2141,In_355);
nand U2771 (N_2771,In_465,In_2046);
and U2772 (N_2772,In_2194,In_514);
nor U2773 (N_2773,In_740,In_2135);
and U2774 (N_2774,In_2158,In_722);
xor U2775 (N_2775,In_1124,In_2131);
xor U2776 (N_2776,In_919,In_1547);
or U2777 (N_2777,In_1441,In_2140);
nor U2778 (N_2778,In_464,In_1819);
and U2779 (N_2779,In_876,In_2310);
nand U2780 (N_2780,In_2296,In_2166);
and U2781 (N_2781,In_1874,In_1038);
or U2782 (N_2782,In_1774,In_1342);
nand U2783 (N_2783,In_2248,In_38);
nor U2784 (N_2784,In_93,In_1330);
xnor U2785 (N_2785,In_513,In_436);
and U2786 (N_2786,In_1405,In_2474);
and U2787 (N_2787,In_1985,In_1560);
nand U2788 (N_2788,In_982,In_1431);
xnor U2789 (N_2789,In_43,In_1997);
or U2790 (N_2790,In_2309,In_1762);
xnor U2791 (N_2791,In_14,In_1714);
nand U2792 (N_2792,In_2386,In_1227);
nand U2793 (N_2793,In_2393,In_1804);
xnor U2794 (N_2794,In_407,In_1364);
and U2795 (N_2795,In_1086,In_1631);
xor U2796 (N_2796,In_842,In_865);
or U2797 (N_2797,In_45,In_1898);
or U2798 (N_2798,In_1655,In_2452);
nor U2799 (N_2799,In_539,In_86);
nor U2800 (N_2800,In_1403,In_2190);
or U2801 (N_2801,In_897,In_655);
or U2802 (N_2802,In_2265,In_2082);
nand U2803 (N_2803,In_1495,In_2023);
nand U2804 (N_2804,In_844,In_858);
nand U2805 (N_2805,In_802,In_473);
nor U2806 (N_2806,In_85,In_1207);
or U2807 (N_2807,In_1902,In_278);
nor U2808 (N_2808,In_2049,In_59);
nand U2809 (N_2809,In_1883,In_1166);
xor U2810 (N_2810,In_1364,In_1948);
xnor U2811 (N_2811,In_797,In_2403);
and U2812 (N_2812,In_2176,In_1053);
or U2813 (N_2813,In_1189,In_1745);
nor U2814 (N_2814,In_1371,In_253);
xnor U2815 (N_2815,In_165,In_2240);
nor U2816 (N_2816,In_1263,In_7);
nand U2817 (N_2817,In_2390,In_33);
and U2818 (N_2818,In_2428,In_1546);
and U2819 (N_2819,In_2209,In_668);
nor U2820 (N_2820,In_1681,In_1809);
and U2821 (N_2821,In_1899,In_564);
or U2822 (N_2822,In_1893,In_2003);
nor U2823 (N_2823,In_1788,In_1973);
or U2824 (N_2824,In_1857,In_22);
nor U2825 (N_2825,In_1400,In_2335);
nand U2826 (N_2826,In_156,In_2201);
xnor U2827 (N_2827,In_2042,In_1486);
and U2828 (N_2828,In_2063,In_2044);
or U2829 (N_2829,In_1343,In_1504);
nand U2830 (N_2830,In_998,In_1965);
or U2831 (N_2831,In_1938,In_2174);
nand U2832 (N_2832,In_1841,In_2122);
nor U2833 (N_2833,In_1865,In_2124);
nor U2834 (N_2834,In_931,In_1243);
or U2835 (N_2835,In_1779,In_1838);
and U2836 (N_2836,In_1830,In_1999);
and U2837 (N_2837,In_1810,In_1304);
nor U2838 (N_2838,In_84,In_1461);
xnor U2839 (N_2839,In_312,In_95);
xor U2840 (N_2840,In_1949,In_1491);
or U2841 (N_2841,In_1959,In_552);
and U2842 (N_2842,In_371,In_769);
nand U2843 (N_2843,In_884,In_2445);
or U2844 (N_2844,In_604,In_1299);
nor U2845 (N_2845,In_2282,In_885);
and U2846 (N_2846,In_1295,In_2362);
nand U2847 (N_2847,In_732,In_1669);
and U2848 (N_2848,In_1075,In_1689);
nor U2849 (N_2849,In_579,In_2289);
or U2850 (N_2850,In_277,In_2058);
nand U2851 (N_2851,In_381,In_1026);
or U2852 (N_2852,In_1611,In_1084);
nand U2853 (N_2853,In_79,In_482);
and U2854 (N_2854,In_355,In_2183);
nand U2855 (N_2855,In_2319,In_100);
nor U2856 (N_2856,In_346,In_1105);
xor U2857 (N_2857,In_768,In_1521);
xor U2858 (N_2858,In_1035,In_1127);
or U2859 (N_2859,In_1504,In_1148);
and U2860 (N_2860,In_785,In_1985);
nand U2861 (N_2861,In_2342,In_1326);
or U2862 (N_2862,In_1870,In_1945);
and U2863 (N_2863,In_469,In_2431);
nor U2864 (N_2864,In_519,In_2348);
xnor U2865 (N_2865,In_277,In_1821);
nand U2866 (N_2866,In_2089,In_2213);
and U2867 (N_2867,In_423,In_1683);
nor U2868 (N_2868,In_1999,In_1813);
or U2869 (N_2869,In_2060,In_744);
nor U2870 (N_2870,In_993,In_1381);
xnor U2871 (N_2871,In_2252,In_145);
nand U2872 (N_2872,In_1768,In_1380);
nand U2873 (N_2873,In_1108,In_265);
or U2874 (N_2874,In_1823,In_2034);
and U2875 (N_2875,In_368,In_1913);
nand U2876 (N_2876,In_1095,In_469);
or U2877 (N_2877,In_1884,In_1492);
xnor U2878 (N_2878,In_1200,In_313);
xnor U2879 (N_2879,In_1605,In_307);
or U2880 (N_2880,In_1722,In_1925);
nor U2881 (N_2881,In_1863,In_1048);
nor U2882 (N_2882,In_1778,In_1439);
xor U2883 (N_2883,In_1567,In_1608);
nor U2884 (N_2884,In_1562,In_645);
and U2885 (N_2885,In_1274,In_1329);
or U2886 (N_2886,In_2092,In_690);
or U2887 (N_2887,In_1821,In_264);
and U2888 (N_2888,In_1635,In_1643);
or U2889 (N_2889,In_117,In_1865);
and U2890 (N_2890,In_562,In_912);
nor U2891 (N_2891,In_2204,In_1043);
and U2892 (N_2892,In_161,In_32);
nor U2893 (N_2893,In_2088,In_1714);
nor U2894 (N_2894,In_1829,In_786);
xor U2895 (N_2895,In_2346,In_1552);
or U2896 (N_2896,In_964,In_152);
xor U2897 (N_2897,In_335,In_321);
nand U2898 (N_2898,In_755,In_526);
xnor U2899 (N_2899,In_626,In_1286);
and U2900 (N_2900,In_1987,In_895);
xor U2901 (N_2901,In_1701,In_318);
and U2902 (N_2902,In_398,In_1415);
and U2903 (N_2903,In_2378,In_1619);
and U2904 (N_2904,In_2244,In_1901);
xor U2905 (N_2905,In_1933,In_2488);
or U2906 (N_2906,In_2264,In_1656);
xnor U2907 (N_2907,In_352,In_144);
xor U2908 (N_2908,In_344,In_1249);
and U2909 (N_2909,In_2469,In_892);
and U2910 (N_2910,In_481,In_1572);
xor U2911 (N_2911,In_148,In_1641);
nand U2912 (N_2912,In_2066,In_2147);
or U2913 (N_2913,In_261,In_940);
xnor U2914 (N_2914,In_1145,In_1428);
nor U2915 (N_2915,In_1803,In_231);
or U2916 (N_2916,In_1310,In_1315);
nor U2917 (N_2917,In_2433,In_981);
nor U2918 (N_2918,In_2280,In_139);
xnor U2919 (N_2919,In_1246,In_522);
nor U2920 (N_2920,In_196,In_2267);
nand U2921 (N_2921,In_2372,In_1785);
or U2922 (N_2922,In_2329,In_670);
and U2923 (N_2923,In_1258,In_1587);
and U2924 (N_2924,In_545,In_738);
and U2925 (N_2925,In_451,In_418);
or U2926 (N_2926,In_1728,In_1794);
nand U2927 (N_2927,In_2240,In_1308);
nand U2928 (N_2928,In_1761,In_2489);
nand U2929 (N_2929,In_468,In_1751);
nand U2930 (N_2930,In_1476,In_1300);
nand U2931 (N_2931,In_708,In_2407);
nand U2932 (N_2932,In_1504,In_571);
and U2933 (N_2933,In_2305,In_215);
nand U2934 (N_2934,In_96,In_1800);
nor U2935 (N_2935,In_2232,In_25);
or U2936 (N_2936,In_1699,In_911);
or U2937 (N_2937,In_290,In_1212);
xor U2938 (N_2938,In_264,In_727);
and U2939 (N_2939,In_1696,In_1857);
nor U2940 (N_2940,In_4,In_1260);
nor U2941 (N_2941,In_150,In_1785);
nor U2942 (N_2942,In_116,In_1315);
nand U2943 (N_2943,In_1895,In_162);
nand U2944 (N_2944,In_1384,In_1504);
nand U2945 (N_2945,In_1235,In_1960);
xor U2946 (N_2946,In_2367,In_1967);
xor U2947 (N_2947,In_2260,In_766);
and U2948 (N_2948,In_1188,In_2073);
or U2949 (N_2949,In_61,In_1184);
and U2950 (N_2950,In_1950,In_2098);
xor U2951 (N_2951,In_1412,In_1694);
or U2952 (N_2952,In_733,In_1340);
or U2953 (N_2953,In_2196,In_1752);
xor U2954 (N_2954,In_153,In_2083);
and U2955 (N_2955,In_1427,In_2461);
or U2956 (N_2956,In_293,In_551);
nand U2957 (N_2957,In_1572,In_1682);
xor U2958 (N_2958,In_1611,In_2180);
nand U2959 (N_2959,In_280,In_1206);
or U2960 (N_2960,In_223,In_1354);
nand U2961 (N_2961,In_2237,In_547);
xnor U2962 (N_2962,In_923,In_2240);
and U2963 (N_2963,In_1997,In_2443);
or U2964 (N_2964,In_947,In_817);
nand U2965 (N_2965,In_1475,In_1511);
nand U2966 (N_2966,In_88,In_1788);
nand U2967 (N_2967,In_758,In_573);
and U2968 (N_2968,In_2217,In_837);
and U2969 (N_2969,In_1194,In_272);
xor U2970 (N_2970,In_1079,In_1331);
nand U2971 (N_2971,In_1290,In_998);
nor U2972 (N_2972,In_750,In_1663);
and U2973 (N_2973,In_2393,In_578);
nand U2974 (N_2974,In_1317,In_799);
xnor U2975 (N_2975,In_99,In_1248);
or U2976 (N_2976,In_1713,In_385);
nand U2977 (N_2977,In_2151,In_1828);
or U2978 (N_2978,In_1028,In_449);
nand U2979 (N_2979,In_245,In_1926);
nand U2980 (N_2980,In_1490,In_1067);
or U2981 (N_2981,In_1097,In_840);
or U2982 (N_2982,In_1301,In_2300);
nor U2983 (N_2983,In_1454,In_2430);
nand U2984 (N_2984,In_812,In_159);
or U2985 (N_2985,In_907,In_590);
xnor U2986 (N_2986,In_353,In_2327);
nand U2987 (N_2987,In_1044,In_1435);
xnor U2988 (N_2988,In_1831,In_1459);
nand U2989 (N_2989,In_2035,In_965);
nor U2990 (N_2990,In_578,In_1164);
and U2991 (N_2991,In_2248,In_2102);
and U2992 (N_2992,In_1866,In_1986);
and U2993 (N_2993,In_2429,In_1872);
xnor U2994 (N_2994,In_750,In_1629);
or U2995 (N_2995,In_726,In_2162);
or U2996 (N_2996,In_1669,In_2208);
xnor U2997 (N_2997,In_1955,In_1916);
xor U2998 (N_2998,In_2233,In_203);
nand U2999 (N_2999,In_1071,In_2152);
and U3000 (N_3000,In_575,In_180);
nand U3001 (N_3001,In_793,In_1097);
or U3002 (N_3002,In_1985,In_355);
and U3003 (N_3003,In_2037,In_1619);
xnor U3004 (N_3004,In_2400,In_2496);
and U3005 (N_3005,In_2402,In_2261);
nor U3006 (N_3006,In_1272,In_112);
and U3007 (N_3007,In_2229,In_1266);
nand U3008 (N_3008,In_452,In_357);
or U3009 (N_3009,In_1548,In_348);
or U3010 (N_3010,In_849,In_924);
nand U3011 (N_3011,In_1742,In_2024);
xor U3012 (N_3012,In_2456,In_1562);
nor U3013 (N_3013,In_2405,In_333);
and U3014 (N_3014,In_1043,In_1009);
nand U3015 (N_3015,In_114,In_1773);
and U3016 (N_3016,In_225,In_1757);
nand U3017 (N_3017,In_90,In_1610);
nand U3018 (N_3018,In_1479,In_1654);
nor U3019 (N_3019,In_1732,In_2278);
nor U3020 (N_3020,In_2221,In_264);
nand U3021 (N_3021,In_180,In_1784);
and U3022 (N_3022,In_1167,In_1682);
or U3023 (N_3023,In_1240,In_478);
xor U3024 (N_3024,In_166,In_1353);
xor U3025 (N_3025,In_2168,In_1416);
nand U3026 (N_3026,In_1966,In_114);
and U3027 (N_3027,In_150,In_170);
nor U3028 (N_3028,In_301,In_2317);
nor U3029 (N_3029,In_2071,In_1147);
and U3030 (N_3030,In_2073,In_1901);
nor U3031 (N_3031,In_805,In_370);
or U3032 (N_3032,In_183,In_1737);
xor U3033 (N_3033,In_2309,In_327);
and U3034 (N_3034,In_1868,In_2461);
and U3035 (N_3035,In_1363,In_547);
xor U3036 (N_3036,In_642,In_1867);
or U3037 (N_3037,In_813,In_80);
xnor U3038 (N_3038,In_398,In_650);
xor U3039 (N_3039,In_1662,In_85);
nor U3040 (N_3040,In_1960,In_1365);
or U3041 (N_3041,In_1446,In_1077);
or U3042 (N_3042,In_2198,In_394);
xor U3043 (N_3043,In_1070,In_679);
nand U3044 (N_3044,In_1875,In_2327);
and U3045 (N_3045,In_748,In_17);
xnor U3046 (N_3046,In_190,In_168);
and U3047 (N_3047,In_1623,In_1760);
and U3048 (N_3048,In_1294,In_250);
nor U3049 (N_3049,In_12,In_1068);
xnor U3050 (N_3050,In_1511,In_156);
xnor U3051 (N_3051,In_1201,In_172);
and U3052 (N_3052,In_1677,In_1814);
or U3053 (N_3053,In_981,In_586);
xnor U3054 (N_3054,In_2026,In_1681);
xor U3055 (N_3055,In_295,In_89);
nor U3056 (N_3056,In_813,In_1981);
and U3057 (N_3057,In_733,In_2222);
nand U3058 (N_3058,In_218,In_361);
or U3059 (N_3059,In_2455,In_874);
nand U3060 (N_3060,In_387,In_2281);
nor U3061 (N_3061,In_596,In_2220);
and U3062 (N_3062,In_949,In_1844);
nand U3063 (N_3063,In_1313,In_72);
or U3064 (N_3064,In_487,In_111);
xor U3065 (N_3065,In_548,In_2097);
or U3066 (N_3066,In_1616,In_183);
and U3067 (N_3067,In_2262,In_2426);
xor U3068 (N_3068,In_1363,In_117);
nor U3069 (N_3069,In_2446,In_1194);
nor U3070 (N_3070,In_1278,In_2469);
and U3071 (N_3071,In_1736,In_1433);
xor U3072 (N_3072,In_1851,In_630);
and U3073 (N_3073,In_2373,In_2460);
xor U3074 (N_3074,In_1035,In_1197);
nand U3075 (N_3075,In_363,In_733);
or U3076 (N_3076,In_305,In_534);
and U3077 (N_3077,In_2066,In_2465);
or U3078 (N_3078,In_1198,In_1225);
and U3079 (N_3079,In_2433,In_685);
xor U3080 (N_3080,In_1436,In_1963);
or U3081 (N_3081,In_1239,In_1429);
xor U3082 (N_3082,In_1263,In_586);
xor U3083 (N_3083,In_2381,In_130);
nand U3084 (N_3084,In_2215,In_948);
nor U3085 (N_3085,In_1921,In_1597);
or U3086 (N_3086,In_2032,In_2188);
or U3087 (N_3087,In_781,In_720);
xor U3088 (N_3088,In_47,In_1924);
xnor U3089 (N_3089,In_442,In_2274);
nand U3090 (N_3090,In_1971,In_1691);
and U3091 (N_3091,In_2052,In_262);
xnor U3092 (N_3092,In_1502,In_2483);
nor U3093 (N_3093,In_2049,In_2295);
nand U3094 (N_3094,In_1277,In_201);
nand U3095 (N_3095,In_516,In_1927);
and U3096 (N_3096,In_580,In_89);
nand U3097 (N_3097,In_1625,In_437);
nor U3098 (N_3098,In_891,In_2259);
xnor U3099 (N_3099,In_735,In_701);
and U3100 (N_3100,In_659,In_2320);
and U3101 (N_3101,In_610,In_1628);
or U3102 (N_3102,In_1877,In_1953);
nand U3103 (N_3103,In_1931,In_117);
xor U3104 (N_3104,In_98,In_2281);
and U3105 (N_3105,In_166,In_933);
or U3106 (N_3106,In_1685,In_705);
xnor U3107 (N_3107,In_1215,In_1368);
or U3108 (N_3108,In_2074,In_745);
nor U3109 (N_3109,In_1863,In_2437);
xnor U3110 (N_3110,In_799,In_786);
nor U3111 (N_3111,In_1255,In_1627);
and U3112 (N_3112,In_765,In_1721);
and U3113 (N_3113,In_1585,In_1259);
or U3114 (N_3114,In_1009,In_1428);
nand U3115 (N_3115,In_352,In_2447);
nand U3116 (N_3116,In_2258,In_1481);
and U3117 (N_3117,In_1531,In_809);
or U3118 (N_3118,In_1627,In_2127);
and U3119 (N_3119,In_1714,In_810);
nand U3120 (N_3120,In_553,In_1021);
nor U3121 (N_3121,In_1811,In_1647);
xnor U3122 (N_3122,In_943,In_2095);
nand U3123 (N_3123,In_870,In_2293);
and U3124 (N_3124,In_2202,In_264);
xnor U3125 (N_3125,In_759,In_699);
nand U3126 (N_3126,In_1880,In_971);
or U3127 (N_3127,In_674,In_2060);
or U3128 (N_3128,In_1490,In_1452);
nand U3129 (N_3129,In_2225,In_2023);
nor U3130 (N_3130,In_1218,In_2403);
xor U3131 (N_3131,In_304,In_1019);
and U3132 (N_3132,In_150,In_1123);
and U3133 (N_3133,In_718,In_706);
nand U3134 (N_3134,In_1524,In_1096);
or U3135 (N_3135,In_447,In_1840);
nor U3136 (N_3136,In_46,In_2486);
nor U3137 (N_3137,In_662,In_2333);
or U3138 (N_3138,In_1857,In_2267);
nor U3139 (N_3139,In_2439,In_573);
or U3140 (N_3140,In_2198,In_21);
xnor U3141 (N_3141,In_206,In_739);
nor U3142 (N_3142,In_1293,In_1098);
and U3143 (N_3143,In_822,In_1282);
nor U3144 (N_3144,In_702,In_651);
xor U3145 (N_3145,In_2387,In_1110);
nor U3146 (N_3146,In_889,In_533);
nor U3147 (N_3147,In_1415,In_82);
or U3148 (N_3148,In_2294,In_1208);
nand U3149 (N_3149,In_898,In_860);
or U3150 (N_3150,In_1913,In_1495);
xnor U3151 (N_3151,In_1809,In_303);
xor U3152 (N_3152,In_1544,In_85);
and U3153 (N_3153,In_1779,In_711);
xor U3154 (N_3154,In_1202,In_2348);
nand U3155 (N_3155,In_2013,In_1405);
xor U3156 (N_3156,In_76,In_1338);
nor U3157 (N_3157,In_1996,In_168);
nor U3158 (N_3158,In_1833,In_395);
and U3159 (N_3159,In_1894,In_2266);
nand U3160 (N_3160,In_449,In_735);
xor U3161 (N_3161,In_157,In_15);
and U3162 (N_3162,In_2119,In_216);
nand U3163 (N_3163,In_1991,In_37);
xor U3164 (N_3164,In_1341,In_2369);
and U3165 (N_3165,In_1542,In_79);
nand U3166 (N_3166,In_601,In_1909);
or U3167 (N_3167,In_1329,In_703);
or U3168 (N_3168,In_576,In_104);
xor U3169 (N_3169,In_1841,In_1987);
xor U3170 (N_3170,In_1222,In_1716);
xor U3171 (N_3171,In_1636,In_1552);
xnor U3172 (N_3172,In_523,In_1947);
nand U3173 (N_3173,In_2102,In_2178);
nand U3174 (N_3174,In_1206,In_755);
nand U3175 (N_3175,In_873,In_1734);
nor U3176 (N_3176,In_1628,In_690);
and U3177 (N_3177,In_335,In_621);
xor U3178 (N_3178,In_1354,In_1174);
or U3179 (N_3179,In_963,In_82);
or U3180 (N_3180,In_1093,In_1708);
and U3181 (N_3181,In_422,In_803);
and U3182 (N_3182,In_1219,In_899);
nand U3183 (N_3183,In_347,In_2352);
xor U3184 (N_3184,In_279,In_1211);
nor U3185 (N_3185,In_2476,In_2339);
and U3186 (N_3186,In_145,In_1390);
nand U3187 (N_3187,In_1416,In_359);
nand U3188 (N_3188,In_2411,In_350);
xnor U3189 (N_3189,In_493,In_818);
xor U3190 (N_3190,In_400,In_1452);
and U3191 (N_3191,In_179,In_1720);
nand U3192 (N_3192,In_962,In_851);
or U3193 (N_3193,In_1094,In_1620);
nand U3194 (N_3194,In_1069,In_965);
or U3195 (N_3195,In_664,In_1489);
nand U3196 (N_3196,In_1899,In_1723);
xnor U3197 (N_3197,In_1892,In_1206);
nor U3198 (N_3198,In_772,In_1829);
nor U3199 (N_3199,In_435,In_918);
or U3200 (N_3200,In_315,In_1118);
nor U3201 (N_3201,In_1318,In_2153);
and U3202 (N_3202,In_444,In_558);
nor U3203 (N_3203,In_1756,In_1282);
and U3204 (N_3204,In_1117,In_1621);
nand U3205 (N_3205,In_1230,In_1910);
nor U3206 (N_3206,In_963,In_2184);
nor U3207 (N_3207,In_410,In_2477);
and U3208 (N_3208,In_1322,In_335);
or U3209 (N_3209,In_1597,In_2236);
xor U3210 (N_3210,In_408,In_1820);
nor U3211 (N_3211,In_169,In_1956);
or U3212 (N_3212,In_90,In_2148);
xor U3213 (N_3213,In_2282,In_783);
nor U3214 (N_3214,In_1929,In_2019);
and U3215 (N_3215,In_2162,In_1342);
nor U3216 (N_3216,In_320,In_842);
nand U3217 (N_3217,In_144,In_909);
nor U3218 (N_3218,In_163,In_801);
or U3219 (N_3219,In_1183,In_2239);
or U3220 (N_3220,In_820,In_440);
and U3221 (N_3221,In_693,In_2184);
nand U3222 (N_3222,In_495,In_908);
or U3223 (N_3223,In_1689,In_611);
or U3224 (N_3224,In_495,In_1860);
nand U3225 (N_3225,In_2352,In_2488);
nor U3226 (N_3226,In_415,In_1678);
nand U3227 (N_3227,In_300,In_1121);
or U3228 (N_3228,In_176,In_2169);
or U3229 (N_3229,In_47,In_2463);
nor U3230 (N_3230,In_2174,In_298);
and U3231 (N_3231,In_303,In_1397);
nand U3232 (N_3232,In_315,In_2262);
xor U3233 (N_3233,In_397,In_709);
or U3234 (N_3234,In_1579,In_2461);
or U3235 (N_3235,In_136,In_821);
or U3236 (N_3236,In_299,In_2327);
or U3237 (N_3237,In_1756,In_42);
xor U3238 (N_3238,In_443,In_2212);
or U3239 (N_3239,In_1339,In_108);
nor U3240 (N_3240,In_430,In_390);
or U3241 (N_3241,In_2493,In_865);
or U3242 (N_3242,In_2456,In_2347);
nor U3243 (N_3243,In_891,In_2293);
and U3244 (N_3244,In_389,In_1197);
xnor U3245 (N_3245,In_1349,In_1947);
nand U3246 (N_3246,In_1816,In_1035);
nor U3247 (N_3247,In_2419,In_1777);
nand U3248 (N_3248,In_93,In_341);
nor U3249 (N_3249,In_2363,In_1858);
xor U3250 (N_3250,In_2097,In_498);
or U3251 (N_3251,In_1056,In_453);
nor U3252 (N_3252,In_1629,In_1553);
nand U3253 (N_3253,In_1080,In_373);
or U3254 (N_3254,In_2154,In_339);
xnor U3255 (N_3255,In_103,In_390);
and U3256 (N_3256,In_1772,In_638);
and U3257 (N_3257,In_1832,In_2328);
xor U3258 (N_3258,In_1166,In_1171);
nor U3259 (N_3259,In_470,In_469);
nor U3260 (N_3260,In_32,In_1580);
or U3261 (N_3261,In_2473,In_1695);
xor U3262 (N_3262,In_2463,In_1434);
or U3263 (N_3263,In_1666,In_2196);
nor U3264 (N_3264,In_2026,In_244);
or U3265 (N_3265,In_455,In_76);
or U3266 (N_3266,In_1701,In_1743);
xnor U3267 (N_3267,In_709,In_1328);
xor U3268 (N_3268,In_1314,In_862);
or U3269 (N_3269,In_1970,In_866);
nor U3270 (N_3270,In_282,In_865);
nand U3271 (N_3271,In_2199,In_1471);
xnor U3272 (N_3272,In_328,In_601);
or U3273 (N_3273,In_1379,In_1710);
nand U3274 (N_3274,In_1854,In_1401);
or U3275 (N_3275,In_326,In_628);
nand U3276 (N_3276,In_2478,In_452);
nor U3277 (N_3277,In_1753,In_1217);
or U3278 (N_3278,In_1895,In_1270);
or U3279 (N_3279,In_464,In_887);
or U3280 (N_3280,In_1465,In_115);
nor U3281 (N_3281,In_2400,In_2391);
and U3282 (N_3282,In_1033,In_800);
nor U3283 (N_3283,In_1884,In_596);
nand U3284 (N_3284,In_273,In_1314);
or U3285 (N_3285,In_877,In_1975);
or U3286 (N_3286,In_995,In_988);
and U3287 (N_3287,In_1681,In_1510);
nor U3288 (N_3288,In_909,In_665);
nor U3289 (N_3289,In_645,In_261);
xor U3290 (N_3290,In_980,In_362);
and U3291 (N_3291,In_297,In_539);
xor U3292 (N_3292,In_1915,In_90);
nor U3293 (N_3293,In_2289,In_2447);
or U3294 (N_3294,In_730,In_479);
xor U3295 (N_3295,In_341,In_322);
or U3296 (N_3296,In_108,In_2487);
nand U3297 (N_3297,In_2272,In_1198);
nand U3298 (N_3298,In_538,In_1466);
xnor U3299 (N_3299,In_1625,In_1787);
nand U3300 (N_3300,In_946,In_313);
nor U3301 (N_3301,In_2427,In_132);
nand U3302 (N_3302,In_1604,In_2040);
nand U3303 (N_3303,In_1808,In_1448);
nor U3304 (N_3304,In_984,In_2156);
xnor U3305 (N_3305,In_2172,In_228);
nand U3306 (N_3306,In_1001,In_710);
xor U3307 (N_3307,In_2302,In_644);
nor U3308 (N_3308,In_261,In_392);
nand U3309 (N_3309,In_988,In_1657);
or U3310 (N_3310,In_101,In_1394);
or U3311 (N_3311,In_2388,In_2437);
xor U3312 (N_3312,In_2299,In_1689);
and U3313 (N_3313,In_1360,In_813);
xor U3314 (N_3314,In_1624,In_1764);
xnor U3315 (N_3315,In_1322,In_1203);
nor U3316 (N_3316,In_2052,In_1583);
and U3317 (N_3317,In_817,In_415);
or U3318 (N_3318,In_2342,In_142);
xnor U3319 (N_3319,In_746,In_172);
nand U3320 (N_3320,In_379,In_2081);
nor U3321 (N_3321,In_2248,In_823);
nor U3322 (N_3322,In_2419,In_51);
or U3323 (N_3323,In_166,In_76);
or U3324 (N_3324,In_1673,In_271);
xor U3325 (N_3325,In_1548,In_1935);
nor U3326 (N_3326,In_517,In_1776);
xnor U3327 (N_3327,In_1239,In_994);
and U3328 (N_3328,In_2481,In_881);
xor U3329 (N_3329,In_1961,In_653);
nor U3330 (N_3330,In_337,In_759);
and U3331 (N_3331,In_858,In_2112);
xnor U3332 (N_3332,In_293,In_1977);
or U3333 (N_3333,In_2447,In_1492);
or U3334 (N_3334,In_1595,In_994);
xnor U3335 (N_3335,In_1341,In_2246);
nor U3336 (N_3336,In_72,In_1717);
or U3337 (N_3337,In_1667,In_2136);
or U3338 (N_3338,In_617,In_773);
nor U3339 (N_3339,In_626,In_1896);
xor U3340 (N_3340,In_652,In_643);
nand U3341 (N_3341,In_1507,In_1972);
nor U3342 (N_3342,In_246,In_2190);
and U3343 (N_3343,In_2284,In_1439);
and U3344 (N_3344,In_2043,In_2123);
xor U3345 (N_3345,In_1353,In_230);
and U3346 (N_3346,In_2329,In_1132);
or U3347 (N_3347,In_1706,In_1478);
xnor U3348 (N_3348,In_1614,In_148);
nand U3349 (N_3349,In_973,In_790);
xor U3350 (N_3350,In_41,In_1416);
or U3351 (N_3351,In_801,In_1399);
or U3352 (N_3352,In_2424,In_720);
nor U3353 (N_3353,In_1997,In_843);
and U3354 (N_3354,In_2232,In_576);
or U3355 (N_3355,In_124,In_1517);
xor U3356 (N_3356,In_1595,In_1559);
xnor U3357 (N_3357,In_535,In_1703);
and U3358 (N_3358,In_437,In_2321);
xnor U3359 (N_3359,In_159,In_412);
nor U3360 (N_3360,In_624,In_319);
and U3361 (N_3361,In_762,In_1783);
and U3362 (N_3362,In_1716,In_2152);
nor U3363 (N_3363,In_1963,In_1699);
nand U3364 (N_3364,In_2197,In_1911);
nand U3365 (N_3365,In_511,In_1361);
nor U3366 (N_3366,In_952,In_2383);
or U3367 (N_3367,In_1499,In_374);
or U3368 (N_3368,In_1200,In_1685);
xor U3369 (N_3369,In_1830,In_367);
and U3370 (N_3370,In_586,In_263);
xnor U3371 (N_3371,In_1044,In_2290);
nand U3372 (N_3372,In_2498,In_931);
nand U3373 (N_3373,In_938,In_1042);
nor U3374 (N_3374,In_268,In_443);
and U3375 (N_3375,In_339,In_668);
xnor U3376 (N_3376,In_366,In_833);
or U3377 (N_3377,In_693,In_2253);
xnor U3378 (N_3378,In_1286,In_1252);
xnor U3379 (N_3379,In_255,In_1871);
and U3380 (N_3380,In_450,In_668);
xnor U3381 (N_3381,In_197,In_1471);
nand U3382 (N_3382,In_34,In_761);
nand U3383 (N_3383,In_1550,In_577);
and U3384 (N_3384,In_1977,In_417);
nor U3385 (N_3385,In_611,In_1160);
xnor U3386 (N_3386,In_1731,In_344);
and U3387 (N_3387,In_135,In_2258);
or U3388 (N_3388,In_1984,In_2342);
nor U3389 (N_3389,In_1736,In_989);
xor U3390 (N_3390,In_1665,In_733);
nor U3391 (N_3391,In_1616,In_2277);
nand U3392 (N_3392,In_27,In_1668);
and U3393 (N_3393,In_2303,In_1339);
and U3394 (N_3394,In_396,In_1963);
nor U3395 (N_3395,In_1462,In_537);
and U3396 (N_3396,In_767,In_1780);
xnor U3397 (N_3397,In_309,In_2014);
xnor U3398 (N_3398,In_894,In_1770);
nor U3399 (N_3399,In_696,In_1199);
and U3400 (N_3400,In_1488,In_1535);
and U3401 (N_3401,In_699,In_489);
nand U3402 (N_3402,In_345,In_412);
and U3403 (N_3403,In_0,In_1222);
or U3404 (N_3404,In_2279,In_1134);
xor U3405 (N_3405,In_728,In_2027);
xnor U3406 (N_3406,In_477,In_807);
and U3407 (N_3407,In_2382,In_712);
and U3408 (N_3408,In_155,In_1071);
nor U3409 (N_3409,In_165,In_1395);
xor U3410 (N_3410,In_564,In_1183);
or U3411 (N_3411,In_1870,In_1439);
nand U3412 (N_3412,In_73,In_1533);
nand U3413 (N_3413,In_1916,In_560);
nor U3414 (N_3414,In_1671,In_1724);
or U3415 (N_3415,In_1245,In_744);
nand U3416 (N_3416,In_1704,In_2202);
nor U3417 (N_3417,In_777,In_4);
nand U3418 (N_3418,In_2006,In_421);
and U3419 (N_3419,In_492,In_1756);
xnor U3420 (N_3420,In_237,In_2021);
or U3421 (N_3421,In_322,In_1037);
xnor U3422 (N_3422,In_1545,In_1838);
nor U3423 (N_3423,In_1111,In_1605);
nor U3424 (N_3424,In_437,In_1371);
nor U3425 (N_3425,In_1888,In_1532);
xnor U3426 (N_3426,In_1675,In_889);
and U3427 (N_3427,In_2493,In_555);
nand U3428 (N_3428,In_1524,In_426);
nor U3429 (N_3429,In_511,In_590);
nand U3430 (N_3430,In_2010,In_2166);
and U3431 (N_3431,In_869,In_1148);
or U3432 (N_3432,In_1880,In_968);
xor U3433 (N_3433,In_1587,In_742);
or U3434 (N_3434,In_1250,In_512);
xnor U3435 (N_3435,In_2175,In_2271);
xnor U3436 (N_3436,In_548,In_1902);
xor U3437 (N_3437,In_1551,In_1610);
nand U3438 (N_3438,In_2161,In_1810);
and U3439 (N_3439,In_918,In_2159);
and U3440 (N_3440,In_1909,In_1933);
and U3441 (N_3441,In_1414,In_2415);
xor U3442 (N_3442,In_441,In_1567);
nand U3443 (N_3443,In_931,In_799);
nor U3444 (N_3444,In_652,In_367);
xor U3445 (N_3445,In_1917,In_1209);
and U3446 (N_3446,In_768,In_742);
xnor U3447 (N_3447,In_872,In_1275);
or U3448 (N_3448,In_1747,In_2224);
nand U3449 (N_3449,In_131,In_810);
xor U3450 (N_3450,In_781,In_2225);
xor U3451 (N_3451,In_1933,In_642);
nand U3452 (N_3452,In_1323,In_1516);
xnor U3453 (N_3453,In_2048,In_1151);
and U3454 (N_3454,In_2345,In_1975);
or U3455 (N_3455,In_1791,In_358);
xor U3456 (N_3456,In_1397,In_2100);
nand U3457 (N_3457,In_1476,In_1756);
or U3458 (N_3458,In_1707,In_1006);
nand U3459 (N_3459,In_1575,In_1132);
or U3460 (N_3460,In_264,In_1598);
or U3461 (N_3461,In_2139,In_802);
nand U3462 (N_3462,In_563,In_2058);
or U3463 (N_3463,In_2466,In_939);
or U3464 (N_3464,In_1092,In_520);
or U3465 (N_3465,In_1101,In_1873);
nor U3466 (N_3466,In_724,In_1411);
nor U3467 (N_3467,In_426,In_1946);
nand U3468 (N_3468,In_760,In_549);
nor U3469 (N_3469,In_1161,In_1393);
xnor U3470 (N_3470,In_1148,In_1089);
and U3471 (N_3471,In_1323,In_678);
nand U3472 (N_3472,In_24,In_1381);
xnor U3473 (N_3473,In_1771,In_869);
nand U3474 (N_3474,In_1192,In_1093);
xnor U3475 (N_3475,In_1987,In_1528);
or U3476 (N_3476,In_312,In_2046);
nor U3477 (N_3477,In_1469,In_1715);
nand U3478 (N_3478,In_225,In_1719);
nand U3479 (N_3479,In_933,In_482);
and U3480 (N_3480,In_246,In_1957);
xnor U3481 (N_3481,In_140,In_2297);
and U3482 (N_3482,In_480,In_2233);
or U3483 (N_3483,In_1650,In_1067);
or U3484 (N_3484,In_2346,In_432);
nor U3485 (N_3485,In_85,In_791);
nor U3486 (N_3486,In_1101,In_427);
xor U3487 (N_3487,In_495,In_2454);
xnor U3488 (N_3488,In_2347,In_1347);
nand U3489 (N_3489,In_1522,In_264);
nand U3490 (N_3490,In_1129,In_2254);
xnor U3491 (N_3491,In_1661,In_434);
nand U3492 (N_3492,In_2497,In_577);
xnor U3493 (N_3493,In_1268,In_974);
nor U3494 (N_3494,In_312,In_387);
nand U3495 (N_3495,In_672,In_1644);
xor U3496 (N_3496,In_1974,In_1221);
nor U3497 (N_3497,In_207,In_868);
nand U3498 (N_3498,In_25,In_1848);
and U3499 (N_3499,In_1756,In_157);
xor U3500 (N_3500,In_2363,In_474);
xor U3501 (N_3501,In_551,In_1846);
nor U3502 (N_3502,In_86,In_1337);
nor U3503 (N_3503,In_1158,In_542);
nor U3504 (N_3504,In_961,In_2360);
and U3505 (N_3505,In_1551,In_1111);
nand U3506 (N_3506,In_381,In_560);
nor U3507 (N_3507,In_1686,In_358);
nand U3508 (N_3508,In_861,In_730);
or U3509 (N_3509,In_760,In_2269);
nor U3510 (N_3510,In_630,In_2435);
or U3511 (N_3511,In_2031,In_150);
or U3512 (N_3512,In_2320,In_486);
and U3513 (N_3513,In_360,In_209);
nor U3514 (N_3514,In_1235,In_1401);
nor U3515 (N_3515,In_231,In_1838);
and U3516 (N_3516,In_233,In_2147);
or U3517 (N_3517,In_573,In_2080);
or U3518 (N_3518,In_1479,In_1334);
and U3519 (N_3519,In_1184,In_2209);
nor U3520 (N_3520,In_766,In_522);
nand U3521 (N_3521,In_925,In_2181);
or U3522 (N_3522,In_2113,In_1184);
and U3523 (N_3523,In_1479,In_328);
and U3524 (N_3524,In_861,In_85);
and U3525 (N_3525,In_744,In_2438);
nand U3526 (N_3526,In_875,In_706);
or U3527 (N_3527,In_417,In_1214);
or U3528 (N_3528,In_321,In_1205);
or U3529 (N_3529,In_2383,In_2259);
and U3530 (N_3530,In_450,In_156);
xor U3531 (N_3531,In_2204,In_2245);
nand U3532 (N_3532,In_2116,In_37);
and U3533 (N_3533,In_2172,In_2061);
or U3534 (N_3534,In_2184,In_1567);
nand U3535 (N_3535,In_371,In_548);
nand U3536 (N_3536,In_2046,In_2129);
nand U3537 (N_3537,In_2049,In_999);
or U3538 (N_3538,In_988,In_879);
nor U3539 (N_3539,In_295,In_1108);
and U3540 (N_3540,In_2345,In_1340);
xor U3541 (N_3541,In_1277,In_2297);
and U3542 (N_3542,In_631,In_2088);
and U3543 (N_3543,In_2194,In_1481);
nand U3544 (N_3544,In_1537,In_1540);
or U3545 (N_3545,In_1485,In_243);
nand U3546 (N_3546,In_1799,In_1198);
xor U3547 (N_3547,In_1269,In_271);
nor U3548 (N_3548,In_1953,In_373);
or U3549 (N_3549,In_1392,In_1119);
nor U3550 (N_3550,In_1302,In_2400);
nor U3551 (N_3551,In_1971,In_630);
nor U3552 (N_3552,In_529,In_649);
and U3553 (N_3553,In_1912,In_2144);
nand U3554 (N_3554,In_1960,In_1675);
xor U3555 (N_3555,In_1171,In_824);
xor U3556 (N_3556,In_630,In_750);
nand U3557 (N_3557,In_820,In_898);
and U3558 (N_3558,In_1858,In_822);
xnor U3559 (N_3559,In_2323,In_975);
or U3560 (N_3560,In_2369,In_2457);
xor U3561 (N_3561,In_2369,In_1161);
or U3562 (N_3562,In_940,In_1824);
nor U3563 (N_3563,In_1872,In_1151);
xnor U3564 (N_3564,In_288,In_534);
nand U3565 (N_3565,In_2369,In_553);
nand U3566 (N_3566,In_684,In_1415);
nor U3567 (N_3567,In_1431,In_628);
and U3568 (N_3568,In_1606,In_1462);
nand U3569 (N_3569,In_961,In_2353);
xnor U3570 (N_3570,In_1972,In_513);
and U3571 (N_3571,In_170,In_1240);
nor U3572 (N_3572,In_1642,In_503);
nand U3573 (N_3573,In_799,In_1371);
nor U3574 (N_3574,In_15,In_855);
and U3575 (N_3575,In_2465,In_926);
nand U3576 (N_3576,In_1688,In_240);
nor U3577 (N_3577,In_368,In_316);
nand U3578 (N_3578,In_2444,In_223);
or U3579 (N_3579,In_1565,In_999);
and U3580 (N_3580,In_1728,In_1677);
and U3581 (N_3581,In_484,In_2361);
nand U3582 (N_3582,In_160,In_1252);
xor U3583 (N_3583,In_2300,In_779);
xor U3584 (N_3584,In_267,In_1081);
and U3585 (N_3585,In_667,In_103);
nand U3586 (N_3586,In_2354,In_1442);
xnor U3587 (N_3587,In_1266,In_2098);
xor U3588 (N_3588,In_1226,In_1705);
and U3589 (N_3589,In_763,In_2260);
xor U3590 (N_3590,In_116,In_939);
or U3591 (N_3591,In_1645,In_1565);
nor U3592 (N_3592,In_2361,In_1650);
and U3593 (N_3593,In_957,In_1571);
nand U3594 (N_3594,In_1287,In_2053);
and U3595 (N_3595,In_2224,In_1761);
xor U3596 (N_3596,In_1816,In_1440);
xor U3597 (N_3597,In_1418,In_925);
nor U3598 (N_3598,In_863,In_1428);
nand U3599 (N_3599,In_726,In_1487);
xor U3600 (N_3600,In_272,In_2296);
nor U3601 (N_3601,In_1209,In_1222);
nand U3602 (N_3602,In_902,In_1257);
nor U3603 (N_3603,In_307,In_2022);
nor U3604 (N_3604,In_200,In_1755);
and U3605 (N_3605,In_2268,In_15);
and U3606 (N_3606,In_1341,In_480);
nor U3607 (N_3607,In_424,In_98);
nand U3608 (N_3608,In_428,In_1426);
nor U3609 (N_3609,In_590,In_1322);
and U3610 (N_3610,In_2206,In_374);
xor U3611 (N_3611,In_818,In_2115);
nand U3612 (N_3612,In_539,In_2492);
nor U3613 (N_3613,In_1104,In_1681);
nor U3614 (N_3614,In_305,In_627);
nor U3615 (N_3615,In_2324,In_597);
or U3616 (N_3616,In_894,In_642);
nand U3617 (N_3617,In_2485,In_1012);
or U3618 (N_3618,In_898,In_772);
or U3619 (N_3619,In_552,In_1838);
nand U3620 (N_3620,In_2322,In_721);
nor U3621 (N_3621,In_786,In_1371);
nand U3622 (N_3622,In_539,In_1089);
and U3623 (N_3623,In_1855,In_915);
xnor U3624 (N_3624,In_1380,In_1947);
nor U3625 (N_3625,In_1769,In_310);
and U3626 (N_3626,In_169,In_1221);
or U3627 (N_3627,In_1882,In_346);
nor U3628 (N_3628,In_1693,In_423);
and U3629 (N_3629,In_2261,In_928);
or U3630 (N_3630,In_2114,In_1388);
nor U3631 (N_3631,In_2004,In_1512);
nand U3632 (N_3632,In_2056,In_1554);
or U3633 (N_3633,In_1046,In_2057);
nand U3634 (N_3634,In_1013,In_876);
and U3635 (N_3635,In_1383,In_363);
and U3636 (N_3636,In_659,In_2255);
nand U3637 (N_3637,In_245,In_1962);
or U3638 (N_3638,In_1631,In_632);
or U3639 (N_3639,In_66,In_1513);
and U3640 (N_3640,In_354,In_1438);
nor U3641 (N_3641,In_1012,In_27);
or U3642 (N_3642,In_779,In_822);
and U3643 (N_3643,In_2261,In_2219);
and U3644 (N_3644,In_1816,In_229);
and U3645 (N_3645,In_2097,In_180);
and U3646 (N_3646,In_69,In_184);
xnor U3647 (N_3647,In_1290,In_891);
nor U3648 (N_3648,In_1298,In_1453);
nand U3649 (N_3649,In_6,In_1655);
or U3650 (N_3650,In_2131,In_420);
nor U3651 (N_3651,In_754,In_226);
nor U3652 (N_3652,In_125,In_599);
nor U3653 (N_3653,In_44,In_1543);
or U3654 (N_3654,In_1988,In_1300);
or U3655 (N_3655,In_1407,In_753);
nand U3656 (N_3656,In_1269,In_727);
nand U3657 (N_3657,In_2237,In_1176);
and U3658 (N_3658,In_379,In_32);
nand U3659 (N_3659,In_1932,In_2406);
and U3660 (N_3660,In_1691,In_2149);
xor U3661 (N_3661,In_1640,In_96);
or U3662 (N_3662,In_1540,In_1882);
nor U3663 (N_3663,In_2192,In_820);
nor U3664 (N_3664,In_1934,In_2324);
and U3665 (N_3665,In_1179,In_1351);
or U3666 (N_3666,In_1357,In_2314);
or U3667 (N_3667,In_1658,In_710);
xnor U3668 (N_3668,In_483,In_1807);
xor U3669 (N_3669,In_675,In_500);
xnor U3670 (N_3670,In_313,In_819);
or U3671 (N_3671,In_1866,In_1242);
nand U3672 (N_3672,In_2096,In_1395);
or U3673 (N_3673,In_877,In_999);
and U3674 (N_3674,In_1995,In_603);
nand U3675 (N_3675,In_603,In_822);
and U3676 (N_3676,In_1567,In_1229);
nand U3677 (N_3677,In_1875,In_322);
xnor U3678 (N_3678,In_532,In_1657);
nand U3679 (N_3679,In_1719,In_1455);
nor U3680 (N_3680,In_394,In_743);
nor U3681 (N_3681,In_1052,In_1297);
xor U3682 (N_3682,In_2194,In_1911);
nand U3683 (N_3683,In_2273,In_229);
and U3684 (N_3684,In_942,In_2264);
nand U3685 (N_3685,In_126,In_148);
and U3686 (N_3686,In_1044,In_2010);
nor U3687 (N_3687,In_1813,In_1658);
and U3688 (N_3688,In_1998,In_1461);
or U3689 (N_3689,In_1609,In_194);
or U3690 (N_3690,In_1574,In_1698);
and U3691 (N_3691,In_740,In_1301);
xor U3692 (N_3692,In_1333,In_1600);
and U3693 (N_3693,In_1529,In_674);
xor U3694 (N_3694,In_1298,In_944);
and U3695 (N_3695,In_1609,In_558);
and U3696 (N_3696,In_1123,In_2402);
xor U3697 (N_3697,In_2422,In_2063);
nand U3698 (N_3698,In_62,In_786);
nand U3699 (N_3699,In_1732,In_32);
or U3700 (N_3700,In_664,In_338);
nor U3701 (N_3701,In_145,In_233);
nor U3702 (N_3702,In_285,In_1209);
nor U3703 (N_3703,In_576,In_1721);
nor U3704 (N_3704,In_1566,In_1216);
or U3705 (N_3705,In_1741,In_110);
xnor U3706 (N_3706,In_71,In_860);
xor U3707 (N_3707,In_117,In_1172);
xor U3708 (N_3708,In_1957,In_257);
nor U3709 (N_3709,In_849,In_1659);
and U3710 (N_3710,In_923,In_494);
and U3711 (N_3711,In_1482,In_635);
nand U3712 (N_3712,In_2154,In_2404);
nand U3713 (N_3713,In_999,In_2193);
nor U3714 (N_3714,In_1524,In_415);
xor U3715 (N_3715,In_374,In_1822);
xnor U3716 (N_3716,In_1440,In_2213);
xnor U3717 (N_3717,In_1238,In_720);
nor U3718 (N_3718,In_142,In_1586);
or U3719 (N_3719,In_1253,In_1273);
or U3720 (N_3720,In_221,In_678);
xor U3721 (N_3721,In_1190,In_896);
and U3722 (N_3722,In_942,In_1222);
and U3723 (N_3723,In_320,In_936);
and U3724 (N_3724,In_935,In_972);
or U3725 (N_3725,In_149,In_50);
nand U3726 (N_3726,In_1011,In_251);
nand U3727 (N_3727,In_2280,In_1095);
or U3728 (N_3728,In_1621,In_1832);
nand U3729 (N_3729,In_612,In_2217);
and U3730 (N_3730,In_1768,In_1508);
or U3731 (N_3731,In_1498,In_2311);
nor U3732 (N_3732,In_15,In_1627);
xnor U3733 (N_3733,In_997,In_953);
nand U3734 (N_3734,In_2142,In_687);
and U3735 (N_3735,In_1189,In_1346);
and U3736 (N_3736,In_2293,In_872);
or U3737 (N_3737,In_2345,In_2228);
nor U3738 (N_3738,In_2020,In_816);
nor U3739 (N_3739,In_2273,In_1654);
nand U3740 (N_3740,In_1379,In_1132);
or U3741 (N_3741,In_1185,In_1651);
xor U3742 (N_3742,In_1020,In_2370);
nand U3743 (N_3743,In_1429,In_1053);
nand U3744 (N_3744,In_1191,In_655);
nor U3745 (N_3745,In_135,In_2210);
nor U3746 (N_3746,In_1214,In_2007);
xnor U3747 (N_3747,In_1502,In_2032);
and U3748 (N_3748,In_2020,In_1947);
nor U3749 (N_3749,In_1572,In_2101);
or U3750 (N_3750,In_1691,In_144);
nand U3751 (N_3751,In_689,In_1995);
nor U3752 (N_3752,In_1149,In_2107);
xor U3753 (N_3753,In_1190,In_1154);
nor U3754 (N_3754,In_1308,In_1858);
or U3755 (N_3755,In_822,In_578);
nand U3756 (N_3756,In_1282,In_1760);
nand U3757 (N_3757,In_1303,In_422);
or U3758 (N_3758,In_177,In_2222);
and U3759 (N_3759,In_100,In_665);
xor U3760 (N_3760,In_905,In_686);
xor U3761 (N_3761,In_1097,In_1405);
nor U3762 (N_3762,In_1590,In_473);
and U3763 (N_3763,In_1985,In_1605);
xor U3764 (N_3764,In_649,In_966);
and U3765 (N_3765,In_784,In_1602);
nor U3766 (N_3766,In_1495,In_88);
or U3767 (N_3767,In_1868,In_1558);
and U3768 (N_3768,In_1520,In_1220);
or U3769 (N_3769,In_641,In_45);
nor U3770 (N_3770,In_1924,In_998);
xor U3771 (N_3771,In_2389,In_1175);
or U3772 (N_3772,In_121,In_859);
nor U3773 (N_3773,In_1134,In_1445);
or U3774 (N_3774,In_128,In_1178);
nand U3775 (N_3775,In_2380,In_2449);
or U3776 (N_3776,In_1548,In_1176);
xnor U3777 (N_3777,In_2175,In_223);
or U3778 (N_3778,In_1880,In_2202);
and U3779 (N_3779,In_953,In_2294);
nor U3780 (N_3780,In_1309,In_1856);
nand U3781 (N_3781,In_1668,In_2497);
nand U3782 (N_3782,In_1813,In_45);
nor U3783 (N_3783,In_1173,In_2108);
nand U3784 (N_3784,In_1801,In_457);
nor U3785 (N_3785,In_942,In_1293);
xnor U3786 (N_3786,In_1467,In_1934);
nor U3787 (N_3787,In_1539,In_2114);
and U3788 (N_3788,In_1557,In_2496);
nor U3789 (N_3789,In_272,In_1441);
xnor U3790 (N_3790,In_2434,In_1781);
or U3791 (N_3791,In_714,In_526);
or U3792 (N_3792,In_1359,In_125);
and U3793 (N_3793,In_1803,In_2264);
and U3794 (N_3794,In_1618,In_867);
nand U3795 (N_3795,In_2285,In_284);
and U3796 (N_3796,In_87,In_1450);
xnor U3797 (N_3797,In_1235,In_1422);
and U3798 (N_3798,In_1753,In_1512);
xor U3799 (N_3799,In_934,In_1931);
and U3800 (N_3800,In_59,In_2216);
and U3801 (N_3801,In_1950,In_1909);
xor U3802 (N_3802,In_360,In_359);
nand U3803 (N_3803,In_1588,In_1152);
xor U3804 (N_3804,In_2377,In_1131);
nand U3805 (N_3805,In_131,In_1535);
xor U3806 (N_3806,In_1346,In_182);
and U3807 (N_3807,In_81,In_1782);
nand U3808 (N_3808,In_2324,In_1019);
nor U3809 (N_3809,In_419,In_1359);
nand U3810 (N_3810,In_2043,In_1849);
nand U3811 (N_3811,In_1437,In_1161);
xnor U3812 (N_3812,In_102,In_250);
or U3813 (N_3813,In_662,In_1273);
and U3814 (N_3814,In_977,In_182);
and U3815 (N_3815,In_2216,In_252);
and U3816 (N_3816,In_2354,In_1275);
xor U3817 (N_3817,In_1709,In_1538);
nor U3818 (N_3818,In_1490,In_276);
nand U3819 (N_3819,In_1113,In_206);
nand U3820 (N_3820,In_2259,In_463);
xnor U3821 (N_3821,In_2487,In_1530);
nor U3822 (N_3822,In_306,In_2251);
and U3823 (N_3823,In_644,In_1563);
xnor U3824 (N_3824,In_2383,In_827);
nor U3825 (N_3825,In_973,In_278);
nor U3826 (N_3826,In_391,In_1221);
nor U3827 (N_3827,In_581,In_905);
or U3828 (N_3828,In_240,In_1971);
or U3829 (N_3829,In_1845,In_378);
nand U3830 (N_3830,In_1237,In_1249);
or U3831 (N_3831,In_1406,In_272);
nor U3832 (N_3832,In_1492,In_2060);
or U3833 (N_3833,In_1616,In_139);
xnor U3834 (N_3834,In_2199,In_1267);
and U3835 (N_3835,In_1458,In_1949);
xnor U3836 (N_3836,In_512,In_1821);
nand U3837 (N_3837,In_2224,In_272);
nand U3838 (N_3838,In_1014,In_1905);
or U3839 (N_3839,In_2350,In_653);
nor U3840 (N_3840,In_287,In_2183);
nand U3841 (N_3841,In_2282,In_179);
and U3842 (N_3842,In_215,In_1623);
nand U3843 (N_3843,In_1972,In_2464);
xor U3844 (N_3844,In_688,In_2090);
xnor U3845 (N_3845,In_1611,In_2473);
nand U3846 (N_3846,In_1666,In_1993);
nand U3847 (N_3847,In_1199,In_2140);
or U3848 (N_3848,In_501,In_1253);
nor U3849 (N_3849,In_2162,In_509);
xnor U3850 (N_3850,In_2111,In_2345);
nand U3851 (N_3851,In_211,In_614);
nand U3852 (N_3852,In_792,In_258);
xnor U3853 (N_3853,In_1814,In_1505);
and U3854 (N_3854,In_327,In_2263);
or U3855 (N_3855,In_996,In_2245);
nor U3856 (N_3856,In_1100,In_1673);
nand U3857 (N_3857,In_1521,In_2080);
nor U3858 (N_3858,In_347,In_111);
and U3859 (N_3859,In_2492,In_1585);
or U3860 (N_3860,In_910,In_949);
nand U3861 (N_3861,In_780,In_1470);
and U3862 (N_3862,In_434,In_1197);
xnor U3863 (N_3863,In_328,In_2028);
and U3864 (N_3864,In_10,In_1938);
nand U3865 (N_3865,In_121,In_2110);
or U3866 (N_3866,In_334,In_803);
xnor U3867 (N_3867,In_1542,In_65);
or U3868 (N_3868,In_1151,In_190);
or U3869 (N_3869,In_964,In_1514);
and U3870 (N_3870,In_2312,In_1970);
xor U3871 (N_3871,In_623,In_545);
and U3872 (N_3872,In_2024,In_1674);
xnor U3873 (N_3873,In_558,In_1151);
or U3874 (N_3874,In_618,In_189);
nand U3875 (N_3875,In_163,In_62);
nor U3876 (N_3876,In_2071,In_964);
and U3877 (N_3877,In_2160,In_2157);
nor U3878 (N_3878,In_2476,In_293);
xor U3879 (N_3879,In_1626,In_2402);
nand U3880 (N_3880,In_245,In_681);
or U3881 (N_3881,In_271,In_1873);
and U3882 (N_3882,In_631,In_664);
xor U3883 (N_3883,In_2030,In_1308);
nand U3884 (N_3884,In_528,In_2166);
xnor U3885 (N_3885,In_955,In_2041);
or U3886 (N_3886,In_562,In_1729);
or U3887 (N_3887,In_1229,In_1885);
or U3888 (N_3888,In_41,In_79);
xnor U3889 (N_3889,In_1579,In_640);
and U3890 (N_3890,In_1322,In_555);
and U3891 (N_3891,In_1203,In_1847);
nand U3892 (N_3892,In_435,In_2345);
xnor U3893 (N_3893,In_948,In_207);
or U3894 (N_3894,In_724,In_495);
xor U3895 (N_3895,In_2025,In_1925);
or U3896 (N_3896,In_930,In_971);
xor U3897 (N_3897,In_1146,In_2195);
or U3898 (N_3898,In_363,In_457);
xnor U3899 (N_3899,In_1351,In_1309);
nand U3900 (N_3900,In_1717,In_24);
and U3901 (N_3901,In_228,In_1380);
xnor U3902 (N_3902,In_710,In_222);
nand U3903 (N_3903,In_1097,In_290);
nor U3904 (N_3904,In_2367,In_177);
nand U3905 (N_3905,In_1698,In_646);
nor U3906 (N_3906,In_492,In_1222);
nor U3907 (N_3907,In_1503,In_1018);
or U3908 (N_3908,In_1086,In_2125);
and U3909 (N_3909,In_1252,In_2427);
nand U3910 (N_3910,In_738,In_650);
nand U3911 (N_3911,In_2058,In_1583);
and U3912 (N_3912,In_1195,In_993);
and U3913 (N_3913,In_2257,In_2476);
or U3914 (N_3914,In_1438,In_1926);
or U3915 (N_3915,In_1466,In_119);
or U3916 (N_3916,In_1116,In_942);
and U3917 (N_3917,In_1570,In_508);
or U3918 (N_3918,In_1887,In_2392);
or U3919 (N_3919,In_391,In_434);
xor U3920 (N_3920,In_1359,In_154);
nand U3921 (N_3921,In_170,In_144);
nor U3922 (N_3922,In_2001,In_1233);
or U3923 (N_3923,In_32,In_2043);
and U3924 (N_3924,In_2386,In_1534);
or U3925 (N_3925,In_112,In_1596);
or U3926 (N_3926,In_58,In_1003);
nand U3927 (N_3927,In_616,In_1537);
nor U3928 (N_3928,In_2138,In_2035);
or U3929 (N_3929,In_114,In_703);
nand U3930 (N_3930,In_1299,In_806);
and U3931 (N_3931,In_1497,In_982);
nor U3932 (N_3932,In_1211,In_2388);
xor U3933 (N_3933,In_2181,In_621);
nand U3934 (N_3934,In_2279,In_405);
and U3935 (N_3935,In_911,In_599);
nor U3936 (N_3936,In_1884,In_2345);
nor U3937 (N_3937,In_1736,In_1746);
xor U3938 (N_3938,In_1314,In_1086);
xnor U3939 (N_3939,In_1371,In_2202);
or U3940 (N_3940,In_1352,In_1279);
or U3941 (N_3941,In_1464,In_1335);
xor U3942 (N_3942,In_1847,In_1722);
and U3943 (N_3943,In_499,In_1945);
and U3944 (N_3944,In_1843,In_2091);
xnor U3945 (N_3945,In_1923,In_1245);
or U3946 (N_3946,In_1741,In_1749);
or U3947 (N_3947,In_1998,In_1817);
and U3948 (N_3948,In_1631,In_2202);
xnor U3949 (N_3949,In_761,In_2466);
or U3950 (N_3950,In_244,In_1971);
xnor U3951 (N_3951,In_119,In_16);
and U3952 (N_3952,In_797,In_580);
and U3953 (N_3953,In_1370,In_944);
nor U3954 (N_3954,In_1749,In_2377);
nand U3955 (N_3955,In_2329,In_367);
nand U3956 (N_3956,In_292,In_2467);
nor U3957 (N_3957,In_889,In_1893);
nand U3958 (N_3958,In_936,In_503);
nand U3959 (N_3959,In_2333,In_1221);
xor U3960 (N_3960,In_2065,In_2304);
or U3961 (N_3961,In_529,In_314);
or U3962 (N_3962,In_840,In_1309);
nand U3963 (N_3963,In_1191,In_344);
xnor U3964 (N_3964,In_1251,In_453);
nor U3965 (N_3965,In_1231,In_1904);
xnor U3966 (N_3966,In_1167,In_1520);
or U3967 (N_3967,In_1595,In_2116);
and U3968 (N_3968,In_372,In_841);
nor U3969 (N_3969,In_2085,In_1547);
nor U3970 (N_3970,In_2414,In_1228);
and U3971 (N_3971,In_1904,In_2088);
and U3972 (N_3972,In_1374,In_1600);
and U3973 (N_3973,In_2337,In_96);
xor U3974 (N_3974,In_273,In_1501);
xor U3975 (N_3975,In_2184,In_701);
nor U3976 (N_3976,In_1409,In_1553);
and U3977 (N_3977,In_2273,In_20);
and U3978 (N_3978,In_897,In_1122);
xor U3979 (N_3979,In_2213,In_526);
and U3980 (N_3980,In_1865,In_1614);
or U3981 (N_3981,In_98,In_2181);
xor U3982 (N_3982,In_1045,In_219);
or U3983 (N_3983,In_1718,In_1079);
nor U3984 (N_3984,In_2268,In_458);
nand U3985 (N_3985,In_1528,In_1382);
xnor U3986 (N_3986,In_2439,In_1138);
or U3987 (N_3987,In_624,In_59);
or U3988 (N_3988,In_501,In_1555);
nand U3989 (N_3989,In_2386,In_45);
and U3990 (N_3990,In_612,In_1254);
nor U3991 (N_3991,In_53,In_2046);
and U3992 (N_3992,In_1797,In_772);
nand U3993 (N_3993,In_875,In_1349);
and U3994 (N_3994,In_560,In_2159);
xnor U3995 (N_3995,In_1226,In_966);
nor U3996 (N_3996,In_2052,In_2309);
nor U3997 (N_3997,In_791,In_18);
nor U3998 (N_3998,In_930,In_2196);
xnor U3999 (N_3999,In_1479,In_2061);
nor U4000 (N_4000,In_1292,In_624);
nand U4001 (N_4001,In_1613,In_2251);
xor U4002 (N_4002,In_1320,In_971);
nand U4003 (N_4003,In_970,In_1821);
nor U4004 (N_4004,In_210,In_2442);
and U4005 (N_4005,In_1185,In_442);
or U4006 (N_4006,In_593,In_2257);
nand U4007 (N_4007,In_1547,In_355);
and U4008 (N_4008,In_1628,In_87);
and U4009 (N_4009,In_338,In_1169);
and U4010 (N_4010,In_2277,In_263);
nor U4011 (N_4011,In_2020,In_2090);
or U4012 (N_4012,In_632,In_1359);
or U4013 (N_4013,In_1029,In_1140);
or U4014 (N_4014,In_365,In_1814);
xor U4015 (N_4015,In_559,In_844);
nor U4016 (N_4016,In_2242,In_2041);
nand U4017 (N_4017,In_504,In_1396);
nand U4018 (N_4018,In_1674,In_2408);
nor U4019 (N_4019,In_1814,In_2431);
nand U4020 (N_4020,In_370,In_725);
nand U4021 (N_4021,In_1467,In_2189);
and U4022 (N_4022,In_1528,In_851);
and U4023 (N_4023,In_1557,In_1990);
xnor U4024 (N_4024,In_1549,In_755);
nor U4025 (N_4025,In_934,In_213);
nor U4026 (N_4026,In_1792,In_1892);
nand U4027 (N_4027,In_2267,In_1045);
or U4028 (N_4028,In_1149,In_2046);
nand U4029 (N_4029,In_2061,In_2484);
nor U4030 (N_4030,In_1456,In_297);
xnor U4031 (N_4031,In_55,In_550);
nor U4032 (N_4032,In_955,In_1595);
and U4033 (N_4033,In_1335,In_526);
nor U4034 (N_4034,In_1642,In_941);
and U4035 (N_4035,In_426,In_134);
and U4036 (N_4036,In_747,In_561);
or U4037 (N_4037,In_1861,In_249);
and U4038 (N_4038,In_2341,In_2283);
nor U4039 (N_4039,In_684,In_79);
nand U4040 (N_4040,In_1247,In_466);
nor U4041 (N_4041,In_1317,In_1259);
xnor U4042 (N_4042,In_2335,In_1207);
nor U4043 (N_4043,In_2453,In_1977);
nor U4044 (N_4044,In_2301,In_1082);
nand U4045 (N_4045,In_48,In_866);
nor U4046 (N_4046,In_629,In_1097);
nand U4047 (N_4047,In_1044,In_2356);
xor U4048 (N_4048,In_587,In_1182);
nand U4049 (N_4049,In_747,In_2179);
or U4050 (N_4050,In_1515,In_2480);
xnor U4051 (N_4051,In_1660,In_450);
nor U4052 (N_4052,In_1102,In_1680);
or U4053 (N_4053,In_1813,In_265);
or U4054 (N_4054,In_2045,In_631);
xor U4055 (N_4055,In_505,In_810);
nor U4056 (N_4056,In_707,In_268);
nand U4057 (N_4057,In_2082,In_801);
nand U4058 (N_4058,In_770,In_539);
or U4059 (N_4059,In_686,In_1593);
nand U4060 (N_4060,In_2129,In_2455);
nand U4061 (N_4061,In_1826,In_1198);
xor U4062 (N_4062,In_2341,In_1388);
nand U4063 (N_4063,In_2469,In_1335);
nor U4064 (N_4064,In_719,In_890);
or U4065 (N_4065,In_2221,In_884);
or U4066 (N_4066,In_1052,In_555);
nand U4067 (N_4067,In_1215,In_154);
or U4068 (N_4068,In_1407,In_1386);
and U4069 (N_4069,In_954,In_1157);
nand U4070 (N_4070,In_2183,In_1238);
or U4071 (N_4071,In_1882,In_458);
or U4072 (N_4072,In_103,In_1794);
nor U4073 (N_4073,In_1301,In_331);
nand U4074 (N_4074,In_986,In_1470);
xnor U4075 (N_4075,In_1537,In_1982);
nor U4076 (N_4076,In_1169,In_939);
xnor U4077 (N_4077,In_366,In_671);
nor U4078 (N_4078,In_1718,In_1737);
and U4079 (N_4079,In_1683,In_1655);
xnor U4080 (N_4080,In_702,In_1724);
nand U4081 (N_4081,In_1327,In_498);
nor U4082 (N_4082,In_1823,In_1452);
and U4083 (N_4083,In_1465,In_503);
nand U4084 (N_4084,In_222,In_2190);
xnor U4085 (N_4085,In_444,In_1791);
nand U4086 (N_4086,In_2137,In_988);
and U4087 (N_4087,In_194,In_358);
and U4088 (N_4088,In_1520,In_1005);
xor U4089 (N_4089,In_565,In_433);
xor U4090 (N_4090,In_161,In_1692);
and U4091 (N_4091,In_1595,In_1481);
nand U4092 (N_4092,In_589,In_1904);
or U4093 (N_4093,In_2308,In_834);
xor U4094 (N_4094,In_1345,In_1264);
or U4095 (N_4095,In_1051,In_2326);
and U4096 (N_4096,In_330,In_1843);
or U4097 (N_4097,In_227,In_737);
or U4098 (N_4098,In_148,In_356);
or U4099 (N_4099,In_2172,In_493);
xor U4100 (N_4100,In_1560,In_650);
nor U4101 (N_4101,In_2385,In_2360);
nand U4102 (N_4102,In_1085,In_2260);
and U4103 (N_4103,In_1026,In_2435);
nor U4104 (N_4104,In_516,In_1235);
or U4105 (N_4105,In_2254,In_1420);
xor U4106 (N_4106,In_2468,In_2416);
nor U4107 (N_4107,In_399,In_992);
xor U4108 (N_4108,In_1804,In_298);
or U4109 (N_4109,In_1826,In_334);
xor U4110 (N_4110,In_1034,In_100);
and U4111 (N_4111,In_164,In_7);
and U4112 (N_4112,In_2303,In_1492);
or U4113 (N_4113,In_717,In_900);
nand U4114 (N_4114,In_1448,In_5);
and U4115 (N_4115,In_2022,In_756);
and U4116 (N_4116,In_942,In_1692);
xnor U4117 (N_4117,In_152,In_805);
xor U4118 (N_4118,In_556,In_472);
or U4119 (N_4119,In_1984,In_366);
and U4120 (N_4120,In_1858,In_2017);
and U4121 (N_4121,In_2167,In_2497);
nor U4122 (N_4122,In_821,In_517);
and U4123 (N_4123,In_1049,In_421);
nor U4124 (N_4124,In_1509,In_1629);
nand U4125 (N_4125,In_1579,In_1969);
or U4126 (N_4126,In_1376,In_430);
and U4127 (N_4127,In_189,In_2130);
nor U4128 (N_4128,In_466,In_2180);
xor U4129 (N_4129,In_552,In_169);
or U4130 (N_4130,In_1469,In_2359);
xnor U4131 (N_4131,In_1608,In_1125);
or U4132 (N_4132,In_971,In_1777);
nand U4133 (N_4133,In_2144,In_1722);
or U4134 (N_4134,In_792,In_666);
and U4135 (N_4135,In_989,In_1953);
xor U4136 (N_4136,In_321,In_1183);
or U4137 (N_4137,In_2274,In_444);
and U4138 (N_4138,In_617,In_68);
or U4139 (N_4139,In_1391,In_2291);
nor U4140 (N_4140,In_2381,In_1483);
and U4141 (N_4141,In_1645,In_1649);
and U4142 (N_4142,In_86,In_945);
nor U4143 (N_4143,In_629,In_1366);
and U4144 (N_4144,In_2245,In_2270);
and U4145 (N_4145,In_1002,In_2389);
nand U4146 (N_4146,In_2189,In_1924);
xnor U4147 (N_4147,In_211,In_657);
or U4148 (N_4148,In_1764,In_1262);
or U4149 (N_4149,In_484,In_2376);
nand U4150 (N_4150,In_2469,In_1515);
or U4151 (N_4151,In_559,In_2058);
or U4152 (N_4152,In_1766,In_1853);
nand U4153 (N_4153,In_688,In_842);
xnor U4154 (N_4154,In_768,In_1633);
nor U4155 (N_4155,In_1372,In_1052);
nor U4156 (N_4156,In_131,In_2370);
and U4157 (N_4157,In_616,In_1157);
nor U4158 (N_4158,In_16,In_2286);
nand U4159 (N_4159,In_1611,In_1971);
xor U4160 (N_4160,In_302,In_2405);
xnor U4161 (N_4161,In_1547,In_1787);
nor U4162 (N_4162,In_555,In_1910);
nor U4163 (N_4163,In_1270,In_329);
xor U4164 (N_4164,In_1827,In_1545);
or U4165 (N_4165,In_80,In_1034);
and U4166 (N_4166,In_1484,In_473);
nor U4167 (N_4167,In_490,In_2280);
nor U4168 (N_4168,In_1253,In_966);
nor U4169 (N_4169,In_1398,In_1422);
xor U4170 (N_4170,In_1389,In_2025);
nor U4171 (N_4171,In_1106,In_627);
nand U4172 (N_4172,In_103,In_1653);
or U4173 (N_4173,In_2149,In_1107);
and U4174 (N_4174,In_504,In_524);
nand U4175 (N_4175,In_456,In_607);
or U4176 (N_4176,In_1101,In_365);
nand U4177 (N_4177,In_2205,In_1994);
and U4178 (N_4178,In_206,In_713);
nor U4179 (N_4179,In_748,In_2429);
or U4180 (N_4180,In_1934,In_377);
and U4181 (N_4181,In_226,In_2165);
nand U4182 (N_4182,In_1341,In_1242);
or U4183 (N_4183,In_583,In_829);
xor U4184 (N_4184,In_2443,In_2184);
and U4185 (N_4185,In_2408,In_371);
and U4186 (N_4186,In_1902,In_556);
and U4187 (N_4187,In_839,In_1360);
and U4188 (N_4188,In_1726,In_783);
xnor U4189 (N_4189,In_2340,In_545);
or U4190 (N_4190,In_50,In_925);
or U4191 (N_4191,In_2229,In_1807);
nand U4192 (N_4192,In_540,In_1987);
xor U4193 (N_4193,In_1418,In_2107);
nor U4194 (N_4194,In_1035,In_412);
nor U4195 (N_4195,In_43,In_30);
xnor U4196 (N_4196,In_1991,In_328);
and U4197 (N_4197,In_1000,In_1606);
xnor U4198 (N_4198,In_2096,In_1895);
nor U4199 (N_4199,In_2196,In_541);
xor U4200 (N_4200,In_1815,In_1518);
nor U4201 (N_4201,In_81,In_463);
and U4202 (N_4202,In_2161,In_140);
xor U4203 (N_4203,In_1428,In_2057);
and U4204 (N_4204,In_528,In_2140);
nand U4205 (N_4205,In_2089,In_430);
xnor U4206 (N_4206,In_2045,In_1236);
and U4207 (N_4207,In_1354,In_1080);
nor U4208 (N_4208,In_57,In_1327);
nand U4209 (N_4209,In_2134,In_993);
or U4210 (N_4210,In_1089,In_549);
nor U4211 (N_4211,In_952,In_1954);
nor U4212 (N_4212,In_1263,In_1026);
nand U4213 (N_4213,In_684,In_1411);
and U4214 (N_4214,In_1811,In_1232);
xnor U4215 (N_4215,In_1589,In_225);
xor U4216 (N_4216,In_539,In_194);
xor U4217 (N_4217,In_324,In_50);
and U4218 (N_4218,In_1548,In_1155);
xnor U4219 (N_4219,In_2323,In_717);
nor U4220 (N_4220,In_227,In_367);
nand U4221 (N_4221,In_1238,In_56);
nor U4222 (N_4222,In_792,In_1316);
or U4223 (N_4223,In_842,In_1544);
and U4224 (N_4224,In_1520,In_4);
xor U4225 (N_4225,In_1678,In_1614);
nor U4226 (N_4226,In_1537,In_164);
or U4227 (N_4227,In_1474,In_2274);
nor U4228 (N_4228,In_1454,In_975);
and U4229 (N_4229,In_2014,In_348);
nand U4230 (N_4230,In_2078,In_62);
and U4231 (N_4231,In_502,In_2037);
or U4232 (N_4232,In_2161,In_624);
or U4233 (N_4233,In_1441,In_2275);
xor U4234 (N_4234,In_2076,In_123);
nor U4235 (N_4235,In_753,In_1772);
and U4236 (N_4236,In_544,In_1967);
nor U4237 (N_4237,In_338,In_1818);
nand U4238 (N_4238,In_402,In_2081);
nand U4239 (N_4239,In_225,In_669);
xor U4240 (N_4240,In_1367,In_678);
and U4241 (N_4241,In_2315,In_1710);
nand U4242 (N_4242,In_433,In_1612);
nand U4243 (N_4243,In_1615,In_534);
xor U4244 (N_4244,In_2025,In_1878);
and U4245 (N_4245,In_667,In_1613);
nand U4246 (N_4246,In_2056,In_719);
and U4247 (N_4247,In_1857,In_1797);
nor U4248 (N_4248,In_2438,In_1812);
xor U4249 (N_4249,In_974,In_2241);
and U4250 (N_4250,In_985,In_963);
nor U4251 (N_4251,In_1525,In_494);
and U4252 (N_4252,In_2419,In_1000);
or U4253 (N_4253,In_2019,In_1065);
xor U4254 (N_4254,In_1055,In_685);
nor U4255 (N_4255,In_230,In_2093);
xor U4256 (N_4256,In_1242,In_491);
nor U4257 (N_4257,In_2042,In_315);
or U4258 (N_4258,In_1132,In_2227);
nand U4259 (N_4259,In_689,In_64);
and U4260 (N_4260,In_1811,In_2386);
or U4261 (N_4261,In_1265,In_2423);
xor U4262 (N_4262,In_1666,In_2244);
or U4263 (N_4263,In_2174,In_921);
or U4264 (N_4264,In_1195,In_1094);
and U4265 (N_4265,In_1313,In_406);
nand U4266 (N_4266,In_1779,In_550);
or U4267 (N_4267,In_1609,In_869);
or U4268 (N_4268,In_122,In_995);
and U4269 (N_4269,In_195,In_2304);
xor U4270 (N_4270,In_683,In_1497);
nand U4271 (N_4271,In_1452,In_2445);
and U4272 (N_4272,In_1707,In_1909);
or U4273 (N_4273,In_928,In_1198);
nand U4274 (N_4274,In_143,In_890);
nor U4275 (N_4275,In_1471,In_115);
nand U4276 (N_4276,In_1981,In_2105);
and U4277 (N_4277,In_1471,In_2121);
nand U4278 (N_4278,In_1095,In_2462);
nor U4279 (N_4279,In_767,In_902);
nand U4280 (N_4280,In_1656,In_1025);
nor U4281 (N_4281,In_60,In_1415);
nor U4282 (N_4282,In_559,In_1279);
or U4283 (N_4283,In_87,In_589);
nor U4284 (N_4284,In_109,In_566);
nor U4285 (N_4285,In_390,In_1532);
and U4286 (N_4286,In_976,In_95);
nand U4287 (N_4287,In_1417,In_2217);
and U4288 (N_4288,In_127,In_1997);
nand U4289 (N_4289,In_1683,In_682);
xnor U4290 (N_4290,In_1908,In_1566);
xor U4291 (N_4291,In_1341,In_1661);
nor U4292 (N_4292,In_1969,In_2411);
and U4293 (N_4293,In_1069,In_1155);
nand U4294 (N_4294,In_1982,In_2315);
xnor U4295 (N_4295,In_1604,In_351);
or U4296 (N_4296,In_1436,In_1104);
or U4297 (N_4297,In_747,In_2480);
xnor U4298 (N_4298,In_364,In_173);
nand U4299 (N_4299,In_1021,In_1880);
nor U4300 (N_4300,In_1338,In_1591);
and U4301 (N_4301,In_2021,In_1808);
nor U4302 (N_4302,In_272,In_1210);
and U4303 (N_4303,In_543,In_395);
nand U4304 (N_4304,In_1566,In_1386);
or U4305 (N_4305,In_740,In_773);
or U4306 (N_4306,In_888,In_2389);
xor U4307 (N_4307,In_255,In_396);
nor U4308 (N_4308,In_1157,In_2288);
nor U4309 (N_4309,In_1427,In_852);
nor U4310 (N_4310,In_2227,In_1796);
xor U4311 (N_4311,In_1751,In_2236);
nor U4312 (N_4312,In_1151,In_394);
xnor U4313 (N_4313,In_1444,In_1828);
nand U4314 (N_4314,In_1628,In_1983);
nand U4315 (N_4315,In_1612,In_2255);
nand U4316 (N_4316,In_2208,In_1609);
and U4317 (N_4317,In_71,In_2352);
nor U4318 (N_4318,In_2037,In_1022);
and U4319 (N_4319,In_980,In_2294);
nand U4320 (N_4320,In_1336,In_1930);
and U4321 (N_4321,In_899,In_1365);
nor U4322 (N_4322,In_512,In_1364);
and U4323 (N_4323,In_1953,In_936);
nand U4324 (N_4324,In_928,In_97);
nor U4325 (N_4325,In_2376,In_605);
and U4326 (N_4326,In_2120,In_1458);
nand U4327 (N_4327,In_1516,In_49);
or U4328 (N_4328,In_246,In_2169);
nor U4329 (N_4329,In_250,In_2441);
or U4330 (N_4330,In_1416,In_1267);
or U4331 (N_4331,In_1328,In_2081);
or U4332 (N_4332,In_1230,In_1657);
nand U4333 (N_4333,In_348,In_2244);
nor U4334 (N_4334,In_2349,In_951);
xor U4335 (N_4335,In_1832,In_1316);
xnor U4336 (N_4336,In_2334,In_853);
and U4337 (N_4337,In_952,In_2248);
or U4338 (N_4338,In_761,In_2346);
xor U4339 (N_4339,In_1287,In_1396);
and U4340 (N_4340,In_2199,In_1555);
and U4341 (N_4341,In_1074,In_265);
nand U4342 (N_4342,In_622,In_702);
nand U4343 (N_4343,In_2446,In_1208);
or U4344 (N_4344,In_373,In_472);
nor U4345 (N_4345,In_846,In_2423);
or U4346 (N_4346,In_1945,In_582);
nor U4347 (N_4347,In_220,In_1705);
nor U4348 (N_4348,In_263,In_1812);
xor U4349 (N_4349,In_654,In_879);
and U4350 (N_4350,In_876,In_555);
xnor U4351 (N_4351,In_1746,In_775);
or U4352 (N_4352,In_922,In_1600);
nand U4353 (N_4353,In_238,In_1278);
nor U4354 (N_4354,In_1954,In_1264);
nor U4355 (N_4355,In_2488,In_474);
xnor U4356 (N_4356,In_1393,In_1687);
nor U4357 (N_4357,In_38,In_647);
and U4358 (N_4358,In_2096,In_1647);
or U4359 (N_4359,In_2213,In_549);
xor U4360 (N_4360,In_420,In_1943);
nor U4361 (N_4361,In_1425,In_2083);
nand U4362 (N_4362,In_2266,In_1177);
xor U4363 (N_4363,In_2051,In_1029);
nand U4364 (N_4364,In_770,In_1375);
nor U4365 (N_4365,In_1236,In_1265);
and U4366 (N_4366,In_1683,In_692);
or U4367 (N_4367,In_2065,In_51);
nand U4368 (N_4368,In_1895,In_1569);
nand U4369 (N_4369,In_146,In_691);
nand U4370 (N_4370,In_1460,In_1235);
xor U4371 (N_4371,In_1637,In_540);
and U4372 (N_4372,In_696,In_1512);
xor U4373 (N_4373,In_1408,In_95);
nand U4374 (N_4374,In_829,In_78);
or U4375 (N_4375,In_1886,In_711);
nor U4376 (N_4376,In_671,In_2218);
xor U4377 (N_4377,In_1631,In_1275);
nor U4378 (N_4378,In_1019,In_999);
xor U4379 (N_4379,In_1202,In_1959);
nand U4380 (N_4380,In_595,In_146);
or U4381 (N_4381,In_741,In_31);
and U4382 (N_4382,In_2159,In_514);
xor U4383 (N_4383,In_667,In_1616);
nand U4384 (N_4384,In_1990,In_2114);
nor U4385 (N_4385,In_2124,In_1709);
nand U4386 (N_4386,In_594,In_2349);
and U4387 (N_4387,In_1712,In_1199);
nand U4388 (N_4388,In_1816,In_737);
nand U4389 (N_4389,In_1169,In_299);
nand U4390 (N_4390,In_117,In_389);
or U4391 (N_4391,In_935,In_275);
nand U4392 (N_4392,In_1166,In_2422);
xor U4393 (N_4393,In_329,In_147);
nor U4394 (N_4394,In_378,In_1619);
nor U4395 (N_4395,In_322,In_1970);
nor U4396 (N_4396,In_1347,In_1472);
nor U4397 (N_4397,In_1112,In_432);
nand U4398 (N_4398,In_1966,In_1270);
and U4399 (N_4399,In_1701,In_685);
xnor U4400 (N_4400,In_2117,In_280);
nand U4401 (N_4401,In_170,In_2484);
nand U4402 (N_4402,In_583,In_1748);
and U4403 (N_4403,In_1695,In_810);
nand U4404 (N_4404,In_2308,In_335);
or U4405 (N_4405,In_2262,In_2223);
xor U4406 (N_4406,In_2064,In_218);
and U4407 (N_4407,In_1926,In_1143);
nand U4408 (N_4408,In_2358,In_812);
nand U4409 (N_4409,In_550,In_752);
nor U4410 (N_4410,In_576,In_579);
xor U4411 (N_4411,In_185,In_578);
nor U4412 (N_4412,In_2298,In_2324);
nand U4413 (N_4413,In_2015,In_1051);
xor U4414 (N_4414,In_1083,In_2331);
and U4415 (N_4415,In_639,In_823);
nand U4416 (N_4416,In_2213,In_2237);
or U4417 (N_4417,In_1764,In_1691);
or U4418 (N_4418,In_1640,In_634);
nor U4419 (N_4419,In_1411,In_1967);
nand U4420 (N_4420,In_2312,In_1626);
nor U4421 (N_4421,In_969,In_2074);
xor U4422 (N_4422,In_63,In_426);
and U4423 (N_4423,In_334,In_2008);
and U4424 (N_4424,In_805,In_277);
nand U4425 (N_4425,In_1841,In_1835);
nor U4426 (N_4426,In_1174,In_2008);
xor U4427 (N_4427,In_1860,In_609);
nand U4428 (N_4428,In_1103,In_61);
and U4429 (N_4429,In_671,In_953);
or U4430 (N_4430,In_1002,In_1696);
or U4431 (N_4431,In_565,In_505);
or U4432 (N_4432,In_2463,In_642);
xor U4433 (N_4433,In_2302,In_398);
nor U4434 (N_4434,In_367,In_751);
nor U4435 (N_4435,In_211,In_1257);
nand U4436 (N_4436,In_1555,In_2443);
xor U4437 (N_4437,In_2339,In_1097);
nand U4438 (N_4438,In_1979,In_891);
and U4439 (N_4439,In_1403,In_2201);
nor U4440 (N_4440,In_1823,In_1928);
nand U4441 (N_4441,In_538,In_2025);
nand U4442 (N_4442,In_1072,In_860);
nor U4443 (N_4443,In_2441,In_584);
nand U4444 (N_4444,In_2178,In_1459);
xnor U4445 (N_4445,In_1808,In_991);
nand U4446 (N_4446,In_264,In_602);
nand U4447 (N_4447,In_2460,In_1336);
and U4448 (N_4448,In_49,In_1061);
or U4449 (N_4449,In_2447,In_7);
xnor U4450 (N_4450,In_2223,In_823);
nor U4451 (N_4451,In_1456,In_1006);
xnor U4452 (N_4452,In_783,In_1727);
xnor U4453 (N_4453,In_869,In_474);
xor U4454 (N_4454,In_1406,In_398);
nand U4455 (N_4455,In_1855,In_2410);
xor U4456 (N_4456,In_65,In_698);
and U4457 (N_4457,In_2204,In_1180);
nand U4458 (N_4458,In_1429,In_930);
nand U4459 (N_4459,In_1233,In_396);
xnor U4460 (N_4460,In_2239,In_1102);
and U4461 (N_4461,In_73,In_966);
nor U4462 (N_4462,In_307,In_2130);
nand U4463 (N_4463,In_1723,In_1810);
nor U4464 (N_4464,In_1372,In_150);
nand U4465 (N_4465,In_787,In_1667);
xor U4466 (N_4466,In_118,In_658);
or U4467 (N_4467,In_2479,In_2339);
nor U4468 (N_4468,In_1371,In_2145);
xnor U4469 (N_4469,In_1554,In_2479);
nor U4470 (N_4470,In_430,In_367);
and U4471 (N_4471,In_1940,In_1827);
nor U4472 (N_4472,In_169,In_2211);
xnor U4473 (N_4473,In_2048,In_2440);
or U4474 (N_4474,In_2151,In_749);
nor U4475 (N_4475,In_586,In_502);
xnor U4476 (N_4476,In_1929,In_83);
and U4477 (N_4477,In_1167,In_1716);
nor U4478 (N_4478,In_33,In_675);
nand U4479 (N_4479,In_1903,In_1678);
xor U4480 (N_4480,In_1016,In_2211);
and U4481 (N_4481,In_2097,In_1861);
and U4482 (N_4482,In_1070,In_1291);
or U4483 (N_4483,In_1095,In_1775);
nand U4484 (N_4484,In_107,In_1168);
and U4485 (N_4485,In_266,In_1461);
nor U4486 (N_4486,In_2136,In_489);
and U4487 (N_4487,In_985,In_1678);
xor U4488 (N_4488,In_1659,In_1408);
xnor U4489 (N_4489,In_745,In_612);
nand U4490 (N_4490,In_1560,In_444);
or U4491 (N_4491,In_2175,In_1056);
and U4492 (N_4492,In_578,In_2211);
nor U4493 (N_4493,In_1759,In_647);
nand U4494 (N_4494,In_2454,In_1628);
nand U4495 (N_4495,In_442,In_1004);
nor U4496 (N_4496,In_2204,In_606);
nor U4497 (N_4497,In_1179,In_589);
and U4498 (N_4498,In_2353,In_1724);
or U4499 (N_4499,In_2111,In_2438);
nand U4500 (N_4500,In_177,In_821);
nand U4501 (N_4501,In_921,In_83);
and U4502 (N_4502,In_1575,In_2433);
nor U4503 (N_4503,In_368,In_1636);
nand U4504 (N_4504,In_128,In_465);
xnor U4505 (N_4505,In_2294,In_494);
nor U4506 (N_4506,In_145,In_1842);
nand U4507 (N_4507,In_871,In_165);
and U4508 (N_4508,In_1696,In_2070);
xnor U4509 (N_4509,In_373,In_630);
xnor U4510 (N_4510,In_630,In_2494);
nor U4511 (N_4511,In_1194,In_398);
nand U4512 (N_4512,In_1363,In_2392);
nor U4513 (N_4513,In_2130,In_362);
and U4514 (N_4514,In_1519,In_45);
nand U4515 (N_4515,In_1673,In_1721);
nand U4516 (N_4516,In_2239,In_1987);
and U4517 (N_4517,In_1047,In_1898);
nor U4518 (N_4518,In_1297,In_2305);
or U4519 (N_4519,In_2111,In_1523);
and U4520 (N_4520,In_1495,In_596);
nand U4521 (N_4521,In_126,In_211);
nor U4522 (N_4522,In_2436,In_741);
and U4523 (N_4523,In_213,In_1510);
nand U4524 (N_4524,In_1619,In_771);
nor U4525 (N_4525,In_1861,In_634);
xor U4526 (N_4526,In_886,In_827);
nand U4527 (N_4527,In_2151,In_2177);
and U4528 (N_4528,In_2152,In_2096);
or U4529 (N_4529,In_2088,In_909);
nand U4530 (N_4530,In_2405,In_165);
nor U4531 (N_4531,In_1863,In_1966);
nand U4532 (N_4532,In_840,In_1843);
xor U4533 (N_4533,In_1516,In_377);
and U4534 (N_4534,In_1495,In_1707);
nand U4535 (N_4535,In_180,In_2017);
nand U4536 (N_4536,In_324,In_1081);
and U4537 (N_4537,In_1346,In_2125);
xnor U4538 (N_4538,In_2169,In_1218);
nand U4539 (N_4539,In_1656,In_2107);
nand U4540 (N_4540,In_1639,In_576);
nand U4541 (N_4541,In_2271,In_1696);
and U4542 (N_4542,In_989,In_1059);
or U4543 (N_4543,In_1370,In_1256);
nor U4544 (N_4544,In_383,In_740);
nor U4545 (N_4545,In_2148,In_550);
xnor U4546 (N_4546,In_242,In_1404);
and U4547 (N_4547,In_1070,In_1810);
or U4548 (N_4548,In_86,In_2147);
nor U4549 (N_4549,In_941,In_1450);
and U4550 (N_4550,In_1736,In_1206);
xor U4551 (N_4551,In_1443,In_887);
and U4552 (N_4552,In_252,In_183);
and U4553 (N_4553,In_1292,In_1114);
and U4554 (N_4554,In_1872,In_2375);
nand U4555 (N_4555,In_2402,In_1730);
nor U4556 (N_4556,In_2462,In_2164);
nand U4557 (N_4557,In_1892,In_241);
nand U4558 (N_4558,In_1584,In_1440);
or U4559 (N_4559,In_969,In_1303);
or U4560 (N_4560,In_1499,In_948);
or U4561 (N_4561,In_1810,In_815);
nor U4562 (N_4562,In_220,In_1626);
nor U4563 (N_4563,In_804,In_15);
nand U4564 (N_4564,In_2118,In_463);
and U4565 (N_4565,In_1336,In_564);
nor U4566 (N_4566,In_1846,In_40);
nor U4567 (N_4567,In_1639,In_238);
nand U4568 (N_4568,In_1962,In_895);
nand U4569 (N_4569,In_1162,In_2081);
or U4570 (N_4570,In_851,In_374);
or U4571 (N_4571,In_2367,In_512);
and U4572 (N_4572,In_696,In_338);
xnor U4573 (N_4573,In_60,In_445);
or U4574 (N_4574,In_1329,In_681);
and U4575 (N_4575,In_555,In_692);
and U4576 (N_4576,In_148,In_1321);
and U4577 (N_4577,In_1946,In_353);
nor U4578 (N_4578,In_2093,In_2341);
nand U4579 (N_4579,In_1308,In_1482);
nor U4580 (N_4580,In_1403,In_1296);
nor U4581 (N_4581,In_2088,In_2497);
nand U4582 (N_4582,In_373,In_1180);
nor U4583 (N_4583,In_238,In_1256);
xnor U4584 (N_4584,In_422,In_1996);
nand U4585 (N_4585,In_2076,In_612);
and U4586 (N_4586,In_850,In_705);
nor U4587 (N_4587,In_2480,In_2006);
xor U4588 (N_4588,In_1988,In_2372);
or U4589 (N_4589,In_2351,In_1342);
nand U4590 (N_4590,In_1375,In_1996);
nor U4591 (N_4591,In_690,In_32);
xnor U4592 (N_4592,In_653,In_192);
and U4593 (N_4593,In_2216,In_1320);
nor U4594 (N_4594,In_917,In_20);
nand U4595 (N_4595,In_956,In_1169);
nor U4596 (N_4596,In_2,In_1109);
xor U4597 (N_4597,In_1985,In_2318);
nand U4598 (N_4598,In_2458,In_738);
nand U4599 (N_4599,In_1623,In_1515);
and U4600 (N_4600,In_71,In_1965);
and U4601 (N_4601,In_605,In_1570);
nor U4602 (N_4602,In_1916,In_929);
xor U4603 (N_4603,In_660,In_1844);
nor U4604 (N_4604,In_1778,In_2491);
nand U4605 (N_4605,In_2485,In_2279);
or U4606 (N_4606,In_2173,In_1593);
nor U4607 (N_4607,In_1218,In_767);
xor U4608 (N_4608,In_1982,In_1983);
xnor U4609 (N_4609,In_1333,In_47);
or U4610 (N_4610,In_2294,In_1949);
or U4611 (N_4611,In_1452,In_1343);
nand U4612 (N_4612,In_1696,In_1908);
xnor U4613 (N_4613,In_1404,In_2288);
and U4614 (N_4614,In_1944,In_1568);
or U4615 (N_4615,In_679,In_2061);
xor U4616 (N_4616,In_1660,In_1751);
nand U4617 (N_4617,In_2175,In_2106);
and U4618 (N_4618,In_184,In_2058);
xor U4619 (N_4619,In_2274,In_809);
xnor U4620 (N_4620,In_1967,In_503);
or U4621 (N_4621,In_995,In_431);
nand U4622 (N_4622,In_1360,In_490);
and U4623 (N_4623,In_300,In_2013);
or U4624 (N_4624,In_2251,In_251);
nand U4625 (N_4625,In_960,In_658);
or U4626 (N_4626,In_1976,In_738);
and U4627 (N_4627,In_807,In_2016);
nor U4628 (N_4628,In_11,In_2263);
or U4629 (N_4629,In_1697,In_2214);
nand U4630 (N_4630,In_611,In_2355);
xor U4631 (N_4631,In_1355,In_738);
and U4632 (N_4632,In_968,In_1348);
xor U4633 (N_4633,In_2288,In_2308);
or U4634 (N_4634,In_923,In_693);
xor U4635 (N_4635,In_1987,In_2062);
nor U4636 (N_4636,In_748,In_536);
xor U4637 (N_4637,In_123,In_1264);
and U4638 (N_4638,In_2096,In_2390);
nand U4639 (N_4639,In_1376,In_475);
nor U4640 (N_4640,In_1837,In_2068);
or U4641 (N_4641,In_805,In_1154);
and U4642 (N_4642,In_1841,In_1580);
xnor U4643 (N_4643,In_2286,In_785);
nand U4644 (N_4644,In_58,In_703);
xor U4645 (N_4645,In_2483,In_994);
or U4646 (N_4646,In_2024,In_651);
and U4647 (N_4647,In_782,In_2414);
nor U4648 (N_4648,In_1748,In_1858);
or U4649 (N_4649,In_2040,In_2237);
or U4650 (N_4650,In_1844,In_2301);
xnor U4651 (N_4651,In_763,In_1325);
and U4652 (N_4652,In_964,In_1060);
nor U4653 (N_4653,In_539,In_750);
or U4654 (N_4654,In_767,In_2316);
nor U4655 (N_4655,In_1325,In_1258);
or U4656 (N_4656,In_391,In_2217);
and U4657 (N_4657,In_2388,In_1822);
nor U4658 (N_4658,In_1797,In_1184);
nor U4659 (N_4659,In_233,In_2207);
nor U4660 (N_4660,In_1082,In_1254);
xnor U4661 (N_4661,In_1649,In_1773);
or U4662 (N_4662,In_1788,In_2332);
nand U4663 (N_4663,In_322,In_1937);
nand U4664 (N_4664,In_2367,In_171);
nor U4665 (N_4665,In_751,In_1607);
and U4666 (N_4666,In_2321,In_1667);
nand U4667 (N_4667,In_191,In_2129);
nand U4668 (N_4668,In_118,In_1680);
and U4669 (N_4669,In_223,In_1528);
or U4670 (N_4670,In_870,In_163);
nand U4671 (N_4671,In_2234,In_2466);
xor U4672 (N_4672,In_1349,In_1689);
nor U4673 (N_4673,In_486,In_603);
and U4674 (N_4674,In_616,In_860);
or U4675 (N_4675,In_630,In_757);
xor U4676 (N_4676,In_1422,In_1463);
and U4677 (N_4677,In_2459,In_1339);
and U4678 (N_4678,In_527,In_1389);
and U4679 (N_4679,In_2489,In_188);
nand U4680 (N_4680,In_2365,In_839);
xor U4681 (N_4681,In_2423,In_792);
or U4682 (N_4682,In_1645,In_1937);
nor U4683 (N_4683,In_2152,In_111);
or U4684 (N_4684,In_1840,In_215);
or U4685 (N_4685,In_504,In_2324);
nand U4686 (N_4686,In_1327,In_1691);
or U4687 (N_4687,In_22,In_369);
xor U4688 (N_4688,In_836,In_538);
or U4689 (N_4689,In_1562,In_2228);
or U4690 (N_4690,In_341,In_334);
nor U4691 (N_4691,In_2365,In_308);
nor U4692 (N_4692,In_1305,In_1005);
or U4693 (N_4693,In_2436,In_1324);
and U4694 (N_4694,In_1310,In_1279);
nor U4695 (N_4695,In_689,In_1184);
nand U4696 (N_4696,In_1501,In_822);
nor U4697 (N_4697,In_166,In_472);
nand U4698 (N_4698,In_2311,In_1306);
nand U4699 (N_4699,In_1954,In_88);
nor U4700 (N_4700,In_325,In_402);
nor U4701 (N_4701,In_19,In_1806);
and U4702 (N_4702,In_245,In_1813);
nand U4703 (N_4703,In_1972,In_1098);
xor U4704 (N_4704,In_1549,In_483);
nand U4705 (N_4705,In_1432,In_2159);
nand U4706 (N_4706,In_553,In_138);
nand U4707 (N_4707,In_2185,In_1862);
or U4708 (N_4708,In_363,In_1835);
or U4709 (N_4709,In_1683,In_2428);
nor U4710 (N_4710,In_2320,In_2316);
nor U4711 (N_4711,In_2151,In_2235);
or U4712 (N_4712,In_1686,In_1973);
or U4713 (N_4713,In_1605,In_1622);
and U4714 (N_4714,In_1077,In_1267);
nor U4715 (N_4715,In_326,In_862);
and U4716 (N_4716,In_1757,In_478);
nand U4717 (N_4717,In_1299,In_1009);
nor U4718 (N_4718,In_2004,In_2267);
nor U4719 (N_4719,In_1393,In_1809);
nor U4720 (N_4720,In_1526,In_264);
xor U4721 (N_4721,In_1633,In_1987);
nor U4722 (N_4722,In_1618,In_1901);
nand U4723 (N_4723,In_406,In_1719);
nor U4724 (N_4724,In_1769,In_1186);
xor U4725 (N_4725,In_1851,In_2231);
nand U4726 (N_4726,In_1585,In_469);
nor U4727 (N_4727,In_1143,In_1152);
xnor U4728 (N_4728,In_1676,In_1835);
and U4729 (N_4729,In_408,In_291);
nor U4730 (N_4730,In_1085,In_1759);
xor U4731 (N_4731,In_1007,In_2315);
nor U4732 (N_4732,In_569,In_93);
nand U4733 (N_4733,In_2265,In_1624);
nor U4734 (N_4734,In_169,In_2376);
xnor U4735 (N_4735,In_178,In_1056);
or U4736 (N_4736,In_337,In_415);
nand U4737 (N_4737,In_1271,In_2293);
nor U4738 (N_4738,In_159,In_553);
nand U4739 (N_4739,In_652,In_542);
xnor U4740 (N_4740,In_34,In_877);
xnor U4741 (N_4741,In_552,In_2153);
xor U4742 (N_4742,In_649,In_1815);
and U4743 (N_4743,In_960,In_803);
and U4744 (N_4744,In_1050,In_1068);
and U4745 (N_4745,In_2154,In_71);
nand U4746 (N_4746,In_541,In_1379);
nand U4747 (N_4747,In_1304,In_228);
and U4748 (N_4748,In_1734,In_740);
nor U4749 (N_4749,In_469,In_1791);
nor U4750 (N_4750,In_21,In_1509);
xor U4751 (N_4751,In_2141,In_2256);
xor U4752 (N_4752,In_2282,In_1833);
nand U4753 (N_4753,In_986,In_370);
or U4754 (N_4754,In_1699,In_643);
xnor U4755 (N_4755,In_1779,In_2071);
or U4756 (N_4756,In_1719,In_858);
nand U4757 (N_4757,In_133,In_1462);
or U4758 (N_4758,In_19,In_1698);
nand U4759 (N_4759,In_766,In_2271);
xnor U4760 (N_4760,In_2346,In_1159);
and U4761 (N_4761,In_341,In_70);
or U4762 (N_4762,In_764,In_102);
and U4763 (N_4763,In_1563,In_893);
nand U4764 (N_4764,In_1047,In_2334);
nor U4765 (N_4765,In_2308,In_316);
nor U4766 (N_4766,In_653,In_1662);
nor U4767 (N_4767,In_1165,In_1530);
nor U4768 (N_4768,In_932,In_970);
or U4769 (N_4769,In_553,In_2217);
xor U4770 (N_4770,In_179,In_167);
or U4771 (N_4771,In_1756,In_872);
nand U4772 (N_4772,In_131,In_255);
xor U4773 (N_4773,In_1933,In_2482);
nor U4774 (N_4774,In_1212,In_248);
and U4775 (N_4775,In_631,In_347);
or U4776 (N_4776,In_1515,In_651);
xor U4777 (N_4777,In_1578,In_71);
nor U4778 (N_4778,In_1951,In_2362);
xnor U4779 (N_4779,In_114,In_1600);
or U4780 (N_4780,In_1003,In_1918);
nand U4781 (N_4781,In_938,In_2356);
nor U4782 (N_4782,In_2343,In_2497);
xnor U4783 (N_4783,In_785,In_38);
xor U4784 (N_4784,In_1583,In_866);
and U4785 (N_4785,In_70,In_1668);
and U4786 (N_4786,In_2087,In_563);
nand U4787 (N_4787,In_191,In_1392);
nor U4788 (N_4788,In_1658,In_87);
and U4789 (N_4789,In_2151,In_843);
nand U4790 (N_4790,In_2196,In_941);
nor U4791 (N_4791,In_873,In_1102);
nor U4792 (N_4792,In_1118,In_1046);
nor U4793 (N_4793,In_373,In_1071);
xnor U4794 (N_4794,In_2214,In_747);
or U4795 (N_4795,In_181,In_1516);
nor U4796 (N_4796,In_2135,In_2062);
or U4797 (N_4797,In_754,In_637);
nor U4798 (N_4798,In_861,In_1718);
xnor U4799 (N_4799,In_1757,In_2403);
nand U4800 (N_4800,In_1316,In_1667);
xor U4801 (N_4801,In_341,In_485);
nand U4802 (N_4802,In_2203,In_862);
or U4803 (N_4803,In_400,In_542);
or U4804 (N_4804,In_587,In_323);
and U4805 (N_4805,In_2019,In_1154);
xor U4806 (N_4806,In_1676,In_1960);
and U4807 (N_4807,In_2185,In_1549);
nand U4808 (N_4808,In_323,In_2088);
nand U4809 (N_4809,In_523,In_1959);
nor U4810 (N_4810,In_2440,In_411);
nor U4811 (N_4811,In_1572,In_447);
and U4812 (N_4812,In_1900,In_1457);
nand U4813 (N_4813,In_1040,In_428);
and U4814 (N_4814,In_2157,In_1596);
nor U4815 (N_4815,In_1491,In_1514);
xor U4816 (N_4816,In_2478,In_171);
nor U4817 (N_4817,In_1343,In_2005);
and U4818 (N_4818,In_2151,In_507);
nor U4819 (N_4819,In_2259,In_2416);
xor U4820 (N_4820,In_1712,In_1189);
nor U4821 (N_4821,In_396,In_1562);
nand U4822 (N_4822,In_939,In_1697);
or U4823 (N_4823,In_2438,In_1236);
nand U4824 (N_4824,In_1033,In_2237);
xnor U4825 (N_4825,In_1413,In_2485);
nand U4826 (N_4826,In_1156,In_2269);
nand U4827 (N_4827,In_1121,In_1280);
and U4828 (N_4828,In_214,In_1376);
or U4829 (N_4829,In_2348,In_927);
nor U4830 (N_4830,In_745,In_406);
nand U4831 (N_4831,In_2302,In_1486);
and U4832 (N_4832,In_22,In_2234);
nor U4833 (N_4833,In_811,In_2168);
or U4834 (N_4834,In_434,In_1106);
xor U4835 (N_4835,In_1636,In_841);
xor U4836 (N_4836,In_2112,In_1676);
nand U4837 (N_4837,In_366,In_1972);
nand U4838 (N_4838,In_892,In_528);
or U4839 (N_4839,In_1762,In_1206);
or U4840 (N_4840,In_1925,In_1588);
nor U4841 (N_4841,In_1999,In_1080);
nand U4842 (N_4842,In_1882,In_1777);
nor U4843 (N_4843,In_377,In_639);
or U4844 (N_4844,In_1049,In_1634);
and U4845 (N_4845,In_162,In_1752);
nor U4846 (N_4846,In_162,In_508);
nor U4847 (N_4847,In_203,In_860);
and U4848 (N_4848,In_1265,In_489);
nand U4849 (N_4849,In_1289,In_2299);
or U4850 (N_4850,In_790,In_2449);
and U4851 (N_4851,In_1146,In_2130);
and U4852 (N_4852,In_2343,In_2466);
nor U4853 (N_4853,In_668,In_1277);
and U4854 (N_4854,In_948,In_683);
and U4855 (N_4855,In_3,In_459);
nand U4856 (N_4856,In_1987,In_2138);
nand U4857 (N_4857,In_454,In_1738);
nand U4858 (N_4858,In_282,In_867);
nand U4859 (N_4859,In_2487,In_279);
nand U4860 (N_4860,In_1548,In_2086);
nor U4861 (N_4861,In_357,In_2321);
or U4862 (N_4862,In_1185,In_1377);
nand U4863 (N_4863,In_105,In_697);
nor U4864 (N_4864,In_182,In_1123);
nor U4865 (N_4865,In_241,In_516);
or U4866 (N_4866,In_1842,In_2065);
nor U4867 (N_4867,In_541,In_1646);
or U4868 (N_4868,In_810,In_1004);
nor U4869 (N_4869,In_755,In_437);
nand U4870 (N_4870,In_1835,In_256);
or U4871 (N_4871,In_223,In_216);
nand U4872 (N_4872,In_1490,In_1450);
and U4873 (N_4873,In_495,In_715);
nand U4874 (N_4874,In_718,In_1260);
xnor U4875 (N_4875,In_1098,In_1688);
nand U4876 (N_4876,In_2280,In_747);
xor U4877 (N_4877,In_672,In_1846);
nor U4878 (N_4878,In_2055,In_1810);
and U4879 (N_4879,In_842,In_16);
nor U4880 (N_4880,In_2488,In_1056);
nor U4881 (N_4881,In_1646,In_2159);
and U4882 (N_4882,In_924,In_380);
nand U4883 (N_4883,In_842,In_2163);
nor U4884 (N_4884,In_1709,In_1043);
nor U4885 (N_4885,In_1324,In_1820);
and U4886 (N_4886,In_1185,In_2201);
or U4887 (N_4887,In_196,In_1676);
xor U4888 (N_4888,In_2139,In_405);
and U4889 (N_4889,In_2398,In_1645);
xor U4890 (N_4890,In_684,In_1802);
nor U4891 (N_4891,In_1360,In_1839);
nor U4892 (N_4892,In_292,In_1684);
and U4893 (N_4893,In_2348,In_1542);
or U4894 (N_4894,In_883,In_1330);
or U4895 (N_4895,In_131,In_675);
and U4896 (N_4896,In_1034,In_185);
xor U4897 (N_4897,In_370,In_1427);
nor U4898 (N_4898,In_1546,In_198);
nand U4899 (N_4899,In_2493,In_2497);
and U4900 (N_4900,In_1868,In_862);
nand U4901 (N_4901,In_2454,In_1509);
and U4902 (N_4902,In_2090,In_1557);
and U4903 (N_4903,In_1504,In_1573);
or U4904 (N_4904,In_266,In_583);
nor U4905 (N_4905,In_1110,In_1295);
or U4906 (N_4906,In_172,In_120);
nor U4907 (N_4907,In_197,In_45);
nor U4908 (N_4908,In_1578,In_1297);
or U4909 (N_4909,In_660,In_1799);
xor U4910 (N_4910,In_467,In_828);
nor U4911 (N_4911,In_1933,In_79);
xor U4912 (N_4912,In_1859,In_151);
or U4913 (N_4913,In_2416,In_381);
nand U4914 (N_4914,In_2162,In_370);
nor U4915 (N_4915,In_1383,In_1109);
nor U4916 (N_4916,In_175,In_1630);
nand U4917 (N_4917,In_2135,In_2378);
xor U4918 (N_4918,In_2257,In_778);
xnor U4919 (N_4919,In_1675,In_1252);
and U4920 (N_4920,In_2327,In_932);
nor U4921 (N_4921,In_1990,In_864);
nor U4922 (N_4922,In_2052,In_337);
and U4923 (N_4923,In_445,In_255);
or U4924 (N_4924,In_1698,In_692);
nand U4925 (N_4925,In_1053,In_940);
xor U4926 (N_4926,In_2111,In_2431);
and U4927 (N_4927,In_2290,In_1268);
and U4928 (N_4928,In_1109,In_2301);
or U4929 (N_4929,In_147,In_760);
nand U4930 (N_4930,In_1488,In_1830);
nor U4931 (N_4931,In_499,In_324);
xnor U4932 (N_4932,In_787,In_1618);
nand U4933 (N_4933,In_1803,In_2236);
and U4934 (N_4934,In_971,In_1282);
nand U4935 (N_4935,In_959,In_1197);
nand U4936 (N_4936,In_777,In_730);
or U4937 (N_4937,In_2370,In_1283);
or U4938 (N_4938,In_1711,In_1156);
nor U4939 (N_4939,In_2366,In_456);
or U4940 (N_4940,In_243,In_1731);
nand U4941 (N_4941,In_2154,In_393);
nand U4942 (N_4942,In_650,In_2009);
xor U4943 (N_4943,In_1792,In_1327);
nand U4944 (N_4944,In_695,In_1506);
nor U4945 (N_4945,In_1863,In_438);
xnor U4946 (N_4946,In_757,In_1203);
xnor U4947 (N_4947,In_2178,In_736);
xor U4948 (N_4948,In_1790,In_1723);
nand U4949 (N_4949,In_44,In_1242);
and U4950 (N_4950,In_1458,In_2452);
nor U4951 (N_4951,In_157,In_2478);
xor U4952 (N_4952,In_538,In_1820);
nand U4953 (N_4953,In_312,In_299);
nand U4954 (N_4954,In_2052,In_2470);
nand U4955 (N_4955,In_1138,In_1506);
xor U4956 (N_4956,In_1135,In_574);
nor U4957 (N_4957,In_508,In_1795);
or U4958 (N_4958,In_2276,In_2121);
and U4959 (N_4959,In_167,In_711);
nor U4960 (N_4960,In_2042,In_636);
and U4961 (N_4961,In_1148,In_198);
or U4962 (N_4962,In_554,In_1662);
and U4963 (N_4963,In_2425,In_394);
nor U4964 (N_4964,In_482,In_643);
nand U4965 (N_4965,In_1909,In_899);
and U4966 (N_4966,In_121,In_1714);
nand U4967 (N_4967,In_1981,In_781);
xor U4968 (N_4968,In_1070,In_867);
xor U4969 (N_4969,In_419,In_131);
or U4970 (N_4970,In_97,In_1259);
nor U4971 (N_4971,In_2461,In_878);
or U4972 (N_4972,In_1255,In_2270);
xnor U4973 (N_4973,In_2435,In_2425);
or U4974 (N_4974,In_79,In_1205);
or U4975 (N_4975,In_642,In_546);
and U4976 (N_4976,In_911,In_2275);
and U4977 (N_4977,In_2250,In_874);
xor U4978 (N_4978,In_53,In_1866);
xor U4979 (N_4979,In_66,In_1199);
or U4980 (N_4980,In_2150,In_694);
or U4981 (N_4981,In_454,In_1578);
or U4982 (N_4982,In_1732,In_2157);
or U4983 (N_4983,In_2014,In_529);
and U4984 (N_4984,In_66,In_2330);
nand U4985 (N_4985,In_2464,In_1791);
or U4986 (N_4986,In_2039,In_2310);
xnor U4987 (N_4987,In_1926,In_201);
nand U4988 (N_4988,In_2380,In_719);
xnor U4989 (N_4989,In_208,In_204);
nor U4990 (N_4990,In_1134,In_1299);
nor U4991 (N_4991,In_1012,In_1821);
xor U4992 (N_4992,In_879,In_1579);
nor U4993 (N_4993,In_2339,In_784);
and U4994 (N_4994,In_96,In_2120);
and U4995 (N_4995,In_575,In_1712);
or U4996 (N_4996,In_51,In_1196);
or U4997 (N_4997,In_434,In_1644);
nor U4998 (N_4998,In_69,In_1815);
and U4999 (N_4999,In_2066,In_1057);
or U5000 (N_5000,N_1140,N_1354);
nor U5001 (N_5001,N_749,N_3267);
xnor U5002 (N_5002,N_2379,N_150);
nand U5003 (N_5003,N_2959,N_906);
nand U5004 (N_5004,N_3298,N_4442);
nor U5005 (N_5005,N_4264,N_2180);
and U5006 (N_5006,N_2672,N_198);
nand U5007 (N_5007,N_4836,N_615);
or U5008 (N_5008,N_3436,N_2851);
or U5009 (N_5009,N_4583,N_1529);
and U5010 (N_5010,N_1746,N_2441);
nor U5011 (N_5011,N_2384,N_3212);
or U5012 (N_5012,N_3447,N_4184);
or U5013 (N_5013,N_2288,N_2267);
or U5014 (N_5014,N_3577,N_1032);
and U5015 (N_5015,N_3557,N_4538);
and U5016 (N_5016,N_2277,N_2624);
nand U5017 (N_5017,N_548,N_3857);
or U5018 (N_5018,N_1146,N_3337);
nand U5019 (N_5019,N_4979,N_874);
or U5020 (N_5020,N_4699,N_1420);
or U5021 (N_5021,N_1644,N_4429);
xor U5022 (N_5022,N_3314,N_1607);
and U5023 (N_5023,N_1907,N_2720);
or U5024 (N_5024,N_2114,N_764);
or U5025 (N_5025,N_592,N_4320);
and U5026 (N_5026,N_2460,N_3560);
xnor U5027 (N_5027,N_1669,N_3444);
nor U5028 (N_5028,N_2902,N_1360);
xor U5029 (N_5029,N_1627,N_3978);
and U5030 (N_5030,N_480,N_1443);
xor U5031 (N_5031,N_4797,N_1473);
or U5032 (N_5032,N_2066,N_420);
or U5033 (N_5033,N_308,N_1348);
xnor U5034 (N_5034,N_2370,N_3156);
xnor U5035 (N_5035,N_2047,N_3083);
nor U5036 (N_5036,N_2589,N_335);
or U5037 (N_5037,N_2548,N_3986);
nand U5038 (N_5038,N_4052,N_128);
nand U5039 (N_5039,N_805,N_948);
and U5040 (N_5040,N_4448,N_3047);
and U5041 (N_5041,N_1173,N_3705);
or U5042 (N_5042,N_4917,N_2286);
nor U5043 (N_5043,N_3433,N_2103);
or U5044 (N_5044,N_4072,N_850);
xor U5045 (N_5045,N_1616,N_3663);
nor U5046 (N_5046,N_4712,N_3606);
or U5047 (N_5047,N_216,N_2917);
xnor U5048 (N_5048,N_732,N_13);
nor U5049 (N_5049,N_1688,N_3654);
nor U5050 (N_5050,N_2898,N_713);
nand U5051 (N_5051,N_1500,N_3332);
xnor U5052 (N_5052,N_2492,N_233);
and U5053 (N_5053,N_3140,N_291);
nor U5054 (N_5054,N_2542,N_2651);
and U5055 (N_5055,N_529,N_4819);
or U5056 (N_5056,N_1437,N_4507);
or U5057 (N_5057,N_4952,N_998);
nand U5058 (N_5058,N_750,N_2366);
nor U5059 (N_5059,N_3991,N_4643);
xor U5060 (N_5060,N_2049,N_3266);
nand U5061 (N_5061,N_1301,N_1612);
and U5062 (N_5062,N_309,N_3116);
or U5063 (N_5063,N_481,N_1101);
nand U5064 (N_5064,N_4898,N_3859);
nand U5065 (N_5065,N_465,N_3272);
and U5066 (N_5066,N_984,N_63);
or U5067 (N_5067,N_1536,N_3133);
xor U5068 (N_5068,N_2852,N_2376);
nand U5069 (N_5069,N_3067,N_2044);
and U5070 (N_5070,N_390,N_2075);
nand U5071 (N_5071,N_28,N_3515);
and U5072 (N_5072,N_4417,N_3791);
nor U5073 (N_5073,N_2887,N_1608);
and U5074 (N_5074,N_441,N_25);
nand U5075 (N_5075,N_2908,N_4906);
nand U5076 (N_5076,N_2239,N_342);
xnor U5077 (N_5077,N_1753,N_2298);
or U5078 (N_5078,N_56,N_4639);
or U5079 (N_5079,N_1454,N_1047);
and U5080 (N_5080,N_859,N_4598);
xnor U5081 (N_5081,N_1458,N_1187);
nor U5082 (N_5082,N_3412,N_1105);
or U5083 (N_5083,N_2956,N_4081);
and U5084 (N_5084,N_1363,N_606);
xor U5085 (N_5085,N_3463,N_3462);
nor U5086 (N_5086,N_2979,N_2778);
and U5087 (N_5087,N_313,N_3699);
nand U5088 (N_5088,N_3366,N_1957);
and U5089 (N_5089,N_458,N_74);
xor U5090 (N_5090,N_1118,N_2832);
nand U5091 (N_5091,N_2782,N_2743);
and U5092 (N_5092,N_2570,N_1809);
nand U5093 (N_5093,N_4347,N_1453);
or U5094 (N_5094,N_973,N_3346);
or U5095 (N_5095,N_3260,N_3510);
nand U5096 (N_5096,N_1048,N_92);
xor U5097 (N_5097,N_2304,N_4541);
and U5098 (N_5098,N_2718,N_4140);
and U5099 (N_5099,N_4933,N_1569);
nor U5100 (N_5100,N_2178,N_4312);
nand U5101 (N_5101,N_536,N_11);
or U5102 (N_5102,N_3860,N_4469);
xor U5103 (N_5103,N_1748,N_453);
nand U5104 (N_5104,N_4498,N_4694);
nand U5105 (N_5105,N_3851,N_3293);
or U5106 (N_5106,N_392,N_559);
nand U5107 (N_5107,N_272,N_4609);
and U5108 (N_5108,N_2777,N_2265);
or U5109 (N_5109,N_2390,N_1252);
xor U5110 (N_5110,N_2000,N_2164);
xor U5111 (N_5111,N_1883,N_642);
xor U5112 (N_5112,N_2546,N_774);
nand U5113 (N_5113,N_2061,N_3007);
nand U5114 (N_5114,N_1787,N_1046);
and U5115 (N_5115,N_1027,N_1729);
or U5116 (N_5116,N_2190,N_617);
and U5117 (N_5117,N_3232,N_3820);
and U5118 (N_5118,N_2791,N_3564);
and U5119 (N_5119,N_3279,N_4311);
xnor U5120 (N_5120,N_588,N_681);
nor U5121 (N_5121,N_3052,N_719);
and U5122 (N_5122,N_4341,N_3525);
and U5123 (N_5123,N_2412,N_3565);
or U5124 (N_5124,N_3159,N_4578);
nor U5125 (N_5125,N_789,N_4087);
or U5126 (N_5126,N_1094,N_2395);
xor U5127 (N_5127,N_1342,N_274);
nand U5128 (N_5128,N_4229,N_4503);
nor U5129 (N_5129,N_4099,N_4425);
nand U5130 (N_5130,N_4431,N_2312);
or U5131 (N_5131,N_1509,N_3947);
xor U5132 (N_5132,N_1582,N_3530);
and U5133 (N_5133,N_1829,N_1001);
nor U5134 (N_5134,N_1516,N_171);
xor U5135 (N_5135,N_1735,N_2358);
and U5136 (N_5136,N_936,N_3326);
and U5137 (N_5137,N_3828,N_621);
nand U5138 (N_5138,N_682,N_2435);
nor U5139 (N_5139,N_2580,N_3782);
or U5140 (N_5140,N_4905,N_464);
xnor U5141 (N_5141,N_1738,N_4562);
nor U5142 (N_5142,N_3125,N_1479);
nor U5143 (N_5143,N_1137,N_4406);
nand U5144 (N_5144,N_1990,N_2954);
nand U5145 (N_5145,N_1179,N_1546);
nor U5146 (N_5146,N_769,N_4056);
xnor U5147 (N_5147,N_2499,N_2176);
or U5148 (N_5148,N_4915,N_2163);
nand U5149 (N_5149,N_4049,N_1310);
xor U5150 (N_5150,N_12,N_2708);
xor U5151 (N_5151,N_3531,N_3364);
nor U5152 (N_5152,N_389,N_4703);
nor U5153 (N_5153,N_594,N_2889);
and U5154 (N_5154,N_649,N_3248);
nor U5155 (N_5155,N_268,N_4157);
and U5156 (N_5156,N_3069,N_1042);
and U5157 (N_5157,N_4983,N_634);
or U5158 (N_5158,N_4165,N_3186);
and U5159 (N_5159,N_3546,N_628);
and U5160 (N_5160,N_3679,N_3922);
or U5161 (N_5161,N_1244,N_4494);
nor U5162 (N_5162,N_3055,N_3384);
xnor U5163 (N_5163,N_1398,N_3599);
nor U5164 (N_5164,N_2881,N_4337);
or U5165 (N_5165,N_4810,N_4856);
nand U5166 (N_5166,N_4768,N_1138);
and U5167 (N_5167,N_4127,N_3465);
xor U5168 (N_5168,N_1532,N_4092);
nor U5169 (N_5169,N_1507,N_2269);
xor U5170 (N_5170,N_3704,N_4739);
nor U5171 (N_5171,N_4829,N_1562);
and U5172 (N_5172,N_1391,N_1452);
nand U5173 (N_5173,N_314,N_1873);
and U5174 (N_5174,N_921,N_3862);
xor U5175 (N_5175,N_1341,N_157);
and U5176 (N_5176,N_1395,N_807);
or U5177 (N_5177,N_2783,N_1606);
xor U5178 (N_5178,N_1543,N_4727);
and U5179 (N_5179,N_386,N_3655);
nand U5180 (N_5180,N_3349,N_2330);
or U5181 (N_5181,N_3905,N_3363);
nand U5182 (N_5182,N_4624,N_4849);
and U5183 (N_5183,N_2968,N_3075);
or U5184 (N_5184,N_4997,N_48);
nor U5185 (N_5185,N_1570,N_188);
nor U5186 (N_5186,N_2209,N_506);
and U5187 (N_5187,N_2745,N_1949);
xnor U5188 (N_5188,N_2194,N_4658);
nand U5189 (N_5189,N_1598,N_3498);
and U5190 (N_5190,N_2165,N_3111);
or U5191 (N_5191,N_3220,N_3446);
nor U5192 (N_5192,N_1920,N_3027);
or U5193 (N_5193,N_4508,N_1216);
nor U5194 (N_5194,N_352,N_2811);
nor U5195 (N_5195,N_951,N_876);
and U5196 (N_5196,N_840,N_4622);
nor U5197 (N_5197,N_2955,N_4991);
nor U5198 (N_5198,N_1793,N_3509);
or U5199 (N_5199,N_3755,N_4053);
or U5200 (N_5200,N_4126,N_426);
or U5201 (N_5201,N_3386,N_1228);
and U5202 (N_5202,N_1298,N_1899);
xnor U5203 (N_5203,N_3089,N_4423);
xnor U5204 (N_5204,N_2696,N_328);
nor U5205 (N_5205,N_2644,N_980);
xor U5206 (N_5206,N_1139,N_757);
and U5207 (N_5207,N_4599,N_1767);
xnor U5208 (N_5208,N_4945,N_86);
and U5209 (N_5209,N_89,N_4141);
nor U5210 (N_5210,N_2767,N_2903);
nor U5211 (N_5211,N_3304,N_1963);
nor U5212 (N_5212,N_4100,N_401);
nor U5213 (N_5213,N_1280,N_3985);
and U5214 (N_5214,N_3473,N_2030);
or U5215 (N_5215,N_2995,N_98);
or U5216 (N_5216,N_992,N_4512);
nor U5217 (N_5217,N_1923,N_4851);
nand U5218 (N_5218,N_4524,N_2346);
xnor U5219 (N_5219,N_4963,N_2661);
xnor U5220 (N_5220,N_2162,N_1867);
xor U5221 (N_5221,N_4247,N_2508);
or U5222 (N_5222,N_81,N_3439);
and U5223 (N_5223,N_3382,N_2815);
and U5224 (N_5224,N_3099,N_3683);
and U5225 (N_5225,N_1799,N_2910);
and U5226 (N_5226,N_4616,N_3927);
nor U5227 (N_5227,N_563,N_1534);
and U5228 (N_5228,N_515,N_21);
nand U5229 (N_5229,N_4890,N_164);
nand U5230 (N_5230,N_614,N_1700);
nand U5231 (N_5231,N_1387,N_2700);
nor U5232 (N_5232,N_4964,N_3664);
nor U5233 (N_5233,N_0,N_4394);
nor U5234 (N_5234,N_1895,N_1750);
and U5235 (N_5235,N_3270,N_912);
nand U5236 (N_5236,N_1851,N_1429);
and U5237 (N_5237,N_738,N_4894);
nand U5238 (N_5238,N_4793,N_4885);
or U5239 (N_5239,N_42,N_144);
and U5240 (N_5240,N_817,N_2757);
xor U5241 (N_5241,N_1369,N_678);
or U5242 (N_5242,N_2630,N_1441);
or U5243 (N_5243,N_2120,N_3290);
nand U5244 (N_5244,N_2347,N_2220);
or U5245 (N_5245,N_4491,N_4802);
and U5246 (N_5246,N_4168,N_3201);
nand U5247 (N_5247,N_2985,N_323);
nor U5248 (N_5248,N_744,N_2318);
xnor U5249 (N_5249,N_3628,N_3477);
xor U5250 (N_5250,N_1205,N_15);
xor U5251 (N_5251,N_1567,N_4065);
xnor U5252 (N_5252,N_3211,N_1067);
nor U5253 (N_5253,N_3792,N_1407);
xor U5254 (N_5254,N_4880,N_4718);
or U5255 (N_5255,N_3231,N_2989);
and U5256 (N_5256,N_2270,N_382);
xnor U5257 (N_5257,N_455,N_910);
or U5258 (N_5258,N_3144,N_4611);
xor U5259 (N_5259,N_4232,N_297);
nand U5260 (N_5260,N_4471,N_1970);
nand U5261 (N_5261,N_3800,N_1684);
or U5262 (N_5262,N_849,N_1075);
nor U5263 (N_5263,N_4683,N_240);
nand U5264 (N_5264,N_1351,N_2256);
or U5265 (N_5265,N_1977,N_1227);
and U5266 (N_5266,N_2951,N_4742);
nor U5267 (N_5267,N_3360,N_707);
nor U5268 (N_5268,N_121,N_3632);
xor U5269 (N_5269,N_1497,N_2603);
nor U5270 (N_5270,N_2714,N_2566);
and U5271 (N_5271,N_4369,N_3464);
or U5272 (N_5272,N_3318,N_2876);
xnor U5273 (N_5273,N_1226,N_900);
and U5274 (N_5274,N_3773,N_3846);
nor U5275 (N_5275,N_893,N_55);
and U5276 (N_5276,N_264,N_149);
nand U5277 (N_5277,N_4198,N_1590);
or U5278 (N_5278,N_1039,N_4877);
nor U5279 (N_5279,N_122,N_1715);
or U5280 (N_5280,N_456,N_1069);
and U5281 (N_5281,N_2524,N_2663);
or U5282 (N_5282,N_4286,N_3919);
or U5283 (N_5283,N_4020,N_2486);
nor U5284 (N_5284,N_444,N_4004);
and U5285 (N_5285,N_1359,N_2410);
nand U5286 (N_5286,N_4452,N_2141);
nor U5287 (N_5287,N_289,N_886);
nand U5288 (N_5288,N_1053,N_4543);
xnor U5289 (N_5289,N_4123,N_2930);
and U5290 (N_5290,N_2958,N_3692);
or U5291 (N_5291,N_4695,N_1832);
nor U5292 (N_5292,N_3086,N_1115);
nor U5293 (N_5293,N_3423,N_4527);
xor U5294 (N_5294,N_3355,N_100);
xnor U5295 (N_5295,N_4958,N_194);
nand U5296 (N_5296,N_2128,N_101);
nand U5297 (N_5297,N_2890,N_3540);
nor U5298 (N_5298,N_4843,N_2242);
or U5299 (N_5299,N_4159,N_902);
nand U5300 (N_5300,N_2879,N_1708);
and U5301 (N_5301,N_3484,N_257);
xnor U5302 (N_5302,N_535,N_1149);
and U5303 (N_5303,N_4091,N_4928);
or U5304 (N_5304,N_3380,N_94);
or U5305 (N_5305,N_3954,N_4641);
and U5306 (N_5306,N_2752,N_4392);
nor U5307 (N_5307,N_3284,N_1637);
nand U5308 (N_5308,N_4661,N_3091);
xor U5309 (N_5309,N_4651,N_3119);
and U5310 (N_5310,N_1585,N_371);
nand U5311 (N_5311,N_2833,N_2801);
xnor U5312 (N_5312,N_2203,N_3649);
nand U5313 (N_5313,N_784,N_4256);
nor U5314 (N_5314,N_4236,N_4054);
xor U5315 (N_5315,N_1112,N_1558);
nand U5316 (N_5316,N_1299,N_2258);
or U5317 (N_5317,N_320,N_4164);
and U5318 (N_5318,N_1595,N_2212);
and U5319 (N_5319,N_3402,N_1021);
or U5320 (N_5320,N_1082,N_199);
or U5321 (N_5321,N_4119,N_3812);
nand U5322 (N_5322,N_4818,N_2402);
nor U5323 (N_5323,N_1087,N_654);
and U5324 (N_5324,N_2079,N_252);
and U5325 (N_5325,N_485,N_761);
and U5326 (N_5326,N_1026,N_1872);
nor U5327 (N_5327,N_2799,N_3994);
nand U5328 (N_5328,N_4937,N_3299);
nor U5329 (N_5329,N_4096,N_3652);
xor U5330 (N_5330,N_4441,N_4191);
and U5331 (N_5331,N_1822,N_1820);
nor U5332 (N_5332,N_4947,N_1905);
or U5333 (N_5333,N_2919,N_2505);
and U5334 (N_5334,N_613,N_3345);
xor U5335 (N_5335,N_3131,N_1326);
nor U5336 (N_5336,N_2363,N_4131);
nor U5337 (N_5337,N_3440,N_2003);
and U5338 (N_5338,N_1005,N_4528);
nand U5339 (N_5339,N_4211,N_3177);
or U5340 (N_5340,N_2215,N_570);
and U5341 (N_5341,N_2986,N_2117);
and U5342 (N_5342,N_3840,N_1857);
and U5343 (N_5343,N_2259,N_4863);
nor U5344 (N_5344,N_126,N_2448);
and U5345 (N_5345,N_1704,N_4380);
or U5346 (N_5346,N_76,N_740);
xor U5347 (N_5347,N_1992,N_2763);
and U5348 (N_5348,N_2598,N_891);
or U5349 (N_5349,N_373,N_1763);
nand U5350 (N_5350,N_332,N_2762);
xnor U5351 (N_5351,N_4653,N_4909);
nand U5352 (N_5352,N_4201,N_2734);
nor U5353 (N_5353,N_4241,N_958);
nor U5354 (N_5354,N_1916,N_4035);
and U5355 (N_5355,N_4032,N_1460);
nor U5356 (N_5356,N_304,N_4308);
nand U5357 (N_5357,N_1667,N_3527);
xor U5358 (N_5358,N_1661,N_138);
and U5359 (N_5359,N_2244,N_4602);
nor U5360 (N_5360,N_3145,N_2321);
nor U5361 (N_5361,N_1756,N_4722);
nor U5362 (N_5362,N_3584,N_2130);
or U5363 (N_5363,N_3287,N_3148);
or U5364 (N_5364,N_4563,N_2357);
nor U5365 (N_5365,N_3114,N_4350);
and U5366 (N_5366,N_700,N_96);
or U5367 (N_5367,N_2011,N_2817);
nor U5368 (N_5368,N_4996,N_2314);
or U5369 (N_5369,N_3990,N_2138);
xnor U5370 (N_5370,N_4105,N_3230);
nand U5371 (N_5371,N_4064,N_2257);
nand U5372 (N_5372,N_3497,N_491);
nand U5373 (N_5373,N_2681,N_1631);
and U5374 (N_5374,N_1827,N_1223);
nand U5375 (N_5375,N_2015,N_4177);
and U5376 (N_5376,N_3969,N_3513);
or U5377 (N_5377,N_1199,N_688);
nor U5378 (N_5378,N_1498,N_2249);
xnor U5379 (N_5379,N_1331,N_2529);
nand U5380 (N_5380,N_2892,N_1225);
xnor U5381 (N_5381,N_3639,N_3740);
or U5382 (N_5382,N_1523,N_940);
nand U5383 (N_5383,N_1050,N_2795);
nand U5384 (N_5384,N_4190,N_1493);
or U5385 (N_5385,N_3499,N_1769);
xor U5386 (N_5386,N_2587,N_1980);
nand U5387 (N_5387,N_3657,N_1133);
nor U5388 (N_5388,N_4342,N_861);
nand U5389 (N_5389,N_3372,N_887);
and U5390 (N_5390,N_3835,N_2429);
nor U5391 (N_5391,N_1613,N_301);
xor U5392 (N_5392,N_2994,N_3357);
and U5393 (N_5393,N_4948,N_2362);
and U5394 (N_5394,N_697,N_3039);
and U5395 (N_5395,N_3154,N_826);
or U5396 (N_5396,N_4574,N_3925);
xor U5397 (N_5397,N_4440,N_3173);
nand U5398 (N_5398,N_225,N_3889);
nor U5399 (N_5399,N_1200,N_4869);
and U5400 (N_5400,N_1488,N_2210);
or U5401 (N_5401,N_90,N_1698);
nand U5402 (N_5402,N_2020,N_1400);
xnor U5403 (N_5403,N_2248,N_528);
nor U5404 (N_5404,N_3648,N_3613);
nand U5405 (N_5405,N_3523,N_1685);
nor U5406 (N_5406,N_993,N_4531);
nand U5407 (N_5407,N_1903,N_2013);
xor U5408 (N_5408,N_1323,N_265);
xnor U5409 (N_5409,N_2888,N_1235);
and U5410 (N_5410,N_4990,N_4390);
nor U5411 (N_5411,N_484,N_556);
or U5412 (N_5412,N_1858,N_2731);
or U5413 (N_5413,N_3271,N_2711);
and U5414 (N_5414,N_3968,N_181);
or U5415 (N_5415,N_8,N_246);
xor U5416 (N_5416,N_146,N_1538);
nand U5417 (N_5417,N_1882,N_119);
nor U5418 (N_5418,N_1571,N_168);
and U5419 (N_5419,N_2620,N_2206);
and U5420 (N_5420,N_4940,N_1390);
xnor U5421 (N_5421,N_877,N_4373);
nor U5422 (N_5422,N_2073,N_2147);
nand U5423 (N_5423,N_3795,N_3064);
nor U5424 (N_5424,N_2452,N_3614);
nand U5425 (N_5425,N_2975,N_279);
and U5426 (N_5426,N_1514,N_1104);
and U5427 (N_5427,N_2525,N_213);
nor U5428 (N_5428,N_2843,N_3771);
nor U5429 (N_5429,N_558,N_3658);
xor U5430 (N_5430,N_516,N_4405);
nor U5431 (N_5431,N_1031,N_660);
xnor U5432 (N_5432,N_3597,N_2864);
nand U5433 (N_5433,N_1183,N_3623);
or U5434 (N_5434,N_1918,N_3722);
and U5435 (N_5435,N_4741,N_50);
xnor U5436 (N_5436,N_1761,N_1754);
and U5437 (N_5437,N_1783,N_3899);
nor U5438 (N_5438,N_116,N_1003);
xor U5439 (N_5439,N_4411,N_3320);
or U5440 (N_5440,N_1328,N_1213);
nand U5441 (N_5441,N_1000,N_2590);
nand U5442 (N_5442,N_552,N_4181);
and U5443 (N_5443,N_2649,N_1935);
and U5444 (N_5444,N_4956,N_3831);
and U5445 (N_5445,N_1164,N_4867);
nor U5446 (N_5446,N_4566,N_1239);
nand U5447 (N_5447,N_2113,N_1165);
or U5448 (N_5448,N_4263,N_2633);
or U5449 (N_5449,N_61,N_1691);
or U5450 (N_5450,N_3167,N_2940);
nand U5451 (N_5451,N_1655,N_249);
xnor U5452 (N_5452,N_3070,N_3003);
nor U5453 (N_5453,N_276,N_834);
nor U5454 (N_5454,N_1871,N_2901);
nor U5455 (N_5455,N_2650,N_1615);
and U5456 (N_5456,N_2948,N_593);
xnor U5457 (N_5457,N_4738,N_3431);
nand U5458 (N_5458,N_2058,N_2907);
nor U5459 (N_5459,N_3108,N_3785);
and U5460 (N_5460,N_3913,N_2884);
nor U5461 (N_5461,N_4640,N_2);
and U5462 (N_5462,N_448,N_495);
or U5463 (N_5463,N_2271,N_2846);
xor U5464 (N_5464,N_2076,N_2159);
nand U5465 (N_5465,N_3480,N_830);
nor U5466 (N_5466,N_1772,N_2828);
nor U5467 (N_5467,N_2476,N_2472);
nor U5468 (N_5468,N_565,N_610);
and U5469 (N_5469,N_5,N_605);
and U5470 (N_5470,N_487,N_4774);
nand U5471 (N_5471,N_3383,N_211);
nand U5472 (N_5472,N_4366,N_1641);
or U5473 (N_5473,N_2569,N_3434);
or U5474 (N_5474,N_4914,N_1713);
or U5475 (N_5475,N_3716,N_1196);
xor U5476 (N_5476,N_997,N_2132);
and U5477 (N_5477,N_4755,N_1791);
nor U5478 (N_5478,N_2722,N_4179);
xnor U5479 (N_5479,N_4214,N_3482);
and U5480 (N_5480,N_2422,N_1581);
nor U5481 (N_5481,N_801,N_4475);
nor U5482 (N_5482,N_4057,N_1120);
xor U5483 (N_5483,N_935,N_3236);
xnor U5484 (N_5484,N_1161,N_1975);
xor U5485 (N_5485,N_2554,N_846);
xnor U5486 (N_5486,N_968,N_2759);
nor U5487 (N_5487,N_160,N_1130);
and U5488 (N_5488,N_4459,N_2139);
nor U5489 (N_5489,N_437,N_2671);
nor U5490 (N_5490,N_4519,N_4);
xor U5491 (N_5491,N_1719,N_2909);
xor U5492 (N_5492,N_1801,N_3146);
nand U5493 (N_5493,N_638,N_3801);
nand U5494 (N_5494,N_83,N_4169);
nand U5495 (N_5495,N_3082,N_4955);
xnor U5496 (N_5496,N_2241,N_3200);
xnor U5497 (N_5497,N_3682,N_4876);
xor U5498 (N_5498,N_4857,N_2738);
or U5499 (N_5499,N_991,N_4708);
nor U5500 (N_5500,N_2385,N_1405);
and U5501 (N_5501,N_2285,N_4844);
nor U5502 (N_5502,N_2170,N_2538);
or U5503 (N_5503,N_2035,N_4912);
or U5504 (N_5504,N_1218,N_1547);
xor U5505 (N_5505,N_3912,N_1678);
xnor U5506 (N_5506,N_2666,N_1663);
xnor U5507 (N_5507,N_3742,N_3926);
xor U5508 (N_5508,N_3894,N_2871);
or U5509 (N_5509,N_2418,N_3883);
xnor U5510 (N_5510,N_496,N_1505);
xor U5511 (N_5511,N_3595,N_4024);
nor U5512 (N_5512,N_1086,N_4553);
and U5513 (N_5513,N_177,N_2097);
nand U5514 (N_5514,N_4172,N_870);
xnor U5515 (N_5515,N_1270,N_123);
xnor U5516 (N_5516,N_489,N_3958);
nor U5517 (N_5517,N_4546,N_686);
or U5518 (N_5518,N_3467,N_2024);
and U5519 (N_5519,N_1106,N_325);
nand U5520 (N_5520,N_4590,N_350);
nor U5521 (N_5521,N_2949,N_4754);
or U5522 (N_5522,N_3694,N_221);
xnor U5523 (N_5523,N_4677,N_4745);
nor U5524 (N_5524,N_1784,N_2420);
nand U5525 (N_5525,N_278,N_4597);
xnor U5526 (N_5526,N_4446,N_3294);
or U5527 (N_5527,N_1459,N_3541);
nor U5528 (N_5528,N_3256,N_2517);
nor U5529 (N_5529,N_2845,N_778);
and U5530 (N_5530,N_2092,N_1512);
nand U5531 (N_5531,N_362,N_1922);
xor U5532 (N_5532,N_2557,N_1413);
and U5533 (N_5533,N_4561,N_693);
or U5534 (N_5534,N_2012,N_675);
or U5535 (N_5535,N_2697,N_2198);
nor U5536 (N_5536,N_1645,N_4686);
or U5537 (N_5537,N_324,N_3807);
or U5538 (N_5538,N_1914,N_3435);
or U5539 (N_5539,N_2576,N_667);
nor U5540 (N_5540,N_3367,N_994);
or U5541 (N_5541,N_3319,N_1506);
and U5542 (N_5542,N_3538,N_2856);
nor U5543 (N_5543,N_4359,N_2056);
nand U5544 (N_5544,N_4815,N_2389);
nand U5545 (N_5545,N_2150,N_4505);
and U5546 (N_5546,N_3330,N_1257);
nand U5547 (N_5547,N_4669,N_1765);
xor U5548 (N_5548,N_4162,N_1579);
or U5549 (N_5549,N_3414,N_545);
nand U5550 (N_5550,N_4432,N_258);
nand U5551 (N_5551,N_1024,N_2808);
nor U5552 (N_5552,N_2126,N_3617);
and U5553 (N_5553,N_3077,N_192);
xnor U5554 (N_5554,N_2497,N_4438);
nor U5555 (N_5555,N_4549,N_854);
or U5556 (N_5556,N_2217,N_4648);
nand U5557 (N_5557,N_31,N_3693);
nand U5558 (N_5558,N_3180,N_3504);
xnor U5559 (N_5559,N_1088,N_1399);
nand U5560 (N_5560,N_3936,N_909);
nor U5561 (N_5561,N_2374,N_2513);
or U5562 (N_5562,N_4697,N_2143);
nor U5563 (N_5563,N_3456,N_2514);
or U5564 (N_5564,N_3908,N_3128);
nand U5565 (N_5565,N_1156,N_471);
xor U5566 (N_5566,N_3873,N_66);
nor U5567 (N_5567,N_2054,N_38);
xnor U5568 (N_5568,N_2245,N_212);
nand U5569 (N_5569,N_2642,N_4231);
nand U5570 (N_5570,N_247,N_3754);
nor U5571 (N_5571,N_2996,N_4367);
nor U5572 (N_5572,N_2036,N_4804);
nand U5573 (N_5573,N_1648,N_2834);
nor U5574 (N_5574,N_1710,N_4479);
xor U5575 (N_5575,N_3646,N_2192);
nor U5576 (N_5576,N_2118,N_4610);
or U5577 (N_5577,N_715,N_1484);
and U5578 (N_5578,N_3620,N_1446);
or U5579 (N_5579,N_3861,N_2100);
nor U5580 (N_5580,N_4580,N_939);
and U5581 (N_5581,N_2792,N_4782);
xnor U5582 (N_5582,N_1275,N_4865);
nor U5583 (N_5583,N_622,N_3223);
xnor U5584 (N_5584,N_4923,N_4671);
xnor U5585 (N_5585,N_640,N_3733);
nand U5586 (N_5586,N_1313,N_337);
xnor U5587 (N_5587,N_4633,N_1815);
nor U5588 (N_5588,N_929,N_3732);
nor U5589 (N_5589,N_209,N_1508);
or U5590 (N_5590,N_214,N_4552);
xnor U5591 (N_5591,N_1526,N_4679);
xor U5592 (N_5592,N_1816,N_3668);
or U5593 (N_5593,N_3660,N_403);
nor U5594 (N_5594,N_1861,N_4250);
nand U5595 (N_5595,N_2766,N_3225);
or U5596 (N_5596,N_3176,N_2183);
or U5597 (N_5597,N_4399,N_1076);
nor U5598 (N_5598,N_1690,N_3344);
or U5599 (N_5599,N_1201,N_1167);
or U5600 (N_5600,N_1015,N_4949);
or U5601 (N_5601,N_2835,N_1766);
nand U5602 (N_5602,N_3001,N_1163);
and U5603 (N_5603,N_1074,N_3457);
xor U5604 (N_5604,N_340,N_1083);
xnor U5605 (N_5605,N_2461,N_3579);
and U5606 (N_5606,N_4501,N_4737);
xnor U5607 (N_5607,N_4137,N_34);
or U5608 (N_5608,N_3459,N_3377);
nor U5609 (N_5609,N_9,N_2515);
xnor U5610 (N_5610,N_833,N_1960);
xnor U5611 (N_5611,N_2935,N_1185);
or U5612 (N_5612,N_4757,N_3512);
and U5613 (N_5613,N_4850,N_4267);
or U5614 (N_5614,N_1382,N_1885);
xnor U5615 (N_5615,N_2637,N_1467);
nand U5616 (N_5616,N_91,N_3891);
or U5617 (N_5617,N_3667,N_2600);
nand U5618 (N_5618,N_4726,N_4920);
nor U5619 (N_5619,N_3252,N_1560);
or U5620 (N_5620,N_1633,N_2438);
and U5621 (N_5621,N_2065,N_855);
and U5622 (N_5622,N_1073,N_1373);
and U5623 (N_5623,N_2562,N_765);
or U5624 (N_5624,N_3629,N_4285);
xnor U5625 (N_5625,N_3678,N_2479);
nand U5626 (N_5626,N_3825,N_424);
and U5627 (N_5627,N_721,N_3245);
nand U5628 (N_5628,N_3940,N_2810);
and U5629 (N_5629,N_3600,N_2482);
or U5630 (N_5630,N_922,N_2068);
and U5631 (N_5631,N_2825,N_1717);
nor U5632 (N_5632,N_2425,N_4638);
xnor U5633 (N_5633,N_3898,N_2659);
and U5634 (N_5634,N_59,N_300);
or U5635 (N_5635,N_3002,N_2741);
and U5636 (N_5636,N_3858,N_2311);
xnor U5637 (N_5637,N_2161,N_3814);
nor U5638 (N_5638,N_811,N_4764);
or U5639 (N_5639,N_2102,N_979);
nand U5640 (N_5640,N_1554,N_40);
and U5641 (N_5641,N_587,N_273);
or U5642 (N_5642,N_393,N_3103);
and U5643 (N_5643,N_142,N_3505);
nor U5644 (N_5644,N_2952,N_1397);
nor U5645 (N_5645,N_3714,N_1762);
or U5646 (N_5646,N_4893,N_103);
nor U5647 (N_5647,N_1238,N_2933);
and U5648 (N_5648,N_2614,N_2184);
xnor U5649 (N_5649,N_159,N_1170);
xor U5650 (N_5650,N_666,N_2308);
nor U5651 (N_5651,N_1921,N_4318);
xnor U5652 (N_5652,N_3552,N_235);
or U5653 (N_5653,N_2648,N_2317);
nand U5654 (N_5654,N_639,N_1951);
xnor U5655 (N_5655,N_624,N_2342);
or U5656 (N_5656,N_1521,N_2408);
and U5657 (N_5657,N_4930,N_2485);
or U5658 (N_5658,N_2096,N_2480);
nor U5659 (N_5659,N_1386,N_2280);
nor U5660 (N_5660,N_1230,N_2676);
xor U5661 (N_5661,N_223,N_1927);
or U5662 (N_5662,N_2033,N_1136);
xor U5663 (N_5663,N_271,N_1415);
xnor U5664 (N_5664,N_2310,N_815);
nand U5665 (N_5665,N_4904,N_1284);
and U5666 (N_5666,N_4756,N_3263);
or U5667 (N_5667,N_894,N_3244);
or U5668 (N_5668,N_723,N_1157);
nand U5669 (N_5669,N_1591,N_844);
or U5670 (N_5670,N_684,N_1879);
nor U5671 (N_5671,N_2939,N_3876);
or U5672 (N_5672,N_4288,N_3411);
and U5673 (N_5673,N_745,N_3331);
nor U5674 (N_5674,N_2218,N_736);
nand U5675 (N_5675,N_1711,N_2140);
and U5676 (N_5676,N_4360,N_2431);
xor U5677 (N_5677,N_2523,N_3181);
nand U5678 (N_5678,N_3938,N_4852);
or U5679 (N_5679,N_3612,N_1195);
nor U5680 (N_5680,N_1864,N_4626);
or U5681 (N_5681,N_978,N_3677);
or U5682 (N_5682,N_656,N_1819);
nor U5683 (N_5683,N_1478,N_3813);
and U5684 (N_5684,N_2225,N_185);
or U5685 (N_5685,N_4104,N_3586);
and U5686 (N_5686,N_971,N_3442);
xor U5687 (N_5687,N_2787,N_4007);
nand U5688 (N_5688,N_2507,N_4973);
or U5689 (N_5689,N_3142,N_2904);
nand U5690 (N_5690,N_3479,N_4873);
nor U5691 (N_5691,N_4345,N_1610);
nand U5692 (N_5692,N_635,N_1327);
or U5693 (N_5693,N_1312,N_4860);
and U5694 (N_5694,N_1709,N_4978);
nand U5695 (N_5695,N_2673,N_1463);
or U5696 (N_5696,N_2842,N_1414);
nor U5697 (N_5697,N_4710,N_4061);
nor U5698 (N_5698,N_795,N_454);
or U5699 (N_5699,N_1853,N_2167);
nor U5700 (N_5700,N_1274,N_3118);
xor U5701 (N_5701,N_1666,N_4664);
nand U5702 (N_5702,N_1950,N_366);
and U5703 (N_5703,N_2123,N_1271);
xnor U5704 (N_5704,N_3427,N_2819);
nand U5705 (N_5705,N_158,N_2401);
or U5706 (N_5706,N_4233,N_3596);
nand U5707 (N_5707,N_2293,N_1742);
or U5708 (N_5708,N_1811,N_425);
or U5709 (N_5709,N_4705,N_1564);
nand U5710 (N_5710,N_3162,N_322);
nor U5711 (N_5711,N_3291,N_3671);
or U5712 (N_5712,N_1776,N_4066);
nor U5713 (N_5713,N_2247,N_4496);
nand U5714 (N_5714,N_3511,N_4146);
or U5715 (N_5715,N_2717,N_4070);
and U5716 (N_5716,N_1942,N_644);
and U5717 (N_5717,N_49,N_3347);
nand U5718 (N_5718,N_2530,N_2124);
or U5719 (N_5719,N_4344,N_241);
xnor U5720 (N_5720,N_2227,N_2037);
nand U5721 (N_5721,N_3283,N_3235);
xor U5722 (N_5722,N_2473,N_4328);
xnor U5723 (N_5723,N_1556,N_3904);
xor U5724 (N_5724,N_4696,N_3574);
nand U5725 (N_5725,N_2657,N_1652);
xor U5726 (N_5726,N_1596,N_69);
or U5727 (N_5727,N_3500,N_4334);
nor U5728 (N_5728,N_2038,N_4167);
nand U5729 (N_5729,N_4352,N_4921);
xnor U5730 (N_5730,N_1696,N_129);
nand U5731 (N_5731,N_1679,N_4777);
or U5732 (N_5732,N_1465,N_2803);
and U5733 (N_5733,N_1826,N_1281);
or U5734 (N_5734,N_1097,N_2334);
nor U5735 (N_5735,N_2426,N_4965);
xor U5736 (N_5736,N_4116,N_3400);
or U5737 (N_5737,N_137,N_2387);
and U5738 (N_5738,N_2214,N_1629);
or U5739 (N_5739,N_1798,N_3009);
xor U5740 (N_5740,N_1148,N_3713);
or U5741 (N_5741,N_838,N_14);
nor U5742 (N_5742,N_2135,N_3381);
nor U5743 (N_5743,N_1214,N_1055);
nor U5744 (N_5744,N_413,N_1152);
xnor U5745 (N_5745,N_493,N_2539);
nand U5746 (N_5746,N_1525,N_3603);
nand U5747 (N_5747,N_3685,N_4003);
nor U5748 (N_5748,N_3955,N_2827);
xnor U5749 (N_5749,N_269,N_357);
nor U5750 (N_5750,N_2965,N_2800);
nor U5751 (N_5751,N_1981,N_423);
xor U5752 (N_5752,N_4969,N_3254);
nand U5753 (N_5753,N_1744,N_3329);
and U5754 (N_5754,N_1034,N_3952);
and U5755 (N_5755,N_2521,N_4470);
xnor U5756 (N_5756,N_2458,N_2193);
nor U5757 (N_5757,N_4194,N_4050);
and U5758 (N_5758,N_4284,N_3419);
or U5759 (N_5759,N_3798,N_1974);
and U5760 (N_5760,N_4684,N_4577);
nor U5761 (N_5761,N_4031,N_2484);
nor U5762 (N_5762,N_3971,N_3247);
or U5763 (N_5763,N_759,N_2303);
and U5764 (N_5764,N_938,N_4277);
xor U5765 (N_5765,N_691,N_2960);
and U5766 (N_5766,N_2083,N_4227);
and U5767 (N_5767,N_945,N_1670);
nand U5768 (N_5768,N_4237,N_2339);
nand U5769 (N_5769,N_1499,N_1866);
nor U5770 (N_5770,N_1419,N_2726);
xnor U5771 (N_5771,N_1366,N_2101);
nor U5772 (N_5772,N_1256,N_4725);
or U5773 (N_5773,N_2586,N_4193);
and U5774 (N_5774,N_3643,N_1600);
nor U5775 (N_5775,N_3915,N_4205);
or U5776 (N_5776,N_2338,N_3516);
xor U5777 (N_5777,N_1266,N_111);
nand U5778 (N_5778,N_2207,N_577);
nand U5779 (N_5779,N_32,N_2691);
xnor U5780 (N_5780,N_4176,N_2577);
xor U5781 (N_5781,N_57,N_2231);
nand U5782 (N_5782,N_4207,N_380);
nor U5783 (N_5783,N_1603,N_2629);
xor U5784 (N_5784,N_4403,N_1030);
xnor U5785 (N_5785,N_2632,N_3534);
and U5786 (N_5786,N_1665,N_3351);
nor U5787 (N_5787,N_2836,N_2850);
nand U5788 (N_5788,N_1743,N_714);
nor U5789 (N_5789,N_1236,N_396);
and U5790 (N_5790,N_4259,N_4370);
nor U5791 (N_5791,N_4296,N_974);
xor U5792 (N_5792,N_763,N_4079);
nand U5793 (N_5793,N_2913,N_943);
and U5794 (N_5794,N_333,N_4206);
or U5795 (N_5795,N_1045,N_1731);
xnor U5796 (N_5796,N_3551,N_117);
or U5797 (N_5797,N_118,N_3729);
and U5798 (N_5798,N_4750,N_1456);
xnor U5799 (N_5799,N_3397,N_4809);
and U5800 (N_5800,N_97,N_155);
and U5801 (N_5801,N_1318,N_2496);
nor U5802 (N_5802,N_4827,N_1723);
or U5803 (N_5803,N_869,N_1640);
and U5804 (N_5804,N_2639,N_955);
nand U5805 (N_5805,N_627,N_1939);
or U5806 (N_5806,N_2551,N_3452);
nor U5807 (N_5807,N_1989,N_2307);
xnor U5808 (N_5808,N_3886,N_4871);
or U5809 (N_5809,N_93,N_2646);
or U5810 (N_5810,N_224,N_1158);
nor U5811 (N_5811,N_3956,N_3751);
nor U5812 (N_5812,N_4321,N_937);
or U5813 (N_5813,N_3703,N_1889);
or U5814 (N_5814,N_4451,N_3206);
nand U5815 (N_5815,N_2383,N_4115);
nand U5816 (N_5816,N_2263,N_925);
or U5817 (N_5817,N_2894,N_4587);
nand U5818 (N_5818,N_692,N_1422);
nand U5819 (N_5819,N_3897,N_3097);
nand U5820 (N_5820,N_1909,N_4239);
nor U5821 (N_5821,N_319,N_3253);
nand U5822 (N_5822,N_4011,N_439);
nand U5823 (N_5823,N_3622,N_1707);
nor U5824 (N_5824,N_791,N_538);
nand U5825 (N_5825,N_1893,N_3393);
and U5826 (N_5826,N_355,N_3917);
nor U5827 (N_5827,N_3450,N_3443);
or U5828 (N_5828,N_2709,N_1278);
or U5829 (N_5829,N_2488,N_1081);
nor U5830 (N_5830,N_3816,N_4642);
and U5831 (N_5831,N_753,N_970);
nand U5832 (N_5832,N_4382,N_2857);
and U5833 (N_5833,N_237,N_88);
nor U5834 (N_5834,N_2744,N_2274);
xor U5835 (N_5835,N_4970,N_2070);
or U5836 (N_5836,N_932,N_2179);
nor U5837 (N_5837,N_3420,N_571);
xnor U5838 (N_5838,N_2392,N_1125);
nor U5839 (N_5839,N_4270,N_2540);
and U5840 (N_5840,N_2961,N_1878);
nand U5841 (N_5841,N_4224,N_381);
nor U5842 (N_5842,N_4314,N_3687);
xor U5843 (N_5843,N_783,N_4634);
and U5844 (N_5844,N_2254,N_3033);
or U5845 (N_5845,N_1211,N_395);
nand U5846 (N_5846,N_2371,N_4882);
or U5847 (N_5847,N_1355,N_3741);
and U5848 (N_5848,N_3503,N_4346);
nand U5849 (N_5849,N_2477,N_2765);
nor U5850 (N_5850,N_1314,N_4666);
and U5851 (N_5851,N_598,N_2112);
or U5852 (N_5852,N_4048,N_3080);
or U5853 (N_5853,N_1008,N_702);
or U5854 (N_5854,N_3185,N_3918);
nand U5855 (N_5855,N_2423,N_3633);
or U5856 (N_5856,N_904,N_709);
xnor U5857 (N_5857,N_4569,N_3265);
and U5858 (N_5858,N_2283,N_4763);
or U5859 (N_5859,N_2186,N_1210);
nor U5860 (N_5860,N_825,N_4200);
or U5861 (N_5861,N_4173,N_3977);
xor U5862 (N_5862,N_1113,N_3013);
nand U5863 (N_5863,N_65,N_3460);
nor U5864 (N_5864,N_2559,N_596);
or U5865 (N_5865,N_478,N_776);
or U5866 (N_5866,N_4082,N_2773);
xor U5867 (N_5867,N_287,N_3406);
nand U5868 (N_5868,N_1378,N_4655);
nor U5869 (N_5869,N_842,N_4875);
or U5870 (N_5870,N_1969,N_1184);
xor U5871 (N_5871,N_500,N_3618);
nand U5872 (N_5872,N_3429,N_204);
or U5873 (N_5873,N_2204,N_2638);
or U5874 (N_5874,N_2906,N_4223);
xnor U5875 (N_5875,N_2737,N_226);
nor U5876 (N_5876,N_942,N_1502);
nand U5877 (N_5877,N_1282,N_4150);
or U5878 (N_5878,N_3902,N_892);
or U5879 (N_5879,N_3259,N_4838);
nand U5880 (N_5880,N_1997,N_3354);
nand U5881 (N_5881,N_1071,N_1589);
nor U5882 (N_5882,N_3988,N_1431);
and U5883 (N_5883,N_2886,N_1495);
nor U5884 (N_5884,N_569,N_1643);
nand U5885 (N_5885,N_2052,N_2273);
or U5886 (N_5886,N_4588,N_1194);
nor U5887 (N_5887,N_263,N_4391);
xnor U5888 (N_5888,N_712,N_1852);
and U5889 (N_5889,N_2352,N_1123);
nand U5890 (N_5890,N_800,N_1965);
or U5891 (N_5891,N_1423,N_1427);
nand U5892 (N_5892,N_3237,N_1470);
or U5893 (N_5893,N_3489,N_4951);
xnor U5894 (N_5894,N_1605,N_4926);
nand U5895 (N_5895,N_3983,N_2976);
and U5896 (N_5896,N_2173,N_24);
xnor U5897 (N_5897,N_1455,N_881);
nor U5898 (N_5898,N_474,N_3789);
or U5899 (N_5899,N_244,N_4545);
xor U5900 (N_5900,N_1982,N_54);
and U5901 (N_5901,N_3656,N_312);
or U5902 (N_5902,N_1741,N_3634);
or U5903 (N_5903,N_2158,N_2885);
nor U5904 (N_5904,N_4585,N_1430);
nand U5905 (N_5905,N_1542,N_798);
nor U5906 (N_5906,N_2855,N_1790);
nand U5907 (N_5907,N_39,N_4636);
nand U5908 (N_5908,N_1734,N_1424);
or U5909 (N_5909,N_523,N_1785);
and U5910 (N_5910,N_3735,N_2812);
xor U5911 (N_5911,N_1865,N_756);
and U5912 (N_5912,N_2282,N_2243);
nor U5913 (N_5913,N_4047,N_2434);
nor U5914 (N_5914,N_4086,N_37);
xor U5915 (N_5915,N_2838,N_3031);
and U5916 (N_5916,N_2937,N_989);
nor U5917 (N_5917,N_3853,N_4784);
and U5918 (N_5918,N_459,N_2897);
nor U5919 (N_5919,N_10,N_2095);
nor U5920 (N_5920,N_1316,N_303);
and U5921 (N_5921,N_3208,N_4258);
and U5922 (N_5922,N_792,N_1066);
xnor U5923 (N_5923,N_134,N_2382);
xnor U5924 (N_5924,N_4591,N_4175);
xnor U5925 (N_5925,N_670,N_705);
nand U5926 (N_5926,N_4808,N_2626);
nor U5927 (N_5927,N_4845,N_4045);
xor U5928 (N_5928,N_2927,N_1340);
nor U5929 (N_5929,N_4509,N_3746);
nor U5930 (N_5930,N_2349,N_4794);
xnor U5931 (N_5931,N_4160,N_995);
xnor U5932 (N_5932,N_1445,N_431);
xor U5933 (N_5933,N_4650,N_944);
xnor U5934 (N_5934,N_3453,N_4823);
and U5935 (N_5935,N_2451,N_875);
xnor U5936 (N_5936,N_3192,N_2983);
or U5937 (N_5937,N_760,N_2463);
or U5938 (N_5938,N_3666,N_726);
nor U5939 (N_5939,N_4523,N_4866);
or U5940 (N_5940,N_3818,N_2615);
nor U5941 (N_5941,N_2878,N_1796);
nor U5942 (N_5942,N_1721,N_4424);
and U5943 (N_5943,N_3698,N_696);
xor U5944 (N_5944,N_3852,N_3257);
nor U5945 (N_5945,N_3110,N_3827);
and U5946 (N_5946,N_1006,N_1285);
xor U5947 (N_5947,N_2848,N_449);
xnor U5948 (N_5948,N_766,N_4526);
or U5949 (N_5949,N_3760,N_4707);
and U5950 (N_5950,N_1817,N_3823);
nand U5951 (N_5951,N_599,N_1561);
or U5952 (N_5952,N_4723,N_2545);
nand U5953 (N_5953,N_3398,N_2617);
or U5954 (N_5954,N_3582,N_4811);
nor U5955 (N_5955,N_983,N_934);
nand U5956 (N_5956,N_2373,N_2475);
and U5957 (N_5957,N_3310,N_2761);
and U5958 (N_5958,N_4628,N_4002);
and U5959 (N_5959,N_283,N_1855);
nand U5960 (N_5960,N_2656,N_3975);
or U5961 (N_5961,N_3553,N_4515);
or U5962 (N_5962,N_2026,N_1860);
nand U5963 (N_5963,N_2287,N_433);
and U5964 (N_5964,N_2427,N_3630);
or U5965 (N_5965,N_4068,N_907);
xnor U5966 (N_5966,N_4307,N_3521);
nand U5967 (N_5967,N_3112,N_1911);
nor U5968 (N_5968,N_3847,N_4998);
nor U5969 (N_5969,N_4299,N_3416);
or U5970 (N_5970,N_928,N_1092);
and U5971 (N_5971,N_1565,N_3478);
or U5972 (N_5972,N_4499,N_680);
nand U5973 (N_5973,N_4465,N_3215);
xnor U5974 (N_5974,N_4230,N_4798);
nand U5975 (N_5975,N_183,N_3998);
and U5976 (N_5976,N_3526,N_4306);
and U5977 (N_5977,N_3981,N_2221);
and U5978 (N_5978,N_1411,N_748);
nor U5979 (N_5979,N_1563,N_3624);
nand U5980 (N_5980,N_2921,N_3924);
nand U5981 (N_5981,N_1098,N_1372);
xor U5982 (N_5982,N_2865,N_1335);
or U5983 (N_5983,N_1160,N_3261);
and U5984 (N_5984,N_4789,N_1971);
xor U5985 (N_5985,N_486,N_501);
nand U5986 (N_5986,N_427,N_3076);
nand U5987 (N_5987,N_4833,N_4946);
or U5988 (N_5988,N_1056,N_579);
nor U5989 (N_5989,N_4027,N_4529);
xnor U5990 (N_5990,N_3626,N_631);
or U5991 (N_5991,N_2086,N_1300);
or U5992 (N_5992,N_2350,N_2232);
and U5993 (N_5993,N_4257,N_3387);
xnor U5994 (N_5994,N_2359,N_578);
nand U5995 (N_5995,N_3428,N_1986);
and U5996 (N_5996,N_2622,N_141);
or U5997 (N_5997,N_4396,N_4058);
nor U5998 (N_5998,N_3696,N_2388);
xnor U5999 (N_5999,N_4030,N_3931);
nor U6000 (N_6000,N_1653,N_554);
and U6001 (N_6001,N_2665,N_3147);
and U6002 (N_6002,N_3020,N_3501);
nor U6003 (N_6003,N_3421,N_2987);
xnor U6004 (N_6004,N_1469,N_4217);
and U6005 (N_6005,N_3280,N_4542);
nand U6006 (N_6006,N_4556,N_483);
or U6007 (N_6007,N_2478,N_1028);
nand U6008 (N_6008,N_2367,N_3188);
nor U6009 (N_6009,N_1191,N_2157);
and U6010 (N_6010,N_3556,N_1973);
or U6011 (N_6011,N_4073,N_3392);
and U6012 (N_6012,N_2246,N_2252);
or U6013 (N_6013,N_2670,N_1812);
or U6014 (N_6014,N_41,N_4118);
and U6015 (N_6015,N_3779,N_4460);
and U6016 (N_6016,N_277,N_2730);
or U6017 (N_6017,N_1259,N_282);
xor U6018 (N_6018,N_176,N_1597);
or U6019 (N_6019,N_777,N_182);
xnor U6020 (N_6020,N_901,N_3153);
nand U6021 (N_6021,N_4435,N_251);
nand U6022 (N_6022,N_2290,N_3018);
xnor U6023 (N_6023,N_4128,N_1375);
xor U6024 (N_6024,N_4426,N_551);
nor U6025 (N_6025,N_2943,N_2916);
and U6026 (N_6026,N_284,N_586);
xnor U6027 (N_6027,N_1254,N_908);
and U6028 (N_6028,N_821,N_1660);
nand U6029 (N_6029,N_1288,N_1630);
and U6030 (N_6030,N_370,N_3418);
nor U6031 (N_6031,N_3833,N_4620);
nor U6032 (N_6032,N_1494,N_3469);
nand U6033 (N_6033,N_1434,N_292);
nor U6034 (N_6034,N_4693,N_1192);
nand U6035 (N_6035,N_215,N_636);
or U6036 (N_6036,N_3702,N_293);
or U6037 (N_6037,N_4576,N_1588);
or U6038 (N_6038,N_336,N_4606);
or U6039 (N_6039,N_447,N_1129);
nand U6040 (N_6040,N_3717,N_4878);
nand U6041 (N_6041,N_2771,N_2874);
and U6042 (N_6042,N_1813,N_4575);
or U6043 (N_6043,N_3794,N_581);
or U6044 (N_6044,N_4153,N_2583);
nor U6045 (N_6045,N_451,N_4338);
xnor U6046 (N_6046,N_3550,N_1077);
xor U6047 (N_6047,N_3745,N_1870);
xnor U6048 (N_6048,N_3216,N_2770);
xor U6049 (N_6049,N_2419,N_518);
xor U6050 (N_6050,N_2802,N_4687);
xnor U6051 (N_6051,N_2168,N_2699);
nand U6052 (N_6052,N_4266,N_1492);
nand U6053 (N_6053,N_2667,N_3580);
or U6054 (N_6054,N_1956,N_4907);
or U6055 (N_6055,N_2612,N_919);
nand U6056 (N_6056,N_3545,N_866);
and U6057 (N_6057,N_2146,N_1322);
or U6058 (N_6058,N_1178,N_3374);
or U6059 (N_6059,N_2764,N_1023);
xor U6060 (N_6060,N_2361,N_4961);
or U6061 (N_6061,N_4111,N_773);
and U6062 (N_6062,N_1656,N_4467);
nor U6063 (N_6063,N_4076,N_2153);
or U6064 (N_6064,N_2635,N_1229);
nand U6065 (N_6065,N_3736,N_2145);
xor U6066 (N_6066,N_1198,N_422);
and U6067 (N_6067,N_1029,N_1025);
xnor U6068 (N_6068,N_4180,N_4151);
nand U6069 (N_6069,N_1311,N_743);
or U6070 (N_6070,N_1732,N_298);
or U6071 (N_6071,N_2449,N_3023);
and U6072 (N_6072,N_2440,N_4393);
xnor U6073 (N_6073,N_2658,N_3616);
and U6074 (N_6074,N_3838,N_3910);
nor U6075 (N_6075,N_2018,N_3549);
or U6076 (N_6076,N_3262,N_4594);
nand U6077 (N_6077,N_1068,N_562);
or U6078 (N_6078,N_4495,N_2820);
nand U6079 (N_6079,N_804,N_2702);
or U6080 (N_6080,N_256,N_4202);
nor U6081 (N_6081,N_1408,N_4999);
nand U6082 (N_6082,N_4155,N_3605);
or U6083 (N_6083,N_853,N_4572);
nor U6084 (N_6084,N_540,N_16);
and U6085 (N_6085,N_3766,N_3029);
nor U6086 (N_6086,N_2946,N_290);
nand U6087 (N_6087,N_4101,N_1084);
nor U6088 (N_6088,N_1242,N_1150);
nand U6089 (N_6089,N_1329,N_4281);
or U6090 (N_6090,N_1448,N_1231);
xor U6091 (N_6091,N_2182,N_4174);
or U6092 (N_6092,N_4942,N_3944);
xor U6093 (N_6093,N_3749,N_3036);
or U6094 (N_6094,N_3026,N_1246);
or U6095 (N_6095,N_2432,N_1622);
nor U6096 (N_6096,N_2160,N_310);
nand U6097 (N_6097,N_1180,N_2674);
and U6098 (N_6098,N_1553,N_508);
nor U6099 (N_6099,N_3753,N_4824);
or U6100 (N_6100,N_4825,N_1007);
nand U6101 (N_6101,N_1122,N_1384);
nand U6102 (N_6102,N_4746,N_331);
or U6103 (N_6103,N_3471,N_1539);
and U6104 (N_6104,N_3043,N_411);
xnor U6105 (N_6105,N_1241,N_2326);
or U6106 (N_6106,N_1304,N_3570);
or U6107 (N_6107,N_2584,N_1888);
nand U6108 (N_6108,N_1043,N_3034);
and U6109 (N_6109,N_4853,N_3061);
or U6110 (N_6110,N_4733,N_1037);
nor U6111 (N_6111,N_513,N_4274);
nor U6112 (N_6112,N_1789,N_2313);
or U6113 (N_6113,N_3323,N_4078);
xnor U6114 (N_6114,N_3143,N_384);
or U6115 (N_6115,N_286,N_4881);
or U6116 (N_6116,N_2196,N_600);
xor U6117 (N_6117,N_1444,N_4589);
and U6118 (N_6118,N_1464,N_4567);
or U6119 (N_6119,N_1141,N_2760);
and U6120 (N_6120,N_1013,N_4276);
nor U6121 (N_6121,N_2302,N_2467);
and U6122 (N_6122,N_1671,N_3723);
or U6123 (N_6123,N_3092,N_3368);
nor U6124 (N_6124,N_1093,N_2686);
or U6125 (N_6125,N_1548,N_2294);
nand U6126 (N_6126,N_4335,N_4326);
xnor U6127 (N_6127,N_1983,N_4478);
and U6128 (N_6128,N_3790,N_4680);
nor U6129 (N_6129,N_3424,N_1686);
xor U6130 (N_6130,N_3403,N_1);
nor U6131 (N_6131,N_1070,N_758);
and U6132 (N_6132,N_1912,N_2055);
and U6133 (N_6133,N_3370,N_1786);
or U6134 (N_6134,N_2595,N_1472);
nor U6135 (N_6135,N_3413,N_376);
xnor U6136 (N_6136,N_1412,N_166);
nand U6137 (N_6137,N_4688,N_3011);
xor U6138 (N_6138,N_195,N_2608);
nand U6139 (N_6139,N_288,N_2253);
nor U6140 (N_6140,N_1800,N_819);
and U6141 (N_6141,N_3062,N_2511);
xnor U6142 (N_6142,N_2944,N_3758);
nor U6143 (N_6143,N_679,N_3032);
xnor U6144 (N_6144,N_3491,N_3333);
nor U6145 (N_6145,N_2406,N_4443);
nand U6146 (N_6146,N_1555,N_4371);
nor U6147 (N_6147,N_4463,N_2365);
xnor U6148 (N_6148,N_4098,N_1253);
nor U6149 (N_6149,N_2609,N_82);
or U6150 (N_6150,N_735,N_1515);
nand U6151 (N_6151,N_3309,N_3461);
or U6152 (N_6152,N_3065,N_1269);
and U6153 (N_6153,N_4614,N_1283);
nor U6154 (N_6154,N_786,N_3865);
or U6155 (N_6155,N_4608,N_4124);
nand U6156 (N_6156,N_3341,N_2354);
and U6157 (N_6157,N_1782,N_1078);
nand U6158 (N_6158,N_2436,N_2704);
nor U6159 (N_6159,N_4944,N_2502);
nand U6160 (N_6160,N_4547,N_490);
xnor U6161 (N_6161,N_2859,N_404);
xnor U6162 (N_6162,N_1794,N_2858);
and U6163 (N_6163,N_4437,N_2500);
nand U6164 (N_6164,N_530,N_2999);
xor U6165 (N_6165,N_897,N_3976);
or U6166 (N_6166,N_2223,N_3399);
and U6167 (N_6167,N_374,N_1249);
nor U6168 (N_6168,N_3084,N_4918);
and U6169 (N_6169,N_361,N_4170);
and U6170 (N_6170,N_3226,N_1181);
nor U6171 (N_6171,N_4803,N_360);
xor U6172 (N_6172,N_2623,N_818);
xor U6173 (N_6173,N_1626,N_3496);
xor U6174 (N_6174,N_884,N_280);
xnor U6175 (N_6175,N_787,N_3506);
nand U6176 (N_6176,N_3900,N_3537);
xor U6177 (N_6177,N_397,N_1726);
nor U6178 (N_6178,N_4565,N_1967);
nor U6179 (N_6179,N_2464,N_4899);
nor U6180 (N_6180,N_2604,N_1273);
nor U6181 (N_6181,N_541,N_3659);
and U6182 (N_6182,N_1673,N_2377);
nand U6183 (N_6183,N_747,N_3041);
nand U6184 (N_6184,N_4927,N_3765);
nor U6185 (N_6185,N_4536,N_1850);
nand U6186 (N_6186,N_1759,N_3644);
xnor U6187 (N_6187,N_2369,N_2900);
nor U6188 (N_6188,N_2250,N_4766);
or U6189 (N_6189,N_3104,N_574);
and U6190 (N_6190,N_3157,N_2345);
xor U6191 (N_6191,N_2050,N_3324);
xor U6192 (N_6192,N_2605,N_3040);
nand U6193 (N_6193,N_3042,N_1370);
nand U6194 (N_6194,N_1520,N_2072);
nand U6195 (N_6195,N_1874,N_1552);
or U6196 (N_6196,N_3066,N_3709);
xor U6197 (N_6197,N_4618,N_3528);
or U6198 (N_6198,N_890,N_1142);
and U6199 (N_6199,N_1752,N_1135);
and U6200 (N_6200,N_2353,N_2687);
and U6201 (N_6201,N_443,N_4673);
xnor U6202 (N_6202,N_2336,N_4761);
and U6203 (N_6203,N_1755,N_1768);
xnor U6204 (N_6204,N_1063,N_741);
nor U6205 (N_6205,N_2360,N_172);
xor U6206 (N_6206,N_4088,N_1108);
and U6207 (N_6207,N_3451,N_653);
xnor U6208 (N_6208,N_3522,N_1646);
nand U6209 (N_6209,N_3343,N_4799);
nand U6210 (N_6210,N_492,N_3817);
and U6211 (N_6211,N_270,N_3422);
nor U6212 (N_6212,N_2348,N_4038);
nor U6213 (N_6213,N_775,N_4713);
and U6214 (N_6214,N_1305,N_377);
or U6215 (N_6215,N_618,N_4372);
nor U6216 (N_6216,N_3774,N_611);
xor U6217 (N_6217,N_4895,N_862);
nand U6218 (N_6218,N_4994,N_2034);
nor U6219 (N_6219,N_4925,N_1847);
nor U6220 (N_6220,N_4069,N_889);
nand U6221 (N_6221,N_4612,N_3845);
xnor U6222 (N_6222,N_3019,N_3950);
xnor U6223 (N_6223,N_652,N_1421);
and U6224 (N_6224,N_4540,N_576);
xor U6225 (N_6225,N_3673,N_2045);
and U6226 (N_6226,N_4485,N_1592);
nor U6227 (N_6227,N_988,N_560);
and U6228 (N_6228,N_3158,N_191);
nor U6229 (N_6229,N_1836,N_3198);
xor U6230 (N_6230,N_3875,N_3044);
xor U6231 (N_6231,N_4787,N_3719);
xor U6232 (N_6232,N_4584,N_539);
and U6233 (N_6233,N_4010,N_1307);
nor U6234 (N_6234,N_3598,N_4225);
or U6235 (N_6235,N_2640,N_1680);
xnor U6236 (N_6236,N_4631,N_4892);
nor U6237 (N_6237,N_3134,N_2082);
nand U6238 (N_6238,N_3054,N_1051);
nor U6239 (N_6239,N_162,N_3989);
and U6240 (N_6240,N_475,N_2641);
nor U6241 (N_6241,N_1774,N_1890);
and U6242 (N_6242,N_1797,N_4189);
and U6243 (N_6243,N_4579,N_4208);
xor U6244 (N_6244,N_3854,N_3190);
nand U6245 (N_6245,N_2725,N_526);
xor U6246 (N_6246,N_2543,N_398);
and U6247 (N_6247,N_725,N_2090);
nor U6248 (N_6248,N_1915,N_4982);
nand U6249 (N_6249,N_193,N_2534);
xor U6250 (N_6250,N_1035,N_1062);
nand U6251 (N_6251,N_4043,N_267);
and U6252 (N_6252,N_4532,N_2495);
nand U6253 (N_6253,N_3535,N_829);
xnor U6254 (N_6254,N_167,N_412);
and U6255 (N_6255,N_1703,N_4163);
xnor U6256 (N_6256,N_473,N_1374);
nand U6257 (N_6257,N_4786,N_1972);
nand U6258 (N_6258,N_4234,N_860);
xnor U6259 (N_6259,N_2645,N_1379);
or U6260 (N_6260,N_1578,N_2080);
nor U6261 (N_6261,N_4349,N_4412);
xor U6262 (N_6262,N_4269,N_623);
nand U6263 (N_6263,N_442,N_1016);
nand U6264 (N_6264,N_2297,N_3965);
or U6265 (N_6265,N_926,N_58);
and U6266 (N_6266,N_813,N_2001);
or U6267 (N_6267,N_547,N_4759);
nand U6268 (N_6268,N_3276,N_3770);
xnor U6269 (N_6269,N_4149,N_2947);
nand U6270 (N_6270,N_2692,N_1212);
xor U6271 (N_6271,N_2490,N_4522);
or U6272 (N_6272,N_4698,N_2882);
xnor U6273 (N_6273,N_2187,N_1289);
nor U6274 (N_6274,N_4897,N_205);
nor U6275 (N_6275,N_1131,N_2031);
nand U6276 (N_6276,N_1689,N_3164);
nor U6277 (N_6277,N_519,N_3224);
nand U6278 (N_6278,N_4839,N_1681);
and U6279 (N_6279,N_2027,N_1647);
xor U6280 (N_6280,N_2133,N_4339);
nand U6281 (N_6281,N_1823,N_3661);
nor U6282 (N_6282,N_898,N_2255);
or U6283 (N_6283,N_718,N_3937);
xnor U6284 (N_6284,N_2591,N_428);
and U6285 (N_6285,N_663,N_3350);
and U6286 (N_6286,N_3213,N_2428);
nor U6287 (N_6287,N_3669,N_963);
nor U6288 (N_6288,N_3869,N_1091);
and U6289 (N_6289,N_29,N_1121);
or U6290 (N_6290,N_2111,N_3585);
nor U6291 (N_6291,N_3893,N_1019);
xor U6292 (N_6292,N_3476,N_1720);
xor U6293 (N_6293,N_3569,N_1725);
xor U6294 (N_6294,N_4652,N_1524);
and U6295 (N_6295,N_4790,N_2009);
nor U6296 (N_6296,N_3189,N_4297);
or U6297 (N_6297,N_3161,N_1634);
nor U6298 (N_6298,N_3373,N_4444);
or U6299 (N_6299,N_3205,N_2575);
xnor U6300 (N_6300,N_3285,N_208);
nand U6301 (N_6301,N_2918,N_4752);
and U6302 (N_6302,N_3686,N_243);
nor U6303 (N_6303,N_3995,N_4776);
xor U6304 (N_6304,N_4013,N_1447);
xor U6305 (N_6305,N_2213,N_3301);
xor U6306 (N_6306,N_1758,N_1770);
xnor U6307 (N_6307,N_4272,N_585);
and U6308 (N_6308,N_3046,N_1040);
nor U6309 (N_6309,N_1193,N_3942);
and U6310 (N_6310,N_1207,N_4196);
nor U6311 (N_6311,N_4740,N_607);
or U6312 (N_6312,N_3100,N_2309);
nand U6313 (N_6313,N_4604,N_3053);
nand U6314 (N_6314,N_4090,N_1751);
and U6315 (N_6315,N_4000,N_4715);
and U6316 (N_6316,N_3957,N_4278);
or U6317 (N_6317,N_2870,N_2375);
nor U6318 (N_6318,N_2625,N_4883);
xnor U6319 (N_6319,N_1334,N_537);
and U6320 (N_6320,N_3941,N_1944);
or U6321 (N_6321,N_1061,N_3385);
xor U6322 (N_6322,N_2715,N_1293);
and U6323 (N_6323,N_1657,N_4089);
xnor U6324 (N_6324,N_1126,N_4672);
and U6325 (N_6325,N_2205,N_1834);
and U6326 (N_6326,N_1856,N_824);
or U6327 (N_6327,N_2526,N_4535);
nor U6328 (N_6328,N_981,N_296);
nand U6329 (N_6329,N_3490,N_4807);
and U6330 (N_6330,N_4586,N_2596);
or U6331 (N_6331,N_4388,N_3829);
or U6332 (N_6332,N_1440,N_2397);
nand U6333 (N_6333,N_2710,N_127);
nand U6334 (N_6334,N_3302,N_488);
xnor U6335 (N_6335,N_1052,N_2226);
or U6336 (N_6336,N_4074,N_4778);
nor U6337 (N_6337,N_4171,N_4213);
or U6338 (N_6338,N_3591,N_3315);
nand U6339 (N_6339,N_746,N_4014);
and U6340 (N_6340,N_1215,N_2197);
xor U6341 (N_6341,N_4244,N_931);
nor U6342 (N_6342,N_27,N_4859);
and U6343 (N_6343,N_4788,N_84);
and U6344 (N_6344,N_2789,N_1432);
and U6345 (N_6345,N_2899,N_3627);
nand U6346 (N_6346,N_468,N_3824);
xnor U6347 (N_6347,N_1486,N_4132);
and U6348 (N_6348,N_2915,N_2724);
xor U6349 (N_6349,N_2268,N_1111);
and U6350 (N_6350,N_2854,N_2853);
or U6351 (N_6351,N_1694,N_299);
nor U6352 (N_6352,N_4067,N_4462);
nor U6353 (N_6353,N_2087,N_4409);
nor U6354 (N_6354,N_4251,N_3615);
xnor U6355 (N_6355,N_1303,N_3592);
xnor U6356 (N_6356,N_4521,N_4678);
and U6357 (N_6357,N_4770,N_985);
and U6358 (N_6358,N_2785,N_752);
nor U6359 (N_6359,N_186,N_1664);
nand U6360 (N_6360,N_3834,N_4916);
xnor U6361 (N_6361,N_4830,N_751);
nor U6362 (N_6362,N_1892,N_3507);
and U6363 (N_6363,N_3074,N_254);
or U6364 (N_6364,N_3127,N_3028);
nand U6365 (N_6365,N_4077,N_1649);
xor U6366 (N_6366,N_810,N_1575);
nand U6367 (N_6367,N_2891,N_987);
or U6368 (N_6368,N_2156,N_512);
nand U6369 (N_6369,N_4212,N_532);
nor U6370 (N_6370,N_4129,N_1468);
nand U6371 (N_6371,N_1530,N_843);
or U6372 (N_6372,N_4289,N_620);
nor U6373 (N_6373,N_4293,N_2487);
and U6374 (N_6374,N_110,N_3879);
nor U6375 (N_6375,N_4421,N_561);
nand U6376 (N_6376,N_4325,N_4422);
nand U6377 (N_6377,N_369,N_4209);
nand U6378 (N_6378,N_4021,N_3485);
nand U6379 (N_6379,N_4185,N_3920);
xnor U6380 (N_6380,N_1594,N_1604);
xnor U6381 (N_6381,N_1096,N_2260);
nor U6382 (N_6382,N_1901,N_4046);
nand U6383 (N_6383,N_3214,N_3165);
nand U6384 (N_6384,N_3227,N_4931);
or U6385 (N_6385,N_3072,N_2866);
or U6386 (N_6386,N_3849,N_3438);
or U6387 (N_6387,N_4953,N_2019);
xor U6388 (N_6388,N_4889,N_3718);
nor U6389 (N_6389,N_4760,N_1477);
xnor U6390 (N_6390,N_67,N_255);
xnor U6391 (N_6391,N_950,N_2335);
nor U6392 (N_6392,N_227,N_1154);
or U6393 (N_6393,N_1343,N_4122);
and U6394 (N_6394,N_2912,N_1675);
nand U6395 (N_6395,N_1439,N_4758);
and U6396 (N_6396,N_3607,N_4242);
and U6397 (N_6397,N_73,N_3589);
or U6398 (N_6398,N_156,N_330);
nand U6399 (N_6399,N_1224,N_4295);
or U6400 (N_6400,N_1609,N_2071);
or U6401 (N_6401,N_364,N_47);
nor U6402 (N_6402,N_3763,N_3711);
or U6403 (N_6403,N_920,N_3024);
nand U6404 (N_6404,N_4062,N_2929);
or U6405 (N_6405,N_4330,N_79);
or U6406 (N_6406,N_4490,N_1825);
nor U6407 (N_6407,N_648,N_3611);
xor U6408 (N_6408,N_637,N_3573);
and U6409 (N_6409,N_4051,N_4813);
nand U6410 (N_6410,N_3102,N_1999);
nand U6411 (N_6411,N_2236,N_3239);
and U6412 (N_6412,N_1535,N_1795);
and U6413 (N_6413,N_1760,N_1262);
nand U6414 (N_6414,N_228,N_580);
nand U6415 (N_6415,N_2981,N_4238);
nor U6416 (N_6416,N_4083,N_4518);
xor U6417 (N_6417,N_2621,N_2437);
nand U6418 (N_6418,N_4667,N_318);
and U6419 (N_6419,N_4343,N_4581);
nand U6420 (N_6420,N_3035,N_3137);
and U6421 (N_6421,N_4450,N_3187);
and U6422 (N_6422,N_3850,N_3645);
and U6423 (N_6423,N_339,N_409);
xnor U6424 (N_6424,N_1306,N_2006);
xor U6425 (N_6425,N_601,N_3772);
nor U6426 (N_6426,N_4458,N_3608);
xor U6427 (N_6427,N_4466,N_3268);
nor U6428 (N_6428,N_4282,N_3984);
nor U6429 (N_6429,N_1255,N_4922);
xnor U6430 (N_6430,N_124,N_2585);
nor U6431 (N_6431,N_3021,N_3135);
nor U6432 (N_6432,N_1176,N_498);
xor U6433 (N_6433,N_2155,N_4313);
nand U6434 (N_6434,N_3811,N_3621);
xnor U6435 (N_6435,N_665,N_2860);
or U6436 (N_6436,N_3038,N_1802);
xnor U6437 (N_6437,N_4747,N_879);
xnor U6438 (N_6438,N_1821,N_2104);
nand U6439 (N_6439,N_402,N_275);
nor U6440 (N_6440,N_3468,N_956);
and U6441 (N_6441,N_1336,N_2057);
nor U6442 (N_6442,N_3404,N_3348);
or U6443 (N_6443,N_2175,N_1296);
nor U6444 (N_6444,N_3483,N_2719);
nand U6445 (N_6445,N_806,N_2690);
and U6446 (N_6446,N_1654,N_1147);
nand U6447 (N_6447,N_4262,N_4142);
nor U6448 (N_6448,N_2685,N_930);
and U6449 (N_6449,N_30,N_466);
and U6450 (N_6450,N_1302,N_772);
xor U6451 (N_6451,N_2378,N_2868);
or U6452 (N_6452,N_3193,N_2728);
and U6453 (N_6453,N_197,N_1722);
nor U6454 (N_6454,N_2550,N_1934);
and U6455 (N_6455,N_1702,N_3430);
nand U6456 (N_6456,N_2925,N_2668);
xor U6457 (N_6457,N_2048,N_2688);
or U6458 (N_6458,N_2698,N_1279);
nand U6459 (N_6459,N_3953,N_2980);
nor U6460 (N_6460,N_1337,N_1220);
and U6461 (N_6461,N_903,N_722);
and U6462 (N_6462,N_3495,N_4936);
nor U6463 (N_6463,N_3228,N_3972);
and U6464 (N_6464,N_4701,N_1868);
nor U6465 (N_6465,N_1730,N_3842);
and U6466 (N_6466,N_3258,N_4647);
nand U6467 (N_6467,N_1737,N_785);
and U6468 (N_6468,N_450,N_2772);
nor U6469 (N_6469,N_187,N_1320);
or U6470 (N_6470,N_4654,N_3863);
nand U6471 (N_6471,N_3759,N_1854);
or U6472 (N_6472,N_4502,N_3063);
and U6473 (N_6473,N_4063,N_2679);
xnor U6474 (N_6474,N_643,N_2149);
xor U6475 (N_6475,N_2594,N_2967);
nand U6476 (N_6476,N_2510,N_4445);
nor U6477 (N_6477,N_3405,N_3979);
nor U6478 (N_6478,N_4957,N_1859);
nand U6479 (N_6479,N_3642,N_4291);
xnor U6480 (N_6480,N_511,N_2705);
and U6481 (N_6481,N_3068,N_23);
nor U6482 (N_6482,N_2736,N_3150);
or U6483 (N_6483,N_3017,N_3514);
nor U6484 (N_6484,N_1017,N_568);
or U6485 (N_6485,N_3964,N_4220);
nor U6486 (N_6486,N_2110,N_3255);
xnor U6487 (N_6487,N_1676,N_1841);
xor U6488 (N_6488,N_1993,N_2682);
or U6489 (N_6489,N_1736,N_590);
xor U6490 (N_6490,N_120,N_2784);
xnor U6491 (N_6491,N_4416,N_2695);
nor U6492 (N_6492,N_248,N_1962);
nor U6493 (N_6493,N_1368,N_2806);
xor U6494 (N_6494,N_1745,N_2634);
and U6495 (N_6495,N_4472,N_4094);
xor U6496 (N_6496,N_651,N_626);
nor U6497 (N_6497,N_3706,N_3594);
or U6498 (N_6498,N_2969,N_1217);
and U6499 (N_6499,N_4828,N_4771);
nor U6500 (N_6500,N_4735,N_4743);
or U6501 (N_6501,N_46,N_4186);
nand U6502 (N_6502,N_2556,N_4993);
and U6503 (N_6503,N_3139,N_2010);
xnor U6504 (N_6504,N_3194,N_2932);
and U6505 (N_6505,N_3870,N_812);
nor U6506 (N_6506,N_734,N_674);
or U6507 (N_6507,N_2351,N_2706);
or U6508 (N_6508,N_3651,N_3172);
and U6509 (N_6509,N_1706,N_4657);
and U6510 (N_6510,N_1145,N_1551);
nor U6511 (N_6511,N_3277,N_3688);
and U6512 (N_6512,N_3743,N_2895);
xnor U6513 (N_6513,N_1204,N_566);
xnor U6514 (N_6514,N_4704,N_629);
or U6515 (N_6515,N_4413,N_2924);
xor U6516 (N_6516,N_2064,N_2074);
and U6517 (N_6517,N_3004,N_1941);
or U6518 (N_6518,N_793,N_4340);
nor U6519 (N_6519,N_3708,N_3095);
nand U6520 (N_6520,N_2571,N_219);
nor U6521 (N_6521,N_3151,N_2327);
and U6522 (N_6522,N_520,N_3079);
nand U6523 (N_6523,N_1435,N_2748);
xnor U6524 (N_6524,N_4842,N_3539);
nor U6525 (N_6525,N_1936,N_1994);
xor U6526 (N_6526,N_2998,N_1346);
or U6527 (N_6527,N_589,N_3126);
and U6528 (N_6528,N_2818,N_477);
or U6529 (N_6529,N_730,N_4434);
xor U6530 (N_6530,N_1747,N_1887);
xnor U6531 (N_6531,N_2498,N_1919);
and U6532 (N_6532,N_2867,N_3289);
or U6533 (N_6533,N_2315,N_2107);
nand U6534 (N_6534,N_1740,N_2664);
nor U6535 (N_6535,N_4034,N_534);
nand U6536 (N_6536,N_3057,N_1839);
and U6537 (N_6537,N_4309,N_3921);
nor U6538 (N_6538,N_1243,N_33);
or U6539 (N_6539,N_3334,N_3784);
nor U6540 (N_6540,N_2826,N_1576);
or U6541 (N_6541,N_3359,N_1573);
or U6542 (N_6542,N_4188,N_1347);
or U6543 (N_6543,N_1701,N_1932);
nand U6544 (N_6544,N_1295,N_4037);
nand U6545 (N_6545,N_4145,N_3769);
nand U6546 (N_6546,N_1687,N_841);
or U6547 (N_6547,N_1727,N_828);
xor U6548 (N_6548,N_1065,N_4943);
and U6549 (N_6549,N_4071,N_1662);
nor U6550 (N_6550,N_1677,N_1659);
nor U6551 (N_6551,N_4564,N_4573);
or U6552 (N_6552,N_476,N_609);
nor U6553 (N_6553,N_2407,N_3929);
or U6554 (N_6554,N_1522,N_2564);
and U6555 (N_6555,N_4846,N_2610);
and U6556 (N_6556,N_4516,N_3048);
nand U6557 (N_6557,N_2970,N_2662);
and U6558 (N_6558,N_1172,N_2454);
xnor U6559 (N_6559,N_1188,N_77);
xor U6560 (N_6560,N_1175,N_112);
and U6561 (N_6561,N_329,N_1428);
and U6562 (N_6562,N_1012,N_3890);
and U6563 (N_6563,N_1014,N_2942);
and U6564 (N_6564,N_3078,N_72);
and U6565 (N_6565,N_3777,N_896);
nand U6566 (N_6566,N_3191,N_4316);
or U6567 (N_6567,N_4363,N_3458);
xor U6568 (N_6568,N_871,N_1771);
or U6569 (N_6569,N_4486,N_3096);
and U6570 (N_6570,N_941,N_3060);
xnor U6571 (N_6571,N_814,N_2749);
and U6572 (N_6572,N_790,N_1550);
nand U6573 (N_6573,N_394,N_1409);
xor U6574 (N_6574,N_1955,N_4348);
and U6575 (N_6575,N_2518,N_4702);
nor U6576 (N_6576,N_1635,N_462);
and U6577 (N_6577,N_109,N_1072);
nand U6578 (N_6578,N_1248,N_767);
nand U6579 (N_6579,N_365,N_1442);
or U6580 (N_6580,N_1309,N_2266);
nand U6581 (N_6581,N_953,N_2535);
nor U6582 (N_6582,N_2549,N_1401);
nor U6583 (N_6583,N_1474,N_1263);
nand U6584 (N_6584,N_3210,N_924);
nor U6585 (N_6585,N_4407,N_3415);
or U6586 (N_6586,N_2875,N_4480);
xnor U6587 (N_6587,N_4615,N_3250);
nor U6588 (N_6588,N_4929,N_344);
nor U6589 (N_6589,N_3939,N_4433);
nand U6590 (N_6590,N_2296,N_4886);
nand U6591 (N_6591,N_4468,N_2129);
xor U6592 (N_6592,N_3448,N_4714);
nand U6593 (N_6593,N_2532,N_3378);
nand U6594 (N_6594,N_2751,N_2847);
nor U6595 (N_6595,N_334,N_3997);
and U6596 (N_6596,N_2560,N_1127);
and U6597 (N_6597,N_104,N_3543);
nand U6598 (N_6598,N_1968,N_3691);
xor U6599 (N_6599,N_2300,N_913);
xnor U6600 (N_6600,N_1638,N_1264);
or U6601 (N_6601,N_1773,N_2941);
nand U6602 (N_6602,N_1103,N_1396);
nand U6603 (N_6603,N_4026,N_60);
nor U6604 (N_6604,N_1294,N_1518);
or U6605 (N_6605,N_1966,N_2380);
or U6606 (N_6606,N_4075,N_3243);
xnor U6607 (N_6607,N_4613,N_4812);
xnor U6608 (N_6608,N_2329,N_2520);
nor U6609 (N_6609,N_143,N_658);
nand U6610 (N_6610,N_1353,N_3120);
xor U6611 (N_6611,N_3094,N_3306);
or U6612 (N_6612,N_3581,N_2445);
or U6613 (N_6613,N_3425,N_3050);
nand U6614 (N_6614,N_694,N_3568);
nand U6615 (N_6615,N_2729,N_788);
nor U6616 (N_6616,N_3731,N_1830);
and U6617 (N_6617,N_1831,N_2316);
nand U6618 (N_6618,N_1392,N_3281);
nand U6619 (N_6619,N_452,N_4322);
nand U6620 (N_6620,N_914,N_2042);
and U6621 (N_6621,N_4260,N_1240);
and U6622 (N_6622,N_3536,N_4005);
or U6623 (N_6623,N_1394,N_429);
and U6624 (N_6624,N_3967,N_852);
nor U6625 (N_6625,N_1924,N_3264);
or U6626 (N_6626,N_326,N_3328);
nor U6627 (N_6627,N_1987,N_1632);
nor U6628 (N_6628,N_250,N_3635);
nand U6629 (N_6629,N_266,N_1583);
nor U6630 (N_6630,N_768,N_210);
and U6631 (N_6631,N_1080,N_125);
xor U6632 (N_6632,N_1389,N_4966);
xnor U6633 (N_6633,N_3352,N_4975);
and U6634 (N_6634,N_4428,N_3848);
and U6635 (N_6635,N_4039,N_661);
or U6636 (N_6636,N_4968,N_1511);
xnor U6637 (N_6637,N_1022,N_2991);
or U6638 (N_6638,N_51,N_647);
xnor U6639 (N_6639,N_4019,N_3014);
nor U6640 (N_6640,N_2573,N_4500);
nor U6641 (N_6641,N_1371,N_3085);
nor U6642 (N_6642,N_4728,N_3488);
nor U6643 (N_6643,N_2025,N_2953);
xor U6644 (N_6644,N_2004,N_4559);
xor U6645 (N_6645,N_4246,N_3884);
and U6646 (N_6646,N_4265,N_3221);
and U6647 (N_6647,N_2689,N_1349);
or U6648 (N_6648,N_2014,N_179);
nor U6649 (N_6649,N_3980,N_4368);
or U6650 (N_6650,N_1058,N_2653);
or U6651 (N_6651,N_2977,N_4158);
or U6652 (N_6652,N_823,N_2416);
and U6653 (N_6653,N_1107,N_3012);
nand U6654 (N_6654,N_522,N_2172);
and U6655 (N_6655,N_2950,N_438);
nor U6656 (N_6656,N_2189,N_975);
and U6657 (N_6657,N_1805,N_4006);
xnor U6658 (N_6658,N_2863,N_4732);
and U6659 (N_6659,N_676,N_986);
and U6660 (N_6660,N_1844,N_3508);
or U6661 (N_6661,N_1466,N_2703);
nand U6662 (N_6662,N_867,N_990);
or U6663 (N_6663,N_3005,N_2169);
xor U6664 (N_6664,N_4477,N_3662);
and U6665 (N_6665,N_1602,N_234);
and U6666 (N_6666,N_2468,N_1272);
xor U6667 (N_6667,N_4183,N_1842);
or U6668 (N_6668,N_2914,N_3138);
nor U6669 (N_6669,N_2821,N_4197);
xnor U6670 (N_6670,N_1504,N_4600);
and U6671 (N_6671,N_1559,N_4910);
nand U6672 (N_6672,N_2462,N_1377);
nor U6673 (N_6673,N_1117,N_1674);
nand U6674 (N_6674,N_2470,N_2796);
nor U6675 (N_6675,N_4492,N_1450);
nor U6676 (N_6676,N_3844,N_1566);
and U6677 (N_6677,N_1258,N_1619);
xor U6678 (N_6678,N_3183,N_4934);
or U6679 (N_6679,N_2131,N_4240);
and U6680 (N_6680,N_3601,N_2450);
nor U6681 (N_6681,N_645,N_3449);
and U6682 (N_6682,N_4395,N_2928);
or U6683 (N_6683,N_827,N_3796);
nand U6684 (N_6684,N_1436,N_4055);
and U6685 (N_6685,N_2344,N_3123);
or U6686 (N_6686,N_1948,N_1803);
nand U6687 (N_6687,N_379,N_685);
xor U6688 (N_6688,N_4059,N_2115);
or U6689 (N_6689,N_933,N_2405);
nor U6690 (N_6690,N_2394,N_1572);
and U6691 (N_6691,N_794,N_3712);
xnor U6692 (N_6692,N_4919,N_4571);
xnor U6693 (N_6693,N_1237,N_4332);
or U6694 (N_6694,N_2337,N_3609);
nor U6695 (N_6695,N_836,N_3388);
or U6696 (N_6696,N_1580,N_4582);
xor U6697 (N_6697,N_4791,N_832);
or U6698 (N_6698,N_1403,N_1517);
nand U6699 (N_6699,N_1471,N_3006);
nor U6700 (N_6700,N_200,N_946);
nand U6701 (N_6701,N_3335,N_4734);
nor U6702 (N_6702,N_3030,N_3356);
nor U6703 (N_6703,N_2228,N_2963);
xnor U6704 (N_6704,N_106,N_1614);
nor U6705 (N_6705,N_4365,N_3336);
nor U6706 (N_6706,N_4216,N_3775);
nor U6707 (N_6707,N_2768,N_689);
nor U6708 (N_6708,N_2137,N_3567);
or U6709 (N_6709,N_2988,N_3738);
nor U6710 (N_6710,N_3987,N_2537);
and U6711 (N_6711,N_1380,N_2067);
nand U6712 (N_6712,N_4977,N_4489);
or U6713 (N_6713,N_1350,N_2421);
nand U6714 (N_6714,N_2171,N_4182);
nor U6715 (N_6715,N_1724,N_4436);
xor U6716 (N_6716,N_3650,N_4139);
xnor U6717 (N_6717,N_1208,N_4555);
and U6718 (N_6718,N_711,N_217);
or U6719 (N_6719,N_2340,N_4249);
nand U6720 (N_6720,N_4806,N_353);
nor U6721 (N_6721,N_1358,N_201);
xnor U6722 (N_6722,N_4554,N_3375);
or U6723 (N_6723,N_1433,N_2399);
or U6724 (N_6724,N_1362,N_2453);
and U6725 (N_6725,N_728,N_3376);
nand U6726 (N_6726,N_2191,N_3701);
or U6727 (N_6727,N_1457,N_378);
xnor U6728 (N_6728,N_3787,N_4817);
and U6729 (N_6729,N_1693,N_1996);
nand U6730 (N_6730,N_701,N_1174);
xor U6731 (N_6731,N_2862,N_650);
and U6732 (N_6732,N_1808,N_2780);
nor U6733 (N_6733,N_4971,N_4029);
xor U6734 (N_6734,N_4887,N_3203);
and U6735 (N_6735,N_1584,N_835);
nor U6736 (N_6736,N_3282,N_3951);
xor U6737 (N_6737,N_236,N_2105);
or U6738 (N_6738,N_178,N_1036);
nor U6739 (N_6739,N_4870,N_2089);
nor U6740 (N_6740,N_4689,N_4780);
or U6741 (N_6741,N_4950,N_2655);
or U6742 (N_6742,N_1545,N_3561);
nand U6743 (N_6743,N_2028,N_387);
or U6744 (N_6744,N_865,N_3170);
and U6745 (N_6745,N_4161,N_3653);
xor U6746 (N_6746,N_2430,N_2883);
nor U6747 (N_6747,N_4248,N_4826);
nor U6748 (N_6748,N_294,N_3672);
or U6749 (N_6749,N_2411,N_261);
or U6750 (N_6750,N_4855,N_4414);
xor U6751 (N_6751,N_4386,N_2262);
nand U6752 (N_6752,N_2993,N_457);
or U6753 (N_6753,N_1877,N_3767);
nand U6754 (N_6754,N_4517,N_1338);
or U6755 (N_6755,N_687,N_2747);
and U6756 (N_6756,N_2433,N_820);
nand U6757 (N_6757,N_3207,N_1190);
nand U6758 (N_6758,N_2109,N_2393);
nor U6759 (N_6759,N_2880,N_4676);
or U6760 (N_6760,N_4985,N_2813);
or U6761 (N_6761,N_206,N_4261);
nor U6762 (N_6762,N_4427,N_3234);
and U6763 (N_6763,N_4785,N_672);
nor U6764 (N_6764,N_4398,N_2148);
xnor U6765 (N_6765,N_3195,N_1020);
nor U6766 (N_6766,N_4534,N_4570);
nand U6767 (N_6767,N_4025,N_4692);
and U6768 (N_6768,N_222,N_482);
or U6769 (N_6769,N_3107,N_1958);
xnor U6770 (N_6770,N_87,N_3724);
nand U6771 (N_6771,N_1621,N_4753);
and U6772 (N_6772,N_2804,N_4840);
xnor U6773 (N_6773,N_3432,N_1587);
xnor U6774 (N_6774,N_238,N_4497);
and U6775 (N_6775,N_1102,N_302);
and U6776 (N_6776,N_1913,N_2240);
nand U6777 (N_6777,N_1933,N_3121);
and U6778 (N_6778,N_802,N_4864);
xnor U6779 (N_6779,N_4731,N_2417);
nand U6780 (N_6780,N_4868,N_3197);
nand U6781 (N_6781,N_3502,N_1182);
xor U6782 (N_6782,N_1085,N_3880);
and U6783 (N_6783,N_4558,N_349);
xnor U6784 (N_6784,N_1527,N_947);
nor U6785 (N_6785,N_3454,N_1209);
or U6786 (N_6786,N_3690,N_549);
nand U6787 (N_6787,N_2936,N_4987);
nand U6788 (N_6788,N_321,N_4138);
xor U6789 (N_6789,N_3524,N_1952);
nand U6790 (N_6790,N_2152,N_708);
xnor U6791 (N_6791,N_3832,N_2125);
or U6792 (N_6792,N_4632,N_1620);
or U6793 (N_6793,N_4222,N_3241);
nand U6794 (N_6794,N_1875,N_4831);
xnor U6795 (N_6795,N_1089,N_1625);
or U6796 (N_6796,N_2177,N_4835);
xnor U6797 (N_6797,N_4044,N_3961);
xnor U6798 (N_6798,N_4218,N_816);
nor U6799 (N_6799,N_2200,N_239);
xor U6800 (N_6800,N_502,N_2541);
nand U6801 (N_6801,N_964,N_113);
nor U6802 (N_6802,N_1900,N_1651);
and U6803 (N_6803,N_3000,N_1757);
and U6804 (N_6804,N_4401,N_4033);
and U6805 (N_6805,N_2331,N_1330);
nand U6806 (N_6806,N_2281,N_2391);
and U6807 (N_6807,N_3992,N_1044);
or U6808 (N_6808,N_436,N_232);
nor U6809 (N_6809,N_2447,N_2456);
xnor U6810 (N_6810,N_1041,N_4354);
and U6811 (N_6811,N_1261,N_4329);
and U6812 (N_6812,N_4719,N_799);
or U6813 (N_6813,N_3303,N_3472);
nor U6814 (N_6814,N_3999,N_690);
xnor U6815 (N_6815,N_3930,N_3481);
nand U6816 (N_6816,N_3871,N_591);
nand U6817 (N_6817,N_4682,N_4355);
or U6818 (N_6818,N_4361,N_2023);
and U6819 (N_6819,N_3275,N_53);
and U6820 (N_6820,N_2251,N_2041);
xnor U6821 (N_6821,N_430,N_1586);
or U6822 (N_6822,N_1416,N_2974);
xor U6823 (N_6823,N_954,N_3321);
and U6824 (N_6824,N_2134,N_3342);
xnor U6825 (N_6825,N_17,N_3202);
and U6826 (N_6826,N_3292,N_4080);
nor U6827 (N_6827,N_510,N_2579);
xor U6828 (N_6828,N_2945,N_3129);
or U6829 (N_6829,N_3209,N_130);
and U6830 (N_6830,N_3680,N_2084);
xor U6831 (N_6831,N_4290,N_4456);
or U6832 (N_6832,N_2122,N_3786);
or U6833 (N_6833,N_3750,N_1846);
nand U6834 (N_6834,N_3401,N_1848);
and U6835 (N_6835,N_1333,N_3305);
nand U6836 (N_6836,N_432,N_3274);
nand U6837 (N_6837,N_4273,N_435);
nor U6838 (N_6838,N_4691,N_2341);
and U6839 (N_6839,N_2046,N_1155);
and U6840 (N_6840,N_1611,N_3841);
and U6841 (N_6841,N_4102,N_3160);
xnor U6842 (N_6842,N_1406,N_3493);
or U6843 (N_6843,N_1321,N_2807);
xnor U6844 (N_6844,N_3695,N_2333);
xnor U6845 (N_6845,N_3441,N_4635);
xor U6846 (N_6846,N_3175,N_4504);
xnor U6847 (N_6847,N_3288,N_3993);
or U6848 (N_6848,N_961,N_729);
nor U6849 (N_6849,N_3394,N_4109);
and U6850 (N_6850,N_2716,N_2032);
nand U6851 (N_6851,N_6,N_3707);
nand U6852 (N_6852,N_4143,N_868);
xnor U6853 (N_6853,N_4121,N_180);
nand U6854 (N_6854,N_147,N_2786);
nand U6855 (N_6855,N_4967,N_716);
nand U6856 (N_6856,N_1090,N_3396);
xor U6857 (N_6857,N_1683,N_2088);
or U6858 (N_6858,N_4769,N_2413);
or U6859 (N_6859,N_2202,N_2552);
or U6860 (N_6860,N_1503,N_4981);
xor U6861 (N_6861,N_1902,N_4001);
xnor U6862 (N_6862,N_808,N_960);
nor U6863 (N_6863,N_3776,N_1906);
nand U6864 (N_6864,N_1481,N_3590);
nand U6865 (N_6865,N_3768,N_1978);
nand U6866 (N_6866,N_3588,N_18);
nor U6867 (N_6867,N_1286,N_2558);
xor U6868 (N_6868,N_3748,N_3409);
and U6869 (N_6869,N_4012,N_727);
and U6870 (N_6870,N_3297,N_2323);
nor U6871 (N_6871,N_543,N_4913);
xnor U6872 (N_6872,N_132,N_4199);
xor U6873 (N_6873,N_2563,N_4514);
or U6874 (N_6874,N_1060,N_1840);
xnor U6875 (N_6875,N_3179,N_2091);
nor U6876 (N_6876,N_3222,N_3881);
xnor U6877 (N_6877,N_1268,N_2356);
or U6878 (N_6878,N_880,N_4801);
or U6879 (N_6879,N_4989,N_1234);
and U6880 (N_6880,N_646,N_4110);
nor U6881 (N_6881,N_2790,N_4112);
xnor U6882 (N_6882,N_4972,N_4924);
or U6883 (N_6883,N_4858,N_2754);
xnor U6884 (N_6884,N_4779,N_4938);
nand U6885 (N_6885,N_1461,N_3578);
nand U6886 (N_6886,N_531,N_306);
nor U6887 (N_6887,N_1049,N_873);
xnor U6888 (N_6888,N_3962,N_4255);
or U6889 (N_6889,N_1203,N_1010);
xor U6890 (N_6890,N_4113,N_1833);
or U6891 (N_6891,N_469,N_2872);
xnor U6892 (N_6892,N_3963,N_4862);
xnor U6893 (N_6893,N_3960,N_3238);
xnor U6894 (N_6894,N_4879,N_2677);
or U6895 (N_6895,N_2753,N_1143);
or U6896 (N_6896,N_3109,N_1114);
and U6897 (N_6897,N_731,N_4195);
and U6898 (N_6898,N_4783,N_2501);
and U6899 (N_6899,N_4662,N_1931);
or U6900 (N_6900,N_2652,N_612);
nand U6901 (N_6901,N_677,N_546);
nor U6902 (N_6902,N_3322,N_3700);
and U6903 (N_6903,N_1151,N_2289);
nand U6904 (N_6904,N_4848,N_2755);
nor U6905 (N_6905,N_2578,N_2233);
xnor U6906 (N_6906,N_1233,N_114);
nor U6907 (N_6907,N_3867,N_4331);
or U6908 (N_6908,N_4323,N_445);
nand U6909 (N_6909,N_1365,N_2216);
and U6910 (N_6910,N_4720,N_1862);
nand U6911 (N_6911,N_3636,N_1639);
nand U6912 (N_6912,N_4623,N_4245);
xnor U6913 (N_6913,N_4336,N_2491);
xor U6914 (N_6914,N_153,N_770);
or U6915 (N_6915,N_1544,N_1728);
xnor U6916 (N_6916,N_3949,N_4533);
or U6917 (N_6917,N_1079,N_338);
nor U6918 (N_6918,N_1489,N_3684);
nand U6919 (N_6919,N_3761,N_2607);
nor U6920 (N_6920,N_3313,N_2469);
nand U6921 (N_6921,N_1352,N_619);
nand U6922 (N_6922,N_4627,N_1928);
xor U6923 (N_6923,N_1383,N_4721);
xnor U6924 (N_6924,N_737,N_1410);
nor U6925 (N_6925,N_899,N_3896);
and U6926 (N_6926,N_3071,N_1002);
nor U6927 (N_6927,N_3783,N_2742);
or U6928 (N_6928,N_3217,N_514);
xnor U6929 (N_6929,N_2211,N_3492);
nor U6930 (N_6930,N_4304,N_2099);
xnor U6931 (N_6931,N_2840,N_2029);
nor U6932 (N_6932,N_2053,N_4117);
xnor U6933 (N_6933,N_781,N_1247);
or U6934 (N_6934,N_683,N_305);
nand U6935 (N_6935,N_1186,N_1739);
and U6936 (N_6936,N_504,N_2982);
nand U6937 (N_6937,N_2188,N_3806);
nor U6938 (N_6938,N_3826,N_2474);
and U6939 (N_6939,N_4800,N_3710);
nor U6940 (N_6940,N_4557,N_262);
nand U6941 (N_6941,N_616,N_2060);
xor U6942 (N_6942,N_4665,N_3115);
nor U6943 (N_6943,N_3715,N_3101);
nand U6944 (N_6944,N_847,N_1623);
xnor U6945 (N_6945,N_417,N_3056);
and U6946 (N_6946,N_3572,N_782);
nand U6947 (N_6947,N_4637,N_3379);
nor U6948 (N_6948,N_1222,N_4992);
and U6949 (N_6949,N_4625,N_3756);
xnor U6950 (N_6950,N_2707,N_2721);
nor U6951 (N_6951,N_2533,N_4976);
and U6952 (N_6952,N_1593,N_3295);
nand U6953 (N_6953,N_3317,N_2531);
and U6954 (N_6954,N_544,N_2992);
xor U6955 (N_6955,N_3872,N_4385);
xnor U6956 (N_6956,N_3311,N_2694);
nand U6957 (N_6957,N_2051,N_3390);
nor U6958 (N_6958,N_1487,N_1930);
nand U6959 (N_6959,N_3529,N_2746);
nor U6960 (N_6960,N_4795,N_4279);
xnor U6961 (N_6961,N_260,N_573);
and U6962 (N_6962,N_699,N_2582);
or U6963 (N_6963,N_2522,N_1528);
nor U6964 (N_6964,N_4775,N_460);
nand U6965 (N_6965,N_2106,N_3174);
xor U6966 (N_6966,N_203,N_1926);
and U6967 (N_6967,N_3269,N_2142);
xor U6968 (N_6968,N_1937,N_2926);
xor U6969 (N_6969,N_2506,N_148);
xor U6970 (N_6970,N_1124,N_317);
nor U6971 (N_6971,N_2234,N_2093);
and U6972 (N_6972,N_809,N_4792);
and U6973 (N_6973,N_2195,N_3934);
nand U6974 (N_6974,N_242,N_1749);
or U6975 (N_6975,N_4106,N_1880);
xor U6976 (N_6976,N_3928,N_2798);
nor U6977 (N_6977,N_363,N_3395);
and U6978 (N_6978,N_1959,N_2923);
nand U6979 (N_6979,N_2750,N_3619);
xnor U6980 (N_6980,N_720,N_2230);
xnor U6981 (N_6981,N_133,N_3744);
or U6982 (N_6982,N_4988,N_4103);
or U6983 (N_6983,N_2873,N_4357);
nor U6984 (N_6984,N_4487,N_4036);
and U6985 (N_6985,N_154,N_3797);
and U6986 (N_6986,N_864,N_2568);
and U6987 (N_6987,N_3602,N_4268);
or U6988 (N_6988,N_3878,N_4210);
xnor U6989 (N_6989,N_2059,N_4156);
xnor U6990 (N_6990,N_878,N_3822);
nand U6991 (N_6991,N_915,N_245);
nor U6992 (N_6992,N_4041,N_102);
nand U6993 (N_6993,N_4854,N_406);
nor U6994 (N_6994,N_3025,N_1712);
nor U6995 (N_6995,N_4568,N_315);
nor U6996 (N_6996,N_597,N_4252);
nor U6997 (N_6997,N_1777,N_1385);
nor U6998 (N_6998,N_4539,N_4040);
nor U6999 (N_6999,N_1568,N_755);
or U7000 (N_7000,N_4410,N_3229);
xor U7001 (N_7001,N_3136,N_4716);
xnor U7002 (N_7002,N_408,N_2775);
nor U7003 (N_7003,N_4730,N_724);
or U7004 (N_7004,N_4324,N_4805);
nand U7005 (N_7005,N_3517,N_4136);
xnor U7006 (N_7006,N_2444,N_7);
xnor U7007 (N_7007,N_4488,N_3273);
nand U7008 (N_7008,N_3948,N_45);
nand U7009 (N_7009,N_4028,N_1162);
and U7010 (N_7010,N_20,N_3725);
or U7011 (N_7011,N_4364,N_4292);
xor U7012 (N_7012,N_527,N_1908);
and U7013 (N_7013,N_3885,N_419);
or U7014 (N_7014,N_1339,N_1491);
xnor U7015 (N_7015,N_4959,N_602);
or U7016 (N_7016,N_4960,N_1361);
or U7017 (N_7017,N_1599,N_1119);
nor U7018 (N_7018,N_1290,N_1780);
nor U7019 (N_7019,N_1881,N_1402);
xor U7020 (N_7020,N_1998,N_3887);
and U7021 (N_7021,N_4351,N_2516);
xor U7022 (N_7022,N_4203,N_1132);
nor U7023 (N_7023,N_4482,N_1011);
and U7024 (N_7024,N_4872,N_3610);
or U7025 (N_7025,N_1100,N_595);
and U7026 (N_7026,N_3547,N_1482);
or U7027 (N_7027,N_95,N_2465);
nor U7028 (N_7028,N_2536,N_2660);
xor U7029 (N_7029,N_1159,N_2647);
xnor U7030 (N_7030,N_1462,N_4430);
and U7031 (N_7031,N_4645,N_3124);
nor U7032 (N_7032,N_1292,N_1425);
and U7033 (N_7033,N_2372,N_3371);
nor U7034 (N_7034,N_771,N_4134);
xnor U7035 (N_7035,N_2185,N_2284);
or U7036 (N_7036,N_220,N_4147);
xnor U7037 (N_7037,N_1778,N_259);
or U7038 (N_7038,N_3532,N_2404);
nand U7039 (N_7039,N_2581,N_152);
xor U7040 (N_7040,N_1189,N_3959);
nand U7041 (N_7041,N_3583,N_1171);
nand U7042 (N_7042,N_3182,N_1485);
nand U7043 (N_7043,N_2136,N_966);
nor U7044 (N_7044,N_281,N_3426);
or U7045 (N_7045,N_3903,N_3587);
nand U7046 (N_7046,N_3558,N_131);
nor U7047 (N_7047,N_3059,N_2222);
nor U7048 (N_7048,N_2512,N_671);
nor U7049 (N_7049,N_839,N_1984);
or U7050 (N_7050,N_1947,N_1781);
xor U7051 (N_7051,N_669,N_1483);
or U7052 (N_7052,N_2208,N_3246);
and U7053 (N_7053,N_2555,N_905);
and U7054 (N_7054,N_2606,N_2527);
or U7055 (N_7055,N_1672,N_2466);
nand U7056 (N_7056,N_2368,N_3689);
xnor U7057 (N_7057,N_2306,N_4816);
or U7058 (N_7058,N_2797,N_4837);
or U7059 (N_7059,N_2229,N_2062);
xnor U7060 (N_7060,N_3196,N_3780);
and U7061 (N_7061,N_2275,N_4603);
nor U7062 (N_7062,N_2446,N_410);
nor U7063 (N_7063,N_4841,N_4659);
nand U7064 (N_7064,N_415,N_3152);
nor U7065 (N_7065,N_3037,N_4093);
or U7066 (N_7066,N_3799,N_4375);
nor U7067 (N_7067,N_4408,N_3788);
nand U7068 (N_7068,N_1219,N_2733);
and U7069 (N_7069,N_2069,N_2439);
and U7070 (N_7070,N_2119,N_3090);
nand U7071 (N_7071,N_1806,N_754);
or U7072 (N_7072,N_3559,N_4060);
nand U7073 (N_7073,N_4493,N_2094);
nor U7074 (N_7074,N_4896,N_4751);
nor U7075 (N_7075,N_2779,N_4418);
nand U7076 (N_7076,N_1917,N_857);
nor U7077 (N_7077,N_2973,N_3966);
nand U7078 (N_7078,N_550,N_797);
nand U7079 (N_7079,N_4095,N_3130);
xor U7080 (N_7080,N_4954,N_1144);
nor U7081 (N_7081,N_1792,N_2503);
or U7082 (N_7082,N_3327,N_1064);
or U7083 (N_7083,N_421,N_1828);
nor U7084 (N_7084,N_982,N_3518);
or U7085 (N_7085,N_173,N_1128);
xnor U7086 (N_7086,N_3935,N_4294);
xnor U7087 (N_7087,N_3892,N_4537);
nor U7088 (N_7088,N_4130,N_4690);
nand U7089 (N_7089,N_917,N_1202);
xnor U7090 (N_7090,N_2272,N_26);
nand U7091 (N_7091,N_572,N_2816);
and U7092 (N_7092,N_1116,N_625);
nand U7093 (N_7093,N_499,N_2494);
nor U7094 (N_7094,N_704,N_2292);
and U7095 (N_7095,N_3901,N_2831);
or U7096 (N_7096,N_3466,N_4287);
nor U7097 (N_7097,N_4980,N_3542);
nor U7098 (N_7098,N_1733,N_4144);
nand U7099 (N_7099,N_1574,N_231);
and U7100 (N_7100,N_3105,N_1904);
xor U7101 (N_7101,N_863,N_1697);
nor U7102 (N_7102,N_1624,N_4660);
or U7103 (N_7103,N_2264,N_4939);
nand U7104 (N_7104,N_521,N_4900);
nor U7105 (N_7105,N_68,N_3819);
and U7106 (N_7106,N_962,N_4821);
xnor U7107 (N_7107,N_1849,N_2565);
or U7108 (N_7108,N_1519,N_3805);
xor U7109 (N_7109,N_2920,N_3647);
or U7110 (N_7110,N_2098,N_2519);
and U7111 (N_7111,N_161,N_345);
or U7112 (N_7112,N_2457,N_3637);
xor U7113 (N_7113,N_3670,N_1367);
xor U7114 (N_7114,N_3087,N_3417);
or U7115 (N_7115,N_3296,N_1894);
or U7116 (N_7116,N_4681,N_316);
xor U7117 (N_7117,N_1658,N_4107);
and U7118 (N_7118,N_1898,N_2844);
or U7119 (N_7119,N_3,N_4108);
nand U7120 (N_7120,N_1033,N_4908);
or U7121 (N_7121,N_4275,N_2680);
xor U7122 (N_7122,N_3982,N_3204);
nor U7123 (N_7123,N_1277,N_1814);
nand U7124 (N_7124,N_3911,N_4226);
nand U7125 (N_7125,N_1869,N_1287);
xnor U7126 (N_7126,N_1476,N_641);
or U7127 (N_7127,N_4114,N_3802);
nand U7128 (N_7128,N_3781,N_4796);
xor U7129 (N_7129,N_4605,N_2324);
or U7130 (N_7130,N_4974,N_3916);
xnor U7131 (N_7131,N_2442,N_3391);
nor U7132 (N_7132,N_4675,N_207);
nor U7133 (N_7133,N_911,N_1357);
and U7134 (N_7134,N_1319,N_2504);
xnor U7135 (N_7135,N_1245,N_3728);
and U7136 (N_7136,N_2301,N_4148);
xor U7137 (N_7137,N_1642,N_1876);
nor U7138 (N_7138,N_3681,N_1636);
and U7139 (N_7139,N_4204,N_659);
xnor U7140 (N_7140,N_4663,N_2794);
nand U7141 (N_7141,N_2593,N_4383);
nor U7142 (N_7142,N_1961,N_2396);
xnor U7143 (N_7143,N_1650,N_4765);
and U7144 (N_7144,N_4271,N_3533);
nor U7145 (N_7145,N_2299,N_3361);
or U7146 (N_7146,N_4457,N_4042);
nand U7147 (N_7147,N_3946,N_399);
nor U7148 (N_7148,N_4656,N_4744);
and U7149 (N_7149,N_64,N_2081);
or U7150 (N_7150,N_2295,N_3307);
or U7151 (N_7151,N_509,N_2493);
xor U7152 (N_7152,N_3178,N_4300);
nor U7153 (N_7153,N_2043,N_4387);
or U7154 (N_7154,N_1418,N_359);
nand U7155 (N_7155,N_4454,N_3631);
or U7156 (N_7156,N_3010,N_3747);
or U7157 (N_7157,N_2984,N_4932);
and U7158 (N_7158,N_1356,N_584);
nand U7159 (N_7159,N_2291,N_4995);
nand U7160 (N_7160,N_99,N_3408);
and U7161 (N_7161,N_3132,N_1897);
nor U7162 (N_7162,N_1345,N_2964);
xor U7163 (N_7163,N_1250,N_4748);
nand U7164 (N_7164,N_3874,N_1910);
nor U7165 (N_7165,N_2022,N_368);
nor U7166 (N_7166,N_4548,N_2636);
nor U7167 (N_7167,N_311,N_3494);
and U7168 (N_7168,N_2861,N_3752);
nor U7169 (N_7169,N_1388,N_327);
nand U7170 (N_7170,N_2592,N_3073);
nor U7171 (N_7171,N_4903,N_4133);
or U7172 (N_7172,N_4228,N_1886);
or U7173 (N_7173,N_4221,N_1617);
xnor U7174 (N_7174,N_418,N_2788);
or U7175 (N_7175,N_4619,N_4015);
nor U7176 (N_7176,N_4402,N_4834);
xor U7177 (N_7177,N_2017,N_4601);
and U7178 (N_7178,N_3810,N_851);
nand U7179 (N_7179,N_3249,N_967);
nor U7180 (N_7180,N_3625,N_2016);
and U7181 (N_7181,N_230,N_494);
xor U7182 (N_7182,N_348,N_36);
nor U7183 (N_7183,N_4506,N_4476);
nor U7184 (N_7184,N_4473,N_1038);
or U7185 (N_7185,N_695,N_1549);
nor U7186 (N_7186,N_1845,N_2732);
nor U7187 (N_7187,N_1979,N_3544);
xnor U7188 (N_7188,N_4415,N_3554);
or U7189 (N_7189,N_4767,N_4986);
xor U7190 (N_7190,N_3163,N_70);
or U7191 (N_7191,N_2328,N_4253);
and U7192 (N_7192,N_407,N_959);
or U7193 (N_7193,N_1824,N_3251);
nor U7194 (N_7194,N_2922,N_2758);
and U7195 (N_7195,N_2077,N_3839);
nor U7196 (N_7196,N_4592,N_4419);
xnor U7197 (N_7197,N_2822,N_4772);
xor U7198 (N_7198,N_2572,N_2181);
or U7199 (N_7199,N_2567,N_4874);
xor U7200 (N_7200,N_2528,N_151);
or U7201 (N_7201,N_4008,N_189);
nor U7202 (N_7202,N_472,N_2116);
xor U7203 (N_7203,N_3169,N_3815);
and U7204 (N_7204,N_2278,N_2962);
or U7205 (N_7205,N_2002,N_71);
and U7206 (N_7206,N_533,N_140);
xnor U7207 (N_7207,N_4154,N_3122);
xnor U7208 (N_7208,N_4717,N_3734);
nand U7209 (N_7209,N_372,N_2483);
and U7210 (N_7210,N_2713,N_4283);
xor U7211 (N_7211,N_3081,N_969);
nor U7212 (N_7212,N_1946,N_3821);
and U7213 (N_7213,N_1775,N_1943);
nand U7214 (N_7214,N_4513,N_779);
nor U7215 (N_7215,N_3168,N_972);
nand U7216 (N_7216,N_4888,N_2489);
or U7217 (N_7217,N_525,N_3914);
xor U7218 (N_7218,N_3149,N_2837);
nor U7219 (N_7219,N_2781,N_2398);
or U7220 (N_7220,N_3088,N_75);
xor U7221 (N_7221,N_952,N_3674);
and U7222 (N_7222,N_2544,N_2415);
xor U7223 (N_7223,N_2509,N_43);
xnor U7224 (N_7224,N_2631,N_582);
and U7225 (N_7225,N_1232,N_3571);
and U7226 (N_7226,N_3793,N_4374);
or U7227 (N_7227,N_796,N_1449);
nand U7228 (N_7228,N_3474,N_4595);
and U7229 (N_7229,N_1059,N_85);
or U7230 (N_7230,N_2997,N_2261);
nor U7231 (N_7231,N_603,N_354);
and U7232 (N_7232,N_4749,N_3675);
xnor U7233 (N_7233,N_4016,N_497);
nor U7234 (N_7234,N_229,N_4593);
nand U7235 (N_7235,N_343,N_3830);
nor U7236 (N_7236,N_3475,N_1541);
nor U7237 (N_7237,N_4178,N_3974);
nor U7238 (N_7238,N_555,N_657);
or U7239 (N_7239,N_2619,N_170);
nor U7240 (N_7240,N_4474,N_4219);
and U7241 (N_7241,N_1267,N_4781);
or U7242 (N_7242,N_202,N_4378);
xnor U7243 (N_7243,N_2877,N_698);
xnor U7244 (N_7244,N_3338,N_2931);
and U7245 (N_7245,N_3739,N_2971);
nand U7246 (N_7246,N_2386,N_883);
nor U7247 (N_7247,N_4356,N_1938);
nand U7248 (N_7248,N_3730,N_3369);
and U7249 (N_7249,N_4560,N_3641);
nor U7250 (N_7250,N_4550,N_3973);
and U7251 (N_7251,N_356,N_1843);
xor U7252 (N_7252,N_416,N_4303);
or U7253 (N_7253,N_916,N_4596);
nor U7254 (N_7254,N_2701,N_2481);
or U7255 (N_7255,N_1206,N_2403);
nand U7256 (N_7256,N_4389,N_1705);
nor U7257 (N_7257,N_2654,N_2319);
and U7258 (N_7258,N_608,N_1884);
xor U7259 (N_7259,N_4736,N_2905);
and U7260 (N_7260,N_4317,N_4301);
and U7261 (N_7261,N_4420,N_1364);
or U7262 (N_7262,N_1940,N_1838);
nor U7263 (N_7263,N_3640,N_4832);
nand U7264 (N_7264,N_3199,N_2343);
nor U7265 (N_7265,N_4333,N_1835);
and U7266 (N_7266,N_3856,N_845);
xnor U7267 (N_7267,N_414,N_3051);
xnor U7268 (N_7268,N_872,N_3445);
nor U7269 (N_7269,N_1317,N_2238);
xor U7270 (N_7270,N_2443,N_2723);
or U7271 (N_7271,N_1451,N_2424);
xnor U7272 (N_7272,N_62,N_4084);
nor U7273 (N_7273,N_1810,N_2332);
and U7274 (N_7274,N_2776,N_4711);
and U7275 (N_7275,N_2547,N_4674);
and U7276 (N_7276,N_2911,N_2938);
or U7277 (N_7277,N_3242,N_346);
and U7278 (N_7278,N_4298,N_2599);
nand U7279 (N_7279,N_2841,N_4302);
and U7280 (N_7280,N_341,N_4120);
or U7281 (N_7281,N_803,N_2613);
xor U7282 (N_7282,N_3548,N_4551);
xor U7283 (N_7283,N_4670,N_2869);
or U7284 (N_7284,N_4901,N_3410);
and U7285 (N_7285,N_4305,N_762);
or U7286 (N_7286,N_3555,N_2739);
nor U7287 (N_7287,N_391,N_3389);
nor U7288 (N_7288,N_4166,N_3353);
nor U7289 (N_7289,N_400,N_673);
and U7290 (N_7290,N_4962,N_604);
nand U7291 (N_7291,N_4235,N_4187);
or U7292 (N_7292,N_2127,N_3923);
nor U7293 (N_7293,N_3325,N_4649);
and U7294 (N_7294,N_2735,N_1718);
nor U7295 (N_7295,N_4447,N_2793);
or U7296 (N_7296,N_3868,N_4510);
and U7297 (N_7297,N_3358,N_2740);
xnor U7298 (N_7298,N_19,N_3312);
or U7299 (N_7299,N_4525,N_3117);
or U7300 (N_7300,N_3697,N_2008);
or U7301 (N_7301,N_4310,N_2675);
nand U7302 (N_7302,N_80,N_4381);
or U7303 (N_7303,N_1480,N_3726);
xnor U7304 (N_7304,N_564,N_1557);
or U7305 (N_7305,N_3906,N_4097);
and U7306 (N_7306,N_4511,N_4254);
xnor U7307 (N_7307,N_307,N_1018);
or U7308 (N_7308,N_706,N_3015);
xnor U7309 (N_7309,N_388,N_1929);
nand U7310 (N_7310,N_4762,N_4017);
and U7311 (N_7311,N_2618,N_4152);
nand U7312 (N_7312,N_105,N_3576);
xor U7313 (N_7313,N_837,N_2151);
nand U7314 (N_7314,N_4358,N_463);
and U7315 (N_7315,N_1540,N_1533);
or U7316 (N_7316,N_4022,N_2774);
xnor U7317 (N_7317,N_557,N_174);
nor U7318 (N_7318,N_1668,N_2814);
nor U7319 (N_7319,N_3455,N_2553);
xnor U7320 (N_7320,N_2325,N_4362);
and U7321 (N_7321,N_135,N_3778);
or U7322 (N_7322,N_2601,N_4215);
xor U7323 (N_7323,N_1896,N_1714);
xnor U7324 (N_7324,N_3008,N_375);
or U7325 (N_7325,N_3762,N_1964);
and U7326 (N_7326,N_2400,N_3233);
nand U7327 (N_7327,N_2305,N_3520);
or U7328 (N_7328,N_3665,N_4439);
nand U7329 (N_7329,N_949,N_3016);
or U7330 (N_7330,N_383,N_1945);
nor U7331 (N_7331,N_4377,N_461);
and U7332 (N_7332,N_2144,N_3098);
or U7333 (N_7333,N_3339,N_505);
and U7334 (N_7334,N_1991,N_1417);
nand U7335 (N_7335,N_1315,N_2355);
nor U7336 (N_7336,N_1376,N_1054);
nor U7337 (N_7337,N_3365,N_3757);
and U7338 (N_7338,N_1344,N_1221);
xnor U7339 (N_7339,N_2727,N_2063);
or U7340 (N_7340,N_2224,N_848);
or U7341 (N_7341,N_668,N_2805);
or U7342 (N_7342,N_3113,N_2829);
and U7343 (N_7343,N_4481,N_1276);
and U7344 (N_7344,N_2684,N_2809);
nand U7345 (N_7345,N_4847,N_4397);
nand U7346 (N_7346,N_1393,N_856);
xnor U7347 (N_7347,N_2166,N_1153);
nor U7348 (N_7348,N_4319,N_3895);
and U7349 (N_7349,N_575,N_1404);
or U7350 (N_7350,N_3316,N_2823);
xnor U7351 (N_7351,N_2364,N_2108);
xor U7352 (N_7352,N_3764,N_1988);
nor U7353 (N_7353,N_703,N_583);
xnor U7354 (N_7354,N_1426,N_1381);
nand U7355 (N_7355,N_4724,N_358);
and U7356 (N_7356,N_2279,N_4617);
or U7357 (N_7357,N_1976,N_1057);
nor U7358 (N_7358,N_1995,N_553);
xor U7359 (N_7359,N_2769,N_4464);
xnor U7360 (N_7360,N_1490,N_999);
nand U7361 (N_7361,N_2978,N_4984);
or U7362 (N_7362,N_1251,N_1325);
or U7363 (N_7363,N_35,N_3593);
nor U7364 (N_7364,N_3184,N_4018);
xor U7365 (N_7365,N_163,N_3809);
and U7366 (N_7366,N_2174,N_3437);
xor U7367 (N_7367,N_3888,N_1804);
xor U7368 (N_7368,N_4453,N_4023);
xor U7369 (N_7369,N_3575,N_145);
nor U7370 (N_7370,N_4544,N_78);
nor U7371 (N_7371,N_1168,N_3093);
xor U7372 (N_7372,N_3970,N_2471);
nand U7373 (N_7373,N_1891,N_4668);
nand U7374 (N_7374,N_1807,N_2966);
xnor U7375 (N_7375,N_1513,N_218);
nand U7376 (N_7376,N_190,N_385);
and U7377 (N_7377,N_1618,N_1577);
nor U7378 (N_7378,N_1716,N_3932);
xor U7379 (N_7379,N_2455,N_1110);
and U7380 (N_7380,N_1099,N_4327);
nor U7381 (N_7381,N_957,N_976);
xnor U7382 (N_7382,N_3340,N_3022);
nand U7383 (N_7383,N_4379,N_3470);
nand U7384 (N_7384,N_3604,N_542);
or U7385 (N_7385,N_3362,N_2957);
or U7386 (N_7386,N_3218,N_2712);
nand U7387 (N_7387,N_108,N_4884);
nor U7388 (N_7388,N_3278,N_2201);
nor U7389 (N_7389,N_1692,N_4773);
nand U7390 (N_7390,N_4861,N_2409);
nor U7391 (N_7391,N_115,N_169);
xor U7392 (N_7392,N_524,N_3486);
and U7393 (N_7393,N_184,N_4820);
or U7394 (N_7394,N_1009,N_4630);
or U7395 (N_7395,N_4404,N_2597);
nor U7396 (N_7396,N_2611,N_1985);
nand U7397 (N_7397,N_923,N_3943);
and U7398 (N_7398,N_4629,N_2078);
or U7399 (N_7399,N_434,N_888);
nor U7400 (N_7400,N_405,N_2235);
and U7401 (N_7401,N_22,N_1863);
nor U7402 (N_7402,N_3562,N_4911);
nand U7403 (N_7403,N_1699,N_3933);
and U7404 (N_7404,N_2007,N_4902);
or U7405 (N_7405,N_440,N_1291);
nor U7406 (N_7406,N_2237,N_3638);
nand U7407 (N_7407,N_733,N_4729);
and U7408 (N_7408,N_1109,N_1134);
or U7409 (N_7409,N_2627,N_4530);
and U7410 (N_7410,N_3049,N_2849);
and U7411 (N_7411,N_4700,N_3240);
nor U7412 (N_7412,N_196,N_479);
or U7413 (N_7413,N_4461,N_3877);
or U7414 (N_7414,N_4891,N_3155);
nor U7415 (N_7415,N_2643,N_717);
and U7416 (N_7416,N_1438,N_996);
nand U7417 (N_7417,N_3882,N_517);
and U7418 (N_7418,N_2320,N_1779);
xnor U7419 (N_7419,N_2039,N_4935);
or U7420 (N_7420,N_567,N_3300);
xor U7421 (N_7421,N_1925,N_3836);
nor U7422 (N_7422,N_3855,N_1501);
and U7423 (N_7423,N_1788,N_831);
and U7424 (N_7424,N_3727,N_4483);
xnor U7425 (N_7425,N_507,N_3563);
xnor U7426 (N_7426,N_4280,N_3909);
xor U7427 (N_7427,N_2005,N_1531);
nand U7428 (N_7428,N_3907,N_1818);
xor U7429 (N_7429,N_885,N_1537);
nand U7430 (N_7430,N_2561,N_3141);
xor U7431 (N_7431,N_4009,N_1837);
and U7432 (N_7432,N_3058,N_858);
or U7433 (N_7433,N_139,N_822);
and U7434 (N_7434,N_2322,N_3945);
nor U7435 (N_7435,N_1953,N_1510);
and U7436 (N_7436,N_3737,N_4709);
nor U7437 (N_7437,N_3106,N_4822);
xnor U7438 (N_7438,N_977,N_2276);
or U7439 (N_7439,N_4353,N_446);
xnor U7440 (N_7440,N_4125,N_4400);
xor U7441 (N_7441,N_1297,N_4384);
nor U7442 (N_7442,N_1601,N_3171);
xnor U7443 (N_7443,N_2602,N_4085);
or U7444 (N_7444,N_4607,N_2085);
nand U7445 (N_7445,N_4376,N_351);
and U7446 (N_7446,N_1260,N_2896);
and U7447 (N_7447,N_175,N_4484);
nand U7448 (N_7448,N_1169,N_739);
nand U7449 (N_7449,N_710,N_3720);
nor U7450 (N_7450,N_3487,N_4135);
and U7451 (N_7451,N_742,N_632);
xnor U7452 (N_7452,N_1764,N_4646);
xor U7453 (N_7453,N_1166,N_165);
and U7454 (N_7454,N_927,N_2893);
nor U7455 (N_7455,N_1475,N_2588);
and U7456 (N_7456,N_367,N_285);
nand U7457 (N_7457,N_2616,N_780);
nand U7458 (N_7458,N_4192,N_633);
nor U7459 (N_7459,N_3219,N_3866);
or U7460 (N_7460,N_4520,N_253);
nand U7461 (N_7461,N_895,N_295);
or U7462 (N_7462,N_4621,N_3566);
nand U7463 (N_7463,N_3808,N_3803);
nand U7464 (N_7464,N_2574,N_107);
nor U7465 (N_7465,N_467,N_630);
nor U7466 (N_7466,N_4685,N_1496);
or U7467 (N_7467,N_4814,N_4941);
nor U7468 (N_7468,N_2040,N_2683);
or U7469 (N_7469,N_2756,N_1308);
or U7470 (N_7470,N_2381,N_1197);
xor U7471 (N_7471,N_1682,N_4243);
or U7472 (N_7472,N_3308,N_3837);
nand U7473 (N_7473,N_2669,N_3864);
and U7474 (N_7474,N_3407,N_347);
or U7475 (N_7475,N_2990,N_2021);
and U7476 (N_7476,N_3045,N_2678);
nand U7477 (N_7477,N_2839,N_2972);
or U7478 (N_7478,N_3996,N_1177);
nor U7479 (N_7479,N_2934,N_1004);
nand U7480 (N_7480,N_2219,N_4644);
nor U7481 (N_7481,N_918,N_664);
or U7482 (N_7482,N_965,N_1628);
and U7483 (N_7483,N_2199,N_1265);
nand U7484 (N_7484,N_2121,N_2414);
xnor U7485 (N_7485,N_4315,N_662);
or U7486 (N_7486,N_3843,N_3519);
nand U7487 (N_7487,N_136,N_655);
xor U7488 (N_7488,N_4455,N_1954);
xor U7489 (N_7489,N_52,N_44);
nand U7490 (N_7490,N_1332,N_3166);
or U7491 (N_7491,N_1095,N_4706);
nand U7492 (N_7492,N_2459,N_882);
nand U7493 (N_7493,N_2830,N_1695);
nand U7494 (N_7494,N_3804,N_2628);
or U7495 (N_7495,N_4449,N_503);
and U7496 (N_7496,N_3721,N_2693);
nor U7497 (N_7497,N_1324,N_2154);
and U7498 (N_7498,N_2824,N_3286);
nand U7499 (N_7499,N_470,N_3676);
and U7500 (N_7500,N_543,N_1611);
and U7501 (N_7501,N_2735,N_3285);
nand U7502 (N_7502,N_3001,N_3897);
nor U7503 (N_7503,N_2156,N_1847);
and U7504 (N_7504,N_3124,N_1863);
nor U7505 (N_7505,N_767,N_1061);
or U7506 (N_7506,N_539,N_3);
nor U7507 (N_7507,N_1775,N_2925);
and U7508 (N_7508,N_1300,N_3577);
xor U7509 (N_7509,N_252,N_4360);
and U7510 (N_7510,N_1414,N_2298);
xor U7511 (N_7511,N_1054,N_3519);
xor U7512 (N_7512,N_3736,N_2668);
nand U7513 (N_7513,N_4874,N_3170);
xnor U7514 (N_7514,N_2988,N_1489);
and U7515 (N_7515,N_399,N_1624);
or U7516 (N_7516,N_281,N_2621);
nand U7517 (N_7517,N_667,N_182);
nor U7518 (N_7518,N_2336,N_4596);
nor U7519 (N_7519,N_1120,N_2546);
or U7520 (N_7520,N_879,N_2496);
or U7521 (N_7521,N_2024,N_3849);
nor U7522 (N_7522,N_4412,N_1323);
and U7523 (N_7523,N_2383,N_2838);
nor U7524 (N_7524,N_185,N_1055);
and U7525 (N_7525,N_4171,N_3656);
nor U7526 (N_7526,N_772,N_4221);
nor U7527 (N_7527,N_3307,N_2660);
or U7528 (N_7528,N_4036,N_2337);
xnor U7529 (N_7529,N_2069,N_3454);
nand U7530 (N_7530,N_2914,N_650);
nand U7531 (N_7531,N_4698,N_1907);
nor U7532 (N_7532,N_3067,N_2337);
and U7533 (N_7533,N_4046,N_379);
or U7534 (N_7534,N_4133,N_1720);
or U7535 (N_7535,N_3567,N_318);
xor U7536 (N_7536,N_1728,N_3486);
or U7537 (N_7537,N_2623,N_2113);
and U7538 (N_7538,N_1442,N_4137);
or U7539 (N_7539,N_57,N_3077);
xor U7540 (N_7540,N_4177,N_1821);
xor U7541 (N_7541,N_1677,N_391);
and U7542 (N_7542,N_4601,N_2630);
nor U7543 (N_7543,N_4339,N_853);
and U7544 (N_7544,N_1159,N_2300);
and U7545 (N_7545,N_1110,N_2669);
nor U7546 (N_7546,N_2577,N_2891);
and U7547 (N_7547,N_883,N_2949);
xnor U7548 (N_7548,N_45,N_1570);
or U7549 (N_7549,N_4429,N_3427);
nand U7550 (N_7550,N_4208,N_2565);
or U7551 (N_7551,N_868,N_572);
or U7552 (N_7552,N_4221,N_1117);
xnor U7553 (N_7553,N_1837,N_3267);
xor U7554 (N_7554,N_4902,N_1634);
nand U7555 (N_7555,N_2332,N_1715);
nand U7556 (N_7556,N_4054,N_510);
xor U7557 (N_7557,N_997,N_1519);
nand U7558 (N_7558,N_4986,N_2212);
and U7559 (N_7559,N_2260,N_1816);
nor U7560 (N_7560,N_4448,N_2326);
nor U7561 (N_7561,N_229,N_2042);
and U7562 (N_7562,N_4319,N_2716);
or U7563 (N_7563,N_679,N_4112);
or U7564 (N_7564,N_1321,N_416);
or U7565 (N_7565,N_1339,N_1994);
xor U7566 (N_7566,N_4582,N_3778);
and U7567 (N_7567,N_2703,N_1002);
nor U7568 (N_7568,N_4130,N_418);
xnor U7569 (N_7569,N_671,N_149);
nand U7570 (N_7570,N_2555,N_1778);
nand U7571 (N_7571,N_3419,N_3940);
xnor U7572 (N_7572,N_4153,N_4229);
nand U7573 (N_7573,N_2956,N_2022);
and U7574 (N_7574,N_2354,N_3085);
and U7575 (N_7575,N_197,N_3825);
or U7576 (N_7576,N_2004,N_968);
xnor U7577 (N_7577,N_209,N_4870);
xor U7578 (N_7578,N_465,N_17);
nor U7579 (N_7579,N_4142,N_3230);
and U7580 (N_7580,N_3833,N_1963);
nor U7581 (N_7581,N_2871,N_626);
or U7582 (N_7582,N_3435,N_3592);
nand U7583 (N_7583,N_1575,N_4247);
or U7584 (N_7584,N_3092,N_645);
xnor U7585 (N_7585,N_3683,N_3837);
xnor U7586 (N_7586,N_4916,N_1798);
and U7587 (N_7587,N_4329,N_1027);
or U7588 (N_7588,N_4667,N_4301);
or U7589 (N_7589,N_2917,N_1817);
and U7590 (N_7590,N_3728,N_2366);
and U7591 (N_7591,N_4672,N_2443);
nor U7592 (N_7592,N_2592,N_2493);
nand U7593 (N_7593,N_1011,N_900);
nor U7594 (N_7594,N_2896,N_387);
nor U7595 (N_7595,N_555,N_4851);
and U7596 (N_7596,N_785,N_2998);
and U7597 (N_7597,N_518,N_1408);
nand U7598 (N_7598,N_4476,N_2754);
nand U7599 (N_7599,N_1837,N_3113);
and U7600 (N_7600,N_3163,N_3137);
or U7601 (N_7601,N_1450,N_1780);
nor U7602 (N_7602,N_539,N_3320);
nor U7603 (N_7603,N_2959,N_796);
xnor U7604 (N_7604,N_1417,N_4386);
xnor U7605 (N_7605,N_3996,N_4394);
nand U7606 (N_7606,N_1506,N_3627);
and U7607 (N_7607,N_4202,N_3868);
nand U7608 (N_7608,N_4093,N_2219);
or U7609 (N_7609,N_3648,N_2695);
nand U7610 (N_7610,N_4768,N_1202);
nand U7611 (N_7611,N_1543,N_2330);
xor U7612 (N_7612,N_4103,N_3727);
nand U7613 (N_7613,N_2790,N_531);
xnor U7614 (N_7614,N_4047,N_3698);
and U7615 (N_7615,N_2599,N_2891);
and U7616 (N_7616,N_3670,N_2426);
or U7617 (N_7617,N_4239,N_198);
nor U7618 (N_7618,N_1494,N_2343);
nand U7619 (N_7619,N_4378,N_3320);
and U7620 (N_7620,N_108,N_2290);
and U7621 (N_7621,N_4704,N_633);
or U7622 (N_7622,N_343,N_176);
and U7623 (N_7623,N_4235,N_3212);
nand U7624 (N_7624,N_798,N_2192);
xnor U7625 (N_7625,N_1904,N_2546);
and U7626 (N_7626,N_4050,N_4775);
and U7627 (N_7627,N_4412,N_3301);
and U7628 (N_7628,N_3387,N_4533);
xnor U7629 (N_7629,N_1339,N_1020);
nor U7630 (N_7630,N_3075,N_4966);
or U7631 (N_7631,N_1921,N_51);
nor U7632 (N_7632,N_4250,N_2318);
and U7633 (N_7633,N_652,N_748);
nor U7634 (N_7634,N_2957,N_3345);
nor U7635 (N_7635,N_493,N_3077);
or U7636 (N_7636,N_4570,N_2281);
nand U7637 (N_7637,N_2397,N_2865);
nor U7638 (N_7638,N_3710,N_3594);
or U7639 (N_7639,N_2893,N_4953);
or U7640 (N_7640,N_4174,N_1574);
xor U7641 (N_7641,N_4909,N_3417);
nor U7642 (N_7642,N_96,N_948);
and U7643 (N_7643,N_3992,N_4337);
nand U7644 (N_7644,N_1989,N_4842);
nor U7645 (N_7645,N_123,N_4404);
nor U7646 (N_7646,N_2493,N_2164);
xor U7647 (N_7647,N_869,N_2862);
and U7648 (N_7648,N_2446,N_1318);
nand U7649 (N_7649,N_773,N_3876);
xnor U7650 (N_7650,N_4187,N_2925);
xor U7651 (N_7651,N_2662,N_2888);
nor U7652 (N_7652,N_908,N_2709);
or U7653 (N_7653,N_233,N_4333);
nand U7654 (N_7654,N_2316,N_4283);
or U7655 (N_7655,N_254,N_3984);
nor U7656 (N_7656,N_380,N_2676);
or U7657 (N_7657,N_2291,N_2067);
xnor U7658 (N_7658,N_2484,N_3362);
nor U7659 (N_7659,N_3562,N_455);
and U7660 (N_7660,N_3117,N_702);
and U7661 (N_7661,N_3626,N_3420);
or U7662 (N_7662,N_172,N_467);
nor U7663 (N_7663,N_693,N_2217);
nand U7664 (N_7664,N_1695,N_4381);
nand U7665 (N_7665,N_4487,N_365);
and U7666 (N_7666,N_4353,N_506);
and U7667 (N_7667,N_1929,N_4872);
xnor U7668 (N_7668,N_4350,N_4160);
nor U7669 (N_7669,N_4461,N_4742);
xor U7670 (N_7670,N_1636,N_4718);
nand U7671 (N_7671,N_3852,N_1276);
or U7672 (N_7672,N_3208,N_2214);
nand U7673 (N_7673,N_735,N_293);
xor U7674 (N_7674,N_499,N_2506);
or U7675 (N_7675,N_4929,N_4117);
or U7676 (N_7676,N_2438,N_4137);
and U7677 (N_7677,N_409,N_1798);
and U7678 (N_7678,N_618,N_2372);
nand U7679 (N_7679,N_3371,N_3683);
and U7680 (N_7680,N_186,N_299);
or U7681 (N_7681,N_3376,N_1266);
nor U7682 (N_7682,N_1245,N_2417);
nand U7683 (N_7683,N_4096,N_1982);
xnor U7684 (N_7684,N_4813,N_432);
nand U7685 (N_7685,N_366,N_1302);
nor U7686 (N_7686,N_1918,N_1066);
and U7687 (N_7687,N_400,N_4973);
nand U7688 (N_7688,N_4219,N_4635);
or U7689 (N_7689,N_4740,N_327);
xor U7690 (N_7690,N_2212,N_4523);
xor U7691 (N_7691,N_2780,N_99);
nand U7692 (N_7692,N_914,N_3139);
nand U7693 (N_7693,N_449,N_1409);
or U7694 (N_7694,N_3168,N_4221);
and U7695 (N_7695,N_4655,N_3618);
nor U7696 (N_7696,N_1917,N_157);
and U7697 (N_7697,N_3404,N_913);
or U7698 (N_7698,N_1197,N_4065);
nand U7699 (N_7699,N_2353,N_4720);
xnor U7700 (N_7700,N_35,N_676);
and U7701 (N_7701,N_1181,N_4720);
or U7702 (N_7702,N_4107,N_4801);
and U7703 (N_7703,N_4324,N_2733);
or U7704 (N_7704,N_3354,N_2181);
nor U7705 (N_7705,N_992,N_3439);
xnor U7706 (N_7706,N_1772,N_2689);
nor U7707 (N_7707,N_3713,N_3502);
xor U7708 (N_7708,N_220,N_4653);
and U7709 (N_7709,N_672,N_2105);
nor U7710 (N_7710,N_51,N_2655);
or U7711 (N_7711,N_1080,N_830);
and U7712 (N_7712,N_3713,N_4842);
nand U7713 (N_7713,N_3566,N_1584);
and U7714 (N_7714,N_1462,N_1816);
or U7715 (N_7715,N_130,N_709);
and U7716 (N_7716,N_3254,N_2844);
and U7717 (N_7717,N_2712,N_345);
nor U7718 (N_7718,N_3263,N_1768);
and U7719 (N_7719,N_1446,N_4);
nand U7720 (N_7720,N_1957,N_1054);
nand U7721 (N_7721,N_1672,N_3254);
and U7722 (N_7722,N_4677,N_2884);
nor U7723 (N_7723,N_4547,N_1060);
and U7724 (N_7724,N_961,N_1182);
or U7725 (N_7725,N_1060,N_115);
xor U7726 (N_7726,N_4251,N_1102);
nand U7727 (N_7727,N_1537,N_1660);
nand U7728 (N_7728,N_3773,N_4862);
nand U7729 (N_7729,N_1016,N_4928);
or U7730 (N_7730,N_2350,N_3705);
and U7731 (N_7731,N_3906,N_3791);
nor U7732 (N_7732,N_3929,N_2642);
or U7733 (N_7733,N_3812,N_2906);
or U7734 (N_7734,N_4160,N_3117);
nor U7735 (N_7735,N_2934,N_4297);
xor U7736 (N_7736,N_3863,N_1086);
nand U7737 (N_7737,N_4208,N_2475);
nand U7738 (N_7738,N_1384,N_2958);
xnor U7739 (N_7739,N_1423,N_1709);
and U7740 (N_7740,N_4822,N_441);
nand U7741 (N_7741,N_573,N_1257);
or U7742 (N_7742,N_4997,N_4600);
and U7743 (N_7743,N_3906,N_3482);
and U7744 (N_7744,N_1974,N_3378);
nor U7745 (N_7745,N_3757,N_3468);
xor U7746 (N_7746,N_650,N_4107);
or U7747 (N_7747,N_3526,N_4297);
and U7748 (N_7748,N_1919,N_2590);
nor U7749 (N_7749,N_3063,N_3672);
or U7750 (N_7750,N_2,N_4165);
and U7751 (N_7751,N_1587,N_3559);
xnor U7752 (N_7752,N_1901,N_3669);
and U7753 (N_7753,N_3262,N_2899);
or U7754 (N_7754,N_4235,N_4160);
or U7755 (N_7755,N_1612,N_3295);
nand U7756 (N_7756,N_4814,N_2047);
or U7757 (N_7757,N_4463,N_4451);
nand U7758 (N_7758,N_1607,N_3770);
or U7759 (N_7759,N_4817,N_3674);
and U7760 (N_7760,N_2069,N_3034);
xor U7761 (N_7761,N_4310,N_1496);
and U7762 (N_7762,N_783,N_4362);
or U7763 (N_7763,N_1751,N_1168);
xnor U7764 (N_7764,N_4014,N_1772);
nand U7765 (N_7765,N_4339,N_1712);
nor U7766 (N_7766,N_2295,N_2381);
or U7767 (N_7767,N_3613,N_580);
xor U7768 (N_7768,N_3824,N_977);
nand U7769 (N_7769,N_4863,N_2424);
nor U7770 (N_7770,N_1256,N_1091);
and U7771 (N_7771,N_1199,N_3486);
nand U7772 (N_7772,N_998,N_564);
or U7773 (N_7773,N_3932,N_1336);
xnor U7774 (N_7774,N_693,N_716);
and U7775 (N_7775,N_3572,N_1081);
nor U7776 (N_7776,N_514,N_2940);
or U7777 (N_7777,N_2042,N_3401);
nor U7778 (N_7778,N_2803,N_3786);
xor U7779 (N_7779,N_3228,N_1015);
or U7780 (N_7780,N_1465,N_494);
and U7781 (N_7781,N_2193,N_660);
xor U7782 (N_7782,N_219,N_658);
or U7783 (N_7783,N_493,N_3097);
xnor U7784 (N_7784,N_4370,N_644);
nor U7785 (N_7785,N_1528,N_3924);
and U7786 (N_7786,N_2541,N_516);
xor U7787 (N_7787,N_3886,N_3327);
nand U7788 (N_7788,N_822,N_3145);
nor U7789 (N_7789,N_3816,N_1912);
xnor U7790 (N_7790,N_1111,N_1604);
xnor U7791 (N_7791,N_2434,N_2900);
and U7792 (N_7792,N_4461,N_4050);
xnor U7793 (N_7793,N_585,N_1733);
nor U7794 (N_7794,N_3636,N_794);
nor U7795 (N_7795,N_1632,N_3241);
nand U7796 (N_7796,N_4000,N_4433);
nor U7797 (N_7797,N_2786,N_2577);
nor U7798 (N_7798,N_4606,N_4920);
nand U7799 (N_7799,N_4440,N_4051);
and U7800 (N_7800,N_2500,N_3115);
nand U7801 (N_7801,N_3698,N_4881);
and U7802 (N_7802,N_2337,N_4307);
nand U7803 (N_7803,N_31,N_4378);
nor U7804 (N_7804,N_61,N_3321);
nand U7805 (N_7805,N_3066,N_75);
nor U7806 (N_7806,N_1125,N_3859);
xnor U7807 (N_7807,N_697,N_3101);
nand U7808 (N_7808,N_3744,N_1943);
nor U7809 (N_7809,N_2087,N_2160);
and U7810 (N_7810,N_4212,N_3605);
nand U7811 (N_7811,N_2208,N_3326);
nand U7812 (N_7812,N_1337,N_4219);
nand U7813 (N_7813,N_1859,N_4712);
nor U7814 (N_7814,N_3985,N_742);
nand U7815 (N_7815,N_2172,N_3090);
xor U7816 (N_7816,N_637,N_3415);
nor U7817 (N_7817,N_1877,N_400);
xnor U7818 (N_7818,N_1069,N_353);
nor U7819 (N_7819,N_2303,N_4103);
or U7820 (N_7820,N_4664,N_287);
xnor U7821 (N_7821,N_4921,N_2404);
nand U7822 (N_7822,N_4374,N_4004);
xnor U7823 (N_7823,N_576,N_4789);
and U7824 (N_7824,N_4761,N_487);
and U7825 (N_7825,N_1735,N_4949);
nand U7826 (N_7826,N_1020,N_4248);
nor U7827 (N_7827,N_1332,N_2314);
or U7828 (N_7828,N_1645,N_3906);
nor U7829 (N_7829,N_3255,N_928);
nand U7830 (N_7830,N_4580,N_3071);
and U7831 (N_7831,N_2009,N_4664);
and U7832 (N_7832,N_2565,N_4479);
and U7833 (N_7833,N_2358,N_4463);
xor U7834 (N_7834,N_2858,N_4389);
and U7835 (N_7835,N_3090,N_2853);
nor U7836 (N_7836,N_1237,N_1220);
xor U7837 (N_7837,N_4526,N_2608);
xor U7838 (N_7838,N_3648,N_3790);
or U7839 (N_7839,N_2933,N_2844);
and U7840 (N_7840,N_379,N_3826);
xnor U7841 (N_7841,N_775,N_154);
nand U7842 (N_7842,N_3785,N_2832);
xor U7843 (N_7843,N_193,N_2220);
or U7844 (N_7844,N_1042,N_4752);
or U7845 (N_7845,N_2631,N_1353);
or U7846 (N_7846,N_3985,N_3215);
nor U7847 (N_7847,N_1487,N_1725);
nor U7848 (N_7848,N_390,N_1840);
xor U7849 (N_7849,N_3212,N_3724);
nand U7850 (N_7850,N_4920,N_2580);
or U7851 (N_7851,N_1600,N_2212);
xor U7852 (N_7852,N_4343,N_4501);
nor U7853 (N_7853,N_2234,N_2022);
nand U7854 (N_7854,N_850,N_1941);
nor U7855 (N_7855,N_82,N_3365);
nand U7856 (N_7856,N_2807,N_392);
nor U7857 (N_7857,N_3290,N_3198);
or U7858 (N_7858,N_1160,N_3090);
or U7859 (N_7859,N_3839,N_4844);
or U7860 (N_7860,N_2585,N_1843);
nor U7861 (N_7861,N_2478,N_3143);
xor U7862 (N_7862,N_3111,N_78);
nor U7863 (N_7863,N_1151,N_187);
or U7864 (N_7864,N_4614,N_2668);
and U7865 (N_7865,N_3036,N_2094);
xor U7866 (N_7866,N_665,N_1855);
nor U7867 (N_7867,N_1048,N_2848);
nand U7868 (N_7868,N_4717,N_3389);
or U7869 (N_7869,N_339,N_1654);
nand U7870 (N_7870,N_978,N_1898);
xor U7871 (N_7871,N_1215,N_873);
xor U7872 (N_7872,N_1320,N_135);
and U7873 (N_7873,N_2116,N_3952);
nand U7874 (N_7874,N_2623,N_2488);
or U7875 (N_7875,N_988,N_2705);
or U7876 (N_7876,N_2878,N_3896);
nand U7877 (N_7877,N_560,N_23);
nand U7878 (N_7878,N_370,N_4331);
nand U7879 (N_7879,N_3825,N_2407);
nor U7880 (N_7880,N_1056,N_3034);
or U7881 (N_7881,N_1242,N_4733);
and U7882 (N_7882,N_3378,N_4145);
nand U7883 (N_7883,N_2963,N_522);
or U7884 (N_7884,N_2206,N_1311);
nand U7885 (N_7885,N_3373,N_148);
nor U7886 (N_7886,N_1254,N_3270);
and U7887 (N_7887,N_4198,N_912);
and U7888 (N_7888,N_1488,N_214);
and U7889 (N_7889,N_310,N_268);
nand U7890 (N_7890,N_1453,N_2300);
xnor U7891 (N_7891,N_2734,N_905);
xnor U7892 (N_7892,N_2017,N_1141);
xnor U7893 (N_7893,N_2432,N_1870);
and U7894 (N_7894,N_1997,N_4153);
xor U7895 (N_7895,N_2557,N_3945);
or U7896 (N_7896,N_185,N_795);
xnor U7897 (N_7897,N_1922,N_2095);
xnor U7898 (N_7898,N_2190,N_3995);
or U7899 (N_7899,N_2416,N_3856);
and U7900 (N_7900,N_628,N_1449);
xnor U7901 (N_7901,N_2314,N_1923);
xor U7902 (N_7902,N_1841,N_730);
xor U7903 (N_7903,N_2097,N_388);
xor U7904 (N_7904,N_2854,N_2746);
and U7905 (N_7905,N_4837,N_1501);
or U7906 (N_7906,N_1637,N_1580);
nand U7907 (N_7907,N_165,N_2350);
nand U7908 (N_7908,N_3198,N_2917);
and U7909 (N_7909,N_3769,N_2250);
xor U7910 (N_7910,N_2872,N_4856);
and U7911 (N_7911,N_3645,N_1516);
nor U7912 (N_7912,N_1725,N_983);
nand U7913 (N_7913,N_1462,N_4666);
xnor U7914 (N_7914,N_115,N_2120);
nor U7915 (N_7915,N_3480,N_693);
nor U7916 (N_7916,N_13,N_2766);
or U7917 (N_7917,N_3967,N_4214);
and U7918 (N_7918,N_3851,N_1789);
and U7919 (N_7919,N_500,N_4276);
or U7920 (N_7920,N_770,N_1132);
nor U7921 (N_7921,N_3842,N_3725);
nor U7922 (N_7922,N_442,N_3271);
nand U7923 (N_7923,N_2866,N_245);
nand U7924 (N_7924,N_3778,N_3757);
nor U7925 (N_7925,N_757,N_2710);
nor U7926 (N_7926,N_1048,N_523);
nor U7927 (N_7927,N_883,N_3440);
xor U7928 (N_7928,N_1273,N_2494);
or U7929 (N_7929,N_594,N_4999);
nor U7930 (N_7930,N_4703,N_4868);
nor U7931 (N_7931,N_1174,N_4069);
nor U7932 (N_7932,N_1609,N_4917);
nor U7933 (N_7933,N_4600,N_1754);
nor U7934 (N_7934,N_472,N_3112);
nor U7935 (N_7935,N_3338,N_4881);
xnor U7936 (N_7936,N_4933,N_4795);
xor U7937 (N_7937,N_3905,N_4773);
xnor U7938 (N_7938,N_1526,N_3988);
and U7939 (N_7939,N_3319,N_708);
nor U7940 (N_7940,N_2733,N_3017);
and U7941 (N_7941,N_210,N_806);
and U7942 (N_7942,N_7,N_4006);
or U7943 (N_7943,N_4454,N_3724);
nand U7944 (N_7944,N_454,N_2545);
and U7945 (N_7945,N_1511,N_2863);
nand U7946 (N_7946,N_2704,N_860);
and U7947 (N_7947,N_795,N_336);
or U7948 (N_7948,N_1265,N_711);
nand U7949 (N_7949,N_3560,N_4326);
or U7950 (N_7950,N_4587,N_1326);
xor U7951 (N_7951,N_3492,N_4442);
nor U7952 (N_7952,N_566,N_110);
nand U7953 (N_7953,N_1555,N_4192);
or U7954 (N_7954,N_2542,N_328);
nand U7955 (N_7955,N_1818,N_1655);
or U7956 (N_7956,N_2831,N_599);
xnor U7957 (N_7957,N_4968,N_2301);
and U7958 (N_7958,N_3678,N_2318);
xnor U7959 (N_7959,N_1435,N_4773);
xnor U7960 (N_7960,N_816,N_856);
and U7961 (N_7961,N_888,N_2402);
nand U7962 (N_7962,N_2187,N_4213);
nor U7963 (N_7963,N_1106,N_342);
and U7964 (N_7964,N_387,N_2830);
nor U7965 (N_7965,N_4945,N_2942);
or U7966 (N_7966,N_3896,N_3365);
nor U7967 (N_7967,N_4328,N_3358);
and U7968 (N_7968,N_3666,N_577);
xor U7969 (N_7969,N_268,N_3762);
or U7970 (N_7970,N_4482,N_3807);
xnor U7971 (N_7971,N_1182,N_3260);
xor U7972 (N_7972,N_3531,N_3479);
or U7973 (N_7973,N_1900,N_2561);
xnor U7974 (N_7974,N_666,N_2339);
or U7975 (N_7975,N_3725,N_67);
xnor U7976 (N_7976,N_3733,N_2528);
nand U7977 (N_7977,N_2331,N_3488);
or U7978 (N_7978,N_2078,N_3207);
and U7979 (N_7979,N_4934,N_3286);
or U7980 (N_7980,N_1917,N_2499);
nor U7981 (N_7981,N_457,N_1968);
xnor U7982 (N_7982,N_4555,N_636);
xnor U7983 (N_7983,N_4147,N_4052);
xor U7984 (N_7984,N_3772,N_1954);
xnor U7985 (N_7985,N_4155,N_685);
or U7986 (N_7986,N_742,N_77);
nand U7987 (N_7987,N_3974,N_1116);
xnor U7988 (N_7988,N_331,N_2948);
nor U7989 (N_7989,N_203,N_2297);
xnor U7990 (N_7990,N_2917,N_119);
and U7991 (N_7991,N_2561,N_3025);
xnor U7992 (N_7992,N_4833,N_3170);
xnor U7993 (N_7993,N_1106,N_3145);
or U7994 (N_7994,N_35,N_1142);
nor U7995 (N_7995,N_2709,N_4550);
nand U7996 (N_7996,N_1340,N_150);
and U7997 (N_7997,N_2784,N_3361);
nand U7998 (N_7998,N_2628,N_2140);
nor U7999 (N_7999,N_2192,N_941);
or U8000 (N_8000,N_1488,N_132);
xnor U8001 (N_8001,N_1200,N_3155);
xor U8002 (N_8002,N_4149,N_4142);
xnor U8003 (N_8003,N_4121,N_3231);
xor U8004 (N_8004,N_1303,N_4409);
nand U8005 (N_8005,N_1256,N_4600);
xor U8006 (N_8006,N_3208,N_2167);
nand U8007 (N_8007,N_2225,N_2553);
nor U8008 (N_8008,N_4471,N_4409);
xnor U8009 (N_8009,N_2802,N_277);
nor U8010 (N_8010,N_844,N_2495);
or U8011 (N_8011,N_150,N_484);
and U8012 (N_8012,N_3857,N_3636);
and U8013 (N_8013,N_3664,N_2352);
nor U8014 (N_8014,N_4969,N_2527);
xnor U8015 (N_8015,N_228,N_3462);
or U8016 (N_8016,N_1475,N_4433);
or U8017 (N_8017,N_2491,N_715);
nand U8018 (N_8018,N_1143,N_4867);
or U8019 (N_8019,N_392,N_2373);
or U8020 (N_8020,N_3972,N_3475);
xnor U8021 (N_8021,N_2555,N_4192);
and U8022 (N_8022,N_3553,N_364);
and U8023 (N_8023,N_1692,N_2752);
or U8024 (N_8024,N_4997,N_4148);
nor U8025 (N_8025,N_3682,N_2445);
nor U8026 (N_8026,N_3786,N_2356);
xor U8027 (N_8027,N_1312,N_3652);
or U8028 (N_8028,N_2739,N_1524);
nor U8029 (N_8029,N_3799,N_3366);
nor U8030 (N_8030,N_191,N_3741);
nor U8031 (N_8031,N_4037,N_3256);
nand U8032 (N_8032,N_2822,N_2151);
xnor U8033 (N_8033,N_4515,N_4284);
xnor U8034 (N_8034,N_1793,N_1717);
or U8035 (N_8035,N_1486,N_1472);
nand U8036 (N_8036,N_1854,N_1578);
nor U8037 (N_8037,N_1856,N_733);
nand U8038 (N_8038,N_2600,N_3538);
or U8039 (N_8039,N_4663,N_3620);
nand U8040 (N_8040,N_795,N_1213);
nor U8041 (N_8041,N_1499,N_1190);
or U8042 (N_8042,N_421,N_2975);
nand U8043 (N_8043,N_2770,N_2960);
or U8044 (N_8044,N_1516,N_1671);
and U8045 (N_8045,N_883,N_4441);
xnor U8046 (N_8046,N_4934,N_1587);
nor U8047 (N_8047,N_657,N_900);
nand U8048 (N_8048,N_3035,N_4827);
and U8049 (N_8049,N_3414,N_1791);
nand U8050 (N_8050,N_221,N_3962);
xor U8051 (N_8051,N_793,N_602);
nor U8052 (N_8052,N_1534,N_1454);
or U8053 (N_8053,N_4618,N_488);
xor U8054 (N_8054,N_982,N_2558);
or U8055 (N_8055,N_4928,N_771);
and U8056 (N_8056,N_3864,N_4920);
nand U8057 (N_8057,N_4076,N_840);
xor U8058 (N_8058,N_3239,N_2204);
nand U8059 (N_8059,N_621,N_2661);
nor U8060 (N_8060,N_1570,N_2209);
nand U8061 (N_8061,N_4859,N_854);
nand U8062 (N_8062,N_1291,N_469);
nor U8063 (N_8063,N_4588,N_537);
xor U8064 (N_8064,N_987,N_1950);
and U8065 (N_8065,N_1470,N_1120);
xor U8066 (N_8066,N_2174,N_4314);
and U8067 (N_8067,N_3083,N_1950);
and U8068 (N_8068,N_4473,N_3906);
nand U8069 (N_8069,N_2977,N_1044);
nor U8070 (N_8070,N_3323,N_3329);
nand U8071 (N_8071,N_4987,N_3140);
or U8072 (N_8072,N_648,N_2477);
or U8073 (N_8073,N_2910,N_4110);
and U8074 (N_8074,N_4184,N_2089);
nand U8075 (N_8075,N_646,N_4014);
and U8076 (N_8076,N_4540,N_1999);
or U8077 (N_8077,N_3059,N_4071);
xor U8078 (N_8078,N_1215,N_3288);
nor U8079 (N_8079,N_2115,N_2916);
and U8080 (N_8080,N_4501,N_4044);
and U8081 (N_8081,N_3173,N_3369);
nand U8082 (N_8082,N_331,N_3362);
or U8083 (N_8083,N_2922,N_3991);
xnor U8084 (N_8084,N_4848,N_597);
xnor U8085 (N_8085,N_2697,N_3394);
nor U8086 (N_8086,N_431,N_1227);
nand U8087 (N_8087,N_3,N_2075);
and U8088 (N_8088,N_2786,N_173);
nand U8089 (N_8089,N_4026,N_2643);
and U8090 (N_8090,N_2115,N_3308);
or U8091 (N_8091,N_4856,N_2455);
xor U8092 (N_8092,N_1768,N_2014);
nand U8093 (N_8093,N_4851,N_1446);
xor U8094 (N_8094,N_1597,N_134);
nor U8095 (N_8095,N_4693,N_4258);
nand U8096 (N_8096,N_3445,N_2907);
nand U8097 (N_8097,N_461,N_4577);
or U8098 (N_8098,N_4550,N_4826);
xor U8099 (N_8099,N_145,N_3703);
or U8100 (N_8100,N_1466,N_165);
xor U8101 (N_8101,N_2705,N_2032);
xnor U8102 (N_8102,N_4672,N_905);
nand U8103 (N_8103,N_4804,N_762);
nor U8104 (N_8104,N_3459,N_3415);
and U8105 (N_8105,N_3503,N_1524);
nand U8106 (N_8106,N_2281,N_4114);
nor U8107 (N_8107,N_966,N_4627);
or U8108 (N_8108,N_4680,N_2341);
xor U8109 (N_8109,N_2033,N_800);
and U8110 (N_8110,N_728,N_2693);
xor U8111 (N_8111,N_3336,N_156);
nand U8112 (N_8112,N_1515,N_3952);
xnor U8113 (N_8113,N_4384,N_172);
or U8114 (N_8114,N_4354,N_794);
nand U8115 (N_8115,N_4807,N_3951);
or U8116 (N_8116,N_1609,N_1362);
xnor U8117 (N_8117,N_2518,N_4653);
and U8118 (N_8118,N_1438,N_783);
xor U8119 (N_8119,N_348,N_4818);
nand U8120 (N_8120,N_3862,N_3250);
xor U8121 (N_8121,N_4132,N_1046);
and U8122 (N_8122,N_3190,N_128);
nor U8123 (N_8123,N_1838,N_3213);
or U8124 (N_8124,N_4486,N_818);
xor U8125 (N_8125,N_2502,N_1419);
and U8126 (N_8126,N_3319,N_2387);
nor U8127 (N_8127,N_3139,N_2355);
nor U8128 (N_8128,N_1100,N_2598);
nor U8129 (N_8129,N_1650,N_4664);
and U8130 (N_8130,N_3939,N_84);
or U8131 (N_8131,N_1313,N_4702);
nand U8132 (N_8132,N_2757,N_3630);
nor U8133 (N_8133,N_4130,N_1295);
nor U8134 (N_8134,N_1873,N_2484);
and U8135 (N_8135,N_2212,N_3341);
and U8136 (N_8136,N_1608,N_1511);
nor U8137 (N_8137,N_4293,N_3824);
nand U8138 (N_8138,N_3965,N_173);
nor U8139 (N_8139,N_4534,N_4296);
or U8140 (N_8140,N_2765,N_4995);
or U8141 (N_8141,N_637,N_4723);
or U8142 (N_8142,N_3771,N_2051);
and U8143 (N_8143,N_2057,N_4118);
or U8144 (N_8144,N_2474,N_1391);
xnor U8145 (N_8145,N_2701,N_3584);
xnor U8146 (N_8146,N_4602,N_648);
and U8147 (N_8147,N_1882,N_2323);
and U8148 (N_8148,N_2107,N_577);
or U8149 (N_8149,N_3684,N_4345);
nor U8150 (N_8150,N_1197,N_1921);
nor U8151 (N_8151,N_3431,N_3908);
or U8152 (N_8152,N_495,N_1878);
nand U8153 (N_8153,N_2587,N_4891);
and U8154 (N_8154,N_980,N_2782);
nor U8155 (N_8155,N_4169,N_1139);
nor U8156 (N_8156,N_1413,N_3798);
and U8157 (N_8157,N_2947,N_3918);
xor U8158 (N_8158,N_282,N_4168);
and U8159 (N_8159,N_391,N_1741);
and U8160 (N_8160,N_1010,N_2057);
nand U8161 (N_8161,N_4802,N_4175);
and U8162 (N_8162,N_3413,N_614);
nor U8163 (N_8163,N_3884,N_4023);
xnor U8164 (N_8164,N_1186,N_2320);
nor U8165 (N_8165,N_503,N_398);
or U8166 (N_8166,N_3078,N_3582);
or U8167 (N_8167,N_3391,N_3127);
nor U8168 (N_8168,N_1420,N_1477);
or U8169 (N_8169,N_2424,N_3919);
and U8170 (N_8170,N_1250,N_2059);
nor U8171 (N_8171,N_3449,N_459);
nand U8172 (N_8172,N_2677,N_2535);
or U8173 (N_8173,N_4963,N_439);
xnor U8174 (N_8174,N_3368,N_4244);
or U8175 (N_8175,N_2973,N_4039);
nor U8176 (N_8176,N_1761,N_1778);
nor U8177 (N_8177,N_4104,N_4821);
nor U8178 (N_8178,N_4445,N_1059);
xnor U8179 (N_8179,N_2947,N_988);
and U8180 (N_8180,N_2610,N_4117);
nand U8181 (N_8181,N_2448,N_2339);
nor U8182 (N_8182,N_657,N_3153);
xnor U8183 (N_8183,N_4252,N_3920);
and U8184 (N_8184,N_412,N_1548);
and U8185 (N_8185,N_4650,N_82);
or U8186 (N_8186,N_3863,N_4402);
and U8187 (N_8187,N_2896,N_4621);
and U8188 (N_8188,N_1479,N_2740);
nor U8189 (N_8189,N_3210,N_1618);
or U8190 (N_8190,N_2134,N_3857);
nand U8191 (N_8191,N_1411,N_1175);
nor U8192 (N_8192,N_1304,N_3782);
or U8193 (N_8193,N_2393,N_2362);
nand U8194 (N_8194,N_1367,N_388);
nor U8195 (N_8195,N_3548,N_2384);
nand U8196 (N_8196,N_3311,N_1315);
nand U8197 (N_8197,N_729,N_3567);
or U8198 (N_8198,N_1101,N_1278);
or U8199 (N_8199,N_69,N_1497);
nor U8200 (N_8200,N_622,N_3799);
and U8201 (N_8201,N_642,N_2976);
nand U8202 (N_8202,N_1817,N_1636);
nand U8203 (N_8203,N_3144,N_424);
nand U8204 (N_8204,N_4563,N_2590);
and U8205 (N_8205,N_1801,N_4274);
or U8206 (N_8206,N_1735,N_4658);
nor U8207 (N_8207,N_763,N_4558);
nor U8208 (N_8208,N_1352,N_3110);
or U8209 (N_8209,N_998,N_4115);
nor U8210 (N_8210,N_900,N_3743);
and U8211 (N_8211,N_2750,N_858);
or U8212 (N_8212,N_2719,N_1500);
nor U8213 (N_8213,N_2355,N_1146);
and U8214 (N_8214,N_1320,N_4521);
or U8215 (N_8215,N_1572,N_4922);
and U8216 (N_8216,N_152,N_814);
xor U8217 (N_8217,N_459,N_1480);
nand U8218 (N_8218,N_4520,N_2818);
nand U8219 (N_8219,N_782,N_2708);
or U8220 (N_8220,N_4956,N_2995);
and U8221 (N_8221,N_1915,N_3656);
and U8222 (N_8222,N_2868,N_4971);
nand U8223 (N_8223,N_1556,N_4201);
nor U8224 (N_8224,N_170,N_2544);
and U8225 (N_8225,N_113,N_3885);
nor U8226 (N_8226,N_3932,N_3765);
nor U8227 (N_8227,N_4510,N_2349);
and U8228 (N_8228,N_1947,N_3427);
xnor U8229 (N_8229,N_3524,N_3172);
xor U8230 (N_8230,N_794,N_2994);
and U8231 (N_8231,N_1213,N_1622);
nand U8232 (N_8232,N_3383,N_4074);
xnor U8233 (N_8233,N_1183,N_4305);
nand U8234 (N_8234,N_4488,N_3224);
and U8235 (N_8235,N_3728,N_642);
xnor U8236 (N_8236,N_1678,N_3528);
nand U8237 (N_8237,N_372,N_1663);
nand U8238 (N_8238,N_2539,N_1092);
and U8239 (N_8239,N_4197,N_2355);
xnor U8240 (N_8240,N_2178,N_4982);
nor U8241 (N_8241,N_4426,N_3052);
xor U8242 (N_8242,N_488,N_4315);
or U8243 (N_8243,N_3630,N_1804);
or U8244 (N_8244,N_3940,N_4584);
xor U8245 (N_8245,N_2804,N_4944);
and U8246 (N_8246,N_2474,N_4642);
xor U8247 (N_8247,N_1643,N_1421);
nor U8248 (N_8248,N_201,N_1880);
and U8249 (N_8249,N_221,N_469);
or U8250 (N_8250,N_4145,N_4257);
xnor U8251 (N_8251,N_2039,N_1965);
nand U8252 (N_8252,N_1929,N_2291);
or U8253 (N_8253,N_4449,N_1586);
and U8254 (N_8254,N_3418,N_802);
or U8255 (N_8255,N_796,N_173);
or U8256 (N_8256,N_975,N_4620);
nand U8257 (N_8257,N_4332,N_577);
nand U8258 (N_8258,N_2027,N_20);
xor U8259 (N_8259,N_3396,N_4940);
xor U8260 (N_8260,N_1696,N_1224);
and U8261 (N_8261,N_3477,N_1781);
nand U8262 (N_8262,N_1383,N_4120);
xor U8263 (N_8263,N_4606,N_3934);
xnor U8264 (N_8264,N_4814,N_1906);
nand U8265 (N_8265,N_4204,N_4461);
nor U8266 (N_8266,N_4195,N_1787);
xnor U8267 (N_8267,N_36,N_1169);
nand U8268 (N_8268,N_2410,N_883);
and U8269 (N_8269,N_3839,N_344);
nor U8270 (N_8270,N_544,N_3180);
nor U8271 (N_8271,N_934,N_2485);
xnor U8272 (N_8272,N_42,N_2939);
nand U8273 (N_8273,N_4287,N_3388);
nand U8274 (N_8274,N_4921,N_1860);
or U8275 (N_8275,N_2038,N_2394);
or U8276 (N_8276,N_3823,N_69);
nand U8277 (N_8277,N_4869,N_394);
and U8278 (N_8278,N_683,N_1530);
nand U8279 (N_8279,N_2092,N_2026);
and U8280 (N_8280,N_3698,N_4913);
or U8281 (N_8281,N_1848,N_3837);
xor U8282 (N_8282,N_1993,N_2302);
nand U8283 (N_8283,N_102,N_827);
or U8284 (N_8284,N_1905,N_378);
and U8285 (N_8285,N_1169,N_123);
xnor U8286 (N_8286,N_2944,N_2046);
nor U8287 (N_8287,N_821,N_1123);
nand U8288 (N_8288,N_4545,N_1480);
xor U8289 (N_8289,N_3003,N_2243);
xnor U8290 (N_8290,N_2210,N_2155);
nand U8291 (N_8291,N_198,N_1843);
and U8292 (N_8292,N_4267,N_1214);
xor U8293 (N_8293,N_2856,N_2966);
xor U8294 (N_8294,N_3726,N_2680);
nor U8295 (N_8295,N_2459,N_497);
nand U8296 (N_8296,N_379,N_4861);
and U8297 (N_8297,N_953,N_28);
and U8298 (N_8298,N_2195,N_500);
or U8299 (N_8299,N_1435,N_3569);
nor U8300 (N_8300,N_1721,N_4099);
xor U8301 (N_8301,N_4650,N_1867);
and U8302 (N_8302,N_4532,N_885);
and U8303 (N_8303,N_1588,N_4716);
xor U8304 (N_8304,N_2752,N_1960);
or U8305 (N_8305,N_4264,N_856);
and U8306 (N_8306,N_2095,N_603);
nor U8307 (N_8307,N_3375,N_4424);
nor U8308 (N_8308,N_2633,N_259);
xnor U8309 (N_8309,N_1586,N_4049);
xor U8310 (N_8310,N_1374,N_4886);
nor U8311 (N_8311,N_2509,N_3193);
or U8312 (N_8312,N_4230,N_1201);
xor U8313 (N_8313,N_378,N_3521);
or U8314 (N_8314,N_2119,N_4080);
and U8315 (N_8315,N_1570,N_519);
xor U8316 (N_8316,N_4973,N_520);
or U8317 (N_8317,N_3465,N_1425);
or U8318 (N_8318,N_3050,N_2946);
xor U8319 (N_8319,N_2918,N_3223);
or U8320 (N_8320,N_4614,N_3375);
and U8321 (N_8321,N_657,N_215);
and U8322 (N_8322,N_2774,N_906);
and U8323 (N_8323,N_684,N_2138);
xor U8324 (N_8324,N_4192,N_2191);
nor U8325 (N_8325,N_4201,N_3387);
and U8326 (N_8326,N_2146,N_580);
nand U8327 (N_8327,N_2702,N_1900);
nor U8328 (N_8328,N_4797,N_1846);
nand U8329 (N_8329,N_2460,N_914);
nand U8330 (N_8330,N_2032,N_2741);
nor U8331 (N_8331,N_744,N_3180);
or U8332 (N_8332,N_4084,N_3271);
nor U8333 (N_8333,N_3888,N_2236);
or U8334 (N_8334,N_2575,N_376);
and U8335 (N_8335,N_2172,N_1902);
xor U8336 (N_8336,N_3318,N_3891);
xnor U8337 (N_8337,N_3258,N_1960);
nor U8338 (N_8338,N_1641,N_3983);
nand U8339 (N_8339,N_1657,N_12);
nand U8340 (N_8340,N_3965,N_2285);
nor U8341 (N_8341,N_988,N_3418);
nor U8342 (N_8342,N_2181,N_1110);
nand U8343 (N_8343,N_4218,N_4408);
xnor U8344 (N_8344,N_4556,N_1235);
xnor U8345 (N_8345,N_1814,N_3193);
nand U8346 (N_8346,N_198,N_2147);
nand U8347 (N_8347,N_2957,N_2627);
xnor U8348 (N_8348,N_3881,N_2759);
or U8349 (N_8349,N_510,N_4898);
and U8350 (N_8350,N_2323,N_4063);
and U8351 (N_8351,N_2151,N_40);
or U8352 (N_8352,N_661,N_4572);
nand U8353 (N_8353,N_1297,N_1877);
and U8354 (N_8354,N_4332,N_3590);
or U8355 (N_8355,N_4811,N_3251);
xor U8356 (N_8356,N_1209,N_649);
or U8357 (N_8357,N_3808,N_3203);
or U8358 (N_8358,N_3993,N_2325);
nand U8359 (N_8359,N_3712,N_4402);
nand U8360 (N_8360,N_4764,N_2661);
nor U8361 (N_8361,N_3656,N_2925);
and U8362 (N_8362,N_227,N_581);
nand U8363 (N_8363,N_4255,N_1280);
nand U8364 (N_8364,N_1719,N_4370);
nor U8365 (N_8365,N_1690,N_2820);
and U8366 (N_8366,N_3680,N_4721);
nand U8367 (N_8367,N_62,N_2202);
or U8368 (N_8368,N_4075,N_2887);
xor U8369 (N_8369,N_681,N_98);
xor U8370 (N_8370,N_509,N_3303);
nand U8371 (N_8371,N_1979,N_1753);
xor U8372 (N_8372,N_2575,N_779);
nor U8373 (N_8373,N_2469,N_479);
nand U8374 (N_8374,N_225,N_1995);
or U8375 (N_8375,N_2381,N_3648);
and U8376 (N_8376,N_3759,N_1437);
nand U8377 (N_8377,N_2986,N_2725);
xor U8378 (N_8378,N_1869,N_1585);
nor U8379 (N_8379,N_204,N_1437);
nand U8380 (N_8380,N_3859,N_3856);
nand U8381 (N_8381,N_2953,N_487);
or U8382 (N_8382,N_1480,N_1712);
and U8383 (N_8383,N_705,N_241);
and U8384 (N_8384,N_4250,N_4387);
or U8385 (N_8385,N_1107,N_3750);
nor U8386 (N_8386,N_2859,N_2332);
nand U8387 (N_8387,N_2844,N_1166);
nand U8388 (N_8388,N_2578,N_3923);
xnor U8389 (N_8389,N_768,N_2737);
and U8390 (N_8390,N_2193,N_1750);
nor U8391 (N_8391,N_3935,N_350);
nor U8392 (N_8392,N_668,N_2093);
nand U8393 (N_8393,N_8,N_2117);
or U8394 (N_8394,N_1588,N_1167);
nand U8395 (N_8395,N_718,N_3947);
xor U8396 (N_8396,N_576,N_3200);
nor U8397 (N_8397,N_1507,N_4907);
or U8398 (N_8398,N_1483,N_4655);
nor U8399 (N_8399,N_1898,N_64);
xnor U8400 (N_8400,N_116,N_3216);
or U8401 (N_8401,N_998,N_4465);
and U8402 (N_8402,N_1058,N_3007);
nand U8403 (N_8403,N_2913,N_3363);
nor U8404 (N_8404,N_1970,N_2762);
and U8405 (N_8405,N_50,N_151);
or U8406 (N_8406,N_2827,N_4717);
nor U8407 (N_8407,N_2622,N_3815);
nand U8408 (N_8408,N_1792,N_75);
and U8409 (N_8409,N_3184,N_2732);
or U8410 (N_8410,N_1040,N_3927);
or U8411 (N_8411,N_1331,N_1044);
nor U8412 (N_8412,N_2763,N_3405);
and U8413 (N_8413,N_4098,N_3246);
nand U8414 (N_8414,N_3074,N_2944);
and U8415 (N_8415,N_2044,N_2858);
nor U8416 (N_8416,N_1651,N_4749);
xor U8417 (N_8417,N_3825,N_3591);
and U8418 (N_8418,N_3280,N_2227);
xnor U8419 (N_8419,N_3190,N_3437);
xor U8420 (N_8420,N_2774,N_4596);
or U8421 (N_8421,N_1438,N_4994);
and U8422 (N_8422,N_3021,N_61);
and U8423 (N_8423,N_2313,N_3606);
or U8424 (N_8424,N_837,N_10);
or U8425 (N_8425,N_4310,N_3191);
xor U8426 (N_8426,N_2918,N_2816);
xnor U8427 (N_8427,N_2099,N_3897);
or U8428 (N_8428,N_2543,N_2693);
xnor U8429 (N_8429,N_1677,N_2757);
xnor U8430 (N_8430,N_2352,N_924);
xnor U8431 (N_8431,N_4416,N_4577);
and U8432 (N_8432,N_2005,N_1677);
nand U8433 (N_8433,N_3132,N_1823);
or U8434 (N_8434,N_2512,N_4119);
and U8435 (N_8435,N_1943,N_2227);
nor U8436 (N_8436,N_3512,N_4362);
nand U8437 (N_8437,N_4511,N_339);
nand U8438 (N_8438,N_2953,N_2372);
nor U8439 (N_8439,N_2337,N_2908);
or U8440 (N_8440,N_952,N_3720);
or U8441 (N_8441,N_4518,N_3753);
nor U8442 (N_8442,N_2418,N_2927);
nor U8443 (N_8443,N_3635,N_444);
xnor U8444 (N_8444,N_2,N_1868);
nor U8445 (N_8445,N_1044,N_3304);
or U8446 (N_8446,N_4633,N_2314);
nand U8447 (N_8447,N_979,N_3443);
nor U8448 (N_8448,N_2033,N_964);
nor U8449 (N_8449,N_4644,N_195);
or U8450 (N_8450,N_255,N_1448);
nand U8451 (N_8451,N_2194,N_4778);
and U8452 (N_8452,N_4367,N_4489);
xnor U8453 (N_8453,N_4936,N_4845);
or U8454 (N_8454,N_3134,N_4281);
xnor U8455 (N_8455,N_950,N_1834);
and U8456 (N_8456,N_4003,N_2651);
nand U8457 (N_8457,N_3333,N_2469);
and U8458 (N_8458,N_1516,N_1740);
and U8459 (N_8459,N_4938,N_3987);
and U8460 (N_8460,N_444,N_1344);
nand U8461 (N_8461,N_2247,N_1323);
xnor U8462 (N_8462,N_884,N_2281);
nand U8463 (N_8463,N_427,N_4823);
nand U8464 (N_8464,N_4300,N_2242);
nand U8465 (N_8465,N_238,N_1851);
and U8466 (N_8466,N_3887,N_3298);
nand U8467 (N_8467,N_4745,N_3547);
and U8468 (N_8468,N_2907,N_1266);
xor U8469 (N_8469,N_2014,N_4038);
nor U8470 (N_8470,N_268,N_3068);
nor U8471 (N_8471,N_1817,N_1650);
and U8472 (N_8472,N_2688,N_1318);
and U8473 (N_8473,N_3195,N_695);
nand U8474 (N_8474,N_4516,N_3498);
xor U8475 (N_8475,N_1111,N_1243);
xor U8476 (N_8476,N_4444,N_2842);
or U8477 (N_8477,N_2458,N_2505);
nand U8478 (N_8478,N_2187,N_2552);
nand U8479 (N_8479,N_2064,N_1938);
and U8480 (N_8480,N_1373,N_3357);
xnor U8481 (N_8481,N_3801,N_911);
nor U8482 (N_8482,N_1413,N_484);
xnor U8483 (N_8483,N_1234,N_2633);
nor U8484 (N_8484,N_1298,N_4690);
and U8485 (N_8485,N_2133,N_3971);
nor U8486 (N_8486,N_168,N_1464);
or U8487 (N_8487,N_3792,N_4811);
xnor U8488 (N_8488,N_1424,N_2805);
and U8489 (N_8489,N_3053,N_3011);
and U8490 (N_8490,N_1014,N_2242);
xor U8491 (N_8491,N_1097,N_1771);
or U8492 (N_8492,N_4889,N_2550);
xnor U8493 (N_8493,N_3057,N_2028);
nor U8494 (N_8494,N_255,N_4300);
or U8495 (N_8495,N_351,N_2782);
or U8496 (N_8496,N_4439,N_3404);
xor U8497 (N_8497,N_2666,N_1853);
xor U8498 (N_8498,N_3628,N_4133);
and U8499 (N_8499,N_4550,N_1595);
nand U8500 (N_8500,N_1187,N_3611);
or U8501 (N_8501,N_3304,N_4471);
xnor U8502 (N_8502,N_647,N_3089);
or U8503 (N_8503,N_1538,N_4715);
or U8504 (N_8504,N_284,N_3697);
xor U8505 (N_8505,N_2540,N_2815);
xnor U8506 (N_8506,N_770,N_4200);
nand U8507 (N_8507,N_3070,N_2763);
or U8508 (N_8508,N_783,N_1206);
or U8509 (N_8509,N_621,N_2263);
xor U8510 (N_8510,N_1518,N_4308);
or U8511 (N_8511,N_3281,N_2338);
xnor U8512 (N_8512,N_1372,N_4218);
nor U8513 (N_8513,N_4600,N_2549);
and U8514 (N_8514,N_3270,N_4729);
nor U8515 (N_8515,N_2679,N_7);
and U8516 (N_8516,N_242,N_4317);
nor U8517 (N_8517,N_974,N_1526);
or U8518 (N_8518,N_4206,N_1741);
and U8519 (N_8519,N_3387,N_2710);
nor U8520 (N_8520,N_110,N_2193);
or U8521 (N_8521,N_2913,N_2998);
or U8522 (N_8522,N_4948,N_957);
nor U8523 (N_8523,N_1248,N_1116);
nand U8524 (N_8524,N_618,N_3304);
nand U8525 (N_8525,N_3627,N_263);
or U8526 (N_8526,N_1283,N_4500);
and U8527 (N_8527,N_1370,N_893);
or U8528 (N_8528,N_3941,N_4284);
nand U8529 (N_8529,N_3496,N_4995);
nand U8530 (N_8530,N_1505,N_4953);
and U8531 (N_8531,N_4476,N_2297);
nor U8532 (N_8532,N_1942,N_2341);
xnor U8533 (N_8533,N_970,N_1090);
and U8534 (N_8534,N_1584,N_94);
xor U8535 (N_8535,N_3221,N_497);
nand U8536 (N_8536,N_932,N_3989);
nor U8537 (N_8537,N_2417,N_2243);
nand U8538 (N_8538,N_2803,N_185);
or U8539 (N_8539,N_2206,N_2548);
and U8540 (N_8540,N_475,N_1366);
nand U8541 (N_8541,N_214,N_1825);
nand U8542 (N_8542,N_3517,N_566);
nand U8543 (N_8543,N_2967,N_1786);
nand U8544 (N_8544,N_2760,N_3997);
and U8545 (N_8545,N_3371,N_3135);
xor U8546 (N_8546,N_2041,N_974);
or U8547 (N_8547,N_1119,N_4380);
nor U8548 (N_8548,N_2217,N_1796);
or U8549 (N_8549,N_811,N_4128);
xnor U8550 (N_8550,N_4623,N_3277);
nand U8551 (N_8551,N_72,N_4286);
and U8552 (N_8552,N_4034,N_4158);
nor U8553 (N_8553,N_3160,N_1441);
nand U8554 (N_8554,N_2339,N_1576);
xnor U8555 (N_8555,N_331,N_4464);
xor U8556 (N_8556,N_4663,N_1178);
or U8557 (N_8557,N_4083,N_2806);
xnor U8558 (N_8558,N_4568,N_3900);
and U8559 (N_8559,N_4511,N_2114);
or U8560 (N_8560,N_4013,N_3753);
nand U8561 (N_8561,N_556,N_2221);
nor U8562 (N_8562,N_3138,N_877);
and U8563 (N_8563,N_2926,N_2628);
xnor U8564 (N_8564,N_293,N_3087);
nand U8565 (N_8565,N_3420,N_191);
nor U8566 (N_8566,N_1891,N_2709);
or U8567 (N_8567,N_479,N_237);
and U8568 (N_8568,N_844,N_2025);
xor U8569 (N_8569,N_636,N_227);
or U8570 (N_8570,N_1630,N_2438);
nand U8571 (N_8571,N_3606,N_4805);
xor U8572 (N_8572,N_4886,N_3582);
and U8573 (N_8573,N_505,N_276);
or U8574 (N_8574,N_4942,N_2596);
or U8575 (N_8575,N_4704,N_3027);
and U8576 (N_8576,N_4626,N_3045);
nand U8577 (N_8577,N_3396,N_3842);
nand U8578 (N_8578,N_3537,N_4009);
nand U8579 (N_8579,N_3160,N_4608);
nor U8580 (N_8580,N_3167,N_150);
or U8581 (N_8581,N_2709,N_3116);
nor U8582 (N_8582,N_2364,N_4596);
nand U8583 (N_8583,N_4401,N_2825);
and U8584 (N_8584,N_3050,N_4773);
nor U8585 (N_8585,N_2417,N_3705);
nand U8586 (N_8586,N_4070,N_2689);
or U8587 (N_8587,N_244,N_3904);
or U8588 (N_8588,N_1453,N_1999);
and U8589 (N_8589,N_1305,N_2974);
or U8590 (N_8590,N_1204,N_3707);
nor U8591 (N_8591,N_2001,N_3191);
nand U8592 (N_8592,N_612,N_1007);
or U8593 (N_8593,N_61,N_18);
nor U8594 (N_8594,N_3794,N_1640);
nand U8595 (N_8595,N_2535,N_3330);
nand U8596 (N_8596,N_3575,N_4409);
or U8597 (N_8597,N_4010,N_4882);
nor U8598 (N_8598,N_4356,N_4576);
and U8599 (N_8599,N_2603,N_4596);
nand U8600 (N_8600,N_4966,N_4041);
nand U8601 (N_8601,N_4812,N_1121);
xnor U8602 (N_8602,N_877,N_3976);
nor U8603 (N_8603,N_792,N_1308);
and U8604 (N_8604,N_1441,N_4621);
or U8605 (N_8605,N_3377,N_2759);
or U8606 (N_8606,N_2238,N_3962);
and U8607 (N_8607,N_2563,N_2514);
and U8608 (N_8608,N_1705,N_1405);
or U8609 (N_8609,N_1021,N_1062);
nor U8610 (N_8610,N_1262,N_3790);
xnor U8611 (N_8611,N_1983,N_291);
xor U8612 (N_8612,N_875,N_2470);
or U8613 (N_8613,N_3637,N_2170);
nor U8614 (N_8614,N_2675,N_895);
or U8615 (N_8615,N_1118,N_1355);
and U8616 (N_8616,N_2142,N_337);
xor U8617 (N_8617,N_774,N_471);
or U8618 (N_8618,N_4026,N_1473);
and U8619 (N_8619,N_1222,N_2282);
xor U8620 (N_8620,N_4972,N_2496);
nand U8621 (N_8621,N_515,N_4941);
and U8622 (N_8622,N_689,N_2450);
or U8623 (N_8623,N_3905,N_1275);
nor U8624 (N_8624,N_2607,N_4247);
nor U8625 (N_8625,N_1371,N_1384);
nor U8626 (N_8626,N_4939,N_3132);
nand U8627 (N_8627,N_4368,N_733);
and U8628 (N_8628,N_2419,N_1580);
nor U8629 (N_8629,N_2908,N_1574);
nand U8630 (N_8630,N_4285,N_2441);
nand U8631 (N_8631,N_1752,N_4887);
or U8632 (N_8632,N_3936,N_4869);
xnor U8633 (N_8633,N_4039,N_3604);
xor U8634 (N_8634,N_5,N_2312);
nand U8635 (N_8635,N_265,N_849);
nand U8636 (N_8636,N_2565,N_3240);
xor U8637 (N_8637,N_1029,N_3379);
or U8638 (N_8638,N_1990,N_3153);
nand U8639 (N_8639,N_4853,N_4173);
nor U8640 (N_8640,N_737,N_4113);
and U8641 (N_8641,N_918,N_4673);
and U8642 (N_8642,N_3911,N_4078);
xor U8643 (N_8643,N_3319,N_1367);
and U8644 (N_8644,N_2998,N_760);
and U8645 (N_8645,N_4533,N_1247);
nor U8646 (N_8646,N_1719,N_4323);
or U8647 (N_8647,N_458,N_2245);
nand U8648 (N_8648,N_977,N_1955);
or U8649 (N_8649,N_2265,N_1609);
nor U8650 (N_8650,N_161,N_4293);
nand U8651 (N_8651,N_3676,N_3285);
nand U8652 (N_8652,N_4736,N_2411);
and U8653 (N_8653,N_2184,N_1525);
or U8654 (N_8654,N_1811,N_195);
or U8655 (N_8655,N_4546,N_3604);
or U8656 (N_8656,N_2458,N_733);
or U8657 (N_8657,N_3906,N_1253);
nand U8658 (N_8658,N_4988,N_4428);
nand U8659 (N_8659,N_2593,N_3822);
nand U8660 (N_8660,N_4410,N_2440);
or U8661 (N_8661,N_4044,N_3500);
nand U8662 (N_8662,N_1832,N_4831);
xor U8663 (N_8663,N_27,N_289);
or U8664 (N_8664,N_4894,N_2589);
xnor U8665 (N_8665,N_1300,N_2289);
xnor U8666 (N_8666,N_1814,N_2094);
or U8667 (N_8667,N_1631,N_4407);
and U8668 (N_8668,N_936,N_1811);
or U8669 (N_8669,N_4342,N_3626);
or U8670 (N_8670,N_4169,N_539);
or U8671 (N_8671,N_4195,N_3741);
or U8672 (N_8672,N_4324,N_510);
or U8673 (N_8673,N_1835,N_2449);
or U8674 (N_8674,N_459,N_2816);
and U8675 (N_8675,N_4125,N_4717);
nor U8676 (N_8676,N_1997,N_1241);
nor U8677 (N_8677,N_4626,N_3944);
nor U8678 (N_8678,N_4245,N_506);
nand U8679 (N_8679,N_3314,N_4457);
nor U8680 (N_8680,N_4136,N_100);
nor U8681 (N_8681,N_3072,N_3763);
xor U8682 (N_8682,N_66,N_560);
xor U8683 (N_8683,N_2924,N_4995);
nor U8684 (N_8684,N_2648,N_769);
or U8685 (N_8685,N_4628,N_4414);
and U8686 (N_8686,N_1550,N_2980);
xnor U8687 (N_8687,N_1720,N_3735);
nand U8688 (N_8688,N_3570,N_3692);
and U8689 (N_8689,N_1760,N_1624);
and U8690 (N_8690,N_2082,N_4903);
and U8691 (N_8691,N_2018,N_2407);
or U8692 (N_8692,N_296,N_2976);
xor U8693 (N_8693,N_4675,N_118);
nor U8694 (N_8694,N_2878,N_1635);
or U8695 (N_8695,N_202,N_966);
and U8696 (N_8696,N_55,N_2824);
and U8697 (N_8697,N_3395,N_3840);
and U8698 (N_8698,N_380,N_2301);
and U8699 (N_8699,N_2875,N_904);
and U8700 (N_8700,N_4938,N_3247);
nor U8701 (N_8701,N_1702,N_2598);
or U8702 (N_8702,N_4089,N_2271);
and U8703 (N_8703,N_2,N_1410);
nand U8704 (N_8704,N_1307,N_3403);
nand U8705 (N_8705,N_572,N_2815);
nand U8706 (N_8706,N_3339,N_4479);
or U8707 (N_8707,N_2006,N_2547);
nand U8708 (N_8708,N_3308,N_2335);
nor U8709 (N_8709,N_1952,N_3941);
nor U8710 (N_8710,N_2974,N_4772);
xnor U8711 (N_8711,N_3408,N_1947);
xnor U8712 (N_8712,N_1230,N_2545);
and U8713 (N_8713,N_3473,N_2474);
and U8714 (N_8714,N_2088,N_2058);
xnor U8715 (N_8715,N_3215,N_819);
or U8716 (N_8716,N_1462,N_3383);
or U8717 (N_8717,N_2194,N_2659);
nor U8718 (N_8718,N_1097,N_4076);
and U8719 (N_8719,N_3566,N_3253);
or U8720 (N_8720,N_121,N_3692);
nor U8721 (N_8721,N_2253,N_454);
xnor U8722 (N_8722,N_2151,N_725);
or U8723 (N_8723,N_1991,N_4979);
or U8724 (N_8724,N_2167,N_3120);
and U8725 (N_8725,N_385,N_1761);
nor U8726 (N_8726,N_2199,N_1548);
nor U8727 (N_8727,N_2185,N_1653);
or U8728 (N_8728,N_2180,N_4961);
or U8729 (N_8729,N_4128,N_3226);
nor U8730 (N_8730,N_3231,N_2171);
or U8731 (N_8731,N_3791,N_2368);
or U8732 (N_8732,N_4928,N_4850);
xnor U8733 (N_8733,N_4262,N_4972);
and U8734 (N_8734,N_4501,N_1208);
nor U8735 (N_8735,N_620,N_4026);
and U8736 (N_8736,N_3484,N_90);
nor U8737 (N_8737,N_3389,N_4614);
nor U8738 (N_8738,N_3398,N_771);
and U8739 (N_8739,N_4121,N_2950);
nor U8740 (N_8740,N_2252,N_3577);
nand U8741 (N_8741,N_3164,N_1642);
or U8742 (N_8742,N_3911,N_2868);
and U8743 (N_8743,N_1249,N_2276);
and U8744 (N_8744,N_1537,N_629);
and U8745 (N_8745,N_536,N_4856);
and U8746 (N_8746,N_2988,N_3809);
xnor U8747 (N_8747,N_3349,N_2746);
nor U8748 (N_8748,N_4310,N_3151);
and U8749 (N_8749,N_1210,N_2841);
nand U8750 (N_8750,N_2984,N_4330);
xor U8751 (N_8751,N_2173,N_393);
xor U8752 (N_8752,N_1774,N_4909);
nand U8753 (N_8753,N_3434,N_1123);
nand U8754 (N_8754,N_4329,N_4276);
xnor U8755 (N_8755,N_1341,N_114);
nor U8756 (N_8756,N_2900,N_3023);
xor U8757 (N_8757,N_471,N_4943);
and U8758 (N_8758,N_342,N_3278);
and U8759 (N_8759,N_80,N_859);
nand U8760 (N_8760,N_631,N_1095);
nor U8761 (N_8761,N_3413,N_4313);
nand U8762 (N_8762,N_2116,N_3741);
and U8763 (N_8763,N_2146,N_2361);
and U8764 (N_8764,N_1338,N_4327);
nor U8765 (N_8765,N_4956,N_3637);
and U8766 (N_8766,N_1227,N_2203);
nor U8767 (N_8767,N_2091,N_325);
nand U8768 (N_8768,N_4963,N_3443);
xor U8769 (N_8769,N_860,N_1326);
xor U8770 (N_8770,N_917,N_3617);
nand U8771 (N_8771,N_2890,N_1797);
and U8772 (N_8772,N_2057,N_3468);
nand U8773 (N_8773,N_4767,N_3535);
nand U8774 (N_8774,N_3848,N_1392);
nor U8775 (N_8775,N_14,N_2542);
or U8776 (N_8776,N_678,N_4933);
and U8777 (N_8777,N_4655,N_4463);
xor U8778 (N_8778,N_221,N_1806);
nor U8779 (N_8779,N_3030,N_3387);
nand U8780 (N_8780,N_1328,N_4032);
xor U8781 (N_8781,N_3766,N_2903);
xnor U8782 (N_8782,N_2320,N_2821);
or U8783 (N_8783,N_1926,N_486);
or U8784 (N_8784,N_1650,N_3046);
nand U8785 (N_8785,N_4222,N_28);
nand U8786 (N_8786,N_1624,N_2044);
nor U8787 (N_8787,N_3757,N_107);
nand U8788 (N_8788,N_1585,N_935);
nand U8789 (N_8789,N_232,N_4129);
nand U8790 (N_8790,N_3713,N_1395);
and U8791 (N_8791,N_3617,N_380);
and U8792 (N_8792,N_3784,N_1751);
and U8793 (N_8793,N_4233,N_2226);
nor U8794 (N_8794,N_1002,N_3034);
nand U8795 (N_8795,N_4592,N_3288);
and U8796 (N_8796,N_3529,N_242);
xnor U8797 (N_8797,N_3910,N_4821);
nor U8798 (N_8798,N_1448,N_698);
and U8799 (N_8799,N_2320,N_2947);
nor U8800 (N_8800,N_2550,N_3890);
nor U8801 (N_8801,N_2276,N_2291);
or U8802 (N_8802,N_2913,N_4578);
nor U8803 (N_8803,N_4895,N_992);
or U8804 (N_8804,N_3768,N_3723);
nor U8805 (N_8805,N_4531,N_4411);
nor U8806 (N_8806,N_1363,N_1144);
nor U8807 (N_8807,N_3276,N_3400);
nor U8808 (N_8808,N_1105,N_2375);
or U8809 (N_8809,N_1621,N_4018);
and U8810 (N_8810,N_1096,N_1933);
xnor U8811 (N_8811,N_2195,N_2052);
nor U8812 (N_8812,N_1878,N_1320);
or U8813 (N_8813,N_1605,N_3890);
nor U8814 (N_8814,N_1288,N_1587);
xnor U8815 (N_8815,N_3409,N_1220);
and U8816 (N_8816,N_3090,N_3679);
and U8817 (N_8817,N_1257,N_3832);
nor U8818 (N_8818,N_2147,N_508);
xor U8819 (N_8819,N_228,N_1646);
nand U8820 (N_8820,N_527,N_1438);
nor U8821 (N_8821,N_239,N_3247);
nand U8822 (N_8822,N_1734,N_3480);
nor U8823 (N_8823,N_2880,N_2220);
nor U8824 (N_8824,N_801,N_2396);
or U8825 (N_8825,N_1517,N_646);
nand U8826 (N_8826,N_3479,N_4449);
nand U8827 (N_8827,N_1895,N_3725);
nand U8828 (N_8828,N_3833,N_1181);
or U8829 (N_8829,N_2389,N_334);
nor U8830 (N_8830,N_697,N_331);
nand U8831 (N_8831,N_384,N_4418);
or U8832 (N_8832,N_2951,N_4012);
nand U8833 (N_8833,N_984,N_3643);
xnor U8834 (N_8834,N_3495,N_3766);
or U8835 (N_8835,N_1049,N_3907);
nand U8836 (N_8836,N_686,N_1877);
nor U8837 (N_8837,N_236,N_298);
xnor U8838 (N_8838,N_1201,N_2097);
or U8839 (N_8839,N_390,N_669);
and U8840 (N_8840,N_3736,N_1984);
xnor U8841 (N_8841,N_1326,N_3021);
nand U8842 (N_8842,N_3794,N_1028);
and U8843 (N_8843,N_2370,N_1822);
and U8844 (N_8844,N_2084,N_2898);
nor U8845 (N_8845,N_4687,N_3917);
or U8846 (N_8846,N_2052,N_1239);
or U8847 (N_8847,N_2482,N_3383);
nand U8848 (N_8848,N_408,N_1204);
nand U8849 (N_8849,N_1879,N_4843);
or U8850 (N_8850,N_2901,N_3317);
nand U8851 (N_8851,N_1132,N_1760);
and U8852 (N_8852,N_4312,N_2834);
or U8853 (N_8853,N_2144,N_3877);
nor U8854 (N_8854,N_1209,N_2705);
xnor U8855 (N_8855,N_3017,N_1070);
nand U8856 (N_8856,N_1543,N_122);
xor U8857 (N_8857,N_2762,N_3212);
xnor U8858 (N_8858,N_3695,N_3036);
and U8859 (N_8859,N_4811,N_687);
and U8860 (N_8860,N_3961,N_4274);
nand U8861 (N_8861,N_4395,N_428);
nor U8862 (N_8862,N_87,N_1634);
nor U8863 (N_8863,N_3665,N_485);
and U8864 (N_8864,N_3675,N_1337);
nand U8865 (N_8865,N_3730,N_3904);
xnor U8866 (N_8866,N_1107,N_2307);
nand U8867 (N_8867,N_1143,N_3305);
or U8868 (N_8868,N_2725,N_1101);
nor U8869 (N_8869,N_3416,N_1220);
or U8870 (N_8870,N_3241,N_3875);
or U8871 (N_8871,N_547,N_283);
xor U8872 (N_8872,N_156,N_3133);
nor U8873 (N_8873,N_4910,N_2990);
and U8874 (N_8874,N_3004,N_3806);
and U8875 (N_8875,N_4753,N_1582);
xor U8876 (N_8876,N_4006,N_4917);
xor U8877 (N_8877,N_2330,N_4820);
xnor U8878 (N_8878,N_2085,N_3909);
or U8879 (N_8879,N_3437,N_3781);
and U8880 (N_8880,N_3946,N_4447);
nand U8881 (N_8881,N_4379,N_4825);
or U8882 (N_8882,N_1380,N_3719);
nor U8883 (N_8883,N_4991,N_605);
xnor U8884 (N_8884,N_4494,N_4929);
or U8885 (N_8885,N_4139,N_4579);
nand U8886 (N_8886,N_2990,N_2295);
nand U8887 (N_8887,N_2562,N_2676);
and U8888 (N_8888,N_165,N_4190);
and U8889 (N_8889,N_2120,N_1634);
and U8890 (N_8890,N_3099,N_467);
nand U8891 (N_8891,N_1912,N_2367);
xnor U8892 (N_8892,N_4215,N_1985);
nor U8893 (N_8893,N_3078,N_2134);
or U8894 (N_8894,N_1340,N_721);
xor U8895 (N_8895,N_2609,N_3346);
or U8896 (N_8896,N_4817,N_3104);
nor U8897 (N_8897,N_1157,N_1069);
nand U8898 (N_8898,N_1437,N_1153);
or U8899 (N_8899,N_4712,N_4655);
and U8900 (N_8900,N_380,N_3200);
nand U8901 (N_8901,N_4208,N_36);
xnor U8902 (N_8902,N_4183,N_4743);
nand U8903 (N_8903,N_3154,N_499);
and U8904 (N_8904,N_443,N_425);
nor U8905 (N_8905,N_4193,N_3407);
and U8906 (N_8906,N_4186,N_3037);
xor U8907 (N_8907,N_4474,N_2906);
and U8908 (N_8908,N_1114,N_486);
and U8909 (N_8909,N_455,N_3708);
and U8910 (N_8910,N_2295,N_1046);
or U8911 (N_8911,N_1129,N_2464);
and U8912 (N_8912,N_165,N_1247);
and U8913 (N_8913,N_2804,N_3426);
xor U8914 (N_8914,N_2578,N_4018);
nor U8915 (N_8915,N_4413,N_3670);
and U8916 (N_8916,N_3689,N_2898);
xor U8917 (N_8917,N_4960,N_4151);
nor U8918 (N_8918,N_472,N_3554);
or U8919 (N_8919,N_1795,N_4941);
or U8920 (N_8920,N_3807,N_4212);
and U8921 (N_8921,N_3724,N_4440);
nand U8922 (N_8922,N_1680,N_3134);
nand U8923 (N_8923,N_2012,N_4545);
nand U8924 (N_8924,N_3442,N_1717);
and U8925 (N_8925,N_3170,N_628);
nand U8926 (N_8926,N_4434,N_3083);
or U8927 (N_8927,N_2055,N_71);
xnor U8928 (N_8928,N_3869,N_2435);
and U8929 (N_8929,N_4109,N_3220);
nand U8930 (N_8930,N_811,N_3312);
xnor U8931 (N_8931,N_280,N_289);
nand U8932 (N_8932,N_2775,N_3118);
or U8933 (N_8933,N_1864,N_2178);
and U8934 (N_8934,N_4435,N_161);
and U8935 (N_8935,N_820,N_414);
nand U8936 (N_8936,N_4336,N_1895);
nor U8937 (N_8937,N_1542,N_1376);
and U8938 (N_8938,N_621,N_2650);
nor U8939 (N_8939,N_1385,N_1355);
or U8940 (N_8940,N_3909,N_915);
xnor U8941 (N_8941,N_1038,N_1894);
or U8942 (N_8942,N_1881,N_3614);
nand U8943 (N_8943,N_852,N_1672);
nand U8944 (N_8944,N_3024,N_4829);
or U8945 (N_8945,N_4702,N_2666);
nor U8946 (N_8946,N_1645,N_1655);
and U8947 (N_8947,N_4334,N_386);
or U8948 (N_8948,N_810,N_2601);
xor U8949 (N_8949,N_4895,N_928);
or U8950 (N_8950,N_682,N_3192);
or U8951 (N_8951,N_1119,N_607);
nand U8952 (N_8952,N_309,N_1804);
xnor U8953 (N_8953,N_4698,N_2901);
nor U8954 (N_8954,N_4766,N_2755);
and U8955 (N_8955,N_3660,N_4263);
xnor U8956 (N_8956,N_3328,N_2477);
xor U8957 (N_8957,N_1470,N_546);
or U8958 (N_8958,N_3180,N_828);
nor U8959 (N_8959,N_1365,N_4774);
or U8960 (N_8960,N_2479,N_2987);
or U8961 (N_8961,N_3501,N_4292);
xnor U8962 (N_8962,N_4113,N_3661);
xor U8963 (N_8963,N_4240,N_3349);
or U8964 (N_8964,N_3545,N_1026);
nor U8965 (N_8965,N_3607,N_2534);
and U8966 (N_8966,N_2234,N_1719);
and U8967 (N_8967,N_935,N_3349);
xor U8968 (N_8968,N_4511,N_3588);
nand U8969 (N_8969,N_1990,N_2835);
and U8970 (N_8970,N_761,N_1189);
and U8971 (N_8971,N_1811,N_1284);
xor U8972 (N_8972,N_3868,N_4959);
nand U8973 (N_8973,N_1149,N_1883);
xor U8974 (N_8974,N_3427,N_616);
xor U8975 (N_8975,N_1670,N_433);
nand U8976 (N_8976,N_3289,N_4241);
nor U8977 (N_8977,N_3232,N_1038);
nand U8978 (N_8978,N_1092,N_4889);
nor U8979 (N_8979,N_505,N_2855);
nand U8980 (N_8980,N_864,N_4090);
xor U8981 (N_8981,N_1760,N_2713);
xor U8982 (N_8982,N_4359,N_2528);
nor U8983 (N_8983,N_2372,N_4595);
nand U8984 (N_8984,N_476,N_1078);
or U8985 (N_8985,N_3984,N_4758);
nor U8986 (N_8986,N_4924,N_2157);
xor U8987 (N_8987,N_4967,N_2650);
nor U8988 (N_8988,N_127,N_2129);
or U8989 (N_8989,N_1358,N_4714);
nand U8990 (N_8990,N_585,N_2490);
nor U8991 (N_8991,N_4147,N_2960);
xor U8992 (N_8992,N_818,N_506);
nor U8993 (N_8993,N_2386,N_57);
or U8994 (N_8994,N_2551,N_4976);
or U8995 (N_8995,N_3469,N_1554);
or U8996 (N_8996,N_3552,N_11);
xnor U8997 (N_8997,N_3037,N_1094);
and U8998 (N_8998,N_1464,N_105);
nand U8999 (N_8999,N_2420,N_3319);
nor U9000 (N_9000,N_4313,N_1507);
xor U9001 (N_9001,N_1298,N_4172);
xor U9002 (N_9002,N_636,N_2390);
nor U9003 (N_9003,N_1330,N_3445);
nand U9004 (N_9004,N_3300,N_2231);
nand U9005 (N_9005,N_1934,N_4459);
or U9006 (N_9006,N_1109,N_4044);
xnor U9007 (N_9007,N_1947,N_1883);
xor U9008 (N_9008,N_3294,N_870);
and U9009 (N_9009,N_2567,N_4422);
nor U9010 (N_9010,N_4983,N_4521);
xor U9011 (N_9011,N_3135,N_3737);
xor U9012 (N_9012,N_1492,N_221);
nand U9013 (N_9013,N_3139,N_3483);
or U9014 (N_9014,N_1509,N_2077);
or U9015 (N_9015,N_4028,N_4588);
xor U9016 (N_9016,N_283,N_3021);
nand U9017 (N_9017,N_430,N_3518);
or U9018 (N_9018,N_4913,N_4773);
nor U9019 (N_9019,N_903,N_4969);
xnor U9020 (N_9020,N_4354,N_2986);
nand U9021 (N_9021,N_3348,N_2709);
and U9022 (N_9022,N_4860,N_3865);
nor U9023 (N_9023,N_385,N_4195);
nor U9024 (N_9024,N_2588,N_3521);
nor U9025 (N_9025,N_1879,N_4578);
xnor U9026 (N_9026,N_3889,N_1613);
or U9027 (N_9027,N_1296,N_4580);
nor U9028 (N_9028,N_769,N_1098);
or U9029 (N_9029,N_232,N_4145);
nand U9030 (N_9030,N_3703,N_3347);
or U9031 (N_9031,N_2173,N_2787);
nor U9032 (N_9032,N_3527,N_1513);
or U9033 (N_9033,N_3695,N_3547);
nand U9034 (N_9034,N_1640,N_4016);
and U9035 (N_9035,N_247,N_2266);
xnor U9036 (N_9036,N_1196,N_793);
nand U9037 (N_9037,N_4553,N_466);
nor U9038 (N_9038,N_4967,N_4986);
xor U9039 (N_9039,N_232,N_2541);
and U9040 (N_9040,N_1762,N_3286);
and U9041 (N_9041,N_166,N_2499);
xnor U9042 (N_9042,N_4514,N_3593);
or U9043 (N_9043,N_4012,N_3703);
or U9044 (N_9044,N_2119,N_864);
nand U9045 (N_9045,N_1114,N_1462);
nor U9046 (N_9046,N_4711,N_1960);
and U9047 (N_9047,N_4107,N_4644);
or U9048 (N_9048,N_3002,N_3444);
nor U9049 (N_9049,N_612,N_4866);
nand U9050 (N_9050,N_2232,N_1438);
nor U9051 (N_9051,N_3780,N_1941);
xnor U9052 (N_9052,N_1037,N_3524);
nand U9053 (N_9053,N_1549,N_103);
nor U9054 (N_9054,N_4031,N_418);
nor U9055 (N_9055,N_2051,N_2474);
and U9056 (N_9056,N_4479,N_1930);
nand U9057 (N_9057,N_1977,N_1702);
or U9058 (N_9058,N_4936,N_2094);
xor U9059 (N_9059,N_209,N_1301);
or U9060 (N_9060,N_929,N_2417);
nand U9061 (N_9061,N_1146,N_1873);
nand U9062 (N_9062,N_3808,N_4666);
or U9063 (N_9063,N_3071,N_2567);
nand U9064 (N_9064,N_4199,N_348);
nor U9065 (N_9065,N_1885,N_1410);
nor U9066 (N_9066,N_3042,N_4470);
or U9067 (N_9067,N_4606,N_1298);
or U9068 (N_9068,N_4355,N_4430);
and U9069 (N_9069,N_4698,N_1569);
and U9070 (N_9070,N_692,N_3028);
or U9071 (N_9071,N_3231,N_4182);
nand U9072 (N_9072,N_4543,N_2673);
or U9073 (N_9073,N_2222,N_1027);
nor U9074 (N_9074,N_453,N_1869);
or U9075 (N_9075,N_1266,N_4827);
nor U9076 (N_9076,N_1785,N_3958);
xor U9077 (N_9077,N_2955,N_2127);
nand U9078 (N_9078,N_994,N_628);
xor U9079 (N_9079,N_869,N_2449);
nor U9080 (N_9080,N_4336,N_2479);
or U9081 (N_9081,N_435,N_4245);
and U9082 (N_9082,N_4289,N_4602);
or U9083 (N_9083,N_1441,N_1556);
and U9084 (N_9084,N_3535,N_2482);
or U9085 (N_9085,N_4592,N_2951);
or U9086 (N_9086,N_1174,N_1577);
nand U9087 (N_9087,N_1173,N_3979);
nand U9088 (N_9088,N_2362,N_2565);
nand U9089 (N_9089,N_672,N_342);
nor U9090 (N_9090,N_1025,N_3873);
nand U9091 (N_9091,N_1436,N_98);
nand U9092 (N_9092,N_4520,N_4616);
nand U9093 (N_9093,N_3279,N_1385);
xor U9094 (N_9094,N_2759,N_2924);
xor U9095 (N_9095,N_2971,N_4674);
xor U9096 (N_9096,N_2707,N_3826);
nor U9097 (N_9097,N_1810,N_3160);
nand U9098 (N_9098,N_3850,N_4893);
and U9099 (N_9099,N_4784,N_3834);
and U9100 (N_9100,N_1159,N_3437);
xnor U9101 (N_9101,N_4045,N_80);
xor U9102 (N_9102,N_1838,N_4235);
nand U9103 (N_9103,N_4094,N_2181);
and U9104 (N_9104,N_2008,N_3362);
and U9105 (N_9105,N_3630,N_2635);
xor U9106 (N_9106,N_4591,N_2506);
nand U9107 (N_9107,N_2912,N_1758);
nand U9108 (N_9108,N_2420,N_2780);
nand U9109 (N_9109,N_3313,N_3498);
and U9110 (N_9110,N_2082,N_3416);
nand U9111 (N_9111,N_4379,N_3631);
xor U9112 (N_9112,N_1127,N_351);
or U9113 (N_9113,N_1904,N_4639);
or U9114 (N_9114,N_1798,N_4610);
xor U9115 (N_9115,N_2442,N_1211);
or U9116 (N_9116,N_2013,N_839);
xor U9117 (N_9117,N_4129,N_2565);
nand U9118 (N_9118,N_4476,N_1883);
nor U9119 (N_9119,N_4557,N_2605);
nor U9120 (N_9120,N_2673,N_378);
xor U9121 (N_9121,N_4198,N_2940);
nand U9122 (N_9122,N_3467,N_1720);
nor U9123 (N_9123,N_939,N_898);
nor U9124 (N_9124,N_4119,N_3727);
xor U9125 (N_9125,N_543,N_353);
and U9126 (N_9126,N_3331,N_4200);
xnor U9127 (N_9127,N_4247,N_923);
xnor U9128 (N_9128,N_4734,N_396);
or U9129 (N_9129,N_2285,N_4707);
xor U9130 (N_9130,N_2278,N_2977);
xor U9131 (N_9131,N_3307,N_1062);
or U9132 (N_9132,N_2077,N_4483);
nor U9133 (N_9133,N_4956,N_581);
or U9134 (N_9134,N_1168,N_1672);
or U9135 (N_9135,N_2440,N_688);
or U9136 (N_9136,N_118,N_682);
nand U9137 (N_9137,N_1343,N_4685);
and U9138 (N_9138,N_1299,N_924);
nand U9139 (N_9139,N_4880,N_1885);
nand U9140 (N_9140,N_918,N_3698);
or U9141 (N_9141,N_593,N_2100);
or U9142 (N_9142,N_691,N_50);
nor U9143 (N_9143,N_4765,N_4399);
nor U9144 (N_9144,N_1443,N_4146);
xnor U9145 (N_9145,N_2506,N_2706);
and U9146 (N_9146,N_3526,N_1703);
nand U9147 (N_9147,N_3789,N_2758);
xnor U9148 (N_9148,N_3629,N_2289);
nand U9149 (N_9149,N_2999,N_47);
or U9150 (N_9150,N_4308,N_1862);
or U9151 (N_9151,N_1228,N_898);
and U9152 (N_9152,N_2565,N_451);
or U9153 (N_9153,N_3471,N_4067);
nand U9154 (N_9154,N_2236,N_4965);
nand U9155 (N_9155,N_3351,N_644);
xor U9156 (N_9156,N_4179,N_2189);
or U9157 (N_9157,N_4587,N_3152);
or U9158 (N_9158,N_146,N_3614);
and U9159 (N_9159,N_4231,N_3881);
xor U9160 (N_9160,N_3230,N_1353);
nor U9161 (N_9161,N_3461,N_1179);
or U9162 (N_9162,N_2762,N_2023);
nor U9163 (N_9163,N_3246,N_4929);
xor U9164 (N_9164,N_4549,N_2356);
and U9165 (N_9165,N_2734,N_386);
nor U9166 (N_9166,N_4792,N_3850);
xor U9167 (N_9167,N_1528,N_4673);
xnor U9168 (N_9168,N_1459,N_4718);
or U9169 (N_9169,N_945,N_1709);
and U9170 (N_9170,N_1718,N_4153);
and U9171 (N_9171,N_4090,N_2755);
or U9172 (N_9172,N_3095,N_1866);
or U9173 (N_9173,N_907,N_3897);
and U9174 (N_9174,N_2887,N_3326);
xor U9175 (N_9175,N_2604,N_4937);
nand U9176 (N_9176,N_1088,N_387);
and U9177 (N_9177,N_4499,N_266);
nor U9178 (N_9178,N_3537,N_128);
nor U9179 (N_9179,N_3564,N_1026);
nor U9180 (N_9180,N_1940,N_2095);
nand U9181 (N_9181,N_642,N_4638);
nor U9182 (N_9182,N_481,N_4793);
nor U9183 (N_9183,N_4913,N_3719);
nand U9184 (N_9184,N_4321,N_3121);
nor U9185 (N_9185,N_4421,N_355);
xor U9186 (N_9186,N_2100,N_3117);
or U9187 (N_9187,N_1395,N_656);
or U9188 (N_9188,N_4675,N_716);
or U9189 (N_9189,N_2429,N_551);
and U9190 (N_9190,N_663,N_3794);
and U9191 (N_9191,N_4432,N_851);
nand U9192 (N_9192,N_3707,N_4126);
xnor U9193 (N_9193,N_2352,N_4056);
or U9194 (N_9194,N_2405,N_415);
nand U9195 (N_9195,N_3461,N_1538);
xnor U9196 (N_9196,N_3942,N_2445);
and U9197 (N_9197,N_365,N_3080);
nor U9198 (N_9198,N_130,N_4482);
and U9199 (N_9199,N_2318,N_4221);
xnor U9200 (N_9200,N_212,N_753);
and U9201 (N_9201,N_1525,N_1976);
and U9202 (N_9202,N_4556,N_1029);
nor U9203 (N_9203,N_4052,N_2059);
xnor U9204 (N_9204,N_2784,N_914);
or U9205 (N_9205,N_136,N_4884);
and U9206 (N_9206,N_3205,N_1370);
nor U9207 (N_9207,N_4019,N_3462);
nand U9208 (N_9208,N_3238,N_3440);
and U9209 (N_9209,N_2102,N_739);
or U9210 (N_9210,N_4685,N_3248);
nand U9211 (N_9211,N_1188,N_3547);
nand U9212 (N_9212,N_3110,N_1938);
and U9213 (N_9213,N_233,N_2623);
and U9214 (N_9214,N_1555,N_2047);
and U9215 (N_9215,N_60,N_2392);
or U9216 (N_9216,N_2159,N_1755);
nor U9217 (N_9217,N_833,N_1849);
nor U9218 (N_9218,N_434,N_4582);
or U9219 (N_9219,N_349,N_2894);
or U9220 (N_9220,N_2667,N_1671);
and U9221 (N_9221,N_3727,N_561);
nor U9222 (N_9222,N_4809,N_2042);
and U9223 (N_9223,N_1734,N_1025);
xor U9224 (N_9224,N_3879,N_2548);
xnor U9225 (N_9225,N_3876,N_1791);
nor U9226 (N_9226,N_175,N_4227);
nor U9227 (N_9227,N_4193,N_3930);
nor U9228 (N_9228,N_3408,N_1858);
nor U9229 (N_9229,N_4791,N_4363);
and U9230 (N_9230,N_2860,N_60);
nor U9231 (N_9231,N_4410,N_1627);
or U9232 (N_9232,N_2219,N_3485);
xnor U9233 (N_9233,N_4532,N_2836);
nand U9234 (N_9234,N_3359,N_1850);
xnor U9235 (N_9235,N_2083,N_3576);
xnor U9236 (N_9236,N_4337,N_4067);
xor U9237 (N_9237,N_4418,N_4183);
or U9238 (N_9238,N_149,N_3267);
and U9239 (N_9239,N_1115,N_1077);
nor U9240 (N_9240,N_2237,N_184);
nor U9241 (N_9241,N_1987,N_1841);
xnor U9242 (N_9242,N_2090,N_3932);
or U9243 (N_9243,N_2527,N_2928);
xnor U9244 (N_9244,N_2639,N_2305);
xnor U9245 (N_9245,N_465,N_3411);
nor U9246 (N_9246,N_3546,N_4003);
nand U9247 (N_9247,N_1470,N_2015);
or U9248 (N_9248,N_3720,N_249);
nand U9249 (N_9249,N_3359,N_4791);
or U9250 (N_9250,N_1303,N_3169);
or U9251 (N_9251,N_3994,N_4424);
or U9252 (N_9252,N_1290,N_1462);
nor U9253 (N_9253,N_2056,N_1805);
xnor U9254 (N_9254,N_2340,N_4686);
and U9255 (N_9255,N_2531,N_135);
and U9256 (N_9256,N_4739,N_3355);
xor U9257 (N_9257,N_1403,N_835);
and U9258 (N_9258,N_3458,N_3337);
nand U9259 (N_9259,N_1554,N_3959);
and U9260 (N_9260,N_2633,N_1238);
or U9261 (N_9261,N_3148,N_1538);
or U9262 (N_9262,N_1215,N_3103);
nor U9263 (N_9263,N_4688,N_4545);
xor U9264 (N_9264,N_3046,N_3334);
nand U9265 (N_9265,N_615,N_1314);
nor U9266 (N_9266,N_692,N_2805);
xor U9267 (N_9267,N_2132,N_4248);
nor U9268 (N_9268,N_3608,N_902);
nand U9269 (N_9269,N_1920,N_3956);
and U9270 (N_9270,N_4615,N_928);
or U9271 (N_9271,N_2651,N_2530);
and U9272 (N_9272,N_2064,N_1950);
or U9273 (N_9273,N_1003,N_4227);
or U9274 (N_9274,N_1571,N_1443);
nor U9275 (N_9275,N_3861,N_4539);
and U9276 (N_9276,N_4382,N_1340);
or U9277 (N_9277,N_3110,N_2140);
nor U9278 (N_9278,N_1807,N_2164);
or U9279 (N_9279,N_1487,N_4540);
xnor U9280 (N_9280,N_223,N_101);
nor U9281 (N_9281,N_3330,N_1268);
nor U9282 (N_9282,N_2886,N_2922);
nand U9283 (N_9283,N_2678,N_1263);
or U9284 (N_9284,N_2086,N_4028);
nor U9285 (N_9285,N_3948,N_2468);
nand U9286 (N_9286,N_2155,N_4480);
and U9287 (N_9287,N_624,N_1997);
xor U9288 (N_9288,N_2589,N_1658);
xor U9289 (N_9289,N_4424,N_3753);
nor U9290 (N_9290,N_3201,N_2485);
nor U9291 (N_9291,N_3723,N_4103);
xnor U9292 (N_9292,N_1627,N_1761);
and U9293 (N_9293,N_133,N_2774);
and U9294 (N_9294,N_3561,N_3219);
and U9295 (N_9295,N_1841,N_836);
nand U9296 (N_9296,N_3653,N_4181);
nand U9297 (N_9297,N_182,N_3307);
nand U9298 (N_9298,N_3835,N_1868);
and U9299 (N_9299,N_326,N_3476);
or U9300 (N_9300,N_2961,N_2364);
or U9301 (N_9301,N_843,N_4500);
xor U9302 (N_9302,N_2194,N_2962);
nand U9303 (N_9303,N_1260,N_2905);
and U9304 (N_9304,N_4259,N_4703);
nor U9305 (N_9305,N_2132,N_4276);
and U9306 (N_9306,N_2599,N_1831);
or U9307 (N_9307,N_89,N_1764);
nand U9308 (N_9308,N_3637,N_4006);
xor U9309 (N_9309,N_4118,N_2834);
nand U9310 (N_9310,N_4999,N_4928);
and U9311 (N_9311,N_2895,N_2464);
and U9312 (N_9312,N_482,N_2009);
nand U9313 (N_9313,N_3037,N_2185);
and U9314 (N_9314,N_2553,N_4286);
or U9315 (N_9315,N_257,N_794);
and U9316 (N_9316,N_553,N_4472);
nor U9317 (N_9317,N_4504,N_4844);
nand U9318 (N_9318,N_2925,N_4385);
or U9319 (N_9319,N_4462,N_4667);
xnor U9320 (N_9320,N_2541,N_3478);
or U9321 (N_9321,N_498,N_3728);
nor U9322 (N_9322,N_4280,N_3584);
and U9323 (N_9323,N_3792,N_588);
nor U9324 (N_9324,N_1655,N_4394);
xnor U9325 (N_9325,N_1022,N_1360);
or U9326 (N_9326,N_4872,N_1131);
or U9327 (N_9327,N_1410,N_3901);
and U9328 (N_9328,N_1539,N_4484);
or U9329 (N_9329,N_1084,N_2377);
nor U9330 (N_9330,N_847,N_2657);
or U9331 (N_9331,N_730,N_552);
nor U9332 (N_9332,N_1131,N_1374);
nor U9333 (N_9333,N_2139,N_3020);
xor U9334 (N_9334,N_4543,N_4148);
and U9335 (N_9335,N_4294,N_4883);
nand U9336 (N_9336,N_998,N_69);
xor U9337 (N_9337,N_3138,N_1308);
nor U9338 (N_9338,N_3842,N_4196);
xor U9339 (N_9339,N_993,N_4244);
xor U9340 (N_9340,N_100,N_3575);
and U9341 (N_9341,N_4912,N_3845);
and U9342 (N_9342,N_4575,N_832);
xor U9343 (N_9343,N_4024,N_1302);
or U9344 (N_9344,N_4103,N_2407);
or U9345 (N_9345,N_1370,N_2388);
and U9346 (N_9346,N_2909,N_2536);
xor U9347 (N_9347,N_1965,N_1502);
nand U9348 (N_9348,N_190,N_3311);
and U9349 (N_9349,N_2335,N_1861);
or U9350 (N_9350,N_1269,N_3868);
or U9351 (N_9351,N_1866,N_3513);
nand U9352 (N_9352,N_1699,N_3527);
nor U9353 (N_9353,N_4721,N_1430);
nand U9354 (N_9354,N_1689,N_519);
nor U9355 (N_9355,N_810,N_4233);
xor U9356 (N_9356,N_4721,N_324);
or U9357 (N_9357,N_4884,N_360);
and U9358 (N_9358,N_3911,N_4668);
nor U9359 (N_9359,N_3596,N_1209);
nor U9360 (N_9360,N_4781,N_3601);
and U9361 (N_9361,N_4447,N_1512);
nor U9362 (N_9362,N_4157,N_113);
or U9363 (N_9363,N_3244,N_2105);
and U9364 (N_9364,N_2223,N_3752);
xnor U9365 (N_9365,N_3855,N_1070);
nand U9366 (N_9366,N_288,N_480);
or U9367 (N_9367,N_1821,N_386);
nand U9368 (N_9368,N_2405,N_1542);
or U9369 (N_9369,N_914,N_1041);
xor U9370 (N_9370,N_3254,N_818);
xnor U9371 (N_9371,N_4580,N_1686);
and U9372 (N_9372,N_1812,N_3168);
or U9373 (N_9373,N_125,N_2735);
nor U9374 (N_9374,N_3683,N_1150);
or U9375 (N_9375,N_4376,N_774);
xnor U9376 (N_9376,N_3657,N_4433);
xor U9377 (N_9377,N_2050,N_4853);
or U9378 (N_9378,N_220,N_4771);
xor U9379 (N_9379,N_1103,N_1960);
nand U9380 (N_9380,N_3549,N_2097);
nand U9381 (N_9381,N_1935,N_696);
nand U9382 (N_9382,N_4380,N_2185);
nand U9383 (N_9383,N_4800,N_825);
or U9384 (N_9384,N_3898,N_3969);
xnor U9385 (N_9385,N_2157,N_393);
and U9386 (N_9386,N_226,N_2348);
nor U9387 (N_9387,N_1776,N_3233);
and U9388 (N_9388,N_2656,N_3394);
xnor U9389 (N_9389,N_1191,N_2775);
nor U9390 (N_9390,N_4961,N_4528);
xnor U9391 (N_9391,N_4341,N_2275);
or U9392 (N_9392,N_805,N_1841);
or U9393 (N_9393,N_3922,N_911);
or U9394 (N_9394,N_2388,N_874);
and U9395 (N_9395,N_2492,N_670);
nand U9396 (N_9396,N_2013,N_3522);
nand U9397 (N_9397,N_4238,N_356);
or U9398 (N_9398,N_613,N_2629);
nor U9399 (N_9399,N_2432,N_955);
and U9400 (N_9400,N_4519,N_3069);
or U9401 (N_9401,N_4025,N_578);
and U9402 (N_9402,N_3892,N_4814);
nand U9403 (N_9403,N_3198,N_605);
nor U9404 (N_9404,N_893,N_3177);
or U9405 (N_9405,N_3721,N_1033);
or U9406 (N_9406,N_4561,N_2006);
nand U9407 (N_9407,N_1641,N_3813);
nor U9408 (N_9408,N_3583,N_579);
nor U9409 (N_9409,N_3794,N_616);
nand U9410 (N_9410,N_2654,N_2603);
nand U9411 (N_9411,N_2957,N_4776);
nor U9412 (N_9412,N_2726,N_280);
nor U9413 (N_9413,N_1790,N_3203);
xnor U9414 (N_9414,N_303,N_4638);
nand U9415 (N_9415,N_4414,N_1442);
and U9416 (N_9416,N_3957,N_1981);
nor U9417 (N_9417,N_1522,N_2909);
or U9418 (N_9418,N_149,N_10);
xor U9419 (N_9419,N_2489,N_916);
or U9420 (N_9420,N_60,N_3274);
and U9421 (N_9421,N_1422,N_4170);
and U9422 (N_9422,N_204,N_2407);
and U9423 (N_9423,N_1245,N_811);
nor U9424 (N_9424,N_3875,N_2940);
and U9425 (N_9425,N_1396,N_167);
and U9426 (N_9426,N_2285,N_1512);
or U9427 (N_9427,N_3693,N_1101);
xnor U9428 (N_9428,N_2272,N_2469);
and U9429 (N_9429,N_1498,N_4588);
or U9430 (N_9430,N_2896,N_4633);
nor U9431 (N_9431,N_2105,N_715);
xor U9432 (N_9432,N_1289,N_4154);
xor U9433 (N_9433,N_3084,N_2271);
xnor U9434 (N_9434,N_3306,N_3907);
and U9435 (N_9435,N_4682,N_605);
or U9436 (N_9436,N_845,N_1768);
or U9437 (N_9437,N_4447,N_47);
and U9438 (N_9438,N_4235,N_906);
and U9439 (N_9439,N_461,N_4300);
nand U9440 (N_9440,N_1203,N_31);
nor U9441 (N_9441,N_2091,N_2550);
or U9442 (N_9442,N_1165,N_4534);
nor U9443 (N_9443,N_4368,N_1537);
xnor U9444 (N_9444,N_3345,N_2203);
nor U9445 (N_9445,N_3953,N_1857);
nand U9446 (N_9446,N_4718,N_3204);
and U9447 (N_9447,N_1328,N_4004);
xor U9448 (N_9448,N_2037,N_1582);
nand U9449 (N_9449,N_4899,N_2856);
nand U9450 (N_9450,N_3871,N_3397);
nand U9451 (N_9451,N_152,N_2282);
xnor U9452 (N_9452,N_3942,N_1123);
nor U9453 (N_9453,N_274,N_1551);
and U9454 (N_9454,N_3361,N_929);
xor U9455 (N_9455,N_2633,N_3334);
or U9456 (N_9456,N_2188,N_4499);
xor U9457 (N_9457,N_1343,N_1757);
xnor U9458 (N_9458,N_191,N_2654);
nor U9459 (N_9459,N_3221,N_602);
or U9460 (N_9460,N_383,N_910);
or U9461 (N_9461,N_2988,N_1677);
nand U9462 (N_9462,N_4177,N_4485);
nor U9463 (N_9463,N_1793,N_1603);
or U9464 (N_9464,N_1223,N_866);
nand U9465 (N_9465,N_383,N_4941);
or U9466 (N_9466,N_4382,N_317);
and U9467 (N_9467,N_3544,N_4523);
and U9468 (N_9468,N_1209,N_133);
or U9469 (N_9469,N_4578,N_796);
or U9470 (N_9470,N_1253,N_3624);
xnor U9471 (N_9471,N_2390,N_3595);
or U9472 (N_9472,N_3330,N_2281);
nor U9473 (N_9473,N_272,N_1844);
and U9474 (N_9474,N_4300,N_1385);
nor U9475 (N_9475,N_2432,N_2084);
nand U9476 (N_9476,N_2050,N_762);
xor U9477 (N_9477,N_4865,N_3319);
and U9478 (N_9478,N_591,N_1214);
xnor U9479 (N_9479,N_4271,N_4354);
or U9480 (N_9480,N_271,N_4867);
xor U9481 (N_9481,N_354,N_4919);
nor U9482 (N_9482,N_3734,N_4802);
or U9483 (N_9483,N_2358,N_2514);
nor U9484 (N_9484,N_970,N_2447);
nand U9485 (N_9485,N_2548,N_662);
nand U9486 (N_9486,N_4571,N_3530);
and U9487 (N_9487,N_991,N_4985);
nor U9488 (N_9488,N_2904,N_3996);
nand U9489 (N_9489,N_4458,N_3885);
xor U9490 (N_9490,N_4278,N_1826);
nor U9491 (N_9491,N_4317,N_3646);
and U9492 (N_9492,N_4041,N_1486);
xor U9493 (N_9493,N_4300,N_1812);
and U9494 (N_9494,N_2367,N_4712);
nor U9495 (N_9495,N_3345,N_1671);
xor U9496 (N_9496,N_3361,N_2764);
nor U9497 (N_9497,N_286,N_187);
xnor U9498 (N_9498,N_3326,N_3223);
and U9499 (N_9499,N_1206,N_3141);
nand U9500 (N_9500,N_3917,N_2753);
or U9501 (N_9501,N_2242,N_2337);
xor U9502 (N_9502,N_3623,N_3219);
or U9503 (N_9503,N_4189,N_4805);
nand U9504 (N_9504,N_3556,N_53);
xnor U9505 (N_9505,N_1002,N_1988);
nand U9506 (N_9506,N_4846,N_18);
nor U9507 (N_9507,N_4745,N_1923);
or U9508 (N_9508,N_4788,N_4351);
and U9509 (N_9509,N_3480,N_4312);
nand U9510 (N_9510,N_519,N_4029);
xnor U9511 (N_9511,N_3016,N_3211);
xnor U9512 (N_9512,N_1848,N_4975);
nand U9513 (N_9513,N_2582,N_3200);
and U9514 (N_9514,N_3388,N_2932);
or U9515 (N_9515,N_1667,N_3007);
nor U9516 (N_9516,N_3871,N_144);
or U9517 (N_9517,N_1675,N_1913);
nor U9518 (N_9518,N_98,N_2361);
and U9519 (N_9519,N_3984,N_4020);
xnor U9520 (N_9520,N_1710,N_3740);
and U9521 (N_9521,N_2195,N_4540);
nand U9522 (N_9522,N_3560,N_579);
or U9523 (N_9523,N_3054,N_4797);
xnor U9524 (N_9524,N_1750,N_4402);
xnor U9525 (N_9525,N_2939,N_1761);
and U9526 (N_9526,N_3896,N_539);
or U9527 (N_9527,N_3505,N_2839);
and U9528 (N_9528,N_1857,N_4346);
nor U9529 (N_9529,N_311,N_2438);
nand U9530 (N_9530,N_3835,N_230);
nor U9531 (N_9531,N_2630,N_1951);
and U9532 (N_9532,N_4664,N_4423);
or U9533 (N_9533,N_3189,N_819);
or U9534 (N_9534,N_1886,N_867);
or U9535 (N_9535,N_3495,N_3001);
nand U9536 (N_9536,N_4226,N_3431);
nor U9537 (N_9537,N_1617,N_1451);
or U9538 (N_9538,N_900,N_1396);
nand U9539 (N_9539,N_3725,N_3270);
or U9540 (N_9540,N_1773,N_4085);
nand U9541 (N_9541,N_1866,N_1201);
nand U9542 (N_9542,N_4277,N_414);
nand U9543 (N_9543,N_1615,N_1451);
xnor U9544 (N_9544,N_3982,N_4281);
xnor U9545 (N_9545,N_366,N_1187);
nor U9546 (N_9546,N_1237,N_2948);
xnor U9547 (N_9547,N_4983,N_1417);
nand U9548 (N_9548,N_2337,N_3561);
nor U9549 (N_9549,N_1613,N_1386);
and U9550 (N_9550,N_618,N_2172);
nor U9551 (N_9551,N_4399,N_366);
or U9552 (N_9552,N_717,N_3279);
nand U9553 (N_9553,N_659,N_297);
or U9554 (N_9554,N_2807,N_1956);
xnor U9555 (N_9555,N_501,N_3647);
nand U9556 (N_9556,N_4375,N_4710);
and U9557 (N_9557,N_3276,N_4075);
nor U9558 (N_9558,N_4462,N_3287);
or U9559 (N_9559,N_186,N_1316);
nand U9560 (N_9560,N_897,N_668);
xnor U9561 (N_9561,N_4402,N_525);
nand U9562 (N_9562,N_3569,N_2157);
or U9563 (N_9563,N_2962,N_1580);
xor U9564 (N_9564,N_3390,N_952);
xnor U9565 (N_9565,N_3305,N_1954);
and U9566 (N_9566,N_3971,N_3172);
or U9567 (N_9567,N_1781,N_1336);
xor U9568 (N_9568,N_4338,N_2950);
nand U9569 (N_9569,N_346,N_4706);
nand U9570 (N_9570,N_3715,N_52);
or U9571 (N_9571,N_4357,N_507);
nor U9572 (N_9572,N_4824,N_708);
nand U9573 (N_9573,N_1045,N_1545);
or U9574 (N_9574,N_745,N_4139);
xor U9575 (N_9575,N_2123,N_4196);
xnor U9576 (N_9576,N_2793,N_3693);
xnor U9577 (N_9577,N_3815,N_1163);
and U9578 (N_9578,N_1131,N_3970);
nand U9579 (N_9579,N_2198,N_864);
and U9580 (N_9580,N_3345,N_967);
nor U9581 (N_9581,N_1724,N_30);
xnor U9582 (N_9582,N_437,N_2168);
xnor U9583 (N_9583,N_745,N_3062);
nor U9584 (N_9584,N_2560,N_929);
xnor U9585 (N_9585,N_384,N_1199);
xnor U9586 (N_9586,N_150,N_1729);
xor U9587 (N_9587,N_1394,N_610);
nor U9588 (N_9588,N_2307,N_1183);
and U9589 (N_9589,N_1729,N_3501);
nor U9590 (N_9590,N_2141,N_2893);
or U9591 (N_9591,N_4071,N_1053);
nor U9592 (N_9592,N_4383,N_331);
nand U9593 (N_9593,N_2328,N_1632);
nand U9594 (N_9594,N_3346,N_1699);
nor U9595 (N_9595,N_2914,N_4863);
nor U9596 (N_9596,N_3361,N_2623);
or U9597 (N_9597,N_3223,N_1192);
and U9598 (N_9598,N_3960,N_749);
or U9599 (N_9599,N_1172,N_2883);
and U9600 (N_9600,N_3314,N_4891);
xnor U9601 (N_9601,N_1177,N_4104);
and U9602 (N_9602,N_4406,N_4947);
and U9603 (N_9603,N_4354,N_4568);
and U9604 (N_9604,N_765,N_4110);
or U9605 (N_9605,N_2842,N_3405);
or U9606 (N_9606,N_1496,N_1943);
or U9607 (N_9607,N_3974,N_1189);
xnor U9608 (N_9608,N_4269,N_3133);
nor U9609 (N_9609,N_4366,N_2744);
nand U9610 (N_9610,N_1041,N_496);
or U9611 (N_9611,N_1871,N_248);
nor U9612 (N_9612,N_1254,N_302);
or U9613 (N_9613,N_752,N_200);
nand U9614 (N_9614,N_2012,N_3805);
xnor U9615 (N_9615,N_1618,N_1300);
or U9616 (N_9616,N_3457,N_1693);
xor U9617 (N_9617,N_3179,N_1123);
xnor U9618 (N_9618,N_792,N_2733);
nand U9619 (N_9619,N_2247,N_1743);
nor U9620 (N_9620,N_2676,N_4558);
and U9621 (N_9621,N_3892,N_3702);
nor U9622 (N_9622,N_4376,N_339);
or U9623 (N_9623,N_3629,N_3538);
or U9624 (N_9624,N_1726,N_1966);
xnor U9625 (N_9625,N_905,N_569);
nand U9626 (N_9626,N_2144,N_916);
and U9627 (N_9627,N_2632,N_2876);
nor U9628 (N_9628,N_3830,N_3853);
nand U9629 (N_9629,N_4234,N_4256);
or U9630 (N_9630,N_2776,N_813);
xor U9631 (N_9631,N_4850,N_2820);
nor U9632 (N_9632,N_2524,N_4366);
xor U9633 (N_9633,N_1989,N_4681);
xor U9634 (N_9634,N_4660,N_4201);
or U9635 (N_9635,N_1904,N_4972);
and U9636 (N_9636,N_1331,N_1406);
nand U9637 (N_9637,N_3548,N_2351);
nand U9638 (N_9638,N_3451,N_3050);
nand U9639 (N_9639,N_2571,N_650);
and U9640 (N_9640,N_3988,N_2222);
and U9641 (N_9641,N_3849,N_4924);
nand U9642 (N_9642,N_112,N_3701);
nand U9643 (N_9643,N_1983,N_4750);
or U9644 (N_9644,N_1963,N_931);
nor U9645 (N_9645,N_666,N_4742);
and U9646 (N_9646,N_574,N_4380);
and U9647 (N_9647,N_683,N_2796);
xor U9648 (N_9648,N_4510,N_4700);
xor U9649 (N_9649,N_2142,N_3221);
and U9650 (N_9650,N_2125,N_917);
and U9651 (N_9651,N_812,N_4874);
or U9652 (N_9652,N_666,N_847);
and U9653 (N_9653,N_2125,N_806);
nor U9654 (N_9654,N_1461,N_1620);
or U9655 (N_9655,N_3374,N_872);
or U9656 (N_9656,N_265,N_4826);
nor U9657 (N_9657,N_3633,N_2736);
or U9658 (N_9658,N_3787,N_4937);
xnor U9659 (N_9659,N_3148,N_4222);
nand U9660 (N_9660,N_4434,N_1084);
nand U9661 (N_9661,N_1666,N_3985);
nor U9662 (N_9662,N_2845,N_2969);
xor U9663 (N_9663,N_3032,N_2643);
and U9664 (N_9664,N_1605,N_2248);
nor U9665 (N_9665,N_3501,N_1736);
and U9666 (N_9666,N_1159,N_3351);
nand U9667 (N_9667,N_3254,N_3770);
and U9668 (N_9668,N_2682,N_1745);
or U9669 (N_9669,N_3964,N_1968);
or U9670 (N_9670,N_4308,N_219);
xnor U9671 (N_9671,N_147,N_2804);
or U9672 (N_9672,N_410,N_2004);
nand U9673 (N_9673,N_1362,N_1089);
nor U9674 (N_9674,N_776,N_4406);
and U9675 (N_9675,N_3843,N_3177);
or U9676 (N_9676,N_2637,N_2809);
nor U9677 (N_9677,N_4672,N_3737);
xnor U9678 (N_9678,N_2935,N_4373);
nand U9679 (N_9679,N_3492,N_4966);
nand U9680 (N_9680,N_2091,N_186);
nand U9681 (N_9681,N_4769,N_112);
xor U9682 (N_9682,N_1013,N_3550);
or U9683 (N_9683,N_2629,N_1373);
and U9684 (N_9684,N_4860,N_2062);
nor U9685 (N_9685,N_1521,N_2396);
and U9686 (N_9686,N_3369,N_2085);
or U9687 (N_9687,N_4930,N_2604);
nand U9688 (N_9688,N_242,N_749);
or U9689 (N_9689,N_3212,N_1487);
nor U9690 (N_9690,N_3008,N_1277);
and U9691 (N_9691,N_254,N_1690);
nor U9692 (N_9692,N_2866,N_3290);
and U9693 (N_9693,N_2881,N_785);
and U9694 (N_9694,N_3126,N_1648);
and U9695 (N_9695,N_4966,N_4301);
nand U9696 (N_9696,N_1822,N_1992);
nor U9697 (N_9697,N_4312,N_3642);
and U9698 (N_9698,N_1332,N_1777);
nand U9699 (N_9699,N_2081,N_367);
xnor U9700 (N_9700,N_2919,N_90);
xnor U9701 (N_9701,N_336,N_345);
and U9702 (N_9702,N_680,N_3345);
xor U9703 (N_9703,N_1708,N_1341);
nor U9704 (N_9704,N_246,N_1482);
and U9705 (N_9705,N_3870,N_3940);
nor U9706 (N_9706,N_4919,N_3584);
or U9707 (N_9707,N_1262,N_3805);
xor U9708 (N_9708,N_2555,N_4137);
xor U9709 (N_9709,N_2149,N_2276);
nand U9710 (N_9710,N_58,N_2139);
or U9711 (N_9711,N_405,N_558);
nor U9712 (N_9712,N_2098,N_3566);
nor U9713 (N_9713,N_4144,N_3474);
xor U9714 (N_9714,N_2980,N_44);
and U9715 (N_9715,N_4324,N_444);
xnor U9716 (N_9716,N_3171,N_2194);
and U9717 (N_9717,N_2724,N_4986);
xnor U9718 (N_9718,N_875,N_4467);
nand U9719 (N_9719,N_4259,N_4625);
and U9720 (N_9720,N_1575,N_627);
nor U9721 (N_9721,N_569,N_674);
xnor U9722 (N_9722,N_1280,N_4725);
nor U9723 (N_9723,N_4057,N_931);
nand U9724 (N_9724,N_4331,N_2717);
nand U9725 (N_9725,N_2675,N_3926);
nand U9726 (N_9726,N_1977,N_530);
and U9727 (N_9727,N_213,N_4662);
and U9728 (N_9728,N_1549,N_4933);
and U9729 (N_9729,N_776,N_4615);
nand U9730 (N_9730,N_3093,N_2306);
xnor U9731 (N_9731,N_1491,N_924);
nor U9732 (N_9732,N_417,N_201);
or U9733 (N_9733,N_4015,N_901);
nand U9734 (N_9734,N_2246,N_4731);
and U9735 (N_9735,N_2709,N_1023);
and U9736 (N_9736,N_1483,N_952);
or U9737 (N_9737,N_4364,N_1109);
xor U9738 (N_9738,N_307,N_4132);
and U9739 (N_9739,N_4770,N_3300);
and U9740 (N_9740,N_3690,N_2132);
nand U9741 (N_9741,N_4447,N_1142);
or U9742 (N_9742,N_3548,N_524);
or U9743 (N_9743,N_2239,N_2037);
nor U9744 (N_9744,N_3621,N_4584);
nor U9745 (N_9745,N_4486,N_1487);
xnor U9746 (N_9746,N_846,N_4630);
nor U9747 (N_9747,N_4359,N_4976);
and U9748 (N_9748,N_2106,N_733);
nand U9749 (N_9749,N_1894,N_2012);
and U9750 (N_9750,N_1381,N_979);
nor U9751 (N_9751,N_4902,N_4786);
xor U9752 (N_9752,N_1912,N_4738);
or U9753 (N_9753,N_2581,N_2183);
or U9754 (N_9754,N_1223,N_1344);
or U9755 (N_9755,N_3278,N_3981);
nand U9756 (N_9756,N_1508,N_3046);
xnor U9757 (N_9757,N_4976,N_3590);
or U9758 (N_9758,N_4905,N_2091);
nor U9759 (N_9759,N_3524,N_4298);
xnor U9760 (N_9760,N_787,N_250);
or U9761 (N_9761,N_29,N_1945);
nor U9762 (N_9762,N_3250,N_1048);
and U9763 (N_9763,N_1888,N_1733);
and U9764 (N_9764,N_843,N_2954);
nor U9765 (N_9765,N_2938,N_1148);
nor U9766 (N_9766,N_3840,N_1128);
xor U9767 (N_9767,N_4975,N_2872);
xor U9768 (N_9768,N_4709,N_4147);
xor U9769 (N_9769,N_1468,N_1803);
or U9770 (N_9770,N_4821,N_1500);
xnor U9771 (N_9771,N_3970,N_1520);
or U9772 (N_9772,N_4717,N_4086);
and U9773 (N_9773,N_3126,N_1907);
xor U9774 (N_9774,N_3115,N_2182);
and U9775 (N_9775,N_3232,N_4928);
nor U9776 (N_9776,N_2813,N_1740);
or U9777 (N_9777,N_3024,N_3259);
and U9778 (N_9778,N_2606,N_3689);
nand U9779 (N_9779,N_645,N_4546);
xnor U9780 (N_9780,N_2898,N_4651);
and U9781 (N_9781,N_1290,N_1489);
and U9782 (N_9782,N_3217,N_3142);
nand U9783 (N_9783,N_4184,N_2116);
nand U9784 (N_9784,N_1972,N_3052);
nand U9785 (N_9785,N_4449,N_1507);
nor U9786 (N_9786,N_4320,N_4118);
xor U9787 (N_9787,N_935,N_1187);
nand U9788 (N_9788,N_1711,N_4900);
nor U9789 (N_9789,N_3441,N_2915);
nand U9790 (N_9790,N_4575,N_2177);
and U9791 (N_9791,N_4395,N_1166);
or U9792 (N_9792,N_3891,N_4405);
or U9793 (N_9793,N_2527,N_899);
or U9794 (N_9794,N_594,N_984);
and U9795 (N_9795,N_2391,N_159);
or U9796 (N_9796,N_1000,N_4846);
and U9797 (N_9797,N_3500,N_4899);
and U9798 (N_9798,N_3741,N_2874);
or U9799 (N_9799,N_2471,N_1366);
and U9800 (N_9800,N_4013,N_653);
nand U9801 (N_9801,N_2533,N_3223);
nand U9802 (N_9802,N_120,N_4680);
nor U9803 (N_9803,N_2657,N_4413);
nor U9804 (N_9804,N_2239,N_4526);
or U9805 (N_9805,N_493,N_4961);
nor U9806 (N_9806,N_200,N_431);
nor U9807 (N_9807,N_2568,N_3937);
nand U9808 (N_9808,N_1205,N_2498);
xnor U9809 (N_9809,N_2915,N_815);
xnor U9810 (N_9810,N_4784,N_1953);
nand U9811 (N_9811,N_3887,N_2715);
xor U9812 (N_9812,N_2089,N_3604);
or U9813 (N_9813,N_1934,N_4333);
and U9814 (N_9814,N_738,N_2255);
or U9815 (N_9815,N_278,N_3952);
and U9816 (N_9816,N_106,N_2423);
and U9817 (N_9817,N_4383,N_4910);
nand U9818 (N_9818,N_3544,N_4297);
or U9819 (N_9819,N_580,N_3418);
and U9820 (N_9820,N_2273,N_1734);
nand U9821 (N_9821,N_4486,N_3234);
xor U9822 (N_9822,N_2031,N_402);
and U9823 (N_9823,N_1346,N_4863);
and U9824 (N_9824,N_742,N_1884);
or U9825 (N_9825,N_2034,N_567);
and U9826 (N_9826,N_426,N_3312);
or U9827 (N_9827,N_1190,N_4795);
or U9828 (N_9828,N_1887,N_3712);
and U9829 (N_9829,N_4954,N_3055);
nor U9830 (N_9830,N_4287,N_2846);
xor U9831 (N_9831,N_2004,N_2298);
nand U9832 (N_9832,N_1406,N_3035);
nor U9833 (N_9833,N_4436,N_4207);
nor U9834 (N_9834,N_1997,N_2114);
or U9835 (N_9835,N_2501,N_4007);
nand U9836 (N_9836,N_487,N_4042);
or U9837 (N_9837,N_567,N_663);
xnor U9838 (N_9838,N_4430,N_4444);
and U9839 (N_9839,N_3594,N_1251);
or U9840 (N_9840,N_4927,N_3153);
or U9841 (N_9841,N_489,N_1720);
or U9842 (N_9842,N_2258,N_1349);
nor U9843 (N_9843,N_4019,N_2675);
or U9844 (N_9844,N_2084,N_4216);
and U9845 (N_9845,N_2393,N_4570);
and U9846 (N_9846,N_1328,N_2041);
xor U9847 (N_9847,N_1,N_4237);
and U9848 (N_9848,N_252,N_433);
xor U9849 (N_9849,N_1296,N_3757);
nand U9850 (N_9850,N_1316,N_4142);
nand U9851 (N_9851,N_2473,N_2258);
xor U9852 (N_9852,N_2287,N_4814);
nor U9853 (N_9853,N_1927,N_3964);
or U9854 (N_9854,N_2918,N_4491);
nand U9855 (N_9855,N_3889,N_4634);
xnor U9856 (N_9856,N_228,N_3133);
nand U9857 (N_9857,N_3612,N_2472);
nor U9858 (N_9858,N_0,N_905);
nor U9859 (N_9859,N_4848,N_1564);
or U9860 (N_9860,N_3028,N_3237);
and U9861 (N_9861,N_3968,N_3059);
and U9862 (N_9862,N_3114,N_4532);
nand U9863 (N_9863,N_2709,N_4682);
or U9864 (N_9864,N_1509,N_3274);
and U9865 (N_9865,N_3899,N_1287);
nor U9866 (N_9866,N_3237,N_44);
or U9867 (N_9867,N_64,N_3046);
nor U9868 (N_9868,N_1422,N_2396);
nor U9869 (N_9869,N_2477,N_3803);
nand U9870 (N_9870,N_1414,N_2971);
and U9871 (N_9871,N_1170,N_2672);
nand U9872 (N_9872,N_4297,N_1590);
and U9873 (N_9873,N_561,N_4903);
nand U9874 (N_9874,N_4835,N_3452);
and U9875 (N_9875,N_171,N_4306);
or U9876 (N_9876,N_4511,N_3566);
nor U9877 (N_9877,N_4122,N_2855);
and U9878 (N_9878,N_682,N_1281);
or U9879 (N_9879,N_4451,N_2377);
nor U9880 (N_9880,N_3226,N_3882);
nand U9881 (N_9881,N_837,N_1396);
nor U9882 (N_9882,N_3473,N_4706);
and U9883 (N_9883,N_1009,N_3976);
nor U9884 (N_9884,N_4755,N_1394);
nand U9885 (N_9885,N_4375,N_946);
nand U9886 (N_9886,N_4725,N_3494);
xor U9887 (N_9887,N_369,N_2049);
xor U9888 (N_9888,N_2869,N_2893);
nand U9889 (N_9889,N_3975,N_3330);
and U9890 (N_9890,N_1542,N_4445);
or U9891 (N_9891,N_1000,N_3063);
or U9892 (N_9892,N_686,N_187);
xnor U9893 (N_9893,N_690,N_2391);
xnor U9894 (N_9894,N_3668,N_1761);
or U9895 (N_9895,N_1437,N_215);
and U9896 (N_9896,N_3185,N_1049);
nand U9897 (N_9897,N_4588,N_2160);
xnor U9898 (N_9898,N_1108,N_194);
xnor U9899 (N_9899,N_3400,N_1002);
nor U9900 (N_9900,N_2896,N_1068);
xnor U9901 (N_9901,N_2934,N_4211);
xor U9902 (N_9902,N_3880,N_2567);
xnor U9903 (N_9903,N_1596,N_929);
nor U9904 (N_9904,N_1377,N_3408);
or U9905 (N_9905,N_2167,N_3751);
nand U9906 (N_9906,N_3552,N_2695);
or U9907 (N_9907,N_4930,N_2483);
and U9908 (N_9908,N_4160,N_3965);
nor U9909 (N_9909,N_2999,N_2988);
or U9910 (N_9910,N_561,N_1690);
xor U9911 (N_9911,N_1720,N_3760);
or U9912 (N_9912,N_3689,N_4502);
nand U9913 (N_9913,N_1952,N_1467);
and U9914 (N_9914,N_315,N_3768);
or U9915 (N_9915,N_2886,N_3029);
nand U9916 (N_9916,N_626,N_1867);
and U9917 (N_9917,N_4047,N_2397);
or U9918 (N_9918,N_4460,N_1450);
xnor U9919 (N_9919,N_2518,N_2807);
xnor U9920 (N_9920,N_1621,N_457);
and U9921 (N_9921,N_1707,N_4009);
nor U9922 (N_9922,N_586,N_4690);
nor U9923 (N_9923,N_2379,N_2880);
xnor U9924 (N_9924,N_2035,N_3188);
xor U9925 (N_9925,N_341,N_4946);
nor U9926 (N_9926,N_3248,N_1050);
and U9927 (N_9927,N_1933,N_2621);
and U9928 (N_9928,N_678,N_2611);
xor U9929 (N_9929,N_143,N_4465);
nand U9930 (N_9930,N_1331,N_3245);
nand U9931 (N_9931,N_3280,N_538);
or U9932 (N_9932,N_3698,N_1370);
nand U9933 (N_9933,N_1112,N_584);
nor U9934 (N_9934,N_1418,N_209);
nor U9935 (N_9935,N_277,N_823);
and U9936 (N_9936,N_2915,N_1633);
xnor U9937 (N_9937,N_1669,N_2971);
and U9938 (N_9938,N_3576,N_1733);
nand U9939 (N_9939,N_4611,N_2225);
nand U9940 (N_9940,N_885,N_2508);
and U9941 (N_9941,N_994,N_494);
xnor U9942 (N_9942,N_4978,N_3749);
xnor U9943 (N_9943,N_4692,N_4023);
or U9944 (N_9944,N_3395,N_1917);
nand U9945 (N_9945,N_4563,N_1011);
and U9946 (N_9946,N_2464,N_1300);
xnor U9947 (N_9947,N_1187,N_2542);
or U9948 (N_9948,N_4295,N_4387);
and U9949 (N_9949,N_1132,N_3800);
nand U9950 (N_9950,N_3137,N_3465);
or U9951 (N_9951,N_660,N_1041);
or U9952 (N_9952,N_4453,N_4210);
nor U9953 (N_9953,N_2373,N_879);
or U9954 (N_9954,N_950,N_292);
or U9955 (N_9955,N_3573,N_699);
nand U9956 (N_9956,N_2651,N_3353);
and U9957 (N_9957,N_4930,N_1740);
xor U9958 (N_9958,N_883,N_3543);
nand U9959 (N_9959,N_4608,N_3692);
or U9960 (N_9960,N_4984,N_4232);
nor U9961 (N_9961,N_3076,N_2070);
xor U9962 (N_9962,N_4445,N_1915);
nand U9963 (N_9963,N_3791,N_2347);
xor U9964 (N_9964,N_1752,N_3671);
xor U9965 (N_9965,N_3940,N_4501);
or U9966 (N_9966,N_4085,N_2260);
or U9967 (N_9967,N_3243,N_2082);
and U9968 (N_9968,N_297,N_2697);
or U9969 (N_9969,N_3780,N_391);
and U9970 (N_9970,N_1201,N_583);
nand U9971 (N_9971,N_309,N_2158);
nor U9972 (N_9972,N_608,N_879);
and U9973 (N_9973,N_992,N_4798);
xnor U9974 (N_9974,N_947,N_1450);
and U9975 (N_9975,N_4333,N_861);
nor U9976 (N_9976,N_3196,N_935);
xor U9977 (N_9977,N_2602,N_2692);
xor U9978 (N_9978,N_1467,N_4282);
or U9979 (N_9979,N_3462,N_1786);
and U9980 (N_9980,N_1771,N_3570);
xor U9981 (N_9981,N_4675,N_4007);
xor U9982 (N_9982,N_2967,N_3282);
xnor U9983 (N_9983,N_4277,N_1699);
nand U9984 (N_9984,N_1857,N_2579);
xnor U9985 (N_9985,N_1583,N_86);
nor U9986 (N_9986,N_3885,N_850);
nor U9987 (N_9987,N_3961,N_2161);
or U9988 (N_9988,N_4746,N_1587);
and U9989 (N_9989,N_3120,N_4750);
nand U9990 (N_9990,N_3260,N_4336);
and U9991 (N_9991,N_4591,N_4935);
xnor U9992 (N_9992,N_1473,N_3652);
and U9993 (N_9993,N_3449,N_1556);
xor U9994 (N_9994,N_2821,N_1924);
nand U9995 (N_9995,N_4301,N_2876);
nor U9996 (N_9996,N_3124,N_2062);
and U9997 (N_9997,N_3109,N_1918);
or U9998 (N_9998,N_1271,N_1911);
nor U9999 (N_9999,N_227,N_3485);
or U10000 (N_10000,N_6197,N_9685);
or U10001 (N_10001,N_7100,N_9905);
nand U10002 (N_10002,N_5151,N_7161);
and U10003 (N_10003,N_8803,N_8374);
nor U10004 (N_10004,N_9638,N_8731);
nor U10005 (N_10005,N_9004,N_5883);
nand U10006 (N_10006,N_5892,N_8403);
and U10007 (N_10007,N_6805,N_5962);
nor U10008 (N_10008,N_9272,N_9881);
xor U10009 (N_10009,N_9460,N_9109);
xor U10010 (N_10010,N_7838,N_9558);
nor U10011 (N_10011,N_6516,N_9320);
nor U10012 (N_10012,N_6084,N_7493);
xnor U10013 (N_10013,N_7480,N_7785);
and U10014 (N_10014,N_5040,N_9226);
or U10015 (N_10015,N_7120,N_5495);
nor U10016 (N_10016,N_9151,N_8787);
nand U10017 (N_10017,N_7453,N_6377);
nor U10018 (N_10018,N_5685,N_5445);
and U10019 (N_10019,N_8583,N_5886);
nor U10020 (N_10020,N_7477,N_6741);
and U10021 (N_10021,N_8580,N_5055);
nand U10022 (N_10022,N_6589,N_8231);
or U10023 (N_10023,N_5468,N_6665);
and U10024 (N_10024,N_7526,N_9008);
or U10025 (N_10025,N_5913,N_5382);
or U10026 (N_10026,N_7651,N_6546);
and U10027 (N_10027,N_8571,N_8527);
nand U10028 (N_10028,N_7371,N_8842);
xor U10029 (N_10029,N_8030,N_7322);
or U10030 (N_10030,N_5760,N_9346);
xnor U10031 (N_10031,N_5558,N_8483);
or U10032 (N_10032,N_8261,N_5849);
and U10033 (N_10033,N_7299,N_5416);
or U10034 (N_10034,N_6469,N_8779);
or U10035 (N_10035,N_8558,N_7311);
and U10036 (N_10036,N_9165,N_9943);
and U10037 (N_10037,N_8885,N_7321);
and U10038 (N_10038,N_5260,N_9582);
xnor U10039 (N_10039,N_8427,N_6512);
nand U10040 (N_10040,N_5718,N_9712);
or U10041 (N_10041,N_6398,N_9751);
nor U10042 (N_10042,N_6802,N_5606);
nor U10043 (N_10043,N_8509,N_7255);
nand U10044 (N_10044,N_9794,N_5610);
nand U10045 (N_10045,N_9065,N_6270);
nor U10046 (N_10046,N_5430,N_6700);
or U10047 (N_10047,N_6224,N_7197);
nor U10048 (N_10048,N_9395,N_7714);
and U10049 (N_10049,N_7980,N_8532);
xnor U10050 (N_10050,N_7664,N_7217);
xor U10051 (N_10051,N_6775,N_8931);
xnor U10052 (N_10052,N_8220,N_5620);
or U10053 (N_10053,N_8704,N_8080);
nor U10054 (N_10054,N_7774,N_6427);
and U10055 (N_10055,N_7022,N_5363);
nand U10056 (N_10056,N_8573,N_5028);
or U10057 (N_10057,N_8518,N_7695);
or U10058 (N_10058,N_7642,N_8256);
and U10059 (N_10059,N_8965,N_9351);
and U10060 (N_10060,N_7445,N_5176);
or U10061 (N_10061,N_8912,N_8841);
xor U10062 (N_10062,N_7611,N_7247);
nand U10063 (N_10063,N_8560,N_8901);
and U10064 (N_10064,N_5431,N_7237);
nor U10065 (N_10065,N_8782,N_5941);
and U10066 (N_10066,N_6361,N_5153);
nor U10067 (N_10067,N_9642,N_7124);
and U10068 (N_10068,N_7772,N_9188);
nor U10069 (N_10069,N_9031,N_5821);
nor U10070 (N_10070,N_8250,N_5340);
nor U10071 (N_10071,N_5129,N_5133);
xor U10072 (N_10072,N_8794,N_7581);
nand U10073 (N_10073,N_6479,N_7298);
and U10074 (N_10074,N_6955,N_5180);
nor U10075 (N_10075,N_8380,N_5034);
nor U10076 (N_10076,N_6864,N_5370);
nand U10077 (N_10077,N_8388,N_7518);
nand U10078 (N_10078,N_9365,N_9090);
xor U10079 (N_10079,N_8505,N_7344);
nand U10080 (N_10080,N_5281,N_5599);
nor U10081 (N_10081,N_8165,N_5625);
xor U10082 (N_10082,N_9867,N_5011);
or U10083 (N_10083,N_7674,N_6106);
or U10084 (N_10084,N_6744,N_8740);
or U10085 (N_10085,N_6116,N_9883);
nand U10086 (N_10086,N_5504,N_9451);
and U10087 (N_10087,N_6140,N_5015);
nand U10088 (N_10088,N_5572,N_7656);
xor U10089 (N_10089,N_6129,N_6966);
and U10090 (N_10090,N_9472,N_7576);
nor U10091 (N_10091,N_5778,N_9868);
and U10092 (N_10092,N_5697,N_6482);
or U10093 (N_10093,N_8185,N_7654);
or U10094 (N_10094,N_9717,N_7083);
or U10095 (N_10095,N_6736,N_7448);
xor U10096 (N_10096,N_5613,N_8265);
and U10097 (N_10097,N_5292,N_7349);
xor U10098 (N_10098,N_5768,N_6111);
xnor U10099 (N_10099,N_5698,N_5302);
or U10100 (N_10100,N_9430,N_8125);
xor U10101 (N_10101,N_8923,N_7951);
nand U10102 (N_10102,N_7134,N_7122);
nor U10103 (N_10103,N_5604,N_5914);
and U10104 (N_10104,N_9819,N_8652);
or U10105 (N_10105,N_5319,N_8106);
nor U10106 (N_10106,N_5228,N_7037);
nand U10107 (N_10107,N_9184,N_5870);
or U10108 (N_10108,N_5257,N_9588);
and U10109 (N_10109,N_6010,N_6352);
nand U10110 (N_10110,N_5123,N_9984);
or U10111 (N_10111,N_9982,N_9174);
nand U10112 (N_10112,N_7240,N_7818);
and U10113 (N_10113,N_6356,N_8602);
or U10114 (N_10114,N_8755,N_5071);
nand U10115 (N_10115,N_8835,N_6409);
and U10116 (N_10116,N_6752,N_7092);
or U10117 (N_10117,N_8476,N_5823);
nand U10118 (N_10118,N_9981,N_8371);
and U10119 (N_10119,N_5921,N_5038);
nand U10120 (N_10120,N_6652,N_7854);
nor U10121 (N_10121,N_8605,N_6450);
nor U10122 (N_10122,N_6227,N_9745);
nand U10123 (N_10123,N_7631,N_9670);
or U10124 (N_10124,N_8420,N_5943);
nand U10125 (N_10125,N_9371,N_8205);
and U10126 (N_10126,N_7606,N_9809);
nor U10127 (N_10127,N_7170,N_8541);
nand U10128 (N_10128,N_7814,N_7905);
or U10129 (N_10129,N_6251,N_6827);
and U10130 (N_10130,N_9534,N_5820);
nor U10131 (N_10131,N_6294,N_7175);
and U10132 (N_10132,N_5414,N_7372);
nor U10133 (N_10133,N_8490,N_8921);
nand U10134 (N_10134,N_6598,N_6221);
nor U10135 (N_10135,N_6009,N_7253);
and U10136 (N_10136,N_9185,N_6000);
or U10137 (N_10137,N_5851,N_6202);
nand U10138 (N_10138,N_5749,N_6400);
and U10139 (N_10139,N_8131,N_5701);
nor U10140 (N_10140,N_9650,N_7984);
nor U10141 (N_10141,N_5287,N_9707);
and U10142 (N_10142,N_5835,N_5238);
or U10143 (N_10143,N_7358,N_6017);
xnor U10144 (N_10144,N_7080,N_6036);
xnor U10145 (N_10145,N_6880,N_5764);
nand U10146 (N_10146,N_8300,N_8935);
xor U10147 (N_10147,N_8500,N_9514);
nor U10148 (N_10148,N_6759,N_7140);
xnor U10149 (N_10149,N_6281,N_5312);
or U10150 (N_10150,N_6707,N_7045);
or U10151 (N_10151,N_7435,N_9845);
or U10152 (N_10152,N_8097,N_8723);
nand U10153 (N_10153,N_5479,N_9572);
or U10154 (N_10154,N_6905,N_5376);
nor U10155 (N_10155,N_5113,N_5345);
and U10156 (N_10156,N_9948,N_5237);
or U10157 (N_10157,N_5065,N_8746);
or U10158 (N_10158,N_9166,N_9137);
and U10159 (N_10159,N_5656,N_8273);
nand U10160 (N_10160,N_5548,N_6021);
nor U10161 (N_10161,N_8411,N_9741);
nand U10162 (N_10162,N_5809,N_7455);
xor U10163 (N_10163,N_6088,N_8737);
and U10164 (N_10164,N_5173,N_5608);
or U10165 (N_10165,N_6172,N_8795);
and U10166 (N_10166,N_8089,N_5198);
and U10167 (N_10167,N_8663,N_8710);
xnor U10168 (N_10168,N_7810,N_5958);
xor U10169 (N_10169,N_7213,N_5093);
and U10170 (N_10170,N_6175,N_6881);
xor U10171 (N_10171,N_8175,N_8073);
nor U10172 (N_10172,N_9313,N_8466);
nand U10173 (N_10173,N_6341,N_5513);
or U10174 (N_10174,N_9202,N_8918);
nand U10175 (N_10175,N_7042,N_5806);
xor U10176 (N_10176,N_9789,N_9459);
or U10177 (N_10177,N_9721,N_6349);
nand U10178 (N_10178,N_8075,N_9079);
and U10179 (N_10179,N_6991,N_7306);
xor U10180 (N_10180,N_9263,N_6641);
or U10181 (N_10181,N_8384,N_5702);
nor U10182 (N_10182,N_5137,N_7742);
nand U10183 (N_10183,N_9041,N_5890);
nor U10184 (N_10184,N_8625,N_9220);
and U10185 (N_10185,N_9922,N_5726);
nand U10186 (N_10186,N_6948,N_7797);
and U10187 (N_10187,N_5986,N_8986);
nor U10188 (N_10188,N_7677,N_5374);
xnor U10189 (N_10189,N_6074,N_5236);
and U10190 (N_10190,N_9739,N_9835);
xor U10191 (N_10191,N_6860,N_5335);
xor U10192 (N_10192,N_9468,N_9016);
xor U10193 (N_10193,N_7385,N_5754);
or U10194 (N_10194,N_6166,N_8489);
and U10195 (N_10195,N_9470,N_5649);
xnor U10196 (N_10196,N_6099,N_5089);
nand U10197 (N_10197,N_5163,N_6455);
or U10198 (N_10198,N_9000,N_8517);
xnor U10199 (N_10199,N_9482,N_9139);
nand U10200 (N_10200,N_6280,N_7738);
and U10201 (N_10201,N_8736,N_7062);
or U10202 (N_10202,N_6907,N_7947);
or U10203 (N_10203,N_6984,N_7260);
and U10204 (N_10204,N_6135,N_9034);
xor U10205 (N_10205,N_6149,N_9337);
or U10206 (N_10206,N_5602,N_8285);
and U10207 (N_10207,N_9005,N_6298);
nand U10208 (N_10208,N_6842,N_5868);
xnor U10209 (N_10209,N_5160,N_6791);
nor U10210 (N_10210,N_9306,N_7064);
nand U10211 (N_10211,N_7692,N_8152);
xor U10212 (N_10212,N_6617,N_5574);
or U10213 (N_10213,N_7939,N_7804);
nor U10214 (N_10214,N_5932,N_9528);
nor U10215 (N_10215,N_9757,N_7625);
nor U10216 (N_10216,N_7816,N_9287);
xor U10217 (N_10217,N_6193,N_6345);
xor U10218 (N_10218,N_8648,N_7820);
xor U10219 (N_10219,N_8306,N_7672);
or U10220 (N_10220,N_8393,N_8562);
xor U10221 (N_10221,N_7932,N_6423);
nor U10222 (N_10222,N_5818,N_8790);
xnor U10223 (N_10223,N_5188,N_7317);
or U10224 (N_10224,N_8235,N_6530);
xor U10225 (N_10225,N_6323,N_8099);
nand U10226 (N_10226,N_9780,N_6462);
and U10227 (N_10227,N_7521,N_5234);
xnor U10228 (N_10228,N_7618,N_7351);
nand U10229 (N_10229,N_9094,N_9884);
nand U10230 (N_10230,N_9092,N_8587);
and U10231 (N_10231,N_9555,N_9406);
and U10232 (N_10232,N_5433,N_8513);
and U10233 (N_10233,N_9715,N_8866);
and U10234 (N_10234,N_9942,N_6625);
nand U10235 (N_10235,N_9585,N_8561);
and U10236 (N_10236,N_5109,N_6330);
and U10237 (N_10237,N_9538,N_6695);
nor U10238 (N_10238,N_8879,N_6830);
nor U10239 (N_10239,N_6636,N_6634);
and U10240 (N_10240,N_6336,N_7396);
and U10241 (N_10241,N_9978,N_8654);
nor U10242 (N_10242,N_5664,N_6058);
xnor U10243 (N_10243,N_5589,N_7586);
and U10244 (N_10244,N_7528,N_6900);
nor U10245 (N_10245,N_5810,N_9830);
or U10246 (N_10246,N_9225,N_7730);
xor U10247 (N_10247,N_5797,N_6279);
nor U10248 (N_10248,N_9196,N_8055);
nand U10249 (N_10249,N_7696,N_6366);
or U10250 (N_10250,N_6170,N_5353);
nand U10251 (N_10251,N_9019,N_6396);
or U10252 (N_10252,N_8922,N_6569);
and U10253 (N_10253,N_6571,N_7552);
and U10254 (N_10254,N_8967,N_7953);
and U10255 (N_10255,N_8484,N_8888);
xor U10256 (N_10256,N_6843,N_8753);
or U10257 (N_10257,N_8539,N_5391);
nor U10258 (N_10258,N_5177,N_8785);
xnor U10259 (N_10259,N_5379,N_8357);
nor U10260 (N_10260,N_6039,N_5957);
or U10261 (N_10261,N_6960,N_6774);
nand U10262 (N_10262,N_8014,N_9084);
nand U10263 (N_10263,N_5842,N_8800);
xnor U10264 (N_10264,N_5645,N_9799);
nand U10265 (N_10265,N_6974,N_8398);
or U10266 (N_10266,N_7594,N_6815);
and U10267 (N_10267,N_9127,N_8564);
nor U10268 (N_10268,N_6347,N_7979);
and U10269 (N_10269,N_8680,N_6490);
nor U10270 (N_10270,N_8431,N_5420);
and U10271 (N_10271,N_8662,N_5014);
nand U10272 (N_10272,N_5357,N_6551);
or U10273 (N_10273,N_6342,N_7190);
xor U10274 (N_10274,N_6394,N_8805);
or U10275 (N_10275,N_9875,N_6624);
and U10276 (N_10276,N_8834,N_6586);
xor U10277 (N_10277,N_9211,N_9953);
and U10278 (N_10278,N_8083,N_6656);
nor U10279 (N_10279,N_7621,N_8051);
xor U10280 (N_10280,N_7284,N_7503);
or U10281 (N_10281,N_5317,N_5853);
and U10282 (N_10282,N_7860,N_9015);
and U10283 (N_10283,N_5451,N_7309);
xnor U10284 (N_10284,N_7753,N_8845);
and U10285 (N_10285,N_8091,N_5703);
nand U10286 (N_10286,N_6865,N_9335);
nand U10287 (N_10287,N_7041,N_6504);
xnor U10288 (N_10288,N_7087,N_5386);
nor U10289 (N_10289,N_7595,N_5337);
nor U10290 (N_10290,N_8331,N_9260);
nand U10291 (N_10291,N_6968,N_9857);
or U10292 (N_10292,N_7534,N_7466);
xnor U10293 (N_10293,N_8294,N_9500);
and U10294 (N_10294,N_5767,N_8685);
xor U10295 (N_10295,N_8797,N_5294);
and U10296 (N_10296,N_5593,N_9212);
nor U10297 (N_10297,N_6938,N_7875);
or U10298 (N_10298,N_8038,N_8017);
or U10299 (N_10299,N_7383,N_9673);
nor U10300 (N_10300,N_9098,N_6460);
and U10301 (N_10301,N_8337,N_9114);
xnor U10302 (N_10302,N_7592,N_7866);
and U10303 (N_10303,N_5632,N_8534);
nand U10304 (N_10304,N_8628,N_5023);
nor U10305 (N_10305,N_7963,N_6305);
xnor U10306 (N_10306,N_6710,N_9575);
xor U10307 (N_10307,N_6605,N_6792);
or U10308 (N_10308,N_8581,N_8386);
or U10309 (N_10309,N_8696,N_7990);
nand U10310 (N_10310,N_5159,N_6093);
nand U10311 (N_10311,N_5455,N_5405);
nor U10312 (N_10312,N_7718,N_7883);
xnor U10313 (N_10313,N_6519,N_5979);
or U10314 (N_10314,N_9058,N_9191);
or U10315 (N_10315,N_7290,N_6806);
nor U10316 (N_10316,N_7263,N_6686);
nand U10317 (N_10317,N_5730,N_5240);
or U10318 (N_10318,N_5295,N_7054);
nand U10319 (N_10319,N_6559,N_5575);
xnor U10320 (N_10320,N_9914,N_9949);
nor U10321 (N_10321,N_8498,N_9702);
xor U10322 (N_10322,N_5815,N_6466);
or U10323 (N_10323,N_6867,N_5149);
xnor U10324 (N_10324,N_7388,N_9769);
or U10325 (N_10325,N_9307,N_9615);
and U10326 (N_10326,N_5737,N_5640);
nand U10327 (N_10327,N_9992,N_6260);
or U10328 (N_10328,N_6687,N_6141);
nor U10329 (N_10329,N_8515,N_7110);
or U10330 (N_10330,N_5221,N_6228);
nor U10331 (N_10331,N_5187,N_6034);
nand U10332 (N_10332,N_9125,N_7413);
xor U10333 (N_10333,N_5275,N_8870);
xor U10334 (N_10334,N_6696,N_8546);
xnor U10335 (N_10335,N_6047,N_7359);
nor U10336 (N_10336,N_9694,N_5218);
xnor U10337 (N_10337,N_7365,N_5263);
and U10338 (N_10338,N_6679,N_7826);
nor U10339 (N_10339,N_8228,N_8312);
nand U10340 (N_10340,N_8891,N_9697);
or U10341 (N_10341,N_9327,N_5242);
nand U10342 (N_10342,N_5650,N_7293);
nor U10343 (N_10343,N_5096,N_7376);
xnor U10344 (N_10344,N_5231,N_6085);
xnor U10345 (N_10345,N_5838,N_5529);
xnor U10346 (N_10346,N_9091,N_5799);
nand U10347 (N_10347,N_8166,N_6767);
xnor U10348 (N_10348,N_7015,N_7930);
xnor U10349 (N_10349,N_7747,N_9440);
nor U10350 (N_10350,N_9782,N_9770);
or U10351 (N_10351,N_9726,N_6630);
and U10352 (N_10352,N_8626,N_9837);
xnor U10353 (N_10353,N_9297,N_6526);
nand U10354 (N_10354,N_6233,N_8315);
and U10355 (N_10355,N_5164,N_5659);
nand U10356 (N_10356,N_5333,N_5373);
and U10357 (N_10357,N_6138,N_5887);
nand U10358 (N_10358,N_9783,N_6837);
nand U10359 (N_10359,N_5506,N_8208);
nand U10360 (N_10360,N_6125,N_5443);
nor U10361 (N_10361,N_9804,N_5562);
nor U10362 (N_10362,N_5728,N_8303);
nor U10363 (N_10363,N_8350,N_8467);
xnor U10364 (N_10364,N_5549,N_9827);
nor U10365 (N_10365,N_9577,N_6339);
and U10366 (N_10366,N_5629,N_8807);
and U10367 (N_10367,N_5477,N_7635);
and U10368 (N_10368,N_6650,N_9810);
nand U10369 (N_10369,N_9743,N_9762);
xnor U10370 (N_10370,N_9367,N_5934);
and U10371 (N_10371,N_7439,N_9361);
nand U10372 (N_10372,N_9108,N_8491);
nor U10373 (N_10373,N_7308,N_9885);
nor U10374 (N_10374,N_5980,N_8934);
and U10375 (N_10375,N_8257,N_8748);
xnor U10376 (N_10376,N_5116,N_6614);
or U10377 (N_10377,N_9798,N_6870);
nand U10378 (N_10378,N_9331,N_7637);
nand U10379 (N_10379,N_6936,N_5396);
nand U10380 (N_10380,N_8732,N_9414);
xor U10381 (N_10381,N_9976,N_8137);
nor U10382 (N_10382,N_7301,N_6689);
nor U10383 (N_10383,N_7221,N_6632);
or U10384 (N_10384,N_5812,N_7241);
xnor U10385 (N_10385,N_5582,N_6845);
and U10386 (N_10386,N_7489,N_6970);
xnor U10387 (N_10387,N_8281,N_7395);
xnor U10388 (N_10388,N_9725,N_6405);
nor U10389 (N_10389,N_9687,N_6483);
and U10390 (N_10390,N_8230,N_7823);
and U10391 (N_10391,N_8479,N_9945);
nand U10392 (N_10392,N_7420,N_6829);
or U10393 (N_10393,N_5784,N_8410);
and U10394 (N_10394,N_8872,N_9564);
nor U10395 (N_10395,N_6933,N_6333);
xor U10396 (N_10396,N_8608,N_6131);
and U10397 (N_10397,N_7851,N_9213);
nor U10398 (N_10398,N_9828,N_7848);
xor U10399 (N_10399,N_5465,N_8478);
nor U10400 (N_10400,N_7660,N_6653);
nor U10401 (N_10401,N_9129,N_7833);
and U10402 (N_10402,N_6766,N_8961);
or U10403 (N_10403,N_7381,N_9111);
or U10404 (N_10404,N_5725,N_7176);
nand U10405 (N_10405,N_8013,N_8780);
nand U10406 (N_10406,N_5977,N_7088);
nand U10407 (N_10407,N_5877,N_6676);
nor U10408 (N_10408,N_6848,N_8985);
nor U10409 (N_10409,N_8368,N_9807);
nand U10410 (N_10410,N_9347,N_6242);
nor U10411 (N_10411,N_5794,N_8276);
nor U10412 (N_10412,N_8004,N_5264);
nor U10413 (N_10413,N_6544,N_9877);
xor U10414 (N_10414,N_5253,N_7387);
nor U10415 (N_10415,N_5963,N_7377);
nand U10416 (N_10416,N_7715,N_6668);
nand U10417 (N_10417,N_8118,N_6188);
nand U10418 (N_10418,N_9652,N_6167);
or U10419 (N_10419,N_5834,N_7115);
xnor U10420 (N_10420,N_5285,N_9690);
and U10421 (N_10421,N_9117,N_9434);
or U10422 (N_10422,N_9409,N_6240);
nor U10423 (N_10423,N_7273,N_9369);
xnor U10424 (N_10424,N_7039,N_6846);
or U10425 (N_10425,N_7226,N_5607);
nor U10426 (N_10426,N_5665,N_8438);
and U10427 (N_10427,N_8788,N_6646);
nand U10428 (N_10428,N_6040,N_6749);
or U10429 (N_10429,N_9647,N_7315);
nor U10430 (N_10430,N_6761,N_7220);
and U10431 (N_10431,N_5751,N_5960);
xnor U10432 (N_10432,N_8993,N_7434);
nand U10433 (N_10433,N_5898,N_5419);
xnor U10434 (N_10434,N_9540,N_7961);
nand U10435 (N_10435,N_8656,N_7331);
nand U10436 (N_10436,N_5272,N_5094);
nor U10437 (N_10437,N_5950,N_7871);
nand U10438 (N_10438,N_6165,N_5907);
and U10439 (N_10439,N_5474,N_6939);
nor U10440 (N_10440,N_8799,N_6771);
nor U10441 (N_10441,N_5246,N_9207);
nor U10442 (N_10442,N_7513,N_6631);
nor U10443 (N_10443,N_5587,N_9141);
nor U10444 (N_10444,N_8862,N_8566);
nor U10445 (N_10445,N_7683,N_5306);
or U10446 (N_10446,N_9423,N_9421);
nand U10447 (N_10447,N_6873,N_5761);
xnor U10448 (N_10448,N_7457,N_6524);
nor U10449 (N_10449,N_5889,N_5636);
xor U10450 (N_10450,N_9583,N_8182);
xor U10451 (N_10451,N_8894,N_7770);
or U10452 (N_10452,N_9871,N_5573);
nand U10453 (N_10453,N_5505,N_7225);
or U10454 (N_10454,N_8428,N_7729);
nand U10455 (N_10455,N_7865,N_5298);
nor U10456 (N_10456,N_7974,N_5905);
nor U10457 (N_10457,N_6618,N_9849);
and U10458 (N_10458,N_6130,N_7634);
and U10459 (N_10459,N_6080,N_9961);
nor U10460 (N_10460,N_5392,N_6753);
nor U10461 (N_10461,N_8184,N_9512);
xor U10462 (N_10462,N_6604,N_6282);
nor U10463 (N_10463,N_5808,N_7400);
xor U10464 (N_10464,N_5623,N_7844);
nor U10465 (N_10465,N_8126,N_6346);
nor U10466 (N_10466,N_6082,N_7831);
nor U10467 (N_10467,N_5249,N_7412);
nand U10468 (N_10468,N_7408,N_6916);
nand U10469 (N_10469,N_8859,N_6478);
nor U10470 (N_10470,N_7765,N_8183);
xnor U10471 (N_10471,N_6716,N_6357);
nor U10472 (N_10472,N_9029,N_8878);
and U10473 (N_10473,N_8824,N_6171);
nand U10474 (N_10474,N_7658,N_5781);
xor U10475 (N_10475,N_8000,N_5043);
nor U10476 (N_10476,N_8105,N_6276);
nor U10477 (N_10477,N_9870,N_9539);
xor U10478 (N_10478,N_7855,N_7082);
and U10479 (N_10479,N_6861,N_8069);
or U10480 (N_10480,N_7535,N_5522);
and U10481 (N_10481,N_8122,N_5829);
or U10482 (N_10482,N_6248,N_6390);
nor U10483 (N_10483,N_7196,N_7788);
xor U10484 (N_10484,N_7491,N_8452);
and U10485 (N_10485,N_6541,N_5528);
or U10486 (N_10486,N_9080,N_9918);
and U10487 (N_10487,N_6596,N_6161);
nor U10488 (N_10488,N_6701,N_7962);
xor U10489 (N_10489,N_8147,N_7549);
nand U10490 (N_10490,N_5435,N_5492);
or U10491 (N_10491,N_8128,N_5687);
nor U10492 (N_10492,N_5865,N_9036);
or U10493 (N_10493,N_5598,N_9195);
or U10494 (N_10494,N_6144,N_9462);
or U10495 (N_10495,N_7472,N_5509);
or U10496 (N_10496,N_6959,N_7709);
nand U10497 (N_10497,N_6527,N_8772);
nor U10498 (N_10498,N_6077,N_9505);
or U10499 (N_10499,N_5712,N_9284);
nor U10500 (N_10500,N_5224,N_9850);
xnor U10501 (N_10501,N_8992,N_7274);
and U10502 (N_10502,N_8274,N_6151);
nand U10503 (N_10503,N_9206,N_7428);
or U10504 (N_10504,N_6122,N_6071);
or U10505 (N_10505,N_9456,N_9373);
or U10506 (N_10506,N_5388,N_5987);
xnor U10507 (N_10507,N_8745,N_5178);
or U10508 (N_10508,N_9394,N_8348);
xor U10509 (N_10509,N_7276,N_8497);
xnor U10510 (N_10510,N_5350,N_6379);
nor U10511 (N_10511,N_6708,N_7209);
and U10512 (N_10512,N_9452,N_5365);
or U10513 (N_10513,N_9236,N_6391);
nor U10514 (N_10514,N_7629,N_6418);
or U10515 (N_10515,N_9424,N_9378);
or U10516 (N_10516,N_9076,N_6784);
nor U10517 (N_10517,N_7450,N_7379);
nor U10518 (N_10518,N_7847,N_8382);
or U10519 (N_10519,N_9140,N_8849);
and U10520 (N_10520,N_6354,N_6358);
and U10521 (N_10521,N_7545,N_8336);
nand U10522 (N_10522,N_8375,N_5214);
nand U10523 (N_10523,N_9483,N_9278);
nor U10524 (N_10524,N_6110,N_7666);
or U10525 (N_10525,N_8749,N_9562);
and U10526 (N_10526,N_8044,N_5276);
and U10527 (N_10527,N_9180,N_6557);
nor U10528 (N_10528,N_7697,N_6380);
xor U10529 (N_10529,N_8133,N_5855);
nand U10530 (N_10530,N_7010,N_8098);
nor U10531 (N_10531,N_6152,N_7136);
nand U10532 (N_10532,N_6363,N_6776);
and U10533 (N_10533,N_5923,N_8535);
nor U10534 (N_10534,N_7498,N_6738);
nor U10535 (N_10535,N_5984,N_8271);
nor U10536 (N_10536,N_7159,N_5148);
nand U10537 (N_10537,N_9644,N_8846);
or U10538 (N_10538,N_7127,N_8630);
nand U10539 (N_10539,N_9853,N_5732);
xor U10540 (N_10540,N_5945,N_6016);
and U10541 (N_10541,N_8236,N_7470);
xor U10542 (N_10542,N_7462,N_8511);
or U10543 (N_10543,N_9205,N_6163);
nor U10544 (N_10544,N_7563,N_8358);
or U10545 (N_10545,N_7492,N_6640);
xnor U10546 (N_10546,N_6620,N_6978);
and U10547 (N_10547,N_9197,N_5634);
xnor U10548 (N_10548,N_6496,N_5740);
or U10549 (N_10549,N_8311,N_5667);
nor U10550 (N_10550,N_5867,N_8117);
xor U10551 (N_10551,N_6089,N_6560);
nor U10552 (N_10552,N_9492,N_5271);
xor U10553 (N_10553,N_6733,N_8826);
and U10554 (N_10554,N_8423,N_6879);
or U10555 (N_10555,N_8598,N_8882);
and U10556 (N_10556,N_5939,N_7548);
nand U10557 (N_10557,N_7426,N_6849);
nor U10558 (N_10558,N_5427,N_9648);
and U10559 (N_10559,N_6585,N_7421);
nor U10560 (N_10560,N_7150,N_5777);
nand U10561 (N_10561,N_9131,N_6772);
and U10562 (N_10562,N_5322,N_5301);
nand U10563 (N_10563,N_7070,N_8939);
nand U10564 (N_10564,N_5863,N_7924);
or U10565 (N_10565,N_9262,N_7938);
nor U10566 (N_10566,N_8646,N_8219);
or U10567 (N_10567,N_5220,N_9045);
or U10568 (N_10568,N_9461,N_7517);
and U10569 (N_10569,N_6497,N_8975);
or U10570 (N_10570,N_8189,N_6353);
xnor U10571 (N_10571,N_9716,N_8545);
nor U10572 (N_10572,N_8617,N_6914);
nand U10573 (N_10573,N_9217,N_9023);
and U10574 (N_10574,N_7514,N_7917);
nand U10575 (N_10575,N_6222,N_7725);
and U10576 (N_10576,N_6893,N_8376);
nand U10577 (N_10577,N_8130,N_5377);
or U10578 (N_10578,N_6730,N_6146);
or U10579 (N_10579,N_5434,N_7405);
nand U10580 (N_10580,N_7074,N_5719);
or U10581 (N_10581,N_6112,N_5424);
nor U10582 (N_10582,N_5660,N_8064);
and U10583 (N_10583,N_7890,N_9490);
nor U10584 (N_10584,N_5336,N_8868);
and U10585 (N_10585,N_5284,N_6740);
xor U10586 (N_10586,N_7072,N_6115);
or U10587 (N_10587,N_8252,N_5207);
nor U10588 (N_10588,N_6424,N_7524);
nor U10589 (N_10589,N_9228,N_5611);
xor U10590 (N_10590,N_8195,N_9037);
or U10591 (N_10591,N_7928,N_7460);
xor U10592 (N_10592,N_6857,N_8093);
or U10593 (N_10593,N_6207,N_7766);
or U10594 (N_10594,N_6195,N_8193);
nand U10595 (N_10595,N_7551,N_9866);
and U10596 (N_10596,N_5439,N_9637);
xnor U10597 (N_10597,N_9855,N_5666);
xor U10598 (N_10598,N_8629,N_9679);
or U10599 (N_10599,N_8170,N_9760);
nor U10600 (N_10600,N_8927,N_6403);
xnor U10601 (N_10601,N_5282,N_8495);
nor U10602 (N_10602,N_8255,N_9230);
xnor U10603 (N_10603,N_7945,N_8871);
or U10604 (N_10604,N_9386,N_6518);
or U10605 (N_10605,N_8068,N_6877);
or U10606 (N_10606,N_9887,N_9333);
xnor U10607 (N_10607,N_8355,N_7090);
nand U10608 (N_10608,N_9243,N_7314);
nor U10609 (N_10609,N_9283,N_9764);
xor U10610 (N_10610,N_6495,N_5027);
nor U10611 (N_10611,N_5466,N_6286);
nor U10612 (N_10612,N_5193,N_6392);
and U10613 (N_10613,N_9006,N_7044);
and U10614 (N_10614,N_6608,N_7880);
xor U10615 (N_10615,N_8178,N_5683);
and U10616 (N_10616,N_6012,N_9814);
or U10617 (N_10617,N_9061,N_5491);
xnor U10618 (N_10618,N_8510,N_8461);
nor U10619 (N_10619,N_7556,N_9404);
nor U10620 (N_10620,N_8643,N_5827);
or U10621 (N_10621,N_8504,N_8026);
or U10622 (N_10622,N_5293,N_5947);
or U10623 (N_10623,N_9581,N_9407);
or U10624 (N_10624,N_5568,N_8299);
xor U10625 (N_10625,N_5467,N_8464);
or U10626 (N_10626,N_7936,N_6119);
nor U10627 (N_10627,N_8508,N_7763);
and U10628 (N_10628,N_6364,N_6432);
xnor U10629 (N_10629,N_7337,N_9498);
or U10630 (N_10630,N_7278,N_7566);
and U10631 (N_10631,N_9565,N_8270);
nand U10632 (N_10632,N_7558,N_5063);
xnor U10633 (N_10633,N_7192,N_5179);
nand U10634 (N_10634,N_5901,N_5891);
nor U10635 (N_10635,N_6200,N_7432);
and U10636 (N_10636,N_6734,N_5937);
or U10637 (N_10637,N_5086,N_7812);
nand U10638 (N_10638,N_6909,N_7589);
xor U10639 (N_10639,N_8447,N_8613);
xor U10640 (N_10640,N_6120,N_8424);
or U10641 (N_10641,N_6796,N_5126);
nor U10642 (N_10642,N_6777,N_5291);
nand U10643 (N_10643,N_9517,N_6573);
and U10644 (N_10644,N_8214,N_8033);
nand U10645 (N_10645,N_9720,N_7982);
and U10646 (N_10646,N_9719,N_7320);
and U10647 (N_10647,N_9792,N_7896);
or U10648 (N_10648,N_7895,N_5217);
nand U10649 (N_10649,N_7893,N_8154);
nand U10650 (N_10650,N_5690,N_7892);
nand U10651 (N_10651,N_7649,N_6735);
nand U10652 (N_10652,N_7223,N_9560);
xnor U10653 (N_10653,N_7235,N_9504);
nand U10654 (N_10654,N_8997,N_8190);
nand U10655 (N_10655,N_8387,N_7158);
xor U10656 (N_10656,N_7113,N_5644);
xnor U10657 (N_10657,N_6054,N_8021);
and U10658 (N_10658,N_5552,N_8651);
nor U10659 (N_10659,N_9551,N_9595);
and U10660 (N_10660,N_9677,N_8635);
nor U10661 (N_10661,N_7732,N_9536);
xnor U10662 (N_10662,N_9304,N_6564);
or U10663 (N_10663,N_8283,N_5406);
nand U10664 (N_10664,N_8077,N_6344);
and U10665 (N_10665,N_5299,N_7782);
nor U10666 (N_10666,N_6199,N_9496);
nand U10667 (N_10667,N_6425,N_7008);
and U10668 (N_10668,N_8286,N_6554);
and U10669 (N_10669,N_6958,N_7824);
or U10670 (N_10670,N_8619,N_7940);
or U10671 (N_10671,N_7675,N_5073);
or U10672 (N_10672,N_5503,N_9802);
nand U10673 (N_10673,N_5118,N_8703);
and U10674 (N_10674,N_8092,N_5779);
nand U10675 (N_10675,N_6459,N_5128);
or U10676 (N_10676,N_7475,N_5321);
xnor U10677 (N_10677,N_7347,N_8110);
or U10678 (N_10678,N_8463,N_6831);
xor U10679 (N_10679,N_9357,N_9489);
xnor U10680 (N_10680,N_5711,N_6453);
and U10681 (N_10681,N_9878,N_6997);
or U10682 (N_10682,N_8482,N_6011);
nand U10683 (N_10683,N_9839,N_9649);
xor U10684 (N_10684,N_9224,N_5079);
and U10685 (N_10685,N_5141,N_7474);
xnor U10686 (N_10686,N_6192,N_6320);
xor U10687 (N_10687,N_7531,N_6705);
nand U10688 (N_10688,N_6428,N_8318);
nand U10689 (N_10689,N_9215,N_6779);
xor U10690 (N_10690,N_6386,N_9401);
xnor U10691 (N_10691,N_7809,N_5657);
and U10692 (N_10692,N_7375,N_6301);
nand U10693 (N_10693,N_6862,N_6964);
nand U10694 (N_10694,N_6057,N_9494);
nor U10695 (N_10695,N_7303,N_8359);
nand U10696 (N_10696,N_5054,N_8298);
nor U10697 (N_10697,N_6155,N_6757);
nand U10698 (N_10698,N_5615,N_5841);
nand U10699 (N_10699,N_7084,N_7903);
nor U10700 (N_10700,N_7850,N_9171);
nor U10701 (N_10701,N_6489,N_5935);
or U10702 (N_10702,N_7601,N_5348);
nor U10703 (N_10703,N_6420,N_5830);
or U10704 (N_10704,N_5897,N_5449);
and U10705 (N_10705,N_6990,N_5592);
and U10706 (N_10706,N_9138,N_5597);
xor U10707 (N_10707,N_7338,N_7562);
nand U10708 (N_10708,N_6886,N_6591);
nor U10709 (N_10709,N_6566,N_5328);
nand U10710 (N_10710,N_6723,N_7112);
nand U10711 (N_10711,N_6533,N_8400);
and U10712 (N_10712,N_5541,N_8324);
and U10713 (N_10713,N_7523,N_5145);
or U10714 (N_10714,N_9450,N_9738);
xnor U10715 (N_10715,N_8591,N_7210);
xnor U10716 (N_10716,N_9987,N_5012);
and U10717 (N_10717,N_9477,N_8320);
and U10718 (N_10718,N_6555,N_9022);
or U10719 (N_10719,N_5988,N_7096);
and U10720 (N_10720,N_5642,N_5953);
xnor U10721 (N_10721,N_8015,N_7861);
nand U10722 (N_10722,N_5289,N_8946);
and U10723 (N_10723,N_8307,N_7567);
xnor U10724 (N_10724,N_9891,N_6957);
or U10725 (N_10725,N_7778,N_6456);
and U10726 (N_10726,N_8361,N_5196);
nand U10727 (N_10727,N_6029,N_5507);
and U10728 (N_10728,N_6603,N_7508);
xor U10729 (N_10729,N_5899,N_7997);
and U10730 (N_10730,N_5762,N_9273);
and U10731 (N_10731,N_9251,N_7958);
or U10732 (N_10732,N_5699,N_8101);
xor U10733 (N_10733,N_5501,N_6097);
and U10734 (N_10734,N_5325,N_6924);
or U10735 (N_10735,N_9342,N_7700);
xor U10736 (N_10736,N_5532,N_5423);
nor U10737 (N_10737,N_6156,N_8659);
xor U10738 (N_10738,N_6209,N_7336);
nand U10739 (N_10739,N_8364,N_8906);
xor U10740 (N_10740,N_7780,N_9267);
or U10741 (N_10741,N_8549,N_6577);
nand U10742 (N_10742,N_8186,N_6575);
nor U10743 (N_10743,N_9183,N_9958);
and U10744 (N_10744,N_6259,N_5274);
nor U10745 (N_10745,N_6317,N_6635);
nor U10746 (N_10746,N_7485,N_9748);
xnor U10747 (N_10747,N_7057,N_6765);
xor U10748 (N_10748,N_7733,N_6580);
nor U10749 (N_10749,N_7346,N_9385);
nand U10750 (N_10750,N_9750,N_6712);
or U10751 (N_10751,N_6561,N_5344);
nand U10752 (N_10752,N_8202,N_5744);
xnor U10753 (N_10753,N_8127,N_9400);
nand U10754 (N_10754,N_7031,N_5084);
nor U10755 (N_10755,N_5964,N_6866);
nor U10756 (N_10756,N_9009,N_8568);
and U10757 (N_10757,N_8848,N_5205);
xnor U10758 (N_10758,N_9097,N_8966);
nand U10759 (N_10759,N_5788,N_6697);
nand U10760 (N_10760,N_9838,N_8829);
or U10761 (N_10761,N_8469,N_7720);
and U10762 (N_10762,N_7630,N_5551);
and U10763 (N_10763,N_9145,N_6664);
nand U10764 (N_10764,N_9218,N_8751);
or U10765 (N_10765,N_7570,N_8770);
nand U10766 (N_10766,N_9046,N_7108);
nand U10767 (N_10767,N_5354,N_6521);
and U10768 (N_10768,N_9063,N_9344);
xor U10769 (N_10769,N_9296,N_8565);
and U10770 (N_10770,N_6853,N_6351);
nor U10771 (N_10771,N_6205,N_8239);
and U10772 (N_10772,N_6307,N_6100);
and U10773 (N_10773,N_5502,N_5300);
and U10774 (N_10774,N_6487,N_7258);
and U10775 (N_10775,N_6078,N_6329);
nor U10776 (N_10776,N_5120,N_9634);
or U10777 (N_10777,N_8207,N_9622);
or U10778 (N_10778,N_6331,N_6442);
or U10779 (N_10779,N_5544,N_6001);
nand U10780 (N_10780,N_9654,N_6246);
xnor U10781 (N_10781,N_7538,N_7946);
nand U10782 (N_10782,N_8991,N_8003);
and U10783 (N_10783,N_7191,N_5917);
and U10784 (N_10784,N_8343,N_6124);
nor U10785 (N_10785,N_6467,N_8450);
nand U10786 (N_10786,N_8076,N_6007);
or U10787 (N_10787,N_9453,N_8246);
xnor U10788 (N_10788,N_5339,N_8664);
nor U10789 (N_10789,N_9617,N_7699);
xnor U10790 (N_10790,N_5983,N_6072);
nand U10791 (N_10791,N_8002,N_7511);
or U10792 (N_10792,N_6828,N_6578);
and U10793 (N_10793,N_5792,N_9561);
xnor U10794 (N_10794,N_7109,N_8911);
nand U10795 (N_10795,N_9620,N_7884);
nand U10796 (N_10796,N_7547,N_9940);
nand U10797 (N_10797,N_9641,N_9744);
nor U10798 (N_10798,N_7198,N_5102);
or U10799 (N_10799,N_9775,N_9594);
nand U10800 (N_10800,N_6203,N_8245);
nor U10801 (N_10801,N_5869,N_9027);
and U10802 (N_10802,N_6241,N_9011);
nor U10803 (N_10803,N_7423,N_5858);
nor U10804 (N_10804,N_7271,N_7366);
xnor U10805 (N_10805,N_9806,N_9085);
or U10806 (N_10806,N_8761,N_9675);
and U10807 (N_10807,N_7550,N_7130);
nand U10808 (N_10808,N_8365,N_9426);
and U10809 (N_10809,N_7171,N_6374);
and U10810 (N_10810,N_7792,N_6056);
and U10811 (N_10811,N_8860,N_7013);
or U10812 (N_10812,N_8550,N_5213);
nor U10813 (N_10813,N_8516,N_6299);
or U10814 (N_10814,N_5966,N_6858);
or U10815 (N_10815,N_9057,N_5106);
or U10816 (N_10816,N_5882,N_7616);
nand U10817 (N_10817,N_7886,N_9977);
nand U10818 (N_10818,N_8612,N_9852);
nand U10819 (N_10819,N_7583,N_6023);
nor U10820 (N_10820,N_7891,N_8174);
xnor U10821 (N_10821,N_9547,N_7795);
nand U10822 (N_10822,N_6659,N_6254);
and U10823 (N_10823,N_9952,N_5490);
xnor U10824 (N_10824,N_9305,N_6639);
or U10825 (N_10825,N_9030,N_5082);
or U10826 (N_10826,N_5031,N_9122);
nand U10827 (N_10827,N_6435,N_9737);
nor U10828 (N_10828,N_5733,N_7682);
nor U10829 (N_10829,N_5080,N_8140);
or U10830 (N_10830,N_6316,N_8676);
xor U10831 (N_10831,N_6891,N_5119);
or U10832 (N_10832,N_7238,N_9427);
nand U10833 (N_10833,N_6863,N_6898);
and U10834 (N_10834,N_5545,N_9148);
nor U10835 (N_10835,N_6895,N_7026);
nand U10836 (N_10836,N_6096,N_9755);
and U10837 (N_10837,N_7053,N_9154);
nand U10838 (N_10838,N_9931,N_9486);
and U10839 (N_10839,N_9392,N_7449);
and U10840 (N_10840,N_5619,N_6607);
xor U10841 (N_10841,N_8638,N_5058);
and U10842 (N_10842,N_9842,N_6253);
and U10843 (N_10843,N_8525,N_9182);
or U10844 (N_10844,N_9113,N_6257);
nor U10845 (N_10845,N_8085,N_7758);
and U10846 (N_10846,N_8037,N_8198);
nor U10847 (N_10847,N_7302,N_8825);
or U10848 (N_10848,N_8977,N_9431);
or U10849 (N_10849,N_7702,N_5314);
and U10850 (N_10850,N_9383,N_7495);
xnor U10851 (N_10851,N_7748,N_9797);
xor U10852 (N_10852,N_7264,N_5546);
nand U10853 (N_10853,N_8896,N_7864);
nor U10854 (N_10854,N_5601,N_5398);
nor U10855 (N_10855,N_8577,N_6798);
or U10856 (N_10856,N_9189,N_7948);
nor U10857 (N_10857,N_6514,N_5919);
or U10858 (N_10858,N_7035,N_5695);
xor U10859 (N_10859,N_7204,N_9418);
nor U10860 (N_10860,N_8713,N_6113);
nor U10861 (N_10861,N_5843,N_6327);
xnor U10862 (N_10862,N_7964,N_6989);
or U10863 (N_10863,N_8151,N_7994);
and U10864 (N_10864,N_8048,N_5399);
nand U10865 (N_10865,N_8789,N_7114);
nand U10866 (N_10866,N_5559,N_9682);
nor U10867 (N_10867,N_9355,N_9299);
and U10868 (N_10868,N_6121,N_8066);
nor U10869 (N_10869,N_8957,N_6186);
nor U10870 (N_10870,N_9508,N_6780);
and U10871 (N_10871,N_5239,N_6311);
xnor U10872 (N_10872,N_9341,N_8448);
nand U10873 (N_10873,N_6822,N_6896);
or U10874 (N_10874,N_7398,N_5108);
and U10875 (N_10875,N_7842,N_6008);
or U10876 (N_10876,N_9676,N_7764);
nand U10877 (N_10877,N_8010,N_5250);
and U10878 (N_10878,N_5154,N_8142);
nor U10879 (N_10879,N_6940,N_5753);
and U10880 (N_10880,N_6463,N_7019);
nor U10881 (N_10881,N_6988,N_6053);
nand U10882 (N_10882,N_5876,N_9372);
and U10883 (N_10883,N_8277,N_8747);
and U10884 (N_10884,N_5688,N_9413);
nand U10885 (N_10885,N_9238,N_9158);
nand U10886 (N_10886,N_9429,N_7540);
nand U10887 (N_10887,N_8280,N_9834);
and U10888 (N_10888,N_7006,N_5723);
or U10889 (N_10889,N_6304,N_7468);
nor U10890 (N_10890,N_7712,N_5975);
xor U10891 (N_10891,N_9692,N_5770);
and U10892 (N_10892,N_5375,N_8150);
nor U10893 (N_10893,N_6674,N_6944);
xnor U10894 (N_10894,N_9822,N_9055);
and U10895 (N_10895,N_8572,N_8421);
nor U10896 (N_10896,N_5197,N_7069);
or U10897 (N_10897,N_6382,N_9811);
xnor U10898 (N_10898,N_9607,N_8858);
and U10899 (N_10899,N_6433,N_5859);
and U10900 (N_10900,N_9533,N_7327);
or U10901 (N_10901,N_6615,N_8919);
xnor U10902 (N_10902,N_7968,N_6963);
and U10903 (N_10903,N_9889,N_6643);
or U10904 (N_10904,N_6212,N_7497);
nand U10905 (N_10905,N_7722,N_8310);
nand U10906 (N_10906,N_5976,N_8035);
xor U10907 (N_10907,N_8253,N_5369);
xor U10908 (N_10908,N_5081,N_7754);
xnor U10909 (N_10909,N_5872,N_7541);
nand U10910 (N_10910,N_8486,N_9495);
and U10911 (N_10911,N_5039,N_7232);
and U10912 (N_10912,N_6025,N_8673);
nor U10913 (N_10913,N_6515,N_6803);
nand U10914 (N_10914,N_7603,N_8007);
or U10915 (N_10915,N_7659,N_6894);
nor U10916 (N_10916,N_5338,N_6722);
nand U10917 (N_10917,N_8422,N_9796);
or U10918 (N_10918,N_6621,N_5183);
or U10919 (N_10919,N_9146,N_7281);
nand U10920 (N_10920,N_9364,N_7775);
nand U10921 (N_10921,N_8124,N_7561);
xnor U10922 (N_10922,N_7085,N_6788);
nand U10923 (N_10923,N_6584,N_8153);
nand U10924 (N_10924,N_7655,N_9669);
or U10925 (N_10925,N_6869,N_5618);
and U10926 (N_10926,N_8773,N_8687);
and U10927 (N_10927,N_6292,N_6159);
and U10928 (N_10928,N_5483,N_6694);
and U10929 (N_10929,N_7676,N_5576);
nand U10930 (N_10930,N_8940,N_7544);
xnor U10931 (N_10931,N_5789,N_8792);
xor U10932 (N_10932,N_8333,N_8102);
xnor U10933 (N_10933,N_8081,N_8784);
nand U10934 (N_10934,N_6491,N_9991);
nor U10935 (N_10935,N_5168,N_7689);
xor U10936 (N_10936,N_6503,N_6622);
xor U10937 (N_10937,N_9816,N_9231);
nor U10938 (N_10938,N_7987,N_6685);
nor U10939 (N_10939,N_9204,N_9397);
xnor U10940 (N_10940,N_9475,N_7118);
and U10941 (N_10941,N_7148,N_5315);
nor U10942 (N_10942,N_8199,N_8765);
and U10943 (N_10943,N_8544,N_9823);
xnor U10944 (N_10944,N_6473,N_8810);
or U10945 (N_10945,N_5083,N_7404);
nand U10946 (N_10946,N_7146,N_5381);
or U10947 (N_10947,N_6230,N_9576);
and U10948 (N_10948,N_8976,N_8481);
or U10949 (N_10949,N_8454,N_9473);
and U10950 (N_10950,N_8721,N_8313);
xnor U10951 (N_10951,N_5087,N_5512);
or U10952 (N_10952,N_9039,N_9149);
or U10953 (N_10953,N_7218,N_8268);
xor U10954 (N_10954,N_5482,N_9044);
nor U10955 (N_10955,N_7165,N_6811);
nand U10956 (N_10956,N_9102,N_9626);
nand U10957 (N_10957,N_6231,N_9081);
or U10958 (N_10958,N_9951,N_7431);
or U10959 (N_10959,N_6312,N_5878);
nor U10960 (N_10960,N_7095,N_7125);
and U10961 (N_10961,N_9526,N_8289);
or U10962 (N_10962,N_7215,N_5716);
nand U10963 (N_10963,N_6162,N_9350);
xor U10964 (N_10964,N_6638,N_8576);
or U10965 (N_10965,N_6375,N_8661);
nand U10966 (N_10966,N_7698,N_7688);
nor U10967 (N_10967,N_7815,N_6663);
and U10968 (N_10968,N_9786,N_5216);
nand U10969 (N_10969,N_7007,N_9014);
nand U10970 (N_10970,N_5190,N_7607);
nor U10971 (N_10971,N_7926,N_5252);
or U10972 (N_10972,N_6367,N_8714);
xor U10973 (N_10973,N_6800,N_7482);
and U10974 (N_10974,N_9147,N_8913);
or U10975 (N_10975,N_9201,N_9747);
and U10976 (N_10976,N_9713,N_6549);
xor U10977 (N_10977,N_9598,N_8701);
and U10978 (N_10978,N_7254,N_6899);
nor U10979 (N_10979,N_9548,N_5968);
nand U10980 (N_10980,N_5103,N_9727);
or U10981 (N_10981,N_7755,N_7802);
xor U10982 (N_10982,N_8406,N_7129);
or U10983 (N_10983,N_8455,N_5750);
xnor U10984 (N_10984,N_7836,N_9537);
and U10985 (N_10985,N_9178,N_5461);
nor U10986 (N_10986,N_5803,N_7522);
or U10987 (N_10987,N_8889,N_5857);
and U10988 (N_10988,N_7187,N_6913);
or U10989 (N_10989,N_8413,N_7919);
nand U10990 (N_10990,N_6360,N_8791);
or U10991 (N_10991,N_7704,N_8039);
and U10992 (N_10992,N_5906,N_6808);
and U10993 (N_10993,N_8540,N_9860);
and U10994 (N_10994,N_7048,N_9497);
xor U10995 (N_10995,N_9938,N_6637);
nor U10996 (N_10996,N_7811,N_8215);
nand U10997 (N_10997,N_9087,N_9232);
nand U10998 (N_10998,N_8100,N_8296);
nor U10999 (N_10999,N_6923,N_9443);
nand U11000 (N_11000,N_6658,N_5140);
nor U11001 (N_11001,N_5124,N_6856);
xor U11002 (N_11002,N_7343,N_5211);
xor U11003 (N_11003,N_9192,N_6833);
or U11004 (N_11004,N_5204,N_5101);
xor U11005 (N_11005,N_5170,N_6216);
or U11006 (N_11006,N_5192,N_7203);
or U11007 (N_11007,N_6154,N_6878);
nor U11008 (N_11008,N_5965,N_7706);
xnor U11009 (N_11009,N_9599,N_7862);
or U11010 (N_11010,N_7230,N_5358);
xor U11011 (N_11011,N_7988,N_5773);
and U11012 (N_11012,N_6492,N_9152);
and U11013 (N_11013,N_6092,N_7931);
nor U11014 (N_11014,N_9610,N_8665);
or U11015 (N_11015,N_6015,N_7923);
xnor U11016 (N_11016,N_7325,N_5521);
nand U11017 (N_11017,N_8631,N_7798);
xor U11018 (N_11018,N_8019,N_5580);
and U11019 (N_11019,N_5436,N_5854);
nor U11020 (N_11020,N_5717,N_8370);
and U11021 (N_11021,N_9927,N_8347);
nor U11022 (N_11022,N_7835,N_8340);
or U11023 (N_11023,N_6535,N_9074);
nor U11024 (N_11024,N_5561,N_7416);
nor U11025 (N_11025,N_5729,N_9714);
xnor U11026 (N_11026,N_8802,N_6290);
or U11027 (N_11027,N_8593,N_9264);
nand U11028 (N_11028,N_6683,N_6046);
or U11029 (N_11029,N_8057,N_5836);
nor U11030 (N_11030,N_9454,N_9545);
and U11031 (N_11031,N_8657,N_8970);
and U11032 (N_11032,N_9374,N_6288);
and U11033 (N_11033,N_6925,N_9471);
or U11034 (N_11034,N_5421,N_5722);
or U11035 (N_11035,N_6417,N_8353);
nor U11036 (N_11036,N_7389,N_5481);
and U11037 (N_11037,N_8712,N_6847);
xnor U11038 (N_11038,N_7623,N_7568);
nor U11039 (N_11039,N_7927,N_6543);
xnor U11040 (N_11040,N_8728,N_9833);
or U11041 (N_11041,N_6983,N_6373);
nand U11042 (N_11042,N_6651,N_9103);
nor U11043 (N_11043,N_6550,N_6035);
xnor U11044 (N_11044,N_5452,N_5595);
nor U11045 (N_11045,N_9926,N_9709);
nand U11046 (N_11046,N_7356,N_8950);
and U11047 (N_11047,N_9176,N_9815);
or U11048 (N_11048,N_8405,N_5591);
xnor U11049 (N_11049,N_6885,N_5001);
nand U11050 (N_11050,N_5009,N_7023);
or U11051 (N_11051,N_8229,N_6376);
nor U11052 (N_11052,N_7403,N_7142);
and U11053 (N_11053,N_9908,N_6568);
xnor U11054 (N_11054,N_7691,N_9066);
and U11055 (N_11055,N_8399,N_8941);
or U11056 (N_11056,N_7488,N_9001);
nor U11057 (N_11057,N_5462,N_8050);
or U11058 (N_11058,N_7879,N_9915);
or U11059 (N_11059,N_5990,N_6754);
xor U11060 (N_11060,N_9247,N_6204);
and U11061 (N_11061,N_8874,N_6187);
nand U11062 (N_11062,N_5662,N_5428);
nor U11063 (N_11063,N_6529,N_5048);
or U11064 (N_11064,N_6702,N_8823);
nand U11065 (N_11065,N_5132,N_7024);
and U11066 (N_11066,N_7469,N_6183);
nor U11067 (N_11067,N_7373,N_7713);
nor U11068 (N_11068,N_6179,N_6499);
and U11069 (N_11069,N_6556,N_7350);
nor U11070 (N_11070,N_6642,N_9986);
nor U11071 (N_11071,N_5776,N_5131);
nand U11072 (N_11072,N_8744,N_7353);
or U11073 (N_11073,N_5793,N_9116);
xnor U11074 (N_11074,N_6810,N_6718);
xnor U11075 (N_11075,N_9356,N_5663);
xor U11076 (N_11076,N_7126,N_9618);
nand U11077 (N_11077,N_7796,N_7995);
or U11078 (N_11078,N_8404,N_6817);
nand U11079 (N_11079,N_8813,N_9998);
nand U11080 (N_11080,N_8944,N_5563);
nor U11081 (N_11081,N_8875,N_5948);
and U11082 (N_11082,N_7504,N_9288);
and U11083 (N_11083,N_9089,N_7391);
xor U11084 (N_11084,N_7662,N_7018);
and U11085 (N_11085,N_6839,N_8272);
nand U11086 (N_11086,N_7296,N_5127);
or U11087 (N_11087,N_9522,N_5497);
nor U11088 (N_11088,N_6273,N_8904);
xor U11089 (N_11089,N_8485,N_7231);
or U11090 (N_11090,N_5888,N_9405);
or U11091 (N_11091,N_8192,N_7843);
nand U11092 (N_11092,N_8588,N_7304);
xor U11093 (N_11093,N_7525,N_7425);
or U11094 (N_11094,N_8445,N_6942);
nand U11095 (N_11095,N_7339,N_5280);
or U11096 (N_11096,N_7587,N_6824);
or U11097 (N_11097,N_8067,N_6812);
xor U11098 (N_11098,N_7249,N_9003);
nor U11099 (N_11099,N_6217,N_9847);
xor U11100 (N_11100,N_8243,N_8062);
xnor U11101 (N_11101,N_8200,N_8996);
xnor U11102 (N_11102,N_8158,N_5714);
nand U11103 (N_11103,N_9198,N_8327);
nor U11104 (N_11104,N_9209,N_9119);
xor U11105 (N_11105,N_9699,N_8907);
nor U11106 (N_11106,N_6211,N_7333);
or U11107 (N_11107,N_9621,N_7786);
xnor U11108 (N_11108,N_8644,N_9110);
nor U11109 (N_11109,N_6971,N_9903);
xor U11110 (N_11110,N_9193,N_6795);
nand U11111 (N_11111,N_6182,N_7454);
xor U11112 (N_11112,N_6540,N_5161);
and U11113 (N_11113,N_5571,N_9028);
and U11114 (N_11114,N_5201,N_8179);
or U11115 (N_11115,N_6787,N_9746);
xor U11116 (N_11116,N_6189,N_9115);
xor U11117 (N_11117,N_7330,N_5658);
xor U11118 (N_11118,N_5150,N_9291);
and U11119 (N_11119,N_8910,N_7574);
or U11120 (N_11120,N_6441,N_9854);
xnor U11121 (N_11121,N_8709,N_7467);
and U11122 (N_11122,N_9118,N_8682);
nand U11123 (N_11123,N_8559,N_7001);
nor U11124 (N_11124,N_6105,N_8449);
nand U11125 (N_11125,N_6319,N_9997);
nor U11126 (N_11126,N_5279,N_5756);
nor U11127 (N_11127,N_6031,N_8462);
and U11128 (N_11128,N_6407,N_5951);
nand U11129 (N_11129,N_5985,N_6675);
or U11130 (N_11130,N_5258,N_7179);
xnor U11131 (N_11131,N_7025,N_8502);
and U11132 (N_11132,N_8290,N_9636);
xor U11133 (N_11133,N_8844,N_7361);
nand U11134 (N_11134,N_6050,N_8811);
or U11135 (N_11135,N_6272,N_9557);
xor U11136 (N_11136,N_6476,N_8433);
xnor U11137 (N_11137,N_7918,N_8156);
nand U11138 (N_11138,N_6234,N_5352);
and U11139 (N_11139,N_7584,N_5061);
nand U11140 (N_11140,N_8743,N_5643);
or U11141 (N_11141,N_6825,N_7038);
xor U11142 (N_11142,N_7354,N_8702);
and U11143 (N_11143,N_6768,N_7268);
and U11144 (N_11144,N_8138,N_8434);
nand U11145 (N_11145,N_5833,N_9966);
xor U11146 (N_11146,N_9235,N_8982);
nand U11147 (N_11147,N_8266,N_6365);
nor U11148 (N_11148,N_9897,N_6583);
or U11149 (N_11149,N_6337,N_8221);
or U11150 (N_11150,N_9144,N_9724);
and U11151 (N_11151,N_9389,N_6498);
or U11152 (N_11152,N_6593,N_8191);
or U11153 (N_11153,N_5074,N_9865);
nor U11154 (N_11154,N_8453,N_8847);
or U11155 (N_11155,N_7671,N_6934);
or U11156 (N_11156,N_8611,N_6289);
nand U11157 (N_11157,N_5066,N_6134);
nor U11158 (N_11158,N_7907,N_5138);
and U11159 (N_11159,N_9410,N_8227);
or U11160 (N_11160,N_5864,N_8159);
and U11161 (N_11161,N_5873,N_7139);
and U11162 (N_11162,N_5400,N_8828);
nand U11163 (N_11163,N_9268,N_7542);
or U11164 (N_11164,N_5326,N_9276);
nand U11165 (N_11165,N_7783,N_6443);
nand U11166 (N_11166,N_6903,N_7429);
nand U11167 (N_11167,N_7787,N_7914);
xor U11168 (N_11168,N_5912,N_8942);
and U11169 (N_11169,N_5926,N_7952);
xnor U11170 (N_11170,N_8148,N_8441);
xor U11171 (N_11171,N_6431,N_6486);
and U11172 (N_11172,N_9851,N_9393);
and U11173 (N_11173,N_5994,N_5920);
nand U11174 (N_11174,N_6458,N_7870);
xor U11175 (N_11175,N_9932,N_5100);
nand U11176 (N_11176,N_6198,N_5746);
nor U11177 (N_11177,N_5517,N_7600);
nand U11178 (N_11178,N_7799,N_9608);
and U11179 (N_11179,N_9315,N_9893);
nand U11180 (N_11180,N_8883,N_9695);
xnor U11181 (N_11181,N_6528,N_9784);
xor U11182 (N_11182,N_9067,N_7773);
or U11183 (N_11183,N_7889,N_6945);
xnor U11184 (N_11184,N_7537,N_6444);
and U11185 (N_11185,N_9939,N_7807);
xor U11186 (N_11186,N_7734,N_6892);
or U11187 (N_11187,N_7612,N_6570);
and U11188 (N_11188,N_8389,N_5105);
and U11189 (N_11189,N_6218,N_8948);
nor U11190 (N_11190,N_6851,N_5928);
nand U11191 (N_11191,N_9731,N_9481);
and U11192 (N_11192,N_7305,N_5489);
nand U11193 (N_11193,N_6032,N_6982);
or U11194 (N_11194,N_8776,N_7971);
xnor U11195 (N_11195,N_7701,N_6954);
nor U11196 (N_11196,N_8114,N_5156);
and U11197 (N_11197,N_5334,N_6855);
xnor U11198 (N_11198,N_8240,N_6397);
and U11199 (N_11199,N_7200,N_8297);
and U11200 (N_11200,N_5033,N_7219);
nand U11201 (N_11201,N_5175,N_9579);
and U11202 (N_11202,N_8496,N_7032);
nand U11203 (N_11203,N_6164,N_7808);
and U11204 (N_11204,N_9643,N_7169);
nor U11205 (N_11205,N_5324,N_6303);
nand U11206 (N_11206,N_6107,N_6147);
or U11207 (N_11207,N_8655,N_6136);
or U11208 (N_11208,N_9567,N_8707);
and U11209 (N_11209,N_7265,N_8492);
or U11210 (N_11210,N_6698,N_6859);
nor U11211 (N_11211,N_7003,N_7447);
nand U11212 (N_11212,N_8768,N_9655);
nor U11213 (N_11213,N_9124,N_5002);
or U11214 (N_11214,N_9070,N_8854);
nor U11215 (N_11215,N_5426,N_8209);
xor U11216 (N_11216,N_5470,N_8908);
or U11217 (N_11217,N_7609,N_8342);
xor U11218 (N_11218,N_6908,N_8916);
xnor U11219 (N_11219,N_6927,N_5813);
nand U11220 (N_11220,N_6889,N_9628);
or U11221 (N_11221,N_7628,N_6660);
or U11222 (N_11222,N_5992,N_9324);
or U11223 (N_11223,N_7183,N_5265);
and U11224 (N_11224,N_9705,N_8470);
and U11225 (N_11225,N_7206,N_8984);
nor U11226 (N_11226,N_6359,N_6574);
and U11227 (N_11227,N_6874,N_8394);
nor U11228 (N_11228,N_7841,N_6180);
nand U11229 (N_11229,N_5097,N_5389);
xnor U11230 (N_11230,N_7743,N_5307);
nor U11231 (N_11231,N_6661,N_8063);
nand U11232 (N_11232,N_8963,N_8893);
and U11233 (N_11233,N_7608,N_5110);
nor U11234 (N_11234,N_8523,N_6381);
nand U11235 (N_11235,N_9979,N_9161);
xor U11236 (N_11236,N_9896,N_5796);
xnor U11237 (N_11237,N_9728,N_8582);
nand U11238 (N_11238,N_9733,N_9578);
or U11239 (N_11239,N_6068,N_5480);
nor U11240 (N_11240,N_7887,N_5380);
xnor U11241 (N_11241,N_5067,N_7554);
xnor U11242 (N_11242,N_6326,N_9611);
or U11243 (N_11243,N_9159,N_8839);
nor U11244 (N_11244,N_7229,N_9261);
nand U11245 (N_11245,N_5484,N_5678);
nor U11246 (N_11246,N_5565,N_9971);
nand U11247 (N_11247,N_6388,N_6309);
nand U11248 (N_11248,N_9286,N_6343);
nor U11249 (N_11249,N_5035,N_9902);
or U11250 (N_11250,N_7925,N_7745);
or U11251 (N_11251,N_8082,N_9047);
nand U11252 (N_11252,N_7527,N_7873);
or U11253 (N_11253,N_7123,N_8914);
or U11254 (N_11254,N_7934,N_7509);
nor U11255 (N_11255,N_9874,N_9947);
or U11256 (N_11256,N_6714,N_6818);
or U11257 (N_11257,N_9246,N_5136);
or U11258 (N_11258,N_6534,N_6511);
or U11259 (N_11259,N_5047,N_8036);
xnor U11260 (N_11260,N_6214,N_5057);
nor U11261 (N_11261,N_6547,N_9169);
nor U11262 (N_11262,N_6965,N_8814);
or U11263 (N_11263,N_9895,N_7163);
and U11264 (N_11264,N_9390,N_9403);
nand U11265 (N_11265,N_5633,N_5511);
nor U11266 (N_11266,N_7777,N_9530);
or U11267 (N_11267,N_5364,N_5790);
nor U11268 (N_11268,N_9532,N_6419);
and U11269 (N_11269,N_6448,N_9083);
xnor U11270 (N_11270,N_7736,N_8684);
and U11271 (N_11271,N_5909,N_6932);
or U11272 (N_11272,N_8909,N_8627);
and U11273 (N_11273,N_7355,N_8377);
and U11274 (N_11274,N_5273,N_7294);
or U11275 (N_11275,N_6654,N_7424);
or U11276 (N_11276,N_8609,N_7933);
xor U11277 (N_11277,N_6789,N_5862);
or U11278 (N_11278,N_9302,N_9445);
or U11279 (N_11279,N_7744,N_6481);
and U11280 (N_11280,N_5904,N_5050);
xnor U11281 (N_11281,N_7898,N_8475);
or U11282 (N_11282,N_9742,N_7693);
or U11283 (N_11283,N_6410,N_7486);
nor U11284 (N_11284,N_6079,N_8012);
nor U11285 (N_11285,N_8647,N_8926);
and U11286 (N_11286,N_7262,N_9343);
nor U11287 (N_11287,N_9969,N_7286);
and U11288 (N_11288,N_6783,N_6996);
nand U11289 (N_11289,N_5212,N_5555);
nand U11290 (N_11290,N_5409,N_8538);
nand U11291 (N_11291,N_6315,N_6332);
xor U11292 (N_11292,N_6731,N_9340);
or U11293 (N_11293,N_8670,N_9928);
and U11294 (N_11294,N_5894,N_7619);
xnor U11295 (N_11295,N_8263,N_5359);
nor U11296 (N_11296,N_7500,N_9559);
xnor U11297 (N_11297,N_6876,N_5520);
xnor U11298 (N_11298,N_6493,N_5248);
nand U11299 (N_11299,N_9623,N_6956);
nand U11300 (N_11300,N_7529,N_9756);
nand U11301 (N_11301,N_5757,N_9503);
or U11302 (N_11302,N_5206,N_8777);
and U11303 (N_11303,N_8880,N_8543);
nor U11304 (N_11304,N_8161,N_5801);
nor U11305 (N_11305,N_5403,N_8816);
nor U11306 (N_11306,N_6915,N_7116);
nand U11307 (N_11307,N_5647,N_8129);
nor U11308 (N_11308,N_9829,N_9345);
xnor U11309 (N_11309,N_5189,N_9474);
nand U11310 (N_11310,N_7071,N_8084);
xor U11311 (N_11311,N_9035,N_5397);
xor U11312 (N_11312,N_9568,N_5903);
and U11313 (N_11313,N_9722,N_5068);
and U11314 (N_11314,N_5241,N_9417);
nand U11315 (N_11315,N_9349,N_9018);
and U11316 (N_11316,N_9101,N_9258);
or U11317 (N_11317,N_5880,N_6051);
and U11318 (N_11318,N_6278,N_6906);
nand U11319 (N_11319,N_9379,N_9861);
or U11320 (N_11320,N_6022,N_8734);
nand U11321 (N_11321,N_8640,N_6821);
or U11322 (N_11322,N_8070,N_8514);
or U11323 (N_11323,N_5500,N_9399);
xor U11324 (N_11324,N_7604,N_8123);
nand U11325 (N_11325,N_9479,N_9501);
or U11326 (N_11326,N_9983,N_6918);
and U11327 (N_11327,N_5755,N_9824);
or U11328 (N_11328,N_5371,N_5172);
nor U11329 (N_11329,N_9657,N_9200);
and U11330 (N_11330,N_8668,N_8592);
nand U11331 (N_11331,N_9666,N_9587);
and U11332 (N_11332,N_5682,N_6750);
xor U11333 (N_11333,N_7061,N_8349);
nor U11334 (N_11334,N_5655,N_8902);
xor U11335 (N_11335,N_6883,N_9668);
nor U11336 (N_11336,N_9813,N_9549);
xor U11337 (N_11337,N_5090,N_8642);
nor U11338 (N_11338,N_8947,N_7911);
nor U11339 (N_11339,N_6682,N_5142);
nand U11340 (N_11340,N_7501,N_7502);
xor U11341 (N_11341,N_8146,N_7653);
xor U11342 (N_11342,N_8596,N_9941);
xor U11343 (N_11343,N_8390,N_8855);
nand U11344 (N_11344,N_8339,N_7579);
nand U11345 (N_11345,N_5162,N_9515);
and U11346 (N_11346,N_5453,N_7427);
and U11347 (N_11347,N_5245,N_6813);
nor U11348 (N_11348,N_8308,N_7975);
nand U11349 (N_11349,N_5741,N_7705);
and U11350 (N_11350,N_8843,N_7058);
or U11351 (N_11351,N_6287,N_8317);
or U11352 (N_11352,N_5535,N_8767);
and U11353 (N_11353,N_7461,N_9242);
and U11354 (N_11354,N_8955,N_5758);
nor U11355 (N_11355,N_5464,N_8771);
xnor U11356 (N_11356,N_5184,N_8979);
nor U11357 (N_11357,N_8551,N_7005);
or U11358 (N_11358,N_6013,N_5072);
nand U11359 (N_11359,N_5516,N_7292);
nand U11360 (N_11360,N_9858,N_6037);
nand U11361 (N_11361,N_8507,N_5578);
xnor U11362 (N_11362,N_6943,N_9706);
nor U11363 (N_11363,N_8677,N_6727);
xnor U11364 (N_11364,N_9447,N_8727);
nand U11365 (N_11365,N_9550,N_9510);
nor U11366 (N_11366,N_9237,N_6271);
and U11367 (N_11367,N_8295,N_9060);
and U11368 (N_11368,N_6006,N_7157);
nand U11369 (N_11369,N_9428,N_6118);
nor U11370 (N_11370,N_9768,N_8697);
or U11371 (N_11371,N_8700,N_9135);
nand U11372 (N_11372,N_9121,N_5638);
and U11373 (N_11373,N_6024,N_8397);
xor U11374 (N_11374,N_8812,N_8930);
and U11375 (N_11375,N_7588,N_5791);
or U11376 (N_11376,N_8857,N_7929);
and U11377 (N_11377,N_5412,N_8708);
and U11378 (N_11378,N_6747,N_6778);
nor U11379 (N_11379,N_8232,N_7956);
nor U11380 (N_11380,N_8556,N_6655);
and U11381 (N_11381,N_6882,N_8778);
and U11382 (N_11382,N_7959,N_5229);
xnor U11383 (N_11383,N_5594,N_6123);
or U11384 (N_11384,N_6177,N_9309);
nand U11385 (N_11385,N_6030,N_7382);
and U11386 (N_11386,N_7657,N_8983);
and U11387 (N_11387,N_9208,N_8614);
nand U11388 (N_11388,N_9913,N_7553);
xnor U11389 (N_11389,N_6901,N_9778);
or U11390 (N_11390,N_9221,N_5182);
or U11391 (N_11391,N_6871,N_9487);
nand U11392 (N_11392,N_8725,N_6755);
nor U11393 (N_11393,N_8705,N_9886);
or U11394 (N_11394,N_6310,N_5720);
or U11395 (N_11395,N_6494,N_7207);
and U11396 (N_11396,N_5621,N_8338);
nand U11397 (N_11397,N_9592,N_5684);
nand U11398 (N_11398,N_6553,N_5347);
and U11399 (N_11399,N_8529,N_9334);
xnor U11400 (N_11400,N_7011,N_8432);
and U11401 (N_11401,N_8836,N_6995);
nor U11402 (N_11402,N_7530,N_8840);
nor U11403 (N_11403,N_9832,N_6751);
nor U11404 (N_11404,N_5780,N_8378);
or U11405 (N_11405,N_8563,N_6662);
xor U11406 (N_11406,N_7731,N_5232);
nor U11407 (N_11407,N_8666,N_5493);
and U11408 (N_11408,N_5030,N_8334);
xor U11409 (N_11409,N_6801,N_6979);
or U11410 (N_11410,N_8248,N_7374);
nand U11411 (N_11411,N_6565,N_9975);
or U11412 (N_11412,N_8412,N_5286);
xor U11413 (N_11413,N_7646,N_5277);
xor U11414 (N_11414,N_8672,N_5186);
nand U11415 (N_11415,N_6820,N_6436);
and U11416 (N_11416,N_8181,N_7680);
nand U11417 (N_11417,N_7921,N_8937);
or U11418 (N_11418,N_7295,N_9763);
nand U11419 (N_11419,N_6219,N_5402);
xor U11420 (N_11420,N_8569,N_5902);
nand U11421 (N_11421,N_5437,N_8694);
nor U11422 (N_11422,N_9962,N_9541);
nand U11423 (N_11423,N_8775,N_9112);
or U11424 (N_11424,N_7362,N_9408);
nand U11425 (N_11425,N_5837,N_7414);
xnor U11426 (N_11426,N_9959,N_8029);
or U11427 (N_11427,N_6059,N_7882);
or U11428 (N_11428,N_7091,N_7185);
or U11429 (N_11429,N_9989,N_7670);
xnor U11430 (N_11430,N_6249,N_6711);
nand U11431 (N_11431,N_8960,N_7073);
or U11432 (N_11432,N_6350,N_8863);
nand U11433 (N_11433,N_6972,N_8078);
nor U11434 (N_11434,N_9791,N_7076);
nand U11435 (N_11435,N_9416,N_6758);
and U11436 (N_11436,N_5641,N_7287);
nand U11437 (N_11437,N_7757,N_9899);
or U11438 (N_11438,N_6157,N_5538);
and U11439 (N_11439,N_9446,N_9142);
nand U11440 (N_11440,N_8480,N_8762);
xnor U11441 (N_11441,N_8018,N_8456);
xor U11442 (N_11442,N_6264,N_8726);
or U11443 (N_11443,N_7199,N_9175);
nor U11444 (N_11444,N_7406,N_5078);
and U11445 (N_11445,N_8335,N_5499);
nor U11446 (N_11446,N_8328,N_7960);
xor U11447 (N_11447,N_9075,N_9266);
nand U11448 (N_11448,N_8827,N_9162);
and U11449 (N_11449,N_8223,N_6793);
and U11450 (N_11450,N_7174,N_7089);
nor U11451 (N_11451,N_5844,N_7881);
nor U11452 (N_11452,N_7364,N_5996);
or U11453 (N_11453,N_7270,N_6322);
nor U11454 (N_11454,N_5041,N_6014);
nand U11455 (N_11455,N_5531,N_8796);
or U11456 (N_11456,N_7214,N_5203);
and U11457 (N_11457,N_8418,N_7456);
nor U11458 (N_11458,N_8570,N_7515);
and U11459 (N_11459,N_6109,N_6477);
and U11460 (N_11460,N_9485,N_8011);
and U11461 (N_11461,N_6485,N_8962);
or U11462 (N_11462,N_5567,N_8932);
or U11463 (N_11463,N_8956,N_7164);
nor U11464 (N_11464,N_9661,N_7154);
nand U11465 (N_11465,N_9910,N_5305);
nor U11466 (N_11466,N_9803,N_7079);
nand U11467 (N_11467,N_9660,N_6763);
or U11468 (N_11468,N_7910,N_9937);
nor U11469 (N_11469,N_5929,N_6411);
xor U11470 (N_11470,N_9381,N_6693);
nand U11471 (N_11471,N_7002,N_9259);
nor U11472 (N_11472,N_5052,N_5766);
nand U11473 (N_11473,N_5745,N_8526);
nand U11474 (N_11474,N_7901,N_5456);
and U11475 (N_11475,N_6590,N_8113);
or U11476 (N_11476,N_6902,N_8188);
or U11477 (N_11477,N_8873,N_6454);
or U11478 (N_11478,N_5805,N_8086);
and U11479 (N_11479,N_5016,N_7483);
xnor U11480 (N_11480,N_6770,N_9957);
xor U11481 (N_11481,N_9625,N_7626);
nand U11482 (N_11482,N_8155,N_7602);
or U11483 (N_11483,N_9433,N_9308);
and U11484 (N_11484,N_6434,N_7160);
nand U11485 (N_11485,N_7767,N_6465);
or U11486 (N_11486,N_9604,N_7806);
nor U11487 (N_11487,N_5961,N_8024);
xnor U11488 (N_11488,N_7067,N_8524);
nand U11489 (N_11489,N_7943,N_8116);
and U11490 (N_11490,N_8244,N_7591);
or U11491 (N_11491,N_5407,N_9086);
nand U11492 (N_11492,N_6026,N_5540);
xor U11493 (N_11493,N_6626,N_8711);
xnor U11494 (N_11494,N_9909,N_5534);
xnor U11495 (N_11495,N_8715,N_9326);
or U11496 (N_11496,N_7507,N_6297);
and U11497 (N_11497,N_5772,N_6117);
xnor U11498 (N_11498,N_5251,N_6414);
and U11499 (N_11499,N_7119,N_9153);
xor U11500 (N_11500,N_5814,N_6181);
xnor U11501 (N_11501,N_6910,N_8020);
nand U11502 (N_11502,N_6438,N_7173);
nand U11503 (N_11503,N_8316,N_9696);
nand U11504 (N_11504,N_9601,N_6102);
nor U11505 (N_11505,N_5669,N_8031);
xnor U11506 (N_11506,N_8204,N_7476);
and U11507 (N_11507,N_9396,N_8864);
and U11508 (N_11508,N_8385,N_6623);
or U11509 (N_11509,N_9160,N_6994);
and U11510 (N_11510,N_7610,N_8162);
nor U11511 (N_11511,N_6004,N_6265);
nand U11512 (N_11512,N_6502,N_5707);
nand U11513 (N_11513,N_5415,N_9531);
nand U11514 (N_11514,N_8900,N_8079);
and U11515 (N_11515,N_5861,N_6235);
nand U11516 (N_11516,N_5884,N_9298);
nand U11517 (N_11517,N_5143,N_9974);
and U11518 (N_11518,N_7291,N_8833);
and U11519 (N_11519,N_9049,N_8169);
nor U11520 (N_11520,N_7684,N_8383);
and U11521 (N_11521,N_8837,N_6126);
or U11522 (N_11522,N_8322,N_5752);
and U11523 (N_11523,N_5085,N_9892);
and U11524 (N_11524,N_9093,N_6576);
or U11525 (N_11525,N_6325,N_9700);
and U11526 (N_11526,N_7536,N_8584);
nor U11527 (N_11527,N_5648,N_6647);
xnor U11528 (N_11528,N_9499,N_7332);
nand U11529 (N_11529,N_9955,N_9846);
nand U11530 (N_11530,N_9970,N_9817);
and U11531 (N_11531,N_7822,N_8430);
and U11532 (N_11532,N_7915,N_7639);
and U11533 (N_11533,N_7555,N_6706);
or U11534 (N_11534,N_9325,N_7539);
nor U11535 (N_11535,N_7978,N_8242);
nand U11536 (N_11536,N_7633,N_7661);
and U11537 (N_11537,N_9054,N_8351);
and U11538 (N_11538,N_5646,N_9553);
or U11539 (N_11539,N_9574,N_6897);
nor U11540 (N_11540,N_7759,N_8474);
xnor U11541 (N_11541,N_5494,N_6790);
and U11542 (N_11542,N_8822,N_7867);
or U11543 (N_11543,N_5973,N_6048);
nand U11544 (N_11544,N_7955,N_6318);
xor U11545 (N_11545,N_9234,N_9519);
or U11546 (N_11546,N_6412,N_5384);
nor U11547 (N_11547,N_5095,N_9619);
nor U11548 (N_11548,N_5454,N_7369);
and U11549 (N_11549,N_7212,N_6484);
xnor U11550 (N_11550,N_5422,N_7837);
and U11551 (N_11551,N_9017,N_9380);
and U11552 (N_11552,N_5972,N_8969);
nor U11553 (N_11553,N_7996,N_9825);
nor U11554 (N_11554,N_7016,N_6340);
xnor U11555 (N_11555,N_5918,N_9785);
nand U11556 (N_11556,N_5327,N_8759);
nand U11557 (N_11557,N_9068,N_7749);
or U11558 (N_11558,N_6049,N_7899);
nand U11559 (N_11559,N_7719,N_9631);
and U11560 (N_11560,N_9123,N_5759);
nand U11561 (N_11561,N_8173,N_5588);
nor U11562 (N_11562,N_7794,N_9609);
nor U11563 (N_11563,N_7669,N_6335);
xor U11564 (N_11564,N_6962,N_8304);
and U11565 (N_11565,N_7559,N_9711);
or U11566 (N_11566,N_7834,N_6609);
nand U11567 (N_11567,N_9295,N_8392);
and U11568 (N_11568,N_7762,N_5195);
nand U11569 (N_11569,N_6452,N_5670);
xnor U11570 (N_11570,N_7014,N_7849);
xnor U11571 (N_11571,N_6028,N_8457);
nor U11572 (N_11572,N_6887,N_9051);
nand U11573 (N_11573,N_7520,N_8675);
nor U11574 (N_11574,N_7752,N_9772);
nor U11575 (N_11575,N_6372,N_7741);
and U11576 (N_11576,N_9869,N_7840);
nor U11577 (N_11577,N_9956,N_6139);
nor U11578 (N_11578,N_6081,N_5267);
or U11579 (N_11579,N_7638,N_7051);
and U11580 (N_11580,N_8262,N_6158);
xnor U11581 (N_11581,N_6953,N_8599);
and U11582 (N_11582,N_9518,N_7652);
nand U11583 (N_11583,N_8501,N_8247);
or U11584 (N_11584,N_9150,N_5938);
xnor U11585 (N_11585,N_5949,N_8305);
xor U11586 (N_11586,N_7409,N_6153);
or U11587 (N_11587,N_6215,N_6745);
and U11588 (N_11588,N_7288,N_8326);
xnor U11589 (N_11589,N_7465,N_8446);
nand U11590 (N_11590,N_7909,N_8601);
and U11591 (N_11591,N_6797,N_7256);
and U11592 (N_11592,N_8766,N_5194);
nor U11593 (N_11593,N_5311,N_6704);
nor U11594 (N_11594,N_5982,N_7433);
nand U11595 (N_11595,N_6931,N_6746);
or U11596 (N_11596,N_9425,N_7605);
and U11597 (N_11597,N_6627,N_9128);
nand U11598 (N_11598,N_9614,N_5485);
xor U11599 (N_11599,N_8201,N_7913);
or U11600 (N_11600,N_7821,N_8329);
and U11601 (N_11601,N_5787,N_9352);
nand U11602 (N_11602,N_8345,N_6709);
nand U11603 (N_11603,N_7728,N_6756);
nor U11604 (N_11604,N_5181,N_5583);
or U11605 (N_11605,N_8890,N_9659);
xor U11606 (N_11606,N_8636,N_8325);
nor U11607 (N_11607,N_8180,N_6666);
nor U11608 (N_11608,N_8667,N_8607);
or U11609 (N_11609,N_7647,N_6517);
nor U11610 (N_11610,N_6947,N_8809);
nor U11611 (N_11611,N_8595,N_7075);
nor U11612 (N_11612,N_9795,N_6926);
nand U11613 (N_11613,N_9509,N_8632);
nand U11614 (N_11614,N_9038,N_6488);
and U11615 (N_11615,N_6951,N_7182);
nor U11616 (N_11616,N_9338,N_7106);
nor U11617 (N_11617,N_6229,N_5390);
nand U11618 (N_11618,N_5233,N_9542);
nor U11619 (N_11619,N_7049,N_8757);
or U11620 (N_11620,N_8733,N_9732);
nor U11621 (N_11621,N_9656,N_5222);
and U11622 (N_11622,N_5724,N_7992);
or U11623 (N_11623,N_5832,N_5566);
nor U11624 (N_11624,N_5393,N_8171);
or U11625 (N_11625,N_5879,N_8346);
or U11626 (N_11626,N_8233,N_6748);
nand U11627 (N_11627,N_5332,N_5577);
nand U11628 (N_11628,N_9289,N_8225);
or U11629 (N_11629,N_9674,N_7329);
nor U11630 (N_11630,N_8203,N_7248);
and U11631 (N_11631,N_8695,N_9096);
xor U11632 (N_11632,N_9994,N_8088);
or U11633 (N_11633,N_8738,N_6064);
nand U11634 (N_11634,N_9290,N_9605);
nor U11635 (N_11635,N_9718,N_9820);
nor U11636 (N_11636,N_7801,N_8006);
xnor U11637 (N_11637,N_9126,N_7363);
nor U11638 (N_11638,N_5515,N_8945);
nand U11639 (N_11639,N_5367,N_7590);
and U11640 (N_11640,N_9366,N_5605);
xor U11641 (N_11641,N_8521,N_8282);
nand U11642 (N_11642,N_7479,N_5875);
and U11643 (N_11643,N_7624,N_8354);
nor U11644 (N_11644,N_5585,N_5411);
nor U11645 (N_11645,N_9484,N_6992);
or U11646 (N_11646,N_8395,N_5446);
nand U11647 (N_11647,N_5860,N_9996);
nor U11648 (N_11648,N_8981,N_7312);
and U11649 (N_11649,N_8594,N_8040);
xor U11650 (N_11650,N_5169,N_8053);
and U11651 (N_11651,N_9458,N_5185);
and U11652 (N_11652,N_8440,N_6191);
nor U11653 (N_11653,N_6645,N_5051);
or U11654 (N_11654,N_5590,N_8699);
and U11655 (N_11655,N_8141,N_5115);
xor U11656 (N_11656,N_6468,N_9527);
nor U11657 (N_11657,N_8639,N_7954);
nor U11658 (N_11658,N_5675,N_9480);
nand U11659 (N_11659,N_7769,N_7277);
xnor U11660 (N_11660,N_9012,N_5278);
or U11661 (N_11661,N_7410,N_7569);
nand U11662 (N_11662,N_5997,N_7020);
nor U11663 (N_11663,N_6083,N_8032);
xor U11664 (N_11664,N_5486,N_7643);
xnor U11665 (N_11665,N_7853,N_8506);
xor U11666 (N_11666,N_8681,N_6321);
and U11667 (N_11667,N_9252,N_5681);
and U11668 (N_11668,N_8853,N_8222);
or U11669 (N_11669,N_9919,N_5134);
nand U11670 (N_11670,N_9493,N_8458);
nor U11671 (N_11671,N_5526,N_8719);
or U11672 (N_11672,N_9216,N_9917);
nand U11673 (N_11673,N_9787,N_8407);
or U11674 (N_11674,N_5266,N_6836);
xnor U11675 (N_11675,N_8264,N_8213);
or U11676 (N_11676,N_7093,N_7172);
and U11677 (N_11677,N_5661,N_6998);
or U11678 (N_11678,N_7967,N_5076);
nor U11679 (N_11679,N_6612,N_6726);
or U11680 (N_11680,N_6269,N_6091);
xnor U11681 (N_11681,N_9805,N_5032);
or U11682 (N_11682,N_8439,N_5003);
xor U11683 (N_11683,N_9021,N_8459);
nor U11684 (N_11684,N_8729,N_9294);
or U11685 (N_11685,N_7133,N_7451);
or U11686 (N_11686,N_9134,N_8861);
or U11687 (N_11687,N_5227,N_6480);
and U11688 (N_11688,N_8552,N_7800);
nand U11689 (N_11689,N_6208,N_5637);
nand U11690 (N_11690,N_6610,N_5019);
or U11691 (N_11691,N_7055,N_6239);
xnor U11692 (N_11692,N_6178,N_9776);
or U11693 (N_11693,N_5146,N_8579);
or U11694 (N_11694,N_7166,N_6067);
xor U11695 (N_11695,N_6781,N_7246);
and U11696 (N_11696,N_5254,N_7188);
or U11697 (N_11697,N_6946,N_8752);
xnor U11698 (N_11698,N_7360,N_7768);
or U11699 (N_11699,N_9818,N_8689);
or U11700 (N_11700,N_9801,N_8293);
or U11701 (N_11701,N_9954,N_5147);
nand U11702 (N_11702,N_8436,N_6472);
or U11703 (N_11703,N_9552,N_5000);
nor U11704 (N_11704,N_7496,N_7345);
xor U11705 (N_11705,N_5651,N_7998);
nand U11706 (N_11706,N_7506,N_8090);
or U11707 (N_11707,N_6399,N_9071);
or U11708 (N_11708,N_8603,N_9569);
nor U11709 (N_11709,N_5846,N_6684);
nand U11710 (N_11710,N_7111,N_5925);
xnor U11711 (N_11711,N_9025,N_9422);
nand U11712 (N_11712,N_6422,N_5092);
xor U11713 (N_11713,N_9170,N_7107);
or U11714 (N_11714,N_8838,N_8952);
or U11715 (N_11715,N_5360,N_9761);
xnor U11716 (N_11716,N_5710,N_9449);
or U11717 (N_11717,N_9616,N_6132);
xnor U11718 (N_11718,N_5008,N_5967);
nand U11719 (N_11719,N_6513,N_6890);
xnor U11720 (N_11720,N_7181,N_6539);
and U11721 (N_11721,N_5020,N_9419);
and U11722 (N_11722,N_6295,N_9274);
or U11723 (N_11723,N_6628,N_5686);
xnor U11724 (N_11724,N_8578,N_5469);
nor U11725 (N_11725,N_5476,N_7443);
nand U11726 (N_11726,N_6782,N_7436);
xnor U11727 (N_11727,N_9985,N_7857);
nand U11728 (N_11728,N_6506,N_6003);
nor U11729 (N_11729,N_6742,N_5693);
xor U11730 (N_11730,N_5059,N_9800);
nor U11731 (N_11731,N_5802,N_6302);
xor U11732 (N_11732,N_5361,N_9157);
nand U11733 (N_11733,N_7685,N_5927);
and U11734 (N_11734,N_5037,N_9010);
nor U11735 (N_11735,N_7077,N_5742);
xnor U11736 (N_11736,N_7441,N_6133);
nand U11737 (N_11737,N_8938,N_5554);
and U11738 (N_11738,N_7152,N_9921);
nor U11739 (N_11739,N_6143,N_5586);
nor U11740 (N_11740,N_7724,N_8269);
nand U11741 (N_11741,N_6816,N_7981);
and U11742 (N_11742,N_8678,N_5734);
nor U11743 (N_11743,N_9916,N_6986);
or U11744 (N_11744,N_6044,N_9754);
xor U11745 (N_11745,N_6284,N_7557);
nor U11746 (N_11746,N_9753,N_8959);
nor U11747 (N_11747,N_6581,N_5639);
or U11748 (N_11748,N_5268,N_6362);
or U11749 (N_11749,N_9968,N_7186);
nor U11750 (N_11750,N_8742,N_7195);
and U11751 (N_11751,N_9077,N_6285);
nand U11752 (N_11752,N_8903,N_5525);
xnor U11753 (N_11753,N_8379,N_5989);
nor U11754 (N_11754,N_6673,N_6247);
or U11755 (N_11755,N_8144,N_7906);
and U11756 (N_11756,N_6114,N_6595);
nor U11757 (N_11757,N_8905,N_9042);
or U11758 (N_11758,N_7393,N_9771);
and U11759 (N_11759,N_8022,N_8460);
or U11760 (N_11760,N_5288,N_7380);
xnor U11761 (N_11761,N_8157,N_9683);
and U11762 (N_11762,N_9104,N_8820);
and U11763 (N_11763,N_9836,N_6715);
or U11764 (N_11764,N_7141,N_9688);
or U11765 (N_11765,N_8437,N_8567);
or U11766 (N_11766,N_9048,N_6475);
and U11767 (N_11767,N_6027,N_7334);
nand U11768 (N_11768,N_9257,N_5944);
or U11769 (N_11769,N_7068,N_5013);
or U11770 (N_11770,N_7516,N_9316);
or U11771 (N_11771,N_8045,N_9663);
or U11772 (N_11772,N_9253,N_8793);
nor U11773 (N_11773,N_7167,N_8442);
nor U11774 (N_11774,N_5200,N_8211);
or U11775 (N_11775,N_7105,N_8275);
or U11776 (N_11776,N_8309,N_6334);
nand U11777 (N_11777,N_9317,N_6185);
nand U11778 (N_11778,N_9736,N_6075);
and U11779 (N_11779,N_7275,N_8819);
nor U11780 (N_11780,N_5924,N_5510);
nand U11781 (N_11781,N_9336,N_6922);
and U11782 (N_11782,N_6562,N_8028);
nand U11783 (N_11783,N_5075,N_8164);
or U11784 (N_11784,N_9888,N_6267);
and U11785 (N_11785,N_9363,N_8503);
xnor U11786 (N_11786,N_9544,N_9684);
xor U11787 (N_11787,N_9271,N_6328);
nand U11788 (N_11788,N_5174,N_8895);
and U11789 (N_11789,N_6904,N_7178);
xnor U11790 (N_11790,N_8548,N_7236);
xor U11791 (N_11791,N_5064,N_8292);
xnor U11792 (N_11792,N_9612,N_5782);
nor U11793 (N_11793,N_8653,N_5368);
nor U11794 (N_11794,N_9664,N_5786);
nand U11795 (N_11795,N_5911,N_6508);
and U11796 (N_11796,N_9164,N_6457);
xnor U11797 (N_11797,N_6256,N_9606);
nand U11798 (N_11798,N_7789,N_6430);
nand U11799 (N_11799,N_6033,N_8323);
nor U11800 (N_11800,N_8988,N_5523);
nand U11801 (N_11801,N_7885,N_5045);
or U11802 (N_11802,N_7957,N_7047);
or U11803 (N_11803,N_7446,N_5024);
nand U11804 (N_11804,N_5432,N_6501);
nand U11805 (N_11805,N_8972,N_9329);
nand U11806 (N_11806,N_9172,N_5930);
nand U11807 (N_11807,N_9248,N_9056);
nor U11808 (N_11808,N_7065,N_7687);
xor U11809 (N_11809,N_5536,N_8226);
or U11810 (N_11810,N_8163,N_5612);
and U11811 (N_11811,N_6823,N_5708);
nand U11812 (N_11812,N_8995,N_9950);
and U11813 (N_11813,N_5004,N_9944);
nor U11814 (N_11814,N_5739,N_5121);
or U11815 (N_11815,N_8688,N_8367);
and U11816 (N_11816,N_6052,N_8929);
nand U11817 (N_11817,N_7289,N_8451);
or U11818 (N_11818,N_7614,N_7279);
and U11819 (N_11819,N_7846,N_9632);
nand U11820 (N_11820,N_7665,N_7805);
xnor U11821 (N_11821,N_7316,N_9502);
or U11822 (N_11822,N_5378,N_6875);
xnor U11823 (N_11823,N_9155,N_6324);
xnor U11824 (N_11824,N_8477,N_7620);
xnor U11825 (N_11825,N_6261,N_9311);
nand U11826 (N_11826,N_8149,N_7149);
or U11827 (N_11827,N_6671,N_9774);
or U11828 (N_11828,N_9370,N_6087);
and U11829 (N_11829,N_9229,N_9099);
or U11830 (N_11830,N_9590,N_7102);
xnor U11831 (N_11831,N_9078,N_6920);
nand U11832 (N_11832,N_8698,N_6582);
nand U11833 (N_11833,N_6095,N_6190);
and U11834 (N_11834,N_5936,N_9269);
or U11835 (N_11835,N_9239,N_7593);
and U11836 (N_11836,N_8958,N_8574);
nor U11837 (N_11837,N_8974,N_8111);
xor U11838 (N_11838,N_8027,N_5112);
xor U11839 (N_11839,N_7832,N_9478);
and U11840 (N_11840,N_5680,N_8867);
nand U11841 (N_11841,N_9020,N_6819);
and U11842 (N_11842,N_6250,N_9704);
and U11843 (N_11843,N_6474,N_8258);
nand U11844 (N_11844,N_7121,N_9765);
nor U11845 (N_11845,N_6606,N_9629);
and U11846 (N_11846,N_7272,N_7137);
or U11847 (N_11847,N_8597,N_7097);
xor U11848 (N_11848,N_9219,N_5320);
xor U11849 (N_11849,N_6644,N_8764);
or U11850 (N_11850,N_8487,N_5825);
nor U11851 (N_11851,N_7830,N_5069);
or U11852 (N_11852,N_9136,N_7151);
nand U11853 (N_11853,N_8009,N_8254);
xor U11854 (N_11854,N_7155,N_7686);
xor U11855 (N_11855,N_9934,N_8877);
nor U11856 (N_11856,N_7645,N_8103);
or U11857 (N_11857,N_9698,N_6852);
and U11858 (N_11858,N_7723,N_5709);
or U11859 (N_11859,N_6268,N_5537);
xnor U11860 (N_11860,N_5826,N_8706);
nor U11861 (N_11861,N_9368,N_6395);
nand U11862 (N_11862,N_5959,N_9597);
xor U11863 (N_11863,N_5974,N_7803);
or U11864 (N_11864,N_7259,N_9686);
xor U11865 (N_11865,N_7565,N_8933);
and U11866 (N_11866,N_5394,N_9319);
or U11867 (N_11867,N_5125,N_8804);
and U11868 (N_11868,N_9466,N_8352);
or U11869 (N_11869,N_9573,N_5331);
nor U11870 (N_11870,N_7902,N_7283);
nor U11871 (N_11871,N_8528,N_9911);
or U11872 (N_11872,N_7636,N_8620);
and U11873 (N_11873,N_8134,N_7813);
or U11874 (N_11874,N_9900,N_7153);
or U11875 (N_11875,N_5408,N_5847);
and U11876 (N_11876,N_7228,N_7972);
nor U11877 (N_11877,N_9880,N_6785);
nand U11878 (N_11878,N_8104,N_8781);
or U11879 (N_11879,N_6728,N_9120);
xnor U11880 (N_11880,N_8043,N_7599);
xnor U11881 (N_11881,N_8953,N_8047);
xor U11882 (N_11882,N_9566,N_5626);
or U11883 (N_11883,N_9457,N_6680);
and U11884 (N_11884,N_9681,N_6223);
nor U11885 (N_11885,N_7417,N_9177);
and U11886 (N_11886,N_8557,N_8876);
nor U11887 (N_11887,N_8074,N_9130);
or U11888 (N_11888,N_5165,N_5819);
nor U11889 (N_11889,N_6128,N_6743);
nand U11890 (N_11890,N_7168,N_9250);
xnor U11891 (N_11891,N_6677,N_8720);
and U11892 (N_11892,N_8555,N_7132);
xnor U11893 (N_11893,N_8519,N_5713);
nand U11894 (N_11894,N_6404,N_7564);
xor U11895 (N_11895,N_5668,N_6531);
xnor U11896 (N_11896,N_6552,N_5036);
or U11897 (N_11897,N_9199,N_6160);
nand U11898 (N_11898,N_6413,N_9890);
xor U11899 (N_11899,N_7904,N_7908);
xnor U11900 (N_11900,N_8160,N_5171);
or U11901 (N_11901,N_9766,N_6935);
nand U11902 (N_11902,N_9563,N_6226);
nor U11903 (N_11903,N_9906,N_9186);
xor U11904 (N_11904,N_6293,N_5765);
or U11905 (N_11905,N_7348,N_7519);
xor U11906 (N_11906,N_9233,N_9181);
xnor U11907 (N_11907,N_7746,N_7000);
and U11908 (N_11908,N_5244,N_8499);
and U11909 (N_11909,N_5498,N_5542);
nor U11910 (N_11910,N_7216,N_7572);
and U11911 (N_11911,N_8001,N_9214);
nand U11912 (N_11912,N_6426,N_5017);
xnor U11913 (N_11913,N_8267,N_5856);
nand U11914 (N_11914,N_9990,N_5310);
nor U11915 (N_11915,N_9633,N_6018);
and U11916 (N_11916,N_5557,N_9586);
xor U11917 (N_11917,N_5630,N_7580);
nand U11918 (N_11918,N_9179,N_5355);
nand U11919 (N_11919,N_9740,N_9280);
nand U11920 (N_11920,N_7681,N_7613);
nand U11921 (N_11921,N_7970,N_6461);
xor U11922 (N_11922,N_5547,N_5413);
xnor U11923 (N_11923,N_6244,N_5706);
and U11924 (N_11924,N_5366,N_8679);
nor U11925 (N_11925,N_7859,N_8216);
xor U11926 (N_11926,N_5022,N_5696);
nand U11927 (N_11927,N_5631,N_8512);
xor U11928 (N_11928,N_8381,N_7081);
nand U11929 (N_11929,N_5922,N_9596);
or U11930 (N_11930,N_5471,N_6308);
xnor U11931 (N_11931,N_6370,N_9933);
xnor U11932 (N_11932,N_8095,N_5978);
nand U11933 (N_11933,N_5351,N_5584);
and U11934 (N_11934,N_7627,N_7650);
and U11935 (N_11935,N_8366,N_5463);
nor U11936 (N_11936,N_7858,N_7869);
xor U11937 (N_11937,N_5635,N_7378);
xnor U11938 (N_11938,N_5107,N_8168);
and U11939 (N_11939,N_6523,N_7793);
xnor U11940 (N_11940,N_6225,N_6835);
and U11941 (N_11941,N_5694,N_7368);
nand U11942 (N_11942,N_5822,N_8041);
xor U11943 (N_11943,N_5942,N_6949);
or U11944 (N_11944,N_5062,N_7184);
xnor U11945 (N_11945,N_9879,N_8071);
or U11946 (N_11946,N_7086,N_5210);
nor U11947 (N_11947,N_6721,N_7464);
and U11948 (N_11948,N_9546,N_6061);
xor U11949 (N_11949,N_7056,N_5158);
xor U11950 (N_11950,N_8435,N_5885);
nor U11951 (N_11951,N_8899,N_9375);
and U11952 (N_11952,N_6525,N_9781);
nand U11953 (N_11953,N_5560,N_9662);
or U11954 (N_11954,N_7935,N_9275);
or U11955 (N_11955,N_8468,N_9156);
nand U11956 (N_11956,N_8949,N_8212);
xnor U11957 (N_11957,N_6076,N_9300);
nand U11958 (N_11958,N_9282,N_5473);
or U11959 (N_11959,N_7499,N_7280);
nand U11960 (N_11960,N_9831,N_6258);
and U11961 (N_11961,N_5356,N_8034);
and U11962 (N_11962,N_5042,N_9040);
xor U11963 (N_11963,N_5581,N_8735);
and U11964 (N_11964,N_8968,N_7202);
and U11965 (N_11965,N_9930,N_5596);
and U11966 (N_11966,N_5342,N_5933);
and U11967 (N_11967,N_7459,N_9301);
and U11968 (N_11968,N_5518,N_5624);
nand U11969 (N_11969,N_7342,N_5556);
xor U11970 (N_11970,N_6912,N_6104);
or U11971 (N_11971,N_5410,N_8197);
nor U11972 (N_11972,N_8372,N_6384);
xnor U11973 (N_11973,N_6069,N_5774);
xor U11974 (N_11974,N_7937,N_8059);
and U11975 (N_11975,N_7211,N_9734);
or U11976 (N_11976,N_6672,N_6975);
and U11977 (N_11977,N_9872,N_5122);
nor U11978 (N_11978,N_8136,N_8821);
xor U11979 (N_11979,N_6429,N_9190);
nand U11980 (N_11980,N_8259,N_7438);
nor U11981 (N_11981,N_5243,N_7340);
xnor U11982 (N_11982,N_8850,N_9107);
nand U11983 (N_11983,N_5999,N_5261);
nand U11984 (N_11984,N_7135,N_5991);
or U11985 (N_11985,N_6176,N_5269);
nand U11986 (N_11986,N_6725,N_7411);
or U11987 (N_11987,N_9840,N_7991);
nor U11988 (N_11988,N_5727,N_9967);
xnor U11989 (N_11989,N_7009,N_9469);
nand U11990 (N_11990,N_8196,N_8917);
or U11991 (N_11991,N_7050,N_7760);
nor U11992 (N_11992,N_6917,N_9689);
xnor U11993 (N_11993,N_6930,N_8520);
and U11994 (N_11994,N_7707,N_7250);
or U11995 (N_11995,N_9703,N_6150);
or U11996 (N_11996,N_7028,N_6567);
nor U11997 (N_11997,N_8774,N_7825);
or U11998 (N_11998,N_8691,N_6648);
xnor U11999 (N_11999,N_8971,N_5954);
nor U12000 (N_12000,N_6720,N_5673);
xnor U12001 (N_12001,N_8415,N_8056);
or U12002 (N_12002,N_9749,N_9088);
or U12003 (N_12003,N_5209,N_8641);
and U12004 (N_12004,N_5731,N_5259);
nand U12005 (N_12005,N_7189,N_7863);
nand U12006 (N_12006,N_8241,N_9222);
xor U12007 (N_12007,N_8925,N_6236);
or U12008 (N_12008,N_5208,N_5674);
xor U12009 (N_12009,N_7989,N_7868);
xor U12010 (N_12010,N_6127,N_7966);
xnor U12011 (N_12011,N_6545,N_8341);
nand U12012 (N_12012,N_9773,N_5488);
nand U12013 (N_12013,N_5747,N_7622);
nor U12014 (N_12014,N_9100,N_7644);
and U12015 (N_12015,N_7222,N_8610);
nand U12016 (N_12016,N_8046,N_9524);
nor U12017 (N_12017,N_7442,N_6505);
or U12018 (N_12018,N_7233,N_7319);
nor U12019 (N_12019,N_6691,N_7900);
xor U12020 (N_12020,N_8973,N_9580);
nor U12021 (N_12021,N_9223,N_5457);
nand U12022 (N_12022,N_7252,N_9187);
or U12023 (N_12023,N_8332,N_5871);
and U12024 (N_12024,N_5157,N_9898);
and U12025 (N_12025,N_6090,N_5671);
xor U12026 (N_12026,N_6263,N_9627);
and U12027 (N_12027,N_8218,N_9442);
or U12028 (N_12028,N_8798,N_9082);
nand U12029 (N_12029,N_5866,N_6616);
nand U12030 (N_12030,N_7180,N_6101);
xor U12031 (N_12031,N_9973,N_7505);
nand U12032 (N_12032,N_9935,N_7532);
nor U12033 (N_12033,N_8072,N_7771);
and U12034 (N_12034,N_9249,N_6670);
and U12035 (N_12035,N_5297,N_6415);
and U12036 (N_12036,N_7615,N_5775);
nor U12037 (N_12037,N_6041,N_8621);
nor U12038 (N_12038,N_6739,N_9210);
xor U12039 (N_12039,N_6108,N_9064);
or U12040 (N_12040,N_7481,N_9894);
xnor U12041 (N_12041,N_7751,N_8616);
nand U12042 (N_12042,N_7234,N_5417);
and U12043 (N_12043,N_9026,N_6385);
and U12044 (N_12044,N_6168,N_7244);
and U12045 (N_12045,N_5971,N_6408);
xor U12046 (N_12046,N_9529,N_6378);
or U12047 (N_12047,N_5006,N_6070);
xor U12048 (N_12048,N_8373,N_8633);
xnor U12049 (N_12049,N_9062,N_9420);
or U12050 (N_12050,N_5442,N_8210);
and U12051 (N_12051,N_9723,N_5807);
nor U12052 (N_12052,N_8978,N_9693);
and U12053 (N_12053,N_5564,N_8429);
or U12054 (N_12054,N_5026,N_9844);
nor U12055 (N_12055,N_7478,N_5533);
and U12056 (N_12056,N_5056,N_9640);
or U12057 (N_12057,N_8426,N_8547);
nand U12058 (N_12058,N_8763,N_9281);
nor U12059 (N_12059,N_8396,N_5343);
xor U12060 (N_12060,N_7326,N_5995);
xnor U12061 (N_12061,N_6274,N_9441);
or U12062 (N_12062,N_9603,N_7999);
or U12063 (N_12063,N_7131,N_9227);
xor U12064 (N_12064,N_6717,N_7307);
and U12065 (N_12065,N_8238,N_5395);
or U12066 (N_12066,N_7324,N_8892);
nor U12067 (N_12067,N_8344,N_5539);
or U12068 (N_12068,N_9435,N_5715);
or U12069 (N_12069,N_5459,N_7878);
nand U12070 (N_12070,N_5429,N_7177);
nand U12071 (N_12071,N_9143,N_8553);
nor U12072 (N_12072,N_8414,N_5993);
or U12073 (N_12073,N_5155,N_8115);
and U12074 (N_12074,N_8287,N_5850);
nand U12075 (N_12075,N_9376,N_9904);
xor U12076 (N_12076,N_9882,N_6137);
nand U12077 (N_12077,N_8065,N_8600);
nand U12078 (N_12078,N_7920,N_7678);
and U12079 (N_12079,N_6729,N_8990);
nand U12080 (N_12080,N_8330,N_5622);
and U12081 (N_12081,N_8852,N_8008);
nor U12082 (N_12082,N_6558,N_9759);
nand U12083 (N_12083,N_8139,N_5283);
nand U12084 (N_12084,N_7828,N_7750);
or U12085 (N_12085,N_7817,N_7285);
nor U12086 (N_12086,N_9946,N_7490);
and U12087 (N_12087,N_8465,N_8649);
or U12088 (N_12088,N_9965,N_9438);
and U12089 (N_12089,N_8669,N_5916);
nand U12090 (N_12090,N_7641,N_7282);
xor U12091 (N_12091,N_8409,N_5676);
nand U12092 (N_12092,N_7575,N_7781);
or U12093 (N_12093,N_5845,N_9387);
and U12094 (N_12094,N_6313,N_8754);
nor U12095 (N_12095,N_9995,N_5029);
nand U12096 (N_12096,N_7667,N_9339);
xor U12097 (N_12097,N_8251,N_9613);
or U12098 (N_12098,N_9241,N_9708);
xnor U12099 (N_12099,N_7419,N_6597);
and U12100 (N_12100,N_5848,N_6952);
nand U12101 (N_12101,N_9535,N_8107);
nand U12102 (N_12102,N_7224,N_6401);
and U12103 (N_12103,N_5956,N_6536);
and U12104 (N_12104,N_7585,N_5053);
nor U12105 (N_12105,N_5704,N_9270);
or U12106 (N_12106,N_9507,N_8314);
or U12107 (N_12107,N_5219,N_8869);
nor U12108 (N_12108,N_6840,N_5329);
and U12109 (N_12109,N_8119,N_6447);
and U12110 (N_12110,N_8951,N_8660);
nand U12111 (N_12111,N_8533,N_9767);
xnor U12112 (N_12112,N_8758,N_9570);
or U12113 (N_12113,N_5440,N_5167);
nand U12114 (N_12114,N_8999,N_8321);
and U12115 (N_12115,N_5450,N_5404);
nor U12116 (N_12116,N_9593,N_8291);
nand U12117 (N_12117,N_7597,N_7973);
xnor U12118 (N_12118,N_6929,N_6669);
nor U12119 (N_12119,N_9402,N_7004);
or U12120 (N_12120,N_8693,N_6245);
nand U12121 (N_12121,N_6841,N_5130);
nor U12122 (N_12122,N_9323,N_6086);
xnor U12123 (N_12123,N_5881,N_8472);
xnor U12124 (N_12124,N_8058,N_9043);
nor U12125 (N_12125,N_9132,N_5738);
and U12126 (N_12126,N_7487,N_8674);
or U12127 (N_12127,N_8005,N_6005);
xnor U12128 (N_12128,N_9790,N_8818);
and U12129 (N_12129,N_6657,N_7143);
nor U12130 (N_12130,N_8783,N_9348);
nor U12131 (N_12131,N_7640,N_7310);
nand U12132 (N_12132,N_7494,N_6237);
or U12133 (N_12133,N_7323,N_7471);
nand U12134 (N_12134,N_6142,N_6062);
or U12135 (N_12135,N_8618,N_9265);
nor U12136 (N_12136,N_9292,N_5191);
xnor U12137 (N_12137,N_8143,N_8356);
and U12138 (N_12138,N_8522,N_9624);
nor U12139 (N_12139,N_5135,N_6210);
nor U12140 (N_12140,N_6838,N_6799);
or U12141 (N_12141,N_9069,N_7737);
or U12142 (N_12142,N_9843,N_6911);
xnor U12143 (N_12143,N_5652,N_7437);
or U12144 (N_12144,N_7243,N_5677);
or U12145 (N_12145,N_5524,N_5617);
xnor U12146 (N_12146,N_5679,N_8537);
nand U12147 (N_12147,N_5672,N_7560);
xor U12148 (N_12148,N_8637,N_8369);
or U12149 (N_12149,N_7103,N_5010);
and U12150 (N_12150,N_7739,N_6724);
xnor U12151 (N_12151,N_6769,N_9639);
and U12152 (N_12152,N_9972,N_9993);
xnor U12153 (N_12153,N_8302,N_9358);
nor U12154 (N_12154,N_8542,N_9788);
and U12155 (N_12155,N_5614,N_6060);
and U12156 (N_12156,N_8786,N_7208);
nand U12157 (N_12157,N_5817,N_6065);
xor U12158 (N_12158,N_7942,N_8108);
xnor U12159 (N_12159,N_7673,N_8049);
nand U12160 (N_12160,N_9353,N_5447);
or U12161 (N_12161,N_9710,N_7874);
nor U12162 (N_12162,N_8016,N_9455);
or U12163 (N_12163,N_8615,N_7145);
nor U12164 (N_12164,N_9672,N_9963);
xnor U12165 (N_12165,N_6446,N_9730);
nor U12166 (N_12166,N_8806,N_5736);
nand U12167 (N_12167,N_7117,N_9600);
or U12168 (N_12168,N_6688,N_5839);
nand U12169 (N_12169,N_5691,N_9388);
xnor U12170 (N_12170,N_7852,N_7227);
or U12171 (N_12171,N_8585,N_6985);
nor U12172 (N_12172,N_7993,N_8187);
or U12173 (N_12173,N_5475,N_7418);
and U12174 (N_12174,N_9964,N_8177);
nand U12175 (N_12175,N_8135,N_6563);
nor U12176 (N_12176,N_9912,N_6854);
or U12177 (N_12177,N_8998,N_5769);
and U12178 (N_12178,N_7679,N_6184);
or U12179 (N_12179,N_9359,N_6732);
or U12180 (N_12180,N_9999,N_5349);
xnor U12181 (N_12181,N_8881,N_9658);
nor U12182 (N_12182,N_7458,N_5981);
nand U12183 (N_12183,N_7367,N_7297);
nand U12184 (N_12184,N_9321,N_7761);
and U12185 (N_12185,N_9735,N_7839);
nor U12186 (N_12186,N_6832,N_8278);
and U12187 (N_12187,N_9024,N_9630);
and U12188 (N_12188,N_5262,N_9988);
and U12189 (N_12189,N_9691,N_9050);
or U12190 (N_12190,N_6681,N_9678);
nand U12191 (N_12191,N_5705,N_5800);
nand U12192 (N_12192,N_7300,N_9464);
and U12193 (N_12193,N_5341,N_6592);
xor U12194 (N_12194,N_6437,N_5323);
nand U12195 (N_12195,N_6973,N_5330);
nor U12196 (N_12196,N_8671,N_7430);
nor U12197 (N_12197,N_7784,N_7098);
xnor U12198 (N_12198,N_6737,N_5600);
and U12199 (N_12199,N_6355,N_7571);
nand U12200 (N_12200,N_5077,N_9667);
nand U12201 (N_12201,N_8760,N_6196);
and U12202 (N_12202,N_7632,N_7060);
or U12203 (N_12203,N_7726,N_8172);
and U12204 (N_12204,N_5448,N_5255);
or U12205 (N_12205,N_7710,N_7078);
xnor U12206 (N_12206,N_8924,N_8964);
xnor U12207 (N_12207,N_6667,N_8831);
nand U12208 (N_12208,N_9671,N_9513);
nor U12209 (N_12209,N_7897,N_8920);
and U12210 (N_12210,N_7578,N_6421);
and U12211 (N_12211,N_7027,N_5530);
xor U12212 (N_12212,N_7986,N_6950);
nand U12213 (N_12213,N_6987,N_7138);
nand U12214 (N_12214,N_5152,N_5318);
nor U12215 (N_12215,N_6510,N_5117);
nand U12216 (N_12216,N_7694,N_9571);
nor U12217 (N_12217,N_8623,N_8145);
nor U12218 (N_12218,N_6471,N_7444);
nand U12219 (N_12219,N_8061,N_7617);
xor U12220 (N_12220,N_8634,N_6809);
xor U12221 (N_12221,N_9516,N_6976);
xnor U12222 (N_12222,N_6807,N_7034);
xnor U12223 (N_12223,N_5952,N_5915);
nor U12224 (N_12224,N_9777,N_6371);
xnor U12225 (N_12225,N_6532,N_5304);
and U12226 (N_12226,N_6255,N_6937);
or U12227 (N_12227,N_8443,N_9651);
or U12228 (N_12228,N_9437,N_9826);
nor U12229 (N_12229,N_7390,N_9701);
nor U12230 (N_12230,N_7128,N_9511);
xor U12231 (N_12231,N_7156,N_6928);
nand U12232 (N_12232,N_7543,N_6522);
nand U12233 (N_12233,N_7776,N_6002);
xnor U12234 (N_12234,N_6977,N_5700);
nand U12235 (N_12235,N_5550,N_8284);
nand U12236 (N_12236,N_7341,N_9520);
nand U12237 (N_12237,N_9929,N_8604);
nand U12238 (N_12238,N_5828,N_9163);
xor U12239 (N_12239,N_7791,N_8112);
and U12240 (N_12240,N_8683,N_7147);
nor U12241 (N_12241,N_5007,N_9506);
nor U12242 (N_12242,N_9467,N_6148);
nor U12243 (N_12243,N_9106,N_6020);
xnor U12244 (N_12244,N_7819,N_6572);
or U12245 (N_12245,N_5653,N_9444);
nor U12246 (N_12246,N_7030,N_8493);
nor U12247 (N_12247,N_9303,N_5313);
nor U12248 (N_12248,N_8494,N_5460);
nor U12249 (N_12249,N_8054,N_6402);
nand U12250 (N_12250,N_6266,N_6220);
and U12251 (N_12251,N_7716,N_6509);
nand U12252 (N_12252,N_6043,N_6073);
xor U12253 (N_12253,N_8739,N_7245);
nor U12254 (N_12254,N_9523,N_7533);
and U12255 (N_12255,N_7328,N_7043);
and U12256 (N_12256,N_9105,N_5098);
nand U12257 (N_12257,N_5308,N_7251);
nor U12258 (N_12258,N_7422,N_6252);
xor U12259 (N_12259,N_6019,N_6439);
and U12260 (N_12260,N_6063,N_9901);
and U12261 (N_12261,N_8025,N_8801);
and U12262 (N_12262,N_7577,N_8856);
or U12263 (N_12263,N_7094,N_7040);
nor U12264 (N_12264,N_7950,N_8832);
or U12265 (N_12265,N_7386,N_6283);
nand U12266 (N_12266,N_6594,N_7033);
and U12267 (N_12267,N_8741,N_5627);
nand U12268 (N_12268,N_6814,N_7407);
or U12269 (N_12269,N_5771,N_7596);
and U12270 (N_12270,N_6703,N_7357);
xor U12271 (N_12271,N_7370,N_8686);
xnor U12272 (N_12272,N_7394,N_9848);
xnor U12273 (N_12273,N_5215,N_5487);
or U12274 (N_12274,N_8865,N_5654);
and U12275 (N_12275,N_7648,N_5689);
and U12276 (N_12276,N_9525,N_6713);
nand U12277 (N_12277,N_7266,N_6094);
or U12278 (N_12278,N_6194,N_6464);
or U12279 (N_12279,N_9665,N_5303);
nor U12280 (N_12280,N_8530,N_5383);
nor U12281 (N_12281,N_5247,N_7969);
xor U12282 (N_12282,N_9279,N_6238);
nand U12283 (N_12283,N_5496,N_8590);
or U12284 (N_12284,N_9752,N_8363);
nor U12285 (N_12285,N_7415,N_8288);
or U12286 (N_12286,N_5060,N_6587);
xor U12287 (N_12287,N_7017,N_8575);
nor U12288 (N_12288,N_5005,N_7912);
xor U12289 (N_12289,N_9168,N_5346);
nand U12290 (N_12290,N_6599,N_5570);
nand U12291 (N_12291,N_7827,N_9052);
nand U12292 (N_12292,N_8898,N_5088);
nand U12293 (N_12293,N_7104,N_6389);
and U12294 (N_12294,N_5811,N_7452);
and U12295 (N_12295,N_7512,N_6338);
xnor U12296 (N_12296,N_6588,N_6232);
and U12297 (N_12297,N_9980,N_9863);
or U12298 (N_12298,N_8718,N_9463);
and U12299 (N_12299,N_7790,N_8586);
or U12300 (N_12300,N_9332,N_8408);
nand U12301 (N_12301,N_8488,N_7463);
and U12302 (N_12302,N_5900,N_7205);
and U12303 (N_12303,N_8817,N_9073);
nand U12304 (N_12304,N_8886,N_9556);
xor U12305 (N_12305,N_9864,N_7335);
and U12306 (N_12306,N_5438,N_7894);
xor U12307 (N_12307,N_8401,N_9362);
or U12308 (N_12308,N_6678,N_5824);
nor U12309 (N_12309,N_7965,N_8756);
xnor U12310 (N_12310,N_8023,N_6773);
nor U12311 (N_12311,N_9398,N_6066);
nor U12312 (N_12312,N_9876,N_7194);
and U12313 (N_12313,N_9377,N_9439);
or U12314 (N_12314,N_6038,N_7721);
xor U12315 (N_12315,N_5519,N_9032);
nor U12316 (N_12316,N_7598,N_5946);
nand U12317 (N_12317,N_6921,N_6999);
and U12318 (N_12318,N_9808,N_5472);
nand U12319 (N_12319,N_9925,N_6042);
and U12320 (N_12320,N_6277,N_5111);
nor U12321 (N_12321,N_5044,N_6507);
and U12322 (N_12322,N_8987,N_7856);
or U12323 (N_12323,N_6243,N_5783);
nand U12324 (N_12324,N_7756,N_6275);
xor U12325 (N_12325,N_6451,N_8536);
nand U12326 (N_12326,N_6692,N_7059);
and U12327 (N_12327,N_8928,N_8096);
xor U12328 (N_12328,N_9328,N_9293);
nand U12329 (N_12329,N_9285,N_5908);
xor U12330 (N_12330,N_9330,N_5225);
or U12331 (N_12331,N_9920,N_5139);
xor U12332 (N_12332,N_6173,N_5070);
nor U12333 (N_12333,N_5256,N_5458);
or U12334 (N_12334,N_7029,N_5441);
and U12335 (N_12335,N_5692,N_9033);
nor U12336 (N_12336,N_6369,N_8650);
or U12337 (N_12337,N_6500,N_5478);
xnor U12338 (N_12338,N_8989,N_5798);
nand U12339 (N_12339,N_6291,N_9360);
nor U12340 (N_12340,N_6764,N_7916);
nand U12341 (N_12341,N_9314,N_8830);
xnor U12342 (N_12342,N_9245,N_5816);
nor U12343 (N_12343,N_6629,N_6804);
nor U12344 (N_12344,N_6760,N_5527);
nor U12345 (N_12345,N_8897,N_5235);
or U12346 (N_12346,N_7012,N_8167);
xor U12347 (N_12347,N_6602,N_9923);
or U12348 (N_12348,N_5230,N_9635);
or U12349 (N_12349,N_8717,N_8416);
nand U12350 (N_12350,N_5795,N_8980);
xnor U12351 (N_12351,N_7740,N_8234);
nor U12352 (N_12352,N_7066,N_6969);
or U12353 (N_12353,N_6520,N_9384);
xor U12354 (N_12354,N_7162,N_6611);
nand U12355 (N_12355,N_7021,N_9436);
nand U12356 (N_12356,N_7402,N_5609);
nor U12357 (N_12357,N_7779,N_5385);
xnor U12358 (N_12358,N_6993,N_7063);
or U12359 (N_12359,N_6719,N_9322);
nand U12360 (N_12360,N_7473,N_5721);
and U12361 (N_12361,N_5628,N_7727);
and U12362 (N_12362,N_8622,N_6449);
nor U12363 (N_12363,N_8750,N_6967);
nand U12364 (N_12364,N_9411,N_6045);
nor U12365 (N_12365,N_8224,N_5603);
and U12366 (N_12366,N_9812,N_6314);
and U12367 (N_12367,N_6548,N_7876);
nor U12368 (N_12368,N_7663,N_9277);
and U12369 (N_12369,N_8362,N_9255);
nor U12370 (N_12370,N_7269,N_6690);
nor U12371 (N_12371,N_9758,N_5931);
and U12372 (N_12372,N_7711,N_7036);
xor U12373 (N_12373,N_8769,N_9382);
xor U12374 (N_12374,N_7267,N_7922);
and U12375 (N_12375,N_5804,N_7668);
and U12376 (N_12376,N_9856,N_8425);
or U12377 (N_12377,N_9521,N_8052);
nor U12378 (N_12378,N_7985,N_9254);
or U12379 (N_12379,N_5091,N_9589);
nor U12380 (N_12380,N_5579,N_8690);
nand U12381 (N_12381,N_9936,N_5018);
nand U12382 (N_12382,N_6980,N_9476);
nor U12383 (N_12383,N_8943,N_9859);
nor U12384 (N_12384,N_8589,N_9391);
xor U12385 (N_12385,N_9007,N_7384);
or U12386 (N_12386,N_8444,N_7717);
nand U12387 (N_12387,N_5296,N_7703);
or U12388 (N_12388,N_9415,N_5202);
and U12389 (N_12389,N_7510,N_8884);
xor U12390 (N_12390,N_5543,N_9203);
xor U12391 (N_12391,N_7318,N_5444);
xnor U12392 (N_12392,N_7052,N_6888);
or U12393 (N_12393,N_8419,N_7546);
and U12394 (N_12394,N_5270,N_6103);
xor U12395 (N_12395,N_8360,N_7261);
and U12396 (N_12396,N_7101,N_8915);
xor U12397 (N_12397,N_7872,N_6844);
and U12398 (N_12398,N_9002,N_7690);
xnor U12399 (N_12399,N_5049,N_6213);
xor U12400 (N_12400,N_7242,N_8936);
and U12401 (N_12401,N_9167,N_9591);
or U12402 (N_12402,N_6055,N_9256);
or U12403 (N_12403,N_8722,N_5418);
nand U12404 (N_12404,N_7845,N_8724);
xnor U12405 (N_12405,N_5199,N_6445);
and U12406 (N_12406,N_9448,N_6981);
nor U12407 (N_12407,N_5021,N_5099);
and U12408 (N_12408,N_9821,N_8954);
xor U12409 (N_12409,N_8606,N_6300);
and U12410 (N_12410,N_5896,N_5743);
or U12411 (N_12411,N_6348,N_7193);
or U12412 (N_12412,N_6961,N_6145);
nor U12413 (N_12413,N_5735,N_5840);
or U12414 (N_12414,N_6262,N_7239);
and U12415 (N_12415,N_9924,N_6537);
and U12416 (N_12416,N_6393,N_7484);
nor U12417 (N_12417,N_8730,N_8249);
nand U12418 (N_12418,N_6406,N_6868);
and U12419 (N_12419,N_6296,N_6383);
nor U12420 (N_12420,N_8716,N_8176);
nand U12421 (N_12421,N_5514,N_8237);
and U12422 (N_12422,N_8887,N_8692);
xor U12423 (N_12423,N_6649,N_9729);
or U12424 (N_12424,N_9072,N_7949);
nor U12425 (N_12425,N_6826,N_5046);
xor U12426 (N_12426,N_5785,N_9862);
xnor U12427 (N_12427,N_7099,N_9194);
nand U12428 (N_12428,N_6098,N_8194);
xnor U12429 (N_12429,N_5553,N_5309);
or U12430 (N_12430,N_9554,N_8402);
xor U12431 (N_12431,N_5969,N_7976);
and U12432 (N_12432,N_8554,N_7397);
nor U12433 (N_12433,N_6601,N_5372);
nor U12434 (N_12434,N_7313,N_6387);
xnor U12435 (N_12435,N_6579,N_8120);
nand U12436 (N_12436,N_5226,N_9240);
xnor U12437 (N_12437,N_8531,N_5387);
xnor U12438 (N_12438,N_6201,N_6941);
xnor U12439 (N_12439,N_8301,N_6699);
or U12440 (N_12440,N_6174,N_9412);
or U12441 (N_12441,N_9488,N_5025);
nand U12442 (N_12442,N_7829,N_7941);
nor U12443 (N_12443,N_6368,N_7401);
or U12444 (N_12444,N_9059,N_9602);
nor U12445 (N_12445,N_9465,N_7144);
or U12446 (N_12446,N_8042,N_7399);
nor U12447 (N_12447,N_6850,N_5852);
or U12448 (N_12448,N_8319,N_5569);
nor U12449 (N_12449,N_7440,N_5895);
or U12450 (N_12450,N_6416,N_6206);
or U12451 (N_12451,N_9960,N_6919);
nand U12452 (N_12452,N_8624,N_5290);
xor U12453 (N_12453,N_8094,N_7735);
nor U12454 (N_12454,N_7983,N_5114);
nand U12455 (N_12455,N_8279,N_8121);
xnor U12456 (N_12456,N_7392,N_7888);
and U12457 (N_12457,N_8417,N_8260);
or U12458 (N_12458,N_6169,N_7201);
or U12459 (N_12459,N_5316,N_6600);
and U12460 (N_12460,N_5616,N_6884);
and U12461 (N_12461,N_8132,N_6834);
or U12462 (N_12462,N_5508,N_7352);
or U12463 (N_12463,N_6613,N_5144);
and U12464 (N_12464,N_8658,N_8851);
nor U12465 (N_12465,N_9491,N_5362);
xnor U12466 (N_12466,N_6470,N_5425);
or U12467 (N_12467,N_6619,N_9310);
nor U12468 (N_12468,N_9907,N_9312);
nor U12469 (N_12469,N_7257,N_7977);
or U12470 (N_12470,N_8217,N_6786);
or U12471 (N_12471,N_5223,N_9680);
and U12472 (N_12472,N_8473,N_9095);
xor U12473 (N_12473,N_9646,N_8391);
and U12474 (N_12474,N_6794,N_9318);
xnor U12475 (N_12475,N_5401,N_6538);
xnor U12476 (N_12476,N_9173,N_7582);
nand U12477 (N_12477,N_9873,N_6762);
xor U12478 (N_12478,N_9432,N_9013);
nand U12479 (N_12479,N_6633,N_8060);
or U12480 (N_12480,N_9841,N_5874);
nor U12481 (N_12481,N_8109,N_6306);
nand U12482 (N_12482,N_8645,N_8815);
and U12483 (N_12483,N_9133,N_8808);
and U12484 (N_12484,N_5763,N_9584);
nor U12485 (N_12485,N_9053,N_9793);
and U12486 (N_12486,N_5166,N_5893);
nand U12487 (N_12487,N_7877,N_8994);
nand U12488 (N_12488,N_5104,N_7046);
nor U12489 (N_12489,N_5970,N_5955);
and U12490 (N_12490,N_9653,N_8206);
nor U12491 (N_12491,N_9779,N_5940);
nand U12492 (N_12492,N_7944,N_7708);
xnor U12493 (N_12493,N_9543,N_9354);
and U12494 (N_12494,N_6542,N_8087);
xnor U12495 (N_12495,N_9645,N_5998);
nor U12496 (N_12496,N_5748,N_7573);
and U12497 (N_12497,N_8471,N_5910);
nor U12498 (N_12498,N_5831,N_6440);
nor U12499 (N_12499,N_9244,N_6872);
and U12500 (N_12500,N_6427,N_9676);
and U12501 (N_12501,N_9236,N_9570);
or U12502 (N_12502,N_7504,N_7091);
or U12503 (N_12503,N_6042,N_8401);
nand U12504 (N_12504,N_8532,N_7140);
nor U12505 (N_12505,N_8434,N_5844);
or U12506 (N_12506,N_9296,N_6711);
and U12507 (N_12507,N_6759,N_9970);
or U12508 (N_12508,N_7624,N_8595);
xnor U12509 (N_12509,N_9483,N_8554);
nand U12510 (N_12510,N_9600,N_7872);
nand U12511 (N_12511,N_8386,N_8957);
nand U12512 (N_12512,N_6886,N_6225);
nand U12513 (N_12513,N_9180,N_9261);
and U12514 (N_12514,N_9172,N_7761);
and U12515 (N_12515,N_6830,N_7954);
and U12516 (N_12516,N_5707,N_5923);
or U12517 (N_12517,N_9962,N_5114);
nor U12518 (N_12518,N_5608,N_5707);
or U12519 (N_12519,N_9848,N_9007);
nor U12520 (N_12520,N_6364,N_6354);
nand U12521 (N_12521,N_7419,N_9607);
or U12522 (N_12522,N_5595,N_5644);
nand U12523 (N_12523,N_5481,N_6003);
and U12524 (N_12524,N_5266,N_7100);
nand U12525 (N_12525,N_9014,N_6541);
nand U12526 (N_12526,N_6124,N_5445);
and U12527 (N_12527,N_7570,N_6068);
nor U12528 (N_12528,N_6420,N_6432);
nor U12529 (N_12529,N_8935,N_9818);
nand U12530 (N_12530,N_6825,N_8600);
nand U12531 (N_12531,N_5439,N_6627);
xor U12532 (N_12532,N_9697,N_7839);
xnor U12533 (N_12533,N_8883,N_6056);
nand U12534 (N_12534,N_5268,N_5759);
nand U12535 (N_12535,N_5680,N_5499);
xor U12536 (N_12536,N_9037,N_6656);
nand U12537 (N_12537,N_7703,N_5572);
and U12538 (N_12538,N_6463,N_5045);
and U12539 (N_12539,N_7295,N_5931);
nor U12540 (N_12540,N_7943,N_8362);
nand U12541 (N_12541,N_8049,N_8437);
and U12542 (N_12542,N_5046,N_5019);
or U12543 (N_12543,N_8358,N_6048);
nand U12544 (N_12544,N_6957,N_5787);
xnor U12545 (N_12545,N_8116,N_6934);
or U12546 (N_12546,N_5799,N_9371);
nand U12547 (N_12547,N_7613,N_7596);
xnor U12548 (N_12548,N_6267,N_7758);
and U12549 (N_12549,N_7037,N_8336);
nand U12550 (N_12550,N_9093,N_5302);
nor U12551 (N_12551,N_8205,N_5976);
nand U12552 (N_12552,N_5253,N_9017);
or U12553 (N_12553,N_6517,N_7223);
and U12554 (N_12554,N_7047,N_7915);
or U12555 (N_12555,N_6262,N_6250);
xnor U12556 (N_12556,N_7855,N_7695);
nor U12557 (N_12557,N_5504,N_8589);
and U12558 (N_12558,N_7764,N_5495);
nand U12559 (N_12559,N_5495,N_8516);
nand U12560 (N_12560,N_8433,N_5669);
nand U12561 (N_12561,N_9404,N_5645);
and U12562 (N_12562,N_8033,N_9828);
nor U12563 (N_12563,N_5372,N_7087);
xor U12564 (N_12564,N_7773,N_7880);
xor U12565 (N_12565,N_9713,N_9200);
nor U12566 (N_12566,N_5517,N_9740);
or U12567 (N_12567,N_7577,N_9729);
nor U12568 (N_12568,N_5568,N_9274);
nand U12569 (N_12569,N_7183,N_5035);
nor U12570 (N_12570,N_8411,N_6512);
xnor U12571 (N_12571,N_7273,N_5548);
or U12572 (N_12572,N_5848,N_8761);
or U12573 (N_12573,N_9964,N_8397);
nand U12574 (N_12574,N_8743,N_9883);
or U12575 (N_12575,N_8384,N_7693);
nor U12576 (N_12576,N_6946,N_8409);
or U12577 (N_12577,N_7301,N_7356);
nand U12578 (N_12578,N_5556,N_6415);
nand U12579 (N_12579,N_7108,N_5862);
or U12580 (N_12580,N_9299,N_5780);
nor U12581 (N_12581,N_8531,N_6549);
or U12582 (N_12582,N_8590,N_5189);
xor U12583 (N_12583,N_5242,N_9776);
nand U12584 (N_12584,N_7830,N_5878);
xor U12585 (N_12585,N_9521,N_6953);
nand U12586 (N_12586,N_8504,N_7657);
xnor U12587 (N_12587,N_9080,N_5617);
and U12588 (N_12588,N_5951,N_8837);
or U12589 (N_12589,N_8479,N_8069);
nor U12590 (N_12590,N_5497,N_8865);
nor U12591 (N_12591,N_5988,N_9977);
xor U12592 (N_12592,N_8744,N_5912);
or U12593 (N_12593,N_5094,N_6076);
nor U12594 (N_12594,N_9102,N_9769);
and U12595 (N_12595,N_9500,N_8240);
and U12596 (N_12596,N_5493,N_8919);
and U12597 (N_12597,N_8094,N_8872);
or U12598 (N_12598,N_8620,N_6653);
xnor U12599 (N_12599,N_8730,N_5651);
and U12600 (N_12600,N_8007,N_9507);
or U12601 (N_12601,N_9103,N_6947);
nor U12602 (N_12602,N_9071,N_8248);
or U12603 (N_12603,N_5118,N_7848);
nand U12604 (N_12604,N_5205,N_8997);
and U12605 (N_12605,N_8653,N_5029);
xnor U12606 (N_12606,N_8563,N_7086);
xor U12607 (N_12607,N_9687,N_9292);
xor U12608 (N_12608,N_9672,N_8899);
nor U12609 (N_12609,N_7086,N_6824);
xnor U12610 (N_12610,N_8252,N_6956);
xnor U12611 (N_12611,N_5012,N_9072);
nand U12612 (N_12612,N_5013,N_7415);
nor U12613 (N_12613,N_6862,N_5028);
or U12614 (N_12614,N_7163,N_7775);
or U12615 (N_12615,N_6314,N_5846);
xor U12616 (N_12616,N_7597,N_8651);
nand U12617 (N_12617,N_5522,N_7112);
xor U12618 (N_12618,N_7491,N_6263);
nor U12619 (N_12619,N_8662,N_9408);
nand U12620 (N_12620,N_8102,N_6731);
nand U12621 (N_12621,N_5746,N_6486);
and U12622 (N_12622,N_8588,N_7281);
and U12623 (N_12623,N_6429,N_7262);
or U12624 (N_12624,N_5501,N_5968);
xor U12625 (N_12625,N_5446,N_6929);
nand U12626 (N_12626,N_5758,N_6075);
and U12627 (N_12627,N_5519,N_7340);
and U12628 (N_12628,N_5867,N_6702);
and U12629 (N_12629,N_7290,N_6907);
and U12630 (N_12630,N_7007,N_7137);
and U12631 (N_12631,N_6453,N_5498);
nor U12632 (N_12632,N_9870,N_9701);
or U12633 (N_12633,N_9989,N_5630);
xor U12634 (N_12634,N_9542,N_5929);
or U12635 (N_12635,N_5392,N_7643);
and U12636 (N_12636,N_5352,N_8354);
xor U12637 (N_12637,N_9602,N_8090);
nand U12638 (N_12638,N_7629,N_6377);
nor U12639 (N_12639,N_7735,N_7353);
nand U12640 (N_12640,N_9219,N_7891);
xnor U12641 (N_12641,N_5097,N_8618);
nand U12642 (N_12642,N_9861,N_6324);
or U12643 (N_12643,N_7419,N_8152);
xnor U12644 (N_12644,N_9453,N_6907);
nand U12645 (N_12645,N_8167,N_7440);
nand U12646 (N_12646,N_9444,N_6807);
nor U12647 (N_12647,N_8645,N_8935);
nor U12648 (N_12648,N_8595,N_5559);
nand U12649 (N_12649,N_6724,N_7241);
or U12650 (N_12650,N_7713,N_6877);
or U12651 (N_12651,N_7388,N_9602);
and U12652 (N_12652,N_9421,N_6225);
nand U12653 (N_12653,N_9062,N_8211);
and U12654 (N_12654,N_9294,N_7620);
or U12655 (N_12655,N_8078,N_8084);
nand U12656 (N_12656,N_5705,N_5046);
nor U12657 (N_12657,N_9999,N_9528);
or U12658 (N_12658,N_9674,N_5495);
xnor U12659 (N_12659,N_9418,N_8094);
and U12660 (N_12660,N_5121,N_5062);
or U12661 (N_12661,N_5898,N_7500);
or U12662 (N_12662,N_8926,N_9606);
xnor U12663 (N_12663,N_6641,N_6699);
and U12664 (N_12664,N_9961,N_5951);
nor U12665 (N_12665,N_8125,N_6105);
and U12666 (N_12666,N_7247,N_5276);
and U12667 (N_12667,N_6085,N_5510);
xor U12668 (N_12668,N_7951,N_5872);
xor U12669 (N_12669,N_9634,N_5184);
nor U12670 (N_12670,N_9935,N_9788);
and U12671 (N_12671,N_5339,N_9523);
nor U12672 (N_12672,N_6588,N_6158);
or U12673 (N_12673,N_6233,N_6800);
xnor U12674 (N_12674,N_6287,N_7014);
or U12675 (N_12675,N_6531,N_6483);
and U12676 (N_12676,N_9175,N_8746);
and U12677 (N_12677,N_6340,N_7429);
or U12678 (N_12678,N_6757,N_6292);
xor U12679 (N_12679,N_7896,N_9410);
and U12680 (N_12680,N_5834,N_8310);
nor U12681 (N_12681,N_9127,N_7770);
and U12682 (N_12682,N_5550,N_9285);
and U12683 (N_12683,N_6300,N_6293);
xor U12684 (N_12684,N_6599,N_8554);
and U12685 (N_12685,N_8104,N_9090);
and U12686 (N_12686,N_7672,N_9748);
nor U12687 (N_12687,N_8868,N_5675);
nand U12688 (N_12688,N_6201,N_7644);
nand U12689 (N_12689,N_8473,N_6320);
nand U12690 (N_12690,N_6930,N_7660);
nand U12691 (N_12691,N_8320,N_8494);
and U12692 (N_12692,N_9202,N_7550);
nor U12693 (N_12693,N_7943,N_5585);
nand U12694 (N_12694,N_5015,N_7364);
nand U12695 (N_12695,N_7472,N_8503);
or U12696 (N_12696,N_8996,N_7382);
xor U12697 (N_12697,N_7531,N_5380);
and U12698 (N_12698,N_8875,N_9425);
nor U12699 (N_12699,N_7415,N_6970);
xor U12700 (N_12700,N_8979,N_7564);
and U12701 (N_12701,N_7632,N_9165);
xor U12702 (N_12702,N_9072,N_7498);
nand U12703 (N_12703,N_8466,N_7379);
or U12704 (N_12704,N_6149,N_8147);
nand U12705 (N_12705,N_8918,N_5859);
nor U12706 (N_12706,N_9270,N_8897);
or U12707 (N_12707,N_8789,N_7857);
or U12708 (N_12708,N_6056,N_6239);
or U12709 (N_12709,N_6068,N_8017);
or U12710 (N_12710,N_8280,N_9386);
and U12711 (N_12711,N_9417,N_8248);
and U12712 (N_12712,N_9655,N_9469);
nand U12713 (N_12713,N_6658,N_6322);
and U12714 (N_12714,N_8309,N_7955);
and U12715 (N_12715,N_5723,N_5592);
nor U12716 (N_12716,N_9678,N_9911);
xnor U12717 (N_12717,N_7697,N_9760);
nor U12718 (N_12718,N_9048,N_6988);
and U12719 (N_12719,N_8572,N_5292);
nand U12720 (N_12720,N_5047,N_6008);
xor U12721 (N_12721,N_8358,N_5026);
or U12722 (N_12722,N_6275,N_5380);
xor U12723 (N_12723,N_6722,N_9796);
or U12724 (N_12724,N_6760,N_9961);
or U12725 (N_12725,N_8739,N_5744);
xnor U12726 (N_12726,N_8705,N_5737);
or U12727 (N_12727,N_7755,N_6591);
nor U12728 (N_12728,N_7581,N_8657);
nor U12729 (N_12729,N_5651,N_9562);
nand U12730 (N_12730,N_9844,N_8644);
nand U12731 (N_12731,N_6481,N_6900);
xnor U12732 (N_12732,N_9803,N_6211);
or U12733 (N_12733,N_5274,N_8580);
xor U12734 (N_12734,N_8352,N_8015);
nor U12735 (N_12735,N_9358,N_9202);
nor U12736 (N_12736,N_8892,N_8143);
xnor U12737 (N_12737,N_8279,N_5332);
nor U12738 (N_12738,N_6714,N_6852);
nor U12739 (N_12739,N_8697,N_5634);
nand U12740 (N_12740,N_6173,N_6118);
nand U12741 (N_12741,N_6255,N_5856);
nor U12742 (N_12742,N_6940,N_5860);
nand U12743 (N_12743,N_7817,N_9129);
nor U12744 (N_12744,N_9902,N_8487);
or U12745 (N_12745,N_7957,N_7402);
xnor U12746 (N_12746,N_8340,N_5212);
or U12747 (N_12747,N_5611,N_7056);
xnor U12748 (N_12748,N_8267,N_5551);
or U12749 (N_12749,N_9099,N_9577);
and U12750 (N_12750,N_6558,N_9341);
nand U12751 (N_12751,N_9413,N_6822);
and U12752 (N_12752,N_6878,N_7979);
or U12753 (N_12753,N_7693,N_5096);
xor U12754 (N_12754,N_7373,N_8861);
nand U12755 (N_12755,N_5809,N_7716);
xnor U12756 (N_12756,N_5200,N_6970);
nor U12757 (N_12757,N_9677,N_7484);
nor U12758 (N_12758,N_9593,N_5842);
and U12759 (N_12759,N_8225,N_7753);
or U12760 (N_12760,N_6016,N_8753);
and U12761 (N_12761,N_5473,N_7988);
or U12762 (N_12762,N_7861,N_6520);
or U12763 (N_12763,N_5561,N_6884);
and U12764 (N_12764,N_9659,N_7400);
nor U12765 (N_12765,N_5798,N_5605);
nand U12766 (N_12766,N_6562,N_7666);
and U12767 (N_12767,N_5397,N_6710);
nand U12768 (N_12768,N_9591,N_6843);
and U12769 (N_12769,N_9368,N_5590);
nor U12770 (N_12770,N_8681,N_6919);
nor U12771 (N_12771,N_8120,N_7460);
or U12772 (N_12772,N_8584,N_6694);
and U12773 (N_12773,N_9102,N_8680);
xnor U12774 (N_12774,N_7755,N_6574);
or U12775 (N_12775,N_8651,N_5462);
or U12776 (N_12776,N_9845,N_9671);
and U12777 (N_12777,N_6217,N_8671);
or U12778 (N_12778,N_5033,N_9763);
nand U12779 (N_12779,N_8556,N_9057);
and U12780 (N_12780,N_9092,N_5035);
xor U12781 (N_12781,N_9241,N_8059);
or U12782 (N_12782,N_6559,N_5603);
nand U12783 (N_12783,N_8854,N_9944);
nand U12784 (N_12784,N_5415,N_5998);
and U12785 (N_12785,N_9156,N_6921);
and U12786 (N_12786,N_5569,N_5666);
xnor U12787 (N_12787,N_5673,N_5256);
xnor U12788 (N_12788,N_6982,N_7232);
and U12789 (N_12789,N_5215,N_6790);
nor U12790 (N_12790,N_6677,N_9809);
xnor U12791 (N_12791,N_9163,N_7478);
nor U12792 (N_12792,N_9675,N_5170);
nor U12793 (N_12793,N_5953,N_7402);
or U12794 (N_12794,N_8730,N_6907);
nand U12795 (N_12795,N_8612,N_7176);
nor U12796 (N_12796,N_7175,N_7348);
and U12797 (N_12797,N_6767,N_5922);
xor U12798 (N_12798,N_6751,N_8349);
nand U12799 (N_12799,N_8978,N_6213);
xnor U12800 (N_12800,N_6266,N_7489);
xor U12801 (N_12801,N_6551,N_9974);
nor U12802 (N_12802,N_5840,N_7846);
and U12803 (N_12803,N_9621,N_6127);
nor U12804 (N_12804,N_7862,N_9770);
xnor U12805 (N_12805,N_7502,N_7917);
nor U12806 (N_12806,N_9337,N_8910);
or U12807 (N_12807,N_6516,N_8330);
or U12808 (N_12808,N_7249,N_7624);
xor U12809 (N_12809,N_9802,N_7455);
nand U12810 (N_12810,N_8309,N_7002);
xor U12811 (N_12811,N_5925,N_8757);
nor U12812 (N_12812,N_8434,N_9381);
nor U12813 (N_12813,N_5682,N_8734);
xnor U12814 (N_12814,N_5198,N_5591);
nand U12815 (N_12815,N_9548,N_9892);
nor U12816 (N_12816,N_6801,N_6557);
xor U12817 (N_12817,N_7221,N_6550);
or U12818 (N_12818,N_9700,N_7959);
or U12819 (N_12819,N_9594,N_5197);
nand U12820 (N_12820,N_6728,N_5547);
nand U12821 (N_12821,N_9929,N_8082);
nor U12822 (N_12822,N_8978,N_7430);
nand U12823 (N_12823,N_5136,N_5442);
xnor U12824 (N_12824,N_6446,N_6537);
nor U12825 (N_12825,N_9840,N_6494);
nor U12826 (N_12826,N_7262,N_5256);
nor U12827 (N_12827,N_9555,N_5969);
or U12828 (N_12828,N_5565,N_9370);
xnor U12829 (N_12829,N_5942,N_7444);
xor U12830 (N_12830,N_6092,N_9543);
nand U12831 (N_12831,N_7668,N_5340);
nor U12832 (N_12832,N_5045,N_7299);
or U12833 (N_12833,N_6815,N_8587);
nor U12834 (N_12834,N_7855,N_7698);
xor U12835 (N_12835,N_9942,N_6761);
xor U12836 (N_12836,N_6440,N_9819);
nand U12837 (N_12837,N_7705,N_8027);
xnor U12838 (N_12838,N_9218,N_8440);
xor U12839 (N_12839,N_7317,N_5010);
and U12840 (N_12840,N_7362,N_9637);
nor U12841 (N_12841,N_7792,N_5005);
nand U12842 (N_12842,N_5947,N_5953);
nor U12843 (N_12843,N_5533,N_9545);
and U12844 (N_12844,N_9475,N_8316);
xor U12845 (N_12845,N_6233,N_6048);
nor U12846 (N_12846,N_6661,N_6619);
xor U12847 (N_12847,N_9561,N_7761);
xnor U12848 (N_12848,N_8422,N_8568);
or U12849 (N_12849,N_8305,N_7519);
and U12850 (N_12850,N_7275,N_9975);
nand U12851 (N_12851,N_7431,N_8589);
nor U12852 (N_12852,N_9762,N_5262);
and U12853 (N_12853,N_8291,N_9199);
nand U12854 (N_12854,N_8077,N_5849);
and U12855 (N_12855,N_8480,N_7598);
nor U12856 (N_12856,N_5175,N_5858);
xor U12857 (N_12857,N_7453,N_6748);
or U12858 (N_12858,N_7350,N_7651);
or U12859 (N_12859,N_8387,N_5578);
nand U12860 (N_12860,N_9348,N_5109);
nand U12861 (N_12861,N_9037,N_6517);
nand U12862 (N_12862,N_9535,N_6972);
nand U12863 (N_12863,N_7378,N_6802);
nand U12864 (N_12864,N_9757,N_7629);
xor U12865 (N_12865,N_7006,N_6492);
nand U12866 (N_12866,N_9586,N_7752);
and U12867 (N_12867,N_7850,N_6088);
and U12868 (N_12868,N_5928,N_5568);
nor U12869 (N_12869,N_8413,N_9090);
or U12870 (N_12870,N_6815,N_7750);
xor U12871 (N_12871,N_9644,N_8382);
nor U12872 (N_12872,N_9852,N_7459);
xnor U12873 (N_12873,N_7501,N_9559);
nand U12874 (N_12874,N_5734,N_8513);
or U12875 (N_12875,N_8830,N_7381);
nor U12876 (N_12876,N_6631,N_5005);
xnor U12877 (N_12877,N_8473,N_6062);
and U12878 (N_12878,N_6580,N_6948);
or U12879 (N_12879,N_8283,N_8074);
nand U12880 (N_12880,N_5259,N_8016);
nand U12881 (N_12881,N_5486,N_9457);
nor U12882 (N_12882,N_9588,N_6091);
xor U12883 (N_12883,N_7915,N_7746);
nor U12884 (N_12884,N_8409,N_7036);
and U12885 (N_12885,N_5921,N_9149);
nor U12886 (N_12886,N_5886,N_5948);
or U12887 (N_12887,N_8814,N_8800);
nand U12888 (N_12888,N_6279,N_7400);
nor U12889 (N_12889,N_8710,N_8634);
nand U12890 (N_12890,N_9499,N_9698);
xnor U12891 (N_12891,N_6572,N_9051);
or U12892 (N_12892,N_7642,N_8310);
xor U12893 (N_12893,N_6536,N_6581);
xnor U12894 (N_12894,N_9077,N_5429);
nand U12895 (N_12895,N_7799,N_7845);
and U12896 (N_12896,N_8128,N_8552);
and U12897 (N_12897,N_9062,N_5660);
xor U12898 (N_12898,N_5428,N_6264);
or U12899 (N_12899,N_9336,N_9301);
nor U12900 (N_12900,N_8589,N_6889);
or U12901 (N_12901,N_6625,N_5503);
nor U12902 (N_12902,N_7576,N_9119);
or U12903 (N_12903,N_8390,N_5125);
nor U12904 (N_12904,N_8684,N_7372);
or U12905 (N_12905,N_6279,N_9561);
or U12906 (N_12906,N_6332,N_6699);
and U12907 (N_12907,N_6291,N_5687);
xor U12908 (N_12908,N_5345,N_9577);
nand U12909 (N_12909,N_9772,N_6771);
xnor U12910 (N_12910,N_5355,N_6495);
nor U12911 (N_12911,N_7985,N_5658);
xnor U12912 (N_12912,N_6268,N_6757);
and U12913 (N_12913,N_8090,N_7604);
and U12914 (N_12914,N_7678,N_8032);
nand U12915 (N_12915,N_8927,N_5190);
or U12916 (N_12916,N_6076,N_6827);
nor U12917 (N_12917,N_6498,N_9281);
and U12918 (N_12918,N_9075,N_6119);
and U12919 (N_12919,N_6774,N_9706);
nand U12920 (N_12920,N_7015,N_5144);
and U12921 (N_12921,N_5530,N_6393);
nor U12922 (N_12922,N_8285,N_9742);
or U12923 (N_12923,N_5873,N_9566);
or U12924 (N_12924,N_8406,N_9644);
nand U12925 (N_12925,N_7212,N_5500);
and U12926 (N_12926,N_7821,N_7906);
and U12927 (N_12927,N_8982,N_9489);
xor U12928 (N_12928,N_5280,N_5271);
or U12929 (N_12929,N_9565,N_8376);
nand U12930 (N_12930,N_7586,N_6629);
nand U12931 (N_12931,N_5355,N_8252);
or U12932 (N_12932,N_8114,N_9050);
and U12933 (N_12933,N_6673,N_6126);
xor U12934 (N_12934,N_5774,N_6384);
and U12935 (N_12935,N_5969,N_9470);
nor U12936 (N_12936,N_5978,N_9384);
and U12937 (N_12937,N_7463,N_6544);
nand U12938 (N_12938,N_6521,N_5433);
xor U12939 (N_12939,N_9943,N_9112);
or U12940 (N_12940,N_9381,N_6884);
nand U12941 (N_12941,N_7926,N_7354);
and U12942 (N_12942,N_6159,N_9295);
nand U12943 (N_12943,N_5927,N_5024);
or U12944 (N_12944,N_5473,N_6619);
nand U12945 (N_12945,N_7128,N_6326);
and U12946 (N_12946,N_5595,N_6278);
nand U12947 (N_12947,N_6673,N_8016);
xor U12948 (N_12948,N_5369,N_5768);
xor U12949 (N_12949,N_5831,N_5187);
nor U12950 (N_12950,N_9352,N_6634);
and U12951 (N_12951,N_7695,N_9647);
and U12952 (N_12952,N_5940,N_6573);
nand U12953 (N_12953,N_6816,N_8482);
nand U12954 (N_12954,N_5010,N_7821);
or U12955 (N_12955,N_9638,N_9898);
nor U12956 (N_12956,N_5836,N_6441);
and U12957 (N_12957,N_6297,N_7204);
xor U12958 (N_12958,N_5130,N_7644);
nand U12959 (N_12959,N_8041,N_6029);
and U12960 (N_12960,N_6749,N_9551);
or U12961 (N_12961,N_5487,N_8462);
or U12962 (N_12962,N_5482,N_7351);
xor U12963 (N_12963,N_6903,N_6000);
xnor U12964 (N_12964,N_5778,N_5671);
xor U12965 (N_12965,N_6168,N_7541);
or U12966 (N_12966,N_5158,N_9816);
xnor U12967 (N_12967,N_8154,N_9277);
nand U12968 (N_12968,N_7752,N_7806);
or U12969 (N_12969,N_9713,N_5876);
and U12970 (N_12970,N_7295,N_5394);
nor U12971 (N_12971,N_8010,N_7424);
or U12972 (N_12972,N_9136,N_5112);
nor U12973 (N_12973,N_6275,N_7536);
nor U12974 (N_12974,N_5061,N_5909);
nand U12975 (N_12975,N_7543,N_8776);
xnor U12976 (N_12976,N_8598,N_6006);
and U12977 (N_12977,N_8021,N_8890);
nand U12978 (N_12978,N_6712,N_7392);
and U12979 (N_12979,N_9740,N_7660);
xnor U12980 (N_12980,N_6597,N_8174);
nand U12981 (N_12981,N_7793,N_9692);
or U12982 (N_12982,N_8798,N_9598);
nand U12983 (N_12983,N_5151,N_5120);
nor U12984 (N_12984,N_8623,N_7590);
and U12985 (N_12985,N_9635,N_9645);
and U12986 (N_12986,N_8762,N_7100);
nor U12987 (N_12987,N_9151,N_8037);
nor U12988 (N_12988,N_7582,N_6620);
or U12989 (N_12989,N_7682,N_8198);
or U12990 (N_12990,N_7639,N_7117);
and U12991 (N_12991,N_7781,N_5798);
nand U12992 (N_12992,N_9887,N_8343);
nand U12993 (N_12993,N_7428,N_6216);
and U12994 (N_12994,N_5420,N_9663);
xnor U12995 (N_12995,N_5449,N_7001);
nor U12996 (N_12996,N_5576,N_7602);
or U12997 (N_12997,N_7271,N_5149);
and U12998 (N_12998,N_5286,N_5727);
nand U12999 (N_12999,N_6304,N_7721);
xnor U13000 (N_13000,N_8000,N_8602);
or U13001 (N_13001,N_7744,N_6558);
nor U13002 (N_13002,N_9887,N_6950);
nor U13003 (N_13003,N_5252,N_7658);
xnor U13004 (N_13004,N_6989,N_6794);
and U13005 (N_13005,N_8239,N_5944);
nand U13006 (N_13006,N_7744,N_7881);
or U13007 (N_13007,N_5185,N_5788);
and U13008 (N_13008,N_9615,N_8862);
nor U13009 (N_13009,N_6168,N_5875);
xor U13010 (N_13010,N_6824,N_9076);
xnor U13011 (N_13011,N_7689,N_6607);
nand U13012 (N_13012,N_6900,N_8404);
nand U13013 (N_13013,N_6735,N_9092);
nand U13014 (N_13014,N_7161,N_9096);
or U13015 (N_13015,N_7735,N_8703);
xnor U13016 (N_13016,N_6060,N_7635);
nand U13017 (N_13017,N_5304,N_5023);
xor U13018 (N_13018,N_5972,N_6559);
nor U13019 (N_13019,N_6846,N_6491);
nand U13020 (N_13020,N_8669,N_7294);
xnor U13021 (N_13021,N_6398,N_7543);
nor U13022 (N_13022,N_7276,N_8017);
and U13023 (N_13023,N_6099,N_8967);
nand U13024 (N_13024,N_8053,N_5974);
or U13025 (N_13025,N_8793,N_7731);
and U13026 (N_13026,N_7062,N_7868);
or U13027 (N_13027,N_6750,N_6335);
nor U13028 (N_13028,N_9441,N_8742);
or U13029 (N_13029,N_5456,N_6648);
nor U13030 (N_13030,N_5802,N_9919);
and U13031 (N_13031,N_5621,N_9170);
or U13032 (N_13032,N_6657,N_5372);
nand U13033 (N_13033,N_5089,N_6567);
xor U13034 (N_13034,N_9183,N_8936);
xor U13035 (N_13035,N_5117,N_5056);
or U13036 (N_13036,N_5906,N_9239);
nor U13037 (N_13037,N_8925,N_9739);
xnor U13038 (N_13038,N_9632,N_8154);
xor U13039 (N_13039,N_7535,N_6182);
nor U13040 (N_13040,N_8339,N_9537);
nand U13041 (N_13041,N_8875,N_9106);
nor U13042 (N_13042,N_6924,N_5630);
xor U13043 (N_13043,N_6771,N_6622);
nand U13044 (N_13044,N_9617,N_8303);
xnor U13045 (N_13045,N_5925,N_5024);
or U13046 (N_13046,N_7014,N_5065);
or U13047 (N_13047,N_5563,N_9879);
xor U13048 (N_13048,N_6048,N_7372);
xnor U13049 (N_13049,N_7557,N_7474);
nor U13050 (N_13050,N_9908,N_5325);
and U13051 (N_13051,N_7800,N_6831);
and U13052 (N_13052,N_5538,N_5027);
nor U13053 (N_13053,N_5206,N_8516);
nor U13054 (N_13054,N_8310,N_9314);
and U13055 (N_13055,N_7041,N_5007);
nor U13056 (N_13056,N_8593,N_7258);
xor U13057 (N_13057,N_5646,N_8869);
or U13058 (N_13058,N_7709,N_6966);
and U13059 (N_13059,N_7728,N_9391);
nor U13060 (N_13060,N_6406,N_6084);
nor U13061 (N_13061,N_8528,N_9815);
nand U13062 (N_13062,N_7681,N_5205);
nand U13063 (N_13063,N_6132,N_5544);
and U13064 (N_13064,N_7674,N_5227);
or U13065 (N_13065,N_6176,N_5176);
nand U13066 (N_13066,N_7167,N_5149);
nor U13067 (N_13067,N_7434,N_6365);
xnor U13068 (N_13068,N_7988,N_7239);
nand U13069 (N_13069,N_7304,N_8733);
or U13070 (N_13070,N_9517,N_6134);
nand U13071 (N_13071,N_5565,N_8254);
xnor U13072 (N_13072,N_9662,N_7459);
or U13073 (N_13073,N_5084,N_5102);
and U13074 (N_13074,N_5116,N_7959);
or U13075 (N_13075,N_8940,N_7909);
xnor U13076 (N_13076,N_5505,N_6755);
nor U13077 (N_13077,N_7546,N_6757);
and U13078 (N_13078,N_8549,N_8868);
nor U13079 (N_13079,N_7993,N_5694);
nand U13080 (N_13080,N_9050,N_6747);
or U13081 (N_13081,N_9705,N_6557);
or U13082 (N_13082,N_7918,N_8733);
or U13083 (N_13083,N_6377,N_7420);
or U13084 (N_13084,N_9670,N_7060);
and U13085 (N_13085,N_7771,N_8356);
xnor U13086 (N_13086,N_7797,N_9441);
and U13087 (N_13087,N_9179,N_5710);
nor U13088 (N_13088,N_9531,N_7583);
or U13089 (N_13089,N_5309,N_6963);
xor U13090 (N_13090,N_7870,N_5894);
xnor U13091 (N_13091,N_8173,N_6569);
xor U13092 (N_13092,N_5447,N_5746);
nor U13093 (N_13093,N_9803,N_5585);
nor U13094 (N_13094,N_8555,N_9572);
xor U13095 (N_13095,N_8931,N_8675);
or U13096 (N_13096,N_5463,N_7424);
or U13097 (N_13097,N_5493,N_9836);
or U13098 (N_13098,N_6516,N_6982);
or U13099 (N_13099,N_6382,N_5606);
or U13100 (N_13100,N_9299,N_5617);
or U13101 (N_13101,N_7810,N_5208);
xnor U13102 (N_13102,N_5262,N_6057);
or U13103 (N_13103,N_5823,N_8121);
nand U13104 (N_13104,N_7344,N_5827);
or U13105 (N_13105,N_9015,N_9179);
xor U13106 (N_13106,N_8467,N_6126);
nor U13107 (N_13107,N_6105,N_9504);
and U13108 (N_13108,N_6186,N_5225);
nand U13109 (N_13109,N_5040,N_7720);
xor U13110 (N_13110,N_9868,N_7361);
nand U13111 (N_13111,N_6804,N_8426);
xnor U13112 (N_13112,N_5437,N_7686);
and U13113 (N_13113,N_5975,N_5829);
xor U13114 (N_13114,N_6909,N_7763);
nand U13115 (N_13115,N_9507,N_7516);
nand U13116 (N_13116,N_9089,N_5261);
nor U13117 (N_13117,N_9845,N_8529);
xor U13118 (N_13118,N_9887,N_6148);
nand U13119 (N_13119,N_6789,N_8511);
xnor U13120 (N_13120,N_8295,N_5057);
and U13121 (N_13121,N_6339,N_9474);
xor U13122 (N_13122,N_7513,N_7795);
nor U13123 (N_13123,N_7019,N_9352);
or U13124 (N_13124,N_7553,N_9851);
and U13125 (N_13125,N_5087,N_6781);
xor U13126 (N_13126,N_6036,N_8720);
xor U13127 (N_13127,N_5164,N_6157);
nor U13128 (N_13128,N_9267,N_7208);
and U13129 (N_13129,N_6238,N_7939);
and U13130 (N_13130,N_6740,N_6339);
or U13131 (N_13131,N_6858,N_9325);
nand U13132 (N_13132,N_8860,N_9404);
and U13133 (N_13133,N_5032,N_9520);
or U13134 (N_13134,N_7089,N_5193);
nand U13135 (N_13135,N_5133,N_6276);
xor U13136 (N_13136,N_9754,N_8600);
xor U13137 (N_13137,N_9647,N_9085);
or U13138 (N_13138,N_8361,N_9743);
or U13139 (N_13139,N_8798,N_8373);
or U13140 (N_13140,N_7542,N_8095);
and U13141 (N_13141,N_8076,N_5200);
xnor U13142 (N_13142,N_8015,N_6677);
or U13143 (N_13143,N_6389,N_7070);
nor U13144 (N_13144,N_5627,N_6173);
nand U13145 (N_13145,N_8473,N_6484);
nand U13146 (N_13146,N_8387,N_7404);
xnor U13147 (N_13147,N_7391,N_9785);
or U13148 (N_13148,N_5880,N_6714);
xor U13149 (N_13149,N_5315,N_7533);
nor U13150 (N_13150,N_8504,N_6856);
or U13151 (N_13151,N_6730,N_9588);
or U13152 (N_13152,N_5584,N_7565);
nor U13153 (N_13153,N_7072,N_6952);
or U13154 (N_13154,N_9543,N_8302);
or U13155 (N_13155,N_6100,N_5161);
and U13156 (N_13156,N_8141,N_7427);
and U13157 (N_13157,N_8675,N_5874);
nor U13158 (N_13158,N_9244,N_7593);
nand U13159 (N_13159,N_5616,N_8882);
xnor U13160 (N_13160,N_5989,N_5603);
and U13161 (N_13161,N_6720,N_6273);
xor U13162 (N_13162,N_8126,N_6567);
nor U13163 (N_13163,N_6675,N_7500);
or U13164 (N_13164,N_7908,N_7463);
nand U13165 (N_13165,N_6220,N_9550);
and U13166 (N_13166,N_5568,N_5949);
or U13167 (N_13167,N_8046,N_8676);
or U13168 (N_13168,N_8053,N_5106);
xnor U13169 (N_13169,N_9693,N_6796);
and U13170 (N_13170,N_5278,N_6503);
or U13171 (N_13171,N_8594,N_7868);
or U13172 (N_13172,N_6422,N_5126);
nor U13173 (N_13173,N_8743,N_5715);
or U13174 (N_13174,N_6113,N_8992);
xnor U13175 (N_13175,N_6023,N_6224);
nor U13176 (N_13176,N_5604,N_9053);
and U13177 (N_13177,N_6224,N_6815);
xor U13178 (N_13178,N_7724,N_8576);
or U13179 (N_13179,N_7494,N_6366);
nand U13180 (N_13180,N_7256,N_6990);
and U13181 (N_13181,N_9839,N_7591);
nor U13182 (N_13182,N_5624,N_7621);
nor U13183 (N_13183,N_9451,N_8452);
nand U13184 (N_13184,N_8502,N_8527);
or U13185 (N_13185,N_6260,N_5972);
and U13186 (N_13186,N_9946,N_9437);
nor U13187 (N_13187,N_5386,N_9870);
or U13188 (N_13188,N_9882,N_5044);
or U13189 (N_13189,N_6596,N_7128);
nor U13190 (N_13190,N_6464,N_9664);
or U13191 (N_13191,N_9018,N_8840);
and U13192 (N_13192,N_7655,N_7561);
and U13193 (N_13193,N_6107,N_8295);
nor U13194 (N_13194,N_5721,N_9063);
or U13195 (N_13195,N_6590,N_7203);
xnor U13196 (N_13196,N_9650,N_5296);
nor U13197 (N_13197,N_7392,N_7401);
nand U13198 (N_13198,N_9667,N_9484);
xnor U13199 (N_13199,N_5892,N_5007);
xor U13200 (N_13200,N_7572,N_7625);
xnor U13201 (N_13201,N_6842,N_9504);
xor U13202 (N_13202,N_8967,N_6367);
nand U13203 (N_13203,N_9955,N_8212);
nor U13204 (N_13204,N_6213,N_8279);
and U13205 (N_13205,N_6226,N_9417);
or U13206 (N_13206,N_5724,N_5846);
xor U13207 (N_13207,N_8981,N_5913);
xor U13208 (N_13208,N_6137,N_6994);
nand U13209 (N_13209,N_5369,N_6011);
or U13210 (N_13210,N_9079,N_7531);
nor U13211 (N_13211,N_6489,N_5669);
xnor U13212 (N_13212,N_6660,N_9465);
nor U13213 (N_13213,N_8394,N_6246);
and U13214 (N_13214,N_9889,N_8107);
and U13215 (N_13215,N_8827,N_9627);
nand U13216 (N_13216,N_8746,N_5939);
or U13217 (N_13217,N_9007,N_7478);
and U13218 (N_13218,N_7372,N_8765);
xor U13219 (N_13219,N_6633,N_9991);
nand U13220 (N_13220,N_7522,N_5114);
or U13221 (N_13221,N_7951,N_7961);
nor U13222 (N_13222,N_9762,N_9547);
nand U13223 (N_13223,N_9185,N_9723);
nand U13224 (N_13224,N_6066,N_6800);
and U13225 (N_13225,N_8350,N_5132);
and U13226 (N_13226,N_5644,N_8211);
or U13227 (N_13227,N_7583,N_9365);
or U13228 (N_13228,N_6318,N_6437);
or U13229 (N_13229,N_7354,N_7845);
nor U13230 (N_13230,N_8780,N_9148);
and U13231 (N_13231,N_6866,N_7030);
nor U13232 (N_13232,N_7388,N_6324);
nor U13233 (N_13233,N_6132,N_7511);
nor U13234 (N_13234,N_6236,N_6331);
xor U13235 (N_13235,N_6028,N_8255);
and U13236 (N_13236,N_8051,N_9287);
xnor U13237 (N_13237,N_5063,N_8267);
or U13238 (N_13238,N_5671,N_9184);
or U13239 (N_13239,N_8091,N_9561);
nand U13240 (N_13240,N_5064,N_8065);
nand U13241 (N_13241,N_6973,N_5683);
xnor U13242 (N_13242,N_9615,N_5939);
xor U13243 (N_13243,N_7043,N_5113);
xnor U13244 (N_13244,N_5367,N_9861);
or U13245 (N_13245,N_6094,N_5033);
nor U13246 (N_13246,N_6257,N_9310);
nand U13247 (N_13247,N_8794,N_6111);
xor U13248 (N_13248,N_9423,N_6591);
nor U13249 (N_13249,N_5048,N_6774);
nor U13250 (N_13250,N_5851,N_5537);
nand U13251 (N_13251,N_9079,N_5171);
and U13252 (N_13252,N_7647,N_6096);
and U13253 (N_13253,N_5596,N_7390);
nand U13254 (N_13254,N_5502,N_9276);
xor U13255 (N_13255,N_6889,N_5927);
nor U13256 (N_13256,N_8031,N_8902);
or U13257 (N_13257,N_6877,N_8031);
or U13258 (N_13258,N_5858,N_5111);
and U13259 (N_13259,N_9186,N_8831);
or U13260 (N_13260,N_9668,N_6259);
nor U13261 (N_13261,N_9972,N_9885);
nand U13262 (N_13262,N_7332,N_7072);
nand U13263 (N_13263,N_6413,N_7766);
or U13264 (N_13264,N_6238,N_5420);
xnor U13265 (N_13265,N_6525,N_6586);
nand U13266 (N_13266,N_6674,N_9984);
nor U13267 (N_13267,N_9921,N_5785);
nor U13268 (N_13268,N_8712,N_8026);
and U13269 (N_13269,N_9269,N_7131);
xor U13270 (N_13270,N_9048,N_7856);
and U13271 (N_13271,N_7109,N_8660);
and U13272 (N_13272,N_6798,N_6661);
nor U13273 (N_13273,N_7013,N_9700);
nor U13274 (N_13274,N_5029,N_8896);
nor U13275 (N_13275,N_9533,N_8503);
nand U13276 (N_13276,N_8349,N_7826);
and U13277 (N_13277,N_8392,N_7624);
or U13278 (N_13278,N_5952,N_8798);
or U13279 (N_13279,N_9924,N_8042);
and U13280 (N_13280,N_9877,N_5835);
xor U13281 (N_13281,N_6005,N_6400);
or U13282 (N_13282,N_9136,N_8546);
nand U13283 (N_13283,N_5178,N_5749);
nand U13284 (N_13284,N_6820,N_7294);
and U13285 (N_13285,N_5482,N_6183);
and U13286 (N_13286,N_5066,N_6552);
nand U13287 (N_13287,N_5788,N_9406);
xor U13288 (N_13288,N_8101,N_6752);
or U13289 (N_13289,N_8695,N_9740);
xnor U13290 (N_13290,N_6299,N_5516);
and U13291 (N_13291,N_9687,N_6918);
or U13292 (N_13292,N_8902,N_6798);
nand U13293 (N_13293,N_9867,N_8181);
nor U13294 (N_13294,N_9282,N_5684);
xor U13295 (N_13295,N_8373,N_6056);
nor U13296 (N_13296,N_7383,N_5251);
or U13297 (N_13297,N_6410,N_9343);
and U13298 (N_13298,N_6036,N_8818);
nor U13299 (N_13299,N_8807,N_6836);
xnor U13300 (N_13300,N_9396,N_6566);
nor U13301 (N_13301,N_9352,N_7856);
nor U13302 (N_13302,N_7659,N_7017);
nand U13303 (N_13303,N_5327,N_7724);
nor U13304 (N_13304,N_8076,N_9622);
nand U13305 (N_13305,N_7924,N_5006);
or U13306 (N_13306,N_5521,N_5447);
nor U13307 (N_13307,N_5075,N_8672);
and U13308 (N_13308,N_6582,N_7308);
nand U13309 (N_13309,N_8470,N_5262);
nor U13310 (N_13310,N_8520,N_7100);
nand U13311 (N_13311,N_9296,N_8787);
nor U13312 (N_13312,N_5022,N_6590);
nand U13313 (N_13313,N_6399,N_8104);
and U13314 (N_13314,N_9752,N_9945);
nor U13315 (N_13315,N_6796,N_9827);
xor U13316 (N_13316,N_9918,N_6259);
and U13317 (N_13317,N_7157,N_8868);
nand U13318 (N_13318,N_5132,N_8763);
nor U13319 (N_13319,N_6253,N_7602);
xor U13320 (N_13320,N_8312,N_9064);
nand U13321 (N_13321,N_6895,N_8206);
nand U13322 (N_13322,N_5694,N_9638);
nand U13323 (N_13323,N_9959,N_6863);
or U13324 (N_13324,N_8668,N_8559);
or U13325 (N_13325,N_9014,N_6663);
and U13326 (N_13326,N_9050,N_5726);
nand U13327 (N_13327,N_6962,N_9942);
xor U13328 (N_13328,N_9570,N_6868);
nand U13329 (N_13329,N_7722,N_8577);
and U13330 (N_13330,N_5894,N_7755);
and U13331 (N_13331,N_8418,N_8825);
nor U13332 (N_13332,N_7496,N_5219);
xnor U13333 (N_13333,N_8388,N_9061);
and U13334 (N_13334,N_5082,N_8065);
xor U13335 (N_13335,N_5470,N_5014);
xnor U13336 (N_13336,N_5387,N_9252);
nor U13337 (N_13337,N_9735,N_7059);
and U13338 (N_13338,N_9740,N_7374);
nor U13339 (N_13339,N_9809,N_9656);
and U13340 (N_13340,N_7898,N_7029);
xor U13341 (N_13341,N_8614,N_9053);
xor U13342 (N_13342,N_6162,N_7208);
and U13343 (N_13343,N_9274,N_8375);
nand U13344 (N_13344,N_5079,N_6092);
and U13345 (N_13345,N_9231,N_8166);
xor U13346 (N_13346,N_6280,N_9736);
and U13347 (N_13347,N_9215,N_7538);
nand U13348 (N_13348,N_7883,N_6611);
and U13349 (N_13349,N_6606,N_8571);
nor U13350 (N_13350,N_5861,N_9067);
nor U13351 (N_13351,N_5056,N_8989);
nand U13352 (N_13352,N_6810,N_7478);
or U13353 (N_13353,N_8916,N_5798);
xnor U13354 (N_13354,N_7961,N_8641);
or U13355 (N_13355,N_9412,N_6112);
nand U13356 (N_13356,N_8114,N_9858);
and U13357 (N_13357,N_8643,N_6734);
or U13358 (N_13358,N_7488,N_5987);
nor U13359 (N_13359,N_9965,N_6666);
nand U13360 (N_13360,N_7804,N_5880);
xor U13361 (N_13361,N_7014,N_9058);
nand U13362 (N_13362,N_8675,N_6652);
or U13363 (N_13363,N_7045,N_7329);
and U13364 (N_13364,N_7378,N_7480);
nand U13365 (N_13365,N_6232,N_7443);
and U13366 (N_13366,N_8204,N_5999);
or U13367 (N_13367,N_6241,N_9498);
nor U13368 (N_13368,N_5439,N_9752);
and U13369 (N_13369,N_6797,N_7263);
and U13370 (N_13370,N_5464,N_7682);
nand U13371 (N_13371,N_8040,N_6213);
nor U13372 (N_13372,N_6621,N_8419);
nor U13373 (N_13373,N_8659,N_7518);
nand U13374 (N_13374,N_7090,N_9166);
and U13375 (N_13375,N_5560,N_7564);
or U13376 (N_13376,N_6190,N_8163);
or U13377 (N_13377,N_6896,N_6176);
or U13378 (N_13378,N_8514,N_6068);
xnor U13379 (N_13379,N_5142,N_9135);
nor U13380 (N_13380,N_6458,N_5135);
nor U13381 (N_13381,N_7715,N_7444);
nor U13382 (N_13382,N_5988,N_9025);
nor U13383 (N_13383,N_7940,N_5654);
nor U13384 (N_13384,N_6856,N_9124);
or U13385 (N_13385,N_9559,N_9750);
nor U13386 (N_13386,N_7407,N_8356);
nor U13387 (N_13387,N_6953,N_5258);
nand U13388 (N_13388,N_7834,N_9744);
xor U13389 (N_13389,N_9301,N_6448);
or U13390 (N_13390,N_6386,N_5747);
xor U13391 (N_13391,N_7237,N_6636);
nand U13392 (N_13392,N_9730,N_5633);
nor U13393 (N_13393,N_6119,N_5415);
nand U13394 (N_13394,N_7878,N_9002);
nand U13395 (N_13395,N_8569,N_7983);
or U13396 (N_13396,N_6493,N_9765);
xnor U13397 (N_13397,N_6404,N_6927);
or U13398 (N_13398,N_5698,N_9286);
nand U13399 (N_13399,N_7027,N_8148);
nor U13400 (N_13400,N_6745,N_6237);
nand U13401 (N_13401,N_6441,N_9254);
and U13402 (N_13402,N_8059,N_8318);
nor U13403 (N_13403,N_8771,N_8463);
or U13404 (N_13404,N_9769,N_9741);
and U13405 (N_13405,N_7729,N_8409);
or U13406 (N_13406,N_6973,N_6592);
nand U13407 (N_13407,N_6298,N_5438);
nand U13408 (N_13408,N_5801,N_8637);
and U13409 (N_13409,N_6816,N_5584);
and U13410 (N_13410,N_9574,N_6687);
nand U13411 (N_13411,N_5193,N_5744);
nor U13412 (N_13412,N_8520,N_7541);
nor U13413 (N_13413,N_9297,N_8783);
and U13414 (N_13414,N_6430,N_5858);
nor U13415 (N_13415,N_7390,N_7924);
or U13416 (N_13416,N_5225,N_6093);
xor U13417 (N_13417,N_6645,N_7514);
nand U13418 (N_13418,N_8920,N_8670);
nand U13419 (N_13419,N_9049,N_5636);
xor U13420 (N_13420,N_8548,N_5104);
xnor U13421 (N_13421,N_7853,N_6599);
or U13422 (N_13422,N_8910,N_6875);
nor U13423 (N_13423,N_7206,N_5213);
nor U13424 (N_13424,N_8948,N_7798);
nand U13425 (N_13425,N_8206,N_7470);
nand U13426 (N_13426,N_8412,N_9263);
nor U13427 (N_13427,N_6926,N_5788);
or U13428 (N_13428,N_8334,N_8660);
or U13429 (N_13429,N_8264,N_5909);
nor U13430 (N_13430,N_5265,N_9869);
and U13431 (N_13431,N_7102,N_5874);
xnor U13432 (N_13432,N_5993,N_6354);
xor U13433 (N_13433,N_7214,N_7507);
nand U13434 (N_13434,N_6164,N_9425);
or U13435 (N_13435,N_9709,N_6724);
nor U13436 (N_13436,N_5302,N_9726);
and U13437 (N_13437,N_8430,N_9956);
nand U13438 (N_13438,N_9371,N_5560);
xnor U13439 (N_13439,N_7813,N_9891);
or U13440 (N_13440,N_9287,N_5715);
or U13441 (N_13441,N_5734,N_9423);
xnor U13442 (N_13442,N_8818,N_5916);
and U13443 (N_13443,N_5516,N_5520);
and U13444 (N_13444,N_5301,N_8896);
xnor U13445 (N_13445,N_5272,N_9178);
and U13446 (N_13446,N_6537,N_7261);
xnor U13447 (N_13447,N_9626,N_5427);
nand U13448 (N_13448,N_6037,N_5767);
xnor U13449 (N_13449,N_9186,N_9826);
nand U13450 (N_13450,N_7612,N_6398);
nor U13451 (N_13451,N_7666,N_7723);
nor U13452 (N_13452,N_5223,N_8693);
nand U13453 (N_13453,N_6644,N_9388);
and U13454 (N_13454,N_5396,N_6816);
and U13455 (N_13455,N_8676,N_9178);
xor U13456 (N_13456,N_7794,N_7611);
nor U13457 (N_13457,N_7670,N_8057);
nand U13458 (N_13458,N_5739,N_7169);
nor U13459 (N_13459,N_9515,N_8069);
or U13460 (N_13460,N_8784,N_9246);
and U13461 (N_13461,N_8420,N_5443);
nor U13462 (N_13462,N_6709,N_5963);
xor U13463 (N_13463,N_9524,N_7864);
and U13464 (N_13464,N_6818,N_9085);
nand U13465 (N_13465,N_9302,N_9748);
nand U13466 (N_13466,N_7380,N_6651);
or U13467 (N_13467,N_9473,N_9062);
xor U13468 (N_13468,N_5471,N_6637);
or U13469 (N_13469,N_5326,N_7962);
xnor U13470 (N_13470,N_7966,N_6877);
nor U13471 (N_13471,N_7915,N_8420);
or U13472 (N_13472,N_8236,N_8349);
nand U13473 (N_13473,N_8702,N_9786);
and U13474 (N_13474,N_9044,N_9375);
and U13475 (N_13475,N_8490,N_7780);
nor U13476 (N_13476,N_9446,N_6987);
xnor U13477 (N_13477,N_6087,N_6011);
nor U13478 (N_13478,N_6064,N_8784);
or U13479 (N_13479,N_6073,N_8677);
or U13480 (N_13480,N_6503,N_5608);
or U13481 (N_13481,N_5236,N_6070);
nand U13482 (N_13482,N_7513,N_7579);
nand U13483 (N_13483,N_6909,N_9926);
and U13484 (N_13484,N_8693,N_9535);
nand U13485 (N_13485,N_5547,N_6873);
nor U13486 (N_13486,N_9151,N_5712);
or U13487 (N_13487,N_8240,N_9521);
and U13488 (N_13488,N_7467,N_8214);
and U13489 (N_13489,N_7847,N_7389);
nand U13490 (N_13490,N_6255,N_6813);
or U13491 (N_13491,N_5630,N_6076);
nor U13492 (N_13492,N_7722,N_6294);
nand U13493 (N_13493,N_6258,N_6708);
nand U13494 (N_13494,N_5733,N_7862);
xnor U13495 (N_13495,N_6835,N_9695);
xnor U13496 (N_13496,N_6671,N_5197);
nand U13497 (N_13497,N_9528,N_6444);
and U13498 (N_13498,N_9595,N_6334);
and U13499 (N_13499,N_8807,N_8885);
xnor U13500 (N_13500,N_9848,N_8137);
xor U13501 (N_13501,N_9808,N_8521);
nand U13502 (N_13502,N_8017,N_8518);
xor U13503 (N_13503,N_9651,N_7863);
and U13504 (N_13504,N_9942,N_8009);
or U13505 (N_13505,N_9246,N_9040);
nor U13506 (N_13506,N_8298,N_7402);
and U13507 (N_13507,N_9804,N_7117);
or U13508 (N_13508,N_6201,N_6669);
or U13509 (N_13509,N_8262,N_5997);
nor U13510 (N_13510,N_9618,N_5712);
nor U13511 (N_13511,N_6973,N_9753);
and U13512 (N_13512,N_8920,N_7107);
nor U13513 (N_13513,N_6190,N_7413);
xor U13514 (N_13514,N_7512,N_5027);
and U13515 (N_13515,N_6509,N_8251);
nand U13516 (N_13516,N_7007,N_9494);
nor U13517 (N_13517,N_8149,N_9207);
or U13518 (N_13518,N_5782,N_9688);
or U13519 (N_13519,N_7467,N_5691);
nand U13520 (N_13520,N_8074,N_8320);
xnor U13521 (N_13521,N_9542,N_9553);
and U13522 (N_13522,N_9468,N_8683);
or U13523 (N_13523,N_7162,N_7118);
and U13524 (N_13524,N_6266,N_9844);
or U13525 (N_13525,N_9602,N_9968);
and U13526 (N_13526,N_5761,N_5465);
nor U13527 (N_13527,N_7809,N_8281);
or U13528 (N_13528,N_5644,N_9877);
nor U13529 (N_13529,N_8810,N_5965);
xnor U13530 (N_13530,N_6209,N_6091);
nand U13531 (N_13531,N_6102,N_6600);
or U13532 (N_13532,N_7724,N_7260);
nand U13533 (N_13533,N_9004,N_5510);
nand U13534 (N_13534,N_8427,N_6230);
nor U13535 (N_13535,N_9918,N_9213);
nand U13536 (N_13536,N_6212,N_8924);
and U13537 (N_13537,N_8455,N_7811);
and U13538 (N_13538,N_7070,N_6731);
or U13539 (N_13539,N_6829,N_6885);
xnor U13540 (N_13540,N_5865,N_5906);
nand U13541 (N_13541,N_9348,N_8695);
and U13542 (N_13542,N_8345,N_7542);
nor U13543 (N_13543,N_7162,N_5855);
or U13544 (N_13544,N_5797,N_7535);
xor U13545 (N_13545,N_9565,N_8276);
nor U13546 (N_13546,N_6127,N_5427);
and U13547 (N_13547,N_6930,N_6700);
or U13548 (N_13548,N_8155,N_9265);
xnor U13549 (N_13549,N_6257,N_8507);
xnor U13550 (N_13550,N_5236,N_5193);
nand U13551 (N_13551,N_7489,N_7846);
xor U13552 (N_13552,N_9261,N_7702);
xor U13553 (N_13553,N_7790,N_6828);
and U13554 (N_13554,N_8488,N_9904);
xor U13555 (N_13555,N_9657,N_8111);
xnor U13556 (N_13556,N_5580,N_9840);
or U13557 (N_13557,N_8751,N_7385);
xnor U13558 (N_13558,N_5946,N_9194);
nor U13559 (N_13559,N_8773,N_5946);
and U13560 (N_13560,N_5490,N_6378);
nand U13561 (N_13561,N_6690,N_9094);
and U13562 (N_13562,N_7479,N_6435);
or U13563 (N_13563,N_5389,N_7779);
or U13564 (N_13564,N_5022,N_5830);
xor U13565 (N_13565,N_5214,N_5517);
and U13566 (N_13566,N_9524,N_6183);
or U13567 (N_13567,N_9701,N_5924);
nand U13568 (N_13568,N_9754,N_6085);
nand U13569 (N_13569,N_6420,N_9177);
xnor U13570 (N_13570,N_6548,N_5135);
nand U13571 (N_13571,N_9403,N_8901);
and U13572 (N_13572,N_5619,N_9937);
xor U13573 (N_13573,N_8424,N_5439);
xor U13574 (N_13574,N_8058,N_5697);
or U13575 (N_13575,N_8122,N_5468);
xnor U13576 (N_13576,N_5719,N_6306);
and U13577 (N_13577,N_6193,N_6914);
xnor U13578 (N_13578,N_6538,N_7130);
xor U13579 (N_13579,N_5037,N_8753);
nor U13580 (N_13580,N_6568,N_6119);
xor U13581 (N_13581,N_6000,N_9949);
nand U13582 (N_13582,N_8657,N_9288);
xnor U13583 (N_13583,N_5203,N_7879);
xnor U13584 (N_13584,N_8228,N_8839);
or U13585 (N_13585,N_7628,N_8482);
nand U13586 (N_13586,N_8651,N_7982);
nor U13587 (N_13587,N_8089,N_9733);
or U13588 (N_13588,N_6728,N_5299);
or U13589 (N_13589,N_8250,N_9048);
or U13590 (N_13590,N_5976,N_7800);
xnor U13591 (N_13591,N_6231,N_7178);
nand U13592 (N_13592,N_5520,N_8347);
nand U13593 (N_13593,N_5167,N_7154);
xnor U13594 (N_13594,N_8632,N_9085);
nand U13595 (N_13595,N_6224,N_9323);
or U13596 (N_13596,N_9115,N_9545);
or U13597 (N_13597,N_6637,N_8475);
xnor U13598 (N_13598,N_9088,N_9552);
and U13599 (N_13599,N_6181,N_6379);
xor U13600 (N_13600,N_6600,N_6571);
and U13601 (N_13601,N_5749,N_5057);
xnor U13602 (N_13602,N_8389,N_7098);
nand U13603 (N_13603,N_7182,N_6904);
and U13604 (N_13604,N_6425,N_7548);
nor U13605 (N_13605,N_9158,N_6006);
nand U13606 (N_13606,N_7728,N_5020);
nand U13607 (N_13607,N_5151,N_5228);
or U13608 (N_13608,N_9555,N_6265);
xor U13609 (N_13609,N_8320,N_6031);
nand U13610 (N_13610,N_7067,N_7215);
and U13611 (N_13611,N_7548,N_6730);
or U13612 (N_13612,N_9396,N_5788);
nor U13613 (N_13613,N_6732,N_7826);
or U13614 (N_13614,N_7950,N_9213);
xor U13615 (N_13615,N_7732,N_5471);
nand U13616 (N_13616,N_9856,N_9427);
xnor U13617 (N_13617,N_9401,N_6764);
nand U13618 (N_13618,N_5032,N_5289);
or U13619 (N_13619,N_6393,N_8559);
xor U13620 (N_13620,N_8205,N_8366);
nor U13621 (N_13621,N_9515,N_7324);
or U13622 (N_13622,N_9952,N_9476);
nor U13623 (N_13623,N_5171,N_7436);
or U13624 (N_13624,N_9001,N_8666);
xnor U13625 (N_13625,N_9596,N_9289);
and U13626 (N_13626,N_9025,N_6275);
or U13627 (N_13627,N_5081,N_8327);
nand U13628 (N_13628,N_8794,N_8474);
or U13629 (N_13629,N_7684,N_5548);
nand U13630 (N_13630,N_7261,N_8238);
xor U13631 (N_13631,N_8954,N_8881);
or U13632 (N_13632,N_9066,N_8842);
or U13633 (N_13633,N_9641,N_8324);
and U13634 (N_13634,N_8084,N_6270);
xor U13635 (N_13635,N_8967,N_9179);
nand U13636 (N_13636,N_6421,N_7064);
and U13637 (N_13637,N_8077,N_6749);
xnor U13638 (N_13638,N_5938,N_9869);
or U13639 (N_13639,N_9061,N_6747);
xnor U13640 (N_13640,N_9917,N_8051);
nor U13641 (N_13641,N_8127,N_7506);
nand U13642 (N_13642,N_9695,N_8526);
or U13643 (N_13643,N_9665,N_8540);
nand U13644 (N_13644,N_8376,N_6222);
nor U13645 (N_13645,N_7546,N_8791);
nor U13646 (N_13646,N_5042,N_5121);
xnor U13647 (N_13647,N_7326,N_9119);
nand U13648 (N_13648,N_8975,N_5789);
nand U13649 (N_13649,N_5757,N_6248);
nor U13650 (N_13650,N_6388,N_7018);
nor U13651 (N_13651,N_8242,N_5437);
or U13652 (N_13652,N_8954,N_6987);
nor U13653 (N_13653,N_9347,N_7362);
and U13654 (N_13654,N_7512,N_8679);
xor U13655 (N_13655,N_9008,N_7006);
nor U13656 (N_13656,N_8917,N_9567);
and U13657 (N_13657,N_9714,N_5834);
xnor U13658 (N_13658,N_5491,N_8539);
or U13659 (N_13659,N_5500,N_7473);
xor U13660 (N_13660,N_5221,N_7885);
nor U13661 (N_13661,N_8361,N_8290);
nor U13662 (N_13662,N_6933,N_5849);
or U13663 (N_13663,N_9068,N_7736);
nand U13664 (N_13664,N_6912,N_5689);
and U13665 (N_13665,N_5961,N_9483);
or U13666 (N_13666,N_6407,N_5396);
nand U13667 (N_13667,N_8591,N_6228);
xnor U13668 (N_13668,N_8348,N_6573);
nor U13669 (N_13669,N_5583,N_9285);
or U13670 (N_13670,N_9512,N_5207);
xnor U13671 (N_13671,N_5503,N_6184);
or U13672 (N_13672,N_7914,N_6048);
nor U13673 (N_13673,N_9755,N_7860);
nand U13674 (N_13674,N_5493,N_5748);
xor U13675 (N_13675,N_5402,N_6466);
nor U13676 (N_13676,N_8242,N_7734);
xnor U13677 (N_13677,N_5987,N_7491);
nor U13678 (N_13678,N_9863,N_9345);
and U13679 (N_13679,N_7508,N_5151);
nor U13680 (N_13680,N_7240,N_9688);
nand U13681 (N_13681,N_9260,N_9592);
nand U13682 (N_13682,N_7818,N_8603);
or U13683 (N_13683,N_5989,N_6726);
nor U13684 (N_13684,N_7192,N_5967);
nor U13685 (N_13685,N_8188,N_9973);
xnor U13686 (N_13686,N_8360,N_8477);
or U13687 (N_13687,N_7038,N_5697);
and U13688 (N_13688,N_5974,N_9027);
and U13689 (N_13689,N_6072,N_9867);
and U13690 (N_13690,N_9990,N_6074);
nor U13691 (N_13691,N_9267,N_7071);
and U13692 (N_13692,N_7182,N_5122);
nor U13693 (N_13693,N_9852,N_7901);
or U13694 (N_13694,N_9453,N_9821);
or U13695 (N_13695,N_8059,N_9180);
nor U13696 (N_13696,N_6648,N_8336);
nor U13697 (N_13697,N_5436,N_8960);
and U13698 (N_13698,N_8794,N_9592);
nor U13699 (N_13699,N_6961,N_8437);
nand U13700 (N_13700,N_5733,N_5633);
nand U13701 (N_13701,N_7374,N_6152);
and U13702 (N_13702,N_5556,N_7793);
nor U13703 (N_13703,N_9701,N_7795);
nor U13704 (N_13704,N_5370,N_6062);
and U13705 (N_13705,N_9835,N_5358);
nand U13706 (N_13706,N_6614,N_7549);
xnor U13707 (N_13707,N_5725,N_9427);
and U13708 (N_13708,N_9020,N_9584);
or U13709 (N_13709,N_9992,N_9124);
nand U13710 (N_13710,N_6415,N_6195);
nor U13711 (N_13711,N_9594,N_6943);
xnor U13712 (N_13712,N_5099,N_9050);
nor U13713 (N_13713,N_6612,N_8788);
and U13714 (N_13714,N_7617,N_5607);
or U13715 (N_13715,N_5442,N_9394);
nand U13716 (N_13716,N_7789,N_8717);
nor U13717 (N_13717,N_6085,N_8721);
and U13718 (N_13718,N_6238,N_7907);
and U13719 (N_13719,N_5507,N_9000);
nor U13720 (N_13720,N_9956,N_8085);
nor U13721 (N_13721,N_9092,N_5150);
or U13722 (N_13722,N_6839,N_6501);
or U13723 (N_13723,N_6071,N_5663);
nor U13724 (N_13724,N_9016,N_7280);
nand U13725 (N_13725,N_5762,N_5949);
or U13726 (N_13726,N_6364,N_7095);
xnor U13727 (N_13727,N_5489,N_8286);
or U13728 (N_13728,N_5500,N_7430);
and U13729 (N_13729,N_6694,N_9871);
and U13730 (N_13730,N_7132,N_8222);
or U13731 (N_13731,N_6083,N_9686);
nand U13732 (N_13732,N_6369,N_6996);
nor U13733 (N_13733,N_7744,N_6340);
nand U13734 (N_13734,N_6969,N_8892);
xnor U13735 (N_13735,N_8259,N_8971);
nand U13736 (N_13736,N_8198,N_9182);
and U13737 (N_13737,N_7666,N_9015);
nor U13738 (N_13738,N_8223,N_7697);
nor U13739 (N_13739,N_9399,N_6458);
nor U13740 (N_13740,N_8495,N_9353);
xor U13741 (N_13741,N_6928,N_8213);
and U13742 (N_13742,N_8096,N_9525);
xnor U13743 (N_13743,N_9900,N_5340);
and U13744 (N_13744,N_9818,N_9324);
or U13745 (N_13745,N_9481,N_9582);
nor U13746 (N_13746,N_8744,N_6163);
nand U13747 (N_13747,N_7819,N_6485);
xor U13748 (N_13748,N_8882,N_6410);
or U13749 (N_13749,N_8508,N_5525);
xnor U13750 (N_13750,N_9473,N_8067);
xnor U13751 (N_13751,N_7052,N_5672);
nand U13752 (N_13752,N_6005,N_7386);
xnor U13753 (N_13753,N_8217,N_7204);
or U13754 (N_13754,N_9917,N_6961);
nor U13755 (N_13755,N_5670,N_8255);
nand U13756 (N_13756,N_5122,N_6452);
nor U13757 (N_13757,N_5735,N_5250);
or U13758 (N_13758,N_6179,N_7521);
and U13759 (N_13759,N_9076,N_8741);
and U13760 (N_13760,N_5107,N_7681);
and U13761 (N_13761,N_8160,N_5262);
nor U13762 (N_13762,N_6982,N_5778);
xor U13763 (N_13763,N_6221,N_8061);
or U13764 (N_13764,N_6892,N_8505);
or U13765 (N_13765,N_5583,N_5337);
nand U13766 (N_13766,N_8692,N_7434);
nor U13767 (N_13767,N_6440,N_9453);
xor U13768 (N_13768,N_7725,N_5727);
xor U13769 (N_13769,N_8246,N_9823);
nor U13770 (N_13770,N_6901,N_9851);
or U13771 (N_13771,N_8665,N_8336);
xor U13772 (N_13772,N_8033,N_7725);
nor U13773 (N_13773,N_8803,N_8488);
and U13774 (N_13774,N_7014,N_6888);
nand U13775 (N_13775,N_9655,N_7861);
and U13776 (N_13776,N_8722,N_8644);
and U13777 (N_13777,N_9909,N_9404);
xnor U13778 (N_13778,N_5661,N_7765);
xnor U13779 (N_13779,N_9397,N_7947);
or U13780 (N_13780,N_5600,N_7606);
and U13781 (N_13781,N_6428,N_9384);
xor U13782 (N_13782,N_5858,N_5329);
and U13783 (N_13783,N_9426,N_7431);
nand U13784 (N_13784,N_9804,N_9889);
nand U13785 (N_13785,N_5250,N_9726);
and U13786 (N_13786,N_5650,N_9400);
or U13787 (N_13787,N_5985,N_5202);
or U13788 (N_13788,N_6171,N_8617);
nor U13789 (N_13789,N_5089,N_8743);
and U13790 (N_13790,N_6414,N_8397);
nand U13791 (N_13791,N_6740,N_8516);
or U13792 (N_13792,N_6130,N_6117);
nand U13793 (N_13793,N_5772,N_8085);
and U13794 (N_13794,N_9656,N_8157);
nor U13795 (N_13795,N_7898,N_9254);
and U13796 (N_13796,N_5075,N_7123);
nor U13797 (N_13797,N_7468,N_6423);
xnor U13798 (N_13798,N_5446,N_9595);
nor U13799 (N_13799,N_7635,N_6195);
xnor U13800 (N_13800,N_6536,N_9411);
nor U13801 (N_13801,N_6241,N_6663);
nand U13802 (N_13802,N_8332,N_8286);
nor U13803 (N_13803,N_9351,N_6181);
or U13804 (N_13804,N_9730,N_9909);
nand U13805 (N_13805,N_9450,N_9506);
and U13806 (N_13806,N_7564,N_9991);
xor U13807 (N_13807,N_9610,N_6314);
xor U13808 (N_13808,N_7028,N_8626);
nor U13809 (N_13809,N_8768,N_8015);
nor U13810 (N_13810,N_7660,N_6383);
and U13811 (N_13811,N_8945,N_5854);
nand U13812 (N_13812,N_6755,N_9075);
xnor U13813 (N_13813,N_7918,N_7400);
xnor U13814 (N_13814,N_7063,N_6941);
xor U13815 (N_13815,N_8864,N_7704);
or U13816 (N_13816,N_6484,N_6896);
nor U13817 (N_13817,N_7210,N_9404);
and U13818 (N_13818,N_6821,N_8216);
and U13819 (N_13819,N_9251,N_8367);
and U13820 (N_13820,N_6100,N_6075);
nand U13821 (N_13821,N_7299,N_8946);
nand U13822 (N_13822,N_7536,N_5809);
xnor U13823 (N_13823,N_9362,N_9505);
and U13824 (N_13824,N_6734,N_8845);
and U13825 (N_13825,N_6664,N_9568);
xnor U13826 (N_13826,N_7360,N_8572);
nor U13827 (N_13827,N_7940,N_9418);
xor U13828 (N_13828,N_8992,N_8568);
nor U13829 (N_13829,N_8741,N_6421);
and U13830 (N_13830,N_7789,N_6872);
and U13831 (N_13831,N_9500,N_7951);
or U13832 (N_13832,N_9025,N_8660);
nand U13833 (N_13833,N_8593,N_8213);
and U13834 (N_13834,N_7342,N_7899);
nand U13835 (N_13835,N_6510,N_7629);
nor U13836 (N_13836,N_5355,N_8934);
xor U13837 (N_13837,N_6107,N_5629);
and U13838 (N_13838,N_9308,N_5233);
or U13839 (N_13839,N_6768,N_9286);
or U13840 (N_13840,N_8661,N_7378);
xnor U13841 (N_13841,N_9572,N_9898);
and U13842 (N_13842,N_7230,N_9857);
nor U13843 (N_13843,N_8626,N_6451);
xor U13844 (N_13844,N_5464,N_5874);
or U13845 (N_13845,N_9102,N_5383);
or U13846 (N_13846,N_9810,N_6857);
and U13847 (N_13847,N_7824,N_9212);
nand U13848 (N_13848,N_9254,N_7914);
xor U13849 (N_13849,N_9242,N_6143);
nand U13850 (N_13850,N_7391,N_8884);
and U13851 (N_13851,N_5965,N_6008);
xnor U13852 (N_13852,N_6026,N_8509);
nand U13853 (N_13853,N_6449,N_7320);
or U13854 (N_13854,N_7375,N_8712);
and U13855 (N_13855,N_5345,N_5061);
xor U13856 (N_13856,N_7971,N_6122);
or U13857 (N_13857,N_5541,N_5208);
and U13858 (N_13858,N_7060,N_5865);
or U13859 (N_13859,N_6968,N_5365);
nand U13860 (N_13860,N_6188,N_6771);
and U13861 (N_13861,N_5451,N_6584);
and U13862 (N_13862,N_5548,N_5782);
and U13863 (N_13863,N_8284,N_9298);
nor U13864 (N_13864,N_7791,N_5125);
and U13865 (N_13865,N_6435,N_6294);
and U13866 (N_13866,N_9764,N_8497);
and U13867 (N_13867,N_5778,N_7836);
or U13868 (N_13868,N_5431,N_7697);
nor U13869 (N_13869,N_7388,N_9484);
nand U13870 (N_13870,N_9151,N_7251);
nor U13871 (N_13871,N_8618,N_5345);
nor U13872 (N_13872,N_8370,N_6393);
and U13873 (N_13873,N_8714,N_9719);
and U13874 (N_13874,N_9893,N_6647);
and U13875 (N_13875,N_5106,N_8007);
and U13876 (N_13876,N_5550,N_5247);
or U13877 (N_13877,N_6858,N_8195);
xor U13878 (N_13878,N_7840,N_9222);
nand U13879 (N_13879,N_8851,N_7921);
nor U13880 (N_13880,N_6755,N_5135);
and U13881 (N_13881,N_9162,N_7668);
or U13882 (N_13882,N_9026,N_9202);
and U13883 (N_13883,N_7402,N_6974);
or U13884 (N_13884,N_8592,N_7299);
xnor U13885 (N_13885,N_8591,N_7393);
or U13886 (N_13886,N_9272,N_6411);
nand U13887 (N_13887,N_6263,N_8893);
nand U13888 (N_13888,N_5566,N_6302);
nand U13889 (N_13889,N_5193,N_5501);
nor U13890 (N_13890,N_8849,N_9917);
or U13891 (N_13891,N_5421,N_8424);
or U13892 (N_13892,N_6320,N_8992);
and U13893 (N_13893,N_9979,N_6833);
or U13894 (N_13894,N_9819,N_6242);
and U13895 (N_13895,N_8766,N_5059);
xnor U13896 (N_13896,N_5980,N_5829);
xor U13897 (N_13897,N_7542,N_6006);
xnor U13898 (N_13898,N_8846,N_7329);
or U13899 (N_13899,N_5162,N_8468);
nand U13900 (N_13900,N_8617,N_6692);
xnor U13901 (N_13901,N_9291,N_9818);
or U13902 (N_13902,N_9620,N_7192);
and U13903 (N_13903,N_7019,N_6138);
xnor U13904 (N_13904,N_7275,N_8796);
nor U13905 (N_13905,N_6564,N_8041);
xor U13906 (N_13906,N_9749,N_8681);
and U13907 (N_13907,N_6448,N_7264);
nor U13908 (N_13908,N_7143,N_6878);
or U13909 (N_13909,N_5387,N_6993);
xnor U13910 (N_13910,N_6744,N_9758);
nor U13911 (N_13911,N_7097,N_5351);
and U13912 (N_13912,N_8771,N_9784);
and U13913 (N_13913,N_9736,N_8787);
xnor U13914 (N_13914,N_6385,N_5440);
or U13915 (N_13915,N_7214,N_9808);
xnor U13916 (N_13916,N_6445,N_6841);
nor U13917 (N_13917,N_5246,N_9938);
or U13918 (N_13918,N_9162,N_6756);
nand U13919 (N_13919,N_6918,N_9993);
nor U13920 (N_13920,N_9609,N_5321);
nor U13921 (N_13921,N_6434,N_8482);
and U13922 (N_13922,N_6399,N_6106);
and U13923 (N_13923,N_6155,N_6843);
or U13924 (N_13924,N_6600,N_5024);
nand U13925 (N_13925,N_5675,N_9336);
and U13926 (N_13926,N_5300,N_6596);
and U13927 (N_13927,N_5826,N_5527);
and U13928 (N_13928,N_5444,N_6429);
xor U13929 (N_13929,N_6435,N_7059);
nand U13930 (N_13930,N_9514,N_9849);
and U13931 (N_13931,N_8212,N_7164);
or U13932 (N_13932,N_8743,N_8849);
nor U13933 (N_13933,N_9569,N_6463);
nand U13934 (N_13934,N_7561,N_8354);
nor U13935 (N_13935,N_5398,N_7289);
xnor U13936 (N_13936,N_9577,N_5442);
and U13937 (N_13937,N_9233,N_9893);
and U13938 (N_13938,N_6732,N_7330);
xnor U13939 (N_13939,N_7401,N_7694);
and U13940 (N_13940,N_8975,N_9550);
and U13941 (N_13941,N_6283,N_7815);
and U13942 (N_13942,N_5117,N_8527);
and U13943 (N_13943,N_5291,N_7111);
nand U13944 (N_13944,N_9875,N_5302);
or U13945 (N_13945,N_5185,N_9105);
or U13946 (N_13946,N_6017,N_9856);
or U13947 (N_13947,N_9588,N_5041);
nand U13948 (N_13948,N_9562,N_7231);
nand U13949 (N_13949,N_8017,N_7282);
and U13950 (N_13950,N_5569,N_8479);
and U13951 (N_13951,N_6333,N_7206);
and U13952 (N_13952,N_6380,N_7198);
or U13953 (N_13953,N_7837,N_6928);
or U13954 (N_13954,N_5686,N_7516);
xor U13955 (N_13955,N_6666,N_9546);
xnor U13956 (N_13956,N_9553,N_6350);
or U13957 (N_13957,N_8915,N_6454);
xor U13958 (N_13958,N_9244,N_8228);
nand U13959 (N_13959,N_5261,N_8169);
nand U13960 (N_13960,N_8490,N_6473);
nor U13961 (N_13961,N_6634,N_7503);
nand U13962 (N_13962,N_6379,N_9333);
nand U13963 (N_13963,N_5317,N_7310);
nand U13964 (N_13964,N_8240,N_6856);
nand U13965 (N_13965,N_7549,N_7079);
xnor U13966 (N_13966,N_9379,N_6878);
or U13967 (N_13967,N_5377,N_9752);
nor U13968 (N_13968,N_8172,N_9980);
xnor U13969 (N_13969,N_9457,N_8735);
nand U13970 (N_13970,N_5096,N_7040);
nor U13971 (N_13971,N_7713,N_5491);
xnor U13972 (N_13972,N_9414,N_8127);
nor U13973 (N_13973,N_5548,N_9140);
or U13974 (N_13974,N_9415,N_9959);
xor U13975 (N_13975,N_5774,N_7051);
nand U13976 (N_13976,N_5788,N_5540);
and U13977 (N_13977,N_5494,N_8978);
or U13978 (N_13978,N_8923,N_5546);
nand U13979 (N_13979,N_5968,N_7233);
xor U13980 (N_13980,N_5555,N_8490);
xnor U13981 (N_13981,N_9033,N_9684);
and U13982 (N_13982,N_8047,N_5047);
or U13983 (N_13983,N_6645,N_8627);
or U13984 (N_13984,N_7531,N_6880);
and U13985 (N_13985,N_7270,N_9135);
xnor U13986 (N_13986,N_6277,N_5900);
xnor U13987 (N_13987,N_8841,N_7549);
xnor U13988 (N_13988,N_9317,N_9488);
and U13989 (N_13989,N_5302,N_5764);
nor U13990 (N_13990,N_7826,N_8382);
or U13991 (N_13991,N_8248,N_6797);
and U13992 (N_13992,N_8709,N_7779);
or U13993 (N_13993,N_7222,N_9957);
xor U13994 (N_13994,N_5193,N_7112);
and U13995 (N_13995,N_8880,N_9337);
xnor U13996 (N_13996,N_8330,N_6449);
xnor U13997 (N_13997,N_8243,N_5610);
nand U13998 (N_13998,N_5096,N_9029);
xor U13999 (N_13999,N_5917,N_6947);
xnor U14000 (N_14000,N_9852,N_8733);
and U14001 (N_14001,N_7816,N_8892);
nand U14002 (N_14002,N_9061,N_9706);
and U14003 (N_14003,N_7398,N_5868);
or U14004 (N_14004,N_7379,N_9714);
and U14005 (N_14005,N_9749,N_8840);
nand U14006 (N_14006,N_8729,N_9477);
nand U14007 (N_14007,N_5232,N_9700);
and U14008 (N_14008,N_5272,N_8299);
nand U14009 (N_14009,N_6927,N_8871);
nand U14010 (N_14010,N_8098,N_6189);
nor U14011 (N_14011,N_7833,N_7936);
nor U14012 (N_14012,N_7680,N_6628);
and U14013 (N_14013,N_6294,N_7015);
nand U14014 (N_14014,N_8541,N_6441);
xor U14015 (N_14015,N_6477,N_7486);
nand U14016 (N_14016,N_9290,N_8630);
nand U14017 (N_14017,N_5448,N_7847);
and U14018 (N_14018,N_7721,N_8184);
xor U14019 (N_14019,N_6352,N_6595);
xnor U14020 (N_14020,N_7793,N_7101);
nor U14021 (N_14021,N_9631,N_6576);
nor U14022 (N_14022,N_9079,N_6210);
or U14023 (N_14023,N_6539,N_8521);
nor U14024 (N_14024,N_7423,N_5943);
nor U14025 (N_14025,N_6143,N_9007);
nand U14026 (N_14026,N_6381,N_7074);
nor U14027 (N_14027,N_7299,N_9708);
nand U14028 (N_14028,N_5499,N_9143);
or U14029 (N_14029,N_6998,N_8796);
nand U14030 (N_14030,N_5899,N_9285);
or U14031 (N_14031,N_9798,N_7144);
or U14032 (N_14032,N_7231,N_9777);
nand U14033 (N_14033,N_8711,N_5713);
and U14034 (N_14034,N_8333,N_8164);
or U14035 (N_14035,N_7764,N_5003);
nor U14036 (N_14036,N_5728,N_6066);
xnor U14037 (N_14037,N_9030,N_5827);
xor U14038 (N_14038,N_8804,N_6411);
or U14039 (N_14039,N_5655,N_9018);
and U14040 (N_14040,N_7047,N_9368);
nand U14041 (N_14041,N_7444,N_6043);
or U14042 (N_14042,N_5312,N_8721);
and U14043 (N_14043,N_8632,N_6403);
nor U14044 (N_14044,N_8399,N_9248);
nand U14045 (N_14045,N_6069,N_5285);
and U14046 (N_14046,N_9624,N_5406);
xor U14047 (N_14047,N_5753,N_9648);
and U14048 (N_14048,N_8039,N_5937);
nand U14049 (N_14049,N_5574,N_5795);
xnor U14050 (N_14050,N_5619,N_8849);
or U14051 (N_14051,N_7882,N_7087);
nor U14052 (N_14052,N_6526,N_8889);
nor U14053 (N_14053,N_6102,N_5208);
and U14054 (N_14054,N_5928,N_5890);
nor U14055 (N_14055,N_6622,N_5891);
or U14056 (N_14056,N_6665,N_5919);
nand U14057 (N_14057,N_9503,N_5003);
and U14058 (N_14058,N_8912,N_8577);
or U14059 (N_14059,N_6225,N_6433);
xor U14060 (N_14060,N_6850,N_5483);
nor U14061 (N_14061,N_8667,N_5777);
and U14062 (N_14062,N_6415,N_7784);
nand U14063 (N_14063,N_9854,N_7730);
or U14064 (N_14064,N_5798,N_6989);
or U14065 (N_14065,N_6910,N_5453);
nand U14066 (N_14066,N_5499,N_6278);
or U14067 (N_14067,N_6420,N_6311);
nand U14068 (N_14068,N_6155,N_5918);
and U14069 (N_14069,N_6994,N_8385);
nand U14070 (N_14070,N_5656,N_7660);
and U14071 (N_14071,N_6886,N_6844);
or U14072 (N_14072,N_6444,N_8752);
nor U14073 (N_14073,N_9664,N_9382);
or U14074 (N_14074,N_5888,N_7370);
xnor U14075 (N_14075,N_5282,N_5832);
or U14076 (N_14076,N_8913,N_6523);
and U14077 (N_14077,N_7654,N_6352);
xor U14078 (N_14078,N_8295,N_7391);
nor U14079 (N_14079,N_6967,N_8866);
xnor U14080 (N_14080,N_8914,N_5987);
nor U14081 (N_14081,N_7794,N_5781);
and U14082 (N_14082,N_7831,N_8859);
nor U14083 (N_14083,N_5605,N_9802);
xnor U14084 (N_14084,N_9011,N_5517);
or U14085 (N_14085,N_8129,N_8740);
xor U14086 (N_14086,N_6006,N_7215);
and U14087 (N_14087,N_5254,N_7840);
nor U14088 (N_14088,N_8123,N_8628);
xor U14089 (N_14089,N_7104,N_9263);
xor U14090 (N_14090,N_5061,N_7358);
or U14091 (N_14091,N_8796,N_5495);
xor U14092 (N_14092,N_6294,N_7655);
xor U14093 (N_14093,N_9758,N_5276);
nand U14094 (N_14094,N_6915,N_7082);
nand U14095 (N_14095,N_6940,N_8968);
and U14096 (N_14096,N_8895,N_9077);
xnor U14097 (N_14097,N_9912,N_7886);
and U14098 (N_14098,N_5042,N_8862);
or U14099 (N_14099,N_5103,N_9219);
nor U14100 (N_14100,N_5538,N_5097);
nor U14101 (N_14101,N_5543,N_7734);
nor U14102 (N_14102,N_5610,N_6904);
or U14103 (N_14103,N_8241,N_5429);
nor U14104 (N_14104,N_7387,N_9095);
nand U14105 (N_14105,N_8127,N_8419);
xor U14106 (N_14106,N_9512,N_5861);
and U14107 (N_14107,N_9904,N_7299);
nor U14108 (N_14108,N_8949,N_7765);
xor U14109 (N_14109,N_7767,N_8662);
xor U14110 (N_14110,N_7282,N_9793);
nor U14111 (N_14111,N_6329,N_5814);
and U14112 (N_14112,N_8153,N_6591);
and U14113 (N_14113,N_7466,N_5027);
or U14114 (N_14114,N_9220,N_5802);
or U14115 (N_14115,N_7139,N_8619);
xor U14116 (N_14116,N_6382,N_7465);
xor U14117 (N_14117,N_9907,N_9912);
nor U14118 (N_14118,N_8357,N_5360);
nor U14119 (N_14119,N_8725,N_6419);
xor U14120 (N_14120,N_7469,N_8791);
nor U14121 (N_14121,N_6023,N_9514);
and U14122 (N_14122,N_7899,N_8984);
or U14123 (N_14123,N_8526,N_7513);
and U14124 (N_14124,N_8875,N_7671);
xor U14125 (N_14125,N_7719,N_7100);
or U14126 (N_14126,N_8838,N_8552);
xor U14127 (N_14127,N_9507,N_7911);
or U14128 (N_14128,N_5546,N_8438);
or U14129 (N_14129,N_9096,N_6475);
and U14130 (N_14130,N_8569,N_6489);
nor U14131 (N_14131,N_5232,N_5368);
xnor U14132 (N_14132,N_5932,N_8612);
nor U14133 (N_14133,N_8264,N_9796);
xnor U14134 (N_14134,N_5283,N_7511);
or U14135 (N_14135,N_9402,N_6371);
and U14136 (N_14136,N_8543,N_6134);
nor U14137 (N_14137,N_8285,N_6078);
or U14138 (N_14138,N_9252,N_9460);
and U14139 (N_14139,N_8282,N_8181);
or U14140 (N_14140,N_7693,N_8140);
xor U14141 (N_14141,N_7977,N_9814);
xor U14142 (N_14142,N_7184,N_6119);
nand U14143 (N_14143,N_9285,N_7376);
nand U14144 (N_14144,N_5806,N_8791);
nand U14145 (N_14145,N_7372,N_9824);
and U14146 (N_14146,N_8273,N_9501);
xor U14147 (N_14147,N_6370,N_5012);
or U14148 (N_14148,N_8820,N_9247);
nor U14149 (N_14149,N_6496,N_9417);
and U14150 (N_14150,N_7072,N_8073);
nand U14151 (N_14151,N_6825,N_5210);
and U14152 (N_14152,N_5194,N_8275);
nor U14153 (N_14153,N_7693,N_7609);
and U14154 (N_14154,N_9606,N_6102);
nand U14155 (N_14155,N_5384,N_5162);
or U14156 (N_14156,N_7551,N_6399);
and U14157 (N_14157,N_9821,N_8194);
or U14158 (N_14158,N_8393,N_5420);
and U14159 (N_14159,N_8445,N_5151);
nor U14160 (N_14160,N_7951,N_9505);
xnor U14161 (N_14161,N_6871,N_9589);
or U14162 (N_14162,N_7430,N_8399);
or U14163 (N_14163,N_6853,N_9287);
xnor U14164 (N_14164,N_5071,N_7737);
xor U14165 (N_14165,N_5710,N_5022);
nand U14166 (N_14166,N_5386,N_5615);
nand U14167 (N_14167,N_5183,N_7173);
xnor U14168 (N_14168,N_7565,N_8393);
nor U14169 (N_14169,N_7584,N_9154);
nand U14170 (N_14170,N_9735,N_7978);
and U14171 (N_14171,N_7778,N_7456);
nor U14172 (N_14172,N_9782,N_9120);
nor U14173 (N_14173,N_8345,N_9508);
nor U14174 (N_14174,N_9913,N_6044);
xor U14175 (N_14175,N_7380,N_9777);
xor U14176 (N_14176,N_9164,N_8266);
or U14177 (N_14177,N_8899,N_9705);
nand U14178 (N_14178,N_7757,N_7206);
xnor U14179 (N_14179,N_7917,N_5727);
nor U14180 (N_14180,N_5636,N_8342);
xor U14181 (N_14181,N_9748,N_9107);
xnor U14182 (N_14182,N_7418,N_8622);
nand U14183 (N_14183,N_7834,N_7186);
or U14184 (N_14184,N_5755,N_5600);
nand U14185 (N_14185,N_8630,N_9976);
nand U14186 (N_14186,N_8675,N_5147);
nor U14187 (N_14187,N_7819,N_5230);
and U14188 (N_14188,N_8731,N_5100);
or U14189 (N_14189,N_9298,N_6313);
nor U14190 (N_14190,N_6516,N_7562);
and U14191 (N_14191,N_6380,N_9385);
and U14192 (N_14192,N_6943,N_9670);
nand U14193 (N_14193,N_6012,N_8168);
and U14194 (N_14194,N_5311,N_7860);
xnor U14195 (N_14195,N_7977,N_6856);
nand U14196 (N_14196,N_8500,N_5416);
nand U14197 (N_14197,N_9991,N_7143);
and U14198 (N_14198,N_7227,N_6023);
xnor U14199 (N_14199,N_9181,N_8155);
nand U14200 (N_14200,N_9767,N_7727);
nand U14201 (N_14201,N_5570,N_9643);
and U14202 (N_14202,N_9288,N_6549);
nor U14203 (N_14203,N_7668,N_5647);
nor U14204 (N_14204,N_8322,N_7363);
and U14205 (N_14205,N_6154,N_9125);
xnor U14206 (N_14206,N_8001,N_5035);
nor U14207 (N_14207,N_7255,N_5265);
or U14208 (N_14208,N_7061,N_8258);
xor U14209 (N_14209,N_5971,N_8315);
nor U14210 (N_14210,N_5687,N_5973);
nand U14211 (N_14211,N_6814,N_9534);
or U14212 (N_14212,N_8855,N_9250);
or U14213 (N_14213,N_6244,N_8635);
xnor U14214 (N_14214,N_7954,N_8656);
nand U14215 (N_14215,N_5061,N_5393);
or U14216 (N_14216,N_8877,N_7397);
xnor U14217 (N_14217,N_8337,N_9922);
nor U14218 (N_14218,N_5101,N_9694);
or U14219 (N_14219,N_5268,N_9416);
xor U14220 (N_14220,N_5089,N_8319);
nand U14221 (N_14221,N_5806,N_7433);
nor U14222 (N_14222,N_7938,N_5488);
xor U14223 (N_14223,N_7528,N_8229);
and U14224 (N_14224,N_5513,N_7192);
nand U14225 (N_14225,N_8137,N_6531);
or U14226 (N_14226,N_6523,N_6279);
nor U14227 (N_14227,N_8425,N_6471);
and U14228 (N_14228,N_6230,N_7950);
or U14229 (N_14229,N_9337,N_6265);
nand U14230 (N_14230,N_5700,N_6844);
xor U14231 (N_14231,N_8254,N_5850);
or U14232 (N_14232,N_9105,N_5929);
nand U14233 (N_14233,N_9520,N_7275);
nand U14234 (N_14234,N_7263,N_8391);
xnor U14235 (N_14235,N_7211,N_8326);
and U14236 (N_14236,N_6921,N_7469);
and U14237 (N_14237,N_9726,N_8059);
nand U14238 (N_14238,N_7441,N_6376);
xnor U14239 (N_14239,N_7084,N_7083);
and U14240 (N_14240,N_9385,N_8949);
nor U14241 (N_14241,N_9300,N_8443);
xor U14242 (N_14242,N_7336,N_5802);
or U14243 (N_14243,N_9717,N_6550);
nor U14244 (N_14244,N_8929,N_9555);
nand U14245 (N_14245,N_9167,N_5150);
xor U14246 (N_14246,N_7993,N_7563);
nand U14247 (N_14247,N_6006,N_8078);
nor U14248 (N_14248,N_6366,N_7561);
or U14249 (N_14249,N_6982,N_7426);
nor U14250 (N_14250,N_7036,N_9386);
and U14251 (N_14251,N_8914,N_8218);
nand U14252 (N_14252,N_5797,N_7917);
nand U14253 (N_14253,N_7488,N_6930);
xor U14254 (N_14254,N_8881,N_7458);
xor U14255 (N_14255,N_7889,N_8551);
xnor U14256 (N_14256,N_5415,N_5226);
nor U14257 (N_14257,N_9162,N_9431);
nor U14258 (N_14258,N_8437,N_5323);
nor U14259 (N_14259,N_7987,N_8329);
nor U14260 (N_14260,N_9500,N_5275);
xor U14261 (N_14261,N_8626,N_9272);
nand U14262 (N_14262,N_9818,N_8105);
and U14263 (N_14263,N_8721,N_6943);
and U14264 (N_14264,N_7090,N_5926);
and U14265 (N_14265,N_5976,N_5484);
nor U14266 (N_14266,N_9952,N_6221);
or U14267 (N_14267,N_5185,N_6484);
or U14268 (N_14268,N_8283,N_5236);
xnor U14269 (N_14269,N_8326,N_8145);
xor U14270 (N_14270,N_8796,N_9438);
nand U14271 (N_14271,N_8951,N_6082);
nand U14272 (N_14272,N_6502,N_6934);
nor U14273 (N_14273,N_7673,N_7689);
nand U14274 (N_14274,N_5179,N_9824);
nor U14275 (N_14275,N_8126,N_5424);
xor U14276 (N_14276,N_5771,N_6993);
nor U14277 (N_14277,N_9582,N_6684);
or U14278 (N_14278,N_5079,N_9325);
or U14279 (N_14279,N_5729,N_5062);
nand U14280 (N_14280,N_8989,N_6619);
xor U14281 (N_14281,N_8804,N_7051);
and U14282 (N_14282,N_7492,N_6986);
nor U14283 (N_14283,N_6708,N_7360);
nor U14284 (N_14284,N_7506,N_6271);
nor U14285 (N_14285,N_8909,N_6765);
and U14286 (N_14286,N_9986,N_7187);
nand U14287 (N_14287,N_9361,N_7567);
xor U14288 (N_14288,N_8487,N_5559);
xor U14289 (N_14289,N_6771,N_9185);
nand U14290 (N_14290,N_6419,N_9162);
nand U14291 (N_14291,N_9925,N_5511);
xnor U14292 (N_14292,N_7787,N_7124);
or U14293 (N_14293,N_5916,N_5245);
nor U14294 (N_14294,N_7104,N_6623);
xor U14295 (N_14295,N_8038,N_7413);
and U14296 (N_14296,N_8596,N_6406);
xor U14297 (N_14297,N_7952,N_8591);
or U14298 (N_14298,N_9146,N_6596);
and U14299 (N_14299,N_6557,N_9745);
xnor U14300 (N_14300,N_7114,N_9134);
nand U14301 (N_14301,N_5259,N_6507);
xor U14302 (N_14302,N_9128,N_6216);
nor U14303 (N_14303,N_7569,N_6321);
nor U14304 (N_14304,N_7084,N_9412);
nand U14305 (N_14305,N_9823,N_7162);
nand U14306 (N_14306,N_5322,N_5980);
nand U14307 (N_14307,N_7562,N_6409);
and U14308 (N_14308,N_5758,N_7663);
nor U14309 (N_14309,N_8295,N_8495);
nand U14310 (N_14310,N_8129,N_5581);
xnor U14311 (N_14311,N_6170,N_8876);
xor U14312 (N_14312,N_5198,N_8593);
nand U14313 (N_14313,N_9113,N_7591);
or U14314 (N_14314,N_8176,N_8362);
nor U14315 (N_14315,N_7119,N_5409);
xnor U14316 (N_14316,N_6468,N_8879);
xor U14317 (N_14317,N_9586,N_8286);
and U14318 (N_14318,N_6294,N_7014);
nor U14319 (N_14319,N_8843,N_6377);
or U14320 (N_14320,N_7129,N_6035);
or U14321 (N_14321,N_5632,N_7608);
or U14322 (N_14322,N_8641,N_6591);
xor U14323 (N_14323,N_6515,N_9127);
or U14324 (N_14324,N_7183,N_9583);
nand U14325 (N_14325,N_9169,N_9966);
nor U14326 (N_14326,N_6269,N_8009);
nand U14327 (N_14327,N_9070,N_6244);
and U14328 (N_14328,N_9183,N_5272);
nor U14329 (N_14329,N_5346,N_9123);
nor U14330 (N_14330,N_8829,N_5558);
and U14331 (N_14331,N_5238,N_7291);
or U14332 (N_14332,N_7204,N_5230);
xnor U14333 (N_14333,N_9041,N_5334);
or U14334 (N_14334,N_8304,N_7312);
and U14335 (N_14335,N_9048,N_7509);
nand U14336 (N_14336,N_5356,N_8351);
nand U14337 (N_14337,N_7349,N_5936);
xnor U14338 (N_14338,N_5649,N_6383);
or U14339 (N_14339,N_6542,N_8982);
and U14340 (N_14340,N_8378,N_8089);
nor U14341 (N_14341,N_8326,N_7759);
or U14342 (N_14342,N_7441,N_5854);
xor U14343 (N_14343,N_7737,N_8251);
xnor U14344 (N_14344,N_7018,N_9876);
xor U14345 (N_14345,N_9215,N_6658);
xor U14346 (N_14346,N_9142,N_8221);
or U14347 (N_14347,N_8820,N_5143);
xnor U14348 (N_14348,N_9950,N_5245);
and U14349 (N_14349,N_8998,N_8714);
and U14350 (N_14350,N_9826,N_9227);
nor U14351 (N_14351,N_7173,N_6786);
xnor U14352 (N_14352,N_9627,N_6167);
nor U14353 (N_14353,N_5294,N_5434);
nand U14354 (N_14354,N_5563,N_7593);
or U14355 (N_14355,N_6613,N_9095);
nor U14356 (N_14356,N_9494,N_9004);
and U14357 (N_14357,N_9931,N_5302);
and U14358 (N_14358,N_6741,N_5514);
and U14359 (N_14359,N_6706,N_7877);
xnor U14360 (N_14360,N_6501,N_6980);
xor U14361 (N_14361,N_8563,N_5324);
nand U14362 (N_14362,N_7804,N_7748);
xor U14363 (N_14363,N_7089,N_5138);
xor U14364 (N_14364,N_5842,N_8315);
nor U14365 (N_14365,N_6709,N_9035);
or U14366 (N_14366,N_6421,N_9890);
nor U14367 (N_14367,N_6663,N_5594);
nand U14368 (N_14368,N_9648,N_6323);
or U14369 (N_14369,N_6860,N_6555);
and U14370 (N_14370,N_8389,N_7015);
xnor U14371 (N_14371,N_7244,N_5652);
or U14372 (N_14372,N_6734,N_8469);
nand U14373 (N_14373,N_6000,N_9994);
or U14374 (N_14374,N_7862,N_7993);
nand U14375 (N_14375,N_8658,N_9395);
or U14376 (N_14376,N_9783,N_6559);
or U14377 (N_14377,N_7637,N_5426);
nor U14378 (N_14378,N_9847,N_7856);
nand U14379 (N_14379,N_6088,N_7697);
nor U14380 (N_14380,N_9681,N_7412);
or U14381 (N_14381,N_5516,N_9531);
or U14382 (N_14382,N_7480,N_6894);
nor U14383 (N_14383,N_7345,N_6143);
xor U14384 (N_14384,N_5599,N_5937);
nand U14385 (N_14385,N_6012,N_7822);
or U14386 (N_14386,N_9283,N_7030);
xnor U14387 (N_14387,N_7166,N_8945);
nand U14388 (N_14388,N_7198,N_9019);
or U14389 (N_14389,N_7481,N_9218);
nor U14390 (N_14390,N_7699,N_6118);
nand U14391 (N_14391,N_9624,N_6981);
or U14392 (N_14392,N_5384,N_5845);
or U14393 (N_14393,N_7317,N_6370);
nand U14394 (N_14394,N_8632,N_5873);
and U14395 (N_14395,N_7839,N_5103);
and U14396 (N_14396,N_9711,N_7505);
and U14397 (N_14397,N_6780,N_9470);
or U14398 (N_14398,N_9279,N_6669);
or U14399 (N_14399,N_5663,N_7510);
and U14400 (N_14400,N_9964,N_8795);
nand U14401 (N_14401,N_7599,N_8489);
xnor U14402 (N_14402,N_5817,N_7162);
nand U14403 (N_14403,N_7788,N_7813);
xor U14404 (N_14404,N_6758,N_9820);
nor U14405 (N_14405,N_7475,N_5707);
or U14406 (N_14406,N_5438,N_8685);
xor U14407 (N_14407,N_7127,N_6598);
and U14408 (N_14408,N_6846,N_8845);
or U14409 (N_14409,N_9468,N_5092);
nor U14410 (N_14410,N_6484,N_5320);
or U14411 (N_14411,N_9242,N_9871);
xnor U14412 (N_14412,N_8629,N_7960);
or U14413 (N_14413,N_7889,N_5080);
or U14414 (N_14414,N_9610,N_6982);
or U14415 (N_14415,N_6870,N_9448);
nand U14416 (N_14416,N_7247,N_8284);
nor U14417 (N_14417,N_8098,N_5209);
xnor U14418 (N_14418,N_9503,N_6242);
nand U14419 (N_14419,N_6305,N_6197);
nand U14420 (N_14420,N_6000,N_5136);
xor U14421 (N_14421,N_8270,N_7980);
xnor U14422 (N_14422,N_9183,N_8147);
xor U14423 (N_14423,N_6804,N_8075);
and U14424 (N_14424,N_5741,N_8978);
nor U14425 (N_14425,N_6147,N_6263);
nor U14426 (N_14426,N_9581,N_7215);
nand U14427 (N_14427,N_9385,N_7007);
xnor U14428 (N_14428,N_8005,N_9626);
or U14429 (N_14429,N_5947,N_8119);
nand U14430 (N_14430,N_9897,N_9888);
and U14431 (N_14431,N_5281,N_6528);
nand U14432 (N_14432,N_7917,N_5772);
nand U14433 (N_14433,N_6568,N_7382);
or U14434 (N_14434,N_6072,N_5741);
or U14435 (N_14435,N_5889,N_5368);
nand U14436 (N_14436,N_5306,N_9010);
and U14437 (N_14437,N_5814,N_5935);
or U14438 (N_14438,N_8140,N_6362);
or U14439 (N_14439,N_7218,N_8358);
and U14440 (N_14440,N_6843,N_5651);
nor U14441 (N_14441,N_6963,N_8388);
nand U14442 (N_14442,N_7566,N_6191);
and U14443 (N_14443,N_7164,N_6700);
xnor U14444 (N_14444,N_8948,N_8792);
or U14445 (N_14445,N_8371,N_9916);
or U14446 (N_14446,N_7750,N_7195);
or U14447 (N_14447,N_6566,N_9490);
nand U14448 (N_14448,N_9474,N_5064);
xor U14449 (N_14449,N_6027,N_9795);
nand U14450 (N_14450,N_5544,N_5957);
nand U14451 (N_14451,N_7035,N_9596);
xnor U14452 (N_14452,N_9495,N_9240);
and U14453 (N_14453,N_8927,N_7307);
or U14454 (N_14454,N_5589,N_9773);
and U14455 (N_14455,N_5302,N_6716);
xnor U14456 (N_14456,N_8881,N_5330);
and U14457 (N_14457,N_6105,N_7369);
nand U14458 (N_14458,N_6563,N_7076);
and U14459 (N_14459,N_6883,N_6170);
xnor U14460 (N_14460,N_8836,N_8725);
or U14461 (N_14461,N_6401,N_5913);
and U14462 (N_14462,N_8971,N_9526);
nor U14463 (N_14463,N_7730,N_6994);
nand U14464 (N_14464,N_8048,N_7008);
nor U14465 (N_14465,N_8863,N_7962);
and U14466 (N_14466,N_6614,N_8170);
and U14467 (N_14467,N_8899,N_7492);
and U14468 (N_14468,N_8150,N_6919);
xnor U14469 (N_14469,N_8101,N_9808);
nand U14470 (N_14470,N_7025,N_7982);
nand U14471 (N_14471,N_8780,N_6220);
xnor U14472 (N_14472,N_8663,N_7807);
or U14473 (N_14473,N_9212,N_7942);
xor U14474 (N_14474,N_7075,N_5690);
and U14475 (N_14475,N_7676,N_9712);
nor U14476 (N_14476,N_9112,N_6850);
xnor U14477 (N_14477,N_8609,N_9926);
xor U14478 (N_14478,N_7287,N_9802);
nand U14479 (N_14479,N_9571,N_5431);
nor U14480 (N_14480,N_7886,N_7564);
or U14481 (N_14481,N_8692,N_9225);
nand U14482 (N_14482,N_7743,N_8425);
xor U14483 (N_14483,N_8541,N_7457);
nor U14484 (N_14484,N_6019,N_5855);
nor U14485 (N_14485,N_8263,N_5634);
nand U14486 (N_14486,N_9919,N_9886);
xnor U14487 (N_14487,N_7439,N_5771);
or U14488 (N_14488,N_6476,N_8445);
xnor U14489 (N_14489,N_5486,N_6938);
nor U14490 (N_14490,N_6951,N_7096);
nor U14491 (N_14491,N_5449,N_7036);
and U14492 (N_14492,N_7427,N_5703);
nand U14493 (N_14493,N_7500,N_5021);
or U14494 (N_14494,N_6400,N_5785);
or U14495 (N_14495,N_9072,N_8083);
nand U14496 (N_14496,N_7098,N_6775);
nand U14497 (N_14497,N_8543,N_9390);
nor U14498 (N_14498,N_5122,N_5336);
xor U14499 (N_14499,N_6329,N_9645);
and U14500 (N_14500,N_6841,N_5938);
nand U14501 (N_14501,N_9636,N_9045);
nand U14502 (N_14502,N_7301,N_5303);
nor U14503 (N_14503,N_5814,N_5758);
or U14504 (N_14504,N_5012,N_9366);
nor U14505 (N_14505,N_7939,N_8889);
xnor U14506 (N_14506,N_9368,N_6397);
nor U14507 (N_14507,N_7927,N_9799);
nor U14508 (N_14508,N_7428,N_7595);
nand U14509 (N_14509,N_6306,N_7935);
and U14510 (N_14510,N_6642,N_8596);
and U14511 (N_14511,N_5768,N_6113);
nor U14512 (N_14512,N_6413,N_5949);
and U14513 (N_14513,N_7614,N_9980);
or U14514 (N_14514,N_6330,N_9696);
nor U14515 (N_14515,N_9908,N_7818);
xnor U14516 (N_14516,N_9120,N_5735);
xor U14517 (N_14517,N_7242,N_9063);
and U14518 (N_14518,N_5996,N_8415);
or U14519 (N_14519,N_5523,N_9786);
nand U14520 (N_14520,N_5346,N_6778);
nor U14521 (N_14521,N_8720,N_8518);
nor U14522 (N_14522,N_6640,N_5014);
and U14523 (N_14523,N_7999,N_9004);
and U14524 (N_14524,N_9465,N_9577);
and U14525 (N_14525,N_7658,N_9471);
nand U14526 (N_14526,N_5795,N_8316);
xor U14527 (N_14527,N_6719,N_9108);
xor U14528 (N_14528,N_7281,N_6635);
nor U14529 (N_14529,N_5288,N_8687);
nor U14530 (N_14530,N_5678,N_8888);
and U14531 (N_14531,N_5357,N_7211);
nor U14532 (N_14532,N_9477,N_9232);
nand U14533 (N_14533,N_6130,N_5641);
nand U14534 (N_14534,N_8941,N_8567);
xor U14535 (N_14535,N_9360,N_8972);
and U14536 (N_14536,N_9784,N_8222);
nand U14537 (N_14537,N_8732,N_7656);
xnor U14538 (N_14538,N_5010,N_6717);
or U14539 (N_14539,N_8134,N_7577);
and U14540 (N_14540,N_8670,N_9070);
xor U14541 (N_14541,N_8811,N_7793);
nand U14542 (N_14542,N_5422,N_9647);
nand U14543 (N_14543,N_5395,N_6947);
or U14544 (N_14544,N_8176,N_5417);
xor U14545 (N_14545,N_6343,N_8994);
and U14546 (N_14546,N_5022,N_5909);
nand U14547 (N_14547,N_7684,N_5886);
nand U14548 (N_14548,N_7774,N_8860);
xnor U14549 (N_14549,N_6767,N_7113);
and U14550 (N_14550,N_5320,N_7087);
and U14551 (N_14551,N_8333,N_6327);
and U14552 (N_14552,N_7714,N_9890);
or U14553 (N_14553,N_9786,N_9576);
xnor U14554 (N_14554,N_6597,N_5678);
nor U14555 (N_14555,N_5395,N_6842);
and U14556 (N_14556,N_6332,N_6668);
xor U14557 (N_14557,N_8150,N_5131);
xnor U14558 (N_14558,N_5698,N_6472);
nand U14559 (N_14559,N_5769,N_7940);
and U14560 (N_14560,N_8501,N_9911);
and U14561 (N_14561,N_6157,N_5575);
and U14562 (N_14562,N_9241,N_5782);
xor U14563 (N_14563,N_8008,N_9714);
xnor U14564 (N_14564,N_7411,N_6762);
xnor U14565 (N_14565,N_6329,N_8796);
xnor U14566 (N_14566,N_7732,N_6673);
or U14567 (N_14567,N_7042,N_5975);
or U14568 (N_14568,N_6542,N_5224);
nand U14569 (N_14569,N_7471,N_9835);
xor U14570 (N_14570,N_5167,N_7035);
nand U14571 (N_14571,N_7737,N_5768);
nor U14572 (N_14572,N_9908,N_5340);
nor U14573 (N_14573,N_5065,N_9496);
or U14574 (N_14574,N_9022,N_6352);
or U14575 (N_14575,N_8116,N_5615);
or U14576 (N_14576,N_8955,N_7602);
or U14577 (N_14577,N_6517,N_6134);
or U14578 (N_14578,N_7043,N_7067);
xor U14579 (N_14579,N_9989,N_8938);
and U14580 (N_14580,N_5369,N_6942);
xor U14581 (N_14581,N_8625,N_7712);
nor U14582 (N_14582,N_7107,N_9946);
xnor U14583 (N_14583,N_5320,N_5801);
xnor U14584 (N_14584,N_7657,N_9194);
or U14585 (N_14585,N_5688,N_8728);
nand U14586 (N_14586,N_5113,N_5638);
xor U14587 (N_14587,N_5851,N_6157);
nor U14588 (N_14588,N_6635,N_9049);
or U14589 (N_14589,N_5819,N_6720);
nor U14590 (N_14590,N_9622,N_7029);
nand U14591 (N_14591,N_9761,N_8597);
or U14592 (N_14592,N_5376,N_6648);
or U14593 (N_14593,N_8162,N_7080);
nor U14594 (N_14594,N_6492,N_9910);
and U14595 (N_14595,N_9231,N_5970);
nor U14596 (N_14596,N_5277,N_5468);
and U14597 (N_14597,N_5059,N_5208);
and U14598 (N_14598,N_8617,N_5874);
and U14599 (N_14599,N_7253,N_5434);
nor U14600 (N_14600,N_8634,N_8301);
and U14601 (N_14601,N_7719,N_9807);
nand U14602 (N_14602,N_7103,N_5248);
or U14603 (N_14603,N_6493,N_8384);
and U14604 (N_14604,N_5486,N_9346);
and U14605 (N_14605,N_6698,N_5234);
nor U14606 (N_14606,N_8700,N_7162);
xor U14607 (N_14607,N_9059,N_7495);
nor U14608 (N_14608,N_8598,N_6919);
nor U14609 (N_14609,N_6347,N_5641);
xnor U14610 (N_14610,N_9248,N_9200);
nor U14611 (N_14611,N_9444,N_8103);
nand U14612 (N_14612,N_5801,N_9030);
nand U14613 (N_14613,N_8269,N_8840);
nand U14614 (N_14614,N_8665,N_8515);
nand U14615 (N_14615,N_9540,N_5032);
nor U14616 (N_14616,N_8150,N_5310);
or U14617 (N_14617,N_5030,N_7258);
nor U14618 (N_14618,N_7599,N_6115);
or U14619 (N_14619,N_5786,N_5267);
and U14620 (N_14620,N_5883,N_5685);
nor U14621 (N_14621,N_9472,N_5748);
nand U14622 (N_14622,N_7851,N_7015);
and U14623 (N_14623,N_9538,N_7732);
nand U14624 (N_14624,N_6023,N_8381);
xor U14625 (N_14625,N_6743,N_6336);
or U14626 (N_14626,N_8437,N_9832);
and U14627 (N_14627,N_8308,N_9971);
xor U14628 (N_14628,N_8078,N_5219);
nor U14629 (N_14629,N_6617,N_7498);
and U14630 (N_14630,N_8202,N_5441);
nand U14631 (N_14631,N_6676,N_8265);
nand U14632 (N_14632,N_7765,N_5732);
or U14633 (N_14633,N_5896,N_5621);
nand U14634 (N_14634,N_5819,N_7600);
and U14635 (N_14635,N_8375,N_5476);
nand U14636 (N_14636,N_7986,N_6407);
xor U14637 (N_14637,N_6308,N_7539);
nor U14638 (N_14638,N_7948,N_6437);
nor U14639 (N_14639,N_5719,N_8055);
xor U14640 (N_14640,N_9755,N_8982);
xor U14641 (N_14641,N_8582,N_5158);
xnor U14642 (N_14642,N_7109,N_5460);
nand U14643 (N_14643,N_6749,N_5527);
nor U14644 (N_14644,N_7247,N_7126);
or U14645 (N_14645,N_5964,N_9608);
and U14646 (N_14646,N_5511,N_5040);
xnor U14647 (N_14647,N_5072,N_8751);
xnor U14648 (N_14648,N_8495,N_7847);
and U14649 (N_14649,N_6192,N_9825);
and U14650 (N_14650,N_7943,N_7089);
nand U14651 (N_14651,N_7373,N_5666);
nand U14652 (N_14652,N_9341,N_5565);
or U14653 (N_14653,N_6538,N_5250);
xnor U14654 (N_14654,N_6442,N_5369);
xor U14655 (N_14655,N_8535,N_6887);
nand U14656 (N_14656,N_6185,N_7550);
or U14657 (N_14657,N_9064,N_8307);
nor U14658 (N_14658,N_6969,N_6215);
and U14659 (N_14659,N_9174,N_9722);
xor U14660 (N_14660,N_7702,N_7443);
or U14661 (N_14661,N_9994,N_7437);
and U14662 (N_14662,N_9083,N_7107);
and U14663 (N_14663,N_8676,N_9518);
xor U14664 (N_14664,N_8071,N_8182);
or U14665 (N_14665,N_5324,N_8579);
or U14666 (N_14666,N_8449,N_7484);
nor U14667 (N_14667,N_5517,N_9690);
xnor U14668 (N_14668,N_8588,N_6706);
and U14669 (N_14669,N_5861,N_6463);
or U14670 (N_14670,N_6592,N_8369);
xor U14671 (N_14671,N_7313,N_9244);
xor U14672 (N_14672,N_9647,N_7011);
nor U14673 (N_14673,N_8961,N_6732);
or U14674 (N_14674,N_8498,N_9631);
xor U14675 (N_14675,N_8465,N_9628);
nor U14676 (N_14676,N_7696,N_6846);
and U14677 (N_14677,N_6585,N_9461);
nor U14678 (N_14678,N_8978,N_6983);
nor U14679 (N_14679,N_5827,N_7888);
and U14680 (N_14680,N_5941,N_8695);
xnor U14681 (N_14681,N_9437,N_9284);
nor U14682 (N_14682,N_5293,N_5647);
nand U14683 (N_14683,N_7826,N_5992);
nand U14684 (N_14684,N_6935,N_8914);
nor U14685 (N_14685,N_6537,N_6061);
nand U14686 (N_14686,N_7523,N_5836);
nor U14687 (N_14687,N_9674,N_6969);
and U14688 (N_14688,N_8638,N_5450);
xor U14689 (N_14689,N_7533,N_8459);
nand U14690 (N_14690,N_6972,N_6816);
xor U14691 (N_14691,N_8438,N_8709);
xnor U14692 (N_14692,N_9282,N_7186);
and U14693 (N_14693,N_8764,N_9817);
nand U14694 (N_14694,N_7918,N_9653);
or U14695 (N_14695,N_8185,N_7678);
or U14696 (N_14696,N_6857,N_6690);
xnor U14697 (N_14697,N_9885,N_6920);
and U14698 (N_14698,N_8117,N_9328);
nand U14699 (N_14699,N_5506,N_5645);
nor U14700 (N_14700,N_8495,N_5111);
nor U14701 (N_14701,N_9535,N_5573);
and U14702 (N_14702,N_6120,N_6569);
nand U14703 (N_14703,N_5605,N_6803);
nand U14704 (N_14704,N_5164,N_6496);
or U14705 (N_14705,N_7654,N_5023);
or U14706 (N_14706,N_6041,N_5755);
nor U14707 (N_14707,N_7824,N_5625);
and U14708 (N_14708,N_9833,N_9012);
and U14709 (N_14709,N_9437,N_5943);
nand U14710 (N_14710,N_5591,N_9144);
nand U14711 (N_14711,N_6383,N_6088);
and U14712 (N_14712,N_6405,N_6574);
xnor U14713 (N_14713,N_7702,N_8435);
or U14714 (N_14714,N_7273,N_6183);
nor U14715 (N_14715,N_5212,N_6877);
and U14716 (N_14716,N_8207,N_8906);
nor U14717 (N_14717,N_7713,N_6938);
xor U14718 (N_14718,N_8121,N_5984);
nand U14719 (N_14719,N_7539,N_7496);
nand U14720 (N_14720,N_8351,N_9216);
and U14721 (N_14721,N_7671,N_6437);
nor U14722 (N_14722,N_6830,N_5110);
nand U14723 (N_14723,N_5194,N_9267);
nor U14724 (N_14724,N_6070,N_9922);
and U14725 (N_14725,N_5581,N_9470);
nor U14726 (N_14726,N_7057,N_7452);
xor U14727 (N_14727,N_9286,N_9862);
nor U14728 (N_14728,N_7440,N_9942);
nor U14729 (N_14729,N_7125,N_8975);
nor U14730 (N_14730,N_6444,N_7852);
nor U14731 (N_14731,N_8304,N_7170);
nand U14732 (N_14732,N_8657,N_9505);
or U14733 (N_14733,N_9611,N_9510);
xnor U14734 (N_14734,N_7679,N_5737);
xor U14735 (N_14735,N_6811,N_6864);
and U14736 (N_14736,N_9565,N_8141);
nor U14737 (N_14737,N_9730,N_6475);
or U14738 (N_14738,N_8128,N_9398);
xor U14739 (N_14739,N_9362,N_9587);
nand U14740 (N_14740,N_7595,N_9365);
or U14741 (N_14741,N_5660,N_9567);
and U14742 (N_14742,N_6701,N_5408);
nor U14743 (N_14743,N_7628,N_8604);
xor U14744 (N_14744,N_6857,N_6950);
nand U14745 (N_14745,N_5660,N_8980);
nand U14746 (N_14746,N_5156,N_6716);
nor U14747 (N_14747,N_6112,N_9527);
nand U14748 (N_14748,N_9332,N_5818);
nor U14749 (N_14749,N_7002,N_6370);
nand U14750 (N_14750,N_6444,N_5638);
nor U14751 (N_14751,N_9077,N_7152);
xnor U14752 (N_14752,N_5196,N_6766);
or U14753 (N_14753,N_7323,N_9982);
xor U14754 (N_14754,N_7835,N_6629);
and U14755 (N_14755,N_7303,N_5155);
and U14756 (N_14756,N_6007,N_9973);
nor U14757 (N_14757,N_9812,N_8032);
and U14758 (N_14758,N_8599,N_5781);
or U14759 (N_14759,N_8483,N_8666);
nand U14760 (N_14760,N_6155,N_6107);
xnor U14761 (N_14761,N_8434,N_6909);
nor U14762 (N_14762,N_6775,N_5728);
nor U14763 (N_14763,N_7013,N_6508);
nand U14764 (N_14764,N_5307,N_7282);
nand U14765 (N_14765,N_6900,N_6584);
xnor U14766 (N_14766,N_9941,N_8151);
or U14767 (N_14767,N_9881,N_6254);
or U14768 (N_14768,N_7324,N_5360);
nor U14769 (N_14769,N_6350,N_7910);
and U14770 (N_14770,N_6506,N_9667);
and U14771 (N_14771,N_8527,N_5102);
and U14772 (N_14772,N_8694,N_5236);
or U14773 (N_14773,N_8461,N_6198);
and U14774 (N_14774,N_9653,N_7268);
or U14775 (N_14775,N_7460,N_9247);
or U14776 (N_14776,N_6975,N_8847);
nand U14777 (N_14777,N_5465,N_8117);
nand U14778 (N_14778,N_8505,N_7196);
nand U14779 (N_14779,N_8308,N_6544);
and U14780 (N_14780,N_5257,N_7738);
and U14781 (N_14781,N_9366,N_9330);
xor U14782 (N_14782,N_6816,N_5898);
nor U14783 (N_14783,N_9028,N_5627);
or U14784 (N_14784,N_7717,N_8531);
nand U14785 (N_14785,N_6525,N_6379);
or U14786 (N_14786,N_8390,N_9313);
xor U14787 (N_14787,N_9009,N_5105);
and U14788 (N_14788,N_5632,N_7275);
or U14789 (N_14789,N_8365,N_9019);
and U14790 (N_14790,N_9461,N_5941);
xnor U14791 (N_14791,N_5912,N_6544);
and U14792 (N_14792,N_9336,N_9401);
nand U14793 (N_14793,N_9288,N_9533);
nor U14794 (N_14794,N_7358,N_9886);
xor U14795 (N_14795,N_6449,N_5430);
and U14796 (N_14796,N_9537,N_7202);
nand U14797 (N_14797,N_6145,N_7551);
and U14798 (N_14798,N_9460,N_5845);
nand U14799 (N_14799,N_5225,N_8199);
nor U14800 (N_14800,N_6197,N_7952);
and U14801 (N_14801,N_9911,N_6484);
nor U14802 (N_14802,N_7909,N_5152);
and U14803 (N_14803,N_8783,N_6426);
nor U14804 (N_14804,N_8461,N_7905);
or U14805 (N_14805,N_8510,N_7723);
or U14806 (N_14806,N_8719,N_9441);
xor U14807 (N_14807,N_9565,N_9895);
xor U14808 (N_14808,N_8175,N_7593);
and U14809 (N_14809,N_6757,N_6277);
nor U14810 (N_14810,N_8583,N_8025);
xnor U14811 (N_14811,N_5462,N_6910);
nand U14812 (N_14812,N_8237,N_8189);
or U14813 (N_14813,N_5681,N_9483);
xor U14814 (N_14814,N_9651,N_7698);
xor U14815 (N_14815,N_6443,N_9696);
xor U14816 (N_14816,N_6546,N_9228);
and U14817 (N_14817,N_6474,N_6603);
nor U14818 (N_14818,N_9662,N_6675);
xnor U14819 (N_14819,N_8615,N_8028);
or U14820 (N_14820,N_5256,N_7985);
and U14821 (N_14821,N_7748,N_7291);
and U14822 (N_14822,N_6626,N_5688);
xor U14823 (N_14823,N_9604,N_6322);
nand U14824 (N_14824,N_7081,N_5009);
and U14825 (N_14825,N_9688,N_7805);
or U14826 (N_14826,N_8632,N_5072);
nor U14827 (N_14827,N_9518,N_8088);
or U14828 (N_14828,N_7059,N_7358);
and U14829 (N_14829,N_8332,N_6171);
nand U14830 (N_14830,N_7772,N_9495);
or U14831 (N_14831,N_7126,N_6714);
xor U14832 (N_14832,N_7632,N_5998);
and U14833 (N_14833,N_6546,N_8130);
nand U14834 (N_14834,N_7466,N_9740);
nand U14835 (N_14835,N_8363,N_7083);
xnor U14836 (N_14836,N_6872,N_6375);
nor U14837 (N_14837,N_8129,N_6615);
or U14838 (N_14838,N_5902,N_8359);
xor U14839 (N_14839,N_7975,N_5388);
and U14840 (N_14840,N_9640,N_5643);
nand U14841 (N_14841,N_7761,N_7524);
or U14842 (N_14842,N_6166,N_6170);
or U14843 (N_14843,N_8407,N_8997);
nand U14844 (N_14844,N_8892,N_9113);
xnor U14845 (N_14845,N_5283,N_6455);
nand U14846 (N_14846,N_5356,N_6665);
xor U14847 (N_14847,N_5403,N_5392);
nand U14848 (N_14848,N_8778,N_5379);
nor U14849 (N_14849,N_8222,N_8394);
xnor U14850 (N_14850,N_6297,N_6694);
nor U14851 (N_14851,N_7737,N_9113);
nor U14852 (N_14852,N_5280,N_6870);
nor U14853 (N_14853,N_6444,N_6555);
and U14854 (N_14854,N_7981,N_7609);
or U14855 (N_14855,N_8775,N_8184);
and U14856 (N_14856,N_5223,N_5727);
and U14857 (N_14857,N_7011,N_8347);
or U14858 (N_14858,N_7368,N_7947);
nor U14859 (N_14859,N_5208,N_9675);
and U14860 (N_14860,N_8705,N_6267);
nor U14861 (N_14861,N_5886,N_6951);
nor U14862 (N_14862,N_5625,N_9597);
xnor U14863 (N_14863,N_7561,N_7197);
and U14864 (N_14864,N_7695,N_5383);
nand U14865 (N_14865,N_6738,N_8967);
nor U14866 (N_14866,N_9513,N_5080);
xor U14867 (N_14867,N_5104,N_8774);
and U14868 (N_14868,N_6856,N_7930);
nand U14869 (N_14869,N_8194,N_7731);
nor U14870 (N_14870,N_5701,N_5242);
xor U14871 (N_14871,N_6140,N_9730);
nand U14872 (N_14872,N_8436,N_8705);
and U14873 (N_14873,N_5206,N_5397);
and U14874 (N_14874,N_5697,N_6488);
and U14875 (N_14875,N_9382,N_7423);
xor U14876 (N_14876,N_7404,N_6905);
and U14877 (N_14877,N_8191,N_6902);
xnor U14878 (N_14878,N_7025,N_8113);
nand U14879 (N_14879,N_9138,N_7124);
nand U14880 (N_14880,N_9723,N_8332);
nand U14881 (N_14881,N_5841,N_8382);
or U14882 (N_14882,N_9465,N_5110);
and U14883 (N_14883,N_8129,N_6824);
and U14884 (N_14884,N_9502,N_7587);
xnor U14885 (N_14885,N_7670,N_6470);
xor U14886 (N_14886,N_5864,N_6825);
nor U14887 (N_14887,N_6122,N_7759);
nand U14888 (N_14888,N_9340,N_7345);
xnor U14889 (N_14889,N_6293,N_8706);
nor U14890 (N_14890,N_6463,N_7809);
nand U14891 (N_14891,N_5168,N_8057);
nor U14892 (N_14892,N_9177,N_7824);
nand U14893 (N_14893,N_5656,N_9240);
nand U14894 (N_14894,N_5654,N_6153);
nand U14895 (N_14895,N_5677,N_8158);
and U14896 (N_14896,N_6951,N_8880);
or U14897 (N_14897,N_7591,N_7671);
and U14898 (N_14898,N_8053,N_5457);
nor U14899 (N_14899,N_8932,N_8804);
or U14900 (N_14900,N_5730,N_7812);
xnor U14901 (N_14901,N_8901,N_6889);
nand U14902 (N_14902,N_8612,N_7192);
nand U14903 (N_14903,N_8889,N_5137);
and U14904 (N_14904,N_5648,N_7088);
nor U14905 (N_14905,N_7395,N_8268);
or U14906 (N_14906,N_9237,N_8648);
nand U14907 (N_14907,N_9634,N_9226);
and U14908 (N_14908,N_7961,N_8407);
and U14909 (N_14909,N_7726,N_9898);
nand U14910 (N_14910,N_7737,N_8659);
nor U14911 (N_14911,N_9996,N_6912);
or U14912 (N_14912,N_5676,N_6115);
and U14913 (N_14913,N_5100,N_5967);
xnor U14914 (N_14914,N_8958,N_6880);
or U14915 (N_14915,N_5043,N_7198);
nand U14916 (N_14916,N_9494,N_7895);
and U14917 (N_14917,N_7987,N_5954);
nor U14918 (N_14918,N_8481,N_7969);
nand U14919 (N_14919,N_5645,N_5497);
nand U14920 (N_14920,N_6848,N_6680);
and U14921 (N_14921,N_7288,N_9418);
nor U14922 (N_14922,N_7455,N_8001);
or U14923 (N_14923,N_5759,N_9131);
and U14924 (N_14924,N_7631,N_8766);
nand U14925 (N_14925,N_9360,N_9307);
and U14926 (N_14926,N_9961,N_6770);
nand U14927 (N_14927,N_9567,N_6353);
nor U14928 (N_14928,N_5048,N_6876);
nand U14929 (N_14929,N_8829,N_6746);
and U14930 (N_14930,N_6348,N_8282);
nor U14931 (N_14931,N_8730,N_5784);
nor U14932 (N_14932,N_7218,N_7070);
or U14933 (N_14933,N_8510,N_9092);
nor U14934 (N_14934,N_8533,N_8667);
or U14935 (N_14935,N_6863,N_9484);
nand U14936 (N_14936,N_6566,N_7485);
nor U14937 (N_14937,N_7397,N_5719);
and U14938 (N_14938,N_7202,N_5436);
xnor U14939 (N_14939,N_9262,N_7233);
or U14940 (N_14940,N_8952,N_8893);
nor U14941 (N_14941,N_7288,N_8737);
xnor U14942 (N_14942,N_8618,N_5588);
and U14943 (N_14943,N_6768,N_8577);
nand U14944 (N_14944,N_5978,N_5593);
and U14945 (N_14945,N_5376,N_9944);
nand U14946 (N_14946,N_7448,N_8772);
nor U14947 (N_14947,N_6563,N_8590);
and U14948 (N_14948,N_9196,N_6704);
nor U14949 (N_14949,N_7136,N_7941);
nor U14950 (N_14950,N_5716,N_8804);
or U14951 (N_14951,N_6754,N_7951);
nand U14952 (N_14952,N_8054,N_9086);
or U14953 (N_14953,N_7874,N_8748);
xnor U14954 (N_14954,N_7701,N_7574);
and U14955 (N_14955,N_8308,N_7159);
nor U14956 (N_14956,N_6177,N_6991);
and U14957 (N_14957,N_5139,N_5984);
and U14958 (N_14958,N_7736,N_6271);
xor U14959 (N_14959,N_9147,N_6284);
nand U14960 (N_14960,N_5662,N_9995);
nand U14961 (N_14961,N_5681,N_5103);
or U14962 (N_14962,N_8536,N_6517);
xor U14963 (N_14963,N_7179,N_9709);
nor U14964 (N_14964,N_6006,N_7267);
or U14965 (N_14965,N_9585,N_7964);
or U14966 (N_14966,N_5992,N_5431);
nand U14967 (N_14967,N_7760,N_8114);
or U14968 (N_14968,N_6624,N_6031);
and U14969 (N_14969,N_9302,N_8221);
nand U14970 (N_14970,N_8568,N_7640);
and U14971 (N_14971,N_6794,N_9702);
nand U14972 (N_14972,N_8306,N_5835);
or U14973 (N_14973,N_9422,N_7059);
nor U14974 (N_14974,N_5849,N_6006);
or U14975 (N_14975,N_7247,N_7748);
nand U14976 (N_14976,N_6687,N_5655);
nand U14977 (N_14977,N_5951,N_6583);
and U14978 (N_14978,N_9526,N_6236);
nor U14979 (N_14979,N_8949,N_5989);
nand U14980 (N_14980,N_5112,N_7954);
xor U14981 (N_14981,N_6379,N_9610);
nand U14982 (N_14982,N_9496,N_6338);
xnor U14983 (N_14983,N_7558,N_6875);
nand U14984 (N_14984,N_8262,N_5837);
and U14985 (N_14985,N_8620,N_6305);
xor U14986 (N_14986,N_6683,N_9181);
nand U14987 (N_14987,N_9321,N_5838);
nand U14988 (N_14988,N_5619,N_5158);
nand U14989 (N_14989,N_7926,N_8688);
nor U14990 (N_14990,N_9395,N_7846);
xor U14991 (N_14991,N_7740,N_7035);
and U14992 (N_14992,N_7281,N_8603);
and U14993 (N_14993,N_7152,N_9558);
or U14994 (N_14994,N_5919,N_7568);
xor U14995 (N_14995,N_5326,N_5486);
xor U14996 (N_14996,N_8077,N_9401);
or U14997 (N_14997,N_8705,N_9374);
or U14998 (N_14998,N_9608,N_9067);
and U14999 (N_14999,N_6345,N_8372);
nor U15000 (N_15000,N_14288,N_14779);
and U15001 (N_15001,N_14153,N_13652);
nand U15002 (N_15002,N_14422,N_12487);
nand U15003 (N_15003,N_11739,N_12417);
and U15004 (N_15004,N_11875,N_13856);
nor U15005 (N_15005,N_12680,N_10284);
xnor U15006 (N_15006,N_14594,N_13694);
nor U15007 (N_15007,N_10935,N_11375);
or U15008 (N_15008,N_11422,N_10910);
nand U15009 (N_15009,N_13621,N_14949);
xor U15010 (N_15010,N_10791,N_14404);
or U15011 (N_15011,N_13761,N_14495);
xor U15012 (N_15012,N_13219,N_13014);
or U15013 (N_15013,N_14449,N_13439);
nand U15014 (N_15014,N_14147,N_13682);
xor U15015 (N_15015,N_12084,N_12443);
xor U15016 (N_15016,N_11018,N_14239);
and U15017 (N_15017,N_11929,N_12385);
xor U15018 (N_15018,N_10270,N_12466);
nor U15019 (N_15019,N_12383,N_11295);
nand U15020 (N_15020,N_14666,N_11961);
nor U15021 (N_15021,N_10786,N_11881);
nor U15022 (N_15022,N_12067,N_10522);
or U15023 (N_15023,N_11222,N_12689);
nand U15024 (N_15024,N_11265,N_11564);
nand U15025 (N_15025,N_12713,N_14442);
and U15026 (N_15026,N_13547,N_13985);
xor U15027 (N_15027,N_12145,N_14084);
nor U15028 (N_15028,N_12502,N_13039);
xnor U15029 (N_15029,N_10075,N_10185);
xnor U15030 (N_15030,N_13596,N_11818);
nor U15031 (N_15031,N_11619,N_10829);
xor U15032 (N_15032,N_10821,N_12769);
nor U15033 (N_15033,N_14311,N_13524);
or U15034 (N_15034,N_10517,N_12564);
xor U15035 (N_15035,N_14165,N_14653);
or U15036 (N_15036,N_13667,N_12904);
xnor U15037 (N_15037,N_10255,N_10119);
and U15038 (N_15038,N_12891,N_14646);
or U15039 (N_15039,N_10155,N_10648);
and U15040 (N_15040,N_13375,N_12106);
nor U15041 (N_15041,N_11182,N_11104);
nor U15042 (N_15042,N_13809,N_13755);
and U15043 (N_15043,N_11839,N_10302);
nand U15044 (N_15044,N_14962,N_13297);
nand U15045 (N_15045,N_13277,N_14960);
and U15046 (N_15046,N_13745,N_12806);
nor U15047 (N_15047,N_10693,N_11670);
nor U15048 (N_15048,N_14007,N_13204);
and U15049 (N_15049,N_10236,N_13157);
xor U15050 (N_15050,N_10414,N_10843);
nand U15051 (N_15051,N_13127,N_10232);
and U15052 (N_15052,N_14378,N_12820);
xnor U15053 (N_15053,N_13525,N_12754);
nand U15054 (N_15054,N_13043,N_13666);
and U15055 (N_15055,N_10896,N_10246);
nor U15056 (N_15056,N_13687,N_10895);
or U15057 (N_15057,N_12584,N_12469);
xor U15058 (N_15058,N_12866,N_11299);
nand U15059 (N_15059,N_11856,N_14738);
nand U15060 (N_15060,N_14811,N_10130);
nand U15061 (N_15061,N_10555,N_11046);
and U15062 (N_15062,N_10763,N_13681);
xnor U15063 (N_15063,N_14881,N_13403);
nand U15064 (N_15064,N_14105,N_10881);
xnor U15065 (N_15065,N_14580,N_13427);
nor U15066 (N_15066,N_13728,N_10090);
and U15067 (N_15067,N_11365,N_11951);
nand U15068 (N_15068,N_13925,N_12041);
nand U15069 (N_15069,N_10165,N_11121);
nand U15070 (N_15070,N_11216,N_10887);
nand U15071 (N_15071,N_12932,N_10636);
xnor U15072 (N_15072,N_14461,N_10727);
or U15073 (N_15073,N_10040,N_13217);
nand U15074 (N_15074,N_12222,N_13190);
nand U15075 (N_15075,N_10142,N_10877);
or U15076 (N_15076,N_10469,N_11040);
or U15077 (N_15077,N_14794,N_12353);
and U15078 (N_15078,N_12302,N_10134);
and U15079 (N_15079,N_14188,N_12297);
nor U15080 (N_15080,N_11709,N_13213);
or U15081 (N_15081,N_12532,N_13141);
nor U15082 (N_15082,N_11024,N_11534);
nor U15083 (N_15083,N_13743,N_11538);
nand U15084 (N_15084,N_13600,N_10824);
and U15085 (N_15085,N_12474,N_14205);
and U15086 (N_15086,N_10511,N_13058);
and U15087 (N_15087,N_11447,N_12011);
and U15088 (N_15088,N_14087,N_13706);
and U15089 (N_15089,N_14723,N_11908);
and U15090 (N_15090,N_11398,N_13889);
nand U15091 (N_15091,N_10726,N_11656);
or U15092 (N_15092,N_11631,N_10026);
and U15093 (N_15093,N_13988,N_12803);
nand U15094 (N_15094,N_14874,N_13451);
or U15095 (N_15095,N_12373,N_12351);
xor U15096 (N_15096,N_11136,N_13149);
or U15097 (N_15097,N_14674,N_11033);
or U15098 (N_15098,N_12146,N_10961);
nand U15099 (N_15099,N_13590,N_12986);
nor U15100 (N_15100,N_13983,N_11647);
xnor U15101 (N_15101,N_14108,N_14432);
or U15102 (N_15102,N_14783,N_11554);
or U15103 (N_15103,N_10673,N_13092);
xnor U15104 (N_15104,N_13421,N_10928);
nor U15105 (N_15105,N_11490,N_12020);
and U15106 (N_15106,N_10239,N_14967);
nand U15107 (N_15107,N_12332,N_13876);
xor U15108 (N_15108,N_10374,N_10157);
nor U15109 (N_15109,N_11622,N_14233);
xnor U15110 (N_15110,N_14175,N_10003);
nor U15111 (N_15111,N_11420,N_11871);
nor U15112 (N_15112,N_14324,N_10675);
or U15113 (N_15113,N_12241,N_10558);
nor U15114 (N_15114,N_13036,N_12509);
or U15115 (N_15115,N_10898,N_13046);
nand U15116 (N_15116,N_14510,N_12597);
and U15117 (N_15117,N_13475,N_14560);
nand U15118 (N_15118,N_11518,N_14648);
nor U15119 (N_15119,N_10947,N_10783);
nand U15120 (N_15120,N_12163,N_12093);
xor U15121 (N_15121,N_14937,N_12256);
nor U15122 (N_15122,N_14182,N_13601);
and U15123 (N_15123,N_11456,N_10341);
or U15124 (N_15124,N_14530,N_12666);
nor U15125 (N_15125,N_12733,N_12056);
or U15126 (N_15126,N_11442,N_14193);
nor U15127 (N_15127,N_14715,N_11237);
xor U15128 (N_15128,N_10657,N_14073);
and U15129 (N_15129,N_11700,N_14720);
nor U15130 (N_15130,N_10574,N_10833);
and U15131 (N_15131,N_12157,N_12402);
or U15132 (N_15132,N_14423,N_14200);
nand U15133 (N_15133,N_11096,N_11746);
nand U15134 (N_15134,N_13541,N_13737);
nor U15135 (N_15135,N_10136,N_13026);
or U15136 (N_15136,N_12877,N_13722);
and U15137 (N_15137,N_14312,N_12944);
or U15138 (N_15138,N_11239,N_10544);
or U15139 (N_15139,N_13201,N_10366);
or U15140 (N_15140,N_11982,N_12085);
and U15141 (N_15141,N_10735,N_13919);
and U15142 (N_15142,N_12730,N_12954);
or U15143 (N_15143,N_11783,N_13469);
or U15144 (N_15144,N_14808,N_12508);
nand U15145 (N_15145,N_10269,N_12996);
xor U15146 (N_15146,N_10942,N_11142);
and U15147 (N_15147,N_10547,N_14883);
and U15148 (N_15148,N_11051,N_13772);
and U15149 (N_15149,N_12639,N_11188);
xnor U15150 (N_15150,N_10262,N_12786);
xor U15151 (N_15151,N_11423,N_10656);
xor U15152 (N_15152,N_13620,N_14622);
and U15153 (N_15153,N_13478,N_12071);
and U15154 (N_15154,N_13507,N_11460);
nor U15155 (N_15155,N_11273,N_14730);
or U15156 (N_15156,N_11342,N_10370);
or U15157 (N_15157,N_13680,N_12560);
nand U15158 (N_15158,N_13565,N_13150);
xnor U15159 (N_15159,N_13397,N_12358);
and U15160 (N_15160,N_12831,N_10927);
xnor U15161 (N_15161,N_10061,N_12805);
nor U15162 (N_15162,N_12287,N_14067);
nand U15163 (N_15163,N_10875,N_13206);
nor U15164 (N_15164,N_13227,N_12075);
and U15165 (N_15165,N_10129,N_12655);
nor U15166 (N_15166,N_11771,N_13113);
xnor U15167 (N_15167,N_10295,N_12375);
and U15168 (N_15168,N_10551,N_11812);
and U15169 (N_15169,N_13212,N_13774);
and U15170 (N_15170,N_13707,N_14463);
or U15171 (N_15171,N_11168,N_12717);
xnor U15172 (N_15172,N_11075,N_10036);
nor U15173 (N_15173,N_11047,N_12648);
nor U15174 (N_15174,N_10664,N_11230);
xor U15175 (N_15175,N_14869,N_10987);
and U15176 (N_15176,N_13057,N_13195);
and U15177 (N_15177,N_13029,N_12591);
or U15178 (N_15178,N_10912,N_10752);
xor U15179 (N_15179,N_13518,N_11960);
or U15180 (N_15180,N_11787,N_10449);
nand U15181 (N_15181,N_12814,N_14004);
nor U15182 (N_15182,N_14889,N_13374);
or U15183 (N_15183,N_14186,N_14323);
nand U15184 (N_15184,N_13814,N_12840);
and U15185 (N_15185,N_10808,N_14839);
or U15186 (N_15186,N_13976,N_11226);
nor U15187 (N_15187,N_11515,N_14953);
nand U15188 (N_15188,N_10132,N_12314);
nor U15189 (N_15189,N_14337,N_14824);
nor U15190 (N_15190,N_11574,N_14524);
nand U15191 (N_15191,N_11772,N_12112);
or U15192 (N_15192,N_11860,N_11338);
nand U15193 (N_15193,N_10672,N_13368);
or U15194 (N_15194,N_14245,N_11020);
and U15195 (N_15195,N_13936,N_10353);
nand U15196 (N_15196,N_10765,N_14458);
nand U15197 (N_15197,N_13870,N_14921);
and U15198 (N_15198,N_10327,N_12282);
nor U15199 (N_15199,N_14887,N_13702);
nand U15200 (N_15200,N_14275,N_13658);
nor U15201 (N_15201,N_13691,N_13758);
xor U15202 (N_15202,N_12547,N_10600);
and U15203 (N_15203,N_13330,N_12123);
or U15204 (N_15204,N_14212,N_13114);
nor U15205 (N_15205,N_10968,N_13154);
xnor U15206 (N_15206,N_10851,N_10836);
or U15207 (N_15207,N_13426,N_13588);
nand U15208 (N_15208,N_12337,N_13926);
nand U15209 (N_15209,N_11270,N_12943);
and U15210 (N_15210,N_11737,N_13796);
and U15211 (N_15211,N_13538,N_14799);
xnor U15212 (N_15212,N_13096,N_12037);
or U15213 (N_15213,N_12214,N_14727);
nor U15214 (N_15214,N_10144,N_10103);
nand U15215 (N_15215,N_14521,N_13402);
nand U15216 (N_15216,N_13757,N_13326);
nor U15217 (N_15217,N_12187,N_11571);
nand U15218 (N_15218,N_12772,N_11603);
and U15219 (N_15219,N_13351,N_13136);
and U15220 (N_15220,N_10241,N_11478);
xor U15221 (N_15221,N_13054,N_11093);
xor U15222 (N_15222,N_10623,N_10041);
nand U15223 (N_15223,N_13725,N_11598);
nand U15224 (N_15224,N_11085,N_14904);
nor U15225 (N_15225,N_10461,N_12218);
nor U15226 (N_15226,N_11568,N_13903);
and U15227 (N_15227,N_11890,N_13515);
xor U15228 (N_15228,N_10478,N_13957);
xor U15229 (N_15229,N_10897,N_12078);
nor U15230 (N_15230,N_13465,N_13360);
nor U15231 (N_15231,N_13730,N_12662);
nor U15232 (N_15232,N_10939,N_10434);
xor U15233 (N_15233,N_13429,N_13486);
and U15234 (N_15234,N_11102,N_11319);
nor U15235 (N_15235,N_13408,N_13877);
xnor U15236 (N_15236,N_14013,N_14999);
and U15237 (N_15237,N_14704,N_14425);
and U15238 (N_15238,N_11120,N_14424);
xnor U15239 (N_15239,N_13276,N_13477);
or U15240 (N_15240,N_14788,N_14400);
nand U15241 (N_15241,N_14001,N_11496);
and U15242 (N_15242,N_10224,N_11708);
nand U15243 (N_15243,N_12773,N_10178);
and U15244 (N_15244,N_14229,N_14787);
xor U15245 (N_15245,N_11902,N_12008);
and U15246 (N_15246,N_13854,N_13570);
or U15247 (N_15247,N_13846,N_13754);
or U15248 (N_15248,N_10335,N_11057);
nand U15249 (N_15249,N_12625,N_14637);
nor U15250 (N_15250,N_10689,N_14396);
nor U15251 (N_15251,N_13389,N_11092);
or U15252 (N_15252,N_13193,N_14988);
or U15253 (N_15253,N_14778,N_14011);
or U15254 (N_15254,N_13237,N_10306);
xor U15255 (N_15255,N_14218,N_12215);
nand U15256 (N_15256,N_11770,N_10645);
nor U15257 (N_15257,N_14065,N_11565);
xnor U15258 (N_15258,N_10181,N_14315);
nand U15259 (N_15259,N_11830,N_13683);
and U15260 (N_15260,N_12335,N_14803);
nor U15261 (N_15261,N_13999,N_12993);
xnor U15262 (N_15262,N_14907,N_12143);
nor U15263 (N_15263,N_11048,N_14052);
or U15264 (N_15264,N_13211,N_14393);
nand U15265 (N_15265,N_11337,N_12470);
xor U15266 (N_15266,N_10274,N_12305);
nand U15267 (N_15267,N_12511,N_10499);
and U15268 (N_15268,N_11089,N_10030);
or U15269 (N_15269,N_14349,N_13557);
nor U15270 (N_15270,N_12857,N_12552);
nor U15271 (N_15271,N_14047,N_14252);
and U15272 (N_15272,N_13868,N_11235);
nor U15273 (N_15273,N_12245,N_12912);
or U15274 (N_15274,N_13939,N_10846);
or U15275 (N_15275,N_10100,N_11964);
nor U15276 (N_15276,N_12559,N_10742);
xor U15277 (N_15277,N_14303,N_14161);
or U15278 (N_15278,N_13184,N_11062);
xnor U15279 (N_15279,N_13280,N_12293);
nand U15280 (N_15280,N_10076,N_11191);
or U15281 (N_15281,N_10131,N_14050);
nand U15282 (N_15282,N_12367,N_10339);
and U15283 (N_15283,N_12267,N_10467);
nor U15284 (N_15284,N_11981,N_13175);
nor U15285 (N_15285,N_13715,N_10305);
nor U15286 (N_15286,N_13642,N_13239);
and U15287 (N_15287,N_10744,N_14553);
and U15288 (N_15288,N_12685,N_13312);
or U15289 (N_15289,N_14922,N_13637);
and U15290 (N_15290,N_11035,N_10571);
and U15291 (N_15291,N_11392,N_12251);
nand U15292 (N_15292,N_13632,N_14978);
or U15293 (N_15293,N_11817,N_11227);
and U15294 (N_15294,N_14729,N_11976);
or U15295 (N_15295,N_11627,N_13696);
nor U15296 (N_15296,N_11006,N_12053);
and U15297 (N_15297,N_14115,N_11274);
xor U15298 (N_15298,N_12536,N_13606);
or U15299 (N_15299,N_10694,N_13143);
or U15300 (N_15300,N_11792,N_13468);
and U15301 (N_15301,N_14601,N_11466);
nand U15302 (N_15302,N_10981,N_10159);
nor U15303 (N_15303,N_12600,N_12488);
xnor U15304 (N_15304,N_14016,N_14399);
xnor U15305 (N_15305,N_10330,N_14125);
and U15306 (N_15306,N_14636,N_11693);
nor U15307 (N_15307,N_12530,N_11347);
nand U15308 (N_15308,N_12343,N_11570);
nor U15309 (N_15309,N_12423,N_11986);
or U15310 (N_15310,N_10161,N_12453);
and U15311 (N_15311,N_12098,N_10698);
nand U15312 (N_15312,N_14494,N_13893);
or U15313 (N_15313,N_10776,N_12158);
xnor U15314 (N_15314,N_12963,N_10139);
nand U15315 (N_15315,N_13888,N_11012);
nor U15316 (N_15316,N_14136,N_13921);
xnor U15317 (N_15317,N_14990,N_11155);
and U15318 (N_15318,N_14375,N_14157);
nand U15319 (N_15319,N_13793,N_14818);
and U15320 (N_15320,N_10539,N_13852);
xnor U15321 (N_15321,N_13367,N_14330);
nand U15322 (N_15322,N_12496,N_10622);
nor U15323 (N_15323,N_11997,N_10900);
xnor U15324 (N_15324,N_14512,N_14629);
xor U15325 (N_15325,N_10501,N_10853);
or U15326 (N_15326,N_12190,N_11323);
nand U15327 (N_15327,N_10008,N_13441);
xor U15328 (N_15328,N_11941,N_12882);
and U15329 (N_15329,N_13676,N_10818);
nand U15330 (N_15330,N_11143,N_10415);
xor U15331 (N_15331,N_10117,N_11256);
nand U15332 (N_15332,N_12802,N_11873);
nor U15333 (N_15333,N_14167,N_12339);
and U15334 (N_15334,N_10087,N_10253);
nor U15335 (N_15335,N_13309,N_10223);
and U15336 (N_15336,N_11264,N_11491);
and U15337 (N_15337,N_13533,N_11269);
nand U15338 (N_15338,N_12283,N_10834);
nand U15339 (N_15339,N_10188,N_14583);
xor U15340 (N_15340,N_13260,N_14810);
or U15341 (N_15341,N_13829,N_13984);
nor U15342 (N_15342,N_14112,N_12438);
and U15343 (N_15343,N_11629,N_10596);
xor U15344 (N_15344,N_11896,N_11583);
or U15345 (N_15345,N_13194,N_12664);
nor U15346 (N_15346,N_13315,N_13168);
nand U15347 (N_15347,N_12171,N_11293);
and U15348 (N_15348,N_11829,N_14705);
and U15349 (N_15349,N_11797,N_14682);
or U15350 (N_15350,N_10126,N_12896);
nand U15351 (N_15351,N_14946,N_10731);
or U15352 (N_15352,N_14643,N_10368);
and U15353 (N_15353,N_14260,N_11606);
or U15354 (N_15354,N_12970,N_11301);
or U15355 (N_15355,N_10915,N_11385);
and U15356 (N_15356,N_14526,N_11072);
nor U15357 (N_15357,N_11180,N_14012);
or U15358 (N_15358,N_11632,N_10112);
or U15359 (N_15359,N_14523,N_10050);
xor U15360 (N_15360,N_10802,N_14600);
nand U15361 (N_15361,N_11483,N_11407);
nor U15362 (N_15362,N_14334,N_13423);
nand U15363 (N_15363,N_14414,N_13394);
and U15364 (N_15364,N_11741,N_14620);
xnor U15365 (N_15365,N_11972,N_14710);
xor U15366 (N_15366,N_10867,N_13581);
nor U15367 (N_15367,N_14846,N_13778);
and U15368 (N_15368,N_12299,N_11757);
xnor U15369 (N_15369,N_10708,N_14302);
xor U15370 (N_15370,N_14652,N_11162);
xnor U15371 (N_15371,N_13850,N_12844);
nor U15372 (N_15372,N_12341,N_13004);
and U15373 (N_15373,N_10215,N_13839);
xnor U15374 (N_15374,N_11512,N_13009);
and U15375 (N_15375,N_12686,N_14812);
or U15376 (N_15376,N_14207,N_13544);
or U15377 (N_15377,N_13748,N_14408);
and U15378 (N_15378,N_12001,N_14849);
nor U15379 (N_15379,N_14473,N_10375);
nor U15380 (N_15380,N_12403,N_12650);
xnor U15381 (N_15381,N_10979,N_13585);
and U15382 (N_15382,N_11042,N_10951);
xnor U15383 (N_15383,N_10114,N_11767);
xor U15384 (N_15384,N_10500,N_13678);
or U15385 (N_15385,N_11081,N_12173);
nand U15386 (N_15386,N_14785,N_10143);
nand U15387 (N_15387,N_11831,N_12636);
nand U15388 (N_15388,N_11399,N_13907);
nand U15389 (N_15389,N_13104,N_13236);
nand U15390 (N_15390,N_12981,N_11435);
or U15391 (N_15391,N_11190,N_11516);
xnor U15392 (N_15392,N_14318,N_13434);
or U15393 (N_15393,N_13181,N_11626);
nand U15394 (N_15394,N_14660,N_10201);
nand U15395 (N_15395,N_14603,N_13497);
and U15396 (N_15396,N_12979,N_13035);
and U15397 (N_15397,N_10798,N_12956);
and U15398 (N_15398,N_11586,N_13665);
nor U15399 (N_15399,N_12125,N_12228);
or U15400 (N_15400,N_14750,N_11678);
or U15401 (N_15401,N_11013,N_10465);
nor U15402 (N_15402,N_12038,N_12587);
nor U15403 (N_15403,N_12015,N_14025);
xnor U15404 (N_15404,N_14285,N_12960);
nand U15405 (N_15405,N_14143,N_12871);
nand U15406 (N_15406,N_14587,N_13908);
xor U15407 (N_15407,N_12054,N_13214);
and U15408 (N_15408,N_11223,N_11919);
nor U15409 (N_15409,N_14876,N_12851);
or U15410 (N_15410,N_12259,N_12961);
xor U15411 (N_15411,N_11166,N_10380);
or U15412 (N_15412,N_11010,N_11314);
nor U15413 (N_15413,N_10700,N_13802);
nand U15414 (N_15414,N_10503,N_12752);
nor U15415 (N_15415,N_10360,N_11475);
nand U15416 (N_15416,N_11050,N_11848);
or U15417 (N_15417,N_14462,N_13160);
nor U15418 (N_15418,N_14977,N_11861);
nor U15419 (N_15419,N_14350,N_11887);
or U15420 (N_15420,N_11419,N_11489);
nand U15421 (N_15421,N_12193,N_12200);
nor U15422 (N_15422,N_14697,N_14406);
nor U15423 (N_15423,N_12561,N_14696);
and U15424 (N_15424,N_10250,N_13396);
and U15425 (N_15425,N_14760,N_13945);
nor U15426 (N_15426,N_12018,N_14301);
or U15427 (N_15427,N_12809,N_10587);
or U15428 (N_15428,N_11935,N_14109);
xnor U15429 (N_15429,N_11356,N_13385);
xnor U15430 (N_15430,N_14566,N_13372);
and U15431 (N_15431,N_14925,N_10124);
nand U15432 (N_15432,N_11837,N_14452);
or U15433 (N_15433,N_14886,N_12178);
or U15434 (N_15434,N_12055,N_10485);
nor U15435 (N_15435,N_10472,N_12646);
nand U15436 (N_15436,N_14376,N_13738);
or U15437 (N_15437,N_12966,N_11695);
nand U15438 (N_15438,N_11747,N_12504);
or U15439 (N_15439,N_12997,N_11446);
nor U15440 (N_15440,N_12457,N_10746);
and U15441 (N_15441,N_12434,N_10371);
nand U15442 (N_15442,N_10724,N_13699);
and U15443 (N_15443,N_14854,N_14120);
nand U15444 (N_15444,N_11842,N_13264);
xor U15445 (N_15445,N_10106,N_13205);
xor U15446 (N_15446,N_11304,N_10579);
nand U15447 (N_15447,N_10128,N_10251);
nand U15448 (N_15448,N_10983,N_10231);
xnor U15449 (N_15449,N_13591,N_13117);
xnor U15450 (N_15450,N_12111,N_11441);
nand U15451 (N_15451,N_14641,N_11689);
and U15452 (N_15452,N_13799,N_14247);
nor U15453 (N_15453,N_10823,N_10093);
nor U15454 (N_15454,N_14577,N_13115);
or U15455 (N_15455,N_12617,N_13263);
nand U15456 (N_15456,N_11210,N_12590);
or U15457 (N_15457,N_14257,N_13773);
nand U15458 (N_15458,N_10297,N_13806);
xnor U15459 (N_15459,N_13924,N_12861);
xnor U15460 (N_15460,N_12061,N_12401);
and U15461 (N_15461,N_14806,N_14691);
nand U15462 (N_15462,N_14370,N_12012);
or U15463 (N_15463,N_11421,N_13906);
and U15464 (N_15464,N_12624,N_10717);
nand U15465 (N_15465,N_13897,N_12492);
xor U15466 (N_15466,N_12565,N_10730);
nand U15467 (N_15467,N_13618,N_14561);
nand U15468 (N_15468,N_14329,N_10055);
xor U15469 (N_15469,N_10815,N_14599);
xor U15470 (N_15470,N_12452,N_13882);
nand U15471 (N_15471,N_11903,N_11355);
and U15472 (N_15472,N_12248,N_13086);
xnor U15473 (N_15473,N_13169,N_11203);
nor U15474 (N_15474,N_14278,N_11562);
xnor U15475 (N_15475,N_10358,N_11053);
and U15476 (N_15476,N_12160,N_12948);
and U15477 (N_15477,N_12690,N_11146);
and U15478 (N_15478,N_10513,N_14623);
or U15479 (N_15479,N_11977,N_12042);
nor U15480 (N_15480,N_14293,N_13734);
xor U15481 (N_15481,N_11302,N_11716);
or U15482 (N_15482,N_11867,N_10505);
or U15483 (N_15483,N_10021,N_14507);
or U15484 (N_15484,N_10613,N_11690);
nor U15485 (N_15485,N_14146,N_12129);
nor U15486 (N_15486,N_14997,N_14054);
and U15487 (N_15487,N_13822,N_14743);
nor U15488 (N_15488,N_13502,N_13768);
nand U15489 (N_15489,N_10971,N_14124);
and U15490 (N_15490,N_14477,N_14344);
and U15491 (N_15491,N_13144,N_11756);
or U15492 (N_15492,N_13631,N_13571);
xnor U15493 (N_15493,N_10340,N_13411);
and U15494 (N_15494,N_14281,N_14033);
xnor U15495 (N_15495,N_12150,N_10831);
xnor U15496 (N_15496,N_12300,N_14879);
or U15497 (N_15497,N_10748,N_14138);
or U15498 (N_15498,N_10283,N_12235);
nand U15499 (N_15499,N_10618,N_12778);
or U15500 (N_15500,N_10709,N_13295);
nor U15501 (N_15501,N_14171,N_12295);
or U15502 (N_15502,N_14364,N_10213);
xor U15503 (N_15503,N_12052,N_14619);
nand U15504 (N_15504,N_14127,N_11597);
nor U15505 (N_15505,N_12951,N_12002);
xor U15506 (N_15506,N_12240,N_12294);
xnor U15507 (N_15507,N_10588,N_14763);
and U15508 (N_15508,N_14544,N_11795);
nand U15509 (N_15509,N_12642,N_13657);
xor U15510 (N_15510,N_10680,N_13447);
and U15511 (N_15511,N_11813,N_11165);
and U15512 (N_15512,N_12120,N_14144);
nand U15513 (N_15513,N_13489,N_13320);
nor U15514 (N_15514,N_10492,N_14131);
nor U15515 (N_15515,N_12867,N_13370);
or U15516 (N_15516,N_12783,N_13549);
nand U15517 (N_15517,N_11238,N_13471);
nand U15518 (N_15518,N_11443,N_12188);
or U15519 (N_15519,N_14982,N_13770);
or U15520 (N_15520,N_10212,N_11083);
nor U15521 (N_15521,N_11513,N_14457);
and U15522 (N_15522,N_14361,N_12499);
nand U15523 (N_15523,N_11832,N_11953);
nor U15524 (N_15524,N_13974,N_14397);
nor U15525 (N_15525,N_11476,N_10789);
nand U15526 (N_15526,N_14695,N_12724);
xnor U15527 (N_15527,N_11431,N_12432);
nand U15528 (N_15528,N_10441,N_14426);
nor U15529 (N_15529,N_13284,N_13750);
or U15530 (N_15530,N_13099,N_13386);
nor U15531 (N_15531,N_13042,N_11261);
or U15532 (N_15532,N_13479,N_12837);
nor U15533 (N_15533,N_13094,N_11894);
or U15534 (N_15534,N_12999,N_11956);
or U15535 (N_15535,N_13245,N_14438);
xor U15536 (N_15536,N_12839,N_11877);
or U15537 (N_15537,N_10811,N_12697);
nand U15538 (N_15538,N_11058,N_10840);
xor U15539 (N_15539,N_12782,N_11720);
or U15540 (N_15540,N_14119,N_14228);
and U15541 (N_15541,N_11791,N_11612);
nand U15542 (N_15542,N_12753,N_12035);
or U15543 (N_15543,N_12165,N_12539);
nand U15544 (N_15544,N_12645,N_12813);
nor U15545 (N_15545,N_12716,N_14279);
nor U15546 (N_15546,N_10686,N_14948);
nor U15547 (N_15547,N_11303,N_12381);
xor U15548 (N_15548,N_12166,N_14673);
nand U15549 (N_15549,N_10562,N_10516);
nor U15550 (N_15550,N_13543,N_12682);
xnor U15551 (N_15551,N_10197,N_12026);
or U15552 (N_15552,N_11163,N_14062);
or U15553 (N_15553,N_13294,N_14308);
and U15554 (N_15554,N_10778,N_10950);
and U15555 (N_15555,N_12258,N_12557);
or U15556 (N_15556,N_12291,N_12918);
and U15557 (N_15557,N_13271,N_13440);
and U15558 (N_15558,N_12450,N_10043);
xor U15559 (N_15559,N_14254,N_14545);
xnor U15560 (N_15560,N_11367,N_12962);
xor U15561 (N_15561,N_13953,N_12741);
nor U15562 (N_15562,N_12350,N_11432);
and U15563 (N_15563,N_10257,N_13238);
and U15564 (N_15564,N_10642,N_14875);
xor U15565 (N_15565,N_10652,N_10550);
xnor U15566 (N_15566,N_10300,N_14496);
and U15567 (N_15567,N_10549,N_13065);
nand U15568 (N_15568,N_10498,N_12622);
and U15569 (N_15569,N_10477,N_11241);
xor U15570 (N_15570,N_13955,N_12777);
and U15571 (N_15571,N_11684,N_11029);
nand U15572 (N_15572,N_10922,N_14490);
nand U15573 (N_15573,N_12592,N_14655);
and U15574 (N_15574,N_11635,N_11859);
xnor U15575 (N_15575,N_12974,N_12853);
and U15576 (N_15576,N_11159,N_13222);
and U15577 (N_15577,N_11229,N_10373);
nand U15578 (N_15578,N_12734,N_10907);
and U15579 (N_15579,N_10537,N_13162);
xnor U15580 (N_15580,N_10042,N_12031);
nor U15581 (N_15581,N_13124,N_12497);
nand U15582 (N_15582,N_13167,N_10265);
xor U15583 (N_15583,N_12852,N_10137);
or U15584 (N_15584,N_10870,N_14009);
and U15585 (N_15585,N_14644,N_11589);
or U15586 (N_15586,N_14758,N_12000);
nor U15587 (N_15587,N_14769,N_10661);
nand U15588 (N_15588,N_14965,N_14069);
xor U15589 (N_15589,N_14092,N_10755);
or U15590 (N_15590,N_12412,N_11560);
xor U15591 (N_15591,N_12556,N_13256);
nand U15592 (N_15592,N_12107,N_10479);
xnor U15593 (N_15593,N_14129,N_10483);
nand U15594 (N_15594,N_10409,N_11055);
nand U15595 (N_15595,N_13775,N_12264);
nor U15596 (N_15596,N_12520,N_10518);
or U15597 (N_15597,N_11945,N_13913);
and U15598 (N_15598,N_10010,N_10310);
nand U15599 (N_15599,N_11440,N_11363);
xnor U15600 (N_15600,N_13705,N_13686);
or U15601 (N_15601,N_13739,N_11403);
xnor U15602 (N_15602,N_10929,N_13998);
or U15603 (N_15603,N_10317,N_12775);
and U15604 (N_15604,N_11139,N_13529);
nand U15605 (N_15605,N_14103,N_10298);
xnor U15606 (N_15606,N_12927,N_12903);
and U15607 (N_15607,N_12593,N_11282);
xor U15608 (N_15608,N_12842,N_14356);
and U15609 (N_15609,N_14745,N_11099);
and U15610 (N_15610,N_14489,N_11428);
nor U15611 (N_15611,N_13528,N_11454);
nand U15612 (N_15612,N_13838,N_12428);
nor U15613 (N_15613,N_11211,N_12555);
xor U15614 (N_15614,N_11607,N_14286);
nor U15615 (N_15615,N_14383,N_12524);
and U15616 (N_15616,N_12116,N_14128);
or U15617 (N_15617,N_14341,N_12325);
nor U15618 (N_15618,N_13735,N_10773);
xnor U15619 (N_15619,N_14726,N_14485);
or U15620 (N_15620,N_14746,N_13317);
nor U15621 (N_15621,N_12554,N_14421);
nand U15622 (N_15622,N_14439,N_10245);
nand U15623 (N_15623,N_11610,N_13306);
nor U15624 (N_15624,N_10254,N_11816);
xnor U15625 (N_15625,N_12159,N_14150);
and U15626 (N_15626,N_10590,N_14256);
nor U15627 (N_15627,N_11749,N_14764);
and U15628 (N_15628,N_14217,N_12451);
and U15629 (N_15629,N_11671,N_14481);
nand U15630 (N_15630,N_12315,N_12727);
nand U15631 (N_15631,N_12538,N_11623);
and U15632 (N_15632,N_13537,N_14853);
and U15633 (N_15633,N_12409,N_12301);
or U15634 (N_15634,N_12869,N_10923);
and U15635 (N_15635,N_14068,N_11245);
nor U15636 (N_15636,N_13347,N_14230);
nand U15637 (N_15637,N_13296,N_13671);
nand U15638 (N_15638,N_10383,N_14918);
nor U15639 (N_15639,N_11501,N_10361);
nor U15640 (N_15640,N_13250,N_13381);
or U15641 (N_15641,N_14535,N_10806);
nor U15642 (N_15642,N_11177,N_10379);
nand U15643 (N_15643,N_10614,N_13364);
and U15644 (N_15644,N_11789,N_11488);
xor U15645 (N_15645,N_12312,N_12025);
xor U15646 (N_15646,N_13431,N_13875);
or U15647 (N_15647,N_11572,N_14411);
xnor U15648 (N_15648,N_11885,N_13097);
nor U15649 (N_15649,N_10400,N_11827);
or U15650 (N_15650,N_14761,N_12201);
and U15651 (N_15651,N_10421,N_11853);
or U15652 (N_15652,N_14081,N_10163);
and U15653 (N_15653,N_12616,N_12854);
or U15654 (N_15654,N_13879,N_13119);
or U15655 (N_15655,N_11648,N_12631);
nand U15656 (N_15656,N_13697,N_10631);
and U15657 (N_15657,N_13496,N_14650);
nand U15658 (N_15658,N_10325,N_13266);
xor U15659 (N_15659,N_11185,N_14130);
nor U15660 (N_15660,N_11545,N_11593);
xor U15661 (N_15661,N_12667,N_10905);
xor U15662 (N_15662,N_14692,N_11578);
xnor U15663 (N_15663,N_12507,N_10177);
and U15664 (N_15664,N_10393,N_11911);
or U15665 (N_15665,N_13915,N_13807);
and U15666 (N_15666,N_14661,N_14685);
nand U15667 (N_15667,N_11043,N_14533);
nor U15668 (N_15668,N_13335,N_14232);
nand U15669 (N_15669,N_14101,N_10407);
xor U15670 (N_15670,N_12881,N_10578);
nand U15671 (N_15671,N_13400,N_14639);
xor U15672 (N_15672,N_14472,N_14372);
and U15673 (N_15673,N_14993,N_11221);
nor U15674 (N_15674,N_11343,N_13200);
nor U15675 (N_15675,N_14390,N_10344);
nor U15676 (N_15676,N_10632,N_12759);
nand U15677 (N_15677,N_14118,N_11248);
xor U15678 (N_15678,N_13643,N_10035);
nand U15679 (N_15679,N_11002,N_13719);
nand U15680 (N_15680,N_14259,N_11889);
xor U15681 (N_15681,N_12276,N_10110);
and U15682 (N_15682,N_14844,N_11169);
and U15683 (N_15683,N_11807,N_10918);
and U15684 (N_15684,N_11868,N_14430);
and U15685 (N_15685,N_13063,N_12132);
nand U15686 (N_15686,N_13438,N_13450);
and U15687 (N_15687,N_14548,N_11995);
xnor U15688 (N_15688,N_10244,N_12455);
nand U15689 (N_15689,N_14829,N_10635);
and U15690 (N_15690,N_11731,N_13523);
and U15691 (N_15691,N_12421,N_14454);
xnor U15692 (N_15692,N_11920,N_12313);
and U15693 (N_15693,N_12911,N_12989);
nand U15694 (N_15694,N_10068,N_10666);
or U15695 (N_15695,N_13718,N_11698);
xnor U15696 (N_15696,N_10595,N_11891);
nor U15697 (N_15697,N_10016,N_13087);
xor U15698 (N_15698,N_14640,N_12913);
nor U15699 (N_15699,N_13808,N_10563);
xnor U15700 (N_15700,N_12365,N_12692);
or U15701 (N_15701,N_11415,N_10630);
xor U15702 (N_15702,N_10403,N_13827);
and U15703 (N_15703,N_14564,N_13078);
or U15704 (N_15704,N_14040,N_11322);
nand U15705 (N_15705,N_14072,N_10955);
and U15706 (N_15706,N_14090,N_11878);
or U15707 (N_15707,N_11990,N_12386);
nor U15708 (N_15708,N_13747,N_14017);
or U15709 (N_15709,N_10525,N_11000);
nor U15710 (N_15710,N_11722,N_10019);
nor U15711 (N_15711,N_10790,N_10863);
and U15712 (N_15712,N_13958,N_14647);
nor U15713 (N_15713,N_10183,N_10767);
and U15714 (N_15714,N_12823,N_11815);
or U15715 (N_15715,N_11247,N_14532);
or U15716 (N_15716,N_13644,N_12513);
or U15717 (N_15717,N_14771,N_13061);
and U15718 (N_15718,N_13197,N_11905);
xnor U15719 (N_15719,N_10456,N_14328);
xor U15720 (N_15720,N_10447,N_10612);
nand U15721 (N_15721,N_11027,N_10336);
or U15722 (N_15722,N_13093,N_10653);
and U15723 (N_15723,N_12181,N_10713);
or U15724 (N_15724,N_13244,N_10779);
nor U15725 (N_15725,N_12811,N_13108);
or U15726 (N_15726,N_11581,N_12396);
xor U15727 (N_15727,N_11630,N_14900);
or U15728 (N_15728,N_13714,N_13180);
xor U15729 (N_15729,N_12468,N_14237);
nor U15730 (N_15730,N_11183,N_13625);
and U15731 (N_15731,N_10679,N_14142);
nand U15732 (N_15732,N_14748,N_14348);
or U15733 (N_15733,N_10609,N_14465);
or U15734 (N_15734,N_11391,N_11307);
nor U15735 (N_15735,N_10487,N_10545);
nand U15736 (N_15736,N_14428,N_12633);
and U15737 (N_15737,N_14834,N_12197);
nand U15738 (N_15738,N_11389,N_13388);
or U15739 (N_15739,N_11786,N_14291);
or U15740 (N_15740,N_10025,N_12749);
xnor U15741 (N_15741,N_14220,N_14137);
nor U15742 (N_15742,N_12246,N_13384);
or U15743 (N_15743,N_14194,N_14913);
or U15744 (N_15744,N_13182,N_11339);
xor U15745 (N_15745,N_13516,N_10063);
xor U15746 (N_15746,N_10801,N_13232);
nor U15747 (N_15747,N_14956,N_14113);
or U15748 (N_15748,N_14365,N_11439);
nand U15749 (N_15749,N_12329,N_11500);
and U15750 (N_15750,N_14928,N_10699);
or U15751 (N_15751,N_12462,N_10930);
nand U15752 (N_15752,N_12933,N_12638);
or U15753 (N_15753,N_11077,N_10135);
or U15754 (N_15754,N_10807,N_14455);
nor U15755 (N_15755,N_12371,N_12832);
nor U15756 (N_15756,N_13218,N_10756);
and U15757 (N_15757,N_12841,N_11469);
xor U15758 (N_15758,N_14028,N_10001);
nand U15759 (N_15759,N_11840,N_10446);
or U15760 (N_15760,N_12514,N_13310);
nor U15761 (N_15761,N_12916,N_14316);
nor U15762 (N_15762,N_14100,N_12758);
nand U15763 (N_15763,N_14500,N_10671);
nand U15764 (N_15764,N_13380,N_10780);
or U15765 (N_15765,N_12681,N_13322);
xor U15766 (N_15766,N_13780,N_14531);
and U15767 (N_15767,N_13650,N_10051);
xor U15768 (N_15768,N_13270,N_12045);
nand U15769 (N_15769,N_14804,N_13597);
xor U15770 (N_15770,N_14605,N_10504);
or U15771 (N_15771,N_11128,N_11590);
or U15772 (N_15772,N_11445,N_12710);
nand U15773 (N_15773,N_12525,N_14450);
and U15774 (N_15774,N_12427,N_10646);
nor U15775 (N_15775,N_10203,N_13446);
nor U15776 (N_15776,N_11198,N_11117);
xnor U15777 (N_15777,N_11773,N_11161);
nand U15778 (N_15778,N_12795,N_12420);
nor U15779 (N_15779,N_10795,N_10439);
or U15780 (N_15780,N_12221,N_14321);
nand U15781 (N_15781,N_14043,N_12411);
nor U15782 (N_15782,N_11553,N_11232);
xor U15783 (N_15783,N_14632,N_14309);
and U15784 (N_15784,N_12397,N_13461);
nor U15785 (N_15785,N_11855,N_14569);
or U15786 (N_15786,N_14187,N_10308);
and U15787 (N_15787,N_10480,N_12945);
and U15788 (N_15788,N_11090,N_10326);
and U15789 (N_15789,N_14618,N_12521);
nor U15790 (N_15790,N_13753,N_13977);
nand U15791 (N_15791,N_14110,N_10638);
and U15792 (N_15792,N_11306,N_14255);
and U15793 (N_15793,N_10037,N_13353);
nand U15794 (N_15794,N_10546,N_14850);
or U15795 (N_15795,N_13522,N_11933);
nand U15796 (N_15796,N_12234,N_10083);
and U15797 (N_15797,N_10331,N_13531);
and U15798 (N_15798,N_14055,N_10350);
xor U15799 (N_15799,N_11160,N_13858);
nand U15800 (N_15800,N_13916,N_12822);
and U15801 (N_15801,N_12109,N_11470);
nand U15802 (N_15802,N_13131,N_13365);
nand U15803 (N_15803,N_10538,N_12921);
xnor U15804 (N_15804,N_12261,N_10216);
xnor U15805 (N_15805,N_12134,N_10702);
or U15806 (N_15806,N_13598,N_12605);
nor U15807 (N_15807,N_12449,N_12931);
or U15808 (N_15808,N_12454,N_10323);
xnor U15809 (N_15809,N_11001,N_10880);
nand U15810 (N_15810,N_11328,N_12141);
xnor U15811 (N_15811,N_14005,N_10278);
or U15812 (N_15812,N_12940,N_13901);
or U15813 (N_15813,N_11272,N_13566);
nand U15814 (N_15814,N_11937,N_11373);
nand U15815 (N_15815,N_11189,N_14774);
or U15816 (N_15816,N_12318,N_10872);
nor U15817 (N_15817,N_12715,N_11721);
or U15818 (N_15818,N_14493,N_11156);
and U15819 (N_15819,N_11134,N_13847);
xnor U15820 (N_15820,N_12908,N_11520);
and U15821 (N_15821,N_10312,N_14064);
nand U15822 (N_15822,N_14627,N_11201);
and U15823 (N_15823,N_12523,N_12829);
nor U15824 (N_15824,N_13233,N_13470);
nand U15825 (N_15825,N_11714,N_10828);
nor U15826 (N_15826,N_14121,N_12346);
nand U15827 (N_15827,N_11740,N_10718);
and U15828 (N_15828,N_12021,N_14505);
xor U15829 (N_15829,N_14079,N_10845);
nand U15830 (N_15830,N_11703,N_13506);
xor U15831 (N_15831,N_13147,N_12273);
nor U15832 (N_15832,N_14615,N_10891);
xor U15833 (N_15833,N_13895,N_11939);
or U15834 (N_15834,N_13129,N_14036);
or U15835 (N_15835,N_13821,N_12926);
or U15836 (N_15836,N_12022,N_11987);
xnor U15837 (N_15837,N_14700,N_10190);
xnor U15838 (N_15838,N_12987,N_10732);
or U15839 (N_15839,N_10256,N_12907);
and U15840 (N_15840,N_10803,N_12102);
nand U15841 (N_15841,N_10914,N_12209);
and U15842 (N_15842,N_13301,N_10032);
xor U15843 (N_15843,N_11943,N_10706);
xor U15844 (N_15844,N_13455,N_11150);
nor U15845 (N_15845,N_13698,N_13805);
nor U15846 (N_15846,N_12079,N_13382);
xor U15847 (N_15847,N_13560,N_13592);
and U15848 (N_15848,N_13610,N_13339);
nor U15849 (N_15849,N_13830,N_12637);
nand U15850 (N_15850,N_10000,N_12477);
or U15851 (N_15851,N_11324,N_11341);
and U15852 (N_15852,N_14994,N_10576);
and U15853 (N_15853,N_11493,N_11138);
xor U15854 (N_15854,N_12792,N_11888);
nor U15855 (N_15855,N_10102,N_12430);
and U15856 (N_15856,N_14851,N_13067);
nor U15857 (N_15857,N_10639,N_10997);
or U15858 (N_15858,N_10899,N_10191);
xnor U15859 (N_15859,N_12673,N_10884);
xnor U15860 (N_15860,N_14078,N_11052);
nand U15861 (N_15861,N_14998,N_13900);
xnor U15862 (N_15862,N_13608,N_11425);
or U15863 (N_15863,N_10004,N_13075);
xnor U15864 (N_15864,N_13467,N_11127);
or U15865 (N_15865,N_13948,N_14195);
nand U15866 (N_15866,N_13449,N_14687);
xor U15867 (N_15867,N_13208,N_13865);
nor U15868 (N_15868,N_14014,N_10825);
and U15869 (N_15869,N_11841,N_12598);
nand U15870 (N_15870,N_10261,N_11808);
nand U15871 (N_15871,N_12463,N_10140);
or U15872 (N_15872,N_11318,N_10527);
nand U15873 (N_15873,N_11236,N_13416);
and U15874 (N_15874,N_13638,N_12968);
and U15875 (N_15875,N_14581,N_12744);
nor U15876 (N_15876,N_14649,N_10189);
xor U15877 (N_15877,N_12818,N_11508);
or U15878 (N_15878,N_10382,N_10861);
or U15879 (N_15879,N_11179,N_12720);
xor U15880 (N_15880,N_12522,N_10817);
nor U15881 (N_15881,N_10376,N_13483);
and U15882 (N_15882,N_13762,N_13885);
nand U15883 (N_15883,N_13176,N_14335);
nor U15884 (N_15884,N_10649,N_10433);
nand U15885 (N_15885,N_12304,N_11492);
nand U15886 (N_15886,N_11826,N_14141);
xnor U15887 (N_15887,N_14104,N_13490);
or U15888 (N_15888,N_14271,N_14675);
xor U15889 (N_15889,N_10799,N_12860);
and U15890 (N_15890,N_14775,N_14223);
xnor U15891 (N_15891,N_12582,N_10108);
and U15892 (N_15892,N_13417,N_10311);
xnor U15893 (N_15893,N_13242,N_10670);
nand U15894 (N_15894,N_14773,N_13454);
and U15895 (N_15895,N_11715,N_12657);
xnor U15896 (N_15896,N_10819,N_14441);
xor U15897 (N_15897,N_14961,N_10841);
xnor U15898 (N_15898,N_13359,N_12895);
nand U15899 (N_15899,N_10289,N_10508);
or U15900 (N_15900,N_14389,N_12333);
or U15901 (N_15901,N_10028,N_10557);
xnor U15902 (N_15902,N_13933,N_13059);
or U15903 (N_15903,N_13503,N_12088);
xor U15904 (N_15904,N_14958,N_14718);
or U15905 (N_15905,N_14927,N_13161);
xor U15906 (N_15906,N_12619,N_11184);
nand U15907 (N_15907,N_14719,N_14467);
nand U15908 (N_15908,N_11567,N_10381);
nand U15909 (N_15909,N_12044,N_13183);
nor U15910 (N_15910,N_10535,N_10451);
nand U15911 (N_15911,N_11550,N_12615);
nand U15912 (N_15912,N_11799,N_13103);
or U15913 (N_15913,N_13466,N_12091);
and U15914 (N_15914,N_10430,N_10496);
nor U15915 (N_15915,N_11267,N_11340);
nor U15916 (N_15916,N_11834,N_11748);
xor U15917 (N_15917,N_10848,N_14932);
xor U15918 (N_15918,N_10018,N_12168);
and U15919 (N_15919,N_10976,N_10804);
and U15920 (N_15920,N_13258,N_13371);
or U15921 (N_15921,N_11975,N_12051);
and U15922 (N_15922,N_10677,N_10984);
xor U15923 (N_15923,N_10367,N_10753);
and U15924 (N_15924,N_12279,N_14410);
xor U15925 (N_15925,N_13010,N_10464);
xor U15926 (N_15926,N_10287,N_10548);
nor U15927 (N_15927,N_14570,N_11008);
or U15928 (N_15928,N_12781,N_14606);
nor U15929 (N_15929,N_11803,N_13843);
nor U15930 (N_15930,N_14975,N_10992);
nand U15931 (N_15931,N_14945,N_11776);
and U15932 (N_15932,N_12589,N_13562);
nand U15933 (N_15933,N_12801,N_14339);
nand U15934 (N_15934,N_12957,N_14903);
nand U15935 (N_15935,N_12210,N_12847);
xor U15936 (N_15936,N_14057,N_13172);
nand U15937 (N_15937,N_10837,N_12838);
nor U15938 (N_15938,N_13122,N_14074);
nor U15939 (N_15939,N_13283,N_13148);
nor U15940 (N_15940,N_14616,N_10070);
or U15941 (N_15941,N_11196,N_13185);
nand U15942 (N_15942,N_12220,N_13357);
nor U15943 (N_15943,N_10450,N_12284);
and U15944 (N_15944,N_13032,N_13358);
or U15945 (N_15945,N_13545,N_14847);
and U15946 (N_15946,N_14460,N_13498);
xor U15947 (N_15947,N_14440,N_14817);
or U15948 (N_15948,N_12641,N_13019);
nor U15949 (N_15949,N_10088,N_10240);
nand U15950 (N_15950,N_13418,N_13100);
xor U15951 (N_15951,N_13316,N_13685);
nand U15952 (N_15952,N_11947,N_14197);
nand U15953 (N_15953,N_12949,N_11644);
nor U15954 (N_15954,N_13630,N_12630);
nor U15955 (N_15955,N_13509,N_10925);
nand U15956 (N_15956,N_14908,N_11760);
xor U15957 (N_15957,N_10180,N_14917);
and U15958 (N_15958,N_10053,N_10759);
and U15959 (N_15959,N_14242,N_10328);
nor U15960 (N_15960,N_13302,N_12676);
xor U15961 (N_15961,N_11406,N_11732);
and U15962 (N_15962,N_14445,N_13563);
and U15963 (N_15963,N_13435,N_13851);
nand U15964 (N_15964,N_14501,N_13584);
or U15965 (N_15965,N_13763,N_10741);
nor U15966 (N_15966,N_11628,N_12227);
or U15967 (N_15967,N_13996,N_12859);
and U15968 (N_15968,N_11869,N_11070);
nand U15969 (N_15969,N_14662,N_14819);
nor U15970 (N_15970,N_13060,N_10911);
xnor U15971 (N_15971,N_13800,N_14985);
or U15972 (N_15972,N_12424,N_14003);
and U15973 (N_15973,N_14608,N_10428);
nand U15974 (N_15974,N_11397,N_11857);
nor U15975 (N_15975,N_12345,N_12779);
or U15976 (N_15976,N_13328,N_10046);
and U15977 (N_15977,N_14097,N_13878);
xor U15978 (N_15978,N_12138,N_11573);
nor U15979 (N_15979,N_14676,N_10924);
and U15980 (N_15980,N_12144,N_12456);
xor U15981 (N_15981,N_13051,N_14828);
or U15982 (N_15982,N_13777,N_12425);
xor U15983 (N_15983,N_11330,N_14082);
xor U15984 (N_15984,N_11575,N_14680);
and U15985 (N_15985,N_11228,N_13709);
nand U15986 (N_15986,N_10170,N_12919);
and U15987 (N_15987,N_12140,N_14322);
and U15988 (N_15988,N_10158,N_14456);
xor U15989 (N_15989,N_13378,N_11666);
nand U15990 (N_15990,N_14487,N_14277);
nor U15991 (N_15991,N_10193,N_14044);
xnor U15992 (N_15992,N_14444,N_12289);
or U15993 (N_15993,N_14559,N_14274);
or U15994 (N_15994,N_14742,N_10830);
or U15995 (N_15995,N_11233,N_10669);
and U15996 (N_15996,N_14568,N_12529);
nor U15997 (N_15997,N_11471,N_11814);
nand U15998 (N_15998,N_14722,N_11297);
nand U15999 (N_15999,N_13519,N_11103);
and U16000 (N_16000,N_10723,N_10577);
or U16001 (N_16001,N_14499,N_12774);
xor U16002 (N_16002,N_13946,N_12644);
nand U16003 (N_16003,N_11609,N_14244);
xnor U16004 (N_16004,N_14139,N_12364);
xnor U16005 (N_16005,N_14892,N_10932);
and U16006 (N_16006,N_13980,N_11692);
nor U16007 (N_16007,N_12917,N_11252);
and U16008 (N_16008,N_13619,N_12988);
or U16009 (N_16009,N_14549,N_11662);
or U16010 (N_16010,N_12721,N_12399);
or U16011 (N_16011,N_14049,N_13041);
or U16012 (N_16012,N_11819,N_13629);
nor U16013 (N_16013,N_11963,N_10423);
nor U16014 (N_16014,N_10667,N_14508);
nand U16015 (N_16015,N_11078,N_11351);
nand U16016 (N_16016,N_13937,N_11009);
xor U16017 (N_16017,N_14497,N_11528);
nand U16018 (N_16018,N_11016,N_14679);
and U16019 (N_16019,N_10560,N_12122);
xor U16020 (N_16020,N_14614,N_14955);
or U16021 (N_16021,N_11167,N_12360);
nand U16022 (N_16022,N_14226,N_12572);
nor U16023 (N_16023,N_10166,N_10598);
nor U16024 (N_16024,N_14343,N_10762);
xor U16025 (N_16025,N_12634,N_13030);
and U16026 (N_16026,N_13187,N_11015);
xnor U16027 (N_16027,N_11551,N_13786);
nand U16028 (N_16028,N_10281,N_10399);
nor U16029 (N_16029,N_11381,N_10094);
nor U16030 (N_16030,N_10651,N_11467);
nand U16031 (N_16031,N_11910,N_13812);
nand U16032 (N_16032,N_14571,N_10481);
and U16033 (N_16033,N_13820,N_12243);
xor U16034 (N_16034,N_14369,N_14283);
xnor U16035 (N_16035,N_13736,N_10747);
nand U16036 (N_16036,N_10248,N_14122);
nor U16037 (N_16037,N_10953,N_13341);
or U16038 (N_16038,N_14885,N_13848);
and U16039 (N_16039,N_12519,N_12878);
or U16040 (N_16040,N_10601,N_11359);
nor U16041 (N_16041,N_12472,N_11918);
xnor U16042 (N_16042,N_10766,N_12947);
and U16043 (N_16043,N_13462,N_14941);
and U16044 (N_16044,N_10277,N_12460);
nor U16045 (N_16045,N_11541,N_12048);
or U16046 (N_16046,N_10725,N_10148);
or U16047 (N_16047,N_11255,N_10920);
xor U16048 (N_16048,N_11525,N_12340);
and U16049 (N_16049,N_13918,N_14258);
xor U16050 (N_16050,N_10581,N_12003);
nor U16051 (N_16051,N_14310,N_11879);
nand U16052 (N_16052,N_12155,N_13356);
and U16053 (N_16053,N_13669,N_13321);
xor U16054 (N_16054,N_13716,N_14289);
xor U16055 (N_16055,N_11291,N_13444);
and U16056 (N_16056,N_13488,N_13098);
xor U16057 (N_16057,N_10056,N_10933);
and U16058 (N_16058,N_13179,N_14708);
nand U16059 (N_16059,N_14782,N_13406);
or U16060 (N_16060,N_14269,N_13084);
xor U16061 (N_16061,N_12771,N_10435);
nand U16062 (N_16062,N_11327,N_14690);
and U16063 (N_16063,N_14584,N_10697);
nand U16064 (N_16064,N_10497,N_11332);
nor U16065 (N_16065,N_12036,N_14574);
xor U16066 (N_16066,N_13782,N_13109);
nor U16067 (N_16067,N_12991,N_11707);
nor U16068 (N_16068,N_11779,N_14642);
xnor U16069 (N_16069,N_14954,N_10892);
nor U16070 (N_16070,N_12906,N_11785);
or U16071 (N_16071,N_11112,N_11938);
or U16072 (N_16072,N_12208,N_14360);
nand U16073 (N_16073,N_12113,N_13031);
xnor U16074 (N_16074,N_14836,N_13804);
nand U16075 (N_16075,N_12101,N_10222);
xnor U16076 (N_16076,N_11526,N_13927);
nand U16077 (N_16077,N_11922,N_10176);
and U16078 (N_16078,N_10589,N_14403);
nand U16079 (N_16079,N_14896,N_13419);
or U16080 (N_16080,N_14075,N_10812);
xor U16081 (N_16081,N_14164,N_14371);
nand U16082 (N_16082,N_13202,N_14882);
nand U16083 (N_16083,N_12306,N_14624);
xnor U16084 (N_16084,N_13410,N_13272);
or U16085 (N_16085,N_14536,N_11212);
xnor U16086 (N_16086,N_12812,N_12285);
nand U16087 (N_16087,N_13558,N_12824);
nand U16088 (N_16088,N_13564,N_12902);
xnor U16089 (N_16089,N_12239,N_14333);
nand U16090 (N_16090,N_11828,N_14297);
nor U16091 (N_16091,N_13607,N_13401);
nor U16092 (N_16092,N_10866,N_11395);
or U16093 (N_16093,N_11634,N_14702);
xor U16094 (N_16094,N_10705,N_11523);
and U16095 (N_16095,N_14575,N_13510);
or U16096 (N_16096,N_12269,N_10453);
nand U16097 (N_16097,N_10988,N_10685);
and U16098 (N_16098,N_10816,N_10941);
or U16099 (N_16099,N_12186,N_10493);
nor U16100 (N_16100,N_13711,N_10475);
xor U16101 (N_16101,N_10279,N_10559);
xor U16102 (N_16102,N_14755,N_10228);
xnor U16103 (N_16103,N_13904,N_13604);
and U16104 (N_16104,N_14634,N_12959);
and U16105 (N_16105,N_12694,N_12330);
nor U16106 (N_16106,N_14094,N_10975);
and U16107 (N_16107,N_14749,N_14114);
nor U16108 (N_16108,N_10200,N_11924);
or U16109 (N_16109,N_13343,N_10869);
nor U16110 (N_16110,N_11954,N_14741);
or U16111 (N_16111,N_12043,N_11923);
or U16112 (N_16112,N_14645,N_12394);
and U16113 (N_16113,N_13587,N_10405);
or U16114 (N_16114,N_11463,N_11967);
xnor U16115 (N_16115,N_10619,N_10532);
or U16116 (N_16116,N_12118,N_11548);
and U16117 (N_16117,N_10926,N_11651);
nor U16118 (N_16118,N_10827,N_12489);
xnor U16119 (N_16119,N_10359,N_12086);
nand U16120 (N_16120,N_12083,N_12535);
and U16121 (N_16121,N_13340,N_10473);
and U16122 (N_16122,N_14154,N_14866);
xor U16123 (N_16123,N_10750,N_11621);
nor U16124 (N_16124,N_12292,N_13337);
or U16125 (N_16125,N_11207,N_12005);
nand U16126 (N_16126,N_12249,N_11909);
nor U16127 (N_16127,N_10839,N_11762);
or U16128 (N_16128,N_11333,N_12967);
nor U16129 (N_16129,N_14180,N_13077);
nand U16130 (N_16130,N_10012,N_13954);
nand U16131 (N_16131,N_13689,N_13323);
xnor U16132 (N_16132,N_11101,N_14250);
nor U16133 (N_16133,N_12711,N_11940);
nor U16134 (N_16134,N_13732,N_10458);
nand U16135 (N_16135,N_11485,N_12897);
nor U16136 (N_16136,N_12879,N_14947);
nand U16137 (N_16137,N_14830,N_12825);
and U16138 (N_16138,N_11969,N_10084);
or U16139 (N_16139,N_13605,N_12475);
nor U16140 (N_16140,N_13726,N_10047);
and U16141 (N_16141,N_12127,N_14832);
nor U16142 (N_16142,N_13561,N_12135);
nand U16143 (N_16143,N_12705,N_11370);
or U16144 (N_16144,N_11300,N_12126);
and U16145 (N_16145,N_14797,N_12683);
xor U16146 (N_16146,N_12357,N_11154);
and U16147 (N_16147,N_11312,N_10179);
and U16148 (N_16148,N_10078,N_12230);
nand U16149 (N_16149,N_12446,N_13338);
or U16150 (N_16150,N_12286,N_12512);
nor U16151 (N_16151,N_11068,N_11701);
nor U16152 (N_16152,N_12731,N_14613);
and U16153 (N_16153,N_10484,N_13354);
and U16154 (N_16154,N_10682,N_13942);
nor U16155 (N_16155,N_12791,N_10745);
nand U16156 (N_16156,N_13649,N_13095);
or U16157 (N_16157,N_14859,N_13192);
nor U16158 (N_16158,N_11450,N_14609);
nand U16159 (N_16159,N_10264,N_14688);
nor U16160 (N_16160,N_11147,N_14448);
or U16161 (N_16161,N_13784,N_13329);
and U16162 (N_16162,N_10013,N_12277);
nor U16163 (N_16163,N_12669,N_10696);
and U16164 (N_16164,N_14895,N_13251);
nor U16165 (N_16165,N_12384,N_11284);
or U16166 (N_16166,N_12955,N_12482);
nor U16167 (N_16167,N_10024,N_14475);
or U16168 (N_16168,N_14470,N_10079);
xor U16169 (N_16169,N_12087,N_11730);
and U16170 (N_16170,N_13002,N_10764);
and U16171 (N_16171,N_14099,N_12310);
xor U16172 (N_16172,N_13675,N_13436);
or U16173 (N_16173,N_13404,N_11316);
nor U16174 (N_16174,N_10247,N_10856);
nor U16175 (N_16175,N_13751,N_10389);
nor U16176 (N_16176,N_12204,N_12232);
or U16177 (N_16177,N_10777,N_12868);
nand U16178 (N_16178,N_13073,N_14215);
or U16179 (N_16179,N_10781,N_13554);
xnor U16180 (N_16180,N_12621,N_14721);
and U16181 (N_16181,N_10628,N_12179);
nand U16182 (N_16182,N_11765,N_13668);
xor U16183 (N_16183,N_13034,N_12629);
or U16184 (N_16184,N_13456,N_12039);
and U16185 (N_16185,N_13231,N_10217);
nor U16186 (N_16186,N_12937,N_11186);
nor U16187 (N_16187,N_14145,N_10082);
nor U16188 (N_16188,N_12747,N_14134);
xnor U16189 (N_16189,N_12723,N_11697);
xnor U16190 (N_16190,N_13254,N_10692);
and U16191 (N_16191,N_12114,N_13428);
and U16192 (N_16192,N_11505,N_12486);
nand U16193 (N_16193,N_10345,N_12007);
nand U16194 (N_16194,N_14032,N_12755);
nor U16195 (N_16195,N_11087,N_14234);
nor U16196 (N_16196,N_12108,N_14235);
nand U16197 (N_16197,N_12429,N_13495);
nand U16198 (N_16198,N_13979,N_14677);
or U16199 (N_16199,N_11687,N_11555);
and U16200 (N_16200,N_12652,N_13517);
nand U16201 (N_16201,N_12253,N_11393);
nand U16202 (N_16202,N_10769,N_11681);
nand U16203 (N_16203,N_14933,N_11437);
xnor U16204 (N_16204,N_11674,N_11444);
nand U16205 (N_16205,N_11802,N_10681);
nand U16206 (N_16206,N_13048,N_11038);
nand U16207 (N_16207,N_11122,N_14840);
nand U16208 (N_16208,N_10980,N_14314);
nor U16209 (N_16209,N_13174,N_11844);
and U16210 (N_16210,N_13138,N_12016);
and U16211 (N_16211,N_11752,N_12856);
nand U16212 (N_16212,N_11129,N_14546);
nand U16213 (N_16213,N_14607,N_14295);
xnor U16214 (N_16214,N_12632,N_12581);
nor U16215 (N_16215,N_14757,N_12548);
xor U16216 (N_16216,N_10377,N_14214);
or U16217 (N_16217,N_11646,N_14827);
xor U16218 (N_16218,N_12533,N_14060);
xor U16219 (N_16219,N_11988,N_11615);
and U16220 (N_16220,N_10425,N_13841);
nand U16221 (N_16221,N_12490,N_14588);
or U16222 (N_16222,N_12807,N_14683);
or U16223 (N_16223,N_14759,N_14733);
nor U16224 (N_16224,N_11082,N_13443);
or U16225 (N_16225,N_14191,N_10122);
or U16226 (N_16226,N_11862,N_11744);
nand U16227 (N_16227,N_12019,N_13540);
and U16228 (N_16228,N_10584,N_13145);
xor U16229 (N_16229,N_13640,N_13721);
nor U16230 (N_16230,N_12459,N_13928);
nor U16231 (N_16231,N_12260,N_10101);
and U16232 (N_16232,N_14413,N_12599);
nor U16233 (N_16233,N_11025,N_10044);
nand U16234 (N_16234,N_13886,N_14251);
or U16235 (N_16235,N_12348,N_14000);
nand U16236 (N_16236,N_11928,N_12196);
xnor U16237 (N_16237,N_14914,N_13079);
and U16238 (N_16238,N_11921,N_13082);
nor U16239 (N_16239,N_11011,N_10273);
xor U16240 (N_16240,N_11970,N_14292);
and U16241 (N_16241,N_13399,N_12982);
and U16242 (N_16242,N_11782,N_14058);
nor U16243 (N_16243,N_14969,N_12242);
nand U16244 (N_16244,N_14864,N_13240);
nand U16245 (N_16245,N_11369,N_14728);
nand U16246 (N_16246,N_12735,N_13811);
and U16247 (N_16247,N_10888,N_12046);
nand U16248 (N_16248,N_10655,N_10186);
xor U16249 (N_16249,N_12709,N_13006);
or U16250 (N_16250,N_14712,N_10864);
nand U16251 (N_16251,N_10945,N_13938);
or U16252 (N_16252,N_14514,N_13314);
nor U16253 (N_16253,N_14915,N_12595);
nor U16254 (N_16254,N_14253,N_10440);
and U16255 (N_16255,N_14952,N_14538);
and U16256 (N_16256,N_13832,N_14106);
nor U16257 (N_16257,N_14168,N_12604);
or U16258 (N_16258,N_10444,N_12885);
and U16259 (N_16259,N_11633,N_11576);
and U16260 (N_16260,N_11712,N_10615);
xor U16261 (N_16261,N_11906,N_11457);
nand U16262 (N_16262,N_14916,N_11794);
xnor U16263 (N_16263,N_14172,N_14219);
xnor U16264 (N_16264,N_13056,N_10424);
or U16265 (N_16265,N_10703,N_12543);
nand U16266 (N_16266,N_11852,N_14354);
xnor U16267 (N_16267,N_11482,N_10452);
nor U16268 (N_16268,N_11017,N_12876);
nor U16269 (N_16269,N_11246,N_14338);
or U16270 (N_16270,N_13448,N_12964);
nand U16271 (N_16271,N_10282,N_12183);
nand U16272 (N_16272,N_11173,N_11133);
nand U16273 (N_16273,N_12205,N_11882);
or U16274 (N_16274,N_13759,N_12049);
xor U16275 (N_16275,N_13027,N_12066);
xnor U16276 (N_16276,N_13015,N_13303);
xnor U16277 (N_16277,N_11130,N_13973);
or U16278 (N_16278,N_10209,N_12154);
xnor U16279 (N_16279,N_12379,N_10066);
nand U16280 (N_16280,N_12426,N_11313);
nand U16281 (N_16281,N_10633,N_12316);
xor U16282 (N_16282,N_14939,N_10431);
xor U16283 (N_16283,N_13869,N_14412);
nand U16284 (N_16284,N_13700,N_13101);
nor U16285 (N_16285,N_13844,N_13713);
xnor U16286 (N_16286,N_13076,N_12766);
nor U16287 (N_16287,N_13324,N_13137);
xor U16288 (N_16288,N_12321,N_13020);
and U16289 (N_16289,N_10858,N_14831);
nand U16290 (N_16290,N_12874,N_14347);
and U16291 (N_16291,N_12484,N_11494);
nor U16292 (N_16292,N_11244,N_10978);
nor U16293 (N_16293,N_14132,N_11968);
nand U16294 (N_16294,N_11522,N_13704);
and U16295 (N_16295,N_12737,N_11430);
or U16296 (N_16296,N_10534,N_10459);
nand U16297 (N_16297,N_10291,N_10115);
nor U16298 (N_16298,N_14596,N_12444);
xor U16299 (N_16299,N_11503,N_13298);
and U16300 (N_16300,N_13199,N_10275);
xor U16301 (N_16301,N_10067,N_12148);
or U16302 (N_16302,N_14189,N_10074);
nand U16303 (N_16303,N_13139,N_14802);
nor U16304 (N_16304,N_13305,N_14163);
nand U16305 (N_16305,N_11843,N_10936);
nor U16306 (N_16306,N_14731,N_11546);
nor U16307 (N_16307,N_10958,N_13235);
or U16308 (N_16308,N_14451,N_11532);
and U16309 (N_16309,N_12574,N_11317);
and U16310 (N_16310,N_12363,N_12515);
or U16311 (N_16311,N_10523,N_12746);
or U16312 (N_16312,N_10813,N_11479);
or U16313 (N_16313,N_10507,N_11914);
nor U16314 (N_16314,N_12845,N_12271);
or U16315 (N_16315,N_12265,N_13569);
or U16316 (N_16316,N_12207,N_14752);
or U16317 (N_16317,N_10071,N_12816);
or U16318 (N_16318,N_11793,N_10252);
xor U16319 (N_16319,N_13943,N_13720);
nor U16320 (N_16320,N_10123,N_13672);
nor U16321 (N_16321,N_10524,N_12442);
nor U16322 (N_16322,N_12640,N_10785);
nor U16323 (N_16323,N_13874,N_13102);
or U16324 (N_16324,N_13177,N_10800);
nand U16325 (N_16325,N_11484,N_12950);
or U16326 (N_16326,N_12290,N_11915);
nand U16327 (N_16327,N_10127,N_14930);
nor U16328 (N_16328,N_13085,N_11763);
and U16329 (N_16329,N_10624,N_11719);
or U16330 (N_16330,N_10583,N_12368);
nand U16331 (N_16331,N_11401,N_14707);
or U16332 (N_16332,N_14934,N_11362);
xor U16333 (N_16333,N_13902,N_12760);
nor U16334 (N_16334,N_10737,N_12303);
nand U16335 (N_16335,N_10528,N_13424);
nand U16336 (N_16336,N_13710,N_14612);
nor U16337 (N_16337,N_12834,N_10814);
nor U16338 (N_16338,N_13164,N_12281);
nand U16339 (N_16339,N_10296,N_12119);
xor U16340 (N_16340,N_12464,N_13593);
or U16341 (N_16341,N_12323,N_13556);
nand U16342 (N_16342,N_12338,N_14805);
nand U16343 (N_16343,N_13311,N_11616);
nand U16344 (N_16344,N_14276,N_12924);
nor U16345 (N_16345,N_13022,N_12762);
nor U16346 (N_16346,N_11742,N_11838);
and U16347 (N_16347,N_12620,N_10333);
nor U16348 (N_16348,N_10738,N_13074);
or U16349 (N_16349,N_13178,N_10175);
xnor U16350 (N_16350,N_10023,N_10322);
or U16351 (N_16351,N_10011,N_13949);
and U16352 (N_16352,N_13559,N_13080);
nand U16353 (N_16353,N_12142,N_12328);
nor U16354 (N_16354,N_14331,N_12076);
nor U16355 (N_16355,N_10107,N_11971);
xnor U16356 (N_16356,N_14668,N_10267);
xnor U16357 (N_16357,N_11480,N_14753);
or U16358 (N_16358,N_11396,N_11999);
nand U16359 (N_16359,N_11955,N_10938);
nand U16360 (N_16360,N_14041,N_11418);
nor U16361 (N_16361,N_12319,N_12090);
or U16362 (N_16362,N_12570,N_12014);
nand U16363 (N_16363,N_11625,N_11424);
xor U16364 (N_16364,N_11386,N_11865);
nand U16365 (N_16365,N_10552,N_14433);
and U16366 (N_16366,N_14878,N_13828);
xor U16367 (N_16367,N_12030,N_13017);
xor U16368 (N_16368,N_14183,N_11558);
nor U16369 (N_16369,N_13224,N_11657);
and U16370 (N_16370,N_10303,N_11736);
and U16371 (N_16371,N_10419,N_10650);
and U16372 (N_16372,N_10662,N_10105);
xnor U16373 (N_16373,N_10591,N_14160);
or U16374 (N_16374,N_13366,N_13287);
nor U16375 (N_16375,N_13106,N_12437);
nor U16376 (N_16376,N_14513,N_11276);
or U16377 (N_16377,N_12901,N_12047);
nor U16378 (N_16378,N_12953,N_10520);
or U16379 (N_16379,N_12017,N_10249);
or U16380 (N_16380,N_10334,N_14357);
xnor U16381 (N_16381,N_10736,N_10684);
nand U16382 (N_16382,N_11645,N_10879);
nor U16383 (N_16383,N_11805,N_13534);
xnor U16384 (N_16384,N_11240,N_12984);
xor U16385 (N_16385,N_14899,N_14744);
or U16386 (N_16386,N_12407,N_14539);
xor U16387 (N_16387,N_11511,N_14300);
and U16388 (N_16388,N_10315,N_12761);
or U16389 (N_16389,N_13860,N_10482);
nand U16390 (N_16390,N_14435,N_10659);
nor U16391 (N_16391,N_11754,N_11704);
or U16392 (N_16392,N_13639,N_13083);
xor U16393 (N_16393,N_14006,N_14162);
nor U16394 (N_16394,N_10999,N_10974);
nor U16395 (N_16395,N_13645,N_11585);
or U16396 (N_16396,N_11942,N_14792);
and U16397 (N_16397,N_11892,N_11032);
or U16398 (N_16398,N_10404,N_11073);
or U16399 (N_16399,N_13826,N_11694);
nand U16400 (N_16400,N_12212,N_10085);
nor U16401 (N_16401,N_12740,N_12152);
nor U16402 (N_16402,N_12675,N_10069);
or U16403 (N_16403,N_14387,N_10959);
nand U16404 (N_16404,N_11927,N_11164);
xnor U16405 (N_16405,N_12096,N_11007);
nor U16406 (N_16406,N_10329,N_10220);
xor U16407 (N_16407,N_14902,N_10009);
xor U16408 (N_16408,N_10794,N_10065);
and U16409 (N_16409,N_11289,N_10894);
and U16410 (N_16410,N_12029,N_11400);
nor U16411 (N_16411,N_13133,N_11137);
or U16412 (N_16412,N_10392,N_14686);
nand U16413 (N_16413,N_14176,N_13542);
xor U16414 (N_16414,N_10356,N_14227);
nor U16415 (N_16415,N_11672,N_11349);
and U16416 (N_16416,N_10413,N_11510);
or U16417 (N_16417,N_13577,N_14021);
and U16418 (N_16418,N_13567,N_11187);
nor U16419 (N_16419,N_13947,N_13616);
nand U16420 (N_16420,N_12501,N_12833);
or U16421 (N_16421,N_12136,N_11836);
xor U16422 (N_16422,N_13140,N_14537);
nand U16423 (N_16423,N_12883,N_13580);
or U16424 (N_16424,N_13653,N_13853);
nand U16425 (N_16425,N_10237,N_14669);
and U16426 (N_16426,N_13646,N_14340);
or U16427 (N_16427,N_12130,N_14689);
nand U16428 (N_16428,N_10049,N_10349);
and U16429 (N_16429,N_11948,N_10665);
xnor U16430 (N_16430,N_12651,N_10852);
nor U16431 (N_16431,N_11559,N_13274);
nor U16432 (N_16432,N_11206,N_10238);
or U16433 (N_16433,N_14664,N_12704);
nor U16434 (N_16434,N_11521,N_12653);
nand U16435 (N_16435,N_12137,N_13463);
or U16436 (N_16436,N_14716,N_14699);
nand U16437 (N_16437,N_14420,N_11468);
xnor U16438 (N_16438,N_13005,N_11895);
or U16439 (N_16439,N_11063,N_10707);
and U16440 (N_16440,N_12799,N_11095);
and U16441 (N_16441,N_11308,N_14029);
nor U16442 (N_16442,N_13769,N_11176);
and U16443 (N_16443,N_14789,N_14027);
and U16444 (N_16444,N_11315,N_10893);
xor U16445 (N_16445,N_11643,N_11416);
nor U16446 (N_16446,N_14031,N_12785);
or U16447 (N_16447,N_13040,N_11202);
nand U16448 (N_16448,N_12900,N_10378);
xor U16449 (N_16449,N_11123,N_10427);
and U16450 (N_16450,N_11097,N_13546);
or U16451 (N_16451,N_13935,N_10097);
or U16452 (N_16452,N_10643,N_11780);
nand U16453 (N_16453,N_14198,N_12481);
xnor U16454 (N_16454,N_13526,N_11668);
nand U16455 (N_16455,N_12500,N_14313);
nor U16456 (N_16456,N_11379,N_10772);
or U16457 (N_16457,N_10634,N_14225);
nor U16458 (N_16458,N_12738,N_14076);
nor U16459 (N_16459,N_13273,N_12594);
nand U16460 (N_16460,N_12858,N_14659);
nor U16461 (N_16461,N_12070,N_11801);
nand U16462 (N_16462,N_11465,N_11699);
nand U16463 (N_16463,N_13818,N_11429);
xor U16464 (N_16464,N_14447,N_14159);
nor U16465 (N_16465,N_11849,N_12765);
nand U16466 (N_16466,N_11979,N_13142);
or U16467 (N_16467,N_13278,N_13815);
nor U16468 (N_16468,N_14077,N_14355);
xor U16469 (N_16469,N_10226,N_12391);
or U16470 (N_16470,N_14174,N_14540);
nand U16471 (N_16471,N_12914,N_12830);
nand U16472 (N_16472,N_11925,N_12626);
xnor U16473 (N_16473,N_11215,N_11614);
or U16474 (N_16474,N_14713,N_14089);
nor U16475 (N_16475,N_14737,N_10593);
and U16476 (N_16476,N_12274,N_14070);
and U16477 (N_16477,N_14502,N_12156);
xor U16478 (N_16478,N_14184,N_11833);
and U16479 (N_16479,N_14319,N_10332);
xor U16480 (N_16480,N_13929,N_14766);
nand U16481 (N_16481,N_13492,N_13105);
nand U16482 (N_16482,N_14111,N_13308);
nor U16483 (N_16483,N_10533,N_12177);
and U16484 (N_16484,N_12531,N_11519);
and U16485 (N_16485,N_10637,N_12607);
nand U16486 (N_16486,N_13090,N_14398);
or U16487 (N_16487,N_12934,N_14725);
nor U16488 (N_16488,N_14972,N_13412);
and U16489 (N_16489,N_12153,N_11539);
or U16490 (N_16490,N_13012,N_13532);
nand U16491 (N_16491,N_14152,N_12006);
nor U16492 (N_16492,N_14821,N_10292);
or U16493 (N_16493,N_10854,N_13334);
nor U16494 (N_16494,N_12034,N_14873);
and U16495 (N_16495,N_12170,N_14693);
nand U16496 (N_16496,N_11980,N_14332);
nor U16497 (N_16497,N_14010,N_13207);
nor U16498 (N_16498,N_12736,N_11845);
nor U16499 (N_16499,N_11409,N_14724);
nor U16500 (N_16500,N_13156,N_14431);
and U16501 (N_16501,N_14202,N_11675);
and U16502 (N_16502,N_14525,N_12244);
xor U16503 (N_16503,N_10138,N_12836);
nor U16504 (N_16504,N_14484,N_11151);
or U16505 (N_16505,N_12793,N_11449);
nor U16506 (N_16506,N_11039,N_14905);
or U16507 (N_16507,N_12602,N_13708);
or U16508 (N_16508,N_11983,N_10607);
nor U16509 (N_16509,N_14418,N_12180);
and U16510 (N_16510,N_13016,N_10502);
and U16511 (N_16511,N_12828,N_11617);
xnor U16512 (N_16512,N_10521,N_10986);
or U16513 (N_16513,N_14602,N_12739);
and U16514 (N_16514,N_11066,N_10072);
xor U16515 (N_16515,N_13836,N_12546);
nand U16516 (N_16516,N_14093,N_12668);
or U16517 (N_16517,N_14877,N_14860);
or U16518 (N_16518,N_14663,N_11259);
xor U16519 (N_16519,N_11728,N_14464);
nand U16520 (N_16520,N_11364,N_11059);
xor U16521 (N_16521,N_13485,N_13472);
xnor U16522 (N_16522,N_11608,N_13859);
and U16523 (N_16523,N_11580,N_11175);
or U16524 (N_16524,N_11751,N_12117);
and U16525 (N_16525,N_13627,N_10338);
or U16526 (N_16526,N_14116,N_11547);
xor U16527 (N_16527,N_11436,N_12473);
nand U16528 (N_16528,N_10580,N_13834);
nor U16529 (N_16529,N_14304,N_13291);
nand U16530 (N_16530,N_11711,N_10567);
and U16531 (N_16531,N_10286,N_12628);
nand U16532 (N_16532,N_14880,N_12268);
or U16533 (N_16533,N_12131,N_13586);
nand U16534 (N_16534,N_13383,N_14573);
nor U16535 (N_16535,N_10007,N_10153);
xor U16536 (N_16536,N_12656,N_12887);
xnor U16537 (N_16537,N_14294,N_12169);
nand U16538 (N_16538,N_10169,N_10164);
and U16539 (N_16539,N_14871,N_14901);
xor U16540 (N_16540,N_12923,N_13930);
or U16541 (N_16541,N_10027,N_12028);
nor U16542 (N_16542,N_13123,N_12691);
and U16543 (N_16543,N_12862,N_13674);
or U16544 (N_16544,N_14709,N_14626);
nor U16545 (N_16545,N_13964,N_12748);
xor U16546 (N_16546,N_11119,N_10418);
and U16547 (N_16547,N_11114,N_14698);
xnor U16548 (N_16548,N_12309,N_14976);
nor U16549 (N_16549,N_14591,N_11254);
and U16550 (N_16550,N_14768,N_13892);
nor U16551 (N_16551,N_11552,N_11451);
xnor U16552 (N_16552,N_13348,N_14359);
nor U16553 (N_16553,N_14926,N_13125);
nand U16554 (N_16554,N_12377,N_12495);
and U16555 (N_16555,N_11958,N_11916);
and U16556 (N_16556,N_13230,N_10494);
or U16557 (N_16557,N_11934,N_14405);
nand U16558 (N_16558,N_14633,N_11094);
nand U16559 (N_16559,N_14391,N_10540);
and U16560 (N_16560,N_10470,N_12247);
and U16561 (N_16561,N_13282,N_11676);
and U16562 (N_16562,N_12032,N_11854);
xor U16563 (N_16563,N_12763,N_12094);
nor U16564 (N_16564,N_14943,N_13325);
nor U16565 (N_16565,N_13346,N_13442);
or U16566 (N_16566,N_14654,N_11566);
xnor U16567 (N_16567,N_14703,N_12865);
xor U16568 (N_16568,N_13289,N_11091);
nand U16569 (N_16569,N_12534,N_11811);
or U16570 (N_16570,N_11658,N_12528);
nor U16571 (N_16571,N_14944,N_10515);
nand U16572 (N_16572,N_14362,N_13599);
or U16573 (N_16573,N_10625,N_14867);
nor U16574 (N_16574,N_11257,N_14209);
or U16575 (N_16575,N_11653,N_12224);
or U16576 (N_16576,N_13126,N_14290);
nor U16577 (N_16577,N_11192,N_10146);
and U16578 (N_16578,N_13911,N_13196);
nor U16579 (N_16579,N_14170,N_13198);
or U16580 (N_16580,N_13673,N_12819);
or U16581 (N_16581,N_10620,N_10372);
xnor U16582 (N_16582,N_14117,N_10952);
xor U16583 (N_16583,N_14541,N_14317);
or U16584 (N_16584,N_13576,N_14740);
nand U16585 (N_16585,N_14158,N_12797);
and U16586 (N_16586,N_13064,N_12558);
nor U16587 (N_16587,N_12718,N_11542);
nor U16588 (N_16588,N_10678,N_13491);
and U16589 (N_16589,N_11329,N_12167);
and U16590 (N_16590,N_14204,N_11696);
xnor U16591 (N_16591,N_12027,N_13155);
xnor U16592 (N_16592,N_11957,N_13660);
nand U16593 (N_16593,N_10940,N_11132);
nor U16594 (N_16594,N_14751,N_11344);
and U16595 (N_16595,N_14384,N_10352);
xor U16596 (N_16596,N_12549,N_11717);
nor U16597 (N_16597,N_10462,N_12266);
and U16598 (N_16598,N_10386,N_10346);
xnor U16599 (N_16599,N_14080,N_11266);
xor U16600 (N_16600,N_10768,N_10733);
nor U16601 (N_16601,N_10691,N_11611);
xor U16602 (N_16602,N_12660,N_13369);
nor U16603 (N_16603,N_12362,N_13362);
or U16604 (N_16604,N_10964,N_12920);
and U16605 (N_16605,N_13624,N_10182);
nor U16606 (N_16606,N_14656,N_10962);
xor U16607 (N_16607,N_10202,N_13855);
or U16608 (N_16608,N_14735,N_10617);
and U16609 (N_16609,N_11883,N_12702);
or U16610 (N_16610,N_12757,N_13864);
xor U16611 (N_16611,N_10490,N_12257);
nor U16612 (N_16612,N_11872,N_11071);
and U16613 (N_16613,N_13221,N_12518);
and U16614 (N_16614,N_13899,N_11404);
xnor U16615 (N_16615,N_14083,N_13692);
nor U16616 (N_16616,N_12706,N_12732);
or U16617 (N_16617,N_10886,N_14476);
nor U16618 (N_16618,N_12855,N_12374);
and U16619 (N_16619,N_13779,N_12040);
or U16620 (N_16620,N_12092,N_10210);
or U16621 (N_16621,N_12888,N_10438);
and U16622 (N_16622,N_10229,N_11411);
xnor U16623 (N_16623,N_13473,N_13530);
and U16624 (N_16624,N_14971,N_13920);
nor U16625 (N_16625,N_14822,N_12491);
nand U16626 (N_16626,N_14516,N_10199);
or U16627 (N_16627,N_10363,N_11003);
nand U16628 (N_16628,N_13931,N_11579);
xor U16629 (N_16629,N_12416,N_10509);
and U16630 (N_16630,N_12985,N_10096);
xnor U16631 (N_16631,N_13021,N_11723);
xor U16632 (N_16632,N_10486,N_11618);
nand U16633 (N_16633,N_10967,N_13482);
nor U16634 (N_16634,N_12372,N_11683);
or U16635 (N_16635,N_10712,N_12952);
xor U16636 (N_16636,N_14380,N_14966);
xor U16637 (N_16637,N_12930,N_11258);
nor U16638 (N_16638,N_12413,N_11825);
or U16639 (N_16639,N_10054,N_14542);
or U16640 (N_16640,N_14474,N_12382);
xor U16641 (N_16641,N_10442,N_12563);
nor U16642 (N_16642,N_13024,N_13070);
nor U16643 (N_16643,N_13833,N_11530);
xor U16644 (N_16644,N_10757,N_10536);
nand U16645 (N_16645,N_13173,N_11549);
or U16646 (N_16646,N_13724,N_11372);
nor U16647 (N_16647,N_13392,N_14374);
and U16648 (N_16648,N_14924,N_13991);
xnor U16649 (N_16649,N_10029,N_11507);
or U16650 (N_16650,N_14469,N_14486);
nor U16651 (N_16651,N_13824,N_10033);
nor U16652 (N_16652,N_11641,N_13508);
and U16653 (N_16653,N_12498,N_11390);
xor U16654 (N_16654,N_11044,N_12162);
and U16655 (N_16655,N_11477,N_11249);
and U16656 (N_16656,N_14552,N_13363);
xnor U16657 (N_16657,N_12848,N_13987);
and U16658 (N_16658,N_12569,N_13615);
or U16659 (N_16659,N_10761,N_13505);
nand U16660 (N_16660,N_12875,N_11288);
xor U16661 (N_16661,N_13970,N_12898);
nand U16662 (N_16662,N_10568,N_14386);
nor U16663 (N_16663,N_11870,N_12756);
and U16664 (N_16664,N_14296,N_11864);
xnor U16665 (N_16665,N_12074,N_10782);
nor U16666 (N_16666,N_11899,N_12527);
and U16667 (N_16667,N_13609,N_13018);
nand U16668 (N_16668,N_11384,N_13342);
or U16669 (N_16669,N_11936,N_10225);
and U16670 (N_16670,N_13188,N_13390);
nand U16671 (N_16671,N_10658,N_12596);
nor U16672 (N_16672,N_12864,N_13257);
nor U16673 (N_16673,N_14635,N_13261);
and U16674 (N_16674,N_11145,N_11079);
xnor U16675 (N_16675,N_14395,N_13285);
nor U16676 (N_16676,N_12936,N_14795);
nand U16677 (N_16677,N_10758,N_13514);
and U16678 (N_16678,N_14133,N_11225);
and U16679 (N_16679,N_10116,N_14381);
xor U16680 (N_16680,N_10916,N_14855);
nand U16681 (N_16681,N_14888,N_10398);
and U16682 (N_16682,N_14790,N_11296);
xor U16683 (N_16683,N_12050,N_11851);
and U16684 (N_16684,N_11088,N_10271);
or U16685 (N_16685,N_10471,N_13072);
nand U16686 (N_16686,N_11069,N_13589);
or U16687 (N_16687,N_10443,N_10218);
xnor U16688 (N_16688,N_12216,N_14781);
nor U16689 (N_16689,N_10152,N_10530);
xor U16690 (N_16690,N_13912,N_10294);
or U16691 (N_16691,N_12110,N_14267);
nor U16692 (N_16692,N_13703,N_12151);
nor U16693 (N_16693,N_13997,N_11336);
and U16694 (N_16694,N_10835,N_11368);
and U16695 (N_16695,N_14586,N_14262);
xor U16696 (N_16696,N_14959,N_14964);
and U16697 (N_16697,N_14088,N_13873);
or U16698 (N_16698,N_10318,N_11357);
or U16699 (N_16699,N_14991,N_11691);
or U16700 (N_16700,N_11774,N_14394);
and U16701 (N_16701,N_12703,N_12998);
or U16702 (N_16702,N_10205,N_11499);
or U16703 (N_16703,N_14520,N_12104);
or U16704 (N_16704,N_11193,N_12576);
nor U16705 (N_16705,N_12189,N_11725);
xor U16706 (N_16706,N_13527,N_12356);
and U16707 (N_16707,N_14845,N_13765);
nand U16708 (N_16708,N_11387,N_13111);
or U16709 (N_16709,N_11733,N_10606);
or U16710 (N_16710,N_11064,N_11253);
and U16711 (N_16711,N_12441,N_13771);
or U16712 (N_16712,N_10343,N_14282);
and U16713 (N_16713,N_10260,N_10582);
nand U16714 (N_16714,N_14980,N_11204);
nand U16715 (N_16715,N_14628,N_14798);
and U16716 (N_16716,N_12361,N_14166);
and U16717 (N_16717,N_10944,N_11809);
and U16718 (N_16718,N_12105,N_11004);
nand U16719 (N_16719,N_10445,N_12798);
or U16720 (N_16720,N_12010,N_14807);
xnor U16721 (N_16721,N_10466,N_11677);
and U16722 (N_16722,N_10676,N_12610);
or U16723 (N_16723,N_10934,N_12941);
nor U16724 (N_16724,N_11350,N_10388);
nor U16725 (N_16725,N_11113,N_10592);
nand U16726 (N_16726,N_12404,N_14935);
and U16727 (N_16727,N_10293,N_12238);
xnor U16728 (N_16728,N_11866,N_13766);
and U16729 (N_16729,N_10647,N_10173);
and U16730 (N_16730,N_13300,N_11076);
nor U16731 (N_16731,N_14515,N_12688);
xnor U16732 (N_16732,N_11602,N_11524);
and U16733 (N_16733,N_12419,N_12743);
and U16734 (N_16734,N_13975,N_12929);
and U16735 (N_16735,N_10603,N_14061);
and U16736 (N_16736,N_13025,N_12506);
and U16737 (N_16737,N_14241,N_14852);
or U16738 (N_16738,N_11014,N_10348);
and U16739 (N_16739,N_10095,N_13635);
nor U16740 (N_16740,N_11798,N_11118);
or U16741 (N_16741,N_12579,N_11250);
or U16742 (N_16742,N_12327,N_11172);
nand U16743 (N_16743,N_14249,N_11458);
and U16744 (N_16744,N_11998,N_10850);
nand U16745 (N_16745,N_12577,N_12976);
or U16746 (N_16746,N_14181,N_11893);
or U16747 (N_16747,N_13521,N_10862);
nand U16748 (N_16748,N_12100,N_13457);
nor U16749 (N_16749,N_11514,N_11405);
nor U16750 (N_16750,N_11022,N_14148);
xnor U16751 (N_16751,N_14621,N_10355);
or U16752 (N_16752,N_13234,N_11504);
xnor U16753 (N_16753,N_10111,N_10954);
or U16754 (N_16754,N_10597,N_12568);
nand U16755 (N_16755,N_13965,N_11290);
and U16756 (N_16756,N_11718,N_10908);
nand U16757 (N_16757,N_14528,N_14238);
or U16758 (N_16758,N_10259,N_11260);
nor U16759 (N_16759,N_11788,N_11822);
and U16760 (N_16760,N_10805,N_10627);
nand U16761 (N_16761,N_14377,N_12983);
or U16762 (N_16762,N_12804,N_14363);
nand U16763 (N_16763,N_12815,N_12661);
nand U16764 (N_16764,N_10455,N_11231);
nand U16765 (N_16765,N_10219,N_10572);
nor U16766 (N_16766,N_11408,N_10014);
nand U16767 (N_16767,N_10594,N_13648);
nor U16768 (N_16768,N_10396,N_10787);
or U16769 (N_16769,N_13433,N_11931);
nor U16770 (N_16770,N_11098,N_12663);
nand U16771 (N_16771,N_10309,N_14765);
xnor U16772 (N_16772,N_13134,N_13845);
and U16773 (N_16773,N_11382,N_11106);
nand U16774 (N_16774,N_11374,N_12195);
nor U16775 (N_16775,N_14772,N_12219);
nor U16776 (N_16776,N_10151,N_11034);
and U16777 (N_16777,N_13226,N_10506);
or U16778 (N_16778,N_14342,N_11412);
nand U16779 (N_16779,N_13248,N_10394);
xnor U16780 (N_16780,N_10749,N_14024);
xor U16781 (N_16781,N_13944,N_12436);
xor U16782 (N_16782,N_11115,N_14466);
nor U16783 (N_16783,N_14565,N_13866);
nor U16784 (N_16784,N_13679,N_12115);
nand U16785 (N_16785,N_12004,N_11283);
nand U16786 (N_16786,N_11706,N_14550);
or U16787 (N_16787,N_12336,N_11930);
or U16788 (N_16788,N_13476,N_11753);
nand U16789 (N_16789,N_12992,N_12393);
nor U16790 (N_16790,N_14488,N_10660);
and U16791 (N_16791,N_11601,N_13130);
nor U16792 (N_16792,N_14231,N_11654);
nand U16793 (N_16793,N_12788,N_14071);
or U16794 (N_16794,N_12603,N_12678);
nand U16795 (N_16795,N_12288,N_14095);
or U16796 (N_16796,N_10604,N_14770);
nor U16797 (N_16797,N_11140,N_12608);
and U16798 (N_16798,N_14366,N_14732);
xor U16799 (N_16799,N_12776,N_10243);
or U16800 (N_16800,N_13393,N_14736);
or U16801 (N_16801,N_11170,N_13011);
or U16802 (N_16802,N_10641,N_11686);
xnor U16803 (N_16803,N_13695,N_12894);
nor U16804 (N_16804,N_13917,N_14863);
or U16805 (N_16805,N_13464,N_12977);
nand U16806 (N_16806,N_13318,N_10474);
nor U16807 (N_16807,N_12366,N_12139);
nor U16808 (N_16808,N_13884,N_12938);
and U16809 (N_16809,N_11462,N_10062);
nor U16810 (N_16810,N_10754,N_11850);
or U16811 (N_16811,N_11685,N_11417);
or U16812 (N_16812,N_14443,N_13978);
or U16813 (N_16813,N_11743,N_10149);
xnor U16814 (N_16814,N_13574,N_10710);
nand U16815 (N_16815,N_13269,N_14210);
nor U16816 (N_16816,N_11735,N_11639);
xnor U16817 (N_16817,N_13670,N_13555);
nor U16818 (N_16818,N_13749,N_12206);
nand U16819 (N_16819,N_13001,N_11294);
nor U16820 (N_16820,N_13481,N_11321);
nor U16821 (N_16821,N_11898,N_14096);
or U16822 (N_16822,N_13253,N_14717);
xor U16823 (N_16823,N_13055,N_10585);
xor U16824 (N_16824,N_11353,N_14979);
nand U16825 (N_16825,N_13252,N_13225);
or U16826 (N_16826,N_10204,N_10417);
nor U16827 (N_16827,N_14419,N_14858);
nand U16828 (N_16828,N_13922,N_10901);
xor U16829 (N_16829,N_13760,N_10156);
xor U16830 (N_16830,N_11926,N_12063);
xnor U16831 (N_16831,N_11599,N_11600);
xnor U16832 (N_16832,N_13729,N_14906);
nand U16833 (N_16833,N_12742,N_10797);
xnor U16834 (N_16834,N_11410,N_14002);
nor U16835 (N_16835,N_12194,N_12649);
nor U16836 (N_16836,N_12893,N_13622);
nor U16837 (N_16837,N_11710,N_12213);
nand U16838 (N_16838,N_12354,N_14651);
xnor U16839 (N_16839,N_12745,N_11527);
and U16840 (N_16840,N_14890,N_13940);
xnor U16841 (N_16841,N_12790,N_10272);
nand U16842 (N_16842,N_13459,N_14582);
nand U16843 (N_16843,N_14734,N_13186);
or U16844 (N_16844,N_14809,N_11592);
nand U16845 (N_16845,N_14942,N_13500);
and U16846 (N_16846,N_13425,N_13602);
or U16847 (N_16847,N_10556,N_11876);
and U16848 (N_16848,N_10235,N_13203);
or U16849 (N_16849,N_11030,N_12609);
or U16850 (N_16850,N_14263,N_14098);
and U16851 (N_16851,N_10171,N_10668);
xnor U16852 (N_16852,N_11640,N_14325);
nand U16853 (N_16853,N_10873,N_13881);
xor U16854 (N_16854,N_10426,N_10491);
and U16855 (N_16855,N_12270,N_13787);
and U16856 (N_16856,N_12431,N_13614);
or U16857 (N_16857,N_14373,N_10788);
nand U16858 (N_16858,N_10605,N_11285);
or U16859 (N_16859,N_11413,N_14023);
xnor U16860 (N_16860,N_10826,N_13430);
and U16861 (N_16861,N_11655,N_11726);
xor U16862 (N_16862,N_11965,N_11604);
or U16863 (N_16863,N_14478,N_11178);
xor U16864 (N_16864,N_12060,N_11200);
and U16865 (N_16865,N_13742,N_10871);
and U16866 (N_16866,N_13166,N_12317);
xnor U16867 (N_16867,N_11348,N_14051);
and U16868 (N_16868,N_14379,N_14589);
xor U16869 (N_16869,N_11495,N_12478);
nand U16870 (N_16870,N_12231,N_10715);
nand U16871 (N_16871,N_11219,N_14747);
and U16872 (N_16872,N_12023,N_12768);
nand U16873 (N_16873,N_12280,N_13548);
nor U16874 (N_16874,N_12846,N_13959);
xor U16875 (N_16875,N_12064,N_12571);
or U16876 (N_16876,N_11109,N_12679);
nor U16877 (N_16877,N_13118,N_13575);
xnor U16878 (N_16878,N_11659,N_13923);
nand U16879 (N_16879,N_11531,N_13333);
and U16880 (N_16880,N_10365,N_10991);
xnor U16881 (N_16881,N_12447,N_10553);
nand U16882 (N_16882,N_12695,N_13319);
or U16883 (N_16883,N_10973,N_13071);
nor U16884 (N_16884,N_11060,N_10242);
nand U16885 (N_16885,N_14936,N_12236);
nand U16886 (N_16886,N_12770,N_10073);
xor U16887 (N_16887,N_13994,N_10728);
or U16888 (N_16888,N_10575,N_11820);
or U16889 (N_16889,N_12175,N_13628);
or U16890 (N_16890,N_11242,N_13647);
nor U16891 (N_16891,N_14353,N_13331);
and U16892 (N_16892,N_13693,N_11220);
nor U16893 (N_16893,N_13623,N_13415);
nand U16894 (N_16894,N_13966,N_11989);
nor U16895 (N_16895,N_13223,N_11863);
nand U16896 (N_16896,N_14938,N_12395);
nor U16897 (N_16897,N_10751,N_13228);
and U16898 (N_16898,N_10304,N_12388);
and U16899 (N_16899,N_11065,N_14415);
and U16900 (N_16900,N_10362,N_13891);
and U16901 (N_16901,N_14320,N_13568);
xnor U16902 (N_16902,N_10198,N_10314);
xor U16903 (N_16903,N_10711,N_10195);
nor U16904 (N_16904,N_13336,N_10057);
xor U16905 (N_16905,N_13377,N_10211);
nor U16906 (N_16906,N_12873,N_10058);
nor U16907 (N_16907,N_13216,N_14893);
xor U16908 (N_16908,N_14791,N_13961);
xor U16909 (N_16909,N_11734,N_12009);
or U16910 (N_16910,N_10989,N_12058);
or U16911 (N_16911,N_14479,N_13595);
and U16912 (N_16912,N_11650,N_13045);
nand U16913 (N_16913,N_14352,N_11679);
nand U16914 (N_16914,N_11959,N_10775);
and U16915 (N_16915,N_10233,N_11049);
nand U16916 (N_16916,N_10796,N_10616);
xor U16917 (N_16917,N_14870,N_12928);
or U16918 (N_16918,N_12647,N_12606);
nand U16919 (N_16919,N_13550,N_10048);
and U16920 (N_16920,N_14498,N_14019);
and U16921 (N_16921,N_11966,N_12400);
or U16922 (N_16922,N_10387,N_12623);
xor U16923 (N_16923,N_12870,N_13776);
nand U16924 (N_16924,N_11056,N_12344);
or U16925 (N_16925,N_14345,N_13764);
or U16926 (N_16926,N_12708,N_10150);
nor U16927 (N_16927,N_10977,N_11759);
nand U16928 (N_16928,N_14543,N_11636);
and U16929 (N_16929,N_14968,N_12808);
nor U16930 (N_16930,N_10141,N_11781);
xnor U16931 (N_16931,N_13132,N_11125);
nor U16932 (N_16932,N_14358,N_14865);
or U16933 (N_16933,N_14894,N_11061);
or U16934 (N_16934,N_11652,N_12553);
xnor U16935 (N_16935,N_13116,N_10342);
or U16936 (N_16936,N_12380,N_10561);
nor U16937 (N_16937,N_12693,N_12237);
nand U16938 (N_16938,N_14206,N_14563);
nor U16939 (N_16939,N_11775,N_13819);
xnor U16940 (N_16940,N_11768,N_10998);
and U16941 (N_16941,N_14045,N_10793);
or U16942 (N_16942,N_10099,N_10714);
and U16943 (N_16943,N_12995,N_14388);
and U16944 (N_16944,N_10406,N_11481);
nor U16945 (N_16945,N_14336,N_12406);
nor U16946 (N_16946,N_12378,N_14506);
nor U16947 (N_16947,N_14554,N_13962);
xnor U16948 (N_16948,N_12922,N_10080);
nor U16949 (N_16949,N_12448,N_10876);
or U16950 (N_16950,N_13209,N_12672);
xnor U16951 (N_16951,N_14826,N_10514);
nor U16952 (N_16952,N_10569,N_10463);
nand U16953 (N_16953,N_11280,N_10526);
or U16954 (N_16954,N_12225,N_14578);
or U16955 (N_16955,N_11673,N_13053);
nor U16956 (N_16956,N_10162,N_13659);
nand U16957 (N_16957,N_12544,N_11448);
nor U16958 (N_16958,N_10121,N_12635);
nor U16959 (N_16959,N_12161,N_10883);
and U16960 (N_16960,N_13972,N_13993);
nand U16961 (N_16961,N_12392,N_10002);
nor U16962 (N_16962,N_12073,N_11533);
nor U16963 (N_16963,N_11880,N_13153);
or U16964 (N_16964,N_14190,N_14022);
or U16965 (N_16965,N_10695,N_13781);
or U16966 (N_16966,N_14066,N_14306);
and U16967 (N_16967,N_11582,N_13332);
nor U16968 (N_16968,N_14593,N_13701);
xor U16969 (N_16969,N_14020,N_13038);
and U16970 (N_16970,N_11110,N_10921);
and U16971 (N_16971,N_12410,N_10489);
or U16972 (N_16972,N_12398,N_12880);
nand U16973 (N_16973,N_13752,N_11023);
nand U16974 (N_16974,N_13791,N_11900);
xor U16975 (N_16975,N_14754,N_14786);
and U16976 (N_16976,N_14491,N_10847);
or U16977 (N_16977,N_10519,N_11108);
or U16978 (N_16978,N_14417,N_14592);
or U16979 (N_16979,N_12516,N_13740);
nor U16980 (N_16980,N_13835,N_12483);
xnor U16981 (N_16981,N_13583,N_11126);
nand U16982 (N_16982,N_13862,N_10720);
xor U16983 (N_16983,N_13023,N_13047);
xnor U16984 (N_16984,N_11996,N_10810);
xor U16985 (N_16985,N_14048,N_10288);
nand U16986 (N_16986,N_10077,N_14107);
nand U16987 (N_16987,N_11251,N_12192);
nor U16988 (N_16988,N_10476,N_10385);
and U16989 (N_16989,N_14307,N_12684);
and U16990 (N_16990,N_13731,N_13794);
xnor U16991 (N_16991,N_14213,N_13803);
xnor U16992 (N_16992,N_12687,N_14208);
nor U16993 (N_16993,N_10982,N_11452);
or U16994 (N_16994,N_11755,N_13883);
xor U16995 (N_16995,N_12164,N_13690);
nand U16996 (N_16996,N_12359,N_13950);
xnor U16997 (N_16997,N_14480,N_11777);
or U16998 (N_16998,N_10015,N_13255);
nor U16999 (N_16999,N_13552,N_14919);
nand U17000 (N_17000,N_13405,N_13279);
or U17001 (N_17001,N_10565,N_10640);
nor U17002 (N_17002,N_12203,N_11311);
or U17003 (N_17003,N_10860,N_13220);
xnor U17004 (N_17004,N_11994,N_14833);
nor U17005 (N_17005,N_11149,N_12750);
xor U17006 (N_17006,N_13813,N_11335);
nor U17007 (N_17007,N_14091,N_13299);
and U17008 (N_17008,N_14800,N_12081);
xnor U17009 (N_17009,N_14177,N_11497);
nand U17010 (N_17010,N_12850,N_12614);
and U17011 (N_17011,N_12827,N_11705);
nand U17012 (N_17012,N_10626,N_10045);
xnor U17013 (N_17013,N_11377,N_11806);
and U17014 (N_17014,N_14657,N_14630);
nand U17015 (N_17015,N_14815,N_12719);
nor U17016 (N_17016,N_14776,N_13008);
or U17017 (N_17017,N_10109,N_13189);
nand U17018 (N_17018,N_14981,N_14222);
xnor U17019 (N_17019,N_13493,N_13969);
nor U17020 (N_17020,N_14018,N_13494);
and U17021 (N_17021,N_13487,N_12969);
nand U17022 (N_17022,N_14272,N_14504);
nor U17023 (N_17023,N_11912,N_13810);
xor U17024 (N_17024,N_10316,N_13281);
nand U17025 (N_17025,N_10865,N_13867);
xnor U17026 (N_17026,N_14813,N_10739);
xnor U17027 (N_17027,N_13756,N_13286);
and U17028 (N_17028,N_12059,N_14556);
xnor U17029 (N_17029,N_10531,N_12510);
nor U17030 (N_17030,N_12826,N_11434);
nand U17031 (N_17031,N_13634,N_13013);
nand U17032 (N_17032,N_10022,N_12013);
or U17033 (N_17033,N_10125,N_11784);
or U17034 (N_17034,N_13327,N_13849);
nor U17035 (N_17035,N_11214,N_14848);
or U17036 (N_17036,N_14884,N_12217);
or U17037 (N_17037,N_10913,N_12583);
xor U17038 (N_17038,N_11729,N_14102);
or U17039 (N_17039,N_14280,N_13290);
nor U17040 (N_17040,N_14814,N_10092);
and U17041 (N_17041,N_13373,N_12124);
and U17042 (N_17042,N_13293,N_10985);
nor U17043 (N_17043,N_13971,N_14368);
and U17044 (N_17044,N_13551,N_11991);
and U17045 (N_17045,N_13992,N_12103);
nor U17046 (N_17046,N_12910,N_10885);
or U17047 (N_17047,N_13003,N_12503);
nand U17048 (N_17048,N_13069,N_14796);
and U17049 (N_17049,N_12578,N_11045);
and U17050 (N_17050,N_12618,N_14555);
and U17051 (N_17051,N_12925,N_10154);
nor U17052 (N_17052,N_14950,N_10390);
and U17053 (N_17053,N_10167,N_10227);
and U17054 (N_17054,N_14970,N_11031);
or U17055 (N_17055,N_14701,N_11005);
xnor U17056 (N_17056,N_13816,N_14482);
or U17057 (N_17057,N_13398,N_14392);
and U17058 (N_17058,N_13578,N_13909);
xnor U17059 (N_17059,N_12601,N_13068);
and U17060 (N_17060,N_10006,N_12352);
nand U17061 (N_17061,N_10290,N_13081);
or U17062 (N_17062,N_11897,N_12149);
nand U17063 (N_17063,N_11569,N_12764);
and U17064 (N_17064,N_14670,N_11124);
or U17065 (N_17065,N_11358,N_12674);
nor U17066 (N_17066,N_11978,N_14459);
and U17067 (N_17067,N_10187,N_11305);
xor U17068 (N_17068,N_12320,N_14427);
or U17069 (N_17069,N_12551,N_11217);
and U17070 (N_17070,N_13247,N_11824);
or U17071 (N_17071,N_14784,N_11378);
nand U17072 (N_17072,N_10963,N_12342);
nand U17073 (N_17073,N_10792,N_13151);
nor U17074 (N_17074,N_14547,N_12147);
xnor U17075 (N_17075,N_13613,N_13594);
or U17076 (N_17076,N_10917,N_10868);
xnor U17077 (N_17077,N_12275,N_13890);
nand U17078 (N_17078,N_13582,N_12537);
and U17079 (N_17079,N_13880,N_11962);
and U17080 (N_17080,N_10113,N_13981);
nand U17081 (N_17081,N_11713,N_13062);
nor U17082 (N_17082,N_14059,N_14046);
xor U17083 (N_17083,N_10280,N_10965);
xor U17084 (N_17084,N_10285,N_13249);
and U17085 (N_17085,N_13241,N_11973);
and U17086 (N_17086,N_12226,N_14216);
and U17087 (N_17087,N_11116,N_14940);
and U17088 (N_17088,N_11234,N_11778);
and U17089 (N_17089,N_13898,N_13741);
nor U17090 (N_17090,N_14625,N_13910);
nor U17091 (N_17091,N_13863,N_12080);
nor U17092 (N_17092,N_10020,N_14897);
or U17093 (N_17093,N_11591,N_12540);
nand U17094 (N_17094,N_12915,N_10081);
nand U17095 (N_17095,N_14678,N_10904);
or U17096 (N_17096,N_12439,N_14008);
nand U17097 (N_17097,N_11544,N_10354);
nand U17098 (N_17098,N_13215,N_11152);
nor U17099 (N_17099,N_11669,N_13091);
nor U17100 (N_17100,N_14407,N_14995);
xor U17101 (N_17101,N_10457,N_10701);
xor U17102 (N_17102,N_11472,N_14595);
and U17103 (N_17103,N_14327,N_13307);
nand U17104 (N_17104,N_14201,N_14155);
xor U17105 (N_17105,N_13612,N_12588);
or U17106 (N_17106,N_11517,N_12479);
xor U17107 (N_17107,N_13089,N_13007);
or U17108 (N_17108,N_14986,N_14446);
or U17109 (N_17109,N_12573,N_14856);
xor U17110 (N_17110,N_14261,N_10432);
and U17111 (N_17111,N_12435,N_14604);
nand U17112 (N_17112,N_12972,N_14265);
nor U17113 (N_17113,N_13536,N_10931);
nand U17114 (N_17114,N_13872,N_10488);
nor U17115 (N_17115,N_14983,N_11835);
nor U17116 (N_17116,N_12627,N_12939);
and U17117 (N_17117,N_13553,N_10943);
nor U17118 (N_17118,N_10147,N_14611);
nor U17119 (N_17119,N_11660,N_14471);
xnor U17120 (N_17120,N_10448,N_14126);
nor U17121 (N_17121,N_14558,N_11371);
or U17122 (N_17122,N_14429,N_10890);
and U17123 (N_17123,N_12068,N_12458);
and U17124 (N_17124,N_10005,N_12331);
nand U17125 (N_17125,N_11279,N_14436);
or U17126 (N_17126,N_14246,N_10554);
nand U17127 (N_17127,N_14671,N_10351);
and U17128 (N_17128,N_10644,N_14667);
or U17129 (N_17129,N_13823,N_10120);
and U17130 (N_17130,N_11158,N_10337);
xnor U17131 (N_17131,N_11141,N_10168);
or U17132 (N_17132,N_13663,N_11287);
nand U17133 (N_17133,N_10996,N_14987);
nand U17134 (N_17134,N_13259,N_10734);
and U17135 (N_17135,N_12062,N_11509);
nand U17136 (N_17136,N_12369,N_13088);
or U17137 (N_17137,N_11946,N_13066);
and U17138 (N_17138,N_13840,N_13379);
or U17139 (N_17139,N_14156,N_10543);
and U17140 (N_17140,N_13989,N_12077);
and U17141 (N_17141,N_11642,N_14658);
xnor U17142 (N_17142,N_14891,N_10770);
nand U17143 (N_17143,N_12505,N_11846);
or U17144 (N_17144,N_14793,N_13267);
and U17145 (N_17145,N_12308,N_12223);
or U17146 (N_17146,N_13535,N_10416);
nor U17147 (N_17147,N_14140,N_11080);
nor U17148 (N_17148,N_12229,N_13661);
or U17149 (N_17149,N_11661,N_11535);
or U17150 (N_17150,N_14224,N_12671);
nand U17151 (N_17151,N_14929,N_11563);
and U17152 (N_17152,N_14843,N_11605);
and U17153 (N_17153,N_14135,N_11268);
or U17154 (N_17154,N_13349,N_13801);
nand U17155 (N_17155,N_14931,N_10174);
and U17156 (N_17156,N_12958,N_11195);
xnor U17157 (N_17157,N_13265,N_12405);
or U17158 (N_17158,N_14248,N_13798);
or U17159 (N_17159,N_13611,N_14522);
nand U17160 (N_17160,N_13817,N_14518);
or U17161 (N_17161,N_14509,N_13407);
nand U17162 (N_17162,N_10564,N_11823);
xor U17163 (N_17163,N_14996,N_14149);
or U17164 (N_17164,N_12800,N_11474);
xor U17165 (N_17165,N_14037,N_11985);
or U17166 (N_17166,N_11135,N_10946);
nor U17167 (N_17167,N_12658,N_11111);
xnor U17168 (N_17168,N_13395,N_12729);
or U17169 (N_17169,N_14527,N_10160);
xor U17170 (N_17170,N_12889,N_13662);
nand U17171 (N_17171,N_13262,N_11275);
and U17172 (N_17172,N_12714,N_13603);
and U17173 (N_17173,N_12174,N_11974);
and U17174 (N_17174,N_13345,N_12057);
and U17175 (N_17175,N_12545,N_12072);
xnor U17176 (N_17176,N_10221,N_12821);
nand U17177 (N_17177,N_11796,N_12946);
and U17178 (N_17178,N_10268,N_11587);
xor U17179 (N_17179,N_10740,N_10721);
xor U17180 (N_17180,N_12566,N_13033);
nor U17181 (N_17181,N_14240,N_11197);
or U17182 (N_17182,N_10313,N_11181);
and U17183 (N_17183,N_10608,N_11810);
xor U17184 (N_17184,N_13420,N_11758);
xor U17185 (N_17185,N_12324,N_10086);
nor U17186 (N_17186,N_10822,N_14920);
and U17187 (N_17187,N_13664,N_10172);
nand U17188 (N_17188,N_12843,N_12567);
nor U17189 (N_17189,N_13513,N_13361);
and U17190 (N_17190,N_11402,N_10820);
xor U17191 (N_17191,N_12654,N_13688);
nand U17192 (N_17192,N_12580,N_12712);
nand U17193 (N_17193,N_12980,N_14192);
xnor U17194 (N_17194,N_13831,N_12670);
or U17195 (N_17195,N_13626,N_13163);
and U17196 (N_17196,N_11021,N_13656);
xnor U17197 (N_17197,N_14767,N_10882);
or U17198 (N_17198,N_10621,N_11271);
nor U17199 (N_17199,N_14264,N_11199);
xor U17200 (N_17200,N_12899,N_12349);
nor U17201 (N_17201,N_10889,N_10674);
and U17202 (N_17202,N_12971,N_14038);
or U17203 (N_17203,N_11588,N_11414);
nor U17204 (N_17204,N_14562,N_12465);
nor U17205 (N_17205,N_14590,N_10903);
nand U17206 (N_17206,N_11086,N_11286);
and U17207 (N_17207,N_10990,N_11194);
nand U17208 (N_17208,N_11067,N_14056);
nand U17209 (N_17209,N_13480,N_14416);
nor U17210 (N_17210,N_13246,N_14529);
xnor U17211 (N_17211,N_14169,N_10266);
xnor U17212 (N_17212,N_12185,N_10412);
nand U17213 (N_17213,N_14842,N_14434);
nor U17214 (N_17214,N_13170,N_14714);
or U17215 (N_17215,N_10301,N_10263);
nor U17216 (N_17216,N_10859,N_13268);
nand U17217 (N_17217,N_11388,N_10542);
nor U17218 (N_17218,N_13789,N_10957);
xor U17219 (N_17219,N_11041,N_13746);
and U17220 (N_17220,N_12433,N_13504);
and U17221 (N_17221,N_13539,N_10599);
nor U17222 (N_17222,N_10995,N_11596);
and U17223 (N_17223,N_10960,N_12252);
nand U17224 (N_17224,N_14684,N_10402);
nand U17225 (N_17225,N_10972,N_12541);
nor U17226 (N_17226,N_10347,N_12611);
nor U17227 (N_17227,N_11944,N_13422);
nor U17228 (N_17228,N_14199,N_13995);
or U17229 (N_17229,N_14762,N_10411);
nor U17230 (N_17230,N_13727,N_11100);
and U17231 (N_17231,N_12250,N_12263);
and U17232 (N_17232,N_12176,N_11473);
or U17233 (N_17233,N_13894,N_11345);
xor U17234 (N_17234,N_11913,N_10994);
nand U17235 (N_17235,N_10919,N_14711);
nor U17236 (N_17236,N_11667,N_11556);
and U17237 (N_17237,N_12517,N_12884);
or U17238 (N_17238,N_10878,N_14409);
or U17239 (N_17239,N_11292,N_11506);
nand U17240 (N_17240,N_12550,N_14517);
nand U17241 (N_17241,N_13121,N_13963);
nor U17242 (N_17242,N_12978,N_12296);
xor U17243 (N_17243,N_14511,N_12849);
nand U17244 (N_17244,N_13376,N_11594);
nand U17245 (N_17245,N_11334,N_11680);
nand U17246 (N_17246,N_10874,N_11453);
xnor U17247 (N_17247,N_13044,N_12467);
nand U17248 (N_17248,N_13677,N_12892);
and U17249 (N_17249,N_10743,N_10909);
and U17250 (N_17250,N_10234,N_13572);
xor U17251 (N_17251,N_10849,N_10091);
xnor U17252 (N_17252,N_14385,N_13112);
or U17253 (N_17253,N_12389,N_11907);
xnor U17254 (N_17254,N_13986,N_12440);
and U17255 (N_17255,N_10970,N_11346);
or U17256 (N_17256,N_13990,N_12322);
and U17257 (N_17257,N_13951,N_14857);
and U17258 (N_17258,N_11459,N_13654);
and U17259 (N_17259,N_10495,N_10510);
xor U17260 (N_17260,N_11932,N_13914);
and U17261 (N_17261,N_12665,N_14579);
nor U17262 (N_17262,N_11277,N_12198);
nor U17263 (N_17263,N_14820,N_10039);
xor U17264 (N_17264,N_14305,N_12965);
xor U17265 (N_17265,N_11213,N_13788);
nor U17266 (N_17266,N_13717,N_10704);
xnor U17267 (N_17267,N_14351,N_13120);
nand U17268 (N_17268,N_11036,N_12089);
nor U17269 (N_17269,N_12480,N_14503);
xor U17270 (N_17270,N_10192,N_10064);
nand U17271 (N_17271,N_12493,N_14957);
nand U17272 (N_17272,N_11019,N_11917);
or U17273 (N_17273,N_10034,N_14243);
and U17274 (N_17274,N_12700,N_13932);
nand U17275 (N_17275,N_12699,N_14299);
or U17276 (N_17276,N_13049,N_14053);
nor U17277 (N_17277,N_14298,N_11486);
xor U17278 (N_17278,N_12461,N_14801);
or U17279 (N_17279,N_14492,N_11620);
nor U17280 (N_17280,N_14367,N_12942);
xnor U17281 (N_17281,N_11380,N_12272);
xnor U17282 (N_17282,N_12334,N_10194);
or U17283 (N_17283,N_14898,N_14838);
and U17284 (N_17284,N_11360,N_11309);
and U17285 (N_17285,N_12082,N_13355);
xnor U17286 (N_17286,N_12370,N_11665);
or U17287 (N_17287,N_11952,N_10663);
or U17288 (N_17288,N_13842,N_14694);
or U17289 (N_17289,N_13641,N_14681);
or U17290 (N_17290,N_13941,N_14567);
and U17291 (N_17291,N_13651,N_14401);
nor U17292 (N_17292,N_11208,N_13028);
and U17293 (N_17293,N_11761,N_12728);
or U17294 (N_17294,N_10468,N_12726);
nor U17295 (N_17295,N_11949,N_13579);
xor U17296 (N_17296,N_11426,N_13484);
nand U17297 (N_17297,N_13790,N_14026);
xnor U17298 (N_17298,N_13050,N_12326);
nand U17299 (N_17299,N_11702,N_11804);
and U17300 (N_17300,N_11624,N_13275);
xnor U17301 (N_17301,N_12355,N_12810);
nor U17302 (N_17302,N_10208,N_14823);
or U17303 (N_17303,N_14909,N_13452);
nor U17304 (N_17304,N_11764,N_11171);
nand U17305 (N_17305,N_14483,N_11263);
nor U17306 (N_17306,N_10206,N_10460);
nand U17307 (N_17307,N_11218,N_14638);
nand U17308 (N_17308,N_14034,N_11026);
nand U17309 (N_17309,N_10038,N_12414);
nand U17310 (N_17310,N_12722,N_12973);
or U17311 (N_17311,N_11107,N_14780);
xor U17312 (N_17312,N_11750,N_13982);
nor U17313 (N_17313,N_13511,N_10320);
and U17314 (N_17314,N_10760,N_12835);
nor U17315 (N_17315,N_13414,N_14597);
and U17316 (N_17316,N_12794,N_12202);
or U17317 (N_17317,N_10832,N_12485);
nor U17318 (N_17318,N_11561,N_12298);
and U17319 (N_17319,N_10966,N_10429);
or U17320 (N_17320,N_14284,N_10420);
xor U17321 (N_17321,N_13655,N_10307);
nor U17322 (N_17322,N_12817,N_11131);
and U17323 (N_17323,N_13171,N_10422);
xor U17324 (N_17324,N_10654,N_14576);
nor U17325 (N_17325,N_14665,N_13413);
nand U17326 (N_17326,N_12233,N_14203);
nand U17327 (N_17327,N_10566,N_11536);
xnor U17328 (N_17328,N_12415,N_13165);
and U17329 (N_17329,N_14326,N_10196);
or U17330 (N_17330,N_14266,N_14672);
or U17331 (N_17331,N_10948,N_12542);
nor U17332 (N_17332,N_10729,N_14617);
xnor U17333 (N_17333,N_11054,N_10683);
and U17334 (N_17334,N_11298,N_14534);
xnor U17335 (N_17335,N_10059,N_10089);
nand U17336 (N_17336,N_14551,N_13744);
or U17337 (N_17337,N_13712,N_14173);
and U17338 (N_17338,N_11540,N_13110);
xnor U17339 (N_17339,N_11074,N_11821);
xor U17340 (N_17340,N_10771,N_13684);
and U17341 (N_17341,N_13158,N_13159);
nor U17342 (N_17342,N_14974,N_12262);
nand U17343 (N_17343,N_11028,N_10529);
nand U17344 (N_17344,N_13135,N_12471);
nand U17345 (N_17345,N_12796,N_12886);
nor U17346 (N_17346,N_11326,N_10690);
and U17347 (N_17347,N_10687,N_10357);
and U17348 (N_17348,N_12935,N_10586);
nand U17349 (N_17349,N_14598,N_11464);
nand U17350 (N_17350,N_11638,N_14346);
nand U17351 (N_17351,N_14951,N_11847);
nand U17352 (N_17352,N_12387,N_10906);
nand U17353 (N_17353,N_11727,N_14086);
and U17354 (N_17354,N_14015,N_13474);
and U17355 (N_17355,N_13304,N_12990);
and U17356 (N_17356,N_10118,N_11738);
or U17357 (N_17357,N_12422,N_12095);
and U17358 (N_17358,N_14236,N_11394);
nand U17359 (N_17359,N_13391,N_13797);
or U17360 (N_17360,N_10993,N_13288);
xor U17361 (N_17361,N_14816,N_11663);
nand U17362 (N_17362,N_13191,N_12172);
xor U17363 (N_17363,N_10437,N_13128);
nand U17364 (N_17364,N_13795,N_11950);
or U17365 (N_17365,N_12133,N_10145);
xor U17366 (N_17366,N_14984,N_10319);
nand U17367 (N_17367,N_12585,N_13960);
nor U17368 (N_17368,N_13243,N_12905);
or U17369 (N_17369,N_12069,N_12789);
nand U17370 (N_17370,N_12099,N_14963);
nand U17371 (N_17371,N_14868,N_14382);
xnor U17372 (N_17372,N_11904,N_11153);
or U17373 (N_17373,N_13785,N_12376);
or U17374 (N_17374,N_14063,N_11874);
nand U17375 (N_17375,N_10207,N_14777);
or U17376 (N_17376,N_11427,N_13037);
nand U17377 (N_17377,N_14085,N_13573);
xor U17378 (N_17378,N_14273,N_10391);
and U17379 (N_17379,N_10688,N_10384);
nor U17380 (N_17380,N_14572,N_14872);
xor U17381 (N_17381,N_13409,N_10364);
or U17382 (N_17382,N_10611,N_12024);
and U17383 (N_17383,N_10855,N_13210);
or U17384 (N_17384,N_13896,N_14911);
xnor U17385 (N_17385,N_14270,N_11461);
nand U17386 (N_17386,N_14178,N_12787);
and U17387 (N_17387,N_11037,N_11557);
or U17388 (N_17388,N_14841,N_13956);
xnor U17389 (N_17389,N_11205,N_13344);
or U17390 (N_17390,N_10369,N_10541);
xor U17391 (N_17391,N_12613,N_14923);
xnor U17392 (N_17392,N_14035,N_14756);
nand U17393 (N_17393,N_12701,N_14185);
xnor U17394 (N_17394,N_13146,N_11884);
xor U17395 (N_17395,N_12526,N_11325);
xor U17396 (N_17396,N_10857,N_10436);
nor U17397 (N_17397,N_11745,N_12707);
xor U17398 (N_17398,N_11262,N_12390);
xnor U17399 (N_17399,N_11682,N_13952);
nor U17400 (N_17400,N_11613,N_12677);
and U17401 (N_17401,N_11383,N_14837);
xnor U17402 (N_17402,N_13152,N_11766);
and U17403 (N_17403,N_10395,N_11157);
nor U17404 (N_17404,N_12751,N_13767);
nand U17405 (N_17405,N_14585,N_14835);
nand U17406 (N_17406,N_13292,N_10276);
xnor U17407 (N_17407,N_10031,N_10401);
nor U17408 (N_17408,N_14861,N_13313);
nor U17409 (N_17409,N_13733,N_11543);
nand U17410 (N_17410,N_10410,N_12890);
or U17411 (N_17411,N_11224,N_14402);
xnor U17412 (N_17412,N_12863,N_13871);
xor U17413 (N_17413,N_12347,N_14992);
and U17414 (N_17414,N_10937,N_14196);
nor U17415 (N_17415,N_11148,N_11529);
nand U17416 (N_17416,N_11243,N_13352);
nor U17417 (N_17417,N_11144,N_11281);
nand U17418 (N_17418,N_11993,N_12254);
or U17419 (N_17419,N_10902,N_10844);
or U17420 (N_17420,N_14437,N_11688);
or U17421 (N_17421,N_12725,N_11352);
and U17422 (N_17422,N_10017,N_11310);
nand U17423 (N_17423,N_11637,N_10060);
nand U17424 (N_17424,N_12994,N_13432);
nand U17425 (N_17425,N_12311,N_14910);
and U17426 (N_17426,N_12784,N_12278);
and U17427 (N_17427,N_13633,N_11366);
or U17428 (N_17428,N_12767,N_11790);
nor U17429 (N_17429,N_12872,N_12255);
or U17430 (N_17430,N_10104,N_14268);
nor U17431 (N_17431,N_10629,N_11361);
nor U17432 (N_17432,N_14123,N_13837);
nand U17433 (N_17433,N_13861,N_10133);
or U17434 (N_17434,N_11584,N_13792);
nor U17435 (N_17435,N_11886,N_10774);
xnor U17436 (N_17436,N_10454,N_11800);
nand U17437 (N_17437,N_13512,N_12065);
nor U17438 (N_17438,N_12033,N_10299);
xor U17439 (N_17439,N_14030,N_12612);
nand U17440 (N_17440,N_14912,N_11209);
or U17441 (N_17441,N_10397,N_14519);
xor U17442 (N_17442,N_13458,N_10214);
nand U17443 (N_17443,N_13636,N_10258);
nand U17444 (N_17444,N_14468,N_12780);
and U17445 (N_17445,N_12909,N_12586);
nand U17446 (N_17446,N_11433,N_11331);
or U17447 (N_17447,N_13437,N_13967);
or U17448 (N_17448,N_10838,N_10570);
and U17449 (N_17449,N_11595,N_10722);
xor U17450 (N_17450,N_14039,N_10512);
and U17451 (N_17451,N_12128,N_12643);
and U17452 (N_17452,N_13783,N_14989);
or U17453 (N_17453,N_12476,N_12182);
and U17454 (N_17454,N_12211,N_14287);
xnor U17455 (N_17455,N_12975,N_13387);
and U17456 (N_17456,N_11984,N_14862);
nor U17457 (N_17457,N_12659,N_12418);
and U17458 (N_17458,N_11487,N_13968);
xor U17459 (N_17459,N_10956,N_14631);
xor U17460 (N_17460,N_12698,N_10719);
or U17461 (N_17461,N_14221,N_13000);
nand U17462 (N_17462,N_10969,N_11084);
nand U17463 (N_17463,N_13825,N_10602);
nor U17464 (N_17464,N_11105,N_13723);
or U17465 (N_17465,N_11498,N_14042);
nor U17466 (N_17466,N_14557,N_10573);
and U17467 (N_17467,N_13453,N_14151);
or U17468 (N_17468,N_10949,N_13052);
and U17469 (N_17469,N_10842,N_13499);
or U17470 (N_17470,N_10184,N_12575);
nand U17471 (N_17471,N_13934,N_13107);
nor U17472 (N_17472,N_11502,N_11901);
nor U17473 (N_17473,N_10321,N_13229);
xnor U17474 (N_17474,N_14825,N_13501);
nor U17475 (N_17475,N_11537,N_14973);
and U17476 (N_17476,N_12445,N_10408);
nand U17477 (N_17477,N_10716,N_11438);
and U17478 (N_17478,N_13887,N_11769);
or U17479 (N_17479,N_10610,N_13445);
nand U17480 (N_17480,N_14739,N_13350);
nand U17481 (N_17481,N_11455,N_10230);
xnor U17482 (N_17482,N_14706,N_13460);
xor U17483 (N_17483,N_14453,N_12696);
xor U17484 (N_17484,N_12408,N_10784);
nand U17485 (N_17485,N_14211,N_13905);
xnor U17486 (N_17486,N_10098,N_11320);
or U17487 (N_17487,N_12494,N_14179);
nand U17488 (N_17488,N_11376,N_11354);
and U17489 (N_17489,N_11649,N_10809);
nand U17490 (N_17490,N_11858,N_10052);
or U17491 (N_17491,N_11278,N_12199);
nand U17492 (N_17492,N_11174,N_12097);
and U17493 (N_17493,N_14610,N_12121);
nor U17494 (N_17494,N_12307,N_13520);
or U17495 (N_17495,N_12562,N_11577);
or U17496 (N_17496,N_13617,N_12184);
and U17497 (N_17497,N_11992,N_11724);
nand U17498 (N_17498,N_13857,N_11664);
and U17499 (N_17499,N_12191,N_10324);
xnor U17500 (N_17500,N_11780,N_14745);
xnor U17501 (N_17501,N_12221,N_14914);
and U17502 (N_17502,N_10878,N_13053);
and U17503 (N_17503,N_13278,N_12490);
xor U17504 (N_17504,N_14490,N_14275);
or U17505 (N_17505,N_14122,N_12168);
nor U17506 (N_17506,N_13957,N_10642);
nor U17507 (N_17507,N_11031,N_13182);
nand U17508 (N_17508,N_11369,N_10751);
or U17509 (N_17509,N_10151,N_11174);
xnor U17510 (N_17510,N_12122,N_13136);
xor U17511 (N_17511,N_11808,N_12972);
xor U17512 (N_17512,N_13504,N_12985);
and U17513 (N_17513,N_10729,N_13381);
nand U17514 (N_17514,N_14897,N_11226);
and U17515 (N_17515,N_12352,N_11924);
xor U17516 (N_17516,N_13188,N_13845);
nor U17517 (N_17517,N_14572,N_13096);
nor U17518 (N_17518,N_11302,N_12134);
xor U17519 (N_17519,N_12050,N_10860);
or U17520 (N_17520,N_13065,N_10214);
or U17521 (N_17521,N_11240,N_10661);
nand U17522 (N_17522,N_10306,N_11916);
nand U17523 (N_17523,N_12018,N_10051);
and U17524 (N_17524,N_13846,N_10542);
xor U17525 (N_17525,N_10450,N_14561);
nor U17526 (N_17526,N_14570,N_13077);
xnor U17527 (N_17527,N_13788,N_10319);
xor U17528 (N_17528,N_13275,N_13564);
nand U17529 (N_17529,N_14870,N_12321);
or U17530 (N_17530,N_12960,N_10294);
or U17531 (N_17531,N_13082,N_14337);
xnor U17532 (N_17532,N_13211,N_11965);
nor U17533 (N_17533,N_10914,N_10392);
nor U17534 (N_17534,N_13249,N_10283);
or U17535 (N_17535,N_11032,N_11593);
and U17536 (N_17536,N_13803,N_10798);
nand U17537 (N_17537,N_14173,N_14505);
and U17538 (N_17538,N_11418,N_14052);
or U17539 (N_17539,N_11334,N_10575);
or U17540 (N_17540,N_10780,N_12327);
nand U17541 (N_17541,N_13282,N_10203);
xnor U17542 (N_17542,N_11264,N_14993);
nand U17543 (N_17543,N_14974,N_12390);
nor U17544 (N_17544,N_14955,N_10369);
nor U17545 (N_17545,N_14260,N_14837);
xnor U17546 (N_17546,N_14281,N_11033);
nand U17547 (N_17547,N_10797,N_14082);
xnor U17548 (N_17548,N_14942,N_14259);
nand U17549 (N_17549,N_11720,N_10788);
nand U17550 (N_17550,N_12300,N_14533);
nor U17551 (N_17551,N_14265,N_12727);
xnor U17552 (N_17552,N_14246,N_11443);
nor U17553 (N_17553,N_13167,N_11172);
xor U17554 (N_17554,N_10023,N_14600);
or U17555 (N_17555,N_14900,N_11931);
nand U17556 (N_17556,N_11712,N_10665);
or U17557 (N_17557,N_13869,N_10665);
nand U17558 (N_17558,N_12612,N_12107);
nor U17559 (N_17559,N_11387,N_13206);
xor U17560 (N_17560,N_13706,N_12715);
nor U17561 (N_17561,N_12982,N_11643);
xor U17562 (N_17562,N_14165,N_11734);
nor U17563 (N_17563,N_11711,N_13504);
nor U17564 (N_17564,N_12262,N_11201);
and U17565 (N_17565,N_11186,N_14187);
xor U17566 (N_17566,N_12682,N_13149);
nand U17567 (N_17567,N_10295,N_14322);
and U17568 (N_17568,N_13391,N_14461);
nor U17569 (N_17569,N_14797,N_14563);
nor U17570 (N_17570,N_11330,N_13363);
nor U17571 (N_17571,N_13060,N_14270);
or U17572 (N_17572,N_12607,N_12083);
nand U17573 (N_17573,N_14029,N_10646);
nor U17574 (N_17574,N_14885,N_10394);
xor U17575 (N_17575,N_14741,N_12589);
or U17576 (N_17576,N_12385,N_10329);
nand U17577 (N_17577,N_10193,N_14711);
or U17578 (N_17578,N_13021,N_13770);
xnor U17579 (N_17579,N_14014,N_12147);
nor U17580 (N_17580,N_13517,N_11705);
or U17581 (N_17581,N_14094,N_14468);
nand U17582 (N_17582,N_13215,N_11205);
xor U17583 (N_17583,N_14137,N_10102);
nor U17584 (N_17584,N_14064,N_14754);
nor U17585 (N_17585,N_11170,N_11466);
nor U17586 (N_17586,N_13764,N_14890);
xor U17587 (N_17587,N_12303,N_10061);
or U17588 (N_17588,N_14479,N_14971);
xor U17589 (N_17589,N_10753,N_13503);
or U17590 (N_17590,N_12393,N_10439);
xor U17591 (N_17591,N_12949,N_12326);
xor U17592 (N_17592,N_14906,N_14749);
or U17593 (N_17593,N_12690,N_12663);
or U17594 (N_17594,N_13905,N_13368);
xor U17595 (N_17595,N_14209,N_13807);
nand U17596 (N_17596,N_11054,N_12047);
nand U17597 (N_17597,N_10997,N_13138);
xnor U17598 (N_17598,N_10507,N_14729);
or U17599 (N_17599,N_11717,N_14389);
or U17600 (N_17600,N_11104,N_13768);
or U17601 (N_17601,N_10302,N_14246);
and U17602 (N_17602,N_11437,N_13159);
nand U17603 (N_17603,N_10362,N_11461);
or U17604 (N_17604,N_13223,N_12946);
or U17605 (N_17605,N_13823,N_10855);
and U17606 (N_17606,N_10326,N_14893);
and U17607 (N_17607,N_12935,N_11463);
nor U17608 (N_17608,N_10052,N_12399);
nand U17609 (N_17609,N_12952,N_12412);
and U17610 (N_17610,N_14378,N_13272);
and U17611 (N_17611,N_13371,N_12208);
nand U17612 (N_17612,N_12174,N_11990);
xor U17613 (N_17613,N_10333,N_13896);
xnor U17614 (N_17614,N_13927,N_11761);
xor U17615 (N_17615,N_11947,N_11969);
and U17616 (N_17616,N_13704,N_12977);
xor U17617 (N_17617,N_14261,N_10026);
xor U17618 (N_17618,N_12764,N_10306);
or U17619 (N_17619,N_13663,N_13610);
nor U17620 (N_17620,N_13970,N_13529);
and U17621 (N_17621,N_12430,N_10573);
nor U17622 (N_17622,N_14753,N_10285);
nand U17623 (N_17623,N_11328,N_11786);
nand U17624 (N_17624,N_13082,N_13812);
nand U17625 (N_17625,N_10197,N_11049);
xor U17626 (N_17626,N_13973,N_12636);
nor U17627 (N_17627,N_14174,N_12002);
nor U17628 (N_17628,N_13864,N_11123);
nor U17629 (N_17629,N_10177,N_14982);
xor U17630 (N_17630,N_14942,N_12823);
and U17631 (N_17631,N_14153,N_13630);
xor U17632 (N_17632,N_14585,N_10253);
nand U17633 (N_17633,N_11337,N_11879);
xnor U17634 (N_17634,N_10074,N_10879);
and U17635 (N_17635,N_13483,N_10257);
xor U17636 (N_17636,N_12885,N_11289);
and U17637 (N_17637,N_10777,N_13204);
and U17638 (N_17638,N_11073,N_13764);
or U17639 (N_17639,N_12013,N_12661);
xor U17640 (N_17640,N_11248,N_14541);
nor U17641 (N_17641,N_12144,N_12057);
and U17642 (N_17642,N_12083,N_13709);
nor U17643 (N_17643,N_13321,N_11292);
and U17644 (N_17644,N_14588,N_13110);
or U17645 (N_17645,N_13907,N_13326);
or U17646 (N_17646,N_14728,N_10843);
or U17647 (N_17647,N_11532,N_13749);
xnor U17648 (N_17648,N_11579,N_11796);
nor U17649 (N_17649,N_13876,N_12267);
nor U17650 (N_17650,N_11816,N_14663);
and U17651 (N_17651,N_11949,N_13761);
xnor U17652 (N_17652,N_13202,N_14995);
xor U17653 (N_17653,N_14608,N_11866);
and U17654 (N_17654,N_10485,N_13163);
xor U17655 (N_17655,N_14024,N_14047);
nor U17656 (N_17656,N_10510,N_12155);
and U17657 (N_17657,N_13594,N_14505);
or U17658 (N_17658,N_12974,N_13758);
nor U17659 (N_17659,N_11712,N_13338);
and U17660 (N_17660,N_11627,N_11140);
xor U17661 (N_17661,N_11763,N_13701);
xor U17662 (N_17662,N_14329,N_11847);
nand U17663 (N_17663,N_10416,N_11415);
or U17664 (N_17664,N_12100,N_13803);
nand U17665 (N_17665,N_10045,N_13572);
and U17666 (N_17666,N_12972,N_14428);
or U17667 (N_17667,N_14074,N_14232);
or U17668 (N_17668,N_13787,N_14279);
and U17669 (N_17669,N_13607,N_13982);
and U17670 (N_17670,N_12294,N_13819);
or U17671 (N_17671,N_12113,N_11458);
and U17672 (N_17672,N_13129,N_13912);
and U17673 (N_17673,N_14452,N_10673);
nor U17674 (N_17674,N_11522,N_11462);
and U17675 (N_17675,N_14110,N_12195);
and U17676 (N_17676,N_13300,N_14606);
or U17677 (N_17677,N_10798,N_12450);
nor U17678 (N_17678,N_10771,N_14455);
nand U17679 (N_17679,N_14292,N_13772);
xnor U17680 (N_17680,N_11277,N_10429);
nor U17681 (N_17681,N_13734,N_14173);
and U17682 (N_17682,N_12882,N_13197);
nand U17683 (N_17683,N_14545,N_13936);
and U17684 (N_17684,N_13923,N_12914);
or U17685 (N_17685,N_13148,N_10320);
or U17686 (N_17686,N_14527,N_14036);
nand U17687 (N_17687,N_14930,N_14197);
and U17688 (N_17688,N_10710,N_12203);
xor U17689 (N_17689,N_12223,N_12551);
or U17690 (N_17690,N_12229,N_10374);
nor U17691 (N_17691,N_11554,N_13280);
and U17692 (N_17692,N_12301,N_13027);
or U17693 (N_17693,N_10250,N_12887);
and U17694 (N_17694,N_13840,N_13333);
and U17695 (N_17695,N_11376,N_12603);
nand U17696 (N_17696,N_10678,N_10786);
xor U17697 (N_17697,N_13748,N_11396);
or U17698 (N_17698,N_10439,N_11645);
or U17699 (N_17699,N_12592,N_11730);
or U17700 (N_17700,N_12368,N_12544);
xor U17701 (N_17701,N_12177,N_14108);
nand U17702 (N_17702,N_10035,N_14104);
or U17703 (N_17703,N_10925,N_11450);
and U17704 (N_17704,N_10602,N_14335);
and U17705 (N_17705,N_10267,N_14669);
or U17706 (N_17706,N_14424,N_14429);
xnor U17707 (N_17707,N_11682,N_14218);
or U17708 (N_17708,N_13297,N_12307);
xnor U17709 (N_17709,N_13888,N_14365);
or U17710 (N_17710,N_10495,N_13583);
nor U17711 (N_17711,N_10881,N_14020);
nor U17712 (N_17712,N_14635,N_12964);
or U17713 (N_17713,N_13679,N_10680);
and U17714 (N_17714,N_10398,N_12839);
nand U17715 (N_17715,N_13689,N_14866);
xor U17716 (N_17716,N_13785,N_14135);
and U17717 (N_17717,N_13504,N_12584);
nand U17718 (N_17718,N_14390,N_12261);
xnor U17719 (N_17719,N_12679,N_12071);
or U17720 (N_17720,N_13086,N_10250);
or U17721 (N_17721,N_11840,N_13822);
and U17722 (N_17722,N_11743,N_10189);
nand U17723 (N_17723,N_13265,N_10682);
or U17724 (N_17724,N_11020,N_12514);
nor U17725 (N_17725,N_11484,N_13356);
xor U17726 (N_17726,N_13154,N_10146);
nand U17727 (N_17727,N_12913,N_10702);
nor U17728 (N_17728,N_14484,N_11171);
nor U17729 (N_17729,N_10755,N_11401);
xnor U17730 (N_17730,N_12692,N_11776);
or U17731 (N_17731,N_11939,N_10724);
nor U17732 (N_17732,N_11799,N_13092);
nor U17733 (N_17733,N_12766,N_13252);
nand U17734 (N_17734,N_11022,N_14134);
or U17735 (N_17735,N_13854,N_11085);
xnor U17736 (N_17736,N_10400,N_11169);
or U17737 (N_17737,N_12472,N_12860);
and U17738 (N_17738,N_11865,N_12213);
and U17739 (N_17739,N_10591,N_12508);
and U17740 (N_17740,N_11316,N_10893);
nor U17741 (N_17741,N_14692,N_10595);
nor U17742 (N_17742,N_12592,N_13736);
nand U17743 (N_17743,N_11374,N_12972);
nand U17744 (N_17744,N_13965,N_13820);
and U17745 (N_17745,N_13268,N_11915);
or U17746 (N_17746,N_10963,N_12374);
and U17747 (N_17747,N_14646,N_12430);
nand U17748 (N_17748,N_14279,N_12046);
nor U17749 (N_17749,N_11731,N_14828);
nor U17750 (N_17750,N_14550,N_11332);
nand U17751 (N_17751,N_14869,N_11326);
nor U17752 (N_17752,N_11784,N_11564);
and U17753 (N_17753,N_12964,N_11194);
xnor U17754 (N_17754,N_14488,N_10208);
nand U17755 (N_17755,N_13563,N_13530);
nand U17756 (N_17756,N_11663,N_13438);
nor U17757 (N_17757,N_13885,N_13945);
nand U17758 (N_17758,N_14065,N_12977);
nand U17759 (N_17759,N_14573,N_14306);
nor U17760 (N_17760,N_13084,N_11395);
and U17761 (N_17761,N_10574,N_14513);
nand U17762 (N_17762,N_12425,N_11551);
nand U17763 (N_17763,N_10652,N_14575);
nor U17764 (N_17764,N_12739,N_13984);
and U17765 (N_17765,N_11719,N_13745);
or U17766 (N_17766,N_14873,N_10229);
nand U17767 (N_17767,N_12534,N_13335);
xor U17768 (N_17768,N_13352,N_14707);
xnor U17769 (N_17769,N_12414,N_10416);
xor U17770 (N_17770,N_12201,N_12052);
nor U17771 (N_17771,N_10746,N_13806);
xnor U17772 (N_17772,N_14359,N_14433);
xor U17773 (N_17773,N_14462,N_10196);
nor U17774 (N_17774,N_12111,N_13958);
and U17775 (N_17775,N_11486,N_11000);
nor U17776 (N_17776,N_12627,N_13202);
nor U17777 (N_17777,N_11603,N_14148);
or U17778 (N_17778,N_13324,N_13111);
and U17779 (N_17779,N_14988,N_14423);
xnor U17780 (N_17780,N_10226,N_13319);
nand U17781 (N_17781,N_11039,N_14462);
nand U17782 (N_17782,N_13598,N_10120);
or U17783 (N_17783,N_11723,N_10695);
nand U17784 (N_17784,N_11744,N_10118);
or U17785 (N_17785,N_11520,N_10780);
xnor U17786 (N_17786,N_13868,N_13148);
nand U17787 (N_17787,N_12442,N_12195);
nor U17788 (N_17788,N_11671,N_13755);
nand U17789 (N_17789,N_10247,N_10976);
nand U17790 (N_17790,N_12708,N_10812);
nand U17791 (N_17791,N_10299,N_14158);
or U17792 (N_17792,N_12988,N_14588);
nor U17793 (N_17793,N_14073,N_10690);
nor U17794 (N_17794,N_13366,N_11068);
nor U17795 (N_17795,N_12849,N_10463);
or U17796 (N_17796,N_14995,N_10871);
or U17797 (N_17797,N_13938,N_10662);
or U17798 (N_17798,N_14904,N_14741);
or U17799 (N_17799,N_12175,N_11121);
nor U17800 (N_17800,N_13203,N_13952);
or U17801 (N_17801,N_13516,N_13322);
nand U17802 (N_17802,N_13851,N_11234);
or U17803 (N_17803,N_11412,N_13506);
nor U17804 (N_17804,N_13948,N_12083);
and U17805 (N_17805,N_13858,N_12217);
and U17806 (N_17806,N_12447,N_14312);
and U17807 (N_17807,N_14311,N_13201);
nor U17808 (N_17808,N_10152,N_12897);
nand U17809 (N_17809,N_11517,N_10366);
nor U17810 (N_17810,N_14064,N_14453);
and U17811 (N_17811,N_10039,N_12669);
xor U17812 (N_17812,N_13845,N_13744);
and U17813 (N_17813,N_12233,N_11207);
or U17814 (N_17814,N_14897,N_11122);
nand U17815 (N_17815,N_13869,N_12323);
or U17816 (N_17816,N_14538,N_12382);
and U17817 (N_17817,N_11699,N_12111);
and U17818 (N_17818,N_11773,N_11024);
or U17819 (N_17819,N_14488,N_11757);
nand U17820 (N_17820,N_11029,N_11971);
or U17821 (N_17821,N_13191,N_14123);
nor U17822 (N_17822,N_14500,N_14508);
xnor U17823 (N_17823,N_14360,N_12903);
or U17824 (N_17824,N_14198,N_13020);
or U17825 (N_17825,N_10326,N_10879);
nand U17826 (N_17826,N_12075,N_10989);
xor U17827 (N_17827,N_14684,N_13175);
or U17828 (N_17828,N_12459,N_13119);
nand U17829 (N_17829,N_12798,N_10658);
or U17830 (N_17830,N_13364,N_12541);
or U17831 (N_17831,N_11520,N_13198);
nor U17832 (N_17832,N_14584,N_10559);
nand U17833 (N_17833,N_13059,N_12279);
nor U17834 (N_17834,N_13670,N_10515);
xnor U17835 (N_17835,N_11593,N_10556);
nor U17836 (N_17836,N_11554,N_11821);
nor U17837 (N_17837,N_10880,N_12672);
nor U17838 (N_17838,N_14317,N_14128);
nor U17839 (N_17839,N_11195,N_11715);
xor U17840 (N_17840,N_14783,N_13301);
and U17841 (N_17841,N_11387,N_10598);
nor U17842 (N_17842,N_11294,N_14231);
and U17843 (N_17843,N_11288,N_11556);
xnor U17844 (N_17844,N_12511,N_12093);
xor U17845 (N_17845,N_13177,N_10678);
nand U17846 (N_17846,N_14640,N_13508);
nand U17847 (N_17847,N_12542,N_14087);
xnor U17848 (N_17848,N_10920,N_14125);
nand U17849 (N_17849,N_14963,N_10221);
nand U17850 (N_17850,N_12750,N_11478);
nand U17851 (N_17851,N_12845,N_10335);
nand U17852 (N_17852,N_14153,N_13533);
and U17853 (N_17853,N_10178,N_12349);
or U17854 (N_17854,N_11352,N_12548);
xnor U17855 (N_17855,N_14453,N_14653);
nand U17856 (N_17856,N_12023,N_11505);
or U17857 (N_17857,N_12411,N_10483);
xor U17858 (N_17858,N_10761,N_11401);
or U17859 (N_17859,N_12050,N_11638);
nor U17860 (N_17860,N_12748,N_10341);
or U17861 (N_17861,N_12739,N_12599);
nor U17862 (N_17862,N_14374,N_10028);
and U17863 (N_17863,N_11732,N_14860);
nand U17864 (N_17864,N_12203,N_12294);
or U17865 (N_17865,N_13975,N_12174);
or U17866 (N_17866,N_12100,N_12488);
xnor U17867 (N_17867,N_11142,N_12478);
nor U17868 (N_17868,N_12280,N_13389);
xor U17869 (N_17869,N_14966,N_10934);
nand U17870 (N_17870,N_14186,N_12129);
nand U17871 (N_17871,N_13857,N_10401);
and U17872 (N_17872,N_12329,N_13916);
nand U17873 (N_17873,N_13543,N_13093);
and U17874 (N_17874,N_12919,N_11739);
nand U17875 (N_17875,N_14015,N_14780);
xor U17876 (N_17876,N_12856,N_11724);
or U17877 (N_17877,N_10523,N_14898);
nor U17878 (N_17878,N_14652,N_14843);
and U17879 (N_17879,N_14500,N_10909);
xnor U17880 (N_17880,N_10963,N_10966);
xnor U17881 (N_17881,N_14177,N_13037);
nand U17882 (N_17882,N_13985,N_13683);
and U17883 (N_17883,N_13292,N_11674);
or U17884 (N_17884,N_13433,N_12634);
nand U17885 (N_17885,N_12858,N_13380);
nor U17886 (N_17886,N_11871,N_10425);
or U17887 (N_17887,N_14807,N_12951);
nor U17888 (N_17888,N_12562,N_11720);
and U17889 (N_17889,N_13304,N_10270);
nor U17890 (N_17890,N_10825,N_12543);
nand U17891 (N_17891,N_13108,N_13369);
nand U17892 (N_17892,N_10314,N_14646);
xnor U17893 (N_17893,N_13147,N_14680);
and U17894 (N_17894,N_14599,N_12258);
and U17895 (N_17895,N_13143,N_10835);
or U17896 (N_17896,N_10191,N_10121);
or U17897 (N_17897,N_13521,N_10615);
nor U17898 (N_17898,N_10629,N_13289);
or U17899 (N_17899,N_13495,N_12260);
xor U17900 (N_17900,N_11415,N_12428);
or U17901 (N_17901,N_12267,N_11565);
nand U17902 (N_17902,N_10226,N_10758);
or U17903 (N_17903,N_12866,N_13787);
xnor U17904 (N_17904,N_13411,N_10972);
and U17905 (N_17905,N_10364,N_10590);
or U17906 (N_17906,N_10289,N_11743);
or U17907 (N_17907,N_14033,N_11571);
nor U17908 (N_17908,N_13225,N_11090);
xnor U17909 (N_17909,N_10562,N_10361);
nor U17910 (N_17910,N_13836,N_13573);
nor U17911 (N_17911,N_13631,N_13903);
xnor U17912 (N_17912,N_13612,N_12084);
nor U17913 (N_17913,N_14516,N_10652);
nand U17914 (N_17914,N_11412,N_14997);
nor U17915 (N_17915,N_14056,N_10902);
or U17916 (N_17916,N_11818,N_14243);
or U17917 (N_17917,N_12607,N_13716);
or U17918 (N_17918,N_10271,N_13370);
and U17919 (N_17919,N_11188,N_14683);
and U17920 (N_17920,N_13464,N_11956);
xor U17921 (N_17921,N_12913,N_10466);
or U17922 (N_17922,N_11236,N_14009);
xor U17923 (N_17923,N_11118,N_13764);
xnor U17924 (N_17924,N_12075,N_12096);
xor U17925 (N_17925,N_11897,N_10007);
nor U17926 (N_17926,N_11934,N_10367);
and U17927 (N_17927,N_14589,N_11910);
xor U17928 (N_17928,N_13853,N_14643);
xnor U17929 (N_17929,N_12404,N_13980);
or U17930 (N_17930,N_14791,N_12144);
nand U17931 (N_17931,N_14521,N_10578);
and U17932 (N_17932,N_12072,N_10915);
and U17933 (N_17933,N_13196,N_12787);
nor U17934 (N_17934,N_14350,N_12118);
xnor U17935 (N_17935,N_14403,N_12360);
or U17936 (N_17936,N_12805,N_13484);
xnor U17937 (N_17937,N_13982,N_10591);
nand U17938 (N_17938,N_12776,N_12071);
nor U17939 (N_17939,N_10624,N_11679);
and U17940 (N_17940,N_14554,N_11478);
or U17941 (N_17941,N_11675,N_13367);
nor U17942 (N_17942,N_11109,N_10949);
xnor U17943 (N_17943,N_10689,N_14309);
nor U17944 (N_17944,N_13856,N_13816);
and U17945 (N_17945,N_14973,N_14557);
nor U17946 (N_17946,N_10134,N_13707);
nor U17947 (N_17947,N_11800,N_10178);
nor U17948 (N_17948,N_14544,N_12600);
or U17949 (N_17949,N_13467,N_11325);
nor U17950 (N_17950,N_11259,N_11886);
nand U17951 (N_17951,N_12113,N_13246);
nand U17952 (N_17952,N_12098,N_11044);
and U17953 (N_17953,N_11799,N_10862);
nor U17954 (N_17954,N_10378,N_10104);
or U17955 (N_17955,N_10077,N_12056);
or U17956 (N_17956,N_11032,N_10798);
nor U17957 (N_17957,N_13760,N_13642);
nand U17958 (N_17958,N_12200,N_13100);
xnor U17959 (N_17959,N_11741,N_10903);
or U17960 (N_17960,N_14766,N_11005);
and U17961 (N_17961,N_12209,N_14154);
nand U17962 (N_17962,N_13324,N_10039);
xnor U17963 (N_17963,N_13166,N_14132);
or U17964 (N_17964,N_11296,N_11542);
or U17965 (N_17965,N_14042,N_10005);
nand U17966 (N_17966,N_10094,N_13624);
nand U17967 (N_17967,N_11577,N_13258);
and U17968 (N_17968,N_11766,N_11177);
and U17969 (N_17969,N_14852,N_13960);
or U17970 (N_17970,N_14778,N_10797);
nand U17971 (N_17971,N_10204,N_13725);
nand U17972 (N_17972,N_10545,N_12998);
nand U17973 (N_17973,N_14193,N_10824);
nor U17974 (N_17974,N_14759,N_11046);
xnor U17975 (N_17975,N_10159,N_11334);
nand U17976 (N_17976,N_10279,N_12084);
xnor U17977 (N_17977,N_11750,N_11288);
xor U17978 (N_17978,N_11325,N_11217);
xor U17979 (N_17979,N_13220,N_13228);
xor U17980 (N_17980,N_13011,N_13086);
xnor U17981 (N_17981,N_14843,N_13731);
nor U17982 (N_17982,N_13790,N_12583);
nor U17983 (N_17983,N_11612,N_11567);
nand U17984 (N_17984,N_10543,N_12173);
nor U17985 (N_17985,N_11420,N_11660);
or U17986 (N_17986,N_10781,N_13641);
nor U17987 (N_17987,N_11050,N_12612);
xor U17988 (N_17988,N_11823,N_14361);
nand U17989 (N_17989,N_11094,N_12097);
nand U17990 (N_17990,N_10756,N_12195);
and U17991 (N_17991,N_12354,N_10940);
and U17992 (N_17992,N_11649,N_13715);
nand U17993 (N_17993,N_11882,N_13413);
and U17994 (N_17994,N_10189,N_10818);
nor U17995 (N_17995,N_12749,N_13743);
xnor U17996 (N_17996,N_10108,N_14340);
nor U17997 (N_17997,N_13654,N_12057);
or U17998 (N_17998,N_14430,N_12496);
nand U17999 (N_17999,N_11452,N_13667);
nand U18000 (N_18000,N_13357,N_12081);
or U18001 (N_18001,N_10370,N_11717);
and U18002 (N_18002,N_13489,N_13528);
nor U18003 (N_18003,N_14356,N_10313);
nand U18004 (N_18004,N_13665,N_10065);
xnor U18005 (N_18005,N_12166,N_10465);
xnor U18006 (N_18006,N_12044,N_11904);
or U18007 (N_18007,N_10040,N_13499);
xor U18008 (N_18008,N_13567,N_11190);
xor U18009 (N_18009,N_11354,N_14455);
nand U18010 (N_18010,N_11853,N_13670);
nor U18011 (N_18011,N_14494,N_14278);
nand U18012 (N_18012,N_10894,N_10337);
and U18013 (N_18013,N_12511,N_10209);
xnor U18014 (N_18014,N_12920,N_12131);
nand U18015 (N_18015,N_12098,N_14419);
and U18016 (N_18016,N_11160,N_11273);
xnor U18017 (N_18017,N_14513,N_14891);
nand U18018 (N_18018,N_13774,N_14555);
nand U18019 (N_18019,N_10749,N_11488);
or U18020 (N_18020,N_13415,N_11655);
and U18021 (N_18021,N_10782,N_11018);
or U18022 (N_18022,N_14305,N_13903);
xnor U18023 (N_18023,N_13413,N_11564);
xor U18024 (N_18024,N_13333,N_10519);
nand U18025 (N_18025,N_12048,N_13823);
nor U18026 (N_18026,N_12022,N_10720);
nor U18027 (N_18027,N_11814,N_10043);
nand U18028 (N_18028,N_11258,N_10884);
nor U18029 (N_18029,N_12204,N_13249);
nand U18030 (N_18030,N_11995,N_13880);
and U18031 (N_18031,N_13511,N_11507);
xnor U18032 (N_18032,N_13524,N_11776);
or U18033 (N_18033,N_11628,N_10457);
nor U18034 (N_18034,N_11098,N_13731);
xor U18035 (N_18035,N_14158,N_14128);
or U18036 (N_18036,N_10886,N_10993);
and U18037 (N_18037,N_10457,N_14734);
nand U18038 (N_18038,N_12827,N_11542);
and U18039 (N_18039,N_12752,N_11600);
xor U18040 (N_18040,N_14191,N_10012);
and U18041 (N_18041,N_14553,N_13338);
nor U18042 (N_18042,N_14749,N_11844);
or U18043 (N_18043,N_10973,N_10099);
or U18044 (N_18044,N_11634,N_13168);
nor U18045 (N_18045,N_10211,N_11297);
or U18046 (N_18046,N_13070,N_13654);
nand U18047 (N_18047,N_14508,N_14165);
xnor U18048 (N_18048,N_10884,N_11304);
and U18049 (N_18049,N_13865,N_14066);
and U18050 (N_18050,N_13770,N_13751);
xor U18051 (N_18051,N_11083,N_10795);
or U18052 (N_18052,N_14407,N_11502);
or U18053 (N_18053,N_11792,N_13551);
nand U18054 (N_18054,N_14746,N_10299);
and U18055 (N_18055,N_12612,N_10214);
xor U18056 (N_18056,N_12899,N_10495);
and U18057 (N_18057,N_14370,N_10805);
or U18058 (N_18058,N_13986,N_10998);
nand U18059 (N_18059,N_14883,N_11006);
xnor U18060 (N_18060,N_13890,N_14149);
nand U18061 (N_18061,N_13998,N_12367);
nand U18062 (N_18062,N_13732,N_13590);
or U18063 (N_18063,N_14716,N_10230);
xor U18064 (N_18064,N_14181,N_10532);
or U18065 (N_18065,N_11887,N_13036);
nand U18066 (N_18066,N_13853,N_14762);
nor U18067 (N_18067,N_11527,N_13661);
xor U18068 (N_18068,N_10216,N_11431);
xor U18069 (N_18069,N_11315,N_13879);
and U18070 (N_18070,N_11069,N_11273);
nand U18071 (N_18071,N_14101,N_12370);
nor U18072 (N_18072,N_11037,N_13150);
xnor U18073 (N_18073,N_10091,N_13621);
nand U18074 (N_18074,N_13360,N_11856);
nand U18075 (N_18075,N_10047,N_14077);
or U18076 (N_18076,N_10626,N_13852);
xnor U18077 (N_18077,N_12192,N_14926);
nor U18078 (N_18078,N_10260,N_10873);
and U18079 (N_18079,N_13438,N_12733);
xor U18080 (N_18080,N_10343,N_11548);
nand U18081 (N_18081,N_11611,N_13127);
and U18082 (N_18082,N_14783,N_14243);
and U18083 (N_18083,N_14905,N_13790);
and U18084 (N_18084,N_11386,N_12285);
xor U18085 (N_18085,N_12129,N_13730);
or U18086 (N_18086,N_11531,N_13664);
nand U18087 (N_18087,N_10394,N_13766);
and U18088 (N_18088,N_13979,N_11455);
nor U18089 (N_18089,N_14708,N_10177);
xor U18090 (N_18090,N_14494,N_12600);
nand U18091 (N_18091,N_11397,N_12864);
nor U18092 (N_18092,N_11826,N_13040);
and U18093 (N_18093,N_13507,N_13674);
and U18094 (N_18094,N_11024,N_14600);
xor U18095 (N_18095,N_10805,N_13636);
and U18096 (N_18096,N_11387,N_10120);
nor U18097 (N_18097,N_14915,N_14912);
xnor U18098 (N_18098,N_11252,N_10729);
and U18099 (N_18099,N_12971,N_12373);
nor U18100 (N_18100,N_14225,N_13695);
and U18101 (N_18101,N_14329,N_13334);
xnor U18102 (N_18102,N_12961,N_12453);
and U18103 (N_18103,N_13726,N_10442);
nand U18104 (N_18104,N_13982,N_10414);
or U18105 (N_18105,N_13601,N_14721);
nand U18106 (N_18106,N_10658,N_10920);
xnor U18107 (N_18107,N_13454,N_13287);
and U18108 (N_18108,N_12585,N_14702);
xor U18109 (N_18109,N_10093,N_10946);
and U18110 (N_18110,N_14883,N_13666);
or U18111 (N_18111,N_12872,N_11210);
nor U18112 (N_18112,N_12588,N_14481);
or U18113 (N_18113,N_11525,N_11037);
xnor U18114 (N_18114,N_14544,N_11646);
nor U18115 (N_18115,N_11629,N_11764);
xnor U18116 (N_18116,N_11712,N_10113);
nor U18117 (N_18117,N_14846,N_14185);
nor U18118 (N_18118,N_14750,N_12778);
or U18119 (N_18119,N_13072,N_11943);
xor U18120 (N_18120,N_13521,N_12868);
nor U18121 (N_18121,N_13465,N_11867);
nand U18122 (N_18122,N_13655,N_13626);
or U18123 (N_18123,N_13745,N_13918);
xnor U18124 (N_18124,N_13845,N_11885);
and U18125 (N_18125,N_10479,N_14170);
nor U18126 (N_18126,N_14014,N_13534);
nand U18127 (N_18127,N_10251,N_14699);
nor U18128 (N_18128,N_11812,N_13712);
nor U18129 (N_18129,N_10753,N_14521);
xnor U18130 (N_18130,N_14348,N_14170);
nand U18131 (N_18131,N_11143,N_14822);
and U18132 (N_18132,N_14592,N_11979);
or U18133 (N_18133,N_11733,N_14646);
xnor U18134 (N_18134,N_11999,N_13320);
and U18135 (N_18135,N_11411,N_14177);
xor U18136 (N_18136,N_11501,N_13914);
nand U18137 (N_18137,N_11556,N_13838);
nor U18138 (N_18138,N_13015,N_11000);
and U18139 (N_18139,N_14043,N_14069);
and U18140 (N_18140,N_10209,N_11800);
and U18141 (N_18141,N_13557,N_13192);
and U18142 (N_18142,N_13503,N_11074);
nand U18143 (N_18143,N_11815,N_10825);
and U18144 (N_18144,N_14078,N_13514);
nor U18145 (N_18145,N_11010,N_14521);
xnor U18146 (N_18146,N_12901,N_11831);
and U18147 (N_18147,N_10492,N_13226);
and U18148 (N_18148,N_11494,N_14488);
xnor U18149 (N_18149,N_13796,N_13406);
nand U18150 (N_18150,N_13023,N_11826);
nor U18151 (N_18151,N_14964,N_10129);
nor U18152 (N_18152,N_11759,N_10879);
and U18153 (N_18153,N_13148,N_11192);
or U18154 (N_18154,N_13624,N_11789);
nand U18155 (N_18155,N_14133,N_12906);
nand U18156 (N_18156,N_12146,N_11578);
and U18157 (N_18157,N_12043,N_12738);
nor U18158 (N_18158,N_14606,N_10323);
and U18159 (N_18159,N_13006,N_14096);
nor U18160 (N_18160,N_10061,N_12647);
nand U18161 (N_18161,N_10027,N_14779);
nand U18162 (N_18162,N_13988,N_13531);
nor U18163 (N_18163,N_14539,N_14770);
xor U18164 (N_18164,N_13457,N_12151);
nor U18165 (N_18165,N_10180,N_12446);
or U18166 (N_18166,N_13924,N_13316);
or U18167 (N_18167,N_14660,N_12561);
and U18168 (N_18168,N_12813,N_12067);
or U18169 (N_18169,N_14492,N_12353);
and U18170 (N_18170,N_14578,N_14985);
or U18171 (N_18171,N_10672,N_11672);
xor U18172 (N_18172,N_10078,N_13059);
xnor U18173 (N_18173,N_12007,N_14115);
nor U18174 (N_18174,N_10080,N_11732);
nand U18175 (N_18175,N_11184,N_10314);
nand U18176 (N_18176,N_13631,N_12783);
nand U18177 (N_18177,N_12229,N_14434);
nand U18178 (N_18178,N_13490,N_12899);
and U18179 (N_18179,N_13514,N_13102);
xor U18180 (N_18180,N_14477,N_13565);
nand U18181 (N_18181,N_12060,N_11507);
nor U18182 (N_18182,N_10146,N_12344);
or U18183 (N_18183,N_13684,N_14601);
nor U18184 (N_18184,N_14703,N_12604);
nor U18185 (N_18185,N_10960,N_13438);
nand U18186 (N_18186,N_13675,N_10702);
xnor U18187 (N_18187,N_11959,N_12317);
nand U18188 (N_18188,N_13752,N_13397);
nor U18189 (N_18189,N_11934,N_12132);
nand U18190 (N_18190,N_13984,N_14459);
or U18191 (N_18191,N_14902,N_11010);
nand U18192 (N_18192,N_10697,N_14602);
nor U18193 (N_18193,N_13160,N_11568);
or U18194 (N_18194,N_13676,N_13112);
nor U18195 (N_18195,N_14029,N_11610);
nand U18196 (N_18196,N_14612,N_13299);
or U18197 (N_18197,N_10305,N_12310);
nor U18198 (N_18198,N_13187,N_14443);
and U18199 (N_18199,N_12980,N_14568);
xnor U18200 (N_18200,N_13950,N_12849);
nor U18201 (N_18201,N_11904,N_10471);
nor U18202 (N_18202,N_11172,N_13340);
or U18203 (N_18203,N_13866,N_13878);
nand U18204 (N_18204,N_12326,N_12742);
xor U18205 (N_18205,N_13763,N_12561);
nand U18206 (N_18206,N_10273,N_10635);
and U18207 (N_18207,N_10658,N_14366);
nor U18208 (N_18208,N_10830,N_12036);
xor U18209 (N_18209,N_13330,N_14125);
xor U18210 (N_18210,N_10569,N_13271);
and U18211 (N_18211,N_14365,N_10226);
or U18212 (N_18212,N_10175,N_13589);
and U18213 (N_18213,N_10916,N_14564);
nand U18214 (N_18214,N_14445,N_11635);
and U18215 (N_18215,N_13353,N_11043);
xnor U18216 (N_18216,N_11732,N_11104);
nor U18217 (N_18217,N_11530,N_10491);
nor U18218 (N_18218,N_11186,N_14435);
nand U18219 (N_18219,N_10267,N_13508);
nand U18220 (N_18220,N_12881,N_14556);
xnor U18221 (N_18221,N_13318,N_11945);
and U18222 (N_18222,N_13169,N_10627);
and U18223 (N_18223,N_12538,N_14608);
nor U18224 (N_18224,N_13873,N_14380);
nand U18225 (N_18225,N_12867,N_14792);
or U18226 (N_18226,N_12743,N_10141);
nor U18227 (N_18227,N_12236,N_12904);
xor U18228 (N_18228,N_12469,N_14051);
and U18229 (N_18229,N_12227,N_10225);
nand U18230 (N_18230,N_14303,N_10202);
and U18231 (N_18231,N_12509,N_11224);
or U18232 (N_18232,N_12690,N_11080);
or U18233 (N_18233,N_12012,N_11143);
nor U18234 (N_18234,N_13161,N_12446);
nand U18235 (N_18235,N_14020,N_10454);
nand U18236 (N_18236,N_14960,N_10187);
nor U18237 (N_18237,N_13955,N_13347);
or U18238 (N_18238,N_11222,N_11237);
or U18239 (N_18239,N_13129,N_13664);
nand U18240 (N_18240,N_12809,N_12896);
or U18241 (N_18241,N_10082,N_13520);
or U18242 (N_18242,N_11187,N_14812);
or U18243 (N_18243,N_12304,N_14389);
nor U18244 (N_18244,N_13731,N_13561);
nor U18245 (N_18245,N_11584,N_10448);
nand U18246 (N_18246,N_11682,N_14431);
or U18247 (N_18247,N_10643,N_10086);
nand U18248 (N_18248,N_11067,N_14972);
nand U18249 (N_18249,N_13239,N_12233);
nand U18250 (N_18250,N_10030,N_12821);
nand U18251 (N_18251,N_13838,N_13285);
nand U18252 (N_18252,N_10869,N_12950);
nor U18253 (N_18253,N_13719,N_14469);
or U18254 (N_18254,N_13979,N_10515);
and U18255 (N_18255,N_14231,N_10307);
and U18256 (N_18256,N_13444,N_12816);
nand U18257 (N_18257,N_14448,N_14915);
and U18258 (N_18258,N_14561,N_13591);
or U18259 (N_18259,N_10745,N_11375);
and U18260 (N_18260,N_13670,N_13115);
xnor U18261 (N_18261,N_11344,N_14593);
or U18262 (N_18262,N_10977,N_13609);
or U18263 (N_18263,N_13041,N_13811);
nand U18264 (N_18264,N_10940,N_13896);
and U18265 (N_18265,N_14533,N_10424);
nand U18266 (N_18266,N_11635,N_10768);
or U18267 (N_18267,N_10912,N_10683);
xor U18268 (N_18268,N_14308,N_13762);
nand U18269 (N_18269,N_10465,N_10900);
nor U18270 (N_18270,N_11911,N_13869);
or U18271 (N_18271,N_14038,N_13575);
nand U18272 (N_18272,N_12335,N_14764);
xnor U18273 (N_18273,N_13785,N_11549);
nand U18274 (N_18274,N_10912,N_14262);
nor U18275 (N_18275,N_12902,N_11968);
nor U18276 (N_18276,N_11732,N_11207);
or U18277 (N_18277,N_12417,N_11950);
or U18278 (N_18278,N_12697,N_14884);
xor U18279 (N_18279,N_12311,N_11683);
and U18280 (N_18280,N_13576,N_14043);
xnor U18281 (N_18281,N_10878,N_11059);
or U18282 (N_18282,N_11310,N_13859);
and U18283 (N_18283,N_14797,N_14456);
xor U18284 (N_18284,N_11238,N_12871);
xnor U18285 (N_18285,N_12639,N_11688);
xnor U18286 (N_18286,N_11791,N_12438);
nor U18287 (N_18287,N_13376,N_12810);
and U18288 (N_18288,N_11290,N_14381);
xnor U18289 (N_18289,N_10707,N_13099);
nor U18290 (N_18290,N_10814,N_10882);
and U18291 (N_18291,N_12756,N_10613);
nor U18292 (N_18292,N_12916,N_11224);
or U18293 (N_18293,N_14293,N_10952);
or U18294 (N_18294,N_14971,N_14299);
xnor U18295 (N_18295,N_13892,N_10224);
xnor U18296 (N_18296,N_14596,N_13706);
xor U18297 (N_18297,N_14877,N_10509);
nand U18298 (N_18298,N_12147,N_13819);
and U18299 (N_18299,N_14520,N_11897);
nor U18300 (N_18300,N_13428,N_13733);
nand U18301 (N_18301,N_11719,N_14907);
and U18302 (N_18302,N_13419,N_10045);
or U18303 (N_18303,N_12455,N_14161);
or U18304 (N_18304,N_13853,N_11193);
nor U18305 (N_18305,N_14877,N_10776);
nor U18306 (N_18306,N_14576,N_12317);
nand U18307 (N_18307,N_12903,N_11705);
nand U18308 (N_18308,N_13799,N_12069);
and U18309 (N_18309,N_13077,N_11227);
nor U18310 (N_18310,N_11823,N_10070);
xnor U18311 (N_18311,N_14503,N_14209);
and U18312 (N_18312,N_11971,N_14380);
xor U18313 (N_18313,N_10697,N_11345);
xor U18314 (N_18314,N_10828,N_14617);
xor U18315 (N_18315,N_12696,N_13739);
nand U18316 (N_18316,N_11080,N_12467);
xnor U18317 (N_18317,N_12553,N_11404);
and U18318 (N_18318,N_12268,N_12856);
nor U18319 (N_18319,N_11373,N_11945);
xnor U18320 (N_18320,N_11458,N_14660);
xnor U18321 (N_18321,N_10282,N_12242);
xnor U18322 (N_18322,N_14082,N_12052);
or U18323 (N_18323,N_11076,N_14199);
nor U18324 (N_18324,N_12033,N_10129);
or U18325 (N_18325,N_13002,N_12442);
or U18326 (N_18326,N_11123,N_14955);
xnor U18327 (N_18327,N_12407,N_11890);
nand U18328 (N_18328,N_13783,N_10808);
and U18329 (N_18329,N_14807,N_14124);
or U18330 (N_18330,N_11857,N_13563);
nand U18331 (N_18331,N_10716,N_14128);
nor U18332 (N_18332,N_10112,N_12921);
nor U18333 (N_18333,N_10363,N_11515);
nand U18334 (N_18334,N_10584,N_13639);
and U18335 (N_18335,N_14623,N_10055);
nand U18336 (N_18336,N_13543,N_12834);
xnor U18337 (N_18337,N_14244,N_11872);
nor U18338 (N_18338,N_14240,N_10552);
and U18339 (N_18339,N_11343,N_14657);
nand U18340 (N_18340,N_13464,N_14365);
or U18341 (N_18341,N_10606,N_13828);
nand U18342 (N_18342,N_11080,N_11646);
xor U18343 (N_18343,N_13248,N_12971);
and U18344 (N_18344,N_12764,N_10455);
nand U18345 (N_18345,N_14552,N_10176);
nand U18346 (N_18346,N_10267,N_10649);
and U18347 (N_18347,N_13266,N_13518);
nand U18348 (N_18348,N_13555,N_11999);
nand U18349 (N_18349,N_14452,N_14042);
nand U18350 (N_18350,N_13910,N_13551);
xor U18351 (N_18351,N_12899,N_11634);
nand U18352 (N_18352,N_11449,N_12854);
xnor U18353 (N_18353,N_13707,N_10993);
xnor U18354 (N_18354,N_10807,N_12140);
xor U18355 (N_18355,N_13092,N_13177);
and U18356 (N_18356,N_13741,N_13168);
nand U18357 (N_18357,N_13395,N_12901);
nor U18358 (N_18358,N_14342,N_11693);
nor U18359 (N_18359,N_13325,N_11005);
and U18360 (N_18360,N_10615,N_12430);
xnor U18361 (N_18361,N_10721,N_13760);
or U18362 (N_18362,N_14962,N_10152);
nor U18363 (N_18363,N_10725,N_14336);
nand U18364 (N_18364,N_12336,N_11629);
or U18365 (N_18365,N_12496,N_13259);
xnor U18366 (N_18366,N_12954,N_11781);
xnor U18367 (N_18367,N_11760,N_11080);
nand U18368 (N_18368,N_11073,N_14121);
xor U18369 (N_18369,N_12502,N_11493);
and U18370 (N_18370,N_14221,N_14293);
and U18371 (N_18371,N_11759,N_11361);
xnor U18372 (N_18372,N_10920,N_10836);
or U18373 (N_18373,N_13662,N_12094);
nand U18374 (N_18374,N_10089,N_13018);
xor U18375 (N_18375,N_11078,N_12675);
or U18376 (N_18376,N_11986,N_13045);
xor U18377 (N_18377,N_13467,N_12224);
and U18378 (N_18378,N_12639,N_13722);
xnor U18379 (N_18379,N_13750,N_12331);
and U18380 (N_18380,N_14181,N_13277);
or U18381 (N_18381,N_14249,N_14001);
nor U18382 (N_18382,N_12563,N_14706);
xnor U18383 (N_18383,N_12252,N_10906);
and U18384 (N_18384,N_11758,N_13054);
and U18385 (N_18385,N_10860,N_11370);
and U18386 (N_18386,N_13440,N_12793);
and U18387 (N_18387,N_10365,N_10670);
nand U18388 (N_18388,N_10072,N_11517);
or U18389 (N_18389,N_11553,N_12440);
xnor U18390 (N_18390,N_10807,N_10292);
or U18391 (N_18391,N_11119,N_11466);
xnor U18392 (N_18392,N_13947,N_12602);
or U18393 (N_18393,N_12809,N_13917);
nor U18394 (N_18394,N_11451,N_10077);
nor U18395 (N_18395,N_13689,N_14019);
xor U18396 (N_18396,N_11295,N_13535);
and U18397 (N_18397,N_12686,N_11229);
and U18398 (N_18398,N_14835,N_11946);
xor U18399 (N_18399,N_11666,N_10927);
and U18400 (N_18400,N_13475,N_13676);
or U18401 (N_18401,N_14174,N_13051);
xor U18402 (N_18402,N_11923,N_11121);
and U18403 (N_18403,N_12106,N_14822);
xnor U18404 (N_18404,N_12193,N_12456);
nand U18405 (N_18405,N_11584,N_14623);
and U18406 (N_18406,N_12928,N_12985);
and U18407 (N_18407,N_13844,N_12917);
nand U18408 (N_18408,N_12168,N_11947);
xnor U18409 (N_18409,N_11435,N_13194);
xnor U18410 (N_18410,N_13349,N_10403);
nor U18411 (N_18411,N_14983,N_13760);
nand U18412 (N_18412,N_12043,N_11184);
xnor U18413 (N_18413,N_13621,N_13660);
xor U18414 (N_18414,N_13299,N_12396);
and U18415 (N_18415,N_10145,N_11715);
nor U18416 (N_18416,N_14305,N_10489);
nor U18417 (N_18417,N_10352,N_12095);
or U18418 (N_18418,N_13740,N_13399);
xor U18419 (N_18419,N_10351,N_13376);
and U18420 (N_18420,N_12373,N_14078);
nor U18421 (N_18421,N_12725,N_14859);
and U18422 (N_18422,N_13864,N_12093);
nand U18423 (N_18423,N_12211,N_14894);
and U18424 (N_18424,N_14741,N_11720);
and U18425 (N_18425,N_10801,N_10318);
nand U18426 (N_18426,N_12459,N_14229);
nand U18427 (N_18427,N_10565,N_13546);
and U18428 (N_18428,N_11349,N_11188);
and U18429 (N_18429,N_14495,N_10317);
nor U18430 (N_18430,N_11939,N_11043);
and U18431 (N_18431,N_10530,N_12408);
nand U18432 (N_18432,N_12353,N_11018);
or U18433 (N_18433,N_14706,N_14744);
nor U18434 (N_18434,N_10632,N_11662);
or U18435 (N_18435,N_12850,N_13956);
nor U18436 (N_18436,N_11546,N_13956);
xor U18437 (N_18437,N_12200,N_12229);
and U18438 (N_18438,N_13060,N_14364);
or U18439 (N_18439,N_11106,N_11519);
xnor U18440 (N_18440,N_10013,N_13784);
xor U18441 (N_18441,N_10648,N_11723);
nand U18442 (N_18442,N_13909,N_13170);
nor U18443 (N_18443,N_12058,N_12299);
or U18444 (N_18444,N_14187,N_14959);
nand U18445 (N_18445,N_12351,N_14712);
or U18446 (N_18446,N_12719,N_13948);
or U18447 (N_18447,N_13140,N_10358);
nor U18448 (N_18448,N_13409,N_13901);
or U18449 (N_18449,N_10232,N_14228);
and U18450 (N_18450,N_13520,N_11892);
xnor U18451 (N_18451,N_14013,N_11238);
xor U18452 (N_18452,N_11700,N_10106);
xnor U18453 (N_18453,N_11986,N_12450);
and U18454 (N_18454,N_14574,N_11987);
or U18455 (N_18455,N_13672,N_10889);
xnor U18456 (N_18456,N_12238,N_12499);
and U18457 (N_18457,N_12108,N_12150);
and U18458 (N_18458,N_11645,N_11215);
or U18459 (N_18459,N_11433,N_10751);
nand U18460 (N_18460,N_14297,N_13345);
nand U18461 (N_18461,N_11464,N_10470);
nand U18462 (N_18462,N_13686,N_13238);
or U18463 (N_18463,N_11919,N_12308);
nand U18464 (N_18464,N_14935,N_10745);
nor U18465 (N_18465,N_11721,N_11007);
xor U18466 (N_18466,N_13642,N_13420);
and U18467 (N_18467,N_12353,N_11197);
nor U18468 (N_18468,N_11249,N_14226);
xnor U18469 (N_18469,N_13131,N_11523);
nand U18470 (N_18470,N_12671,N_10427);
or U18471 (N_18471,N_10264,N_13452);
and U18472 (N_18472,N_14983,N_12612);
nand U18473 (N_18473,N_11011,N_11264);
xnor U18474 (N_18474,N_10335,N_14132);
nor U18475 (N_18475,N_14111,N_12606);
and U18476 (N_18476,N_12175,N_13730);
nand U18477 (N_18477,N_12234,N_10272);
or U18478 (N_18478,N_10631,N_13821);
or U18479 (N_18479,N_14387,N_13852);
xor U18480 (N_18480,N_14946,N_10844);
nor U18481 (N_18481,N_11993,N_12852);
or U18482 (N_18482,N_13100,N_10244);
nand U18483 (N_18483,N_11098,N_13242);
xor U18484 (N_18484,N_12648,N_10435);
nand U18485 (N_18485,N_11711,N_13843);
nor U18486 (N_18486,N_10704,N_11208);
xnor U18487 (N_18487,N_13334,N_14723);
nor U18488 (N_18488,N_11621,N_14480);
and U18489 (N_18489,N_11627,N_10410);
and U18490 (N_18490,N_11021,N_13139);
xor U18491 (N_18491,N_14129,N_10146);
and U18492 (N_18492,N_14206,N_14186);
or U18493 (N_18493,N_11981,N_14814);
nand U18494 (N_18494,N_11231,N_12689);
nand U18495 (N_18495,N_12680,N_10535);
nand U18496 (N_18496,N_12264,N_14012);
nand U18497 (N_18497,N_12015,N_12409);
nor U18498 (N_18498,N_10982,N_14004);
or U18499 (N_18499,N_11667,N_14512);
nand U18500 (N_18500,N_12489,N_10019);
nand U18501 (N_18501,N_13189,N_12320);
and U18502 (N_18502,N_11618,N_12768);
xor U18503 (N_18503,N_10694,N_13327);
and U18504 (N_18504,N_13270,N_11310);
xnor U18505 (N_18505,N_11425,N_11576);
and U18506 (N_18506,N_12725,N_14460);
or U18507 (N_18507,N_14298,N_13862);
nor U18508 (N_18508,N_14875,N_11118);
nand U18509 (N_18509,N_10936,N_11229);
nand U18510 (N_18510,N_12453,N_12236);
nand U18511 (N_18511,N_12697,N_11298);
nor U18512 (N_18512,N_10146,N_10424);
or U18513 (N_18513,N_12813,N_12502);
or U18514 (N_18514,N_12628,N_14932);
nor U18515 (N_18515,N_12517,N_14987);
and U18516 (N_18516,N_10413,N_13937);
and U18517 (N_18517,N_11168,N_11620);
or U18518 (N_18518,N_14333,N_10746);
and U18519 (N_18519,N_14975,N_12842);
or U18520 (N_18520,N_10449,N_14109);
and U18521 (N_18521,N_13847,N_11093);
xor U18522 (N_18522,N_13068,N_11337);
nor U18523 (N_18523,N_12016,N_14754);
and U18524 (N_18524,N_14571,N_12585);
and U18525 (N_18525,N_14776,N_12378);
and U18526 (N_18526,N_14704,N_12818);
or U18527 (N_18527,N_14581,N_14970);
or U18528 (N_18528,N_14733,N_11174);
and U18529 (N_18529,N_13456,N_11366);
xnor U18530 (N_18530,N_11612,N_10096);
nor U18531 (N_18531,N_10814,N_11306);
and U18532 (N_18532,N_14707,N_13590);
nand U18533 (N_18533,N_10813,N_12186);
and U18534 (N_18534,N_14799,N_11954);
xor U18535 (N_18535,N_13602,N_10841);
nor U18536 (N_18536,N_13089,N_12056);
nor U18537 (N_18537,N_11727,N_11486);
or U18538 (N_18538,N_14388,N_13535);
xnor U18539 (N_18539,N_13742,N_13940);
and U18540 (N_18540,N_11516,N_11635);
nor U18541 (N_18541,N_14110,N_12969);
or U18542 (N_18542,N_14625,N_13289);
and U18543 (N_18543,N_13099,N_10444);
xor U18544 (N_18544,N_14919,N_10110);
or U18545 (N_18545,N_12987,N_14274);
xor U18546 (N_18546,N_13027,N_12493);
nand U18547 (N_18547,N_12074,N_13398);
xnor U18548 (N_18548,N_11891,N_13903);
and U18549 (N_18549,N_13311,N_14183);
nand U18550 (N_18550,N_10602,N_12745);
or U18551 (N_18551,N_11834,N_12351);
or U18552 (N_18552,N_14684,N_10800);
and U18553 (N_18553,N_12585,N_10111);
xor U18554 (N_18554,N_13751,N_10633);
nand U18555 (N_18555,N_12322,N_11597);
or U18556 (N_18556,N_13014,N_14703);
xnor U18557 (N_18557,N_13665,N_10621);
nand U18558 (N_18558,N_10046,N_14276);
or U18559 (N_18559,N_12012,N_11828);
nand U18560 (N_18560,N_13790,N_14678);
nand U18561 (N_18561,N_14670,N_11456);
nor U18562 (N_18562,N_10489,N_11509);
nor U18563 (N_18563,N_13744,N_10229);
xnor U18564 (N_18564,N_11013,N_12656);
nor U18565 (N_18565,N_11793,N_10525);
and U18566 (N_18566,N_10959,N_10763);
nor U18567 (N_18567,N_10226,N_12844);
nor U18568 (N_18568,N_14411,N_12414);
nor U18569 (N_18569,N_12484,N_10934);
xnor U18570 (N_18570,N_13986,N_14111);
nand U18571 (N_18571,N_14145,N_12784);
and U18572 (N_18572,N_12513,N_12184);
xor U18573 (N_18573,N_11574,N_14812);
or U18574 (N_18574,N_11630,N_10682);
and U18575 (N_18575,N_12167,N_14511);
nand U18576 (N_18576,N_11503,N_14786);
nor U18577 (N_18577,N_14596,N_13476);
nand U18578 (N_18578,N_12410,N_11038);
nor U18579 (N_18579,N_12769,N_13109);
nand U18580 (N_18580,N_11507,N_12850);
xnor U18581 (N_18581,N_13392,N_14231);
nor U18582 (N_18582,N_13612,N_12087);
xnor U18583 (N_18583,N_11280,N_12458);
nor U18584 (N_18584,N_13490,N_11832);
and U18585 (N_18585,N_12360,N_13937);
nand U18586 (N_18586,N_11561,N_10167);
xor U18587 (N_18587,N_11383,N_13217);
or U18588 (N_18588,N_11289,N_14385);
xnor U18589 (N_18589,N_11214,N_10977);
or U18590 (N_18590,N_14794,N_11886);
xnor U18591 (N_18591,N_11869,N_10733);
and U18592 (N_18592,N_11033,N_12737);
or U18593 (N_18593,N_10854,N_13785);
and U18594 (N_18594,N_12885,N_13403);
nand U18595 (N_18595,N_14538,N_11840);
xor U18596 (N_18596,N_14229,N_14572);
and U18597 (N_18597,N_14848,N_14425);
nor U18598 (N_18598,N_11205,N_12116);
nand U18599 (N_18599,N_14151,N_10832);
nand U18600 (N_18600,N_12711,N_13498);
or U18601 (N_18601,N_12805,N_12919);
or U18602 (N_18602,N_12933,N_11041);
and U18603 (N_18603,N_14126,N_14154);
and U18604 (N_18604,N_10759,N_12598);
or U18605 (N_18605,N_13236,N_12515);
xnor U18606 (N_18606,N_13435,N_11780);
nand U18607 (N_18607,N_14384,N_11525);
and U18608 (N_18608,N_10704,N_13946);
xnor U18609 (N_18609,N_12761,N_11360);
and U18610 (N_18610,N_13523,N_11780);
and U18611 (N_18611,N_14856,N_14142);
and U18612 (N_18612,N_10158,N_14821);
nand U18613 (N_18613,N_11775,N_11246);
or U18614 (N_18614,N_10420,N_14057);
nor U18615 (N_18615,N_14600,N_12737);
or U18616 (N_18616,N_13473,N_13523);
nor U18617 (N_18617,N_12217,N_11674);
or U18618 (N_18618,N_11451,N_12881);
xnor U18619 (N_18619,N_12882,N_13155);
or U18620 (N_18620,N_14478,N_12804);
nor U18621 (N_18621,N_12168,N_10221);
or U18622 (N_18622,N_13928,N_11712);
nand U18623 (N_18623,N_13518,N_12113);
nand U18624 (N_18624,N_12314,N_14951);
xnor U18625 (N_18625,N_11712,N_11264);
nand U18626 (N_18626,N_13008,N_11577);
and U18627 (N_18627,N_12835,N_10320);
or U18628 (N_18628,N_11114,N_12515);
xor U18629 (N_18629,N_11815,N_13915);
xor U18630 (N_18630,N_14822,N_11005);
and U18631 (N_18631,N_10802,N_12531);
nor U18632 (N_18632,N_14042,N_13831);
nand U18633 (N_18633,N_12092,N_10481);
xnor U18634 (N_18634,N_12634,N_10701);
nor U18635 (N_18635,N_10445,N_10365);
or U18636 (N_18636,N_12237,N_11638);
nor U18637 (N_18637,N_12600,N_12605);
nor U18638 (N_18638,N_14937,N_14172);
xor U18639 (N_18639,N_14625,N_13544);
nor U18640 (N_18640,N_11428,N_13079);
and U18641 (N_18641,N_12399,N_14546);
nand U18642 (N_18642,N_13272,N_14921);
xor U18643 (N_18643,N_11337,N_14953);
and U18644 (N_18644,N_14359,N_12184);
nor U18645 (N_18645,N_12301,N_12529);
xnor U18646 (N_18646,N_10452,N_10555);
nand U18647 (N_18647,N_10745,N_11249);
or U18648 (N_18648,N_10002,N_10677);
and U18649 (N_18649,N_13165,N_13564);
or U18650 (N_18650,N_14641,N_13779);
or U18651 (N_18651,N_12553,N_10210);
and U18652 (N_18652,N_12709,N_10304);
and U18653 (N_18653,N_13621,N_11265);
nor U18654 (N_18654,N_11674,N_12038);
nor U18655 (N_18655,N_11913,N_13570);
nand U18656 (N_18656,N_12935,N_13388);
and U18657 (N_18657,N_11444,N_14266);
nand U18658 (N_18658,N_11381,N_13365);
nand U18659 (N_18659,N_12784,N_11946);
xnor U18660 (N_18660,N_10052,N_12543);
xnor U18661 (N_18661,N_10525,N_13637);
nand U18662 (N_18662,N_11747,N_10570);
xor U18663 (N_18663,N_13584,N_11292);
xnor U18664 (N_18664,N_10571,N_14136);
and U18665 (N_18665,N_11591,N_13743);
nand U18666 (N_18666,N_14271,N_11143);
nor U18667 (N_18667,N_11051,N_12222);
nor U18668 (N_18668,N_10593,N_10559);
or U18669 (N_18669,N_13344,N_14888);
or U18670 (N_18670,N_11026,N_10336);
and U18671 (N_18671,N_10746,N_13043);
nor U18672 (N_18672,N_11531,N_12521);
and U18673 (N_18673,N_13389,N_10697);
xor U18674 (N_18674,N_14755,N_12575);
and U18675 (N_18675,N_13678,N_13202);
or U18676 (N_18676,N_13724,N_11608);
nand U18677 (N_18677,N_12252,N_12601);
nand U18678 (N_18678,N_11708,N_14149);
xor U18679 (N_18679,N_13877,N_12445);
or U18680 (N_18680,N_13001,N_11372);
nor U18681 (N_18681,N_12255,N_11071);
nand U18682 (N_18682,N_14143,N_10433);
and U18683 (N_18683,N_13826,N_13806);
nor U18684 (N_18684,N_10863,N_14280);
or U18685 (N_18685,N_11753,N_10571);
or U18686 (N_18686,N_10512,N_14932);
xor U18687 (N_18687,N_12460,N_14144);
xnor U18688 (N_18688,N_14659,N_12282);
or U18689 (N_18689,N_10456,N_14347);
or U18690 (N_18690,N_11139,N_13225);
or U18691 (N_18691,N_10348,N_13382);
xor U18692 (N_18692,N_11009,N_14877);
nor U18693 (N_18693,N_12233,N_14552);
nand U18694 (N_18694,N_13727,N_14954);
nand U18695 (N_18695,N_10605,N_10547);
nor U18696 (N_18696,N_11831,N_11587);
xor U18697 (N_18697,N_10842,N_14111);
xor U18698 (N_18698,N_12169,N_10836);
nand U18699 (N_18699,N_12003,N_12697);
or U18700 (N_18700,N_13533,N_14554);
nor U18701 (N_18701,N_13469,N_14723);
nand U18702 (N_18702,N_12136,N_14890);
nand U18703 (N_18703,N_12888,N_12648);
and U18704 (N_18704,N_10011,N_12241);
and U18705 (N_18705,N_10815,N_14377);
and U18706 (N_18706,N_12311,N_12899);
xor U18707 (N_18707,N_11571,N_14380);
xnor U18708 (N_18708,N_10048,N_14750);
xnor U18709 (N_18709,N_12790,N_13543);
nand U18710 (N_18710,N_11369,N_10533);
nand U18711 (N_18711,N_10443,N_14787);
nand U18712 (N_18712,N_10225,N_14775);
or U18713 (N_18713,N_10221,N_13161);
or U18714 (N_18714,N_14091,N_10056);
nand U18715 (N_18715,N_14958,N_11222);
nand U18716 (N_18716,N_10678,N_10335);
and U18717 (N_18717,N_13841,N_13967);
xnor U18718 (N_18718,N_13324,N_13890);
nor U18719 (N_18719,N_10785,N_13545);
xor U18720 (N_18720,N_10762,N_11096);
or U18721 (N_18721,N_14709,N_12578);
xor U18722 (N_18722,N_14880,N_12177);
xor U18723 (N_18723,N_14632,N_11322);
nor U18724 (N_18724,N_10226,N_12750);
nand U18725 (N_18725,N_12905,N_10053);
and U18726 (N_18726,N_14824,N_14649);
nand U18727 (N_18727,N_11876,N_14963);
nor U18728 (N_18728,N_14784,N_14997);
or U18729 (N_18729,N_12690,N_14012);
xor U18730 (N_18730,N_11207,N_13887);
xor U18731 (N_18731,N_10512,N_12326);
nor U18732 (N_18732,N_13176,N_12407);
or U18733 (N_18733,N_11618,N_11397);
xnor U18734 (N_18734,N_14848,N_11488);
nand U18735 (N_18735,N_11332,N_10972);
and U18736 (N_18736,N_11933,N_14489);
nand U18737 (N_18737,N_11131,N_12020);
nand U18738 (N_18738,N_13446,N_11233);
xor U18739 (N_18739,N_12352,N_11945);
or U18740 (N_18740,N_12867,N_12344);
nand U18741 (N_18741,N_14739,N_12344);
nor U18742 (N_18742,N_11651,N_13787);
or U18743 (N_18743,N_12976,N_14009);
nor U18744 (N_18744,N_12936,N_11305);
nand U18745 (N_18745,N_14475,N_10192);
and U18746 (N_18746,N_10553,N_11873);
nand U18747 (N_18747,N_11541,N_14932);
and U18748 (N_18748,N_12954,N_14808);
and U18749 (N_18749,N_12944,N_11157);
nor U18750 (N_18750,N_11250,N_14812);
nor U18751 (N_18751,N_12219,N_12211);
xor U18752 (N_18752,N_12956,N_11935);
and U18753 (N_18753,N_12058,N_14315);
and U18754 (N_18754,N_12302,N_10828);
or U18755 (N_18755,N_11520,N_11658);
or U18756 (N_18756,N_11616,N_10795);
or U18757 (N_18757,N_10092,N_12954);
or U18758 (N_18758,N_13317,N_13619);
xnor U18759 (N_18759,N_12276,N_11288);
nor U18760 (N_18760,N_12859,N_12813);
nor U18761 (N_18761,N_12462,N_12817);
xnor U18762 (N_18762,N_12862,N_13820);
nand U18763 (N_18763,N_10735,N_13856);
nand U18764 (N_18764,N_12095,N_13135);
nand U18765 (N_18765,N_13208,N_14304);
and U18766 (N_18766,N_10992,N_12496);
nand U18767 (N_18767,N_11569,N_13124);
nand U18768 (N_18768,N_13883,N_13174);
xor U18769 (N_18769,N_11470,N_10306);
nor U18770 (N_18770,N_13754,N_12623);
and U18771 (N_18771,N_13611,N_11398);
nand U18772 (N_18772,N_11933,N_11245);
nand U18773 (N_18773,N_11626,N_10025);
xor U18774 (N_18774,N_11087,N_11158);
xnor U18775 (N_18775,N_14054,N_12063);
xor U18776 (N_18776,N_12713,N_10538);
nand U18777 (N_18777,N_14002,N_12215);
nand U18778 (N_18778,N_13779,N_10402);
and U18779 (N_18779,N_11015,N_10601);
or U18780 (N_18780,N_10354,N_13879);
nor U18781 (N_18781,N_12321,N_10493);
and U18782 (N_18782,N_14224,N_14751);
and U18783 (N_18783,N_14496,N_12939);
nand U18784 (N_18784,N_12336,N_11786);
and U18785 (N_18785,N_14018,N_14057);
nand U18786 (N_18786,N_14555,N_10930);
nand U18787 (N_18787,N_12492,N_11152);
xnor U18788 (N_18788,N_12158,N_11266);
xnor U18789 (N_18789,N_12887,N_11555);
and U18790 (N_18790,N_13842,N_10179);
nor U18791 (N_18791,N_12169,N_13400);
and U18792 (N_18792,N_10178,N_13929);
nor U18793 (N_18793,N_12503,N_11735);
xnor U18794 (N_18794,N_10312,N_13297);
and U18795 (N_18795,N_12114,N_11413);
xor U18796 (N_18796,N_14338,N_10172);
nand U18797 (N_18797,N_14056,N_11266);
and U18798 (N_18798,N_13434,N_11018);
nand U18799 (N_18799,N_12365,N_10915);
or U18800 (N_18800,N_12985,N_10834);
nor U18801 (N_18801,N_10899,N_12334);
or U18802 (N_18802,N_10718,N_12221);
nor U18803 (N_18803,N_13506,N_14015);
or U18804 (N_18804,N_11457,N_12519);
nor U18805 (N_18805,N_10405,N_10640);
xnor U18806 (N_18806,N_11680,N_12804);
or U18807 (N_18807,N_13128,N_13059);
xnor U18808 (N_18808,N_11674,N_11812);
or U18809 (N_18809,N_13587,N_14106);
nand U18810 (N_18810,N_14206,N_10725);
or U18811 (N_18811,N_10040,N_10986);
xor U18812 (N_18812,N_11762,N_13332);
or U18813 (N_18813,N_11998,N_13138);
or U18814 (N_18814,N_10644,N_14937);
nand U18815 (N_18815,N_12731,N_14018);
nand U18816 (N_18816,N_10638,N_14804);
xor U18817 (N_18817,N_12633,N_11746);
xor U18818 (N_18818,N_12154,N_13210);
nand U18819 (N_18819,N_14919,N_14962);
or U18820 (N_18820,N_12954,N_13125);
xor U18821 (N_18821,N_13930,N_10950);
nor U18822 (N_18822,N_10115,N_13836);
nor U18823 (N_18823,N_10460,N_12092);
xnor U18824 (N_18824,N_10817,N_13624);
nand U18825 (N_18825,N_10227,N_11710);
and U18826 (N_18826,N_12986,N_14371);
nor U18827 (N_18827,N_11816,N_14267);
or U18828 (N_18828,N_12065,N_11071);
or U18829 (N_18829,N_12091,N_12389);
xor U18830 (N_18830,N_10136,N_11211);
and U18831 (N_18831,N_13862,N_10019);
and U18832 (N_18832,N_12906,N_10853);
nor U18833 (N_18833,N_11518,N_13274);
nor U18834 (N_18834,N_13012,N_14941);
xor U18835 (N_18835,N_10427,N_12408);
and U18836 (N_18836,N_13511,N_11145);
nand U18837 (N_18837,N_10046,N_12141);
nand U18838 (N_18838,N_10228,N_12720);
xnor U18839 (N_18839,N_11095,N_11845);
or U18840 (N_18840,N_14347,N_14463);
nand U18841 (N_18841,N_12365,N_12238);
xnor U18842 (N_18842,N_12838,N_14663);
nor U18843 (N_18843,N_11084,N_14502);
xnor U18844 (N_18844,N_12542,N_13116);
nand U18845 (N_18845,N_10280,N_14137);
and U18846 (N_18846,N_14628,N_10913);
nor U18847 (N_18847,N_12332,N_10446);
or U18848 (N_18848,N_14447,N_12621);
nor U18849 (N_18849,N_14003,N_14170);
or U18850 (N_18850,N_14460,N_10417);
nand U18851 (N_18851,N_10410,N_10433);
nor U18852 (N_18852,N_10835,N_11791);
and U18853 (N_18853,N_13273,N_12775);
nor U18854 (N_18854,N_11180,N_14535);
xnor U18855 (N_18855,N_14621,N_13627);
or U18856 (N_18856,N_13988,N_11359);
or U18857 (N_18857,N_11114,N_12032);
nor U18858 (N_18858,N_14143,N_10566);
nand U18859 (N_18859,N_10545,N_13035);
nand U18860 (N_18860,N_11699,N_11307);
xor U18861 (N_18861,N_10150,N_13801);
or U18862 (N_18862,N_11599,N_13070);
nand U18863 (N_18863,N_11341,N_10734);
nor U18864 (N_18864,N_14171,N_12937);
nor U18865 (N_18865,N_13701,N_12662);
nor U18866 (N_18866,N_11311,N_13922);
and U18867 (N_18867,N_10879,N_11335);
and U18868 (N_18868,N_11215,N_14143);
or U18869 (N_18869,N_12067,N_10389);
and U18870 (N_18870,N_12556,N_11362);
and U18871 (N_18871,N_11258,N_14005);
xnor U18872 (N_18872,N_14073,N_10069);
or U18873 (N_18873,N_13260,N_13427);
xnor U18874 (N_18874,N_10349,N_10968);
xor U18875 (N_18875,N_10142,N_11488);
nand U18876 (N_18876,N_13388,N_14610);
or U18877 (N_18877,N_11312,N_12542);
or U18878 (N_18878,N_14338,N_11055);
xor U18879 (N_18879,N_12311,N_13581);
xor U18880 (N_18880,N_11157,N_14920);
nor U18881 (N_18881,N_14391,N_14101);
and U18882 (N_18882,N_14369,N_12808);
nor U18883 (N_18883,N_12370,N_10092);
and U18884 (N_18884,N_12994,N_10954);
and U18885 (N_18885,N_13775,N_13353);
nor U18886 (N_18886,N_14254,N_14791);
or U18887 (N_18887,N_13734,N_13918);
or U18888 (N_18888,N_10995,N_11473);
or U18889 (N_18889,N_11850,N_14624);
xnor U18890 (N_18890,N_12872,N_14838);
nor U18891 (N_18891,N_11798,N_11632);
xnor U18892 (N_18892,N_12206,N_13337);
or U18893 (N_18893,N_10271,N_11349);
xnor U18894 (N_18894,N_12720,N_13321);
and U18895 (N_18895,N_13437,N_14478);
nand U18896 (N_18896,N_11685,N_13498);
nor U18897 (N_18897,N_14850,N_11404);
nor U18898 (N_18898,N_12367,N_10427);
nand U18899 (N_18899,N_13570,N_10438);
or U18900 (N_18900,N_13880,N_12182);
and U18901 (N_18901,N_13583,N_11601);
and U18902 (N_18902,N_14175,N_12107);
or U18903 (N_18903,N_14098,N_14126);
and U18904 (N_18904,N_10975,N_14026);
xor U18905 (N_18905,N_10018,N_11541);
and U18906 (N_18906,N_12815,N_11721);
and U18907 (N_18907,N_13854,N_13002);
or U18908 (N_18908,N_10472,N_14845);
and U18909 (N_18909,N_13027,N_13994);
and U18910 (N_18910,N_10443,N_11103);
or U18911 (N_18911,N_14664,N_11457);
nand U18912 (N_18912,N_14417,N_10281);
xnor U18913 (N_18913,N_13511,N_12947);
or U18914 (N_18914,N_14639,N_11347);
nor U18915 (N_18915,N_11980,N_12822);
xnor U18916 (N_18916,N_14596,N_13524);
and U18917 (N_18917,N_14882,N_12879);
and U18918 (N_18918,N_11407,N_14362);
xnor U18919 (N_18919,N_13034,N_12442);
and U18920 (N_18920,N_14798,N_13818);
or U18921 (N_18921,N_11807,N_14172);
xnor U18922 (N_18922,N_14001,N_10874);
and U18923 (N_18923,N_14679,N_13319);
and U18924 (N_18924,N_13301,N_14560);
xnor U18925 (N_18925,N_13736,N_11875);
or U18926 (N_18926,N_11727,N_12028);
or U18927 (N_18927,N_11634,N_12669);
nor U18928 (N_18928,N_12047,N_10751);
and U18929 (N_18929,N_10697,N_12265);
xor U18930 (N_18930,N_14717,N_13704);
or U18931 (N_18931,N_12927,N_14623);
nand U18932 (N_18932,N_12859,N_14218);
or U18933 (N_18933,N_14460,N_11326);
nor U18934 (N_18934,N_12241,N_12861);
nand U18935 (N_18935,N_14284,N_10727);
xnor U18936 (N_18936,N_13261,N_10194);
xnor U18937 (N_18937,N_12645,N_12113);
nor U18938 (N_18938,N_12859,N_14663);
and U18939 (N_18939,N_10063,N_13919);
and U18940 (N_18940,N_10107,N_14581);
nand U18941 (N_18941,N_14894,N_13578);
nand U18942 (N_18942,N_11900,N_14132);
nor U18943 (N_18943,N_14958,N_10816);
nor U18944 (N_18944,N_14699,N_11230);
xor U18945 (N_18945,N_14310,N_12343);
xnor U18946 (N_18946,N_11718,N_13098);
and U18947 (N_18947,N_11862,N_12869);
or U18948 (N_18948,N_13775,N_11642);
nand U18949 (N_18949,N_14778,N_10613);
and U18950 (N_18950,N_11485,N_13018);
nand U18951 (N_18951,N_13579,N_14080);
nor U18952 (N_18952,N_14115,N_10591);
nor U18953 (N_18953,N_10490,N_12897);
xnor U18954 (N_18954,N_12464,N_10792);
nor U18955 (N_18955,N_10238,N_13866);
or U18956 (N_18956,N_14609,N_10062);
nand U18957 (N_18957,N_13956,N_10876);
and U18958 (N_18958,N_11673,N_11751);
nand U18959 (N_18959,N_10967,N_12692);
nand U18960 (N_18960,N_11739,N_11954);
nor U18961 (N_18961,N_12519,N_14577);
nor U18962 (N_18962,N_14379,N_14468);
xnor U18963 (N_18963,N_11304,N_12050);
nand U18964 (N_18964,N_11373,N_14794);
or U18965 (N_18965,N_10084,N_10574);
xnor U18966 (N_18966,N_10560,N_11033);
xnor U18967 (N_18967,N_14023,N_10098);
nand U18968 (N_18968,N_12870,N_12644);
nand U18969 (N_18969,N_14192,N_10689);
and U18970 (N_18970,N_13796,N_10053);
xnor U18971 (N_18971,N_11095,N_10688);
nand U18972 (N_18972,N_13241,N_12940);
nor U18973 (N_18973,N_12916,N_13441);
nand U18974 (N_18974,N_11023,N_14322);
nor U18975 (N_18975,N_10459,N_13304);
and U18976 (N_18976,N_10738,N_14080);
xnor U18977 (N_18977,N_10986,N_10353);
xnor U18978 (N_18978,N_14558,N_12291);
nand U18979 (N_18979,N_14777,N_12597);
and U18980 (N_18980,N_11263,N_14308);
and U18981 (N_18981,N_12754,N_12724);
nand U18982 (N_18982,N_14326,N_13277);
xor U18983 (N_18983,N_12431,N_12252);
and U18984 (N_18984,N_11127,N_11738);
or U18985 (N_18985,N_12110,N_12864);
or U18986 (N_18986,N_11991,N_12825);
or U18987 (N_18987,N_10372,N_10939);
or U18988 (N_18988,N_12834,N_14362);
nor U18989 (N_18989,N_13155,N_11610);
or U18990 (N_18990,N_14046,N_14598);
or U18991 (N_18991,N_11906,N_12946);
nor U18992 (N_18992,N_14855,N_13162);
or U18993 (N_18993,N_13682,N_10449);
and U18994 (N_18994,N_12731,N_14566);
or U18995 (N_18995,N_14168,N_11957);
xnor U18996 (N_18996,N_12986,N_12782);
xnor U18997 (N_18997,N_12016,N_12838);
and U18998 (N_18998,N_12283,N_11484);
or U18999 (N_18999,N_13901,N_11477);
or U19000 (N_19000,N_12401,N_14116);
and U19001 (N_19001,N_10897,N_10357);
nor U19002 (N_19002,N_14126,N_11568);
or U19003 (N_19003,N_11563,N_14157);
nand U19004 (N_19004,N_12220,N_11275);
or U19005 (N_19005,N_14114,N_11272);
nor U19006 (N_19006,N_10057,N_14927);
nand U19007 (N_19007,N_10193,N_14077);
nand U19008 (N_19008,N_14840,N_11424);
and U19009 (N_19009,N_14753,N_12051);
or U19010 (N_19010,N_14284,N_11778);
nor U19011 (N_19011,N_12617,N_13916);
nand U19012 (N_19012,N_14090,N_13607);
or U19013 (N_19013,N_14439,N_14009);
nand U19014 (N_19014,N_14234,N_12623);
nand U19015 (N_19015,N_10268,N_13978);
xnor U19016 (N_19016,N_13496,N_12537);
nand U19017 (N_19017,N_10850,N_12415);
nor U19018 (N_19018,N_13793,N_12177);
nor U19019 (N_19019,N_12522,N_11016);
nand U19020 (N_19020,N_10623,N_11741);
nand U19021 (N_19021,N_10267,N_14461);
or U19022 (N_19022,N_13154,N_13238);
nor U19023 (N_19023,N_13226,N_11723);
and U19024 (N_19024,N_12931,N_12977);
xor U19025 (N_19025,N_12894,N_12739);
xor U19026 (N_19026,N_11301,N_12153);
nand U19027 (N_19027,N_12262,N_14500);
xor U19028 (N_19028,N_11753,N_13395);
and U19029 (N_19029,N_14396,N_11523);
and U19030 (N_19030,N_10606,N_13510);
or U19031 (N_19031,N_13409,N_14112);
and U19032 (N_19032,N_14202,N_11595);
and U19033 (N_19033,N_13733,N_11230);
xor U19034 (N_19034,N_13957,N_12876);
nand U19035 (N_19035,N_14882,N_10601);
nor U19036 (N_19036,N_11678,N_11045);
or U19037 (N_19037,N_14490,N_14063);
and U19038 (N_19038,N_14458,N_13348);
xnor U19039 (N_19039,N_10429,N_13144);
or U19040 (N_19040,N_12190,N_14340);
nand U19041 (N_19041,N_10195,N_12245);
xnor U19042 (N_19042,N_11405,N_12221);
xnor U19043 (N_19043,N_13537,N_11706);
nor U19044 (N_19044,N_14446,N_10745);
nor U19045 (N_19045,N_14822,N_11765);
nand U19046 (N_19046,N_11041,N_10167);
and U19047 (N_19047,N_11079,N_14137);
nor U19048 (N_19048,N_14217,N_13343);
and U19049 (N_19049,N_13024,N_11343);
nor U19050 (N_19050,N_10877,N_10076);
and U19051 (N_19051,N_13231,N_14747);
nand U19052 (N_19052,N_10993,N_10924);
and U19053 (N_19053,N_10220,N_11959);
xor U19054 (N_19054,N_11811,N_10294);
nor U19055 (N_19055,N_12565,N_12745);
or U19056 (N_19056,N_10349,N_11884);
or U19057 (N_19057,N_13553,N_11073);
or U19058 (N_19058,N_11167,N_11556);
nor U19059 (N_19059,N_11626,N_13403);
or U19060 (N_19060,N_10979,N_13834);
nand U19061 (N_19061,N_11196,N_10885);
or U19062 (N_19062,N_14279,N_10353);
and U19063 (N_19063,N_12927,N_14531);
or U19064 (N_19064,N_12743,N_10157);
xor U19065 (N_19065,N_12743,N_10379);
and U19066 (N_19066,N_13516,N_14999);
nand U19067 (N_19067,N_12965,N_14802);
or U19068 (N_19068,N_12640,N_14729);
and U19069 (N_19069,N_13701,N_11669);
xor U19070 (N_19070,N_10291,N_12990);
nand U19071 (N_19071,N_11719,N_12608);
and U19072 (N_19072,N_10608,N_10379);
nand U19073 (N_19073,N_12246,N_14790);
and U19074 (N_19074,N_11633,N_12897);
nand U19075 (N_19075,N_13951,N_14182);
xor U19076 (N_19076,N_14573,N_14868);
or U19077 (N_19077,N_12372,N_12413);
nand U19078 (N_19078,N_13649,N_11979);
nor U19079 (N_19079,N_14030,N_13973);
or U19080 (N_19080,N_10268,N_13210);
nor U19081 (N_19081,N_10698,N_12667);
and U19082 (N_19082,N_10055,N_12349);
xnor U19083 (N_19083,N_11972,N_14641);
and U19084 (N_19084,N_10052,N_12188);
or U19085 (N_19085,N_10814,N_11386);
or U19086 (N_19086,N_10613,N_11683);
and U19087 (N_19087,N_13939,N_14569);
or U19088 (N_19088,N_13644,N_10313);
nor U19089 (N_19089,N_11439,N_14175);
xor U19090 (N_19090,N_14710,N_13633);
and U19091 (N_19091,N_14075,N_12134);
xor U19092 (N_19092,N_12842,N_14517);
or U19093 (N_19093,N_11781,N_11968);
and U19094 (N_19094,N_12431,N_11481);
xnor U19095 (N_19095,N_14491,N_12772);
nor U19096 (N_19096,N_12129,N_12814);
nand U19097 (N_19097,N_10711,N_12592);
nor U19098 (N_19098,N_10147,N_11357);
nand U19099 (N_19099,N_12476,N_13358);
or U19100 (N_19100,N_11432,N_11891);
and U19101 (N_19101,N_13335,N_10724);
nand U19102 (N_19102,N_13077,N_14713);
nand U19103 (N_19103,N_10568,N_14807);
xnor U19104 (N_19104,N_13401,N_14030);
nand U19105 (N_19105,N_10493,N_11709);
or U19106 (N_19106,N_13121,N_14392);
nand U19107 (N_19107,N_12872,N_14092);
nand U19108 (N_19108,N_13298,N_11775);
and U19109 (N_19109,N_13685,N_14427);
xor U19110 (N_19110,N_13086,N_14126);
xor U19111 (N_19111,N_11786,N_11450);
or U19112 (N_19112,N_14325,N_14498);
nor U19113 (N_19113,N_11151,N_13067);
or U19114 (N_19114,N_10606,N_14150);
nor U19115 (N_19115,N_11690,N_10507);
and U19116 (N_19116,N_11601,N_11963);
nor U19117 (N_19117,N_10164,N_11997);
and U19118 (N_19118,N_14699,N_11482);
nor U19119 (N_19119,N_10345,N_10122);
or U19120 (N_19120,N_14940,N_14739);
nand U19121 (N_19121,N_11865,N_13518);
xor U19122 (N_19122,N_14787,N_11575);
nand U19123 (N_19123,N_10909,N_12034);
or U19124 (N_19124,N_13429,N_11540);
or U19125 (N_19125,N_10275,N_11987);
xor U19126 (N_19126,N_14274,N_13038);
or U19127 (N_19127,N_14626,N_12500);
xor U19128 (N_19128,N_14586,N_14033);
nand U19129 (N_19129,N_11700,N_14038);
xnor U19130 (N_19130,N_10390,N_11559);
or U19131 (N_19131,N_12475,N_13168);
nand U19132 (N_19132,N_13900,N_12266);
nand U19133 (N_19133,N_12423,N_14050);
xor U19134 (N_19134,N_12048,N_12327);
xnor U19135 (N_19135,N_12205,N_14859);
nand U19136 (N_19136,N_13090,N_14827);
nand U19137 (N_19137,N_13493,N_14006);
or U19138 (N_19138,N_14972,N_14434);
nor U19139 (N_19139,N_11666,N_10088);
xor U19140 (N_19140,N_13184,N_12283);
nand U19141 (N_19141,N_14582,N_12412);
and U19142 (N_19142,N_11482,N_14969);
nand U19143 (N_19143,N_10298,N_13446);
and U19144 (N_19144,N_11045,N_11616);
and U19145 (N_19145,N_14839,N_12481);
and U19146 (N_19146,N_10315,N_12650);
nor U19147 (N_19147,N_11828,N_13932);
and U19148 (N_19148,N_13308,N_14310);
nand U19149 (N_19149,N_10151,N_11718);
or U19150 (N_19150,N_10937,N_10441);
xnor U19151 (N_19151,N_13680,N_10812);
and U19152 (N_19152,N_13052,N_10919);
or U19153 (N_19153,N_12802,N_14581);
and U19154 (N_19154,N_13331,N_10316);
nor U19155 (N_19155,N_10606,N_14066);
xnor U19156 (N_19156,N_10685,N_12438);
xor U19157 (N_19157,N_10469,N_14159);
and U19158 (N_19158,N_10815,N_10813);
nor U19159 (N_19159,N_11407,N_13760);
or U19160 (N_19160,N_14092,N_12606);
and U19161 (N_19161,N_14321,N_12898);
nand U19162 (N_19162,N_12600,N_11801);
xor U19163 (N_19163,N_12136,N_14344);
and U19164 (N_19164,N_14911,N_11677);
or U19165 (N_19165,N_12804,N_12037);
or U19166 (N_19166,N_13345,N_13457);
nand U19167 (N_19167,N_13463,N_13191);
xor U19168 (N_19168,N_10401,N_10068);
nand U19169 (N_19169,N_14034,N_11398);
or U19170 (N_19170,N_12095,N_10874);
xor U19171 (N_19171,N_10469,N_11167);
nor U19172 (N_19172,N_12965,N_10834);
nand U19173 (N_19173,N_11245,N_12411);
nand U19174 (N_19174,N_14724,N_11751);
or U19175 (N_19175,N_14181,N_14072);
nand U19176 (N_19176,N_11480,N_13003);
xnor U19177 (N_19177,N_13510,N_12019);
nand U19178 (N_19178,N_12602,N_10663);
and U19179 (N_19179,N_12918,N_13155);
and U19180 (N_19180,N_12110,N_12192);
or U19181 (N_19181,N_14629,N_10141);
nor U19182 (N_19182,N_11495,N_14255);
nand U19183 (N_19183,N_14336,N_12448);
nand U19184 (N_19184,N_11915,N_14409);
nor U19185 (N_19185,N_14577,N_11935);
or U19186 (N_19186,N_14320,N_14296);
or U19187 (N_19187,N_13792,N_11442);
xnor U19188 (N_19188,N_14926,N_13472);
nor U19189 (N_19189,N_10587,N_13342);
nor U19190 (N_19190,N_14030,N_10274);
nand U19191 (N_19191,N_11627,N_12176);
xor U19192 (N_19192,N_13300,N_13465);
nand U19193 (N_19193,N_13773,N_10372);
xnor U19194 (N_19194,N_11986,N_13321);
and U19195 (N_19195,N_12204,N_10428);
nand U19196 (N_19196,N_12278,N_11009);
and U19197 (N_19197,N_14352,N_10824);
xor U19198 (N_19198,N_13212,N_12889);
and U19199 (N_19199,N_14144,N_12907);
xnor U19200 (N_19200,N_11607,N_14892);
nor U19201 (N_19201,N_14592,N_10112);
or U19202 (N_19202,N_10319,N_10576);
nand U19203 (N_19203,N_12486,N_13628);
nor U19204 (N_19204,N_10243,N_10480);
xor U19205 (N_19205,N_12931,N_13949);
xnor U19206 (N_19206,N_12008,N_13812);
or U19207 (N_19207,N_13810,N_14072);
nor U19208 (N_19208,N_10389,N_11826);
nand U19209 (N_19209,N_11277,N_11075);
nand U19210 (N_19210,N_13807,N_11514);
or U19211 (N_19211,N_10709,N_10484);
nand U19212 (N_19212,N_14956,N_14591);
nor U19213 (N_19213,N_12740,N_10241);
xor U19214 (N_19214,N_14155,N_13248);
or U19215 (N_19215,N_11245,N_11965);
or U19216 (N_19216,N_13602,N_10325);
nand U19217 (N_19217,N_12691,N_14169);
nand U19218 (N_19218,N_12245,N_14372);
or U19219 (N_19219,N_14303,N_13711);
and U19220 (N_19220,N_14379,N_12609);
and U19221 (N_19221,N_14819,N_11892);
xnor U19222 (N_19222,N_13734,N_11109);
and U19223 (N_19223,N_10666,N_10299);
nand U19224 (N_19224,N_10025,N_13000);
nand U19225 (N_19225,N_14446,N_10799);
nand U19226 (N_19226,N_13674,N_10156);
or U19227 (N_19227,N_10308,N_12941);
and U19228 (N_19228,N_10320,N_14312);
or U19229 (N_19229,N_12886,N_10592);
or U19230 (N_19230,N_14039,N_12786);
nor U19231 (N_19231,N_11162,N_14921);
or U19232 (N_19232,N_11403,N_10144);
nor U19233 (N_19233,N_14089,N_12902);
and U19234 (N_19234,N_10469,N_10599);
xnor U19235 (N_19235,N_14471,N_11534);
or U19236 (N_19236,N_11757,N_13149);
nand U19237 (N_19237,N_12447,N_12039);
xnor U19238 (N_19238,N_14122,N_12174);
xor U19239 (N_19239,N_14419,N_13977);
xor U19240 (N_19240,N_10012,N_11260);
nand U19241 (N_19241,N_14767,N_11664);
xor U19242 (N_19242,N_10091,N_11176);
xnor U19243 (N_19243,N_14075,N_13422);
nor U19244 (N_19244,N_13300,N_11235);
nand U19245 (N_19245,N_14604,N_11522);
or U19246 (N_19246,N_14529,N_11229);
nor U19247 (N_19247,N_14671,N_11320);
and U19248 (N_19248,N_14958,N_11379);
and U19249 (N_19249,N_12254,N_10054);
and U19250 (N_19250,N_10104,N_14272);
or U19251 (N_19251,N_11824,N_14555);
and U19252 (N_19252,N_13144,N_11431);
nor U19253 (N_19253,N_11738,N_13098);
and U19254 (N_19254,N_11902,N_13385);
or U19255 (N_19255,N_10984,N_11161);
nand U19256 (N_19256,N_14539,N_12948);
nor U19257 (N_19257,N_14902,N_10204);
and U19258 (N_19258,N_11023,N_14458);
and U19259 (N_19259,N_11944,N_14456);
nand U19260 (N_19260,N_11534,N_14661);
nand U19261 (N_19261,N_13314,N_10223);
and U19262 (N_19262,N_13063,N_13111);
or U19263 (N_19263,N_11734,N_12753);
xnor U19264 (N_19264,N_10672,N_14915);
or U19265 (N_19265,N_13371,N_13029);
nand U19266 (N_19266,N_12698,N_13875);
xnor U19267 (N_19267,N_10721,N_14485);
and U19268 (N_19268,N_10151,N_10682);
xor U19269 (N_19269,N_13717,N_10857);
nand U19270 (N_19270,N_13343,N_11247);
xnor U19271 (N_19271,N_13630,N_13460);
nand U19272 (N_19272,N_11532,N_11804);
nor U19273 (N_19273,N_13508,N_12991);
or U19274 (N_19274,N_11399,N_10726);
and U19275 (N_19275,N_13820,N_11599);
nand U19276 (N_19276,N_14593,N_10473);
or U19277 (N_19277,N_12546,N_10277);
and U19278 (N_19278,N_10018,N_14170);
nand U19279 (N_19279,N_14656,N_13248);
nor U19280 (N_19280,N_12332,N_10680);
xor U19281 (N_19281,N_11977,N_10936);
xnor U19282 (N_19282,N_13122,N_13390);
nor U19283 (N_19283,N_12208,N_11834);
or U19284 (N_19284,N_10416,N_10682);
xor U19285 (N_19285,N_13198,N_10448);
nor U19286 (N_19286,N_13762,N_14474);
nor U19287 (N_19287,N_12306,N_11485);
and U19288 (N_19288,N_14240,N_12797);
or U19289 (N_19289,N_10059,N_13297);
nor U19290 (N_19290,N_14708,N_14938);
nand U19291 (N_19291,N_13356,N_12376);
nor U19292 (N_19292,N_10712,N_10081);
or U19293 (N_19293,N_12442,N_14950);
and U19294 (N_19294,N_10210,N_13636);
xor U19295 (N_19295,N_13720,N_14341);
xor U19296 (N_19296,N_11713,N_12225);
nand U19297 (N_19297,N_10570,N_13777);
nand U19298 (N_19298,N_12780,N_13263);
nor U19299 (N_19299,N_11444,N_11100);
nand U19300 (N_19300,N_10779,N_14996);
nand U19301 (N_19301,N_10976,N_11767);
xor U19302 (N_19302,N_14002,N_11175);
nor U19303 (N_19303,N_12914,N_10006);
or U19304 (N_19304,N_14684,N_10544);
nor U19305 (N_19305,N_13844,N_14283);
and U19306 (N_19306,N_11602,N_12611);
xor U19307 (N_19307,N_10585,N_12209);
nand U19308 (N_19308,N_12068,N_14141);
nor U19309 (N_19309,N_12168,N_10449);
and U19310 (N_19310,N_12504,N_12945);
xor U19311 (N_19311,N_14144,N_14151);
nor U19312 (N_19312,N_12631,N_14008);
nand U19313 (N_19313,N_13765,N_13172);
nand U19314 (N_19314,N_10828,N_12618);
and U19315 (N_19315,N_14732,N_12406);
nor U19316 (N_19316,N_14021,N_11977);
xor U19317 (N_19317,N_14393,N_14468);
nand U19318 (N_19318,N_14300,N_10739);
or U19319 (N_19319,N_12649,N_14439);
xnor U19320 (N_19320,N_14064,N_13607);
or U19321 (N_19321,N_14729,N_13303);
and U19322 (N_19322,N_11558,N_14289);
and U19323 (N_19323,N_12682,N_10183);
nand U19324 (N_19324,N_13666,N_10500);
nor U19325 (N_19325,N_11105,N_12206);
and U19326 (N_19326,N_11333,N_14655);
xor U19327 (N_19327,N_11522,N_13519);
nor U19328 (N_19328,N_11088,N_11857);
or U19329 (N_19329,N_12323,N_12889);
nor U19330 (N_19330,N_10574,N_10744);
xnor U19331 (N_19331,N_13925,N_10523);
or U19332 (N_19332,N_13333,N_11717);
nor U19333 (N_19333,N_10919,N_12588);
nand U19334 (N_19334,N_10762,N_10916);
nor U19335 (N_19335,N_13677,N_12773);
nand U19336 (N_19336,N_12613,N_14763);
nor U19337 (N_19337,N_14092,N_10922);
and U19338 (N_19338,N_11112,N_10493);
xnor U19339 (N_19339,N_13707,N_14868);
nand U19340 (N_19340,N_11311,N_13705);
and U19341 (N_19341,N_13240,N_10968);
nand U19342 (N_19342,N_11244,N_12040);
or U19343 (N_19343,N_11140,N_12382);
or U19344 (N_19344,N_10629,N_14831);
and U19345 (N_19345,N_11628,N_13628);
nor U19346 (N_19346,N_13138,N_12729);
or U19347 (N_19347,N_12698,N_11970);
and U19348 (N_19348,N_14792,N_12071);
nand U19349 (N_19349,N_12012,N_10905);
and U19350 (N_19350,N_13015,N_12774);
or U19351 (N_19351,N_13758,N_12426);
nor U19352 (N_19352,N_14056,N_13906);
or U19353 (N_19353,N_13371,N_10359);
and U19354 (N_19354,N_14469,N_10918);
nand U19355 (N_19355,N_14115,N_14219);
nand U19356 (N_19356,N_12759,N_12211);
nor U19357 (N_19357,N_12614,N_10280);
xnor U19358 (N_19358,N_13791,N_12239);
and U19359 (N_19359,N_12263,N_14826);
or U19360 (N_19360,N_10207,N_12472);
xnor U19361 (N_19361,N_10553,N_13478);
nand U19362 (N_19362,N_11292,N_14104);
or U19363 (N_19363,N_14109,N_14975);
nand U19364 (N_19364,N_11438,N_14421);
xnor U19365 (N_19365,N_10912,N_11191);
or U19366 (N_19366,N_12434,N_14845);
nand U19367 (N_19367,N_13253,N_13783);
nand U19368 (N_19368,N_13872,N_14888);
xor U19369 (N_19369,N_11113,N_14929);
and U19370 (N_19370,N_10638,N_14608);
nor U19371 (N_19371,N_12347,N_13921);
xor U19372 (N_19372,N_14825,N_11657);
or U19373 (N_19373,N_13381,N_14168);
nand U19374 (N_19374,N_11343,N_14431);
and U19375 (N_19375,N_12048,N_11191);
nor U19376 (N_19376,N_10694,N_14020);
or U19377 (N_19377,N_14323,N_12765);
nand U19378 (N_19378,N_14951,N_12371);
xnor U19379 (N_19379,N_10986,N_12025);
xor U19380 (N_19380,N_14170,N_12056);
or U19381 (N_19381,N_13770,N_10858);
and U19382 (N_19382,N_12887,N_14335);
or U19383 (N_19383,N_14657,N_13735);
xnor U19384 (N_19384,N_11838,N_10863);
xor U19385 (N_19385,N_13580,N_10724);
nand U19386 (N_19386,N_13108,N_11381);
xnor U19387 (N_19387,N_13562,N_13983);
xnor U19388 (N_19388,N_10818,N_14648);
nor U19389 (N_19389,N_12573,N_11365);
nand U19390 (N_19390,N_11510,N_11047);
or U19391 (N_19391,N_11162,N_10250);
nand U19392 (N_19392,N_12318,N_12433);
nor U19393 (N_19393,N_12513,N_13327);
or U19394 (N_19394,N_10156,N_10325);
or U19395 (N_19395,N_10942,N_10106);
xnor U19396 (N_19396,N_13051,N_11025);
or U19397 (N_19397,N_13658,N_10463);
nor U19398 (N_19398,N_12566,N_12262);
xor U19399 (N_19399,N_13214,N_13630);
or U19400 (N_19400,N_12793,N_14384);
nand U19401 (N_19401,N_11792,N_13265);
and U19402 (N_19402,N_11398,N_11311);
and U19403 (N_19403,N_11191,N_14657);
and U19404 (N_19404,N_13627,N_10323);
or U19405 (N_19405,N_11757,N_14212);
or U19406 (N_19406,N_12288,N_11418);
or U19407 (N_19407,N_14859,N_11792);
nor U19408 (N_19408,N_13652,N_10225);
and U19409 (N_19409,N_11384,N_12993);
or U19410 (N_19410,N_10569,N_13354);
nand U19411 (N_19411,N_10969,N_12963);
nor U19412 (N_19412,N_12800,N_12088);
nor U19413 (N_19413,N_11889,N_13742);
nor U19414 (N_19414,N_11853,N_14867);
or U19415 (N_19415,N_10406,N_10471);
nor U19416 (N_19416,N_11083,N_13746);
nand U19417 (N_19417,N_11436,N_12752);
or U19418 (N_19418,N_13310,N_10987);
nand U19419 (N_19419,N_14307,N_13962);
nand U19420 (N_19420,N_12662,N_14001);
xnor U19421 (N_19421,N_14099,N_13308);
nand U19422 (N_19422,N_13703,N_14994);
or U19423 (N_19423,N_10877,N_11644);
nor U19424 (N_19424,N_11236,N_12614);
and U19425 (N_19425,N_13538,N_10457);
xor U19426 (N_19426,N_11258,N_11490);
and U19427 (N_19427,N_14172,N_13218);
nor U19428 (N_19428,N_10590,N_14003);
nor U19429 (N_19429,N_10240,N_14389);
and U19430 (N_19430,N_12409,N_14103);
nor U19431 (N_19431,N_13857,N_12815);
nor U19432 (N_19432,N_11930,N_14746);
or U19433 (N_19433,N_13264,N_12100);
or U19434 (N_19434,N_14793,N_13248);
nand U19435 (N_19435,N_10531,N_10177);
and U19436 (N_19436,N_14116,N_14950);
nor U19437 (N_19437,N_13807,N_10639);
or U19438 (N_19438,N_12463,N_12810);
nor U19439 (N_19439,N_12162,N_11975);
or U19440 (N_19440,N_14813,N_12320);
nand U19441 (N_19441,N_14158,N_10590);
nand U19442 (N_19442,N_12415,N_10508);
nand U19443 (N_19443,N_10693,N_12039);
nor U19444 (N_19444,N_10748,N_14201);
xor U19445 (N_19445,N_14360,N_12146);
nand U19446 (N_19446,N_12909,N_10782);
or U19447 (N_19447,N_14068,N_12947);
or U19448 (N_19448,N_10327,N_10016);
xnor U19449 (N_19449,N_10048,N_13124);
and U19450 (N_19450,N_13078,N_12929);
nor U19451 (N_19451,N_11555,N_11926);
and U19452 (N_19452,N_12930,N_11549);
and U19453 (N_19453,N_11475,N_11035);
or U19454 (N_19454,N_14681,N_14527);
and U19455 (N_19455,N_11952,N_11403);
or U19456 (N_19456,N_10981,N_11010);
or U19457 (N_19457,N_14079,N_12986);
nand U19458 (N_19458,N_14473,N_13690);
nor U19459 (N_19459,N_10082,N_11058);
and U19460 (N_19460,N_13301,N_14053);
or U19461 (N_19461,N_13240,N_14476);
nor U19462 (N_19462,N_14559,N_12847);
nand U19463 (N_19463,N_12836,N_14004);
nand U19464 (N_19464,N_13142,N_10203);
nor U19465 (N_19465,N_13891,N_13112);
and U19466 (N_19466,N_11975,N_10834);
xnor U19467 (N_19467,N_13869,N_14030);
nor U19468 (N_19468,N_10557,N_14657);
or U19469 (N_19469,N_10580,N_11196);
nor U19470 (N_19470,N_14317,N_11589);
or U19471 (N_19471,N_14455,N_13475);
or U19472 (N_19472,N_12515,N_10208);
or U19473 (N_19473,N_12674,N_13979);
and U19474 (N_19474,N_14722,N_10051);
or U19475 (N_19475,N_11625,N_10438);
or U19476 (N_19476,N_11470,N_11632);
nand U19477 (N_19477,N_13974,N_11296);
or U19478 (N_19478,N_10288,N_13359);
xor U19479 (N_19479,N_10422,N_13507);
xor U19480 (N_19480,N_14812,N_12894);
nand U19481 (N_19481,N_11728,N_14029);
nor U19482 (N_19482,N_13326,N_12041);
xnor U19483 (N_19483,N_10421,N_11909);
xnor U19484 (N_19484,N_10364,N_10473);
nand U19485 (N_19485,N_13836,N_11428);
nand U19486 (N_19486,N_11726,N_13669);
or U19487 (N_19487,N_11735,N_14489);
nor U19488 (N_19488,N_12037,N_12647);
nor U19489 (N_19489,N_11347,N_13835);
xnor U19490 (N_19490,N_11612,N_12290);
nand U19491 (N_19491,N_11935,N_12673);
nor U19492 (N_19492,N_10466,N_12361);
nor U19493 (N_19493,N_10462,N_12788);
nand U19494 (N_19494,N_10642,N_14198);
or U19495 (N_19495,N_13452,N_13336);
nand U19496 (N_19496,N_14871,N_12627);
and U19497 (N_19497,N_14107,N_13875);
or U19498 (N_19498,N_12630,N_13939);
nor U19499 (N_19499,N_10789,N_12138);
or U19500 (N_19500,N_13974,N_13484);
or U19501 (N_19501,N_10602,N_12592);
xnor U19502 (N_19502,N_13859,N_14855);
nand U19503 (N_19503,N_14354,N_14140);
and U19504 (N_19504,N_13418,N_13624);
xnor U19505 (N_19505,N_12570,N_11038);
nor U19506 (N_19506,N_11931,N_13277);
nand U19507 (N_19507,N_14885,N_11406);
xnor U19508 (N_19508,N_10768,N_14838);
nand U19509 (N_19509,N_13348,N_10890);
nor U19510 (N_19510,N_14859,N_12282);
or U19511 (N_19511,N_12175,N_14697);
nand U19512 (N_19512,N_12557,N_14590);
nor U19513 (N_19513,N_12245,N_14123);
and U19514 (N_19514,N_14782,N_12548);
and U19515 (N_19515,N_13755,N_11831);
xnor U19516 (N_19516,N_10410,N_11764);
nor U19517 (N_19517,N_11924,N_13591);
nor U19518 (N_19518,N_10391,N_11486);
or U19519 (N_19519,N_14153,N_10413);
or U19520 (N_19520,N_13379,N_12525);
and U19521 (N_19521,N_13846,N_12773);
xor U19522 (N_19522,N_11300,N_13087);
and U19523 (N_19523,N_10600,N_14069);
xor U19524 (N_19524,N_10405,N_12507);
nand U19525 (N_19525,N_12539,N_14303);
or U19526 (N_19526,N_14338,N_10995);
nand U19527 (N_19527,N_13884,N_10133);
nor U19528 (N_19528,N_12551,N_13612);
xnor U19529 (N_19529,N_11310,N_14840);
nor U19530 (N_19530,N_14416,N_13218);
xnor U19531 (N_19531,N_11646,N_14888);
nor U19532 (N_19532,N_10171,N_14359);
nor U19533 (N_19533,N_14327,N_14578);
and U19534 (N_19534,N_14215,N_14138);
and U19535 (N_19535,N_10871,N_13043);
nor U19536 (N_19536,N_14941,N_10122);
and U19537 (N_19537,N_10518,N_14182);
and U19538 (N_19538,N_13280,N_11724);
xor U19539 (N_19539,N_13630,N_13806);
and U19540 (N_19540,N_13285,N_12547);
and U19541 (N_19541,N_14212,N_10399);
nor U19542 (N_19542,N_10159,N_12148);
and U19543 (N_19543,N_10878,N_12406);
and U19544 (N_19544,N_11088,N_10585);
nor U19545 (N_19545,N_11105,N_11229);
and U19546 (N_19546,N_14493,N_12665);
xnor U19547 (N_19547,N_12942,N_11225);
nor U19548 (N_19548,N_12275,N_14290);
xor U19549 (N_19549,N_14147,N_12560);
or U19550 (N_19550,N_10202,N_10299);
xnor U19551 (N_19551,N_11824,N_13090);
and U19552 (N_19552,N_12991,N_13125);
nor U19553 (N_19553,N_10632,N_10060);
and U19554 (N_19554,N_10354,N_13747);
nor U19555 (N_19555,N_13047,N_11986);
or U19556 (N_19556,N_14299,N_10054);
nand U19557 (N_19557,N_12237,N_14193);
nor U19558 (N_19558,N_13162,N_14512);
xnor U19559 (N_19559,N_13575,N_14123);
nand U19560 (N_19560,N_14726,N_14507);
nand U19561 (N_19561,N_11144,N_14583);
or U19562 (N_19562,N_13054,N_14059);
nand U19563 (N_19563,N_12962,N_12324);
nor U19564 (N_19564,N_10471,N_11266);
or U19565 (N_19565,N_14330,N_14971);
nor U19566 (N_19566,N_14295,N_12922);
and U19567 (N_19567,N_14092,N_13841);
nor U19568 (N_19568,N_12551,N_13503);
nor U19569 (N_19569,N_14250,N_14112);
xnor U19570 (N_19570,N_11788,N_10411);
nand U19571 (N_19571,N_10519,N_12510);
or U19572 (N_19572,N_13003,N_10186);
nand U19573 (N_19573,N_10898,N_10436);
xor U19574 (N_19574,N_14266,N_10855);
and U19575 (N_19575,N_13818,N_10659);
or U19576 (N_19576,N_13302,N_10780);
or U19577 (N_19577,N_14167,N_11037);
and U19578 (N_19578,N_13789,N_11420);
nand U19579 (N_19579,N_13810,N_11909);
nor U19580 (N_19580,N_14439,N_12268);
nand U19581 (N_19581,N_11262,N_13939);
nand U19582 (N_19582,N_10443,N_11119);
and U19583 (N_19583,N_12081,N_13491);
xor U19584 (N_19584,N_10306,N_13324);
nand U19585 (N_19585,N_11233,N_13828);
and U19586 (N_19586,N_10701,N_14760);
and U19587 (N_19587,N_11664,N_12956);
and U19588 (N_19588,N_14099,N_14881);
or U19589 (N_19589,N_14172,N_12084);
xor U19590 (N_19590,N_10442,N_10465);
or U19591 (N_19591,N_12756,N_11905);
or U19592 (N_19592,N_14508,N_13185);
xnor U19593 (N_19593,N_11336,N_10968);
and U19594 (N_19594,N_14705,N_14837);
xor U19595 (N_19595,N_13326,N_13131);
or U19596 (N_19596,N_13931,N_10815);
nand U19597 (N_19597,N_10123,N_13556);
nor U19598 (N_19598,N_12466,N_12739);
xor U19599 (N_19599,N_11116,N_13893);
nand U19600 (N_19600,N_13369,N_13861);
and U19601 (N_19601,N_10767,N_12818);
xor U19602 (N_19602,N_11781,N_14629);
xnor U19603 (N_19603,N_11672,N_11740);
nand U19604 (N_19604,N_12543,N_10544);
nand U19605 (N_19605,N_13453,N_13213);
nand U19606 (N_19606,N_13463,N_11215);
and U19607 (N_19607,N_12567,N_13016);
nand U19608 (N_19608,N_12958,N_14523);
or U19609 (N_19609,N_13413,N_12845);
nor U19610 (N_19610,N_10850,N_12518);
or U19611 (N_19611,N_12046,N_14971);
nand U19612 (N_19612,N_14581,N_11161);
nor U19613 (N_19613,N_10284,N_13049);
nor U19614 (N_19614,N_11980,N_12385);
xnor U19615 (N_19615,N_10960,N_11870);
and U19616 (N_19616,N_10980,N_10641);
xnor U19617 (N_19617,N_13499,N_11088);
and U19618 (N_19618,N_10079,N_14608);
nor U19619 (N_19619,N_11609,N_11507);
or U19620 (N_19620,N_11505,N_10305);
and U19621 (N_19621,N_14208,N_10850);
nor U19622 (N_19622,N_12425,N_14774);
nor U19623 (N_19623,N_11754,N_10914);
or U19624 (N_19624,N_12220,N_14999);
or U19625 (N_19625,N_11561,N_13341);
nor U19626 (N_19626,N_12664,N_13018);
or U19627 (N_19627,N_11219,N_14245);
nor U19628 (N_19628,N_13044,N_12404);
xnor U19629 (N_19629,N_12926,N_12159);
nor U19630 (N_19630,N_14273,N_10572);
and U19631 (N_19631,N_14177,N_11558);
nor U19632 (N_19632,N_14754,N_10443);
or U19633 (N_19633,N_12365,N_12619);
or U19634 (N_19634,N_13693,N_12660);
or U19635 (N_19635,N_11064,N_13803);
and U19636 (N_19636,N_10732,N_13610);
xor U19637 (N_19637,N_12908,N_12116);
nand U19638 (N_19638,N_14120,N_11775);
nand U19639 (N_19639,N_14169,N_10914);
and U19640 (N_19640,N_10707,N_14659);
nor U19641 (N_19641,N_14431,N_10754);
nor U19642 (N_19642,N_11862,N_13586);
and U19643 (N_19643,N_13938,N_14052);
xnor U19644 (N_19644,N_13760,N_10846);
xor U19645 (N_19645,N_10264,N_10640);
xor U19646 (N_19646,N_11705,N_13889);
nand U19647 (N_19647,N_11704,N_13178);
nand U19648 (N_19648,N_10572,N_11267);
xor U19649 (N_19649,N_14199,N_13918);
nor U19650 (N_19650,N_10474,N_12800);
xnor U19651 (N_19651,N_13435,N_11171);
nor U19652 (N_19652,N_14948,N_14176);
nor U19653 (N_19653,N_14379,N_14914);
xnor U19654 (N_19654,N_12521,N_14749);
nor U19655 (N_19655,N_13613,N_12965);
or U19656 (N_19656,N_10179,N_12376);
nor U19657 (N_19657,N_13289,N_13410);
or U19658 (N_19658,N_13385,N_11606);
nand U19659 (N_19659,N_14506,N_10244);
and U19660 (N_19660,N_10522,N_13326);
nor U19661 (N_19661,N_10851,N_12337);
and U19662 (N_19662,N_11387,N_14083);
or U19663 (N_19663,N_13079,N_10027);
nor U19664 (N_19664,N_10834,N_10485);
nor U19665 (N_19665,N_13259,N_13191);
and U19666 (N_19666,N_12427,N_14289);
xnor U19667 (N_19667,N_14811,N_11412);
nand U19668 (N_19668,N_12247,N_14268);
nor U19669 (N_19669,N_13921,N_10968);
nor U19670 (N_19670,N_12882,N_14401);
xnor U19671 (N_19671,N_14624,N_12580);
or U19672 (N_19672,N_13134,N_13025);
nor U19673 (N_19673,N_13751,N_10900);
xor U19674 (N_19674,N_11320,N_13201);
nand U19675 (N_19675,N_11876,N_12891);
nor U19676 (N_19676,N_12890,N_11519);
nor U19677 (N_19677,N_12083,N_13070);
nor U19678 (N_19678,N_14183,N_14036);
nor U19679 (N_19679,N_13663,N_12259);
and U19680 (N_19680,N_14584,N_12262);
nand U19681 (N_19681,N_10237,N_12067);
nand U19682 (N_19682,N_12373,N_12960);
and U19683 (N_19683,N_11948,N_14747);
nor U19684 (N_19684,N_10989,N_13187);
and U19685 (N_19685,N_10487,N_11416);
nand U19686 (N_19686,N_10044,N_10992);
nand U19687 (N_19687,N_12687,N_12616);
nand U19688 (N_19688,N_11271,N_13958);
and U19689 (N_19689,N_12177,N_10569);
and U19690 (N_19690,N_13847,N_14741);
or U19691 (N_19691,N_14899,N_12917);
xnor U19692 (N_19692,N_13008,N_14360);
nor U19693 (N_19693,N_10363,N_10316);
and U19694 (N_19694,N_11648,N_14151);
nor U19695 (N_19695,N_14293,N_13503);
and U19696 (N_19696,N_13526,N_11004);
and U19697 (N_19697,N_12889,N_12769);
nor U19698 (N_19698,N_10649,N_10203);
and U19699 (N_19699,N_13060,N_12921);
or U19700 (N_19700,N_12650,N_13955);
xnor U19701 (N_19701,N_14143,N_12003);
or U19702 (N_19702,N_13610,N_10854);
nand U19703 (N_19703,N_10955,N_12755);
or U19704 (N_19704,N_12512,N_14792);
and U19705 (N_19705,N_11533,N_11262);
nor U19706 (N_19706,N_14585,N_11603);
nand U19707 (N_19707,N_12613,N_14092);
nand U19708 (N_19708,N_10014,N_10478);
and U19709 (N_19709,N_13210,N_10999);
nand U19710 (N_19710,N_12842,N_13932);
or U19711 (N_19711,N_12324,N_13532);
nor U19712 (N_19712,N_13950,N_10830);
or U19713 (N_19713,N_13847,N_10425);
xnor U19714 (N_19714,N_11047,N_14900);
or U19715 (N_19715,N_10838,N_12061);
nor U19716 (N_19716,N_11506,N_11389);
and U19717 (N_19717,N_10482,N_10917);
and U19718 (N_19718,N_11290,N_10517);
or U19719 (N_19719,N_12807,N_12079);
or U19720 (N_19720,N_10680,N_12506);
and U19721 (N_19721,N_10027,N_11988);
xnor U19722 (N_19722,N_13431,N_14852);
and U19723 (N_19723,N_14698,N_13706);
or U19724 (N_19724,N_10893,N_12217);
xor U19725 (N_19725,N_13695,N_14630);
nor U19726 (N_19726,N_11494,N_11983);
nand U19727 (N_19727,N_12869,N_11160);
nor U19728 (N_19728,N_10083,N_13546);
nand U19729 (N_19729,N_13123,N_11388);
or U19730 (N_19730,N_12871,N_10265);
and U19731 (N_19731,N_14420,N_13224);
nor U19732 (N_19732,N_10403,N_11373);
xnor U19733 (N_19733,N_14045,N_14178);
or U19734 (N_19734,N_14136,N_12845);
xnor U19735 (N_19735,N_12526,N_14377);
nor U19736 (N_19736,N_11204,N_12653);
nand U19737 (N_19737,N_10441,N_11565);
and U19738 (N_19738,N_14024,N_11221);
and U19739 (N_19739,N_11295,N_12573);
or U19740 (N_19740,N_11058,N_11128);
nor U19741 (N_19741,N_10102,N_13745);
xnor U19742 (N_19742,N_12437,N_14889);
or U19743 (N_19743,N_12907,N_10154);
xnor U19744 (N_19744,N_10775,N_12040);
nor U19745 (N_19745,N_14628,N_14274);
or U19746 (N_19746,N_10121,N_10122);
nor U19747 (N_19747,N_14462,N_13700);
nor U19748 (N_19748,N_11201,N_11512);
nand U19749 (N_19749,N_11133,N_12708);
nor U19750 (N_19750,N_10475,N_12148);
nor U19751 (N_19751,N_11953,N_14062);
or U19752 (N_19752,N_14684,N_10179);
and U19753 (N_19753,N_10389,N_10614);
nand U19754 (N_19754,N_12321,N_13163);
xor U19755 (N_19755,N_11216,N_14981);
nand U19756 (N_19756,N_10672,N_13217);
xor U19757 (N_19757,N_10636,N_12805);
and U19758 (N_19758,N_10317,N_10175);
and U19759 (N_19759,N_10398,N_12763);
nor U19760 (N_19760,N_13758,N_14842);
nand U19761 (N_19761,N_14425,N_10835);
xnor U19762 (N_19762,N_12770,N_13075);
and U19763 (N_19763,N_13037,N_11986);
or U19764 (N_19764,N_14653,N_14904);
nor U19765 (N_19765,N_10926,N_11152);
nand U19766 (N_19766,N_12266,N_10461);
nand U19767 (N_19767,N_14358,N_11222);
or U19768 (N_19768,N_13454,N_11383);
nand U19769 (N_19769,N_10563,N_12680);
nor U19770 (N_19770,N_13475,N_12516);
nand U19771 (N_19771,N_11821,N_13570);
and U19772 (N_19772,N_12908,N_14167);
or U19773 (N_19773,N_12199,N_12667);
nand U19774 (N_19774,N_13337,N_13643);
xor U19775 (N_19775,N_11861,N_14607);
or U19776 (N_19776,N_12204,N_11063);
and U19777 (N_19777,N_10192,N_12718);
nand U19778 (N_19778,N_11514,N_11001);
or U19779 (N_19779,N_14061,N_10003);
and U19780 (N_19780,N_12105,N_12493);
or U19781 (N_19781,N_14447,N_10714);
nand U19782 (N_19782,N_10050,N_12455);
or U19783 (N_19783,N_13622,N_14868);
nand U19784 (N_19784,N_11346,N_11058);
or U19785 (N_19785,N_10994,N_14918);
or U19786 (N_19786,N_11797,N_14164);
or U19787 (N_19787,N_13013,N_11862);
nor U19788 (N_19788,N_11480,N_10433);
or U19789 (N_19789,N_10444,N_10363);
nand U19790 (N_19790,N_13917,N_13098);
nor U19791 (N_19791,N_13679,N_11032);
xor U19792 (N_19792,N_13960,N_13776);
xnor U19793 (N_19793,N_14597,N_14272);
xnor U19794 (N_19794,N_13125,N_13189);
or U19795 (N_19795,N_11524,N_12055);
or U19796 (N_19796,N_11221,N_12960);
nor U19797 (N_19797,N_11812,N_10772);
and U19798 (N_19798,N_12982,N_11729);
nor U19799 (N_19799,N_11183,N_13539);
nand U19800 (N_19800,N_11115,N_13552);
nand U19801 (N_19801,N_11650,N_12996);
or U19802 (N_19802,N_12855,N_11169);
xor U19803 (N_19803,N_13224,N_11712);
xor U19804 (N_19804,N_11388,N_14707);
nor U19805 (N_19805,N_14079,N_10632);
nor U19806 (N_19806,N_11775,N_10480);
xnor U19807 (N_19807,N_14090,N_14217);
and U19808 (N_19808,N_10839,N_11821);
nand U19809 (N_19809,N_13977,N_11947);
nand U19810 (N_19810,N_11622,N_10475);
or U19811 (N_19811,N_10841,N_13028);
or U19812 (N_19812,N_11954,N_14398);
and U19813 (N_19813,N_10906,N_13442);
nor U19814 (N_19814,N_12780,N_13978);
nand U19815 (N_19815,N_13774,N_12262);
nand U19816 (N_19816,N_12711,N_12579);
nor U19817 (N_19817,N_11706,N_14479);
and U19818 (N_19818,N_10117,N_10762);
nand U19819 (N_19819,N_11347,N_13853);
nor U19820 (N_19820,N_11050,N_14102);
xnor U19821 (N_19821,N_10591,N_11130);
or U19822 (N_19822,N_11210,N_11072);
and U19823 (N_19823,N_10490,N_10473);
nand U19824 (N_19824,N_12497,N_12581);
nand U19825 (N_19825,N_11659,N_14258);
and U19826 (N_19826,N_14058,N_11230);
and U19827 (N_19827,N_11459,N_10225);
nor U19828 (N_19828,N_13556,N_12649);
xnor U19829 (N_19829,N_11692,N_10207);
and U19830 (N_19830,N_13257,N_10076);
or U19831 (N_19831,N_12772,N_13082);
and U19832 (N_19832,N_10084,N_10291);
and U19833 (N_19833,N_12573,N_14974);
and U19834 (N_19834,N_10783,N_11151);
nor U19835 (N_19835,N_14489,N_13182);
nor U19836 (N_19836,N_11219,N_14819);
xnor U19837 (N_19837,N_13778,N_12576);
or U19838 (N_19838,N_13082,N_10051);
or U19839 (N_19839,N_12824,N_12411);
or U19840 (N_19840,N_14136,N_14941);
nand U19841 (N_19841,N_14665,N_13096);
nand U19842 (N_19842,N_10297,N_14087);
nand U19843 (N_19843,N_13874,N_13134);
xor U19844 (N_19844,N_14946,N_14482);
nor U19845 (N_19845,N_13290,N_14318);
and U19846 (N_19846,N_12561,N_14072);
xor U19847 (N_19847,N_10553,N_13480);
nor U19848 (N_19848,N_12690,N_12497);
nor U19849 (N_19849,N_10087,N_10425);
or U19850 (N_19850,N_13614,N_12764);
xnor U19851 (N_19851,N_12626,N_11649);
xor U19852 (N_19852,N_14535,N_13537);
nor U19853 (N_19853,N_11835,N_14475);
xor U19854 (N_19854,N_13867,N_12755);
or U19855 (N_19855,N_11153,N_10024);
xnor U19856 (N_19856,N_10636,N_11053);
nor U19857 (N_19857,N_12610,N_11982);
nand U19858 (N_19858,N_14093,N_10907);
nand U19859 (N_19859,N_11402,N_13546);
nor U19860 (N_19860,N_14352,N_14501);
nand U19861 (N_19861,N_14507,N_13492);
nor U19862 (N_19862,N_10070,N_14994);
nor U19863 (N_19863,N_14517,N_12113);
or U19864 (N_19864,N_11939,N_14359);
or U19865 (N_19865,N_11836,N_14953);
xor U19866 (N_19866,N_11254,N_13564);
xnor U19867 (N_19867,N_11169,N_14672);
nand U19868 (N_19868,N_10444,N_10995);
or U19869 (N_19869,N_10107,N_12394);
and U19870 (N_19870,N_12477,N_10172);
xnor U19871 (N_19871,N_11751,N_14306);
or U19872 (N_19872,N_14167,N_13176);
xnor U19873 (N_19873,N_12800,N_12023);
xnor U19874 (N_19874,N_13426,N_14722);
nand U19875 (N_19875,N_11562,N_10002);
nor U19876 (N_19876,N_11169,N_12554);
and U19877 (N_19877,N_11032,N_11913);
nor U19878 (N_19878,N_13547,N_10750);
and U19879 (N_19879,N_14714,N_10358);
and U19880 (N_19880,N_13753,N_12791);
nand U19881 (N_19881,N_10298,N_11757);
xnor U19882 (N_19882,N_14992,N_11730);
xor U19883 (N_19883,N_14585,N_10695);
nor U19884 (N_19884,N_13588,N_11176);
nor U19885 (N_19885,N_12742,N_11534);
nand U19886 (N_19886,N_10013,N_13157);
or U19887 (N_19887,N_10394,N_10626);
nand U19888 (N_19888,N_13171,N_13759);
nor U19889 (N_19889,N_10165,N_11006);
and U19890 (N_19890,N_10339,N_10691);
or U19891 (N_19891,N_11032,N_10385);
nor U19892 (N_19892,N_14118,N_11050);
nor U19893 (N_19893,N_10610,N_10583);
nand U19894 (N_19894,N_14631,N_14471);
nand U19895 (N_19895,N_13291,N_12552);
xor U19896 (N_19896,N_13343,N_10393);
nand U19897 (N_19897,N_12457,N_14690);
or U19898 (N_19898,N_12040,N_10055);
nand U19899 (N_19899,N_11119,N_13336);
nand U19900 (N_19900,N_14547,N_13981);
nand U19901 (N_19901,N_14704,N_12792);
or U19902 (N_19902,N_12864,N_13945);
or U19903 (N_19903,N_12006,N_11337);
xor U19904 (N_19904,N_12062,N_11670);
and U19905 (N_19905,N_11971,N_14138);
and U19906 (N_19906,N_13900,N_11535);
nor U19907 (N_19907,N_14524,N_10244);
nand U19908 (N_19908,N_12275,N_14230);
or U19909 (N_19909,N_10112,N_10557);
nand U19910 (N_19910,N_12464,N_13061);
nor U19911 (N_19911,N_14802,N_14112);
nand U19912 (N_19912,N_12808,N_11072);
nand U19913 (N_19913,N_11393,N_10535);
and U19914 (N_19914,N_10830,N_13426);
nor U19915 (N_19915,N_14125,N_10568);
nand U19916 (N_19916,N_13726,N_14158);
or U19917 (N_19917,N_14183,N_14544);
xnor U19918 (N_19918,N_11549,N_13357);
or U19919 (N_19919,N_11017,N_10434);
xnor U19920 (N_19920,N_13919,N_12062);
nand U19921 (N_19921,N_13980,N_14679);
and U19922 (N_19922,N_14332,N_10561);
or U19923 (N_19923,N_13696,N_12305);
xor U19924 (N_19924,N_10815,N_11241);
nor U19925 (N_19925,N_14403,N_11900);
nand U19926 (N_19926,N_12473,N_11551);
nor U19927 (N_19927,N_13898,N_14732);
nand U19928 (N_19928,N_12379,N_14130);
xnor U19929 (N_19929,N_11661,N_12079);
nand U19930 (N_19930,N_12599,N_14310);
nand U19931 (N_19931,N_10647,N_11930);
or U19932 (N_19932,N_14838,N_13005);
nor U19933 (N_19933,N_13185,N_13911);
xnor U19934 (N_19934,N_13633,N_12039);
and U19935 (N_19935,N_10450,N_13238);
xnor U19936 (N_19936,N_10589,N_10053);
nor U19937 (N_19937,N_10721,N_11320);
nor U19938 (N_19938,N_12083,N_11999);
nand U19939 (N_19939,N_14132,N_13890);
nand U19940 (N_19940,N_14426,N_10899);
or U19941 (N_19941,N_14313,N_10158);
or U19942 (N_19942,N_12896,N_14632);
xnor U19943 (N_19943,N_14826,N_14450);
nand U19944 (N_19944,N_14674,N_10677);
or U19945 (N_19945,N_14797,N_12783);
or U19946 (N_19946,N_14288,N_13608);
nand U19947 (N_19947,N_12821,N_14493);
xnor U19948 (N_19948,N_12286,N_11410);
nand U19949 (N_19949,N_10317,N_14412);
nor U19950 (N_19950,N_11780,N_11458);
nor U19951 (N_19951,N_10748,N_11099);
and U19952 (N_19952,N_10403,N_10306);
or U19953 (N_19953,N_11949,N_10302);
xor U19954 (N_19954,N_13234,N_10084);
nor U19955 (N_19955,N_10309,N_11764);
xnor U19956 (N_19956,N_14783,N_11956);
xor U19957 (N_19957,N_14149,N_12363);
nand U19958 (N_19958,N_14339,N_13422);
or U19959 (N_19959,N_14831,N_14803);
xor U19960 (N_19960,N_11972,N_11466);
or U19961 (N_19961,N_11448,N_13811);
nor U19962 (N_19962,N_14433,N_14490);
nor U19963 (N_19963,N_10772,N_12790);
nor U19964 (N_19964,N_14141,N_14060);
nor U19965 (N_19965,N_12297,N_12161);
xnor U19966 (N_19966,N_14649,N_14211);
nor U19967 (N_19967,N_14787,N_10407);
nor U19968 (N_19968,N_10294,N_12122);
xnor U19969 (N_19969,N_11240,N_10330);
and U19970 (N_19970,N_12610,N_10398);
and U19971 (N_19971,N_12838,N_12450);
xnor U19972 (N_19972,N_13121,N_12281);
nand U19973 (N_19973,N_13244,N_10061);
nor U19974 (N_19974,N_10564,N_10586);
or U19975 (N_19975,N_12521,N_10764);
nor U19976 (N_19976,N_13308,N_11324);
nand U19977 (N_19977,N_14565,N_10387);
nand U19978 (N_19978,N_13292,N_14287);
and U19979 (N_19979,N_10457,N_10472);
or U19980 (N_19980,N_10377,N_13197);
and U19981 (N_19981,N_12858,N_14057);
xor U19982 (N_19982,N_11436,N_12442);
and U19983 (N_19983,N_13242,N_14986);
nor U19984 (N_19984,N_12336,N_13559);
nor U19985 (N_19985,N_10730,N_11498);
xnor U19986 (N_19986,N_12035,N_13560);
nand U19987 (N_19987,N_10599,N_11539);
xor U19988 (N_19988,N_10703,N_10572);
xor U19989 (N_19989,N_11162,N_10341);
nand U19990 (N_19990,N_14029,N_11565);
nor U19991 (N_19991,N_11107,N_14611);
or U19992 (N_19992,N_13570,N_12645);
xnor U19993 (N_19993,N_10656,N_14432);
nand U19994 (N_19994,N_12318,N_12503);
or U19995 (N_19995,N_11976,N_12529);
xnor U19996 (N_19996,N_12399,N_13354);
xor U19997 (N_19997,N_13197,N_13738);
and U19998 (N_19998,N_10667,N_14140);
nor U19999 (N_19999,N_12815,N_11028);
nor U20000 (N_20000,N_16040,N_17546);
nand U20001 (N_20001,N_16361,N_15250);
and U20002 (N_20002,N_18582,N_16250);
and U20003 (N_20003,N_16784,N_18690);
or U20004 (N_20004,N_18801,N_18304);
nor U20005 (N_20005,N_16023,N_16923);
or U20006 (N_20006,N_16930,N_17242);
nand U20007 (N_20007,N_17527,N_16936);
or U20008 (N_20008,N_19155,N_15795);
nor U20009 (N_20009,N_15573,N_16215);
or U20010 (N_20010,N_19789,N_18506);
xnor U20011 (N_20011,N_17344,N_15563);
xnor U20012 (N_20012,N_18658,N_15340);
nand U20013 (N_20013,N_16367,N_19392);
nor U20014 (N_20014,N_19169,N_19989);
or U20015 (N_20015,N_15064,N_16920);
or U20016 (N_20016,N_15289,N_19810);
nand U20017 (N_20017,N_19573,N_19150);
nor U20018 (N_20018,N_15155,N_15226);
and U20019 (N_20019,N_17632,N_18025);
nor U20020 (N_20020,N_18300,N_16392);
nor U20021 (N_20021,N_18626,N_16054);
nand U20022 (N_20022,N_17309,N_18662);
and U20023 (N_20023,N_17573,N_16033);
or U20024 (N_20024,N_16173,N_18759);
xnor U20025 (N_20025,N_19553,N_18329);
xnor U20026 (N_20026,N_17924,N_17779);
or U20027 (N_20027,N_19937,N_16551);
nand U20028 (N_20028,N_19233,N_16888);
nor U20029 (N_20029,N_17897,N_15686);
or U20030 (N_20030,N_18008,N_15134);
and U20031 (N_20031,N_15982,N_18598);
and U20032 (N_20032,N_16541,N_17377);
nand U20033 (N_20033,N_18794,N_18800);
and U20034 (N_20034,N_17722,N_15094);
nand U20035 (N_20035,N_17734,N_15277);
xor U20036 (N_20036,N_16430,N_16654);
xor U20037 (N_20037,N_15848,N_18637);
nor U20038 (N_20038,N_19873,N_17379);
or U20039 (N_20039,N_19589,N_17977);
nor U20040 (N_20040,N_16402,N_17757);
xnor U20041 (N_20041,N_16036,N_16427);
nand U20042 (N_20042,N_17305,N_17701);
nand U20043 (N_20043,N_19729,N_16230);
nor U20044 (N_20044,N_18871,N_18572);
nand U20045 (N_20045,N_18490,N_19653);
nand U20046 (N_20046,N_18500,N_18767);
and U20047 (N_20047,N_16295,N_16927);
nor U20048 (N_20048,N_16333,N_15859);
nor U20049 (N_20049,N_18494,N_16415);
or U20050 (N_20050,N_16824,N_16629);
and U20051 (N_20051,N_19707,N_18846);
xnor U20052 (N_20052,N_18864,N_16357);
or U20053 (N_20053,N_18996,N_15488);
nor U20054 (N_20054,N_19166,N_19428);
or U20055 (N_20055,N_16963,N_17611);
nand U20056 (N_20056,N_16907,N_18897);
or U20057 (N_20057,N_15205,N_15577);
and U20058 (N_20058,N_16240,N_17232);
nor U20059 (N_20059,N_19242,N_17851);
and U20060 (N_20060,N_17692,N_17028);
nor U20061 (N_20061,N_19574,N_15156);
xor U20062 (N_20062,N_15310,N_16224);
nand U20063 (N_20063,N_17114,N_18562);
xnor U20064 (N_20064,N_18636,N_18954);
or U20065 (N_20065,N_16309,N_16314);
and U20066 (N_20066,N_18590,N_19028);
xnor U20067 (N_20067,N_18323,N_16089);
and U20068 (N_20068,N_19202,N_18452);
and U20069 (N_20069,N_15805,N_16887);
nor U20070 (N_20070,N_19910,N_18896);
nand U20071 (N_20071,N_15482,N_15548);
xnor U20072 (N_20072,N_17210,N_16535);
and U20073 (N_20073,N_15460,N_16571);
xnor U20074 (N_20074,N_15253,N_17358);
xnor U20075 (N_20075,N_16006,N_18170);
xnor U20076 (N_20076,N_19550,N_15216);
nand U20077 (N_20077,N_17990,N_15063);
nand U20078 (N_20078,N_19737,N_19476);
and U20079 (N_20079,N_15519,N_16220);
xor U20080 (N_20080,N_17254,N_19970);
nand U20081 (N_20081,N_18503,N_18212);
nor U20082 (N_20082,N_19103,N_18442);
and U20083 (N_20083,N_19112,N_15237);
and U20084 (N_20084,N_16441,N_15139);
and U20085 (N_20085,N_19452,N_18236);
and U20086 (N_20086,N_16901,N_16334);
nand U20087 (N_20087,N_16649,N_15481);
nor U20088 (N_20088,N_19631,N_17556);
nand U20089 (N_20089,N_15719,N_15713);
nand U20090 (N_20090,N_17269,N_18963);
or U20091 (N_20091,N_17070,N_15590);
nand U20092 (N_20092,N_15542,N_17748);
xnor U20093 (N_20093,N_15889,N_18475);
nor U20094 (N_20094,N_15832,N_18029);
nor U20095 (N_20095,N_17130,N_19305);
and U20096 (N_20096,N_16792,N_17832);
or U20097 (N_20097,N_18751,N_19814);
nor U20098 (N_20098,N_19416,N_19340);
xor U20099 (N_20099,N_16097,N_16957);
or U20100 (N_20100,N_18695,N_15788);
nor U20101 (N_20101,N_16417,N_17282);
nor U20102 (N_20102,N_19453,N_18938);
and U20103 (N_20103,N_18327,N_18497);
nor U20104 (N_20104,N_15148,N_18021);
nor U20105 (N_20105,N_16422,N_15374);
and U20106 (N_20106,N_15418,N_16911);
xor U20107 (N_20107,N_15341,N_19422);
xnor U20108 (N_20108,N_15305,N_16646);
xnor U20109 (N_20109,N_15407,N_15614);
xnor U20110 (N_20110,N_17158,N_19128);
nand U20111 (N_20111,N_18026,N_17155);
nor U20112 (N_20112,N_17252,N_16491);
and U20113 (N_20113,N_16081,N_18046);
xor U20114 (N_20114,N_15292,N_15397);
xnor U20115 (N_20115,N_16279,N_15712);
xnor U20116 (N_20116,N_18196,N_19558);
xor U20117 (N_20117,N_16436,N_15589);
nand U20118 (N_20118,N_16876,N_19352);
or U20119 (N_20119,N_17142,N_16604);
or U20120 (N_20120,N_15091,N_19885);
nor U20121 (N_20121,N_19827,N_15122);
nor U20122 (N_20122,N_19632,N_19564);
nand U20123 (N_20123,N_18015,N_16517);
nand U20124 (N_20124,N_18863,N_16691);
and U20125 (N_20125,N_15471,N_16530);
and U20126 (N_20126,N_17879,N_18489);
or U20127 (N_20127,N_15746,N_19815);
and U20128 (N_20128,N_15888,N_18734);
nand U20129 (N_20129,N_17886,N_15401);
and U20130 (N_20130,N_19391,N_15348);
and U20131 (N_20131,N_19146,N_19681);
or U20132 (N_20132,N_16159,N_19140);
nor U20133 (N_20133,N_15144,N_17314);
nand U20134 (N_20134,N_18354,N_19670);
and U20135 (N_20135,N_15796,N_19537);
or U20136 (N_20136,N_19967,N_16744);
or U20137 (N_20137,N_18247,N_18701);
nand U20138 (N_20138,N_15120,N_16166);
nand U20139 (N_20139,N_15092,N_15035);
nand U20140 (N_20140,N_17827,N_17217);
nor U20141 (N_20141,N_17316,N_18539);
nand U20142 (N_20142,N_18548,N_16980);
nor U20143 (N_20143,N_18307,N_19843);
nand U20144 (N_20144,N_16924,N_16572);
and U20145 (N_20145,N_19506,N_18530);
nor U20146 (N_20146,N_15818,N_18763);
nor U20147 (N_20147,N_19555,N_16566);
xor U20148 (N_20148,N_15303,N_15753);
nor U20149 (N_20149,N_17050,N_16471);
or U20150 (N_20150,N_18797,N_16725);
nor U20151 (N_20151,N_16763,N_17480);
or U20152 (N_20152,N_17115,N_19257);
and U20153 (N_20153,N_17559,N_18477);
xor U20154 (N_20154,N_17101,N_16741);
and U20155 (N_20155,N_15870,N_19087);
xor U20156 (N_20156,N_15125,N_16047);
or U20157 (N_20157,N_15639,N_15791);
and U20158 (N_20158,N_18264,N_16512);
nand U20159 (N_20159,N_19419,N_18297);
nor U20160 (N_20160,N_15088,N_18331);
xnor U20161 (N_20161,N_16291,N_17589);
nor U20162 (N_20162,N_18145,N_16839);
or U20163 (N_20163,N_17192,N_15017);
or U20164 (N_20164,N_15792,N_16811);
xor U20165 (N_20165,N_18518,N_18730);
or U20166 (N_20166,N_15140,N_18085);
nand U20167 (N_20167,N_15151,N_17520);
xnor U20168 (N_20168,N_17849,N_16620);
nand U20169 (N_20169,N_19861,N_18577);
and U20170 (N_20170,N_19244,N_19241);
nand U20171 (N_20171,N_17249,N_17054);
nor U20172 (N_20172,N_15710,N_15065);
and U20173 (N_20173,N_16434,N_16878);
or U20174 (N_20174,N_19362,N_16598);
nor U20175 (N_20175,N_18524,N_15019);
nor U20176 (N_20176,N_18126,N_19957);
nand U20177 (N_20177,N_18314,N_15533);
xor U20178 (N_20178,N_18423,N_17084);
and U20179 (N_20179,N_16894,N_16752);
nand U20180 (N_20180,N_15555,N_19204);
xor U20181 (N_20181,N_17656,N_17838);
nor U20182 (N_20182,N_19088,N_16149);
nor U20183 (N_20183,N_17129,N_15682);
and U20184 (N_20184,N_19045,N_16626);
and U20185 (N_20185,N_18923,N_18289);
and U20186 (N_20186,N_18727,N_19381);
or U20187 (N_20187,N_19900,N_16938);
xor U20188 (N_20188,N_15838,N_15990);
or U20189 (N_20189,N_15529,N_17161);
or U20190 (N_20190,N_17484,N_17706);
and U20191 (N_20191,N_17374,N_15026);
and U20192 (N_20192,N_16562,N_17756);
nor U20193 (N_20193,N_18336,N_18669);
and U20194 (N_20194,N_17677,N_16852);
nand U20195 (N_20195,N_16380,N_19410);
xnor U20196 (N_20196,N_15324,N_15867);
xnor U20197 (N_20197,N_18228,N_17426);
nand U20198 (N_20198,N_19779,N_16925);
nand U20199 (N_20199,N_17699,N_15335);
xor U20200 (N_20200,N_17200,N_18728);
xnor U20201 (N_20201,N_19254,N_16390);
or U20202 (N_20202,N_17670,N_19064);
or U20203 (N_20203,N_16999,N_18924);
xor U20204 (N_20204,N_16996,N_19968);
xnor U20205 (N_20205,N_19668,N_16001);
xor U20206 (N_20206,N_16729,N_18664);
nor U20207 (N_20207,N_17303,N_15231);
or U20208 (N_20208,N_15517,N_18067);
xor U20209 (N_20209,N_17332,N_19021);
xor U20210 (N_20210,N_17860,N_19748);
or U20211 (N_20211,N_16640,N_15013);
or U20212 (N_20212,N_18592,N_15413);
xnor U20213 (N_20213,N_19136,N_17861);
and U20214 (N_20214,N_16644,N_18213);
nor U20215 (N_20215,N_17820,N_19646);
and U20216 (N_20216,N_18967,N_16102);
or U20217 (N_20217,N_16025,N_17736);
or U20218 (N_20218,N_18507,N_19182);
nand U20219 (N_20219,N_18113,N_17333);
xnor U20220 (N_20220,N_16257,N_16085);
nor U20221 (N_20221,N_16319,N_17328);
and U20222 (N_20222,N_16246,N_17452);
nor U20223 (N_20223,N_19191,N_19542);
or U20224 (N_20224,N_16293,N_17956);
and U20225 (N_20225,N_19421,N_15814);
xor U20226 (N_20226,N_18115,N_19527);
xnor U20227 (N_20227,N_17154,N_15477);
nor U20228 (N_20228,N_15492,N_16856);
or U20229 (N_20229,N_18443,N_19415);
nand U20230 (N_20230,N_17329,N_17319);
and U20231 (N_20231,N_18916,N_18288);
and U20232 (N_20232,N_18855,N_18357);
or U20233 (N_20233,N_17814,N_15044);
or U20234 (N_20234,N_16618,N_15558);
xnor U20235 (N_20235,N_15421,N_15074);
and U20236 (N_20236,N_19418,N_17228);
and U20237 (N_20237,N_15581,N_17761);
nor U20238 (N_20238,N_16477,N_15728);
nand U20239 (N_20239,N_16897,N_18769);
nand U20240 (N_20240,N_16579,N_19304);
nor U20241 (N_20241,N_15207,N_17932);
nand U20242 (N_20242,N_19372,N_18322);
nor U20243 (N_20243,N_18223,N_16711);
xnor U20244 (N_20244,N_18915,N_19909);
or U20245 (N_20245,N_17998,N_15197);
and U20246 (N_20246,N_15905,N_17792);
xnor U20247 (N_20247,N_15702,N_16942);
and U20248 (N_20248,N_16636,N_15613);
xnor U20249 (N_20249,N_19086,N_16099);
xnor U20250 (N_20250,N_19816,N_16867);
or U20251 (N_20251,N_18161,N_17807);
nand U20252 (N_20252,N_18034,N_15009);
nor U20253 (N_20253,N_19120,N_19451);
and U20254 (N_20254,N_15935,N_16128);
xnor U20255 (N_20255,N_16219,N_19890);
or U20256 (N_20256,N_17810,N_18472);
nor U20257 (N_20257,N_18792,N_15766);
nor U20258 (N_20258,N_17816,N_17953);
nand U20259 (N_20259,N_18688,N_17781);
nand U20260 (N_20260,N_17850,N_16408);
or U20261 (N_20261,N_15946,N_16454);
or U20262 (N_20262,N_18546,N_19920);
nor U20263 (N_20263,N_17270,N_18461);
or U20264 (N_20264,N_19509,N_19276);
nand U20265 (N_20265,N_16538,N_19467);
and U20266 (N_20266,N_16709,N_15350);
xnor U20267 (N_20267,N_19007,N_18579);
nor U20268 (N_20268,N_19279,N_17984);
or U20269 (N_20269,N_15055,N_16916);
xnor U20270 (N_20270,N_19343,N_16202);
or U20271 (N_20271,N_16922,N_17620);
nand U20272 (N_20272,N_18258,N_19960);
nand U20273 (N_20273,N_18456,N_19489);
and U20274 (N_20274,N_18717,N_17272);
or U20275 (N_20275,N_19301,N_19867);
xor U20276 (N_20276,N_19565,N_16669);
nand U20277 (N_20277,N_18771,N_17058);
nand U20278 (N_20278,N_17571,N_19863);
and U20279 (N_20279,N_15208,N_16059);
nor U20280 (N_20280,N_19056,N_18144);
xnor U20281 (N_20281,N_19698,N_16391);
or U20282 (N_20282,N_18471,N_15569);
xor U20283 (N_20283,N_19164,N_15451);
or U20284 (N_20284,N_16487,N_16815);
xnor U20285 (N_20285,N_16284,N_19036);
xnor U20286 (N_20286,N_17920,N_17392);
or U20287 (N_20287,N_16420,N_18045);
or U20288 (N_20288,N_17539,N_17411);
xor U20289 (N_20289,N_16882,N_15337);
nand U20290 (N_20290,N_19393,N_16870);
nand U20291 (N_20291,N_15582,N_16675);
and U20292 (N_20292,N_16608,N_17751);
and U20293 (N_20293,N_18062,N_19777);
nand U20294 (N_20294,N_18398,N_15837);
xor U20295 (N_20295,N_19070,N_19434);
or U20296 (N_20296,N_15886,N_19993);
and U20297 (N_20297,N_15104,N_19659);
nand U20298 (N_20298,N_18832,N_17650);
and U20299 (N_20299,N_17443,N_18180);
nand U20300 (N_20300,N_16968,N_18553);
or U20301 (N_20301,N_15704,N_15276);
nor U20302 (N_20302,N_18948,N_18463);
nor U20303 (N_20303,N_15651,N_17691);
xnor U20304 (N_20304,N_18774,N_16414);
nand U20305 (N_20305,N_15857,N_19761);
or U20306 (N_20306,N_19835,N_17967);
or U20307 (N_20307,N_16145,N_18533);
nor U20308 (N_20308,N_17186,N_17408);
and U20309 (N_20309,N_15866,N_16819);
or U20310 (N_20310,N_15745,N_17176);
nand U20311 (N_20311,N_15800,N_16162);
and U20312 (N_20312,N_18110,N_16966);
nand U20313 (N_20313,N_19709,N_19534);
and U20314 (N_20314,N_17466,N_16229);
xnor U20315 (N_20315,N_19980,N_17720);
or U20316 (N_20316,N_15306,N_15621);
and U20317 (N_20317,N_15841,N_18584);
and U20318 (N_20318,N_18284,N_15157);
and U20319 (N_20319,N_17259,N_17899);
and U20320 (N_20320,N_16273,N_18615);
and U20321 (N_20321,N_19445,N_17105);
or U20322 (N_20322,N_16652,N_18775);
or U20323 (N_20323,N_18773,N_19212);
or U20324 (N_20324,N_18057,N_18961);
and U20325 (N_20325,N_16252,N_17640);
xnor U20326 (N_20326,N_16724,N_17774);
and U20327 (N_20327,N_15077,N_15395);
nor U20328 (N_20328,N_19773,N_17870);
nor U20329 (N_20329,N_19610,N_17025);
nand U20330 (N_20330,N_18060,N_16045);
nor U20331 (N_20331,N_19268,N_15115);
nand U20332 (N_20332,N_16207,N_15915);
xor U20333 (N_20333,N_15747,N_16713);
or U20334 (N_20334,N_15992,N_17738);
xor U20335 (N_20335,N_16525,N_17930);
or U20336 (N_20336,N_16854,N_17937);
or U20337 (N_20337,N_17499,N_16733);
or U20338 (N_20338,N_15251,N_17951);
xnor U20339 (N_20339,N_18070,N_16714);
nand U20340 (N_20340,N_18016,N_17618);
xnor U20341 (N_20341,N_15287,N_15833);
or U20342 (N_20342,N_18960,N_16998);
xnor U20343 (N_20343,N_17927,N_18785);
nand U20344 (N_20344,N_19195,N_17241);
xnor U20345 (N_20345,N_17087,N_18493);
xor U20346 (N_20346,N_17045,N_19133);
nor U20347 (N_20347,N_19047,N_16197);
nor U20348 (N_20348,N_18385,N_15811);
or U20349 (N_20349,N_16710,N_15887);
nor U20350 (N_20350,N_18140,N_18515);
and U20351 (N_20351,N_18358,N_18295);
and U20352 (N_20352,N_18901,N_19126);
xnor U20353 (N_20353,N_16090,N_19223);
nor U20354 (N_20354,N_16169,N_19002);
nor U20355 (N_20355,N_18600,N_16032);
or U20356 (N_20356,N_19597,N_18343);
xnor U20357 (N_20357,N_16294,N_17240);
nor U20358 (N_20358,N_19173,N_18977);
or U20359 (N_20359,N_18222,N_18393);
or U20360 (N_20360,N_16198,N_19821);
nand U20361 (N_20361,N_18601,N_15354);
nand U20362 (N_20362,N_17795,N_15427);
or U20363 (N_20363,N_15038,N_19132);
nor U20364 (N_20364,N_16798,N_16952);
nor U20365 (N_20365,N_17788,N_17331);
and U20366 (N_20366,N_15902,N_15076);
or U20367 (N_20367,N_19385,N_16276);
xor U20368 (N_20368,N_16480,N_17726);
xnor U20369 (N_20369,N_18788,N_15945);
or U20370 (N_20370,N_17724,N_19953);
and U20371 (N_20371,N_16504,N_15048);
or U20372 (N_20372,N_18325,N_18912);
and U20373 (N_20373,N_19731,N_18469);
nand U20374 (N_20374,N_15764,N_16835);
nor U20375 (N_20375,N_17223,N_15974);
nand U20376 (N_20376,N_17199,N_17421);
nor U20377 (N_20377,N_15921,N_18849);
xnor U20378 (N_20378,N_15333,N_17409);
xnor U20379 (N_20379,N_15729,N_16437);
or U20380 (N_20380,N_17302,N_19251);
or U20381 (N_20381,N_17271,N_19152);
nand U20382 (N_20382,N_18027,N_17349);
nor U20383 (N_20383,N_18913,N_16795);
and U20384 (N_20384,N_15183,N_17958);
nand U20385 (N_20385,N_17455,N_16774);
and U20386 (N_20386,N_16780,N_16935);
nor U20387 (N_20387,N_15860,N_18277);
nand U20388 (N_20388,N_18652,N_17626);
nand U20389 (N_20389,N_18294,N_19949);
and U20390 (N_20390,N_19762,N_16921);
and U20391 (N_20391,N_18316,N_16425);
nor U20392 (N_20392,N_18704,N_19130);
and U20393 (N_20393,N_15969,N_17026);
nor U20394 (N_20394,N_17008,N_17378);
xor U20395 (N_20395,N_16413,N_16340);
or U20396 (N_20396,N_17423,N_16370);
nor U20397 (N_20397,N_18430,N_16311);
nand U20398 (N_20398,N_15603,N_16289);
or U20399 (N_20399,N_15202,N_15561);
nor U20400 (N_20400,N_16301,N_15808);
and U20401 (N_20401,N_19876,N_15265);
and U20402 (N_20402,N_17195,N_19976);
or U20403 (N_20403,N_19881,N_17030);
xor U20404 (N_20404,N_19101,N_17352);
nor U20405 (N_20405,N_16175,N_17024);
and U20406 (N_20406,N_15005,N_16961);
xnor U20407 (N_20407,N_18829,N_15593);
nand U20408 (N_20408,N_17778,N_19540);
and U20409 (N_20409,N_16558,N_18587);
or U20410 (N_20410,N_15635,N_17918);
xor U20411 (N_20411,N_18899,N_15173);
nor U20412 (N_20412,N_16352,N_17086);
and U20413 (N_20413,N_18966,N_18473);
nand U20414 (N_20414,N_17622,N_18607);
or U20415 (N_20415,N_15378,N_18640);
or U20416 (N_20416,N_15217,N_17363);
xor U20417 (N_20417,N_16786,N_19739);
nor U20418 (N_20418,N_18011,N_18002);
or U20419 (N_20419,N_15431,N_15685);
and U20420 (N_20420,N_15093,N_18361);
or U20421 (N_20421,N_18189,N_16723);
nor U20422 (N_20422,N_16770,N_18382);
or U20423 (N_20423,N_18138,N_19750);
nand U20424 (N_20424,N_19334,N_17554);
or U20425 (N_20425,N_15219,N_19083);
xnor U20426 (N_20426,N_18235,N_15781);
nor U20427 (N_20427,N_17878,N_15135);
nand U20428 (N_20428,N_17880,N_18729);
xnor U20429 (N_20429,N_16179,N_18190);
nor U20430 (N_20430,N_16078,N_15212);
nand U20431 (N_20431,N_18362,N_15632);
nand U20432 (N_20432,N_18981,N_16106);
nand U20433 (N_20433,N_18862,N_17483);
nand U20434 (N_20434,N_15918,N_17887);
xor U20435 (N_20435,N_18187,N_19884);
xor U20436 (N_20436,N_19977,N_17966);
xnor U20437 (N_20437,N_15999,N_15756);
nor U20438 (N_20438,N_19482,N_17601);
nor U20439 (N_20439,N_18203,N_18687);
or U20440 (N_20440,N_19903,N_16893);
nor U20441 (N_20441,N_15986,N_16234);
or U20442 (N_20442,N_16325,N_19231);
nand U20443 (N_20443,N_16242,N_17311);
or U20444 (N_20444,N_17658,N_17822);
and U20445 (N_20445,N_16407,N_15723);
and U20446 (N_20446,N_19644,N_16270);
and U20447 (N_20447,N_16123,N_18135);
and U20448 (N_20448,N_17447,N_17661);
or U20449 (N_20449,N_16737,N_19171);
xnor U20450 (N_20450,N_18697,N_16688);
nand U20451 (N_20451,N_18685,N_19726);
nand U20452 (N_20452,N_19472,N_17401);
xnor U20453 (N_20453,N_17858,N_15272);
nand U20454 (N_20454,N_15379,N_16643);
and U20455 (N_20455,N_19433,N_19662);
nand U20456 (N_20456,N_16528,N_18291);
nor U20457 (N_20457,N_17555,N_17644);
xor U20458 (N_20458,N_17624,N_18158);
nor U20459 (N_20459,N_16842,N_19965);
nand U20460 (N_20460,N_19759,N_16662);
nand U20461 (N_20461,N_15130,N_18675);
xnor U20462 (N_20462,N_17659,N_18875);
nand U20463 (N_20463,N_19775,N_15479);
xnor U20464 (N_20464,N_15942,N_19933);
and U20465 (N_20465,N_18460,N_15317);
nand U20466 (N_20466,N_19669,N_19714);
and U20467 (N_20467,N_15977,N_17204);
nor U20468 (N_20468,N_15973,N_18486);
nor U20469 (N_20469,N_18596,N_18479);
nor U20470 (N_20470,N_19785,N_19066);
or U20471 (N_20471,N_17296,N_16576);
and U20472 (N_20472,N_15608,N_17596);
nor U20473 (N_20473,N_18990,N_18815);
nand U20474 (N_20474,N_17145,N_19655);
and U20475 (N_20475,N_15778,N_16718);
nand U20476 (N_20476,N_15813,N_19295);
and U20477 (N_20477,N_19742,N_16986);
nor U20478 (N_20478,N_19062,N_15996);
nand U20479 (N_20479,N_16153,N_17244);
and U20480 (N_20480,N_15404,N_16762);
xnor U20481 (N_20481,N_15678,N_19671);
or U20482 (N_20482,N_18510,N_15402);
xor U20483 (N_20483,N_17078,N_17638);
or U20484 (N_20484,N_19494,N_18928);
or U20485 (N_20485,N_17356,N_15178);
nor U20486 (N_20486,N_18993,N_15615);
or U20487 (N_20487,N_19262,N_18561);
xnor U20488 (N_20488,N_16611,N_18588);
and U20489 (N_20489,N_15757,N_16540);
or U20490 (N_20490,N_18433,N_15136);
nor U20491 (N_20491,N_15836,N_19973);
xor U20492 (N_20492,N_15062,N_17654);
nor U20493 (N_20493,N_17245,N_17063);
nand U20494 (N_20494,N_15732,N_19134);
nor U20495 (N_20495,N_18455,N_17572);
and U20496 (N_20496,N_18597,N_16868);
xnor U20497 (N_20497,N_15116,N_17742);
xnor U20498 (N_20498,N_19844,N_18129);
or U20499 (N_20499,N_17373,N_16641);
or U20500 (N_20500,N_17564,N_17614);
or U20501 (N_20501,N_19225,N_17915);
nand U20502 (N_20502,N_17741,N_15480);
xor U20503 (N_20503,N_16707,N_18929);
or U20504 (N_20504,N_15290,N_16628);
or U20505 (N_20505,N_16672,N_18655);
and U20506 (N_20506,N_19567,N_15364);
or U20507 (N_20507,N_18256,N_19353);
nand U20508 (N_20508,N_17800,N_19590);
xnor U20509 (N_20509,N_19298,N_17364);
nor U20510 (N_20510,N_18242,N_16989);
xor U20511 (N_20511,N_16549,N_15798);
and U20512 (N_20512,N_18448,N_16561);
nor U20513 (N_20513,N_18866,N_18893);
nor U20514 (N_20514,N_19289,N_16631);
xnor U20515 (N_20515,N_19480,N_16112);
or U20516 (N_20516,N_17926,N_18660);
nor U20517 (N_20517,N_16365,N_17750);
and U20518 (N_20518,N_19598,N_17504);
xnor U20519 (N_20519,N_18851,N_18885);
nand U20520 (N_20520,N_19730,N_15474);
xor U20521 (N_20521,N_16847,N_16326);
nand U20522 (N_20522,N_15770,N_19615);
xnor U20523 (N_20523,N_15663,N_15940);
or U20524 (N_20524,N_18425,N_15114);
and U20525 (N_20525,N_18565,N_19397);
nor U20526 (N_20526,N_18079,N_15295);
nor U20527 (N_20527,N_17921,N_18552);
nand U20528 (N_20528,N_16165,N_16739);
nand U20529 (N_20529,N_15235,N_19364);
nand U20530 (N_20530,N_17188,N_19899);
nor U20531 (N_20531,N_19190,N_16485);
and U20532 (N_20532,N_15232,N_16985);
xor U20533 (N_20533,N_19336,N_17289);
and U20534 (N_20534,N_17570,N_15282);
or U20535 (N_20535,N_19766,N_19280);
nor U20536 (N_20536,N_19074,N_19197);
nor U20537 (N_20537,N_17548,N_18676);
xnor U20538 (N_20538,N_16350,N_18630);
nand U20539 (N_20539,N_15845,N_15768);
and U20540 (N_20540,N_18273,N_16764);
and U20541 (N_20541,N_17684,N_17287);
xnor U20542 (N_20542,N_16262,N_19864);
or U20543 (N_20543,N_18644,N_15662);
xnor U20544 (N_20544,N_19586,N_19915);
and U20545 (N_20545,N_19009,N_18994);
nor U20546 (N_20546,N_18104,N_16185);
xnor U20547 (N_20547,N_18467,N_19384);
or U20548 (N_20548,N_16472,N_16143);
nor U20549 (N_20549,N_18279,N_17317);
xnor U20550 (N_20550,N_17039,N_18483);
nand U20551 (N_20551,N_19717,N_16670);
xnor U20552 (N_20552,N_15047,N_15885);
xor U20553 (N_20553,N_18397,N_18877);
or U20554 (N_20554,N_18714,N_15266);
and U20555 (N_20555,N_18547,N_19210);
nor U20556 (N_20556,N_16183,N_16049);
xor U20557 (N_20557,N_17728,N_16954);
xor U20558 (N_20558,N_16695,N_16969);
or U20559 (N_20559,N_17236,N_19441);
and U20560 (N_20560,N_18853,N_19389);
and U20561 (N_20561,N_18283,N_16138);
xor U20562 (N_20562,N_19077,N_17082);
nor U20563 (N_20563,N_15388,N_18538);
xnor U20564 (N_20564,N_16804,N_19379);
nand U20565 (N_20565,N_15976,N_16605);
xnor U20566 (N_20566,N_15171,N_15527);
nor U20567 (N_20567,N_18069,N_17264);
and U20568 (N_20568,N_18209,N_18904);
xnor U20569 (N_20569,N_16544,N_17168);
xnor U20570 (N_20570,N_15283,N_15929);
nand U20571 (N_20571,N_19570,N_18986);
xnor U20572 (N_20572,N_19093,N_16481);
xor U20573 (N_20573,N_15864,N_18305);
xnor U20574 (N_20574,N_17675,N_18193);
and U20575 (N_20575,N_17588,N_15087);
or U20576 (N_20576,N_16318,N_16354);
nand U20577 (N_20577,N_18957,N_19883);
nand U20578 (N_20578,N_16410,N_17293);
xor U20579 (N_20579,N_16865,N_18137);
and U20580 (N_20580,N_18555,N_19549);
and U20581 (N_20581,N_18198,N_17123);
nor U20582 (N_20582,N_18526,N_16678);
xor U20583 (N_20583,N_15066,N_19278);
xnor U20584 (N_20584,N_19214,N_18947);
and U20585 (N_20585,N_15565,N_18072);
or U20586 (N_20586,N_16875,N_19854);
nor U20587 (N_20587,N_18102,N_16424);
nand U20588 (N_20588,N_16016,N_18204);
and U20589 (N_20589,N_18001,N_17465);
xor U20590 (N_20590,N_17089,N_15680);
nor U20591 (N_20591,N_16514,N_15278);
nor U20592 (N_20592,N_16050,N_18976);
or U20593 (N_20593,N_15597,N_17841);
nor U20594 (N_20594,N_16287,N_15422);
or U20595 (N_20595,N_17371,N_18073);
nand U20596 (N_20596,N_16155,N_18557);
and U20597 (N_20597,N_19250,N_16928);
xnor U20598 (N_20598,N_18860,N_15101);
xor U20599 (N_20599,N_17912,N_16406);
or U20600 (N_20600,N_19918,N_17116);
nor U20601 (N_20601,N_19219,N_18999);
and U20602 (N_20602,N_15203,N_16403);
nand U20603 (N_20603,N_16439,N_19029);
and U20604 (N_20604,N_19265,N_19207);
xnor U20605 (N_20605,N_15557,N_19436);
or U20606 (N_20606,N_18241,N_16794);
xnor U20607 (N_20607,N_15199,N_17298);
xor U20608 (N_20608,N_16621,N_18699);
or U20609 (N_20609,N_16656,N_17746);
xnor U20610 (N_20610,N_15172,N_19677);
nand U20611 (N_20611,N_17459,N_18280);
nand U20612 (N_20612,N_15383,N_16396);
nand U20613 (N_20613,N_15650,N_19363);
xor U20614 (N_20614,N_16046,N_19335);
or U20615 (N_20615,N_16523,N_18694);
and U20616 (N_20616,N_16039,N_18569);
or U20617 (N_20617,N_18513,N_16861);
or U20618 (N_20618,N_16266,N_15744);
nand U20619 (N_20619,N_16885,N_15166);
nor U20620 (N_20620,N_18902,N_15222);
nor U20621 (N_20621,N_15606,N_16731);
xor U20622 (N_20622,N_17709,N_15163);
nand U20623 (N_20623,N_15249,N_17764);
or U20624 (N_20624,N_15693,N_19842);
xor U20625 (N_20625,N_16445,N_19652);
nand U20626 (N_20626,N_16453,N_19922);
nor U20627 (N_20627,N_19601,N_19667);
or U20628 (N_20628,N_16984,N_16880);
and U20629 (N_20629,N_16864,N_15616);
nand U20630 (N_20630,N_16750,N_15201);
or U20631 (N_20631,N_17749,N_17703);
and U20632 (N_20632,N_16448,N_17535);
and U20633 (N_20633,N_15975,N_17273);
and U20634 (N_20634,N_17109,N_17079);
and U20635 (N_20635,N_17980,N_15925);
or U20636 (N_20636,N_16778,N_15551);
nor U20637 (N_20637,N_17137,N_16895);
and U20638 (N_20638,N_18647,N_15997);
and U20639 (N_20639,N_16526,N_19650);
nor U20640 (N_20640,N_16557,N_17587);
or U20641 (N_20641,N_16310,N_16511);
nand U20642 (N_20642,N_18342,N_16694);
xor U20643 (N_20643,N_17925,N_18390);
nand U20644 (N_20644,N_19547,N_19181);
and U20645 (N_20645,N_15737,N_15676);
xnor U20646 (N_20646,N_16940,N_16564);
and U20647 (N_20647,N_15742,N_16962);
nor U20648 (N_20648,N_19751,N_16192);
nand U20649 (N_20649,N_15412,N_17102);
nor U20650 (N_20650,N_19432,N_19503);
nor U20651 (N_20651,N_16681,N_18985);
xnor U20652 (N_20652,N_15968,N_16201);
and U20653 (N_20653,N_15679,N_17577);
xor U20654 (N_20654,N_16281,N_18667);
nand U20655 (N_20655,N_17099,N_15007);
xor U20656 (N_20656,N_18465,N_15611);
or U20657 (N_20657,N_17253,N_17695);
or U20658 (N_20658,N_16247,N_19292);
and U20659 (N_20659,N_16345,N_17657);
and U20660 (N_20660,N_18328,N_19490);
nand U20661 (N_20661,N_18619,N_15020);
nor U20662 (N_20662,N_16747,N_16905);
and U20663 (N_20663,N_17765,N_18594);
nand U20664 (N_20664,N_18650,N_18071);
xnor U20665 (N_20665,N_17010,N_15029);
and U20666 (N_20666,N_16483,N_16109);
xor U20667 (N_20667,N_18337,N_15457);
or U20668 (N_20668,N_17645,N_16509);
xnor U20669 (N_20669,N_18738,N_17542);
nand U20670 (N_20670,N_19333,N_18760);
and U20671 (N_20671,N_16506,N_18634);
nand U20672 (N_20672,N_16163,N_15964);
or U20673 (N_20673,N_17384,N_19312);
and U20674 (N_20674,N_18391,N_15351);
nor U20675 (N_20675,N_17138,N_18381);
nand U20676 (N_20676,N_17674,N_19040);
or U20677 (N_20677,N_19868,N_16363);
or U20678 (N_20678,N_16501,N_19018);
nor U20679 (N_20679,N_18946,N_19907);
and U20680 (N_20680,N_17169,N_15152);
or U20681 (N_20681,N_18953,N_18618);
or U20682 (N_20682,N_18852,N_16965);
or U20683 (N_20683,N_19382,N_18633);
nor U20684 (N_20684,N_16324,N_18840);
xnor U20685 (N_20685,N_17760,N_15966);
nor U20686 (N_20686,N_18514,N_19702);
and U20687 (N_20687,N_18310,N_19995);
nand U20688 (N_20688,N_18686,N_15668);
nand U20689 (N_20689,N_16232,N_18827);
xor U20690 (N_20690,N_15442,N_15141);
nand U20691 (N_20691,N_15755,N_15535);
nor U20692 (N_20692,N_16343,N_19311);
or U20693 (N_20693,N_18881,N_18431);
or U20694 (N_20694,N_19255,N_17255);
xor U20695 (N_20695,N_17237,N_15478);
or U20696 (N_20696,N_16634,N_15826);
xnor U20697 (N_20697,N_15854,N_16404);
nand U20698 (N_20698,N_18534,N_15705);
nor U20699 (N_20699,N_15191,N_19896);
xnor U20700 (N_20700,N_15629,N_16239);
nand U20701 (N_20701,N_15079,N_19521);
and U20702 (N_20702,N_16328,N_15503);
xnor U20703 (N_20703,N_16158,N_18653);
nor U20704 (N_20704,N_19430,N_15499);
nor U20705 (N_20705,N_16676,N_17689);
or U20706 (N_20706,N_17615,N_17177);
and U20707 (N_20707,N_15806,N_19216);
xor U20708 (N_20708,N_15530,N_19656);
or U20709 (N_20709,N_17693,N_18217);
or U20710 (N_20710,N_19638,N_15456);
xnor U20711 (N_20711,N_18502,N_17471);
nand U20712 (N_20712,N_18932,N_17246);
nand U20713 (N_20713,N_19319,N_16196);
nor U20714 (N_20714,N_18925,N_15100);
nor U20715 (N_20715,N_15699,N_17687);
nand U20716 (N_20716,N_15985,N_18648);
nand U20717 (N_20717,N_16248,N_18927);
nand U20718 (N_20718,N_17182,N_15750);
xnor U20719 (N_20719,N_16029,N_17595);
xor U20720 (N_20720,N_18749,N_17583);
and U20721 (N_20721,N_16953,N_16958);
xor U20722 (N_20722,N_19528,N_19693);
or U20723 (N_20723,N_19004,N_17042);
nand U20724 (N_20724,N_17939,N_19478);
xnor U20725 (N_20725,N_16508,N_15630);
nor U20726 (N_20726,N_17609,N_17651);
nor U20727 (N_20727,N_17673,N_15109);
xnor U20728 (N_20728,N_18870,N_18890);
or U20729 (N_20729,N_17785,N_16686);
and U20730 (N_20730,N_17057,N_16467);
or U20731 (N_20731,N_16701,N_16462);
nand U20732 (N_20732,N_19860,N_19053);
or U20733 (N_20733,N_19205,N_19180);
nand U20734 (N_20734,N_17441,N_17478);
nand U20735 (N_20735,N_17388,N_19847);
xor U20736 (N_20736,N_15901,N_16858);
or U20737 (N_20737,N_15592,N_16992);
and U20738 (N_20738,N_17619,N_16323);
xnor U20739 (N_20739,N_16210,N_19371);
and U20740 (N_20740,N_17773,N_18543);
or U20741 (N_20741,N_18542,N_16011);
nor U20742 (N_20742,N_19167,N_18892);
or U20743 (N_20743,N_18311,N_18971);
xor U20744 (N_20744,N_17098,N_17081);
nand U20745 (N_20745,N_15453,N_19772);
and U20746 (N_20746,N_16091,N_18370);
or U20747 (N_20747,N_18949,N_16189);
nand U20748 (N_20748,N_19605,N_18225);
nor U20749 (N_20749,N_17683,N_16451);
xnor U20750 (N_20750,N_18649,N_18639);
nand U20751 (N_20751,N_17140,N_15855);
or U20752 (N_20752,N_18263,N_16693);
and U20753 (N_20753,N_17429,N_15532);
nor U20754 (N_20754,N_17107,N_17610);
nor U20755 (N_20755,N_19648,N_17865);
nand U20756 (N_20756,N_17630,N_15339);
and U20757 (N_20757,N_19706,N_15086);
nor U20758 (N_20758,N_19782,N_17533);
and U20759 (N_20759,N_19753,N_16320);
xor U20760 (N_20760,N_16455,N_19765);
nand U20761 (N_20761,N_16087,N_19249);
nor U20762 (N_20762,N_18713,N_19628);
nand U20763 (N_20763,N_17666,N_15575);
and U20764 (N_20764,N_17929,N_15016);
nor U20765 (N_20765,N_16386,N_18312);
and U20766 (N_20766,N_15910,N_17872);
and U20767 (N_20767,N_19979,N_18260);
or U20768 (N_20768,N_17671,N_17336);
or U20769 (N_20769,N_15708,N_18681);
or U20770 (N_20770,N_16913,N_17961);
and U20771 (N_20771,N_17386,N_18368);
xor U20772 (N_20772,N_16012,N_16758);
and U20773 (N_20773,N_19183,N_15659);
nand U20774 (N_20774,N_18613,N_16405);
and U20775 (N_20775,N_15312,N_19982);
or U20776 (N_20776,N_17708,N_17495);
nor U20777 (N_20777,N_15161,N_16917);
or U20778 (N_20778,N_19634,N_16156);
nand U20779 (N_20779,N_15297,N_19935);
and U20780 (N_20780,N_15146,N_19906);
and U20781 (N_20781,N_18848,N_16037);
xnor U20782 (N_20782,N_17797,N_19008);
nor U20783 (N_20783,N_15928,N_15268);
and U20784 (N_20784,N_17836,N_15835);
nand U20785 (N_20785,N_17983,N_16682);
nand U20786 (N_20786,N_17648,N_17442);
nor U20787 (N_20787,N_15684,N_16660);
or U20788 (N_20788,N_15822,N_19135);
nor U20789 (N_20789,N_16421,N_18369);
xor U20790 (N_20790,N_19676,N_17970);
or U20791 (N_20791,N_16178,N_15807);
nand U20792 (N_20792,N_16020,N_17474);
nand U20793 (N_20793,N_19678,N_19872);
nor U20794 (N_20794,N_16080,N_19701);
or U20795 (N_20795,N_19038,N_18481);
or U20796 (N_20796,N_16374,N_17283);
nand U20797 (N_20797,N_19585,N_15286);
nand U20798 (N_20798,N_15549,N_17565);
or U20799 (N_20799,N_18747,N_15718);
xor U20800 (N_20800,N_17593,N_16253);
nor U20801 (N_20801,N_17381,N_19734);
nand U20802 (N_20802,N_17826,N_15550);
xnor U20803 (N_20803,N_17833,N_16700);
and U20804 (N_20804,N_18835,N_15243);
nand U20805 (N_20805,N_15957,N_17602);
nand U20806 (N_20806,N_19006,N_16100);
nand U20807 (N_20807,N_17541,N_15979);
xnor U20808 (N_20808,N_18367,N_18136);
xor U20809 (N_20809,N_19530,N_19458);
xnor U20810 (N_20810,N_17404,N_17509);
xnor U20811 (N_20811,N_16236,N_17649);
nor U20812 (N_20812,N_16068,N_17162);
xor U20813 (N_20813,N_19518,N_15541);
or U20814 (N_20814,N_19522,N_18380);
nand U20815 (N_20815,N_18012,N_18188);
xor U20816 (N_20816,N_19787,N_18334);
nand U20817 (N_20817,N_16879,N_17514);
or U20818 (N_20818,N_19846,N_16302);
and U20819 (N_20819,N_17007,N_17029);
nand U20820 (N_20820,N_18883,N_16375);
xor U20821 (N_20821,N_19339,N_15600);
or U20822 (N_20822,N_18451,N_16152);
nand U20823 (N_20823,N_18445,N_18048);
nand U20824 (N_20824,N_15142,N_17448);
and U20825 (N_20825,N_15884,N_19768);
nand U20826 (N_20826,N_19893,N_19501);
nor U20827 (N_20827,N_16353,N_18030);
nor U20828 (N_20828,N_16136,N_17536);
or U20829 (N_20829,N_16226,N_19635);
nor U20830 (N_20830,N_17672,N_17906);
or U20831 (N_20831,N_15285,N_17598);
nor U20832 (N_20832,N_19096,N_19095);
nor U20833 (N_20833,N_15057,N_19037);
xor U20834 (N_20834,N_15343,N_16048);
nand U20835 (N_20835,N_17938,N_16015);
xnor U20836 (N_20836,N_16677,N_19222);
or U20837 (N_20837,N_16397,N_18024);
or U20838 (N_20838,N_15033,N_16157);
or U20839 (N_20839,N_19721,N_16217);
nor U20840 (N_20840,N_17231,N_17900);
or U20841 (N_20841,N_15170,N_16161);
or U20842 (N_20842,N_18672,N_18003);
xor U20843 (N_20843,N_16837,N_15126);
nand U20844 (N_20844,N_19981,N_16098);
and U20845 (N_20845,N_17150,N_17324);
and U20846 (N_20846,N_18097,N_17094);
nor U20847 (N_20847,N_19654,N_17635);
and U20848 (N_20848,N_16329,N_15840);
xnor U20849 (N_20849,N_15433,N_16125);
or U20850 (N_20850,N_19465,N_15559);
nand U20851 (N_20851,N_17890,N_19636);
xnor U20852 (N_20852,N_17412,N_18109);
nand U20853 (N_20853,N_18440,N_19321);
or U20854 (N_20854,N_19035,N_16590);
xnor U20855 (N_20855,N_15959,N_18230);
nor U20856 (N_20856,N_17719,N_16520);
xor U20857 (N_20857,N_16010,N_19887);
nand U20858 (N_20858,N_17972,N_17846);
or U20859 (N_20859,N_18700,N_16496);
nand U20860 (N_20860,N_17419,N_16019);
nand U20861 (N_20861,N_18780,N_15024);
nand U20862 (N_20862,N_16053,N_15103);
and U20863 (N_20863,N_16315,N_17784);
xnor U20864 (N_20864,N_18268,N_17859);
or U20865 (N_20865,N_15396,N_17574);
or U20866 (N_20866,N_18192,N_17507);
or U20867 (N_20867,N_18152,N_15252);
nor U20868 (N_20868,N_17558,N_16077);
nor U20869 (N_20869,N_17144,N_19733);
nor U20870 (N_20870,N_16831,N_18179);
and U20871 (N_20871,N_16591,N_15701);
nor U20872 (N_20872,N_19461,N_18360);
and U20873 (N_20873,N_17346,N_17438);
nor U20874 (N_20874,N_15188,N_17286);
nand U20875 (N_20875,N_19215,N_15240);
nand U20876 (N_20876,N_19404,N_17889);
or U20877 (N_20877,N_18078,N_15673);
and U20878 (N_20878,N_16022,N_19532);
nand U20879 (N_20879,N_19849,N_18111);
xor U20880 (N_20880,N_19902,N_15323);
xor U20881 (N_20881,N_17639,N_18726);
nand U20882 (N_20882,N_19402,N_15785);
nor U20883 (N_20883,N_18436,N_19448);
nand U20884 (N_20884,N_19131,N_18014);
nand U20885 (N_20885,N_17376,N_17059);
xor U20886 (N_20886,N_16459,N_19237);
nand U20887 (N_20887,N_17470,N_17325);
nand U20888 (N_20888,N_19629,N_19199);
or U20889 (N_20889,N_16009,N_19329);
and U20890 (N_20890,N_17599,N_15061);
xor U20891 (N_20891,N_19141,N_19780);
nand U20892 (N_20892,N_18076,N_18153);
xor U20893 (N_20893,N_16460,N_18991);
and U20894 (N_20894,N_19300,N_16474);
and U20895 (N_20895,N_18501,N_18563);
nand U20896 (N_20896,N_15720,N_19356);
and U20897 (N_20897,N_15440,N_16991);
nand U20898 (N_20898,N_18405,N_16027);
or U20899 (N_20899,N_18909,N_15776);
or U20900 (N_20900,N_17458,N_18889);
nor U20901 (N_20901,N_17933,N_18703);
xor U20902 (N_20902,N_16181,N_18459);
nand U20903 (N_20903,N_16560,N_17205);
nand U20904 (N_20904,N_18374,N_16255);
nor U20905 (N_20905,N_18559,N_18603);
and U20906 (N_20906,N_15362,N_15176);
xor U20907 (N_20907,N_19187,N_18419);
nand U20908 (N_20908,N_19687,N_18781);
nand U20909 (N_20909,N_17667,N_17268);
xor U20910 (N_20910,N_17125,N_18941);
nor U20911 (N_20911,N_17819,N_15181);
or U20912 (N_20912,N_18591,N_16042);
nor U20913 (N_20913,N_16108,N_16507);
nor U20914 (N_20914,N_17267,N_17403);
xnor U20915 (N_20915,N_18000,N_15578);
nor U20916 (N_20916,N_18417,N_15332);
nand U20917 (N_20917,N_19855,N_19235);
nor U20918 (N_20918,N_15687,N_16184);
or U20919 (N_20919,N_16663,N_19228);
xor U20920 (N_20920,N_15483,N_18789);
or U20921 (N_20921,N_17790,N_17354);
nand U20922 (N_20922,N_15145,N_19637);
xnor U20923 (N_20923,N_15824,N_15912);
and U20924 (N_20924,N_17433,N_17989);
xnor U20925 (N_20925,N_19431,N_15733);
nand U20926 (N_20926,N_19079,N_18013);
or U20927 (N_20927,N_17942,N_19168);
or U20928 (N_20928,N_18776,N_15512);
or U20929 (N_20929,N_19561,N_18721);
nor U20930 (N_20930,N_16431,N_15526);
nor U20931 (N_20931,N_17183,N_19614);
nand U20932 (N_20932,N_17147,N_17340);
xor U20933 (N_20933,N_19529,N_17576);
xor U20934 (N_20934,N_17941,N_18616);
xnor U20935 (N_20935,N_19229,N_16862);
nand U20936 (N_20936,N_16195,N_16630);
nor U20937 (N_20937,N_19836,N_17992);
and U20938 (N_20938,N_15468,N_19493);
or U20939 (N_20939,N_19455,N_15417);
or U20940 (N_20940,N_18651,N_16299);
and U20941 (N_20941,N_17124,N_18165);
and U20942 (N_20942,N_18017,N_17830);
nor U20943 (N_20943,N_16013,N_19865);
and U20944 (N_20944,N_16568,N_17126);
xnor U20945 (N_20945,N_15947,N_18575);
nand U20946 (N_20946,N_15043,N_15298);
nor U20947 (N_20947,N_17234,N_19063);
xor U20948 (N_20948,N_17862,N_16651);
and U20949 (N_20949,N_17417,N_19429);
or U20950 (N_20950,N_18441,N_15491);
xnor U20951 (N_20951,N_17968,N_15774);
or U20952 (N_20952,N_16290,N_15186);
and U20953 (N_20953,N_18505,N_16124);
nor U20954 (N_20954,N_18098,N_15511);
nor U20955 (N_20955,N_18807,N_16449);
or U20956 (N_20956,N_16661,N_19552);
xnor U20957 (N_20957,N_16841,N_16735);
nand U20958 (N_20958,N_19703,N_19679);
and U20959 (N_20959,N_15919,N_19997);
and U20960 (N_20960,N_16716,N_15229);
nor U20961 (N_20961,N_19897,N_18680);
nand U20962 (N_20962,N_16658,N_15331);
nand U20963 (N_20963,N_19496,N_16372);
nand U20964 (N_20964,N_16830,N_19661);
xor U20965 (N_20965,N_18293,N_18298);
xor U20966 (N_20966,N_18668,N_19507);
nand U20967 (N_20967,N_17398,N_16791);
or U20968 (N_20968,N_19548,N_18049);
xnor U20969 (N_20969,N_16978,N_15643);
or U20970 (N_20970,N_18083,N_15470);
or U20971 (N_20971,N_15794,N_16070);
nor U20972 (N_20972,N_15907,N_18689);
nand U20973 (N_20973,N_15241,N_19870);
and U20974 (N_20974,N_17866,N_19837);
and U20975 (N_20975,N_16637,N_17022);
and U20976 (N_20976,N_17540,N_18148);
nor U20977 (N_20977,N_16720,N_16243);
or U20978 (N_20978,N_17936,N_15873);
nor U20979 (N_20979,N_15780,N_19072);
xor U20980 (N_20980,N_16435,N_18921);
xnor U20981 (N_20981,N_15595,N_15513);
and U20982 (N_20982,N_15893,N_17410);
or U20983 (N_20983,N_19080,N_15849);
xnor U20984 (N_20984,N_19987,N_15036);
nand U20985 (N_20985,N_17285,N_17307);
and U20986 (N_20986,N_15715,N_17477);
nor U20987 (N_20987,N_16975,N_18082);
and U20988 (N_20988,N_19368,N_16468);
and U20989 (N_20989,N_17959,N_17383);
nand U20990 (N_20990,N_17730,N_19351);
nand U20991 (N_20991,N_19178,N_15725);
nor U20992 (N_20992,N_18570,N_16465);
or U20993 (N_20993,N_16814,N_18783);
and U20994 (N_20994,N_19365,N_18581);
and U20995 (N_20995,N_17500,N_17112);
and U20996 (N_20996,N_19206,N_17867);
or U20997 (N_20997,N_15748,N_18541);
and U20998 (N_20998,N_15891,N_16756);
and U20999 (N_20999,N_17397,N_15023);
and U21000 (N_21000,N_18439,N_16727);
xnor U21001 (N_21001,N_17327,N_18266);
nor U21002 (N_21002,N_15102,N_18133);
and U21003 (N_21003,N_17811,N_15510);
xnor U21004 (N_21004,N_15762,N_18755);
or U21005 (N_21005,N_19246,N_15620);
nand U21006 (N_21006,N_15495,N_18406);
and U21007 (N_21007,N_15749,N_16394);
xor U21008 (N_21008,N_15084,N_17803);
or U21009 (N_21009,N_18087,N_19084);
xor U21010 (N_21010,N_17482,N_16653);
nor U21011 (N_21011,N_18174,N_15313);
nor U21012 (N_21012,N_17690,N_16121);
nand U21013 (N_21013,N_17772,N_19236);
nor U21014 (N_21014,N_15496,N_16249);
nor U21015 (N_21015,N_16960,N_17717);
xor U21016 (N_21016,N_16533,N_19639);
nand U21017 (N_21017,N_17668,N_16096);
nor U21018 (N_21018,N_17187,N_15896);
nand U21019 (N_21019,N_19158,N_19866);
or U21020 (N_21020,N_16687,N_19664);
nor U21021 (N_21021,N_15399,N_19160);
nand U21022 (N_21022,N_18221,N_19378);
and U21023 (N_21023,N_19952,N_19823);
or U21024 (N_21024,N_16332,N_16586);
and U21025 (N_21025,N_17494,N_15450);
or U21026 (N_21026,N_19332,N_17704);
or U21027 (N_21027,N_16767,N_18269);
xor U21028 (N_21028,N_17856,N_18355);
xor U21029 (N_21029,N_15028,N_15099);
nor U21030 (N_21030,N_18635,N_18054);
or U21031 (N_21031,N_16748,N_16912);
nor U21032 (N_21032,N_18560,N_15714);
or U21033 (N_21033,N_15227,N_17566);
nand U21034 (N_21034,N_16545,N_18937);
or U21035 (N_21035,N_16130,N_17907);
xor U21036 (N_21036,N_15018,N_19481);
nand U21037 (N_21037,N_19722,N_19741);
or U21038 (N_21038,N_18691,N_19069);
or U21039 (N_21039,N_19502,N_16851);
xor U21040 (N_21040,N_18816,N_18096);
or U21041 (N_21041,N_17437,N_18983);
or U21042 (N_21042,N_18545,N_18743);
or U21043 (N_21043,N_17395,N_19499);
nor U21044 (N_21044,N_18585,N_17762);
xor U21045 (N_21045,N_19877,N_17964);
nor U21046 (N_21046,N_19390,N_18100);
and U21047 (N_21047,N_15913,N_19172);
xnor U21048 (N_21048,N_18841,N_15939);
xor U21049 (N_21049,N_18252,N_16003);
nor U21050 (N_21050,N_15220,N_17100);
or U21051 (N_21051,N_18566,N_16180);
xor U21052 (N_21052,N_19969,N_15000);
nand U21053 (N_21053,N_19685,N_16349);
nand U21054 (N_21054,N_16094,N_15466);
nand U21055 (N_21055,N_16783,N_19359);
xor U21056 (N_21056,N_19756,N_19491);
xor U21057 (N_21057,N_18207,N_19144);
xnor U21058 (N_21058,N_17120,N_19019);
nand U21059 (N_21059,N_18876,N_19299);
nand U21060 (N_21060,N_15949,N_18998);
nor U21061 (N_21061,N_19613,N_19622);
or U21062 (N_21062,N_19724,N_17206);
nand U21063 (N_21063,N_18586,N_18411);
or U21064 (N_21064,N_18617,N_18200);
and U21065 (N_21065,N_19424,N_17969);
xor U21066 (N_21066,N_18286,N_16883);
xor U21067 (N_21067,N_19260,N_18711);
xor U21068 (N_21068,N_15952,N_17710);
xor U21069 (N_21069,N_17261,N_19895);
nor U21070 (N_21070,N_16537,N_16429);
nand U21071 (N_21071,N_15539,N_17190);
and U21072 (N_21072,N_17041,N_18372);
or U21073 (N_21073,N_19240,N_17338);
xor U21074 (N_21074,N_15647,N_18628);
or U21075 (N_21075,N_16304,N_15179);
or U21076 (N_21076,N_16031,N_19259);
and U21077 (N_21077,N_15604,N_17523);
or U21078 (N_21078,N_16458,N_15502);
xor U21079 (N_21079,N_19925,N_15382);
and U21080 (N_21080,N_18595,N_19851);
xor U21081 (N_21081,N_17006,N_17834);
and U21082 (N_21082,N_15123,N_16699);
nor U21083 (N_21083,N_17335,N_16785);
xnor U21084 (N_21084,N_16177,N_19326);
or U21085 (N_21085,N_15587,N_18308);
and U21086 (N_21086,N_18347,N_15398);
nor U21087 (N_21087,N_18720,N_18811);
nand U21088 (N_21088,N_19609,N_18944);
and U21089 (N_21089,N_18330,N_19985);
nor U21090 (N_21090,N_17370,N_19271);
xnor U21091 (N_21091,N_16884,N_16275);
nand U21092 (N_21092,N_18413,N_19857);
nor U21093 (N_21093,N_15490,N_16808);
nand U21094 (N_21094,N_18918,N_16187);
nor U21095 (N_21095,N_18253,N_15827);
xnor U21096 (N_21096,N_19122,N_19972);
xnor U21097 (N_21097,N_18777,N_19587);
xor U21098 (N_21098,N_16577,N_19697);
nand U21099 (N_21099,N_15003,N_18130);
or U21100 (N_21100,N_19039,N_17808);
nand U21101 (N_21101,N_19010,N_19539);
or U21102 (N_21102,N_15881,N_16126);
nand U21103 (N_21103,N_15204,N_15160);
xor U21104 (N_21104,N_17439,N_17263);
and U21105 (N_21105,N_18645,N_19091);
nor U21106 (N_21106,N_17092,N_16225);
nor U21107 (N_21107,N_18195,N_15039);
nor U21108 (N_21108,N_15920,N_15081);
nor U21109 (N_21109,N_15879,N_17111);
and U21110 (N_21110,N_15428,N_18974);
or U21111 (N_21111,N_17103,N_15588);
xnor U21112 (N_21112,N_17431,N_18770);
or U21113 (N_21113,N_19185,N_17385);
and U21114 (N_21114,N_18956,N_17214);
nor U21115 (N_21115,N_15124,N_18022);
or U21116 (N_21116,N_18124,N_18164);
nor U21117 (N_21117,N_16199,N_15570);
nor U21118 (N_21118,N_15021,N_19374);
and U21119 (N_21119,N_18061,N_16900);
nand U21120 (N_21120,N_19137,N_16802);
nand U21121 (N_21121,N_15270,N_15829);
nor U21122 (N_21122,N_17065,N_15467);
nand U21123 (N_21123,N_18364,N_19793);
nand U21124 (N_21124,N_19801,N_17464);
nor U21125 (N_21125,N_15610,N_15904);
xnor U21126 (N_21126,N_16995,N_18036);
nand U21127 (N_21127,N_17584,N_16755);
or U21128 (N_21128,N_16305,N_16671);
nand U21129 (N_21129,N_18365,N_16188);
and U21130 (N_21130,N_17148,N_19032);
nor U21131 (N_21131,N_17888,N_15962);
nand U21132 (N_21132,N_17582,N_17971);
xnor U21133 (N_21133,N_19710,N_19297);
and U21134 (N_21134,N_17432,N_15987);
and U21135 (N_21135,N_16044,N_15844);
nor U21136 (N_21136,N_16073,N_15406);
nand U21137 (N_21137,N_19723,N_17525);
and U21138 (N_21138,N_18926,N_18199);
nand U21139 (N_21139,N_15909,N_18303);
nand U21140 (N_21140,N_18255,N_16064);
nand U21141 (N_21141,N_15045,N_15930);
xnor U21142 (N_21142,N_15322,N_19891);
nand U21143 (N_21143,N_16635,N_18718);
and U21144 (N_21144,N_16065,N_19208);
and U21145 (N_21145,N_15544,N_15494);
nor U21146 (N_21146,N_19296,N_19791);
xnor U21147 (N_21147,N_17207,N_15566);
or U21148 (N_21148,N_18379,N_15775);
and U21149 (N_21149,N_16607,N_18420);
nand U21150 (N_21150,N_16789,N_19162);
xor U21151 (N_21151,N_17233,N_18970);
nand U21152 (N_21152,N_19715,N_18151);
xor U21153 (N_21153,N_18134,N_18105);
nor U21154 (N_21154,N_19261,N_18162);
or U21155 (N_21155,N_17997,N_16268);
or U21156 (N_21156,N_17904,N_17170);
xor U21157 (N_21157,N_19904,N_16543);
nor U21158 (N_21158,N_18321,N_19016);
or U21159 (N_21159,N_19771,N_16213);
or U21160 (N_21160,N_18593,N_15352);
or U21161 (N_21161,N_15300,N_18053);
nand U21162 (N_21162,N_19642,N_19769);
or U21163 (N_21163,N_15049,N_18532);
xor U21164 (N_21164,N_15895,N_18088);
xnor U21165 (N_21165,N_15368,N_16934);
xor U21166 (N_21166,N_19194,N_15218);
or U21167 (N_21167,N_17511,N_16909);
and U21168 (N_21168,N_18251,N_17896);
nor U21169 (N_21169,N_15623,N_16918);
xor U21170 (N_21170,N_19147,N_17179);
nor U21171 (N_21171,N_17946,N_19523);
nand U21172 (N_21172,N_19804,N_16083);
or U21173 (N_21173,N_17979,N_16297);
xnor U21174 (N_21174,N_16696,N_19456);
nand U21175 (N_21175,N_15280,N_19853);
nor U21176 (N_21176,N_18573,N_19946);
xnor U21177 (N_21177,N_18243,N_18602);
nand U21178 (N_21178,N_19796,N_15046);
nand U21179 (N_21179,N_15810,N_18992);
or U21180 (N_21180,N_15694,N_19619);
xor U21181 (N_21181,N_16933,N_18959);
nand U21182 (N_21182,N_15001,N_19377);
and U21183 (N_21183,N_19514,N_19916);
xnor U21184 (N_21184,N_16704,N_18872);
and U21185 (N_21185,N_15716,N_19111);
or U21186 (N_21186,N_17608,N_15709);
nand U21187 (N_21187,N_19110,N_17758);
or U21188 (N_21188,N_16127,N_17723);
or U21189 (N_21189,N_18402,N_18895);
and U21190 (N_21190,N_17718,N_16685);
nand U21191 (N_21191,N_15128,N_15958);
xnor U21192 (N_21192,N_16387,N_16648);
nor U21193 (N_21193,N_19674,N_16665);
nor U21194 (N_21194,N_17952,N_19213);
and U21195 (N_21195,N_17014,N_15464);
and U21196 (N_21196,N_17005,N_15640);
and U21197 (N_21197,N_17985,N_18786);
xor U21198 (N_21198,N_17308,N_19468);
or U21199 (N_21199,N_18086,N_15978);
nor U21200 (N_21200,N_15649,N_19833);
nand U21201 (N_21201,N_19930,N_18259);
nor U21202 (N_21202,N_15311,N_17497);
nand U21203 (N_21203,N_16476,N_17852);
xor U21204 (N_21204,N_15627,N_16559);
nand U21205 (N_21205,N_18118,N_18119);
xor U21206 (N_21206,N_17627,N_17375);
xnor U21207 (N_21207,N_17715,N_19705);
nand U21208 (N_21208,N_19417,N_15083);
nor U21209 (N_21209,N_19524,N_19889);
nand U21210 (N_21210,N_16959,N_18733);
xnor U21211 (N_21211,N_16084,N_16826);
nand U21212 (N_21212,N_15389,N_16204);
nand U21213 (N_21213,N_19477,N_17257);
and U21214 (N_21214,N_15954,N_18646);
nor U21215 (N_21215,N_15861,N_19315);
and U21216 (N_21216,N_18033,N_18408);
xnor U21217 (N_21217,N_15294,N_15543);
and U21218 (N_21218,N_16285,N_18031);
nand U21219 (N_21219,N_18748,N_17173);
nand U21220 (N_21220,N_19732,N_17513);
nand U21221 (N_21221,N_18240,N_16101);
or U21222 (N_21222,N_18169,N_18535);
nor U21223 (N_21223,N_19513,N_16359);
nand U21224 (N_21224,N_18287,N_16261);
and U21225 (N_21225,N_16546,N_16623);
nor U21226 (N_21226,N_16775,N_19498);
and U21227 (N_21227,N_15989,N_17791);
xnor U21228 (N_21228,N_16743,N_19790);
or U21229 (N_21229,N_19577,N_16838);
nand U21230 (N_21230,N_17676,N_16575);
nand U21231 (N_21231,N_18746,N_16450);
or U21232 (N_21232,N_18450,N_17175);
or U21233 (N_21233,N_15540,N_16206);
nor U21234 (N_21234,N_16076,N_17842);
nand U21235 (N_21235,N_19383,N_17716);
nand U21236 (N_21236,N_18163,N_18470);
nand U21237 (N_21237,N_15508,N_17119);
or U21238 (N_21238,N_17292,N_19291);
nor U21239 (N_21239,N_18958,N_17775);
xnor U21240 (N_21240,N_15097,N_18568);
xnor U21241 (N_21241,N_18822,N_18121);
or U21242 (N_21242,N_16600,N_18724);
or U21243 (N_21243,N_18047,N_19829);
and U21244 (N_21244,N_17714,N_19470);
and U21245 (N_21245,N_16330,N_16513);
and U21246 (N_21246,N_15771,N_17688);
nand U21247 (N_21247,N_15734,N_18804);
and U21248 (N_21248,N_19680,N_17425);
nand U21249 (N_21249,N_17881,N_17821);
nor U21250 (N_21250,N_16548,N_17422);
or U21251 (N_21251,N_17132,N_18715);
xnor U21252 (N_21252,N_18731,N_16619);
xor U21253 (N_21253,N_15984,N_19665);
nor U21254 (N_21254,N_16147,N_18583);
and U21255 (N_21255,N_17973,N_18940);
and U21256 (N_21256,N_15787,N_16376);
and U21257 (N_21257,N_15602,N_17894);
or U21258 (N_21258,N_19055,N_16757);
nor U21259 (N_21259,N_16288,N_15717);
xnor U21260 (N_21260,N_19983,N_18859);
xor U21261 (N_21261,N_17713,N_19811);
and U21262 (N_21262,N_19566,N_17153);
nor U21263 (N_21263,N_17721,N_19049);
and U21264 (N_21264,N_16176,N_19220);
xor U21265 (N_21265,N_16113,N_18608);
nand U21266 (N_21266,N_15162,N_16850);
or U21267 (N_21267,N_15321,N_16062);
and U21268 (N_21268,N_17628,N_15703);
and U21269 (N_21269,N_15972,N_18156);
or U21270 (N_21270,N_16606,N_15820);
xor U21271 (N_21271,N_15674,N_15591);
and U21272 (N_21272,N_18709,N_16411);
or U21273 (N_21273,N_15391,N_19511);
and U21274 (N_21274,N_17711,N_19495);
nand U21275 (N_21275,N_18244,N_17248);
and U21276 (N_21276,N_18495,N_19423);
xor U21277 (N_21277,N_16254,N_15700);
nor U21278 (N_21278,N_15299,N_15452);
or U21279 (N_21279,N_19978,N_17817);
nor U21280 (N_21280,N_15262,N_17727);
or U21281 (N_21281,N_18831,N_16539);
nor U21282 (N_21282,N_15865,N_17122);
nand U21283 (N_21283,N_19525,N_15572);
and U21284 (N_21284,N_17962,N_17361);
xnor U21285 (N_21285,N_17613,N_17991);
xor U21286 (N_21286,N_18813,N_19620);
and U21287 (N_21287,N_16368,N_18261);
nand U21288 (N_21288,N_19322,N_16321);
or U21289 (N_21289,N_18388,N_19092);
xnor U21290 (N_21290,N_19940,N_19994);
nor U21291 (N_21291,N_19504,N_19054);
nand U21292 (N_21292,N_17035,N_17884);
and U21293 (N_21293,N_18123,N_15872);
xnor U21294 (N_21294,N_19917,N_15175);
xor U21295 (N_21295,N_17901,N_18845);
or U21296 (N_21296,N_16805,N_15233);
xor U21297 (N_21297,N_19186,N_18401);
xnor U21298 (N_21298,N_15690,N_19583);
nor U21299 (N_21299,N_18480,N_19546);
or U21300 (N_21300,N_18020,N_19576);
or U21301 (N_21301,N_17208,N_15738);
and U21302 (N_21302,N_18215,N_16389);
nor U21303 (N_21303,N_15473,N_19044);
and U21304 (N_21304,N_15580,N_16150);
nor U21305 (N_21305,N_19831,N_17617);
nand U21306 (N_21306,N_19275,N_19575);
and U21307 (N_21307,N_15110,N_15522);
and U21308 (N_21308,N_19349,N_15626);
xor U21309 (N_21309,N_15344,N_15825);
or U21310 (N_21310,N_15583,N_18257);
nand U21311 (N_21311,N_17250,N_16556);
nor U21312 (N_21312,N_17201,N_17855);
nor U21313 (N_21313,N_16074,N_17725);
xnor U21314 (N_21314,N_16133,N_16051);
nor U21315 (N_21315,N_19690,N_19302);
and U21316 (N_21316,N_18384,N_18090);
xnor U21317 (N_21317,N_18141,N_16881);
nand U21318 (N_21318,N_16874,N_15137);
nor U21319 (N_21319,N_16521,N_17616);
nor U21320 (N_21320,N_19645,N_19776);
nor U21321 (N_21321,N_16260,N_16278);
and U21322 (N_21322,N_18962,N_16592);
and U21323 (N_21323,N_17009,N_19719);
nor U21324 (N_21324,N_18202,N_17871);
nor U21325 (N_21325,N_16787,N_17021);
nor U21326 (N_21326,N_18906,N_17230);
xor U21327 (N_21327,N_19763,N_17857);
or U21328 (N_21328,N_19407,N_16043);
and U21329 (N_21329,N_16222,N_17359);
or U21330 (N_21330,N_15434,N_19510);
and U21331 (N_21331,N_15455,N_15349);
nor U21332 (N_21332,N_18844,N_17524);
xor U21333 (N_21333,N_19118,N_18191);
nand U21334 (N_21334,N_17913,N_17191);
and U21335 (N_21335,N_15150,N_16379);
nand U21336 (N_21336,N_15027,N_17341);
nand U21337 (N_21337,N_19253,N_19616);
nor U21338 (N_21338,N_19042,N_17184);
and U21339 (N_21339,N_18363,N_18476);
xor U21340 (N_21340,N_15465,N_17529);
or U21341 (N_21341,N_15878,N_16639);
or U21342 (N_21342,N_17828,N_17004);
nand U21343 (N_21343,N_16469,N_17326);
nor U21344 (N_21344,N_16820,N_17393);
xor U21345 (N_21345,N_16316,N_19505);
xor U21346 (N_21346,N_16873,N_16655);
nand U21347 (N_21347,N_15377,N_16267);
xnor U21348 (N_21348,N_17943,N_17420);
nor U21349 (N_21349,N_17196,N_15783);
and U21350 (N_21350,N_15105,N_18018);
or U21351 (N_21351,N_19290,N_17783);
or U21352 (N_21352,N_19663,N_15790);
or U21353 (N_21353,N_16766,N_17829);
nor U21354 (N_21354,N_16730,N_18168);
nor U21355 (N_21355,N_18512,N_15843);
and U21356 (N_21356,N_15894,N_19345);
or U21357 (N_21357,N_16058,N_19115);
or U21358 (N_21358,N_19043,N_16869);
xor U21359 (N_21359,N_17418,N_16812);
nand U21360 (N_21360,N_16351,N_17545);
or U21361 (N_21361,N_17776,N_17212);
or U21362 (N_21362,N_17492,N_15739);
or U21363 (N_21363,N_17508,N_18081);
or U21364 (N_21364,N_18499,N_15877);
nand U21365 (N_21365,N_18787,N_19696);
and U21366 (N_21366,N_18629,N_19153);
nor U21367 (N_21367,N_19984,N_17239);
nand U21368 (N_21368,N_17534,N_15267);
xor U21369 (N_21369,N_18964,N_16570);
xor U21370 (N_21370,N_16937,N_19745);
nand U21371 (N_21371,N_19758,N_18317);
nand U21372 (N_21372,N_18444,N_19041);
xnor U21373 (N_21373,N_17389,N_15677);
and U21374 (N_21374,N_17568,N_16765);
or U21375 (N_21375,N_15917,N_19515);
and U21376 (N_21376,N_16466,N_17786);
nor U21377 (N_21377,N_18407,N_15777);
nor U21378 (N_21378,N_18567,N_17995);
nand U21379 (N_21379,N_15518,N_16719);
and U21380 (N_21380,N_19440,N_18987);
xnor U21381 (N_21381,N_18146,N_17498);
nor U21382 (N_21382,N_15648,N_16848);
nand U21383 (N_21383,N_19347,N_17845);
nor U21384 (N_21384,N_15447,N_19323);
nor U21385 (N_21385,N_16728,N_15269);
nor U21386 (N_21386,N_19256,N_16734);
xnor U21387 (N_21387,N_18219,N_15970);
or U21388 (N_21388,N_17280,N_19802);
nand U21389 (N_21389,N_17700,N_16383);
and U21390 (N_21390,N_19395,N_17118);
and U21391 (N_21391,N_15459,N_19161);
xor U21392 (N_21392,N_19600,N_15660);
and U21393 (N_21393,N_17876,N_16221);
and U21394 (N_21394,N_18670,N_19048);
nor U21395 (N_21395,N_15993,N_17747);
nor U21396 (N_21396,N_17407,N_16452);
nand U21397 (N_21397,N_19806,N_17350);
nand U21398 (N_21398,N_15607,N_15432);
xor U21399 (N_21399,N_16683,N_17759);
xor U21400 (N_21400,N_15839,N_19563);
and U21401 (N_21401,N_16565,N_17919);
nand U21402 (N_21402,N_17002,N_17209);
nand U21403 (N_21403,N_19105,N_19149);
and U21404 (N_21404,N_15437,N_16344);
or U21405 (N_21405,N_17551,N_18005);
nand U21406 (N_21406,N_15121,N_16148);
or U21407 (N_21407,N_15435,N_19497);
nand U21408 (N_21408,N_15653,N_15334);
and U21409 (N_21409,N_18843,N_19956);
or U21410 (N_21410,N_15923,N_17135);
and U21411 (N_21411,N_19306,N_16793);
xnor U21412 (N_21412,N_17794,N_18075);
nand U21413 (N_21413,N_19725,N_19361);
and U21414 (N_21414,N_18166,N_15042);
nand U21415 (N_21415,N_19375,N_15779);
nor U21416 (N_21416,N_15356,N_16647);
xor U21417 (N_21417,N_16356,N_19446);
xnor U21418 (N_21418,N_19928,N_17468);
xnor U21419 (N_21419,N_16489,N_16292);
and U21420 (N_21420,N_18446,N_17343);
and U21421 (N_21421,N_17928,N_15271);
nor U21422 (N_21422,N_16516,N_17224);
or U21423 (N_21423,N_16906,N_17663);
xnor U21424 (N_21424,N_19338,N_18898);
and U21425 (N_21425,N_17436,N_18462);
or U21426 (N_21426,N_16833,N_16114);
xor U21427 (N_21427,N_15244,N_17435);
xor U21428 (N_21428,N_19294,N_15914);
nand U21429 (N_21429,N_16777,N_16373);
nand U21430 (N_21430,N_15797,N_19085);
and U21431 (N_21431,N_19950,N_17681);
nor U21432 (N_21432,N_18606,N_17798);
or U21433 (N_21433,N_18468,N_16844);
and U21434 (N_21434,N_18238,N_18414);
and U21435 (N_21435,N_16061,N_19116);
nor U21436 (N_21436,N_19473,N_19068);
or U21437 (N_21437,N_19568,N_18157);
xor U21438 (N_21438,N_18857,N_19094);
and U21439 (N_21439,N_15329,N_19803);
or U21440 (N_21440,N_15420,N_18296);
or U21441 (N_21441,N_15314,N_19357);
nand U21442 (N_21442,N_18710,N_19005);
or U21443 (N_21443,N_17516,N_18356);
and U21444 (N_21444,N_18080,N_18122);
or U21445 (N_21445,N_19366,N_17055);
and U21446 (N_21446,N_18536,N_18092);
or U21447 (N_21447,N_16832,N_16038);
nor U21448 (N_21448,N_15359,N_18447);
nor U21449 (N_21449,N_17987,N_19695);
and U21450 (N_21450,N_17908,N_17642);
and U21451 (N_21451,N_19175,N_19562);
nand U21452 (N_21452,N_16553,N_16705);
and U21453 (N_21453,N_15631,N_19188);
nand U21454 (N_21454,N_15133,N_15622);
or U21455 (N_21455,N_16227,N_15012);
nand U21456 (N_21456,N_16000,N_15264);
nor U21457 (N_21457,N_16131,N_16186);
nand U21458 (N_21458,N_18735,N_17607);
xor U21459 (N_21459,N_19649,N_15890);
xnor U21460 (N_21460,N_17080,N_18160);
or U21461 (N_21461,N_18220,N_17875);
nor U21462 (N_21462,N_15281,N_17347);
or U21463 (N_21463,N_16510,N_17891);
or U21464 (N_21464,N_18578,N_19996);
nor U21465 (N_21465,N_19076,N_17318);
xnor U21466 (N_21466,N_19964,N_17707);
nand U21467 (N_21467,N_16633,N_19264);
nand U21468 (N_21468,N_18127,N_17247);
xor U21469 (N_21469,N_19273,N_17345);
xor U21470 (N_21470,N_15228,N_15761);
nand U21471 (N_21471,N_19274,N_16944);
and U21472 (N_21472,N_16461,N_17597);
and U21473 (N_21473,N_15711,N_18270);
or U21474 (N_21474,N_15520,N_17770);
and U21475 (N_21475,N_17146,N_18458);
and U21476 (N_21476,N_17117,N_17537);
nor U21477 (N_21477,N_19651,N_16338);
xor U21478 (N_21478,N_15858,N_15741);
and U21479 (N_21479,N_17211,N_17954);
xor U21480 (N_21480,N_15393,N_18867);
and U21481 (N_21481,N_15198,N_16843);
or U21482 (N_21482,N_18205,N_19673);
nand U21483 (N_21483,N_18861,N_15113);
nand U21484 (N_21484,N_15031,N_16769);
and U21485 (N_21485,N_19248,N_17023);
or U21486 (N_21486,N_16951,N_16939);
nand U21487 (N_21487,N_18825,N_16617);
and U21488 (N_21488,N_15638,N_18249);
nand U21489 (N_21489,N_15726,N_19030);
or U21490 (N_21490,N_19189,N_15015);
nand U21491 (N_21491,N_15167,N_16154);
xnor U21492 (N_21492,N_15617,N_16697);
nor U21493 (N_21493,N_18761,N_19760);
xnor U21494 (N_21494,N_17322,N_19943);
nand U21495 (N_21495,N_19346,N_19825);
and U21496 (N_21496,N_17015,N_19579);
and U21497 (N_21497,N_17454,N_17394);
or U21498 (N_21498,N_18052,N_15256);
nand U21499 (N_21499,N_15419,N_18638);
and U21500 (N_21500,N_15531,N_16726);
and U21501 (N_21501,N_17367,N_18183);
nor U21502 (N_21502,N_16759,N_15011);
and U21503 (N_21503,N_18793,N_15740);
or U21504 (N_21504,N_16632,N_15609);
nor U21505 (N_21505,N_18178,N_19708);
and U21506 (N_21506,N_15230,N_19592);
nor U21507 (N_21507,N_16005,N_18418);
and U21508 (N_21508,N_19834,N_16738);
and U21509 (N_21509,N_16603,N_18878);
nor U21510 (N_21510,N_17428,N_16813);
nand U21511 (N_21511,N_18678,N_19165);
nand U21512 (N_21512,N_15804,N_15054);
or U21513 (N_21513,N_15041,N_17456);
nand U21514 (N_21514,N_19832,N_19691);
or U21515 (N_21515,N_15385,N_15504);
and U21516 (N_21516,N_18496,N_17017);
xor U21517 (N_21517,N_18348,N_19666);
nand U21518 (N_21518,N_19469,N_17812);
nor U21519 (N_21519,N_15636,N_19792);
xnor U21520 (N_21520,N_15390,N_16190);
and U21521 (N_21521,N_19196,N_16892);
nor U21522 (N_21522,N_16164,N_19764);
nand U21523 (N_21523,N_16494,N_16233);
xor U21524 (N_21524,N_19812,N_17552);
and U21525 (N_21525,N_16871,N_15403);
and U21526 (N_21526,N_15476,N_18824);
and U21527 (N_21527,N_17669,N_18492);
nand U21528 (N_21528,N_19728,N_19464);
or U21529 (N_21529,N_19408,N_15698);
or U21530 (N_21530,N_18466,N_16531);
and U21531 (N_21531,N_15275,N_19245);
nor U21532 (N_21532,N_16490,N_19894);
nor U21533 (N_21533,N_18732,N_17988);
nor U21534 (N_21534,N_19281,N_16625);
nor U21535 (N_21535,N_17357,N_19531);
xor U21536 (N_21536,N_19822,N_18812);
and U21537 (N_21537,N_17266,N_15852);
xor U21538 (N_21538,N_16362,N_17149);
xor U21539 (N_21539,N_19179,N_17000);
nand U21540 (N_21540,N_17874,N_15408);
nor U21541 (N_21541,N_17993,N_18826);
nand U21542 (N_21542,N_15763,N_19011);
nor U21543 (N_21543,N_19443,N_16668);
xnor U21544 (N_21544,N_15245,N_16499);
nand U21545 (N_21545,N_16929,N_15944);
nor U21546 (N_21546,N_15224,N_15658);
or U21547 (N_21547,N_16231,N_19355);
nor U21548 (N_21548,N_15415,N_17787);
and U21549 (N_21549,N_19571,N_17737);
nand U21550 (N_21550,N_16956,N_17743);
nor U21551 (N_21551,N_15926,N_15469);
and U21552 (N_21552,N_17831,N_19683);
xnor U21553 (N_21553,N_17151,N_16829);
and U21554 (N_21554,N_16355,N_19367);
xor U21555 (N_21555,N_19807,N_18010);
nand U21556 (N_21556,N_16877,N_16614);
or U21557 (N_21557,N_17156,N_16308);
or U21558 (N_21558,N_16366,N_18350);
nor U21559 (N_21559,N_19327,N_17802);
or U21560 (N_21560,N_16503,N_15683);
xnor U21561 (N_21561,N_17557,N_18315);
and U21562 (N_21562,N_18888,N_18386);
or U21563 (N_21563,N_15596,N_16017);
xor U21564 (N_21564,N_19582,N_15260);
nand U21565 (N_21565,N_15069,N_17279);
nand U21566 (N_21566,N_19396,N_17813);
nor U21567 (N_21567,N_17705,N_19938);
and U21568 (N_21568,N_16684,N_16103);
or U21569 (N_21569,N_19580,N_17003);
nor U21570 (N_21570,N_19075,N_18509);
nand U21571 (N_21571,N_17038,N_19824);
nor U21572 (N_21572,N_16067,N_17281);
or U21573 (N_21573,N_15534,N_18834);
xnor U21574 (N_21574,N_16698,N_15255);
or U21575 (N_21575,N_17662,N_19941);
nand U21576 (N_21576,N_16259,N_16007);
nor U21577 (N_21577,N_17510,N_17892);
and U21578 (N_21578,N_18396,N_15073);
and U21579 (N_21579,N_16132,N_19211);
nand U21580 (N_21580,N_18671,N_17848);
nand U21581 (N_21581,N_16890,N_16529);
nor U21582 (N_21582,N_15784,N_17544);
xnor U21583 (N_21583,N_16393,N_16612);
xnor U21584 (N_21584,N_17090,N_19962);
nand U21585 (N_21585,N_18854,N_18833);
nand U21586 (N_21586,N_16426,N_18988);
and U21587 (N_21587,N_17219,N_16208);
or U21588 (N_21588,N_15279,N_18744);
or U21589 (N_21589,N_15347,N_15315);
or U21590 (N_21590,N_17744,N_18782);
xor U21591 (N_21591,N_15400,N_15426);
nand U21592 (N_21592,N_15489,N_18101);
xor U21593 (N_21593,N_16205,N_17165);
or U21594 (N_21594,N_18719,N_16258);
nor U21595 (N_21595,N_15112,N_16272);
nor U21596 (N_21596,N_18077,N_19744);
and U21597 (N_21597,N_17605,N_16761);
or U21598 (N_21598,N_15376,N_18224);
nand U21599 (N_21599,N_16495,N_19308);
nor U21600 (N_21600,N_19125,N_15090);
xnor U21601 (N_21601,N_18064,N_15370);
nand U21602 (N_21602,N_15995,N_16317);
xnor U21603 (N_21603,N_16977,N_15357);
or U21604 (N_21604,N_15085,N_18997);
nor U21605 (N_21605,N_18605,N_18969);
nor U21606 (N_21606,N_15288,N_18907);
or U21607 (N_21607,N_19065,N_16388);
nor U21608 (N_21608,N_19324,N_19675);
and U21609 (N_21609,N_19373,N_18798);
nor U21610 (N_21610,N_19686,N_18059);
and U21611 (N_21611,N_15369,N_15193);
or U21612 (N_21612,N_16082,N_18950);
or U21613 (N_21613,N_16746,N_19871);
xor U21614 (N_21614,N_16597,N_16014);
nand U21615 (N_21615,N_17934,N_19988);
or U21616 (N_21616,N_16360,N_19875);
or U21617 (N_21617,N_15528,N_19684);
and U21618 (N_21618,N_15892,N_16689);
or U21619 (N_21619,N_15815,N_18491);
nand U21620 (N_21620,N_17944,N_16478);
and U21621 (N_21621,N_16974,N_18765);
or U21622 (N_21622,N_19593,N_15429);
and U21623 (N_21623,N_19435,N_16941);
and U21624 (N_21624,N_15553,N_18095);
or U21625 (N_21625,N_15801,N_15174);
or U21626 (N_21626,N_17476,N_19331);
nand U21627 (N_21627,N_15736,N_19104);
and U21628 (N_21628,N_18784,N_17274);
or U21629 (N_21629,N_18028,N_19046);
nand U21630 (N_21630,N_18340,N_18521);
and U21631 (N_21631,N_19914,N_18389);
xor U21632 (N_21632,N_18839,N_18482);
and U21633 (N_21633,N_15108,N_19457);
or U21634 (N_21634,N_16331,N_19057);
xnor U21635 (N_21635,N_17365,N_17789);
or U21636 (N_21636,N_18823,N_18359);
nand U21637 (N_21637,N_15793,N_19460);
xnor U21638 (N_21638,N_18210,N_16857);
nand U21639 (N_21639,N_15080,N_16807);
nand U21640 (N_21640,N_16642,N_19694);
and U21641 (N_21641,N_17563,N_16385);
xor U21642 (N_21642,N_17369,N_18757);
xnor U21643 (N_21643,N_19081,N_17553);
and U21644 (N_21644,N_16827,N_17131);
or U21645 (N_21645,N_19526,N_15963);
nand U21646 (N_21646,N_18186,N_17457);
or U21647 (N_21647,N_18041,N_16271);
nand U21648 (N_21648,N_19014,N_19735);
xor U21649 (N_21649,N_17974,N_19841);
nand U21650 (N_21650,N_15367,N_17752);
xor U21651 (N_21651,N_19459,N_17299);
or U21652 (N_21652,N_19778,N_17506);
xnor U21653 (N_21653,N_17127,N_17043);
nor U21654 (N_21654,N_16666,N_16664);
nand U21655 (N_21655,N_19658,N_19090);
or U21656 (N_21656,N_15722,N_19123);
nand U21657 (N_21657,N_15830,N_15661);
or U21658 (N_21658,N_19612,N_19839);
and U21659 (N_21659,N_18819,N_15899);
xnor U21660 (N_21660,N_17011,N_15816);
nor U21661 (N_21661,N_15165,N_16547);
and U21662 (N_21662,N_18828,N_16191);
nand U21663 (N_21663,N_15514,N_15075);
nor U21664 (N_21664,N_19420,N_16115);
nand U21665 (N_21665,N_19488,N_15472);
nand U21666 (N_21666,N_18387,N_17251);
and U21667 (N_21667,N_15436,N_15961);
and U21668 (N_21668,N_18432,N_16809);
nor U21669 (N_21669,N_15107,N_19508);
xnor U21670 (N_21670,N_15444,N_17178);
nand U21671 (N_21671,N_15991,N_17490);
nor U21672 (N_21672,N_19121,N_17040);
xnor U21673 (N_21673,N_19058,N_16060);
nor U21674 (N_21674,N_19157,N_17869);
nor U21675 (N_21675,N_19405,N_16211);
and U21676 (N_21676,N_18982,N_17391);
and U21677 (N_21677,N_15760,N_19089);
xnor U21678 (N_21678,N_19688,N_15296);
xnor U21679 (N_21679,N_19992,N_16160);
xnor U21680 (N_21680,N_16095,N_15955);
or U21681 (N_21681,N_15669,N_16650);
nand U21682 (N_21682,N_18006,N_17229);
or U21683 (N_21683,N_19082,N_19596);
xor U21684 (N_21684,N_16863,N_16896);
nand U21685 (N_21685,N_18799,N_15342);
or U21686 (N_21686,N_17387,N_19633);
nor U21687 (N_21687,N_16263,N_19805);
and U21688 (N_21688,N_19874,N_17647);
and U21689 (N_21689,N_18683,N_18611);
nand U21690 (N_21690,N_18063,N_19749);
xnor U21691 (N_21691,N_19720,N_16486);
nand U21692 (N_21692,N_19143,N_16859);
xnor U21693 (N_21693,N_18805,N_15034);
nor U21694 (N_21694,N_19647,N_16137);
nor U21695 (N_21695,N_19961,N_19536);
or U21696 (N_21696,N_17194,N_18540);
nor U21697 (N_21697,N_15449,N_16522);
xor U21698 (N_21698,N_16627,N_18936);
nand U21699 (N_21699,N_17399,N_18176);
nor U21700 (N_21700,N_18474,N_15223);
or U21701 (N_21701,N_15634,N_16146);
nor U21702 (N_21702,N_15809,N_15988);
and U21703 (N_21703,N_15903,N_15868);
xnor U21704 (N_21704,N_16610,N_17143);
nor U21705 (N_21705,N_16120,N_18285);
or U21706 (N_21706,N_16645,N_17633);
and U21707 (N_21707,N_17330,N_19127);
and U21708 (N_21708,N_17430,N_16945);
xor U21709 (N_21709,N_19409,N_15180);
nor U21710 (N_21710,N_17905,N_18519);
or U21711 (N_21711,N_16135,N_15185);
xnor U21712 (N_21712,N_15052,N_15394);
xor U21713 (N_21713,N_19626,N_15831);
nor U21714 (N_21714,N_17265,N_19931);
xor U21715 (N_21715,N_17697,N_16817);
nand U21716 (N_21716,N_15619,N_17088);
nor U21717 (N_21717,N_17396,N_19107);
nor U21718 (N_21718,N_16904,N_15067);
nand U21719 (N_21719,N_17337,N_18942);
nand U21720 (N_21720,N_17515,N_18930);
nor U21721 (N_21721,N_15154,N_16550);
xor U21722 (N_21722,N_19543,N_16708);
xor U21723 (N_21723,N_15053,N_17965);
or U21724 (N_21724,N_17427,N_18712);
nor U21725 (N_21725,N_16776,N_18155);
nor U21726 (N_21726,N_18758,N_15515);
or U21727 (N_21727,N_16703,N_19712);
xor U21728 (N_21728,N_16889,N_18737);
xor U21729 (N_21729,N_18766,N_18150);
nand U21730 (N_21730,N_17986,N_19201);
nor U21731 (N_21731,N_18112,N_16433);
or U21732 (N_21732,N_18725,N_18511);
nand U21733 (N_21733,N_17222,N_18508);
or U21734 (N_21734,N_18159,N_15247);
or U21735 (N_21735,N_16891,N_17528);
xor U21736 (N_21736,N_17027,N_17108);
nand U21737 (N_21737,N_16237,N_18693);
nor U21738 (N_21738,N_19738,N_16616);
or U21739 (N_21739,N_15645,N_17637);
nor U21740 (N_21740,N_18201,N_19862);
nor U21741 (N_21741,N_19286,N_19413);
or U21742 (N_21742,N_18376,N_15320);
xor U21743 (N_21743,N_15911,N_15274);
and U21744 (N_21744,N_16567,N_16182);
and U21745 (N_21745,N_15983,N_15111);
nand U21746 (N_21746,N_16742,N_16283);
nand U21747 (N_21747,N_18185,N_18275);
nor U21748 (N_21748,N_15261,N_17133);
nand U21749 (N_21749,N_19061,N_18803);
or U21750 (N_21750,N_17295,N_15325);
xnor U21751 (N_21751,N_19450,N_15131);
xnor U21752 (N_21752,N_15851,N_17581);
nor U21753 (N_21753,N_15521,N_15730);
nand U21754 (N_21754,N_15336,N_18965);
xor U21755 (N_21755,N_18914,N_17491);
nor U21756 (N_21756,N_16168,N_19414);
and U21757 (N_21757,N_17372,N_17592);
or U21758 (N_21758,N_19313,N_16502);
xnor U21759 (N_21759,N_17152,N_15537);
nand U21760 (N_21760,N_19017,N_17013);
nor U21761 (N_21761,N_17740,N_17453);
and U21762 (N_21762,N_15941,N_19794);
or U21763 (N_21763,N_16492,N_17074);
and U21764 (N_21764,N_17203,N_19050);
nor U21765 (N_21765,N_19285,N_18659);
nor U21766 (N_21766,N_16702,N_17288);
nor U21767 (N_21767,N_16444,N_17532);
and U21768 (N_21768,N_19990,N_19437);
nor U21769 (N_21769,N_15599,N_19447);
nand U21770 (N_21770,N_16680,N_15751);
nor U21771 (N_21771,N_15618,N_17479);
nand U21772 (N_21772,N_19544,N_17291);
nor U21773 (N_21773,N_16193,N_15056);
nor U21774 (N_21774,N_16251,N_16950);
or U21775 (N_21775,N_18039,N_18333);
and U21776 (N_21776,N_17449,N_19595);
or U21777 (N_21777,N_17488,N_19177);
and U21778 (N_21778,N_19560,N_19102);
or U21779 (N_21779,N_18309,N_17522);
or U21780 (N_21780,N_19951,N_17110);
or U21781 (N_21781,N_16274,N_15556);
nor U21782 (N_21782,N_16371,N_17434);
xor U21783 (N_21783,N_16423,N_16440);
nor U21784 (N_21784,N_16578,N_19784);
or U21785 (N_21785,N_19071,N_17413);
and U21786 (N_21786,N_17262,N_18438);
nand U21787 (N_21787,N_16574,N_15691);
nor U21788 (N_21788,N_17321,N_17660);
xor U21789 (N_21789,N_16107,N_15506);
xor U21790 (N_21790,N_19287,N_15688);
nand U21791 (N_21791,N_17981,N_19003);
nand U21792 (N_21792,N_15875,N_18074);
or U21793 (N_21793,N_17415,N_18099);
nor U21794 (N_21794,N_17625,N_19727);
xnor U21795 (N_21795,N_16280,N_15689);
and U21796 (N_21796,N_18173,N_19606);
or U21797 (N_21797,N_16223,N_17963);
or U21798 (N_21798,N_17550,N_19317);
and U21799 (N_21799,N_17243,N_16341);
nand U21800 (N_21800,N_18120,N_17868);
and U21801 (N_21801,N_19114,N_18292);
nand U21802 (N_21802,N_17531,N_17680);
xor U21803 (N_21803,N_19203,N_17056);
or U21804 (N_21804,N_19569,N_17873);
or U21805 (N_21805,N_18905,N_16298);
and U21806 (N_21806,N_17481,N_17163);
or U21807 (N_21807,N_17837,N_16347);
nor U21808 (N_21808,N_18009,N_17631);
or U21809 (N_21809,N_16313,N_15953);
nand U21810 (N_21810,N_16518,N_19483);
nand U21811 (N_21811,N_18654,N_19888);
xor U21812 (N_21812,N_16498,N_18206);
and U21813 (N_21813,N_15438,N_16470);
nand U21814 (N_21814,N_17256,N_19073);
or U21815 (N_21815,N_18091,N_19689);
nand U21816 (N_21816,N_18624,N_16967);
xor U21817 (N_21817,N_17646,N_19999);
and U21818 (N_21818,N_18301,N_17227);
nor U21819 (N_21819,N_17157,N_19939);
nor U21820 (N_21820,N_15242,N_19119);
and U21821 (N_21821,N_19602,N_16542);
or U21822 (N_21822,N_15943,N_18599);
xnor U21823 (N_21823,N_19770,N_17362);
xnor U21824 (N_21824,N_18874,N_17485);
and U21825 (N_21825,N_18214,N_16801);
xor U21826 (N_21826,N_18528,N_17202);
xor U21827 (N_21827,N_19401,N_17033);
nor U21828 (N_21828,N_16119,N_16104);
nand U21829 (N_21829,N_19898,N_17754);
and U21830 (N_21830,N_19934,N_18428);
and U21831 (N_21831,N_15153,N_17128);
nand U21832 (N_21832,N_15363,N_17068);
xor U21833 (N_21833,N_17922,N_19113);
nand U21834 (N_21834,N_15880,N_17171);
nand U21835 (N_21835,N_19581,N_19813);
xnor U21836 (N_21836,N_19700,N_15445);
nand U21837 (N_21837,N_16740,N_15908);
xnor U21838 (N_21838,N_16057,N_16908);
nor U21839 (N_21839,N_16122,N_17095);
and U21840 (N_21840,N_17854,N_18740);
nand U21841 (N_21841,N_15032,N_17679);
xor U21842 (N_21842,N_15743,N_18612);
nand U21843 (N_21843,N_19411,N_16997);
xor U21844 (N_21844,N_15584,N_19936);
or U21845 (N_21845,N_18488,N_16657);
nand U21846 (N_21846,N_19230,N_16834);
xnor U21847 (N_21847,N_17796,N_19818);
or U21848 (N_21848,N_18698,N_19643);
or U21849 (N_21849,N_16855,N_17001);
nor U21850 (N_21850,N_15924,N_16602);
or U21851 (N_21851,N_15846,N_17051);
and U21852 (N_21852,N_19328,N_16919);
or U21853 (N_21853,N_18007,N_18232);
and U21854 (N_21854,N_19117,N_19099);
and U21855 (N_21855,N_15384,N_18556);
or U21856 (N_21856,N_19618,N_15239);
and U21857 (N_21857,N_19479,N_17945);
or U21858 (N_21858,N_19588,N_18434);
nand U21859 (N_21859,N_19156,N_18574);
nor U21860 (N_21860,N_16505,N_16244);
xnor U21861 (N_21861,N_16369,N_18549);
nor U21862 (N_21862,N_17603,N_17840);
xor U21863 (N_21863,N_17472,N_18128);
xnor U21864 (N_21864,N_16987,N_17763);
or U21865 (N_21865,N_17020,N_16638);
and U21866 (N_21866,N_16063,N_19282);
or U21867 (N_21867,N_18886,N_18132);
nor U21868 (N_21868,N_18673,N_18504);
nand U21869 (N_21869,N_16706,N_16569);
and U21870 (N_21870,N_17600,N_16624);
nand U21871 (N_21871,N_16482,N_17185);
and U21872 (N_21872,N_17665,N_16659);
nor U21873 (N_21873,N_19394,N_18551);
and U21874 (N_21874,N_19234,N_19174);
and U21875 (N_21875,N_18868,N_19927);
nor U21876 (N_21876,N_18395,N_18952);
nand U21877 (N_21877,N_15759,N_17197);
nor U21878 (N_21878,N_16151,N_18043);
and U21879 (N_21879,N_15948,N_18818);
nor U21880 (N_21880,N_19438,N_18429);
nor U21881 (N_21881,N_18051,N_16484);
or U21882 (N_21882,N_19817,N_18366);
nand U21883 (N_21883,N_18677,N_15960);
xor U21884 (N_21884,N_18891,N_17064);
or U21885 (N_21885,N_18254,N_17049);
and U21886 (N_21886,N_16432,N_17916);
nand U21887 (N_21887,N_18306,N_16947);
or U21888 (N_21888,N_19944,N_17526);
nand U21889 (N_21889,N_15192,N_15411);
and U21890 (N_21890,N_15546,N_15025);
nor U21891 (N_21891,N_17297,N_16732);
xnor U21892 (N_21892,N_16026,N_18290);
nor U21893 (N_21893,N_19991,N_15002);
nand U21894 (N_21894,N_18522,N_17012);
nor U21895 (N_21895,N_15355,N_17104);
xor U21896 (N_21896,N_18632,N_17940);
nand U21897 (N_21897,N_16265,N_19627);
nand U21898 (N_21898,N_15670,N_17072);
xnor U21899 (N_21899,N_18739,N_17044);
or U21900 (N_21900,N_16457,N_19060);
and U21901 (N_21901,N_17629,N_17277);
nand U21902 (N_21902,N_19442,N_17949);
and U21903 (N_21903,N_17215,N_17489);
and U21904 (N_21904,N_19752,N_16286);
xor U21905 (N_21905,N_16899,N_18945);
or U21906 (N_21906,N_15309,N_18415);
nor U21907 (N_21907,N_16840,N_15897);
nor U21908 (N_21908,N_19746,N_18449);
nor U21909 (N_21909,N_15187,N_19942);
nor U21910 (N_21910,N_17060,N_15118);
xnor U21911 (N_21911,N_15291,N_18464);
and U21912 (N_21912,N_19699,N_19608);
xnor U21913 (N_21913,N_16926,N_18880);
nand U21914 (N_21914,N_19097,N_17606);
nor U21915 (N_21915,N_19755,N_18523);
nand U21916 (N_21916,N_19239,N_16055);
nor U21917 (N_21917,N_17682,N_18609);
and U21918 (N_21918,N_18400,N_15416);
and U21919 (N_21919,N_17463,N_16008);
and U21920 (N_21920,N_15655,N_19533);
nand U21921 (N_21921,N_18313,N_16823);
nor U21922 (N_21922,N_17948,N_16588);
nor U21923 (N_21923,N_19859,N_19224);
and U21924 (N_21924,N_19078,N_19908);
and U21925 (N_21925,N_19263,N_15127);
and U21926 (N_21926,N_18842,N_16853);
nor U21927 (N_21927,N_15823,N_18181);
nand U21928 (N_21928,N_17503,N_19023);
or U21929 (N_21929,N_16816,N_18172);
or U21930 (N_21930,N_18233,N_15817);
and U21931 (N_21931,N_15950,N_19556);
and U21932 (N_21932,N_18410,N_18908);
xor U21933 (N_21933,N_15119,N_15568);
or U21934 (N_21934,N_17198,N_18184);
or U21935 (N_21935,N_18989,N_17258);
nand U21936 (N_21936,N_15828,N_15731);
xor U21937 (N_21937,N_15782,N_15143);
and U21938 (N_21938,N_17655,N_19557);
nand U21939 (N_21939,N_15874,N_17604);
xor U21940 (N_21940,N_15463,N_18939);
nor U21941 (N_21941,N_16768,N_15707);
and U21942 (N_21942,N_15132,N_17121);
xor U21943 (N_21943,N_17530,N_18790);
or U21944 (N_21944,N_15922,N_16846);
or U21945 (N_21945,N_18682,N_16021);
nor U21946 (N_21946,N_16582,N_17755);
nor U21947 (N_21947,N_19485,N_15856);
and U21948 (N_21948,N_19283,N_18147);
or U21949 (N_21949,N_17220,N_16035);
or U21950 (N_21950,N_18706,N_19516);
nor U21951 (N_21951,N_18752,N_17853);
nand U21952 (N_21952,N_15487,N_16679);
and U21953 (N_21953,N_18302,N_17276);
and U21954 (N_21954,N_19020,N_17181);
xnor U21955 (N_21955,N_17769,N_17735);
or U21956 (N_21956,N_16209,N_19519);
and U21957 (N_21957,N_15509,N_19232);
nand U21958 (N_21958,N_18656,N_19277);
and U21959 (N_21959,N_15200,N_16717);
and U21960 (N_21960,N_18103,N_16018);
or U21961 (N_21961,N_16342,N_15936);
nand U21962 (N_21962,N_15681,N_18754);
nand U21963 (N_21963,N_17911,N_17549);
nand U21964 (N_21964,N_16563,N_16456);
xor U21965 (N_21965,N_18375,N_17547);
or U21966 (N_21966,N_18865,N_19623);
nor U21967 (N_21967,N_15302,N_15375);
and U21968 (N_21968,N_19184,N_15386);
nor U21969 (N_21969,N_18208,N_19052);
xor U21970 (N_21970,N_19657,N_19269);
xnor U21971 (N_21971,N_17032,N_19747);
nand U21972 (N_21972,N_17315,N_17519);
nor U21973 (N_21973,N_18040,N_18352);
or U21974 (N_21974,N_17067,N_18319);
xor U21975 (N_21975,N_16948,N_17323);
and U21976 (N_21976,N_19783,N_17037);
nor U21977 (N_21977,N_19923,N_15932);
xor U21978 (N_21978,N_15505,N_15234);
and U21979 (N_21979,N_16066,N_17771);
xnor U21980 (N_21980,N_17226,N_19163);
or U21981 (N_21981,N_18299,N_17141);
and U21982 (N_21982,N_16790,N_17097);
nor U21983 (N_21983,N_15554,N_16595);
xnor U21984 (N_21984,N_15696,N_19227);
or U21985 (N_21985,N_17512,N_16910);
nand U21986 (N_21986,N_19247,N_17048);
xor U21987 (N_21987,N_19713,N_15585);
and U21988 (N_21988,N_19427,N_17898);
nand U21989 (N_21989,N_18631,N_19604);
xnor U21990 (N_21990,N_17804,N_15538);
and U21991 (N_21991,N_17382,N_17134);
or U21992 (N_21992,N_19718,N_15752);
or U21993 (N_21993,N_18267,N_19538);
nor U21994 (N_21994,N_16024,N_19330);
xor U21995 (N_21995,N_18421,N_19380);
nand U21996 (N_21996,N_19971,N_17164);
xor U21997 (N_21997,N_15786,N_15159);
xor U21998 (N_21998,N_17636,N_19142);
or U21999 (N_21999,N_16613,N_17910);
nor U22000 (N_22000,N_17955,N_17406);
nor U22001 (N_22001,N_15536,N_16584);
or U22002 (N_22002,N_15998,N_18271);
xnor U22003 (N_22003,N_17745,N_19159);
or U22004 (N_22004,N_15876,N_18197);
or U22005 (N_22005,N_16443,N_18094);
and U22006 (N_22006,N_16398,N_16071);
and U22007 (N_22007,N_19369,N_18529);
or U22008 (N_22008,N_17782,N_18879);
or U22009 (N_22009,N_15586,N_15967);
nor U22010 (N_22010,N_19955,N_19337);
or U22011 (N_22011,N_16412,N_19098);
nand U22012 (N_22012,N_18984,N_15765);
or U22013 (N_22013,N_15461,N_17213);
xor U22014 (N_22014,N_18107,N_15665);
xnor U22015 (N_22015,N_18246,N_16174);
xnor U22016 (N_22016,N_16993,N_16052);
xor U22017 (N_22017,N_16134,N_16142);
and U22018 (N_22018,N_19517,N_15812);
nor U22019 (N_22019,N_17061,N_19354);
and U22020 (N_22020,N_18353,N_18106);
or U22021 (N_22021,N_18665,N_15301);
xor U22022 (N_22022,N_19341,N_17825);
nand U22023 (N_22023,N_19439,N_16519);
or U22024 (N_22024,N_16228,N_19025);
or U22025 (N_22025,N_15425,N_18943);
xnor U22026 (N_22026,N_15819,N_16722);
and U22027 (N_22027,N_18745,N_17446);
and U22028 (N_22028,N_18320,N_19376);
or U22029 (N_22029,N_18177,N_15516);
xor U22030 (N_22030,N_16446,N_16797);
or U22031 (N_22031,N_16536,N_15906);
xnor U22032 (N_22032,N_15601,N_15346);
and U22033 (N_22033,N_16692,N_19022);
nor U22034 (N_22034,N_17678,N_19124);
xnor U22035 (N_22035,N_15547,N_18032);
and U22036 (N_22036,N_16955,N_16715);
nand U22037 (N_22037,N_19929,N_15319);
xor U22038 (N_22038,N_19924,N_17696);
nand U22039 (N_22039,N_16004,N_16438);
or U22040 (N_22040,N_18809,N_18149);
or U22041 (N_22041,N_16194,N_15821);
nor U22042 (N_22042,N_18093,N_18167);
and U22043 (N_22043,N_17046,N_16395);
xor U22044 (N_22044,N_17180,N_16915);
nor U22045 (N_22045,N_15392,N_16337);
xor U22046 (N_22046,N_17766,N_16034);
nand U22047 (N_22047,N_17594,N_17294);
xor U22048 (N_22048,N_16028,N_17031);
and U22049 (N_22049,N_18403,N_16079);
xor U22050 (N_22050,N_16972,N_16463);
or U22051 (N_22051,N_15381,N_19466);
nor U22052 (N_22052,N_16093,N_15956);
nand U22053 (N_22053,N_16580,N_19828);
xor U22054 (N_22054,N_15523,N_15190);
and U22055 (N_22055,N_15071,N_17071);
nor U22056 (N_22056,N_17390,N_17301);
nor U22057 (N_22057,N_15138,N_17976);
nor U22058 (N_22058,N_16264,N_15493);
nand U22059 (N_22059,N_15545,N_17578);
and U22060 (N_22060,N_17768,N_19145);
nand U22061 (N_22061,N_18457,N_16589);
or U22062 (N_22062,N_18779,N_15773);
or U22063 (N_22063,N_18335,N_17069);
or U22064 (N_22064,N_15754,N_17172);
or U22065 (N_22065,N_16532,N_17950);
or U22066 (N_22066,N_17310,N_19858);
and U22067 (N_22067,N_15758,N_15177);
xor U22068 (N_22068,N_18610,N_18911);
nand U22069 (N_22069,N_19034,N_18708);
nor U22070 (N_22070,N_18517,N_18154);
or U22071 (N_22071,N_19288,N_15562);
nand U22072 (N_22072,N_15182,N_17368);
and U22073 (N_22073,N_17400,N_16075);
nand U22074 (N_22074,N_18019,N_18973);
nand U22075 (N_22075,N_15008,N_17505);
and U22076 (N_22076,N_19584,N_19559);
xnor U22077 (N_22077,N_17016,N_16609);
nand U22078 (N_22078,N_18345,N_17077);
nor U22079 (N_22079,N_16932,N_17999);
nand U22080 (N_22080,N_18274,N_18278);
nor U22081 (N_22081,N_19192,N_16200);
xnor U22082 (N_22082,N_18772,N_18498);
nor U22083 (N_22083,N_15409,N_16527);
and U22084 (N_22084,N_15724,N_15628);
xnor U22085 (N_22085,N_15373,N_18422);
nand U22086 (N_22086,N_18858,N_18272);
xnor U22087 (N_22087,N_16555,N_19998);
xor U22088 (N_22088,N_16779,N_15327);
and U22089 (N_22089,N_15883,N_17664);
or U22090 (N_22090,N_19388,N_17643);
xnor U22091 (N_22091,N_15006,N_15304);
nand U22092 (N_22092,N_18282,N_15293);
or U22093 (N_22093,N_17260,N_18919);
nor U22094 (N_22094,N_15213,N_17777);
or U22095 (N_22095,N_19672,N_19226);
xnor U22096 (N_22096,N_15642,N_17450);
xor U22097 (N_22097,N_19462,N_18171);
and U22098 (N_22098,N_16400,N_17360);
or U22099 (N_22099,N_17902,N_18604);
nand U22100 (N_22100,N_18344,N_19033);
or U22101 (N_22101,N_19403,N_18666);
and U22102 (N_22102,N_19318,N_16552);
or U22103 (N_22103,N_18850,N_15646);
or U22104 (N_22104,N_15246,N_17733);
nand U22105 (N_22105,N_19198,N_18229);
xnor U22106 (N_22106,N_19386,N_19138);
nor U22107 (N_22107,N_17923,N_16409);
and U22108 (N_22108,N_17221,N_19310);
nand U22109 (N_22109,N_16821,N_18042);
xnor U22110 (N_22110,N_15644,N_19740);
nand U22111 (N_22111,N_16886,N_17445);
nor U22112 (N_22112,N_17801,N_18808);
nand U22113 (N_22113,N_15194,N_19848);
nor U22114 (N_22114,N_18218,N_15441);
xnor U22115 (N_22115,N_19886,N_18194);
or U22116 (N_22116,N_19799,N_15937);
nand U22117 (N_22117,N_15410,N_15365);
or U22118 (N_22118,N_16690,N_16583);
nand U22119 (N_22119,N_16141,N_19838);
xor U22120 (N_22120,N_19400,N_18951);
nor U22121 (N_22121,N_17823,N_19912);
nor U22122 (N_22122,N_19704,N_16346);
and U22123 (N_22123,N_18211,N_16667);
nor U22124 (N_22124,N_18056,N_17424);
xor U22125 (N_22125,N_18764,N_18806);
nand U22126 (N_22126,N_15458,N_15799);
xnor U22127 (N_22127,N_17893,N_18265);
xnor U22128 (N_22128,N_18371,N_17994);
xor U22129 (N_22129,N_15672,N_16981);
xnor U22130 (N_22130,N_18741,N_16030);
or U22131 (N_22131,N_16674,N_16803);
xnor U22132 (N_22132,N_17290,N_19830);
nor U22133 (N_22133,N_17487,N_15195);
xnor U22134 (N_22134,N_16990,N_16339);
nor U22135 (N_22135,N_19370,N_18404);
and U22136 (N_22136,N_16479,N_16593);
xor U22137 (N_22137,N_15051,N_17809);
and U22138 (N_22138,N_19869,N_16116);
nand U22139 (N_22139,N_19975,N_16475);
xnor U22140 (N_22140,N_19795,N_17355);
and U22141 (N_22141,N_15938,N_16171);
xnor U22142 (N_22142,N_17843,N_19325);
and U22143 (N_22143,N_17623,N_17612);
and U22144 (N_22144,N_16296,N_17767);
and U22145 (N_22145,N_15834,N_19426);
nor U22146 (N_22146,N_17517,N_18873);
and U22147 (N_22147,N_19108,N_15316);
nor U22148 (N_22148,N_16399,N_16377);
or U22149 (N_22149,N_17306,N_16988);
nand U22150 (N_22150,N_15574,N_15258);
or U22151 (N_22151,N_19767,N_19266);
xor U22152 (N_22152,N_16358,N_15934);
nor U22153 (N_22153,N_19463,N_19272);
xnor U22154 (N_22154,N_18416,N_19974);
nor U22155 (N_22155,N_19000,N_18756);
or U22156 (N_22156,N_15096,N_16416);
xnor U22157 (N_22157,N_15951,N_19176);
nand U22158 (N_22158,N_19845,N_18931);
nor U22159 (N_22159,N_16587,N_18394);
nand U22160 (N_22160,N_18226,N_16828);
nand U22161 (N_22161,N_17698,N_18558);
nand U22162 (N_22162,N_16069,N_17284);
nor U22163 (N_22163,N_17561,N_18065);
or U22164 (N_22164,N_19808,N_17053);
nand U22165 (N_22165,N_19551,N_19307);
nor U22166 (N_22166,N_16594,N_16170);
and U22167 (N_22167,N_15641,N_18620);
nand U22168 (N_22168,N_17047,N_19252);
or U22169 (N_22169,N_19743,N_17957);
or U22170 (N_22170,N_18576,N_19024);
and U22171 (N_22171,N_15448,N_15040);
nand U22172 (N_22172,N_18527,N_16754);
nand U22173 (N_22173,N_15576,N_17469);
or U22174 (N_22174,N_18412,N_15318);
nand U22175 (N_22175,N_17093,N_19958);
nor U22176 (N_22176,N_17238,N_19344);
nand U22177 (N_22177,N_16781,N_17652);
xnor U22178 (N_22178,N_17159,N_15657);
and U22179 (N_22179,N_19486,N_19500);
nor U22180 (N_22180,N_18762,N_16931);
xnor U22181 (N_22181,N_16256,N_19027);
nor U22182 (N_22182,N_15862,N_16327);
nor U22183 (N_22183,N_19454,N_17312);
nand U22184 (N_22184,N_16307,N_19218);
and U22185 (N_22185,N_18753,N_18544);
or U22186 (N_22186,N_18050,N_19484);
or U22187 (N_22187,N_16534,N_15206);
or U22188 (N_22188,N_18642,N_19425);
nand U22189 (N_22189,N_17496,N_19270);
and U22190 (N_22190,N_18722,N_16581);
nand U22191 (N_22191,N_15184,N_17461);
and U22192 (N_22192,N_17731,N_15501);
xor U22193 (N_22193,N_17235,N_19621);
or U22194 (N_22194,N_18979,N_17189);
xor U22195 (N_22195,N_15129,N_15594);
or U22196 (N_22196,N_15330,N_19139);
nor U22197 (N_22197,N_16382,N_18796);
xor U22198 (N_22198,N_19387,N_15257);
nor U22199 (N_22199,N_15853,N_18383);
nand U22200 (N_22200,N_18838,N_15098);
or U22201 (N_22201,N_18920,N_15497);
nor U22202 (N_22202,N_16381,N_15423);
nor U22203 (N_22203,N_15789,N_16002);
nor U22204 (N_22204,N_15980,N_18684);
or U22205 (N_22205,N_15353,N_19617);
xnor U22206 (N_22206,N_15263,N_16092);
and U22207 (N_22207,N_15552,N_16898);
and U22208 (N_22208,N_15443,N_16806);
nor U22209 (N_22209,N_15900,N_17475);
and U22210 (N_22210,N_19545,N_19905);
nor U22211 (N_22211,N_19800,N_17083);
nand U22212 (N_22212,N_16418,N_17806);
or U22213 (N_22213,N_16622,N_16312);
nor U22214 (N_22214,N_16303,N_19303);
or U22215 (N_22215,N_19342,N_19682);
xor U22216 (N_22216,N_15605,N_15307);
or U22217 (N_22217,N_18245,N_19948);
nand U22218 (N_22218,N_18231,N_17780);
nor U22219 (N_22219,N_17351,N_18894);
or U22220 (N_22220,N_15158,N_18537);
nor U22221 (N_22221,N_18346,N_15215);
nand U22222 (N_22222,N_18142,N_17567);
or U22223 (N_22223,N_15446,N_19986);
nand U22224 (N_22224,N_16979,N_15211);
nand U22225 (N_22225,N_19541,N_19238);
nand U22226 (N_22226,N_15994,N_15078);
nor U22227 (N_22227,N_19106,N_18972);
and U22228 (N_22228,N_19892,N_18453);
and U22229 (N_22229,N_18435,N_18338);
or U22230 (N_22230,N_17167,N_16943);
xnor U22231 (N_22231,N_16810,N_19840);
nand U22232 (N_22232,N_16946,N_18554);
xor U22233 (N_22233,N_18351,N_16245);
xor U22234 (N_22234,N_18934,N_19716);
or U22235 (N_22235,N_17543,N_16818);
nor U22236 (N_22236,N_15430,N_18068);
or U22237 (N_22237,N_18108,N_19031);
xnor U22238 (N_22238,N_17903,N_16056);
nor U22239 (N_22239,N_15692,N_16745);
nand U22240 (N_22240,N_18066,N_16599);
and U22241 (N_22241,N_18847,N_19474);
nand U22242 (N_22242,N_19963,N_18795);
and U22243 (N_22243,N_16872,N_15666);
or U22244 (N_22244,N_16241,N_17096);
nand U22245 (N_22245,N_19786,N_17560);
nor U22246 (N_22246,N_16428,N_18324);
and U22247 (N_22247,N_18679,N_19200);
and U22248 (N_22248,N_16117,N_15236);
xnor U22249 (N_22249,N_18117,N_15524);
and U22250 (N_22250,N_16277,N_18182);
xnor U22251 (N_22251,N_19954,N_18791);
nand U22252 (N_22252,N_19797,N_17113);
and U22253 (N_22253,N_15361,N_16973);
nor U22254 (N_22254,N_16282,N_16216);
or U22255 (N_22255,N_16500,N_19788);
nand U22256 (N_22256,N_16269,N_15454);
nor U22257 (N_22257,N_17863,N_19243);
nand U22258 (N_22258,N_16903,N_15372);
or U22259 (N_22259,N_15462,N_18349);
xor U22260 (N_22260,N_19850,N_17460);
or U22261 (N_22261,N_18037,N_15380);
nand U22262 (N_22262,N_17844,N_15358);
or U22263 (N_22263,N_19320,N_17883);
nand U22264 (N_22264,N_19170,N_15965);
nor U22265 (N_22265,N_17634,N_17839);
or U22266 (N_22266,N_16348,N_17174);
nand U22267 (N_22267,N_18454,N_17160);
nand U22268 (N_22268,N_17847,N_17440);
xor U22269 (N_22269,N_18657,N_15273);
and U22270 (N_22270,N_19051,N_16335);
nand U22271 (N_22271,N_19781,N_19966);
and U22272 (N_22272,N_16140,N_18516);
and U22273 (N_22273,N_18175,N_16214);
xor U22274 (N_22274,N_16129,N_17405);
xor U22275 (N_22275,N_15850,N_15022);
and U22276 (N_22276,N_17885,N_15571);
xnor U22277 (N_22277,N_18399,N_15014);
nor U22278 (N_22278,N_18484,N_15082);
xnor U22279 (N_22279,N_18339,N_15803);
xnor U22280 (N_22280,N_17653,N_19878);
xnor U22281 (N_22281,N_16788,N_15366);
and U22282 (N_22282,N_19624,N_19591);
nand U22283 (N_22283,N_19882,N_18332);
xnor U22284 (N_22284,N_18622,N_17451);
nand U22285 (N_22285,N_18377,N_18674);
nand U22286 (N_22286,N_19611,N_19129);
nand U22287 (N_22287,N_17621,N_17106);
and U22288 (N_22288,N_16515,N_17799);
xnor U22289 (N_22289,N_18234,N_15149);
xnor U22290 (N_22290,N_16673,N_16401);
xor U22291 (N_22291,N_17835,N_19959);
nand U22292 (N_22292,N_18326,N_19512);
and U22293 (N_22293,N_18661,N_19736);
and U22294 (N_22294,N_18975,N_18723);
nor U22295 (N_22295,N_17579,N_16760);
or U22296 (N_22296,N_17462,N_19809);
and U22297 (N_22297,N_17353,N_15697);
nand U22298 (N_22298,N_15598,N_16849);
nand U22299 (N_22299,N_19314,N_19919);
nand U22300 (N_22300,N_16749,N_18935);
nand U22301 (N_22301,N_16493,N_16144);
nor U22302 (N_22302,N_17590,N_17416);
xor U22303 (N_22303,N_19819,N_16914);
nand U22304 (N_22304,N_19945,N_16111);
or U22305 (N_22305,N_19398,N_15189);
xnor U22306 (N_22306,N_15675,N_19492);
nor U22307 (N_22307,N_18917,N_16721);
and U22308 (N_22308,N_19471,N_15484);
xnor U22309 (N_22309,N_17917,N_15727);
xnor U22310 (N_22310,N_18716,N_15439);
nand U22311 (N_22311,N_16825,N_19217);
and U22312 (N_22312,N_15037,N_19475);
and U22313 (N_22313,N_16088,N_18143);
nand U22314 (N_22314,N_16585,N_18692);
nor U22315 (N_22315,N_18933,N_17062);
nand U22316 (N_22316,N_18978,N_18044);
nor U22317 (N_22317,N_17036,N_16524);
nand U22318 (N_22318,N_18882,N_19444);
and U22319 (N_22319,N_17882,N_17034);
nor U22320 (N_22320,N_18487,N_15050);
or U22321 (N_22321,N_17686,N_17278);
or U22322 (N_22322,N_17066,N_17501);
or U22323 (N_22323,N_15196,N_19820);
nand U22324 (N_22324,N_18643,N_17444);
and U22325 (N_22325,N_18409,N_18856);
nand U22326 (N_22326,N_19067,N_19154);
and U22327 (N_22327,N_18424,N_17960);
and U22328 (N_22328,N_16573,N_15671);
nor U22329 (N_22329,N_15147,N_15863);
nand U22330 (N_22330,N_17580,N_17139);
nor U22331 (N_22331,N_16964,N_15869);
and U22332 (N_22332,N_19284,N_16172);
nor U22333 (N_22333,N_16949,N_15772);
nand U22334 (N_22334,N_18564,N_19572);
and U22335 (N_22335,N_16782,N_17864);
xnor U22336 (N_22336,N_15059,N_15847);
nand U22337 (N_22337,N_18437,N_16772);
and U22338 (N_22338,N_18817,N_17729);
nand U22339 (N_22339,N_17935,N_18520);
nor U22340 (N_22340,N_18531,N_19293);
and U22341 (N_22341,N_17739,N_17585);
xnor U22342 (N_22342,N_15664,N_19309);
xor U22343 (N_22343,N_18837,N_16601);
xnor U22344 (N_22344,N_19316,N_17166);
nand U22345 (N_22345,N_15767,N_16970);
and U22346 (N_22346,N_18884,N_18821);
nor U22347 (N_22347,N_15284,N_18023);
nand U22348 (N_22348,N_18276,N_15010);
xor U22349 (N_22349,N_15004,N_17339);
or U22350 (N_22350,N_16771,N_15248);
and U22351 (N_22351,N_18623,N_18705);
or U22352 (N_22352,N_16822,N_18696);
nand U22353 (N_22353,N_19947,N_16447);
nand U22354 (N_22354,N_16982,N_15326);
xor U22355 (N_22355,N_17073,N_15971);
nand U22356 (N_22356,N_19221,N_15117);
or U22357 (N_22357,N_16773,N_15259);
nand U22358 (N_22358,N_15058,N_15842);
or U22359 (N_22359,N_19798,N_18980);
nor U22360 (N_22360,N_18427,N_19412);
nor U22361 (N_22361,N_17712,N_19630);
xor U22362 (N_22362,N_19487,N_19754);
xnor U22363 (N_22363,N_16322,N_19826);
or U22364 (N_22364,N_16497,N_18131);
nand U22365 (N_22365,N_17732,N_17334);
nor U22366 (N_22366,N_19258,N_15695);
and U22367 (N_22367,N_17575,N_15238);
nor U22368 (N_22368,N_19013,N_16736);
and U22369 (N_22369,N_19926,N_18038);
nor U22370 (N_22370,N_19406,N_17818);
nor U22371 (N_22371,N_17947,N_18035);
nand U22372 (N_22372,N_19100,N_16105);
nor U22373 (N_22373,N_17473,N_17562);
and U22374 (N_22374,N_15210,N_15072);
nor U22375 (N_22375,N_18820,N_18084);
nand U22376 (N_22376,N_16041,N_16212);
and U22377 (N_22377,N_19911,N_17793);
nor U22378 (N_22378,N_15169,N_17075);
nor U22379 (N_22379,N_18116,N_17502);
and U22380 (N_22380,N_17996,N_15214);
or U22381 (N_22381,N_15564,N_17052);
nand U22382 (N_22382,N_16235,N_18621);
nor U22383 (N_22383,N_17702,N_18227);
xor U22384 (N_22384,N_18216,N_16860);
and U22385 (N_22385,N_17136,N_16419);
or U22386 (N_22386,N_16464,N_18250);
and U22387 (N_22387,N_18485,N_15652);
nor U22388 (N_22388,N_15106,N_16384);
xor U22389 (N_22389,N_15360,N_19209);
nor U22390 (N_22390,N_16218,N_15424);
or U22391 (N_22391,N_17091,N_19358);
nand U22392 (N_22392,N_19059,N_18262);
nand U22393 (N_22393,N_18125,N_15095);
nand U22394 (N_22394,N_19852,N_19151);
nor U22395 (N_22395,N_16994,N_15485);
or U22396 (N_22396,N_17486,N_17909);
nand U22397 (N_22397,N_15654,N_17320);
xnor U22398 (N_22398,N_19360,N_17018);
nor U22399 (N_22399,N_18968,N_17694);
and U22400 (N_22400,N_15706,N_18378);
nand U22401 (N_22401,N_19921,N_18089);
xor U22402 (N_22402,N_17193,N_18318);
and U22403 (N_22403,N_17569,N_17300);
or U22404 (N_22404,N_18887,N_17366);
nor U22405 (N_22405,N_17304,N_19267);
xnor U22406 (N_22406,N_15414,N_19001);
and U22407 (N_22407,N_15030,N_17685);
and U22408 (N_22408,N_15981,N_18900);
and U22409 (N_22409,N_18995,N_15164);
nand U22410 (N_22410,N_15898,N_16336);
nand U22411 (N_22411,N_15475,N_16378);
xnor U22412 (N_22412,N_16845,N_15633);
nand U22413 (N_22413,N_17216,N_16866);
or U22414 (N_22414,N_17753,N_16800);
nor U22415 (N_22415,N_19660,N_19641);
or U22416 (N_22416,N_17521,N_15802);
and U22417 (N_22417,N_17975,N_17518);
nor U22418 (N_22418,N_15209,N_18869);
xor U22419 (N_22419,N_15579,N_18750);
or U22420 (N_22420,N_17342,N_18580);
nor U22421 (N_22421,N_19193,N_17467);
xnor U22422 (N_22422,N_15387,N_15931);
xnor U22423 (N_22423,N_17641,N_15060);
and U22424 (N_22424,N_19757,N_15338);
xnor U22425 (N_22425,N_16751,N_19640);
xor U22426 (N_22426,N_17982,N_16072);
nand U22427 (N_22427,N_15308,N_18478);
and U22428 (N_22428,N_15735,N_16976);
or U22429 (N_22429,N_17877,N_15637);
xnor U22430 (N_22430,N_15721,N_17586);
nor U22431 (N_22431,N_18004,N_18814);
xor U22432 (N_22432,N_17076,N_19603);
or U22433 (N_22433,N_18426,N_19932);
nand U22434 (N_22434,N_19554,N_15769);
or U22435 (N_22435,N_19535,N_16238);
xnor U22436 (N_22436,N_19449,N_18058);
or U22437 (N_22437,N_19520,N_15405);
nand U22438 (N_22438,N_15927,N_19599);
xor U22439 (N_22439,N_18627,N_15068);
or U22440 (N_22440,N_19148,N_17380);
xor U22441 (N_22441,N_18239,N_19625);
xnor U22442 (N_22442,N_17815,N_19692);
nor U22443 (N_22443,N_15507,N_18281);
and U22444 (N_22444,N_18373,N_18139);
nor U22445 (N_22445,N_15371,N_17218);
nor U22446 (N_22446,N_16753,N_18055);
nor U22447 (N_22447,N_18702,N_15498);
and U22448 (N_22448,N_16086,N_16596);
or U22449 (N_22449,N_19594,N_17978);
nand U22450 (N_22450,N_17275,N_15667);
nand U22451 (N_22451,N_16488,N_18114);
nor U22452 (N_22452,N_17019,N_16983);
nand U22453 (N_22453,N_16110,N_16364);
nand U22454 (N_22454,N_15328,N_18237);
or U22455 (N_22455,N_15254,N_18802);
and U22456 (N_22456,N_15624,N_18903);
and U22457 (N_22457,N_15225,N_18836);
nand U22458 (N_22458,N_17225,N_19399);
or U22459 (N_22459,N_15933,N_18341);
or U22460 (N_22460,N_15567,N_15221);
xor U22461 (N_22461,N_17085,N_18589);
xnor U22462 (N_22462,N_15612,N_16139);
or U22463 (N_22463,N_15486,N_18778);
or U22464 (N_22464,N_17402,N_16167);
or U22465 (N_22465,N_18736,N_17313);
nor U22466 (N_22466,N_19913,N_16306);
xnor U22467 (N_22467,N_19012,N_18614);
nand U22468 (N_22468,N_18641,N_19015);
xor U22469 (N_22469,N_16203,N_17414);
nand U22470 (N_22470,N_17348,N_17538);
nand U22471 (N_22471,N_15525,N_18625);
xnor U22472 (N_22472,N_18742,N_18571);
xor U22473 (N_22473,N_15168,N_18392);
nor U22474 (N_22474,N_19607,N_19026);
or U22475 (N_22475,N_18922,N_15560);
or U22476 (N_22476,N_19880,N_15070);
and U22477 (N_22477,N_17931,N_18248);
nor U22478 (N_22478,N_19774,N_19109);
or U22479 (N_22479,N_19879,N_17895);
and U22480 (N_22480,N_19348,N_15882);
or U22481 (N_22481,N_19711,N_17805);
nor U22482 (N_22482,N_18663,N_16442);
nand U22483 (N_22483,N_17914,N_15345);
xnor U22484 (N_22484,N_16118,N_19578);
or U22485 (N_22485,N_15625,N_18955);
or U22486 (N_22486,N_17824,N_16615);
or U22487 (N_22487,N_18707,N_15500);
or U22488 (N_22488,N_17493,N_19856);
nor U22489 (N_22489,N_15656,N_18768);
or U22490 (N_22490,N_17591,N_18830);
nor U22491 (N_22491,N_16473,N_15916);
and U22492 (N_22492,N_18910,N_16836);
and U22493 (N_22493,N_16554,N_15871);
or U22494 (N_22494,N_18525,N_15089);
nand U22495 (N_22495,N_19901,N_18810);
nand U22496 (N_22496,N_16799,N_16902);
nor U22497 (N_22497,N_16712,N_18550);
nand U22498 (N_22498,N_16971,N_19350);
and U22499 (N_22499,N_16796,N_16300);
nor U22500 (N_22500,N_18264,N_19081);
and U22501 (N_22501,N_19296,N_19214);
nor U22502 (N_22502,N_18483,N_18390);
xor U22503 (N_22503,N_18516,N_15049);
nor U22504 (N_22504,N_15233,N_18978);
nand U22505 (N_22505,N_19927,N_16908);
nand U22506 (N_22506,N_15143,N_18340);
and U22507 (N_22507,N_19020,N_17254);
and U22508 (N_22508,N_19291,N_15725);
nand U22509 (N_22509,N_17495,N_19176);
and U22510 (N_22510,N_18047,N_17223);
and U22511 (N_22511,N_16653,N_19794);
xnor U22512 (N_22512,N_15807,N_15596);
nor U22513 (N_22513,N_18672,N_19153);
nor U22514 (N_22514,N_16208,N_16607);
nor U22515 (N_22515,N_16170,N_18322);
and U22516 (N_22516,N_15832,N_18380);
or U22517 (N_22517,N_15041,N_16229);
and U22518 (N_22518,N_19130,N_15138);
nor U22519 (N_22519,N_19842,N_17715);
xnor U22520 (N_22520,N_15716,N_19502);
nand U22521 (N_22521,N_16204,N_18606);
nand U22522 (N_22522,N_17419,N_18039);
xor U22523 (N_22523,N_15065,N_15255);
and U22524 (N_22524,N_19796,N_18470);
nand U22525 (N_22525,N_17069,N_17692);
and U22526 (N_22526,N_19647,N_18013);
and U22527 (N_22527,N_18713,N_18734);
nor U22528 (N_22528,N_15500,N_19679);
or U22529 (N_22529,N_16477,N_18435);
xnor U22530 (N_22530,N_19244,N_19816);
nand U22531 (N_22531,N_18451,N_18098);
or U22532 (N_22532,N_18186,N_15122);
xor U22533 (N_22533,N_19847,N_19504);
xnor U22534 (N_22534,N_19782,N_18091);
and U22535 (N_22535,N_16278,N_15663);
or U22536 (N_22536,N_19926,N_15352);
or U22537 (N_22537,N_19608,N_18740);
xor U22538 (N_22538,N_17355,N_16772);
xor U22539 (N_22539,N_15751,N_19736);
or U22540 (N_22540,N_19529,N_19815);
and U22541 (N_22541,N_15103,N_19355);
and U22542 (N_22542,N_19166,N_19684);
nor U22543 (N_22543,N_15427,N_15644);
nor U22544 (N_22544,N_17035,N_18277);
nand U22545 (N_22545,N_15588,N_17779);
nand U22546 (N_22546,N_17861,N_19883);
nand U22547 (N_22547,N_16483,N_17418);
and U22548 (N_22548,N_16511,N_16917);
nor U22549 (N_22549,N_15233,N_19102);
nand U22550 (N_22550,N_17129,N_16569);
xor U22551 (N_22551,N_16400,N_19665);
or U22552 (N_22552,N_15863,N_18528);
nor U22553 (N_22553,N_18199,N_17565);
and U22554 (N_22554,N_18839,N_15570);
and U22555 (N_22555,N_18129,N_15736);
xnor U22556 (N_22556,N_17011,N_17326);
xor U22557 (N_22557,N_15614,N_17483);
xor U22558 (N_22558,N_16308,N_19689);
nor U22559 (N_22559,N_16842,N_16980);
and U22560 (N_22560,N_17147,N_17020);
or U22561 (N_22561,N_15141,N_15040);
nor U22562 (N_22562,N_17297,N_19744);
nor U22563 (N_22563,N_18984,N_15735);
or U22564 (N_22564,N_16476,N_18908);
xor U22565 (N_22565,N_15799,N_15809);
nand U22566 (N_22566,N_15479,N_16490);
and U22567 (N_22567,N_16696,N_17424);
nor U22568 (N_22568,N_15738,N_19683);
nand U22569 (N_22569,N_19320,N_17041);
xor U22570 (N_22570,N_18633,N_18724);
xor U22571 (N_22571,N_16806,N_16404);
nand U22572 (N_22572,N_17401,N_18885);
nand U22573 (N_22573,N_18752,N_15450);
and U22574 (N_22574,N_15889,N_15266);
nor U22575 (N_22575,N_19916,N_18924);
nand U22576 (N_22576,N_17850,N_19127);
nor U22577 (N_22577,N_19694,N_15918);
nand U22578 (N_22578,N_15503,N_16179);
nand U22579 (N_22579,N_17688,N_16432);
nor U22580 (N_22580,N_16194,N_17689);
nand U22581 (N_22581,N_19282,N_16870);
nor U22582 (N_22582,N_15417,N_18002);
nand U22583 (N_22583,N_19392,N_17667);
or U22584 (N_22584,N_18378,N_16876);
and U22585 (N_22585,N_15120,N_16082);
nand U22586 (N_22586,N_16658,N_16176);
xor U22587 (N_22587,N_15729,N_15818);
nand U22588 (N_22588,N_16659,N_17345);
and U22589 (N_22589,N_16481,N_17071);
nand U22590 (N_22590,N_17458,N_15808);
xnor U22591 (N_22591,N_16341,N_19715);
and U22592 (N_22592,N_19175,N_16177);
xor U22593 (N_22593,N_18160,N_18386);
xor U22594 (N_22594,N_19278,N_15566);
xor U22595 (N_22595,N_17610,N_16962);
nand U22596 (N_22596,N_17266,N_15226);
or U22597 (N_22597,N_17445,N_18094);
nor U22598 (N_22598,N_15953,N_16729);
or U22599 (N_22599,N_18992,N_16515);
or U22600 (N_22600,N_17138,N_17949);
nand U22601 (N_22601,N_15568,N_18983);
nand U22602 (N_22602,N_17176,N_17246);
xor U22603 (N_22603,N_15539,N_15773);
nand U22604 (N_22604,N_18709,N_19814);
xnor U22605 (N_22605,N_17001,N_19362);
nor U22606 (N_22606,N_16125,N_17009);
or U22607 (N_22607,N_19794,N_17837);
or U22608 (N_22608,N_19724,N_16856);
or U22609 (N_22609,N_18722,N_19832);
nor U22610 (N_22610,N_19236,N_19103);
nand U22611 (N_22611,N_18363,N_18399);
nor U22612 (N_22612,N_19926,N_17241);
or U22613 (N_22613,N_17421,N_15199);
nor U22614 (N_22614,N_19249,N_15839);
and U22615 (N_22615,N_15538,N_19600);
nand U22616 (N_22616,N_18827,N_16172);
xor U22617 (N_22617,N_15487,N_18895);
nor U22618 (N_22618,N_17535,N_18872);
xnor U22619 (N_22619,N_17202,N_19339);
nor U22620 (N_22620,N_15598,N_18758);
or U22621 (N_22621,N_16646,N_15435);
or U22622 (N_22622,N_15350,N_15110);
and U22623 (N_22623,N_16537,N_18656);
or U22624 (N_22624,N_16398,N_16761);
xor U22625 (N_22625,N_17455,N_15323);
xnor U22626 (N_22626,N_16493,N_15049);
nand U22627 (N_22627,N_17869,N_18363);
or U22628 (N_22628,N_17461,N_17596);
xor U22629 (N_22629,N_17306,N_16696);
and U22630 (N_22630,N_15755,N_18374);
nand U22631 (N_22631,N_19276,N_18993);
nand U22632 (N_22632,N_15585,N_16386);
nor U22633 (N_22633,N_17485,N_16684);
or U22634 (N_22634,N_16432,N_17642);
nor U22635 (N_22635,N_15852,N_15851);
or U22636 (N_22636,N_18276,N_15079);
and U22637 (N_22637,N_18706,N_15420);
or U22638 (N_22638,N_18938,N_18445);
or U22639 (N_22639,N_16941,N_17294);
nor U22640 (N_22640,N_17194,N_15856);
nand U22641 (N_22641,N_16245,N_17245);
xor U22642 (N_22642,N_16963,N_18356);
or U22643 (N_22643,N_19679,N_19863);
xor U22644 (N_22644,N_19344,N_16850);
and U22645 (N_22645,N_19170,N_17089);
nand U22646 (N_22646,N_17690,N_15776);
and U22647 (N_22647,N_16460,N_15451);
xor U22648 (N_22648,N_15281,N_19164);
or U22649 (N_22649,N_15899,N_18159);
and U22650 (N_22650,N_18465,N_15789);
xor U22651 (N_22651,N_17727,N_19694);
xnor U22652 (N_22652,N_17955,N_15648);
or U22653 (N_22653,N_17706,N_19805);
nand U22654 (N_22654,N_15423,N_17640);
or U22655 (N_22655,N_16812,N_16407);
nand U22656 (N_22656,N_19716,N_16295);
nor U22657 (N_22657,N_15781,N_17090);
nor U22658 (N_22658,N_16178,N_15199);
nor U22659 (N_22659,N_17191,N_17175);
nor U22660 (N_22660,N_18858,N_16129);
nand U22661 (N_22661,N_18368,N_19547);
or U22662 (N_22662,N_17462,N_18409);
and U22663 (N_22663,N_19460,N_15761);
nor U22664 (N_22664,N_18061,N_16396);
xor U22665 (N_22665,N_15341,N_17202);
or U22666 (N_22666,N_17886,N_15377);
or U22667 (N_22667,N_16259,N_16574);
xnor U22668 (N_22668,N_15233,N_15799);
xor U22669 (N_22669,N_19848,N_17440);
and U22670 (N_22670,N_15656,N_18396);
xnor U22671 (N_22671,N_18337,N_17258);
and U22672 (N_22672,N_18397,N_17240);
nand U22673 (N_22673,N_16758,N_17560);
or U22674 (N_22674,N_18681,N_17701);
and U22675 (N_22675,N_17413,N_17375);
or U22676 (N_22676,N_18879,N_16214);
nand U22677 (N_22677,N_17993,N_19862);
xor U22678 (N_22678,N_15586,N_19547);
nand U22679 (N_22679,N_18649,N_15009);
or U22680 (N_22680,N_19077,N_19078);
or U22681 (N_22681,N_17144,N_16813);
nand U22682 (N_22682,N_17228,N_15257);
or U22683 (N_22683,N_16031,N_17397);
nand U22684 (N_22684,N_15495,N_15578);
or U22685 (N_22685,N_18104,N_18112);
xor U22686 (N_22686,N_19406,N_15248);
nor U22687 (N_22687,N_18151,N_19051);
nor U22688 (N_22688,N_16701,N_16837);
and U22689 (N_22689,N_17247,N_19006);
xor U22690 (N_22690,N_15217,N_17058);
and U22691 (N_22691,N_17751,N_15265);
nor U22692 (N_22692,N_15101,N_17279);
nor U22693 (N_22693,N_19085,N_17616);
nand U22694 (N_22694,N_18229,N_19421);
nor U22695 (N_22695,N_16530,N_17076);
or U22696 (N_22696,N_16373,N_15432);
nand U22697 (N_22697,N_17801,N_15010);
or U22698 (N_22698,N_19730,N_17346);
nor U22699 (N_22699,N_19325,N_15640);
nand U22700 (N_22700,N_18926,N_19378);
nand U22701 (N_22701,N_16581,N_17503);
or U22702 (N_22702,N_19394,N_18439);
xnor U22703 (N_22703,N_18407,N_18440);
or U22704 (N_22704,N_15367,N_15507);
nand U22705 (N_22705,N_16471,N_15724);
or U22706 (N_22706,N_19894,N_15446);
xnor U22707 (N_22707,N_18360,N_18397);
and U22708 (N_22708,N_19430,N_18507);
nand U22709 (N_22709,N_17972,N_19498);
and U22710 (N_22710,N_15287,N_17659);
nand U22711 (N_22711,N_15231,N_19023);
and U22712 (N_22712,N_15949,N_18799);
or U22713 (N_22713,N_15510,N_18516);
nor U22714 (N_22714,N_17951,N_18760);
or U22715 (N_22715,N_15382,N_19216);
nand U22716 (N_22716,N_19250,N_15723);
or U22717 (N_22717,N_17255,N_19619);
xnor U22718 (N_22718,N_18190,N_19229);
or U22719 (N_22719,N_19622,N_17827);
nand U22720 (N_22720,N_15578,N_15991);
nand U22721 (N_22721,N_16467,N_18059);
and U22722 (N_22722,N_15061,N_18786);
nor U22723 (N_22723,N_17463,N_16865);
xor U22724 (N_22724,N_17033,N_18706);
xor U22725 (N_22725,N_16599,N_17192);
nand U22726 (N_22726,N_19819,N_16458);
nand U22727 (N_22727,N_18050,N_18195);
and U22728 (N_22728,N_17168,N_19956);
or U22729 (N_22729,N_18823,N_16539);
and U22730 (N_22730,N_18066,N_16750);
or U22731 (N_22731,N_19812,N_19142);
nor U22732 (N_22732,N_19125,N_18494);
nor U22733 (N_22733,N_18773,N_15154);
xor U22734 (N_22734,N_18973,N_15879);
and U22735 (N_22735,N_15687,N_18382);
nand U22736 (N_22736,N_18951,N_15711);
xnor U22737 (N_22737,N_16467,N_19126);
or U22738 (N_22738,N_18092,N_18041);
nor U22739 (N_22739,N_16965,N_18126);
and U22740 (N_22740,N_18376,N_16243);
nand U22741 (N_22741,N_19055,N_19445);
or U22742 (N_22742,N_19976,N_19931);
xor U22743 (N_22743,N_19081,N_17780);
and U22744 (N_22744,N_15398,N_16549);
and U22745 (N_22745,N_18948,N_18928);
nor U22746 (N_22746,N_19489,N_17305);
and U22747 (N_22747,N_17974,N_19920);
and U22748 (N_22748,N_18844,N_15841);
nor U22749 (N_22749,N_16441,N_17784);
nand U22750 (N_22750,N_19619,N_19036);
and U22751 (N_22751,N_17976,N_15642);
or U22752 (N_22752,N_15271,N_15964);
or U22753 (N_22753,N_17076,N_16252);
or U22754 (N_22754,N_15570,N_16524);
or U22755 (N_22755,N_16875,N_15068);
and U22756 (N_22756,N_16034,N_15774);
and U22757 (N_22757,N_15534,N_15563);
nand U22758 (N_22758,N_18340,N_15546);
xor U22759 (N_22759,N_15457,N_16202);
and U22760 (N_22760,N_17718,N_16395);
xor U22761 (N_22761,N_17752,N_15146);
xnor U22762 (N_22762,N_19268,N_19841);
or U22763 (N_22763,N_17370,N_17188);
nand U22764 (N_22764,N_16897,N_18627);
or U22765 (N_22765,N_19230,N_18560);
nor U22766 (N_22766,N_18336,N_15952);
or U22767 (N_22767,N_19210,N_18147);
and U22768 (N_22768,N_16700,N_16085);
xor U22769 (N_22769,N_15506,N_16419);
and U22770 (N_22770,N_16291,N_15791);
or U22771 (N_22771,N_19775,N_18724);
xor U22772 (N_22772,N_17629,N_17845);
and U22773 (N_22773,N_15524,N_16683);
or U22774 (N_22774,N_19685,N_17596);
nand U22775 (N_22775,N_16214,N_17101);
nor U22776 (N_22776,N_17458,N_17585);
nor U22777 (N_22777,N_16983,N_17601);
or U22778 (N_22778,N_15638,N_15004);
nand U22779 (N_22779,N_17795,N_17870);
or U22780 (N_22780,N_18051,N_15886);
nor U22781 (N_22781,N_19838,N_19893);
or U22782 (N_22782,N_18438,N_19222);
nor U22783 (N_22783,N_19722,N_17968);
xnor U22784 (N_22784,N_18017,N_15310);
nor U22785 (N_22785,N_18325,N_19423);
or U22786 (N_22786,N_19693,N_19262);
nand U22787 (N_22787,N_17521,N_17750);
xnor U22788 (N_22788,N_17319,N_15964);
nor U22789 (N_22789,N_15547,N_17915);
and U22790 (N_22790,N_15739,N_17766);
or U22791 (N_22791,N_16767,N_19215);
nand U22792 (N_22792,N_16789,N_15675);
nand U22793 (N_22793,N_16891,N_17115);
or U22794 (N_22794,N_16402,N_16321);
nor U22795 (N_22795,N_18849,N_15317);
nor U22796 (N_22796,N_18080,N_16026);
xor U22797 (N_22797,N_16059,N_15598);
xnor U22798 (N_22798,N_15556,N_16828);
nor U22799 (N_22799,N_16608,N_18263);
and U22800 (N_22800,N_16370,N_16374);
nor U22801 (N_22801,N_19625,N_18298);
or U22802 (N_22802,N_17627,N_19751);
and U22803 (N_22803,N_17905,N_17454);
nand U22804 (N_22804,N_15249,N_19074);
and U22805 (N_22805,N_19147,N_15064);
nand U22806 (N_22806,N_16319,N_17186);
xnor U22807 (N_22807,N_18724,N_19169);
or U22808 (N_22808,N_18850,N_19552);
nor U22809 (N_22809,N_15125,N_15535);
nor U22810 (N_22810,N_19358,N_19060);
nor U22811 (N_22811,N_15649,N_17918);
and U22812 (N_22812,N_15440,N_17845);
xor U22813 (N_22813,N_18923,N_19403);
nand U22814 (N_22814,N_19101,N_16267);
xnor U22815 (N_22815,N_19622,N_18430);
or U22816 (N_22816,N_18541,N_17798);
nor U22817 (N_22817,N_19450,N_19642);
or U22818 (N_22818,N_17954,N_15560);
and U22819 (N_22819,N_19306,N_15536);
or U22820 (N_22820,N_19107,N_18118);
xor U22821 (N_22821,N_16287,N_17555);
and U22822 (N_22822,N_15680,N_18135);
xor U22823 (N_22823,N_18317,N_17374);
xor U22824 (N_22824,N_18239,N_19169);
xor U22825 (N_22825,N_15579,N_15130);
nand U22826 (N_22826,N_18688,N_16055);
and U22827 (N_22827,N_18655,N_15991);
nand U22828 (N_22828,N_19536,N_15899);
xor U22829 (N_22829,N_19981,N_16541);
or U22830 (N_22830,N_17106,N_19278);
nand U22831 (N_22831,N_19602,N_17983);
and U22832 (N_22832,N_19649,N_19766);
or U22833 (N_22833,N_16681,N_18182);
and U22834 (N_22834,N_17496,N_18705);
or U22835 (N_22835,N_17272,N_17468);
or U22836 (N_22836,N_15800,N_17232);
and U22837 (N_22837,N_18086,N_16206);
nor U22838 (N_22838,N_19348,N_17590);
nor U22839 (N_22839,N_15524,N_16013);
and U22840 (N_22840,N_15730,N_19031);
and U22841 (N_22841,N_17838,N_17865);
nor U22842 (N_22842,N_19052,N_17734);
nor U22843 (N_22843,N_17416,N_19417);
xnor U22844 (N_22844,N_18130,N_15948);
or U22845 (N_22845,N_18326,N_19650);
nand U22846 (N_22846,N_19470,N_19903);
nor U22847 (N_22847,N_18146,N_18601);
nand U22848 (N_22848,N_15429,N_18293);
nor U22849 (N_22849,N_17980,N_16000);
nand U22850 (N_22850,N_16575,N_17943);
nor U22851 (N_22851,N_18204,N_15503);
or U22852 (N_22852,N_16470,N_17763);
or U22853 (N_22853,N_15704,N_16774);
nor U22854 (N_22854,N_19782,N_18331);
nand U22855 (N_22855,N_18482,N_16064);
xor U22856 (N_22856,N_15933,N_15835);
nand U22857 (N_22857,N_15686,N_17406);
nand U22858 (N_22858,N_17160,N_16534);
or U22859 (N_22859,N_17719,N_15981);
nand U22860 (N_22860,N_15164,N_17616);
and U22861 (N_22861,N_15301,N_19567);
xnor U22862 (N_22862,N_18966,N_19363);
xor U22863 (N_22863,N_17288,N_15098);
or U22864 (N_22864,N_19148,N_17347);
and U22865 (N_22865,N_17200,N_18439);
nand U22866 (N_22866,N_17364,N_15335);
nand U22867 (N_22867,N_19311,N_15271);
nor U22868 (N_22868,N_17503,N_15953);
nor U22869 (N_22869,N_19646,N_19267);
nand U22870 (N_22870,N_18379,N_15092);
nand U22871 (N_22871,N_18463,N_19635);
nand U22872 (N_22872,N_15493,N_19063);
nand U22873 (N_22873,N_18376,N_17940);
or U22874 (N_22874,N_18297,N_18909);
xor U22875 (N_22875,N_18033,N_15303);
and U22876 (N_22876,N_15014,N_16249);
and U22877 (N_22877,N_19861,N_16672);
or U22878 (N_22878,N_18181,N_17353);
xnor U22879 (N_22879,N_18932,N_15106);
xnor U22880 (N_22880,N_17697,N_17204);
nor U22881 (N_22881,N_19661,N_18559);
or U22882 (N_22882,N_19776,N_15099);
and U22883 (N_22883,N_18136,N_16701);
nand U22884 (N_22884,N_17102,N_15066);
nand U22885 (N_22885,N_15608,N_19491);
nand U22886 (N_22886,N_19681,N_18382);
and U22887 (N_22887,N_16118,N_19130);
or U22888 (N_22888,N_17648,N_17969);
nand U22889 (N_22889,N_16017,N_17387);
xor U22890 (N_22890,N_17478,N_16804);
or U22891 (N_22891,N_19637,N_15725);
xnor U22892 (N_22892,N_18149,N_19284);
or U22893 (N_22893,N_19883,N_19220);
or U22894 (N_22894,N_17056,N_15752);
xor U22895 (N_22895,N_19137,N_19016);
and U22896 (N_22896,N_18881,N_19259);
or U22897 (N_22897,N_16193,N_16857);
xnor U22898 (N_22898,N_17297,N_16786);
nand U22899 (N_22899,N_19330,N_18116);
or U22900 (N_22900,N_15883,N_19576);
nand U22901 (N_22901,N_18745,N_18465);
or U22902 (N_22902,N_16701,N_16189);
and U22903 (N_22903,N_15125,N_15621);
and U22904 (N_22904,N_15330,N_17671);
or U22905 (N_22905,N_18518,N_17334);
and U22906 (N_22906,N_16083,N_17114);
xor U22907 (N_22907,N_16359,N_17116);
nor U22908 (N_22908,N_19911,N_15195);
and U22909 (N_22909,N_17378,N_18384);
nand U22910 (N_22910,N_19616,N_15666);
nand U22911 (N_22911,N_19549,N_17765);
and U22912 (N_22912,N_17923,N_18568);
nand U22913 (N_22913,N_15539,N_19327);
nand U22914 (N_22914,N_16423,N_16511);
xnor U22915 (N_22915,N_17507,N_15869);
nand U22916 (N_22916,N_17874,N_16511);
or U22917 (N_22917,N_18453,N_16164);
nor U22918 (N_22918,N_16169,N_19886);
nor U22919 (N_22919,N_15378,N_15738);
nand U22920 (N_22920,N_18078,N_16079);
or U22921 (N_22921,N_17280,N_16799);
and U22922 (N_22922,N_18964,N_16310);
or U22923 (N_22923,N_16855,N_19758);
xor U22924 (N_22924,N_16264,N_18542);
nor U22925 (N_22925,N_16480,N_19808);
nor U22926 (N_22926,N_16876,N_16847);
and U22927 (N_22927,N_15623,N_17877);
xnor U22928 (N_22928,N_16031,N_15554);
xor U22929 (N_22929,N_19939,N_17206);
nand U22930 (N_22930,N_16884,N_19665);
xor U22931 (N_22931,N_15382,N_17183);
and U22932 (N_22932,N_16997,N_15187);
nor U22933 (N_22933,N_15462,N_15595);
and U22934 (N_22934,N_19396,N_18257);
nand U22935 (N_22935,N_16695,N_15191);
xnor U22936 (N_22936,N_19876,N_17963);
or U22937 (N_22937,N_15537,N_17853);
nand U22938 (N_22938,N_19755,N_16419);
nand U22939 (N_22939,N_15358,N_17102);
nand U22940 (N_22940,N_15635,N_16234);
xor U22941 (N_22941,N_16860,N_19455);
nand U22942 (N_22942,N_17997,N_16051);
xor U22943 (N_22943,N_17256,N_17327);
and U22944 (N_22944,N_18327,N_15605);
nor U22945 (N_22945,N_16339,N_16265);
nand U22946 (N_22946,N_19687,N_18825);
and U22947 (N_22947,N_15332,N_15116);
or U22948 (N_22948,N_18760,N_18579);
nand U22949 (N_22949,N_19824,N_18250);
or U22950 (N_22950,N_15355,N_15088);
nor U22951 (N_22951,N_16169,N_15371);
or U22952 (N_22952,N_18222,N_15593);
and U22953 (N_22953,N_15816,N_15710);
nand U22954 (N_22954,N_19567,N_19793);
nor U22955 (N_22955,N_17772,N_17079);
and U22956 (N_22956,N_15545,N_15434);
nor U22957 (N_22957,N_16684,N_17421);
or U22958 (N_22958,N_18954,N_15335);
xnor U22959 (N_22959,N_19867,N_17758);
nor U22960 (N_22960,N_19146,N_17509);
nor U22961 (N_22961,N_18455,N_15255);
or U22962 (N_22962,N_15235,N_17896);
nand U22963 (N_22963,N_19596,N_18019);
nor U22964 (N_22964,N_17027,N_19041);
xnor U22965 (N_22965,N_17221,N_15921);
xor U22966 (N_22966,N_17111,N_19718);
or U22967 (N_22967,N_15649,N_15806);
nand U22968 (N_22968,N_18238,N_18883);
nor U22969 (N_22969,N_16114,N_15617);
nand U22970 (N_22970,N_15174,N_19327);
or U22971 (N_22971,N_15493,N_15708);
nor U22972 (N_22972,N_19084,N_15258);
nor U22973 (N_22973,N_15201,N_17330);
and U22974 (N_22974,N_17130,N_15471);
or U22975 (N_22975,N_17237,N_16513);
xor U22976 (N_22976,N_17638,N_16449);
nand U22977 (N_22977,N_17703,N_16697);
and U22978 (N_22978,N_15517,N_16580);
nand U22979 (N_22979,N_19528,N_18368);
nor U22980 (N_22980,N_17774,N_16561);
and U22981 (N_22981,N_17261,N_18154);
or U22982 (N_22982,N_18549,N_16914);
or U22983 (N_22983,N_17332,N_18252);
nand U22984 (N_22984,N_19760,N_16307);
and U22985 (N_22985,N_15559,N_15982);
nand U22986 (N_22986,N_19564,N_18423);
nor U22987 (N_22987,N_16560,N_18152);
xor U22988 (N_22988,N_17203,N_18083);
or U22989 (N_22989,N_18267,N_15619);
and U22990 (N_22990,N_15646,N_15952);
and U22991 (N_22991,N_16730,N_15924);
nor U22992 (N_22992,N_17947,N_16979);
xor U22993 (N_22993,N_15245,N_18457);
nor U22994 (N_22994,N_17968,N_18302);
nor U22995 (N_22995,N_15282,N_15243);
nand U22996 (N_22996,N_15081,N_15274);
nand U22997 (N_22997,N_16755,N_15800);
and U22998 (N_22998,N_19906,N_18765);
and U22999 (N_22999,N_18691,N_19913);
nand U23000 (N_23000,N_19917,N_15607);
nor U23001 (N_23001,N_17562,N_17245);
or U23002 (N_23002,N_16776,N_18444);
or U23003 (N_23003,N_16966,N_17958);
and U23004 (N_23004,N_16082,N_15032);
xor U23005 (N_23005,N_16175,N_18799);
nor U23006 (N_23006,N_15087,N_16765);
nor U23007 (N_23007,N_15586,N_15224);
nor U23008 (N_23008,N_17363,N_16558);
or U23009 (N_23009,N_19735,N_15524);
or U23010 (N_23010,N_16368,N_16227);
xnor U23011 (N_23011,N_15709,N_18872);
nand U23012 (N_23012,N_15409,N_18612);
nor U23013 (N_23013,N_15039,N_19299);
nor U23014 (N_23014,N_18213,N_16559);
xnor U23015 (N_23015,N_19520,N_16204);
nand U23016 (N_23016,N_17977,N_15586);
nand U23017 (N_23017,N_17762,N_18808);
nor U23018 (N_23018,N_18153,N_17603);
nor U23019 (N_23019,N_19206,N_17740);
nand U23020 (N_23020,N_15742,N_16839);
nand U23021 (N_23021,N_18943,N_18647);
and U23022 (N_23022,N_19879,N_16930);
nor U23023 (N_23023,N_18875,N_16352);
nand U23024 (N_23024,N_17907,N_16664);
or U23025 (N_23025,N_18728,N_19503);
nand U23026 (N_23026,N_16304,N_19063);
and U23027 (N_23027,N_16851,N_19336);
nor U23028 (N_23028,N_19233,N_16293);
and U23029 (N_23029,N_15624,N_15275);
nand U23030 (N_23030,N_19220,N_17186);
nor U23031 (N_23031,N_18940,N_17886);
xnor U23032 (N_23032,N_19971,N_17029);
and U23033 (N_23033,N_15753,N_16029);
and U23034 (N_23034,N_16784,N_15050);
xnor U23035 (N_23035,N_19727,N_18226);
xor U23036 (N_23036,N_16542,N_15914);
nor U23037 (N_23037,N_16533,N_19580);
xnor U23038 (N_23038,N_15564,N_16783);
nor U23039 (N_23039,N_19347,N_18860);
or U23040 (N_23040,N_15893,N_19130);
nor U23041 (N_23041,N_16413,N_15832);
or U23042 (N_23042,N_18246,N_18804);
nor U23043 (N_23043,N_16252,N_16838);
and U23044 (N_23044,N_16236,N_18953);
xnor U23045 (N_23045,N_18274,N_16781);
xor U23046 (N_23046,N_15759,N_15771);
xnor U23047 (N_23047,N_18136,N_19925);
nand U23048 (N_23048,N_16610,N_16313);
nand U23049 (N_23049,N_17260,N_19613);
xnor U23050 (N_23050,N_19757,N_16439);
or U23051 (N_23051,N_15531,N_18651);
and U23052 (N_23052,N_19252,N_18233);
xor U23053 (N_23053,N_16195,N_15200);
xnor U23054 (N_23054,N_15013,N_18051);
and U23055 (N_23055,N_19897,N_19483);
or U23056 (N_23056,N_19482,N_17207);
nand U23057 (N_23057,N_19904,N_18245);
and U23058 (N_23058,N_17707,N_18677);
xnor U23059 (N_23059,N_18801,N_16585);
nand U23060 (N_23060,N_19421,N_15401);
xor U23061 (N_23061,N_17390,N_15894);
and U23062 (N_23062,N_19919,N_16393);
nand U23063 (N_23063,N_15076,N_17826);
and U23064 (N_23064,N_15794,N_16795);
nand U23065 (N_23065,N_17007,N_19211);
or U23066 (N_23066,N_17965,N_17430);
xnor U23067 (N_23067,N_17085,N_17643);
and U23068 (N_23068,N_19869,N_17004);
nor U23069 (N_23069,N_17099,N_19153);
xor U23070 (N_23070,N_15916,N_19408);
or U23071 (N_23071,N_16101,N_16701);
and U23072 (N_23072,N_19010,N_16328);
and U23073 (N_23073,N_17851,N_18150);
nand U23074 (N_23074,N_16622,N_16836);
or U23075 (N_23075,N_17916,N_19410);
and U23076 (N_23076,N_17163,N_19504);
and U23077 (N_23077,N_19278,N_16076);
xor U23078 (N_23078,N_18334,N_15275);
nor U23079 (N_23079,N_15002,N_17767);
or U23080 (N_23080,N_18933,N_18156);
or U23081 (N_23081,N_16605,N_15474);
and U23082 (N_23082,N_16030,N_19187);
or U23083 (N_23083,N_15202,N_17333);
or U23084 (N_23084,N_16646,N_18413);
xor U23085 (N_23085,N_18409,N_15181);
and U23086 (N_23086,N_17981,N_18730);
nor U23087 (N_23087,N_19413,N_15990);
xnor U23088 (N_23088,N_15429,N_15201);
nand U23089 (N_23089,N_18269,N_19387);
nor U23090 (N_23090,N_18579,N_19331);
or U23091 (N_23091,N_19362,N_15391);
and U23092 (N_23092,N_18903,N_18707);
or U23093 (N_23093,N_16945,N_18867);
nand U23094 (N_23094,N_15807,N_19551);
nor U23095 (N_23095,N_15048,N_17668);
nand U23096 (N_23096,N_17635,N_19621);
and U23097 (N_23097,N_17754,N_17009);
or U23098 (N_23098,N_19149,N_18582);
or U23099 (N_23099,N_17929,N_15928);
or U23100 (N_23100,N_15039,N_17335);
nand U23101 (N_23101,N_18464,N_18446);
and U23102 (N_23102,N_17429,N_18946);
and U23103 (N_23103,N_18630,N_19770);
nand U23104 (N_23104,N_17388,N_19372);
or U23105 (N_23105,N_15827,N_15002);
xor U23106 (N_23106,N_16741,N_17272);
nor U23107 (N_23107,N_19165,N_18713);
and U23108 (N_23108,N_16659,N_17238);
nor U23109 (N_23109,N_16738,N_19987);
and U23110 (N_23110,N_17252,N_17522);
xor U23111 (N_23111,N_18840,N_16079);
or U23112 (N_23112,N_19914,N_19274);
nand U23113 (N_23113,N_18703,N_17676);
xor U23114 (N_23114,N_16034,N_19218);
or U23115 (N_23115,N_16806,N_15154);
nor U23116 (N_23116,N_18875,N_16694);
nand U23117 (N_23117,N_18406,N_17782);
nor U23118 (N_23118,N_15033,N_17941);
or U23119 (N_23119,N_16740,N_15867);
nand U23120 (N_23120,N_16430,N_19474);
or U23121 (N_23121,N_17271,N_19494);
nor U23122 (N_23122,N_19804,N_16592);
or U23123 (N_23123,N_16301,N_18426);
xor U23124 (N_23124,N_18137,N_18737);
nor U23125 (N_23125,N_18349,N_16276);
and U23126 (N_23126,N_19027,N_15768);
nor U23127 (N_23127,N_17021,N_18773);
or U23128 (N_23128,N_17162,N_17503);
nand U23129 (N_23129,N_15650,N_17107);
nand U23130 (N_23130,N_15493,N_15372);
or U23131 (N_23131,N_15963,N_17555);
nor U23132 (N_23132,N_18752,N_17235);
or U23133 (N_23133,N_16441,N_17984);
nand U23134 (N_23134,N_19654,N_19463);
or U23135 (N_23135,N_19323,N_19457);
or U23136 (N_23136,N_17719,N_15481);
and U23137 (N_23137,N_18524,N_16818);
and U23138 (N_23138,N_16408,N_17623);
or U23139 (N_23139,N_16958,N_18974);
nand U23140 (N_23140,N_15851,N_18143);
nand U23141 (N_23141,N_18481,N_16971);
xnor U23142 (N_23142,N_19823,N_17183);
nand U23143 (N_23143,N_18615,N_18458);
or U23144 (N_23144,N_15368,N_17106);
nor U23145 (N_23145,N_15351,N_18034);
nand U23146 (N_23146,N_18401,N_16916);
nor U23147 (N_23147,N_19896,N_16998);
and U23148 (N_23148,N_16685,N_18179);
nand U23149 (N_23149,N_17910,N_19631);
nand U23150 (N_23150,N_15233,N_19178);
or U23151 (N_23151,N_15597,N_15255);
or U23152 (N_23152,N_18810,N_16139);
xor U23153 (N_23153,N_17097,N_18630);
nor U23154 (N_23154,N_17847,N_18292);
xnor U23155 (N_23155,N_19003,N_17856);
or U23156 (N_23156,N_16485,N_16069);
and U23157 (N_23157,N_19630,N_18288);
xor U23158 (N_23158,N_17297,N_18177);
xor U23159 (N_23159,N_15123,N_18660);
and U23160 (N_23160,N_18536,N_15688);
or U23161 (N_23161,N_15492,N_15498);
and U23162 (N_23162,N_15706,N_19259);
and U23163 (N_23163,N_18476,N_16991);
or U23164 (N_23164,N_15191,N_15631);
xnor U23165 (N_23165,N_18472,N_15385);
xnor U23166 (N_23166,N_15737,N_19311);
nand U23167 (N_23167,N_18767,N_17115);
and U23168 (N_23168,N_15234,N_19873);
xnor U23169 (N_23169,N_15436,N_18891);
xnor U23170 (N_23170,N_18722,N_18780);
nand U23171 (N_23171,N_15137,N_16555);
nand U23172 (N_23172,N_19828,N_19066);
xnor U23173 (N_23173,N_19473,N_16007);
and U23174 (N_23174,N_16192,N_19255);
and U23175 (N_23175,N_18745,N_15236);
xnor U23176 (N_23176,N_17009,N_16885);
nand U23177 (N_23177,N_16302,N_15844);
nand U23178 (N_23178,N_19656,N_15945);
nor U23179 (N_23179,N_16612,N_15244);
and U23180 (N_23180,N_17592,N_18627);
or U23181 (N_23181,N_16036,N_15950);
nor U23182 (N_23182,N_17438,N_18040);
nor U23183 (N_23183,N_17233,N_16794);
nor U23184 (N_23184,N_19331,N_17608);
and U23185 (N_23185,N_19790,N_17729);
nand U23186 (N_23186,N_16449,N_17977);
and U23187 (N_23187,N_16366,N_15700);
nor U23188 (N_23188,N_18104,N_17647);
and U23189 (N_23189,N_19861,N_17467);
nand U23190 (N_23190,N_16986,N_17555);
nand U23191 (N_23191,N_18829,N_17999);
and U23192 (N_23192,N_18864,N_15818);
and U23193 (N_23193,N_17348,N_16573);
and U23194 (N_23194,N_16744,N_15825);
nor U23195 (N_23195,N_15138,N_17742);
nor U23196 (N_23196,N_16662,N_18916);
xor U23197 (N_23197,N_16871,N_19615);
nand U23198 (N_23198,N_19857,N_17491);
xor U23199 (N_23199,N_18060,N_16058);
nor U23200 (N_23200,N_16218,N_18818);
nand U23201 (N_23201,N_16316,N_19044);
and U23202 (N_23202,N_16626,N_15988);
nand U23203 (N_23203,N_17093,N_19055);
xnor U23204 (N_23204,N_18844,N_17112);
and U23205 (N_23205,N_17447,N_19948);
nand U23206 (N_23206,N_15235,N_16119);
nor U23207 (N_23207,N_18693,N_17040);
or U23208 (N_23208,N_18724,N_15773);
nand U23209 (N_23209,N_17279,N_15170);
nand U23210 (N_23210,N_15257,N_15523);
xnor U23211 (N_23211,N_16360,N_19581);
and U23212 (N_23212,N_16167,N_17972);
and U23213 (N_23213,N_16793,N_16525);
xor U23214 (N_23214,N_19170,N_16439);
nand U23215 (N_23215,N_16879,N_17946);
and U23216 (N_23216,N_19291,N_17754);
xnor U23217 (N_23217,N_16752,N_18612);
nor U23218 (N_23218,N_18272,N_15026);
xnor U23219 (N_23219,N_17291,N_16294);
or U23220 (N_23220,N_18443,N_15476);
or U23221 (N_23221,N_17496,N_18404);
and U23222 (N_23222,N_17081,N_17027);
or U23223 (N_23223,N_17585,N_16795);
or U23224 (N_23224,N_15227,N_16210);
and U23225 (N_23225,N_18121,N_18973);
xor U23226 (N_23226,N_17736,N_15916);
and U23227 (N_23227,N_17002,N_19711);
xor U23228 (N_23228,N_16147,N_17606);
nand U23229 (N_23229,N_15002,N_18378);
nor U23230 (N_23230,N_17752,N_18013);
nand U23231 (N_23231,N_16506,N_18556);
and U23232 (N_23232,N_19920,N_17851);
nand U23233 (N_23233,N_16293,N_17199);
or U23234 (N_23234,N_19433,N_17180);
nand U23235 (N_23235,N_15515,N_16728);
nand U23236 (N_23236,N_16301,N_18272);
or U23237 (N_23237,N_15769,N_16099);
xnor U23238 (N_23238,N_19747,N_16758);
xor U23239 (N_23239,N_18706,N_19560);
and U23240 (N_23240,N_19941,N_19363);
nand U23241 (N_23241,N_17689,N_19314);
or U23242 (N_23242,N_15792,N_18565);
and U23243 (N_23243,N_18308,N_17789);
or U23244 (N_23244,N_19222,N_17176);
nand U23245 (N_23245,N_15990,N_15550);
nand U23246 (N_23246,N_15597,N_18133);
or U23247 (N_23247,N_19956,N_19081);
xor U23248 (N_23248,N_17920,N_19420);
nand U23249 (N_23249,N_15283,N_17108);
nor U23250 (N_23250,N_16896,N_17725);
and U23251 (N_23251,N_16617,N_17218);
xor U23252 (N_23252,N_16459,N_18541);
xnor U23253 (N_23253,N_19581,N_19580);
xnor U23254 (N_23254,N_18406,N_19703);
xor U23255 (N_23255,N_18797,N_17588);
nor U23256 (N_23256,N_18485,N_17148);
xor U23257 (N_23257,N_19118,N_15982);
or U23258 (N_23258,N_18979,N_17421);
or U23259 (N_23259,N_18039,N_16344);
or U23260 (N_23260,N_16471,N_15643);
nand U23261 (N_23261,N_16585,N_19020);
or U23262 (N_23262,N_17639,N_17488);
nor U23263 (N_23263,N_18634,N_15358);
xnor U23264 (N_23264,N_16518,N_19060);
or U23265 (N_23265,N_15180,N_15216);
nand U23266 (N_23266,N_15077,N_18489);
nor U23267 (N_23267,N_15279,N_18081);
xor U23268 (N_23268,N_16009,N_15965);
nand U23269 (N_23269,N_15070,N_18490);
nand U23270 (N_23270,N_19970,N_19561);
nor U23271 (N_23271,N_18693,N_17133);
and U23272 (N_23272,N_19852,N_16084);
nor U23273 (N_23273,N_16721,N_18368);
or U23274 (N_23274,N_19902,N_19598);
xnor U23275 (N_23275,N_19644,N_15544);
and U23276 (N_23276,N_18702,N_19233);
xor U23277 (N_23277,N_17657,N_19927);
nor U23278 (N_23278,N_19715,N_19224);
nand U23279 (N_23279,N_17651,N_17220);
or U23280 (N_23280,N_18900,N_17611);
nor U23281 (N_23281,N_16171,N_17645);
and U23282 (N_23282,N_17279,N_16160);
xnor U23283 (N_23283,N_15048,N_16163);
and U23284 (N_23284,N_18757,N_15599);
xnor U23285 (N_23285,N_18691,N_15607);
xnor U23286 (N_23286,N_19060,N_19284);
and U23287 (N_23287,N_18597,N_18797);
xnor U23288 (N_23288,N_16594,N_16216);
nor U23289 (N_23289,N_15175,N_17285);
nand U23290 (N_23290,N_16727,N_18338);
xor U23291 (N_23291,N_17715,N_16206);
nand U23292 (N_23292,N_19356,N_16666);
xnor U23293 (N_23293,N_16498,N_17845);
nor U23294 (N_23294,N_18057,N_15301);
nand U23295 (N_23295,N_19769,N_18793);
or U23296 (N_23296,N_17240,N_15389);
and U23297 (N_23297,N_16950,N_18758);
or U23298 (N_23298,N_16826,N_17930);
and U23299 (N_23299,N_19008,N_16940);
and U23300 (N_23300,N_15583,N_19420);
or U23301 (N_23301,N_19253,N_16223);
and U23302 (N_23302,N_15668,N_17567);
nor U23303 (N_23303,N_19493,N_17961);
or U23304 (N_23304,N_19062,N_17132);
nand U23305 (N_23305,N_19024,N_19553);
nand U23306 (N_23306,N_19642,N_18682);
and U23307 (N_23307,N_16913,N_17878);
or U23308 (N_23308,N_15483,N_18604);
nand U23309 (N_23309,N_17164,N_18968);
and U23310 (N_23310,N_19108,N_16347);
nand U23311 (N_23311,N_18968,N_17318);
or U23312 (N_23312,N_18582,N_16147);
or U23313 (N_23313,N_19313,N_19341);
or U23314 (N_23314,N_15595,N_17235);
nand U23315 (N_23315,N_15580,N_18631);
and U23316 (N_23316,N_16911,N_16721);
nand U23317 (N_23317,N_17347,N_17788);
nor U23318 (N_23318,N_16029,N_16207);
nor U23319 (N_23319,N_17989,N_16193);
nand U23320 (N_23320,N_18054,N_17567);
nand U23321 (N_23321,N_18787,N_17727);
xnor U23322 (N_23322,N_18603,N_15718);
nand U23323 (N_23323,N_18662,N_19258);
xnor U23324 (N_23324,N_17862,N_15802);
and U23325 (N_23325,N_18622,N_16276);
and U23326 (N_23326,N_17965,N_19115);
or U23327 (N_23327,N_15276,N_19755);
nor U23328 (N_23328,N_16379,N_15550);
and U23329 (N_23329,N_17924,N_17655);
nor U23330 (N_23330,N_18347,N_19037);
and U23331 (N_23331,N_18661,N_18091);
or U23332 (N_23332,N_19310,N_17242);
nand U23333 (N_23333,N_16109,N_19305);
or U23334 (N_23334,N_15441,N_18128);
nor U23335 (N_23335,N_18179,N_16279);
xor U23336 (N_23336,N_15956,N_15090);
and U23337 (N_23337,N_17772,N_16589);
or U23338 (N_23338,N_18825,N_15287);
or U23339 (N_23339,N_19075,N_19204);
nor U23340 (N_23340,N_19556,N_17665);
or U23341 (N_23341,N_15589,N_18800);
xor U23342 (N_23342,N_15715,N_17208);
nand U23343 (N_23343,N_18913,N_18201);
or U23344 (N_23344,N_18838,N_19235);
nor U23345 (N_23345,N_19197,N_17326);
and U23346 (N_23346,N_19055,N_16124);
nand U23347 (N_23347,N_17030,N_16681);
nand U23348 (N_23348,N_18822,N_16220);
and U23349 (N_23349,N_18688,N_17049);
or U23350 (N_23350,N_19710,N_16397);
nor U23351 (N_23351,N_19706,N_19845);
and U23352 (N_23352,N_16679,N_15198);
or U23353 (N_23353,N_16249,N_18204);
nor U23354 (N_23354,N_15600,N_15147);
and U23355 (N_23355,N_17618,N_19434);
xnor U23356 (N_23356,N_17525,N_19912);
nand U23357 (N_23357,N_17805,N_18622);
xor U23358 (N_23358,N_16988,N_18050);
nand U23359 (N_23359,N_15843,N_16951);
nor U23360 (N_23360,N_17932,N_18434);
or U23361 (N_23361,N_16287,N_19383);
nand U23362 (N_23362,N_19597,N_18187);
xnor U23363 (N_23363,N_17209,N_16247);
xnor U23364 (N_23364,N_17767,N_17871);
or U23365 (N_23365,N_19208,N_16894);
nand U23366 (N_23366,N_17547,N_18363);
and U23367 (N_23367,N_19649,N_16156);
xnor U23368 (N_23368,N_18421,N_15708);
or U23369 (N_23369,N_19365,N_15773);
xnor U23370 (N_23370,N_18578,N_16056);
xnor U23371 (N_23371,N_15540,N_17722);
nor U23372 (N_23372,N_16708,N_17225);
nor U23373 (N_23373,N_19175,N_16746);
and U23374 (N_23374,N_18921,N_17815);
nor U23375 (N_23375,N_19480,N_16320);
nor U23376 (N_23376,N_18745,N_19757);
or U23377 (N_23377,N_16574,N_17215);
or U23378 (N_23378,N_18562,N_17491);
nor U23379 (N_23379,N_16880,N_19547);
or U23380 (N_23380,N_19147,N_19285);
xnor U23381 (N_23381,N_15978,N_15476);
nand U23382 (N_23382,N_17896,N_19121);
and U23383 (N_23383,N_15542,N_16559);
xor U23384 (N_23384,N_18030,N_15175);
xor U23385 (N_23385,N_15874,N_15230);
nor U23386 (N_23386,N_18075,N_17690);
or U23387 (N_23387,N_18077,N_19899);
or U23388 (N_23388,N_19963,N_18377);
or U23389 (N_23389,N_19679,N_18763);
nor U23390 (N_23390,N_17496,N_18663);
and U23391 (N_23391,N_16649,N_19318);
nand U23392 (N_23392,N_15260,N_16992);
and U23393 (N_23393,N_19973,N_15108);
xnor U23394 (N_23394,N_19156,N_19313);
nand U23395 (N_23395,N_16959,N_15274);
xor U23396 (N_23396,N_17057,N_17308);
nand U23397 (N_23397,N_18865,N_19121);
or U23398 (N_23398,N_16876,N_15251);
or U23399 (N_23399,N_19477,N_17570);
or U23400 (N_23400,N_18547,N_19931);
xnor U23401 (N_23401,N_18108,N_17173);
nor U23402 (N_23402,N_19779,N_18017);
nor U23403 (N_23403,N_17430,N_18732);
nand U23404 (N_23404,N_15273,N_19845);
xnor U23405 (N_23405,N_19314,N_16664);
xor U23406 (N_23406,N_19490,N_19212);
nor U23407 (N_23407,N_16153,N_15953);
xor U23408 (N_23408,N_19806,N_16347);
xor U23409 (N_23409,N_19924,N_18569);
nand U23410 (N_23410,N_15482,N_17543);
and U23411 (N_23411,N_18537,N_19248);
nand U23412 (N_23412,N_19738,N_18158);
and U23413 (N_23413,N_16825,N_19459);
nor U23414 (N_23414,N_19180,N_15787);
and U23415 (N_23415,N_19674,N_18727);
nand U23416 (N_23416,N_18658,N_15630);
nand U23417 (N_23417,N_18408,N_16875);
nor U23418 (N_23418,N_15795,N_16993);
or U23419 (N_23419,N_18651,N_17871);
or U23420 (N_23420,N_18392,N_17818);
xor U23421 (N_23421,N_17004,N_16862);
xnor U23422 (N_23422,N_19091,N_18150);
nand U23423 (N_23423,N_15972,N_18600);
or U23424 (N_23424,N_16647,N_18102);
or U23425 (N_23425,N_16397,N_16963);
nor U23426 (N_23426,N_19046,N_19957);
and U23427 (N_23427,N_16194,N_15798);
nand U23428 (N_23428,N_16953,N_16548);
xnor U23429 (N_23429,N_19363,N_18411);
and U23430 (N_23430,N_15538,N_18588);
nand U23431 (N_23431,N_15170,N_19789);
xor U23432 (N_23432,N_16128,N_17871);
and U23433 (N_23433,N_16216,N_16437);
nand U23434 (N_23434,N_19499,N_17088);
xor U23435 (N_23435,N_16849,N_19924);
xor U23436 (N_23436,N_17802,N_19160);
or U23437 (N_23437,N_19240,N_15160);
nand U23438 (N_23438,N_19403,N_16145);
xnor U23439 (N_23439,N_19954,N_16670);
nand U23440 (N_23440,N_19558,N_19785);
and U23441 (N_23441,N_18997,N_16035);
nor U23442 (N_23442,N_19500,N_15506);
nand U23443 (N_23443,N_16850,N_16302);
or U23444 (N_23444,N_19432,N_17717);
nand U23445 (N_23445,N_15239,N_17312);
nor U23446 (N_23446,N_19925,N_15069);
xnor U23447 (N_23447,N_17262,N_18785);
nand U23448 (N_23448,N_17190,N_15382);
or U23449 (N_23449,N_15066,N_16322);
xor U23450 (N_23450,N_17159,N_18497);
or U23451 (N_23451,N_17138,N_17222);
nor U23452 (N_23452,N_18313,N_15178);
xnor U23453 (N_23453,N_19590,N_17353);
or U23454 (N_23454,N_18244,N_19478);
and U23455 (N_23455,N_16171,N_17558);
or U23456 (N_23456,N_15533,N_16522);
and U23457 (N_23457,N_18867,N_19496);
or U23458 (N_23458,N_17192,N_17197);
nand U23459 (N_23459,N_17912,N_18869);
and U23460 (N_23460,N_18345,N_19644);
nor U23461 (N_23461,N_19996,N_16714);
and U23462 (N_23462,N_16751,N_19433);
and U23463 (N_23463,N_17988,N_19875);
nand U23464 (N_23464,N_15409,N_19185);
nand U23465 (N_23465,N_15380,N_18473);
nor U23466 (N_23466,N_18591,N_18305);
xor U23467 (N_23467,N_15216,N_15355);
xnor U23468 (N_23468,N_15009,N_15422);
xor U23469 (N_23469,N_15891,N_15758);
xnor U23470 (N_23470,N_16926,N_19492);
nand U23471 (N_23471,N_16883,N_16706);
and U23472 (N_23472,N_18614,N_15821);
or U23473 (N_23473,N_18959,N_15685);
or U23474 (N_23474,N_15373,N_16136);
nand U23475 (N_23475,N_18759,N_16349);
xnor U23476 (N_23476,N_19136,N_18855);
or U23477 (N_23477,N_18766,N_15242);
and U23478 (N_23478,N_19814,N_15564);
or U23479 (N_23479,N_15371,N_18453);
nand U23480 (N_23480,N_18034,N_16285);
xnor U23481 (N_23481,N_19776,N_15705);
nand U23482 (N_23482,N_17325,N_18216);
or U23483 (N_23483,N_18273,N_19446);
xor U23484 (N_23484,N_17282,N_16431);
nor U23485 (N_23485,N_15207,N_16430);
xor U23486 (N_23486,N_19794,N_18227);
and U23487 (N_23487,N_15773,N_19999);
nor U23488 (N_23488,N_17102,N_17632);
nor U23489 (N_23489,N_18467,N_16648);
xnor U23490 (N_23490,N_15640,N_15716);
xor U23491 (N_23491,N_17464,N_15164);
xor U23492 (N_23492,N_19055,N_15171);
and U23493 (N_23493,N_15148,N_18707);
nand U23494 (N_23494,N_16893,N_18966);
xor U23495 (N_23495,N_18883,N_17153);
nor U23496 (N_23496,N_19283,N_17450);
nand U23497 (N_23497,N_17672,N_15765);
nor U23498 (N_23498,N_15589,N_17973);
nor U23499 (N_23499,N_16016,N_18698);
nor U23500 (N_23500,N_19666,N_19078);
and U23501 (N_23501,N_18577,N_17504);
nand U23502 (N_23502,N_18308,N_15413);
and U23503 (N_23503,N_15047,N_19043);
or U23504 (N_23504,N_16354,N_18567);
and U23505 (N_23505,N_16312,N_18432);
and U23506 (N_23506,N_15603,N_18204);
nand U23507 (N_23507,N_17082,N_15777);
and U23508 (N_23508,N_16717,N_19834);
nor U23509 (N_23509,N_15902,N_17506);
and U23510 (N_23510,N_18149,N_16925);
and U23511 (N_23511,N_16857,N_19611);
xor U23512 (N_23512,N_19780,N_17664);
nor U23513 (N_23513,N_17258,N_16232);
or U23514 (N_23514,N_19409,N_15029);
nand U23515 (N_23515,N_16025,N_19229);
nor U23516 (N_23516,N_17018,N_19119);
and U23517 (N_23517,N_15300,N_17479);
and U23518 (N_23518,N_18091,N_18688);
nor U23519 (N_23519,N_17424,N_17013);
or U23520 (N_23520,N_18261,N_19217);
xnor U23521 (N_23521,N_19026,N_15399);
xnor U23522 (N_23522,N_18311,N_17782);
nand U23523 (N_23523,N_19984,N_15222);
nor U23524 (N_23524,N_19706,N_17553);
and U23525 (N_23525,N_16251,N_17376);
or U23526 (N_23526,N_18701,N_18326);
nand U23527 (N_23527,N_15906,N_19981);
and U23528 (N_23528,N_15403,N_17825);
and U23529 (N_23529,N_15060,N_18383);
xor U23530 (N_23530,N_19982,N_17360);
or U23531 (N_23531,N_16200,N_16254);
nand U23532 (N_23532,N_18433,N_19832);
and U23533 (N_23533,N_15319,N_17974);
nand U23534 (N_23534,N_18663,N_19292);
xnor U23535 (N_23535,N_16672,N_17139);
nand U23536 (N_23536,N_16369,N_17231);
and U23537 (N_23537,N_19500,N_16140);
nor U23538 (N_23538,N_17740,N_18102);
or U23539 (N_23539,N_19976,N_17047);
xnor U23540 (N_23540,N_17677,N_16284);
and U23541 (N_23541,N_18094,N_18689);
nor U23542 (N_23542,N_16332,N_15097);
xnor U23543 (N_23543,N_15117,N_15926);
nor U23544 (N_23544,N_16855,N_17895);
or U23545 (N_23545,N_19850,N_17435);
nor U23546 (N_23546,N_16730,N_16009);
or U23547 (N_23547,N_16774,N_17831);
nor U23548 (N_23548,N_17385,N_17710);
xnor U23549 (N_23549,N_19369,N_19552);
nand U23550 (N_23550,N_17505,N_15704);
xor U23551 (N_23551,N_18738,N_18545);
or U23552 (N_23552,N_19757,N_18128);
xnor U23553 (N_23553,N_16861,N_15354);
and U23554 (N_23554,N_15771,N_19694);
nor U23555 (N_23555,N_16769,N_18804);
and U23556 (N_23556,N_17498,N_17869);
nand U23557 (N_23557,N_15869,N_19930);
xor U23558 (N_23558,N_18296,N_17513);
or U23559 (N_23559,N_16978,N_16173);
or U23560 (N_23560,N_18567,N_19932);
or U23561 (N_23561,N_17552,N_19518);
and U23562 (N_23562,N_19024,N_19891);
or U23563 (N_23563,N_17471,N_19362);
nand U23564 (N_23564,N_17779,N_19832);
nand U23565 (N_23565,N_16131,N_16474);
nand U23566 (N_23566,N_15851,N_16671);
nand U23567 (N_23567,N_17111,N_16556);
nor U23568 (N_23568,N_19159,N_18739);
or U23569 (N_23569,N_15456,N_15338);
and U23570 (N_23570,N_19482,N_17804);
nor U23571 (N_23571,N_17700,N_15431);
nor U23572 (N_23572,N_18458,N_19694);
nand U23573 (N_23573,N_17703,N_19014);
nor U23574 (N_23574,N_19207,N_17469);
or U23575 (N_23575,N_18589,N_18874);
nor U23576 (N_23576,N_19535,N_16550);
and U23577 (N_23577,N_18498,N_19499);
and U23578 (N_23578,N_16061,N_16334);
or U23579 (N_23579,N_15096,N_17351);
nor U23580 (N_23580,N_18863,N_15972);
and U23581 (N_23581,N_16582,N_16370);
nor U23582 (N_23582,N_19467,N_18925);
or U23583 (N_23583,N_16430,N_15530);
xnor U23584 (N_23584,N_17180,N_18142);
nand U23585 (N_23585,N_15410,N_19367);
and U23586 (N_23586,N_15806,N_16080);
xnor U23587 (N_23587,N_18541,N_19370);
nor U23588 (N_23588,N_18079,N_15528);
xnor U23589 (N_23589,N_19875,N_15915);
xnor U23590 (N_23590,N_19577,N_16318);
xnor U23591 (N_23591,N_19416,N_17718);
xnor U23592 (N_23592,N_19007,N_19772);
and U23593 (N_23593,N_16122,N_19345);
xnor U23594 (N_23594,N_19739,N_15073);
nand U23595 (N_23595,N_18345,N_19502);
nand U23596 (N_23596,N_17624,N_18464);
nor U23597 (N_23597,N_17477,N_19691);
or U23598 (N_23598,N_15011,N_18964);
and U23599 (N_23599,N_19406,N_18520);
xor U23600 (N_23600,N_16733,N_17683);
nor U23601 (N_23601,N_18161,N_18663);
xor U23602 (N_23602,N_15399,N_16427);
nor U23603 (N_23603,N_16285,N_18157);
nand U23604 (N_23604,N_16292,N_19459);
nand U23605 (N_23605,N_17251,N_19021);
nor U23606 (N_23606,N_17111,N_18381);
or U23607 (N_23607,N_15483,N_16348);
nor U23608 (N_23608,N_16842,N_19896);
nand U23609 (N_23609,N_17048,N_17625);
nor U23610 (N_23610,N_16610,N_19032);
nor U23611 (N_23611,N_19908,N_18746);
and U23612 (N_23612,N_16655,N_19497);
nand U23613 (N_23613,N_16686,N_18565);
or U23614 (N_23614,N_19067,N_17947);
xor U23615 (N_23615,N_17698,N_15904);
and U23616 (N_23616,N_15468,N_17275);
nand U23617 (N_23617,N_17152,N_16943);
xnor U23618 (N_23618,N_16622,N_16489);
nor U23619 (N_23619,N_18676,N_18425);
nand U23620 (N_23620,N_16381,N_17730);
nand U23621 (N_23621,N_16465,N_17668);
nand U23622 (N_23622,N_17446,N_15442);
xor U23623 (N_23623,N_16280,N_19079);
xnor U23624 (N_23624,N_19311,N_15685);
nor U23625 (N_23625,N_17525,N_16785);
or U23626 (N_23626,N_16518,N_19788);
xnor U23627 (N_23627,N_15537,N_18424);
xor U23628 (N_23628,N_18177,N_19473);
nor U23629 (N_23629,N_16746,N_19003);
and U23630 (N_23630,N_15607,N_19152);
nor U23631 (N_23631,N_15887,N_15431);
nor U23632 (N_23632,N_19679,N_17587);
nor U23633 (N_23633,N_16705,N_18388);
xor U23634 (N_23634,N_15849,N_17954);
xnor U23635 (N_23635,N_18626,N_15484);
nand U23636 (N_23636,N_16548,N_15813);
or U23637 (N_23637,N_15668,N_17860);
or U23638 (N_23638,N_16423,N_16922);
nor U23639 (N_23639,N_15473,N_15737);
and U23640 (N_23640,N_19373,N_16274);
and U23641 (N_23641,N_15622,N_18662);
nor U23642 (N_23642,N_16888,N_16916);
and U23643 (N_23643,N_19364,N_16885);
xnor U23644 (N_23644,N_16165,N_18931);
xnor U23645 (N_23645,N_15751,N_17904);
xnor U23646 (N_23646,N_17066,N_15189);
nand U23647 (N_23647,N_18793,N_19987);
nor U23648 (N_23648,N_16695,N_18701);
nand U23649 (N_23649,N_16187,N_17180);
nor U23650 (N_23650,N_15984,N_16413);
and U23651 (N_23651,N_18812,N_19974);
nor U23652 (N_23652,N_18887,N_15291);
nand U23653 (N_23653,N_16343,N_17437);
nor U23654 (N_23654,N_17997,N_18090);
nand U23655 (N_23655,N_18240,N_19614);
nor U23656 (N_23656,N_19016,N_17590);
and U23657 (N_23657,N_16641,N_17543);
or U23658 (N_23658,N_17984,N_18660);
and U23659 (N_23659,N_19247,N_18307);
nor U23660 (N_23660,N_17876,N_17863);
nor U23661 (N_23661,N_16580,N_16069);
nor U23662 (N_23662,N_18120,N_18785);
and U23663 (N_23663,N_16118,N_18070);
xor U23664 (N_23664,N_17576,N_16909);
and U23665 (N_23665,N_18602,N_17498);
or U23666 (N_23666,N_16097,N_15688);
nand U23667 (N_23667,N_15832,N_15941);
or U23668 (N_23668,N_19693,N_18380);
nand U23669 (N_23669,N_15757,N_18596);
or U23670 (N_23670,N_19446,N_17392);
and U23671 (N_23671,N_17951,N_15964);
nor U23672 (N_23672,N_16438,N_15378);
nand U23673 (N_23673,N_19223,N_17181);
and U23674 (N_23674,N_16916,N_16857);
nand U23675 (N_23675,N_19543,N_18648);
xnor U23676 (N_23676,N_19252,N_19746);
xnor U23677 (N_23677,N_17092,N_15604);
xnor U23678 (N_23678,N_18527,N_16131);
xor U23679 (N_23679,N_16603,N_15995);
xor U23680 (N_23680,N_15312,N_19808);
xnor U23681 (N_23681,N_15973,N_16028);
xnor U23682 (N_23682,N_16276,N_19511);
xnor U23683 (N_23683,N_16972,N_17991);
xor U23684 (N_23684,N_15620,N_17744);
and U23685 (N_23685,N_15358,N_17517);
and U23686 (N_23686,N_17361,N_17789);
or U23687 (N_23687,N_16273,N_15813);
or U23688 (N_23688,N_16889,N_15693);
nand U23689 (N_23689,N_15393,N_16073);
and U23690 (N_23690,N_19320,N_19472);
and U23691 (N_23691,N_16769,N_16775);
and U23692 (N_23692,N_18056,N_17537);
or U23693 (N_23693,N_19400,N_16041);
nor U23694 (N_23694,N_19195,N_15785);
or U23695 (N_23695,N_15752,N_17493);
or U23696 (N_23696,N_18954,N_19113);
nor U23697 (N_23697,N_16615,N_15702);
nor U23698 (N_23698,N_17616,N_16016);
xor U23699 (N_23699,N_15276,N_17031);
nor U23700 (N_23700,N_18826,N_15235);
or U23701 (N_23701,N_17134,N_17268);
nand U23702 (N_23702,N_18785,N_19606);
xor U23703 (N_23703,N_15921,N_18890);
xnor U23704 (N_23704,N_19230,N_19803);
nand U23705 (N_23705,N_16499,N_15874);
nor U23706 (N_23706,N_15239,N_19587);
nand U23707 (N_23707,N_17975,N_15280);
or U23708 (N_23708,N_15731,N_18416);
nor U23709 (N_23709,N_19829,N_17007);
xor U23710 (N_23710,N_16471,N_18839);
or U23711 (N_23711,N_18933,N_18644);
xnor U23712 (N_23712,N_18254,N_15265);
xnor U23713 (N_23713,N_16168,N_18832);
or U23714 (N_23714,N_16434,N_15248);
or U23715 (N_23715,N_17812,N_17258);
nand U23716 (N_23716,N_17294,N_17727);
xor U23717 (N_23717,N_19107,N_15997);
and U23718 (N_23718,N_15471,N_17894);
and U23719 (N_23719,N_16375,N_19708);
or U23720 (N_23720,N_16582,N_19284);
xnor U23721 (N_23721,N_16998,N_17716);
xor U23722 (N_23722,N_19962,N_18780);
and U23723 (N_23723,N_19190,N_18483);
nor U23724 (N_23724,N_16943,N_17372);
and U23725 (N_23725,N_18408,N_17806);
and U23726 (N_23726,N_18054,N_16255);
nor U23727 (N_23727,N_17986,N_19067);
nand U23728 (N_23728,N_19917,N_17961);
or U23729 (N_23729,N_16086,N_18385);
xnor U23730 (N_23730,N_16301,N_16760);
nand U23731 (N_23731,N_18727,N_17619);
nor U23732 (N_23732,N_16204,N_17311);
nand U23733 (N_23733,N_16185,N_18400);
xor U23734 (N_23734,N_19517,N_18360);
and U23735 (N_23735,N_15045,N_17162);
xor U23736 (N_23736,N_18250,N_16764);
or U23737 (N_23737,N_15706,N_16905);
nor U23738 (N_23738,N_18024,N_16378);
xnor U23739 (N_23739,N_16779,N_18757);
or U23740 (N_23740,N_17023,N_15176);
or U23741 (N_23741,N_19551,N_16306);
xor U23742 (N_23742,N_17546,N_19809);
or U23743 (N_23743,N_17560,N_19590);
nand U23744 (N_23744,N_19140,N_17139);
xor U23745 (N_23745,N_16325,N_18953);
or U23746 (N_23746,N_16093,N_15958);
nand U23747 (N_23747,N_16203,N_17514);
xor U23748 (N_23748,N_19112,N_17459);
xnor U23749 (N_23749,N_16347,N_18191);
nor U23750 (N_23750,N_16740,N_19416);
or U23751 (N_23751,N_18335,N_18237);
nor U23752 (N_23752,N_18744,N_18890);
nor U23753 (N_23753,N_18956,N_17987);
and U23754 (N_23754,N_17303,N_17966);
and U23755 (N_23755,N_17752,N_18701);
nor U23756 (N_23756,N_17642,N_18908);
or U23757 (N_23757,N_15358,N_17967);
and U23758 (N_23758,N_16315,N_17229);
nand U23759 (N_23759,N_17448,N_17568);
nor U23760 (N_23760,N_18055,N_17063);
xnor U23761 (N_23761,N_15712,N_17321);
nor U23762 (N_23762,N_19179,N_18300);
and U23763 (N_23763,N_16360,N_19171);
and U23764 (N_23764,N_15566,N_16584);
xor U23765 (N_23765,N_15734,N_18330);
or U23766 (N_23766,N_18196,N_19575);
or U23767 (N_23767,N_17484,N_15092);
nand U23768 (N_23768,N_15800,N_16369);
nand U23769 (N_23769,N_15543,N_17379);
xnor U23770 (N_23770,N_16014,N_15292);
nor U23771 (N_23771,N_18093,N_15627);
or U23772 (N_23772,N_15357,N_19013);
nor U23773 (N_23773,N_17219,N_19882);
xnor U23774 (N_23774,N_16107,N_15575);
nor U23775 (N_23775,N_18436,N_19110);
nor U23776 (N_23776,N_15296,N_17981);
nor U23777 (N_23777,N_18207,N_19929);
nand U23778 (N_23778,N_18593,N_15583);
xor U23779 (N_23779,N_18524,N_18567);
or U23780 (N_23780,N_16267,N_19202);
and U23781 (N_23781,N_15101,N_18516);
nand U23782 (N_23782,N_15305,N_16324);
xnor U23783 (N_23783,N_18124,N_15911);
nor U23784 (N_23784,N_16824,N_19758);
xor U23785 (N_23785,N_15167,N_18709);
nand U23786 (N_23786,N_18283,N_19530);
xnor U23787 (N_23787,N_17481,N_19180);
or U23788 (N_23788,N_16086,N_18843);
or U23789 (N_23789,N_19309,N_16129);
nand U23790 (N_23790,N_19493,N_15663);
and U23791 (N_23791,N_15893,N_16996);
and U23792 (N_23792,N_15371,N_17940);
or U23793 (N_23793,N_16316,N_16678);
or U23794 (N_23794,N_15671,N_17847);
nand U23795 (N_23795,N_15079,N_18703);
nor U23796 (N_23796,N_18156,N_19062);
xor U23797 (N_23797,N_18561,N_19822);
xnor U23798 (N_23798,N_16907,N_19980);
xnor U23799 (N_23799,N_16356,N_16950);
xor U23800 (N_23800,N_19483,N_17377);
nand U23801 (N_23801,N_19101,N_15513);
xnor U23802 (N_23802,N_15153,N_18187);
xor U23803 (N_23803,N_17981,N_18232);
nor U23804 (N_23804,N_18590,N_15165);
xnor U23805 (N_23805,N_16774,N_16554);
xor U23806 (N_23806,N_16483,N_15782);
and U23807 (N_23807,N_19521,N_15655);
nor U23808 (N_23808,N_19951,N_17224);
nor U23809 (N_23809,N_16936,N_19623);
or U23810 (N_23810,N_15249,N_18978);
and U23811 (N_23811,N_18484,N_17165);
and U23812 (N_23812,N_16997,N_18641);
xnor U23813 (N_23813,N_16891,N_18275);
xor U23814 (N_23814,N_19547,N_15958);
nor U23815 (N_23815,N_18415,N_18655);
or U23816 (N_23816,N_17803,N_18023);
xor U23817 (N_23817,N_16081,N_16682);
nand U23818 (N_23818,N_18976,N_19784);
or U23819 (N_23819,N_19749,N_19500);
xnor U23820 (N_23820,N_15910,N_16615);
and U23821 (N_23821,N_19147,N_18765);
or U23822 (N_23822,N_16439,N_16137);
nand U23823 (N_23823,N_17284,N_18578);
or U23824 (N_23824,N_17785,N_15711);
nor U23825 (N_23825,N_16406,N_15166);
or U23826 (N_23826,N_16680,N_19083);
and U23827 (N_23827,N_15018,N_17266);
xor U23828 (N_23828,N_19793,N_16277);
nand U23829 (N_23829,N_19405,N_19142);
nor U23830 (N_23830,N_17320,N_18318);
nand U23831 (N_23831,N_18850,N_19409);
nand U23832 (N_23832,N_16335,N_19790);
xnor U23833 (N_23833,N_18475,N_18211);
xnor U23834 (N_23834,N_18790,N_19404);
nand U23835 (N_23835,N_18122,N_17154);
and U23836 (N_23836,N_18211,N_16208);
or U23837 (N_23837,N_17703,N_18455);
and U23838 (N_23838,N_15970,N_16355);
or U23839 (N_23839,N_15125,N_19513);
or U23840 (N_23840,N_19308,N_18771);
nand U23841 (N_23841,N_17735,N_16702);
or U23842 (N_23842,N_16538,N_17653);
and U23843 (N_23843,N_15964,N_17728);
nor U23844 (N_23844,N_17280,N_18036);
and U23845 (N_23845,N_18981,N_19008);
nor U23846 (N_23846,N_16886,N_17252);
nand U23847 (N_23847,N_19029,N_19172);
and U23848 (N_23848,N_16073,N_18429);
and U23849 (N_23849,N_19411,N_17581);
and U23850 (N_23850,N_19981,N_19674);
or U23851 (N_23851,N_15919,N_17700);
and U23852 (N_23852,N_16923,N_17588);
xor U23853 (N_23853,N_17927,N_16775);
and U23854 (N_23854,N_17006,N_16817);
xnor U23855 (N_23855,N_15458,N_16273);
or U23856 (N_23856,N_16819,N_16577);
or U23857 (N_23857,N_19239,N_15756);
xnor U23858 (N_23858,N_18874,N_15259);
nor U23859 (N_23859,N_18134,N_16372);
xor U23860 (N_23860,N_15653,N_16285);
nand U23861 (N_23861,N_16696,N_15515);
and U23862 (N_23862,N_18961,N_17878);
xnor U23863 (N_23863,N_15416,N_17766);
nor U23864 (N_23864,N_15811,N_19689);
xor U23865 (N_23865,N_19411,N_19031);
and U23866 (N_23866,N_18616,N_15679);
and U23867 (N_23867,N_18914,N_15666);
nor U23868 (N_23868,N_16551,N_18944);
nor U23869 (N_23869,N_18019,N_17777);
xor U23870 (N_23870,N_15048,N_18237);
xnor U23871 (N_23871,N_15923,N_17891);
nand U23872 (N_23872,N_18818,N_17293);
nand U23873 (N_23873,N_17644,N_17079);
xor U23874 (N_23874,N_19637,N_16730);
nand U23875 (N_23875,N_18382,N_17820);
nand U23876 (N_23876,N_16051,N_15633);
nand U23877 (N_23877,N_16715,N_16071);
nand U23878 (N_23878,N_16119,N_18840);
nor U23879 (N_23879,N_16706,N_16343);
xnor U23880 (N_23880,N_15320,N_19691);
and U23881 (N_23881,N_19107,N_17323);
xnor U23882 (N_23882,N_17489,N_17334);
nand U23883 (N_23883,N_18341,N_17199);
xor U23884 (N_23884,N_15222,N_17932);
or U23885 (N_23885,N_19385,N_15957);
and U23886 (N_23886,N_19834,N_17976);
and U23887 (N_23887,N_17358,N_16225);
or U23888 (N_23888,N_19671,N_16507);
and U23889 (N_23889,N_18474,N_18356);
and U23890 (N_23890,N_18366,N_17785);
nor U23891 (N_23891,N_16862,N_17596);
or U23892 (N_23892,N_15675,N_17025);
and U23893 (N_23893,N_16762,N_16531);
and U23894 (N_23894,N_15816,N_16328);
or U23895 (N_23895,N_17396,N_16830);
nor U23896 (N_23896,N_18205,N_16439);
nor U23897 (N_23897,N_17862,N_19848);
nor U23898 (N_23898,N_18863,N_15429);
nor U23899 (N_23899,N_16763,N_16421);
or U23900 (N_23900,N_17346,N_19079);
xnor U23901 (N_23901,N_17679,N_19394);
nand U23902 (N_23902,N_17457,N_18077);
nand U23903 (N_23903,N_17604,N_18978);
nand U23904 (N_23904,N_15051,N_18036);
nor U23905 (N_23905,N_19428,N_16908);
or U23906 (N_23906,N_16224,N_15407);
nand U23907 (N_23907,N_15209,N_15394);
nand U23908 (N_23908,N_18830,N_18993);
or U23909 (N_23909,N_17095,N_16766);
and U23910 (N_23910,N_16992,N_15917);
nand U23911 (N_23911,N_17264,N_16871);
nor U23912 (N_23912,N_17817,N_19517);
xor U23913 (N_23913,N_16681,N_16889);
or U23914 (N_23914,N_17924,N_15728);
and U23915 (N_23915,N_18915,N_18339);
xnor U23916 (N_23916,N_16730,N_15122);
and U23917 (N_23917,N_15587,N_16351);
or U23918 (N_23918,N_18010,N_19825);
nor U23919 (N_23919,N_17241,N_15929);
and U23920 (N_23920,N_17687,N_17354);
and U23921 (N_23921,N_19609,N_18062);
nand U23922 (N_23922,N_15974,N_17991);
nor U23923 (N_23923,N_18689,N_17766);
and U23924 (N_23924,N_19361,N_15832);
nor U23925 (N_23925,N_19952,N_17682);
and U23926 (N_23926,N_18072,N_15468);
nor U23927 (N_23927,N_17290,N_16557);
and U23928 (N_23928,N_18918,N_19152);
nand U23929 (N_23929,N_18364,N_19226);
nand U23930 (N_23930,N_18846,N_18405);
and U23931 (N_23931,N_16792,N_15260);
nand U23932 (N_23932,N_18293,N_18349);
xor U23933 (N_23933,N_15535,N_15615);
and U23934 (N_23934,N_17618,N_15029);
nor U23935 (N_23935,N_18705,N_16264);
and U23936 (N_23936,N_15293,N_16576);
and U23937 (N_23937,N_18273,N_17289);
nor U23938 (N_23938,N_19543,N_19731);
and U23939 (N_23939,N_18225,N_18938);
and U23940 (N_23940,N_17421,N_16646);
and U23941 (N_23941,N_17229,N_18181);
nor U23942 (N_23942,N_15280,N_19464);
nand U23943 (N_23943,N_18127,N_15952);
or U23944 (N_23944,N_18003,N_19740);
nand U23945 (N_23945,N_15760,N_16602);
and U23946 (N_23946,N_16306,N_18298);
nand U23947 (N_23947,N_17013,N_18057);
or U23948 (N_23948,N_19949,N_19573);
xnor U23949 (N_23949,N_16482,N_15785);
or U23950 (N_23950,N_18940,N_17140);
xnor U23951 (N_23951,N_18708,N_16487);
nor U23952 (N_23952,N_17232,N_15687);
xor U23953 (N_23953,N_15297,N_16446);
nor U23954 (N_23954,N_15662,N_15035);
or U23955 (N_23955,N_16572,N_17448);
and U23956 (N_23956,N_19627,N_17129);
nor U23957 (N_23957,N_18270,N_18588);
and U23958 (N_23958,N_17137,N_17273);
or U23959 (N_23959,N_18280,N_18921);
or U23960 (N_23960,N_16119,N_18619);
xor U23961 (N_23961,N_16225,N_19969);
nor U23962 (N_23962,N_19579,N_19304);
nor U23963 (N_23963,N_17560,N_17718);
xnor U23964 (N_23964,N_17942,N_16769);
or U23965 (N_23965,N_17826,N_18188);
or U23966 (N_23966,N_19982,N_15971);
xnor U23967 (N_23967,N_18029,N_18861);
xnor U23968 (N_23968,N_16812,N_15045);
xnor U23969 (N_23969,N_16759,N_19275);
and U23970 (N_23970,N_19116,N_18176);
xor U23971 (N_23971,N_19841,N_19142);
nor U23972 (N_23972,N_17447,N_16058);
and U23973 (N_23973,N_16073,N_19888);
nor U23974 (N_23974,N_17926,N_17554);
and U23975 (N_23975,N_18550,N_17237);
xor U23976 (N_23976,N_17828,N_18865);
nor U23977 (N_23977,N_19194,N_17096);
and U23978 (N_23978,N_18762,N_17076);
nor U23979 (N_23979,N_16144,N_15925);
or U23980 (N_23980,N_16556,N_15343);
nor U23981 (N_23981,N_17095,N_15190);
nor U23982 (N_23982,N_15888,N_16619);
or U23983 (N_23983,N_17221,N_17634);
and U23984 (N_23984,N_17692,N_17357);
xnor U23985 (N_23985,N_18900,N_15996);
and U23986 (N_23986,N_19954,N_18670);
and U23987 (N_23987,N_16711,N_17906);
and U23988 (N_23988,N_18962,N_17834);
or U23989 (N_23989,N_17337,N_16325);
nand U23990 (N_23990,N_19839,N_16531);
xnor U23991 (N_23991,N_15546,N_16152);
and U23992 (N_23992,N_19616,N_18620);
nand U23993 (N_23993,N_18020,N_17148);
nand U23994 (N_23994,N_19354,N_17397);
xor U23995 (N_23995,N_16977,N_17898);
and U23996 (N_23996,N_17234,N_18869);
xor U23997 (N_23997,N_16422,N_16474);
or U23998 (N_23998,N_16125,N_17116);
nor U23999 (N_23999,N_18294,N_19339);
and U24000 (N_24000,N_17064,N_17736);
nand U24001 (N_24001,N_16454,N_18481);
xnor U24002 (N_24002,N_18522,N_15472);
or U24003 (N_24003,N_19503,N_17080);
and U24004 (N_24004,N_19816,N_15583);
nor U24005 (N_24005,N_19177,N_16471);
nand U24006 (N_24006,N_15821,N_15421);
nand U24007 (N_24007,N_18161,N_17888);
xor U24008 (N_24008,N_15910,N_17050);
and U24009 (N_24009,N_16381,N_19156);
xnor U24010 (N_24010,N_16729,N_17004);
or U24011 (N_24011,N_16366,N_18062);
or U24012 (N_24012,N_15148,N_19107);
and U24013 (N_24013,N_17559,N_19575);
or U24014 (N_24014,N_15361,N_16929);
or U24015 (N_24015,N_18165,N_17689);
nor U24016 (N_24016,N_15665,N_16772);
or U24017 (N_24017,N_16524,N_17143);
nand U24018 (N_24018,N_17902,N_19995);
or U24019 (N_24019,N_15079,N_15400);
and U24020 (N_24020,N_17960,N_16496);
xnor U24021 (N_24021,N_19978,N_16189);
and U24022 (N_24022,N_19170,N_17398);
xor U24023 (N_24023,N_17976,N_19229);
nand U24024 (N_24024,N_17608,N_19070);
and U24025 (N_24025,N_19035,N_18178);
and U24026 (N_24026,N_15371,N_18736);
xnor U24027 (N_24027,N_17642,N_15827);
nor U24028 (N_24028,N_17543,N_17077);
or U24029 (N_24029,N_15740,N_19500);
and U24030 (N_24030,N_15810,N_15539);
or U24031 (N_24031,N_18704,N_18040);
xor U24032 (N_24032,N_18235,N_19942);
nor U24033 (N_24033,N_15650,N_15638);
nor U24034 (N_24034,N_17870,N_15472);
nand U24035 (N_24035,N_15706,N_19920);
nor U24036 (N_24036,N_16890,N_18839);
xnor U24037 (N_24037,N_15682,N_19779);
nor U24038 (N_24038,N_17799,N_17434);
nand U24039 (N_24039,N_15774,N_16998);
xor U24040 (N_24040,N_15390,N_19616);
nor U24041 (N_24041,N_18659,N_16513);
xnor U24042 (N_24042,N_18647,N_15247);
and U24043 (N_24043,N_18771,N_19579);
xnor U24044 (N_24044,N_19947,N_16594);
or U24045 (N_24045,N_18593,N_18343);
nand U24046 (N_24046,N_15874,N_16235);
or U24047 (N_24047,N_16481,N_18085);
nor U24048 (N_24048,N_19279,N_17557);
or U24049 (N_24049,N_15729,N_17686);
nor U24050 (N_24050,N_15670,N_17186);
nor U24051 (N_24051,N_19173,N_16772);
nor U24052 (N_24052,N_16979,N_16212);
nand U24053 (N_24053,N_16721,N_19606);
and U24054 (N_24054,N_19499,N_19599);
nand U24055 (N_24055,N_18304,N_16389);
xnor U24056 (N_24056,N_18465,N_18002);
nand U24057 (N_24057,N_17871,N_16272);
xnor U24058 (N_24058,N_15137,N_19180);
nor U24059 (N_24059,N_17147,N_16405);
and U24060 (N_24060,N_18137,N_18158);
nand U24061 (N_24061,N_18782,N_15020);
xor U24062 (N_24062,N_17286,N_18094);
nor U24063 (N_24063,N_15280,N_19384);
xor U24064 (N_24064,N_18306,N_16320);
nand U24065 (N_24065,N_16379,N_19714);
xor U24066 (N_24066,N_17172,N_18255);
nor U24067 (N_24067,N_19044,N_15661);
nand U24068 (N_24068,N_15059,N_18520);
nand U24069 (N_24069,N_17143,N_19367);
xnor U24070 (N_24070,N_18608,N_18103);
and U24071 (N_24071,N_16925,N_18819);
nand U24072 (N_24072,N_15958,N_19948);
xor U24073 (N_24073,N_16442,N_16683);
nor U24074 (N_24074,N_18964,N_15083);
and U24075 (N_24075,N_15946,N_16685);
nand U24076 (N_24076,N_17032,N_17214);
nor U24077 (N_24077,N_16090,N_17268);
xor U24078 (N_24078,N_17659,N_19873);
nand U24079 (N_24079,N_15847,N_17454);
or U24080 (N_24080,N_18208,N_16112);
nor U24081 (N_24081,N_17636,N_17066);
nand U24082 (N_24082,N_17237,N_18134);
xor U24083 (N_24083,N_15814,N_19378);
nor U24084 (N_24084,N_17435,N_18515);
nor U24085 (N_24085,N_19533,N_17745);
xor U24086 (N_24086,N_17309,N_16196);
and U24087 (N_24087,N_15245,N_18092);
or U24088 (N_24088,N_17453,N_16213);
nand U24089 (N_24089,N_15420,N_16620);
nor U24090 (N_24090,N_16762,N_15430);
or U24091 (N_24091,N_15288,N_16660);
nor U24092 (N_24092,N_15550,N_16863);
xor U24093 (N_24093,N_16681,N_18200);
or U24094 (N_24094,N_15451,N_16269);
xor U24095 (N_24095,N_16049,N_15633);
or U24096 (N_24096,N_17068,N_18273);
xnor U24097 (N_24097,N_16115,N_18818);
or U24098 (N_24098,N_15799,N_16134);
xnor U24099 (N_24099,N_17213,N_19479);
xnor U24100 (N_24100,N_17752,N_15296);
xor U24101 (N_24101,N_17704,N_15626);
nand U24102 (N_24102,N_18783,N_17778);
or U24103 (N_24103,N_15158,N_18157);
nand U24104 (N_24104,N_18438,N_17005);
xor U24105 (N_24105,N_19996,N_17119);
nor U24106 (N_24106,N_18161,N_17821);
nand U24107 (N_24107,N_16022,N_15629);
and U24108 (N_24108,N_17420,N_16334);
xor U24109 (N_24109,N_17039,N_15206);
nand U24110 (N_24110,N_15363,N_17867);
xnor U24111 (N_24111,N_16118,N_18399);
and U24112 (N_24112,N_15409,N_17002);
nor U24113 (N_24113,N_15843,N_18232);
nor U24114 (N_24114,N_15537,N_15316);
or U24115 (N_24115,N_16749,N_15805);
nor U24116 (N_24116,N_17330,N_19152);
and U24117 (N_24117,N_18160,N_18232);
or U24118 (N_24118,N_18992,N_18129);
xnor U24119 (N_24119,N_19054,N_19810);
nor U24120 (N_24120,N_18841,N_16835);
or U24121 (N_24121,N_19477,N_15870);
and U24122 (N_24122,N_18509,N_18437);
nor U24123 (N_24123,N_18978,N_18958);
xnor U24124 (N_24124,N_17195,N_19552);
and U24125 (N_24125,N_18276,N_17803);
and U24126 (N_24126,N_17111,N_18885);
nand U24127 (N_24127,N_15047,N_15783);
xor U24128 (N_24128,N_17646,N_17629);
xnor U24129 (N_24129,N_15274,N_16454);
or U24130 (N_24130,N_16645,N_19666);
or U24131 (N_24131,N_18104,N_16433);
nor U24132 (N_24132,N_15159,N_16178);
and U24133 (N_24133,N_16924,N_16979);
xor U24134 (N_24134,N_18799,N_17694);
xor U24135 (N_24135,N_16244,N_16299);
or U24136 (N_24136,N_17783,N_16454);
nand U24137 (N_24137,N_19223,N_19136);
or U24138 (N_24138,N_18062,N_17238);
nor U24139 (N_24139,N_17747,N_19163);
nor U24140 (N_24140,N_18123,N_15577);
and U24141 (N_24141,N_19653,N_16619);
xnor U24142 (N_24142,N_19099,N_17794);
xor U24143 (N_24143,N_17939,N_17032);
nor U24144 (N_24144,N_19768,N_17184);
nand U24145 (N_24145,N_16931,N_15304);
and U24146 (N_24146,N_16387,N_15875);
nor U24147 (N_24147,N_19919,N_19244);
or U24148 (N_24148,N_18724,N_17001);
nor U24149 (N_24149,N_19443,N_17058);
and U24150 (N_24150,N_16954,N_19589);
xor U24151 (N_24151,N_18449,N_16804);
nand U24152 (N_24152,N_19792,N_15119);
xor U24153 (N_24153,N_15559,N_18565);
nand U24154 (N_24154,N_19742,N_18513);
nand U24155 (N_24155,N_15220,N_18970);
nor U24156 (N_24156,N_16552,N_18774);
xnor U24157 (N_24157,N_19486,N_16536);
nor U24158 (N_24158,N_16668,N_15998);
nor U24159 (N_24159,N_16028,N_15627);
and U24160 (N_24160,N_17016,N_16697);
nor U24161 (N_24161,N_19339,N_19532);
or U24162 (N_24162,N_18655,N_19559);
or U24163 (N_24163,N_16085,N_15888);
xnor U24164 (N_24164,N_15302,N_16981);
nand U24165 (N_24165,N_19011,N_17442);
or U24166 (N_24166,N_15154,N_18419);
and U24167 (N_24167,N_19093,N_15756);
or U24168 (N_24168,N_16558,N_19557);
and U24169 (N_24169,N_16251,N_19822);
xnor U24170 (N_24170,N_15083,N_18459);
nor U24171 (N_24171,N_15098,N_18922);
nor U24172 (N_24172,N_17215,N_16845);
nor U24173 (N_24173,N_15407,N_18823);
and U24174 (N_24174,N_17015,N_17203);
and U24175 (N_24175,N_17425,N_17530);
nor U24176 (N_24176,N_16963,N_16330);
nand U24177 (N_24177,N_19204,N_17371);
xor U24178 (N_24178,N_18654,N_16315);
xor U24179 (N_24179,N_15430,N_19604);
xor U24180 (N_24180,N_17975,N_15376);
or U24181 (N_24181,N_18009,N_17740);
xor U24182 (N_24182,N_16201,N_15394);
xnor U24183 (N_24183,N_15935,N_18682);
nand U24184 (N_24184,N_18172,N_19136);
nand U24185 (N_24185,N_17485,N_19038);
or U24186 (N_24186,N_18675,N_18249);
or U24187 (N_24187,N_17007,N_18734);
nor U24188 (N_24188,N_17529,N_18514);
xnor U24189 (N_24189,N_15677,N_16886);
nand U24190 (N_24190,N_19179,N_15867);
and U24191 (N_24191,N_19021,N_19617);
nor U24192 (N_24192,N_15514,N_16803);
nand U24193 (N_24193,N_19548,N_17215);
xnor U24194 (N_24194,N_19602,N_17951);
or U24195 (N_24195,N_18096,N_18773);
and U24196 (N_24196,N_18630,N_16558);
xor U24197 (N_24197,N_17811,N_15896);
xnor U24198 (N_24198,N_17723,N_19499);
and U24199 (N_24199,N_15160,N_17096);
nor U24200 (N_24200,N_15654,N_19496);
nand U24201 (N_24201,N_15753,N_15469);
or U24202 (N_24202,N_19409,N_19784);
nor U24203 (N_24203,N_16103,N_18594);
nor U24204 (N_24204,N_15408,N_18316);
and U24205 (N_24205,N_15485,N_19456);
xnor U24206 (N_24206,N_15508,N_15349);
nand U24207 (N_24207,N_16876,N_19254);
and U24208 (N_24208,N_16585,N_18388);
xnor U24209 (N_24209,N_15529,N_18100);
and U24210 (N_24210,N_17223,N_19452);
nor U24211 (N_24211,N_17440,N_15107);
and U24212 (N_24212,N_19019,N_16087);
nor U24213 (N_24213,N_16507,N_19183);
xor U24214 (N_24214,N_15760,N_16683);
and U24215 (N_24215,N_16317,N_19241);
nand U24216 (N_24216,N_15021,N_16520);
nor U24217 (N_24217,N_19006,N_19916);
or U24218 (N_24218,N_19271,N_17878);
nand U24219 (N_24219,N_15951,N_17472);
or U24220 (N_24220,N_19026,N_16218);
and U24221 (N_24221,N_18284,N_15630);
nor U24222 (N_24222,N_15840,N_16543);
and U24223 (N_24223,N_19632,N_17868);
or U24224 (N_24224,N_17461,N_19705);
nor U24225 (N_24225,N_18833,N_16217);
xnor U24226 (N_24226,N_15140,N_19355);
or U24227 (N_24227,N_18496,N_16273);
and U24228 (N_24228,N_18901,N_19429);
and U24229 (N_24229,N_18394,N_15292);
nand U24230 (N_24230,N_16796,N_16971);
nor U24231 (N_24231,N_17249,N_18695);
and U24232 (N_24232,N_16797,N_19053);
and U24233 (N_24233,N_18645,N_17207);
or U24234 (N_24234,N_16079,N_17685);
xor U24235 (N_24235,N_18330,N_15893);
or U24236 (N_24236,N_16774,N_16732);
and U24237 (N_24237,N_17790,N_17969);
and U24238 (N_24238,N_19372,N_17095);
xnor U24239 (N_24239,N_19927,N_17976);
xnor U24240 (N_24240,N_16834,N_18627);
nor U24241 (N_24241,N_15476,N_15752);
and U24242 (N_24242,N_17655,N_19053);
nor U24243 (N_24243,N_15920,N_19978);
or U24244 (N_24244,N_17042,N_17963);
or U24245 (N_24245,N_15303,N_16430);
or U24246 (N_24246,N_18477,N_19126);
xor U24247 (N_24247,N_15094,N_17780);
or U24248 (N_24248,N_18544,N_16579);
nor U24249 (N_24249,N_15935,N_19529);
or U24250 (N_24250,N_16006,N_17373);
and U24251 (N_24251,N_16793,N_16328);
nand U24252 (N_24252,N_19070,N_17043);
or U24253 (N_24253,N_16090,N_18329);
nor U24254 (N_24254,N_19038,N_17247);
and U24255 (N_24255,N_16766,N_19493);
xnor U24256 (N_24256,N_17790,N_17798);
xor U24257 (N_24257,N_18914,N_18333);
nand U24258 (N_24258,N_16350,N_17513);
nand U24259 (N_24259,N_19604,N_17868);
nor U24260 (N_24260,N_17235,N_16005);
nor U24261 (N_24261,N_19769,N_18172);
and U24262 (N_24262,N_16710,N_15397);
xnor U24263 (N_24263,N_17186,N_15311);
nand U24264 (N_24264,N_18932,N_19839);
nand U24265 (N_24265,N_15334,N_15993);
or U24266 (N_24266,N_19470,N_16095);
and U24267 (N_24267,N_16179,N_16824);
xor U24268 (N_24268,N_18284,N_16702);
nor U24269 (N_24269,N_17962,N_17042);
nand U24270 (N_24270,N_18277,N_17457);
nor U24271 (N_24271,N_15044,N_18492);
nand U24272 (N_24272,N_15665,N_18327);
xor U24273 (N_24273,N_18706,N_16658);
nand U24274 (N_24274,N_17915,N_18838);
and U24275 (N_24275,N_15287,N_19198);
xnor U24276 (N_24276,N_15473,N_19593);
or U24277 (N_24277,N_17997,N_19201);
nor U24278 (N_24278,N_19131,N_16066);
xor U24279 (N_24279,N_16468,N_19212);
nand U24280 (N_24280,N_19035,N_19698);
nand U24281 (N_24281,N_19766,N_16717);
xnor U24282 (N_24282,N_16712,N_17237);
nand U24283 (N_24283,N_16431,N_15849);
xor U24284 (N_24284,N_17952,N_18741);
and U24285 (N_24285,N_17355,N_15198);
and U24286 (N_24286,N_17301,N_18120);
nand U24287 (N_24287,N_18351,N_17170);
nand U24288 (N_24288,N_16350,N_16425);
and U24289 (N_24289,N_16848,N_16136);
xnor U24290 (N_24290,N_19283,N_16587);
or U24291 (N_24291,N_16475,N_15099);
nor U24292 (N_24292,N_16701,N_19874);
nor U24293 (N_24293,N_19692,N_16726);
xor U24294 (N_24294,N_19041,N_19010);
nor U24295 (N_24295,N_16072,N_19998);
and U24296 (N_24296,N_16211,N_15115);
xnor U24297 (N_24297,N_16464,N_17469);
nand U24298 (N_24298,N_18567,N_18821);
or U24299 (N_24299,N_19154,N_17335);
nor U24300 (N_24300,N_19879,N_18820);
nand U24301 (N_24301,N_18767,N_15379);
nand U24302 (N_24302,N_15850,N_16457);
nand U24303 (N_24303,N_18973,N_18773);
xor U24304 (N_24304,N_15471,N_17565);
and U24305 (N_24305,N_19316,N_18849);
and U24306 (N_24306,N_18125,N_15897);
nand U24307 (N_24307,N_18771,N_15772);
and U24308 (N_24308,N_17274,N_19419);
xnor U24309 (N_24309,N_17317,N_16654);
xnor U24310 (N_24310,N_19548,N_19699);
nand U24311 (N_24311,N_17587,N_19080);
xnor U24312 (N_24312,N_18163,N_15763);
or U24313 (N_24313,N_15366,N_17541);
nand U24314 (N_24314,N_16725,N_17248);
or U24315 (N_24315,N_19472,N_18587);
xnor U24316 (N_24316,N_17161,N_16511);
nand U24317 (N_24317,N_16123,N_19145);
nor U24318 (N_24318,N_18951,N_17613);
xor U24319 (N_24319,N_15980,N_15988);
nand U24320 (N_24320,N_15164,N_18411);
nor U24321 (N_24321,N_15406,N_19495);
or U24322 (N_24322,N_18699,N_17595);
and U24323 (N_24323,N_16699,N_16696);
nand U24324 (N_24324,N_16215,N_19775);
nor U24325 (N_24325,N_16111,N_18060);
nand U24326 (N_24326,N_19221,N_18612);
and U24327 (N_24327,N_17191,N_18290);
xor U24328 (N_24328,N_19804,N_17526);
nor U24329 (N_24329,N_18342,N_15518);
and U24330 (N_24330,N_19841,N_15982);
xnor U24331 (N_24331,N_15628,N_16339);
and U24332 (N_24332,N_18449,N_18768);
nor U24333 (N_24333,N_16664,N_17714);
or U24334 (N_24334,N_15851,N_16015);
and U24335 (N_24335,N_16253,N_15331);
and U24336 (N_24336,N_18712,N_18861);
and U24337 (N_24337,N_17955,N_17616);
or U24338 (N_24338,N_15535,N_15560);
or U24339 (N_24339,N_16678,N_15893);
xnor U24340 (N_24340,N_17652,N_18532);
and U24341 (N_24341,N_16843,N_17203);
nand U24342 (N_24342,N_16702,N_15825);
nor U24343 (N_24343,N_18280,N_15090);
nand U24344 (N_24344,N_16230,N_15548);
and U24345 (N_24345,N_17649,N_15504);
and U24346 (N_24346,N_18043,N_15703);
nand U24347 (N_24347,N_15208,N_16569);
nand U24348 (N_24348,N_16739,N_19846);
nor U24349 (N_24349,N_18217,N_18938);
and U24350 (N_24350,N_17870,N_17903);
nand U24351 (N_24351,N_15766,N_18716);
nand U24352 (N_24352,N_18650,N_18370);
nand U24353 (N_24353,N_15483,N_19328);
nand U24354 (N_24354,N_16766,N_16860);
nand U24355 (N_24355,N_18853,N_17386);
and U24356 (N_24356,N_17654,N_16834);
and U24357 (N_24357,N_18865,N_17296);
nor U24358 (N_24358,N_17129,N_19533);
or U24359 (N_24359,N_15217,N_17374);
nor U24360 (N_24360,N_18457,N_15750);
xor U24361 (N_24361,N_18310,N_19985);
nand U24362 (N_24362,N_15091,N_15453);
nor U24363 (N_24363,N_15607,N_17293);
or U24364 (N_24364,N_15548,N_18735);
nand U24365 (N_24365,N_17414,N_15985);
xnor U24366 (N_24366,N_18152,N_19962);
xor U24367 (N_24367,N_15947,N_17961);
nor U24368 (N_24368,N_18418,N_15161);
nand U24369 (N_24369,N_16252,N_18996);
or U24370 (N_24370,N_16017,N_16578);
nand U24371 (N_24371,N_19883,N_16424);
nor U24372 (N_24372,N_15304,N_19466);
xnor U24373 (N_24373,N_17219,N_19371);
nand U24374 (N_24374,N_18830,N_19883);
or U24375 (N_24375,N_17345,N_19402);
or U24376 (N_24376,N_18834,N_17033);
or U24377 (N_24377,N_18103,N_16140);
nand U24378 (N_24378,N_16359,N_18270);
nand U24379 (N_24379,N_19734,N_17017);
or U24380 (N_24380,N_17498,N_15122);
nand U24381 (N_24381,N_19333,N_17330);
xor U24382 (N_24382,N_17792,N_16385);
xor U24383 (N_24383,N_15193,N_15057);
xor U24384 (N_24384,N_17744,N_15418);
xnor U24385 (N_24385,N_17164,N_19437);
and U24386 (N_24386,N_16129,N_16028);
xor U24387 (N_24387,N_19975,N_15566);
nand U24388 (N_24388,N_17717,N_18655);
nand U24389 (N_24389,N_18165,N_15094);
nand U24390 (N_24390,N_18893,N_15397);
or U24391 (N_24391,N_18468,N_15877);
and U24392 (N_24392,N_17500,N_19767);
and U24393 (N_24393,N_18286,N_18127);
nor U24394 (N_24394,N_19740,N_18066);
nor U24395 (N_24395,N_16332,N_19694);
or U24396 (N_24396,N_18979,N_17265);
nand U24397 (N_24397,N_15111,N_15013);
nor U24398 (N_24398,N_16298,N_18914);
nor U24399 (N_24399,N_18839,N_19333);
nand U24400 (N_24400,N_15767,N_18058);
or U24401 (N_24401,N_17597,N_19315);
and U24402 (N_24402,N_18483,N_16603);
and U24403 (N_24403,N_19009,N_16498);
and U24404 (N_24404,N_18983,N_15143);
nand U24405 (N_24405,N_19555,N_19772);
nand U24406 (N_24406,N_15129,N_15916);
xor U24407 (N_24407,N_17723,N_16649);
xor U24408 (N_24408,N_19929,N_16021);
xnor U24409 (N_24409,N_15405,N_16683);
xor U24410 (N_24410,N_16569,N_16678);
and U24411 (N_24411,N_18019,N_15226);
nor U24412 (N_24412,N_17985,N_16002);
and U24413 (N_24413,N_15158,N_18624);
nand U24414 (N_24414,N_15981,N_16203);
or U24415 (N_24415,N_17443,N_18875);
nand U24416 (N_24416,N_15437,N_17798);
and U24417 (N_24417,N_16202,N_19393);
or U24418 (N_24418,N_17626,N_18498);
nor U24419 (N_24419,N_19751,N_17998);
or U24420 (N_24420,N_16869,N_19097);
nor U24421 (N_24421,N_19905,N_16935);
xor U24422 (N_24422,N_17476,N_19258);
and U24423 (N_24423,N_16289,N_19624);
or U24424 (N_24424,N_15826,N_19257);
nand U24425 (N_24425,N_15112,N_18461);
nand U24426 (N_24426,N_16442,N_15411);
or U24427 (N_24427,N_16037,N_16708);
xor U24428 (N_24428,N_19059,N_16124);
nand U24429 (N_24429,N_17214,N_15956);
and U24430 (N_24430,N_18438,N_17584);
and U24431 (N_24431,N_17251,N_17614);
nand U24432 (N_24432,N_17836,N_16907);
and U24433 (N_24433,N_17729,N_16187);
nand U24434 (N_24434,N_19385,N_16177);
and U24435 (N_24435,N_19724,N_16705);
xor U24436 (N_24436,N_15688,N_16988);
nor U24437 (N_24437,N_17385,N_17938);
or U24438 (N_24438,N_18427,N_16736);
xor U24439 (N_24439,N_15050,N_16781);
nand U24440 (N_24440,N_15440,N_16905);
xnor U24441 (N_24441,N_16823,N_16771);
or U24442 (N_24442,N_17283,N_15147);
nor U24443 (N_24443,N_15693,N_16028);
xnor U24444 (N_24444,N_19428,N_19816);
or U24445 (N_24445,N_16390,N_19506);
nand U24446 (N_24446,N_18754,N_16683);
xnor U24447 (N_24447,N_15852,N_19023);
xnor U24448 (N_24448,N_18100,N_15509);
nor U24449 (N_24449,N_16296,N_15425);
or U24450 (N_24450,N_16144,N_17977);
or U24451 (N_24451,N_19282,N_15290);
nand U24452 (N_24452,N_17190,N_16411);
and U24453 (N_24453,N_15487,N_17942);
and U24454 (N_24454,N_18549,N_17652);
xnor U24455 (N_24455,N_17753,N_18898);
xnor U24456 (N_24456,N_15126,N_16585);
or U24457 (N_24457,N_18460,N_15444);
or U24458 (N_24458,N_16679,N_17294);
nand U24459 (N_24459,N_16239,N_17051);
and U24460 (N_24460,N_16155,N_18291);
and U24461 (N_24461,N_19645,N_16151);
nand U24462 (N_24462,N_18946,N_17549);
nor U24463 (N_24463,N_19629,N_18683);
xnor U24464 (N_24464,N_15459,N_17155);
nand U24465 (N_24465,N_16917,N_19756);
nand U24466 (N_24466,N_17740,N_18349);
and U24467 (N_24467,N_18924,N_17476);
nand U24468 (N_24468,N_17286,N_17597);
xor U24469 (N_24469,N_17522,N_15767);
and U24470 (N_24470,N_15844,N_15001);
and U24471 (N_24471,N_17973,N_18139);
or U24472 (N_24472,N_16540,N_17061);
nor U24473 (N_24473,N_19326,N_16920);
nor U24474 (N_24474,N_16470,N_15107);
nand U24475 (N_24475,N_18273,N_18149);
nor U24476 (N_24476,N_15573,N_16875);
and U24477 (N_24477,N_19463,N_19054);
nand U24478 (N_24478,N_18301,N_16216);
xor U24479 (N_24479,N_17869,N_16299);
nor U24480 (N_24480,N_18512,N_15260);
nand U24481 (N_24481,N_16718,N_17594);
xor U24482 (N_24482,N_15612,N_18157);
xnor U24483 (N_24483,N_15157,N_17130);
or U24484 (N_24484,N_19875,N_16953);
nand U24485 (N_24485,N_18359,N_18839);
xnor U24486 (N_24486,N_15195,N_16118);
or U24487 (N_24487,N_15241,N_16402);
and U24488 (N_24488,N_15596,N_16165);
and U24489 (N_24489,N_15987,N_19822);
nand U24490 (N_24490,N_19599,N_16419);
or U24491 (N_24491,N_16537,N_16408);
and U24492 (N_24492,N_17496,N_18250);
or U24493 (N_24493,N_19667,N_17131);
xor U24494 (N_24494,N_16076,N_15982);
and U24495 (N_24495,N_18684,N_15501);
and U24496 (N_24496,N_15990,N_17888);
and U24497 (N_24497,N_18008,N_17310);
xnor U24498 (N_24498,N_17946,N_17805);
nor U24499 (N_24499,N_15248,N_15419);
xor U24500 (N_24500,N_15237,N_15881);
or U24501 (N_24501,N_19831,N_15383);
nor U24502 (N_24502,N_18061,N_15471);
and U24503 (N_24503,N_17992,N_17366);
or U24504 (N_24504,N_18905,N_18031);
and U24505 (N_24505,N_18720,N_19279);
xnor U24506 (N_24506,N_17584,N_16201);
nand U24507 (N_24507,N_19760,N_19654);
nand U24508 (N_24508,N_15576,N_17973);
xnor U24509 (N_24509,N_18814,N_16111);
and U24510 (N_24510,N_16228,N_17183);
or U24511 (N_24511,N_19262,N_16878);
xor U24512 (N_24512,N_17766,N_18637);
xor U24513 (N_24513,N_18363,N_18483);
nor U24514 (N_24514,N_17768,N_16539);
or U24515 (N_24515,N_16078,N_18144);
xnor U24516 (N_24516,N_18657,N_16818);
xnor U24517 (N_24517,N_17971,N_19429);
xor U24518 (N_24518,N_15803,N_17483);
nand U24519 (N_24519,N_16056,N_15063);
or U24520 (N_24520,N_18991,N_15929);
and U24521 (N_24521,N_17803,N_16911);
nor U24522 (N_24522,N_17778,N_17622);
nand U24523 (N_24523,N_18782,N_17275);
or U24524 (N_24524,N_16983,N_15632);
nor U24525 (N_24525,N_17740,N_15239);
xor U24526 (N_24526,N_19818,N_19089);
or U24527 (N_24527,N_16048,N_16726);
and U24528 (N_24528,N_19681,N_19255);
nand U24529 (N_24529,N_19582,N_15147);
nand U24530 (N_24530,N_15847,N_16245);
nor U24531 (N_24531,N_18548,N_16248);
nor U24532 (N_24532,N_16168,N_19718);
and U24533 (N_24533,N_19174,N_19910);
and U24534 (N_24534,N_19434,N_19378);
xor U24535 (N_24535,N_19835,N_15944);
nand U24536 (N_24536,N_15119,N_17265);
or U24537 (N_24537,N_15624,N_15777);
nor U24538 (N_24538,N_15363,N_17058);
and U24539 (N_24539,N_16455,N_15832);
and U24540 (N_24540,N_17834,N_19914);
nor U24541 (N_24541,N_17608,N_18671);
and U24542 (N_24542,N_16005,N_17910);
nand U24543 (N_24543,N_17293,N_15444);
xnor U24544 (N_24544,N_16788,N_18146);
nand U24545 (N_24545,N_18456,N_15002);
or U24546 (N_24546,N_18245,N_18581);
or U24547 (N_24547,N_16579,N_15969);
xor U24548 (N_24548,N_18735,N_16607);
nand U24549 (N_24549,N_16159,N_19973);
or U24550 (N_24550,N_18895,N_15342);
nor U24551 (N_24551,N_19658,N_17832);
nand U24552 (N_24552,N_19170,N_17703);
and U24553 (N_24553,N_15045,N_15919);
and U24554 (N_24554,N_15717,N_18933);
xor U24555 (N_24555,N_18440,N_18581);
nand U24556 (N_24556,N_16317,N_18133);
xnor U24557 (N_24557,N_15831,N_16978);
and U24558 (N_24558,N_16676,N_17286);
xor U24559 (N_24559,N_19484,N_18254);
nand U24560 (N_24560,N_16273,N_17866);
and U24561 (N_24561,N_15969,N_15319);
xnor U24562 (N_24562,N_15936,N_19997);
xor U24563 (N_24563,N_16386,N_16282);
nand U24564 (N_24564,N_15794,N_18419);
and U24565 (N_24565,N_16278,N_16919);
and U24566 (N_24566,N_19739,N_16489);
nand U24567 (N_24567,N_17018,N_18875);
xnor U24568 (N_24568,N_15303,N_19710);
and U24569 (N_24569,N_15819,N_16492);
nor U24570 (N_24570,N_17854,N_18412);
or U24571 (N_24571,N_17943,N_18132);
or U24572 (N_24572,N_17322,N_16453);
and U24573 (N_24573,N_19037,N_18876);
or U24574 (N_24574,N_17353,N_18943);
nor U24575 (N_24575,N_17091,N_19986);
nand U24576 (N_24576,N_17105,N_17279);
nor U24577 (N_24577,N_18185,N_18059);
nand U24578 (N_24578,N_18015,N_16221);
nand U24579 (N_24579,N_19323,N_17369);
and U24580 (N_24580,N_17613,N_15639);
and U24581 (N_24581,N_17721,N_15014);
and U24582 (N_24582,N_17836,N_17342);
and U24583 (N_24583,N_16388,N_17186);
nand U24584 (N_24584,N_18380,N_18991);
or U24585 (N_24585,N_18998,N_16136);
or U24586 (N_24586,N_18663,N_19471);
nand U24587 (N_24587,N_17053,N_18596);
xor U24588 (N_24588,N_15760,N_15026);
xnor U24589 (N_24589,N_17731,N_17780);
and U24590 (N_24590,N_15935,N_19781);
and U24591 (N_24591,N_19111,N_19560);
nor U24592 (N_24592,N_16234,N_18601);
nor U24593 (N_24593,N_19963,N_18042);
or U24594 (N_24594,N_15409,N_16681);
and U24595 (N_24595,N_18642,N_17632);
nand U24596 (N_24596,N_15527,N_17740);
or U24597 (N_24597,N_16941,N_16893);
and U24598 (N_24598,N_15540,N_18363);
nor U24599 (N_24599,N_16946,N_17313);
nand U24600 (N_24600,N_18534,N_18083);
or U24601 (N_24601,N_17058,N_16127);
or U24602 (N_24602,N_17510,N_17043);
xnor U24603 (N_24603,N_17258,N_15301);
or U24604 (N_24604,N_15344,N_17831);
nor U24605 (N_24605,N_17275,N_19877);
xor U24606 (N_24606,N_18259,N_18510);
nand U24607 (N_24607,N_15650,N_16933);
nand U24608 (N_24608,N_15850,N_17867);
nand U24609 (N_24609,N_15039,N_18220);
or U24610 (N_24610,N_18890,N_18270);
and U24611 (N_24611,N_19021,N_16264);
xnor U24612 (N_24612,N_17893,N_15860);
nand U24613 (N_24613,N_19313,N_17152);
xor U24614 (N_24614,N_17380,N_17418);
and U24615 (N_24615,N_18088,N_18586);
nor U24616 (N_24616,N_15492,N_19240);
xnor U24617 (N_24617,N_15751,N_18073);
or U24618 (N_24618,N_16049,N_17537);
nor U24619 (N_24619,N_17575,N_18619);
or U24620 (N_24620,N_18889,N_16699);
nand U24621 (N_24621,N_16537,N_15359);
and U24622 (N_24622,N_15765,N_16633);
xor U24623 (N_24623,N_17754,N_18502);
xor U24624 (N_24624,N_17942,N_19697);
or U24625 (N_24625,N_19955,N_16115);
nor U24626 (N_24626,N_17215,N_17511);
xor U24627 (N_24627,N_19751,N_19310);
nand U24628 (N_24628,N_16812,N_16626);
xor U24629 (N_24629,N_17520,N_15280);
xor U24630 (N_24630,N_15481,N_19250);
nand U24631 (N_24631,N_19859,N_17745);
nor U24632 (N_24632,N_16193,N_18994);
xor U24633 (N_24633,N_19015,N_15821);
nand U24634 (N_24634,N_16786,N_16140);
and U24635 (N_24635,N_19047,N_18738);
nor U24636 (N_24636,N_18187,N_18548);
xor U24637 (N_24637,N_17749,N_17738);
nor U24638 (N_24638,N_15244,N_17888);
nor U24639 (N_24639,N_16921,N_17052);
and U24640 (N_24640,N_18104,N_19457);
xnor U24641 (N_24641,N_18783,N_15194);
and U24642 (N_24642,N_17306,N_17414);
xor U24643 (N_24643,N_16636,N_17854);
or U24644 (N_24644,N_18830,N_15031);
and U24645 (N_24645,N_15529,N_18568);
nor U24646 (N_24646,N_19284,N_18119);
nor U24647 (N_24647,N_18466,N_19194);
and U24648 (N_24648,N_19683,N_16989);
nand U24649 (N_24649,N_17090,N_15691);
xnor U24650 (N_24650,N_16544,N_15691);
or U24651 (N_24651,N_18414,N_15752);
or U24652 (N_24652,N_17658,N_17589);
nand U24653 (N_24653,N_15169,N_17230);
and U24654 (N_24654,N_19973,N_19911);
and U24655 (N_24655,N_19305,N_17534);
xor U24656 (N_24656,N_18894,N_19687);
nor U24657 (N_24657,N_18191,N_19554);
and U24658 (N_24658,N_18546,N_19528);
nand U24659 (N_24659,N_16481,N_18247);
or U24660 (N_24660,N_17423,N_17791);
nor U24661 (N_24661,N_17994,N_19248);
nand U24662 (N_24662,N_15730,N_16292);
nor U24663 (N_24663,N_19974,N_19923);
xnor U24664 (N_24664,N_16198,N_15801);
or U24665 (N_24665,N_19335,N_17470);
and U24666 (N_24666,N_18038,N_16352);
nand U24667 (N_24667,N_16492,N_15419);
and U24668 (N_24668,N_18013,N_17460);
nor U24669 (N_24669,N_17033,N_16595);
xnor U24670 (N_24670,N_19427,N_19085);
or U24671 (N_24671,N_17255,N_17854);
or U24672 (N_24672,N_15065,N_16685);
and U24673 (N_24673,N_17644,N_17636);
and U24674 (N_24674,N_17305,N_19814);
and U24675 (N_24675,N_17099,N_15220);
nor U24676 (N_24676,N_17945,N_15683);
or U24677 (N_24677,N_18916,N_16690);
or U24678 (N_24678,N_18938,N_18130);
or U24679 (N_24679,N_18426,N_18554);
nor U24680 (N_24680,N_15238,N_19336);
xnor U24681 (N_24681,N_18837,N_17197);
nand U24682 (N_24682,N_19294,N_19636);
nand U24683 (N_24683,N_16705,N_17110);
or U24684 (N_24684,N_18188,N_19616);
or U24685 (N_24685,N_19301,N_19929);
xor U24686 (N_24686,N_16897,N_15301);
or U24687 (N_24687,N_18156,N_18289);
or U24688 (N_24688,N_18872,N_17757);
nand U24689 (N_24689,N_16579,N_15301);
or U24690 (N_24690,N_15461,N_17549);
nor U24691 (N_24691,N_17684,N_15302);
nor U24692 (N_24692,N_15995,N_19726);
xor U24693 (N_24693,N_15112,N_15766);
nor U24694 (N_24694,N_18079,N_16610);
or U24695 (N_24695,N_16553,N_18801);
and U24696 (N_24696,N_15885,N_15158);
nor U24697 (N_24697,N_18840,N_15601);
nor U24698 (N_24698,N_15610,N_18120);
nand U24699 (N_24699,N_16813,N_18459);
nand U24700 (N_24700,N_18598,N_15054);
nand U24701 (N_24701,N_18768,N_19377);
nand U24702 (N_24702,N_15935,N_19981);
nand U24703 (N_24703,N_15623,N_19747);
xnor U24704 (N_24704,N_17456,N_15446);
xor U24705 (N_24705,N_18886,N_15705);
and U24706 (N_24706,N_17223,N_19834);
and U24707 (N_24707,N_15607,N_18259);
nand U24708 (N_24708,N_19475,N_17448);
nand U24709 (N_24709,N_16825,N_19585);
nor U24710 (N_24710,N_19159,N_15701);
nand U24711 (N_24711,N_18149,N_17319);
xor U24712 (N_24712,N_17290,N_19850);
nand U24713 (N_24713,N_18887,N_15691);
nand U24714 (N_24714,N_18915,N_18439);
and U24715 (N_24715,N_16374,N_15046);
nor U24716 (N_24716,N_19794,N_19248);
nand U24717 (N_24717,N_16061,N_18919);
and U24718 (N_24718,N_18850,N_17424);
or U24719 (N_24719,N_15473,N_15321);
or U24720 (N_24720,N_19674,N_16512);
nand U24721 (N_24721,N_18905,N_15396);
and U24722 (N_24722,N_18975,N_19538);
and U24723 (N_24723,N_16556,N_17350);
and U24724 (N_24724,N_15609,N_18548);
or U24725 (N_24725,N_15918,N_16921);
xor U24726 (N_24726,N_16676,N_16941);
nand U24727 (N_24727,N_18870,N_19957);
or U24728 (N_24728,N_15799,N_17672);
or U24729 (N_24729,N_18740,N_19202);
or U24730 (N_24730,N_19993,N_19281);
or U24731 (N_24731,N_15278,N_15891);
nor U24732 (N_24732,N_17147,N_19740);
nand U24733 (N_24733,N_18861,N_17691);
nor U24734 (N_24734,N_16072,N_18116);
nor U24735 (N_24735,N_19398,N_15289);
nor U24736 (N_24736,N_15139,N_18453);
xor U24737 (N_24737,N_15995,N_18290);
xor U24738 (N_24738,N_17807,N_16603);
nor U24739 (N_24739,N_16937,N_17218);
and U24740 (N_24740,N_17110,N_19031);
or U24741 (N_24741,N_16406,N_19553);
or U24742 (N_24742,N_19059,N_18703);
nor U24743 (N_24743,N_18993,N_18866);
xor U24744 (N_24744,N_15099,N_16282);
nand U24745 (N_24745,N_19679,N_18952);
xnor U24746 (N_24746,N_18732,N_17884);
and U24747 (N_24747,N_17836,N_16479);
nand U24748 (N_24748,N_15851,N_19506);
nor U24749 (N_24749,N_19666,N_17342);
and U24750 (N_24750,N_16969,N_19627);
xnor U24751 (N_24751,N_15570,N_16457);
xor U24752 (N_24752,N_15546,N_16510);
nand U24753 (N_24753,N_18742,N_15864);
and U24754 (N_24754,N_19518,N_16989);
nor U24755 (N_24755,N_16450,N_17964);
nor U24756 (N_24756,N_19105,N_18078);
or U24757 (N_24757,N_18711,N_17098);
or U24758 (N_24758,N_17389,N_16314);
xor U24759 (N_24759,N_17181,N_16200);
xor U24760 (N_24760,N_19183,N_19110);
or U24761 (N_24761,N_18721,N_16208);
xor U24762 (N_24762,N_17934,N_19627);
nand U24763 (N_24763,N_18233,N_17081);
nand U24764 (N_24764,N_16253,N_18830);
and U24765 (N_24765,N_17113,N_17516);
or U24766 (N_24766,N_19348,N_16423);
xor U24767 (N_24767,N_17020,N_16188);
nor U24768 (N_24768,N_15527,N_18544);
nor U24769 (N_24769,N_17581,N_16559);
and U24770 (N_24770,N_16516,N_18505);
xor U24771 (N_24771,N_18203,N_15855);
or U24772 (N_24772,N_17039,N_15184);
or U24773 (N_24773,N_16391,N_16432);
nand U24774 (N_24774,N_17496,N_17981);
nor U24775 (N_24775,N_17256,N_19567);
or U24776 (N_24776,N_19002,N_15782);
xor U24777 (N_24777,N_16578,N_16216);
xnor U24778 (N_24778,N_15413,N_19586);
or U24779 (N_24779,N_15338,N_16861);
or U24780 (N_24780,N_17262,N_16831);
nand U24781 (N_24781,N_19092,N_17020);
or U24782 (N_24782,N_17512,N_17006);
nand U24783 (N_24783,N_15773,N_19525);
and U24784 (N_24784,N_16666,N_18217);
and U24785 (N_24785,N_15923,N_17868);
and U24786 (N_24786,N_18058,N_16568);
nor U24787 (N_24787,N_16521,N_18386);
xor U24788 (N_24788,N_16050,N_18213);
and U24789 (N_24789,N_16393,N_16019);
xnor U24790 (N_24790,N_15950,N_17370);
xor U24791 (N_24791,N_16082,N_19860);
nor U24792 (N_24792,N_15699,N_15258);
nor U24793 (N_24793,N_18221,N_18635);
nand U24794 (N_24794,N_18818,N_19694);
xor U24795 (N_24795,N_18458,N_15426);
nor U24796 (N_24796,N_15067,N_18203);
nor U24797 (N_24797,N_15594,N_18146);
xnor U24798 (N_24798,N_19760,N_16265);
nand U24799 (N_24799,N_18232,N_19355);
nor U24800 (N_24800,N_18579,N_18815);
nor U24801 (N_24801,N_18102,N_17791);
xnor U24802 (N_24802,N_16291,N_18399);
nand U24803 (N_24803,N_19699,N_17120);
or U24804 (N_24804,N_16605,N_17631);
or U24805 (N_24805,N_18594,N_15521);
or U24806 (N_24806,N_19249,N_16136);
xor U24807 (N_24807,N_19978,N_16200);
or U24808 (N_24808,N_15914,N_17199);
or U24809 (N_24809,N_16197,N_15255);
and U24810 (N_24810,N_15134,N_16223);
nand U24811 (N_24811,N_19941,N_19171);
nor U24812 (N_24812,N_17123,N_19309);
or U24813 (N_24813,N_17995,N_17187);
nand U24814 (N_24814,N_15841,N_19538);
or U24815 (N_24815,N_18095,N_18556);
and U24816 (N_24816,N_17204,N_18550);
or U24817 (N_24817,N_17301,N_17169);
or U24818 (N_24818,N_17782,N_19742);
nor U24819 (N_24819,N_16483,N_16627);
nand U24820 (N_24820,N_18079,N_17428);
nor U24821 (N_24821,N_18574,N_15603);
xnor U24822 (N_24822,N_18494,N_17815);
or U24823 (N_24823,N_19879,N_17466);
or U24824 (N_24824,N_18605,N_16776);
nand U24825 (N_24825,N_18253,N_16774);
nor U24826 (N_24826,N_18853,N_19115);
nand U24827 (N_24827,N_18353,N_15460);
or U24828 (N_24828,N_18992,N_16145);
xnor U24829 (N_24829,N_19444,N_15778);
and U24830 (N_24830,N_17735,N_17522);
xnor U24831 (N_24831,N_19485,N_17815);
nor U24832 (N_24832,N_18311,N_15837);
or U24833 (N_24833,N_19225,N_19991);
nor U24834 (N_24834,N_16942,N_19840);
or U24835 (N_24835,N_19320,N_17573);
xnor U24836 (N_24836,N_17889,N_17256);
nand U24837 (N_24837,N_15444,N_15971);
nor U24838 (N_24838,N_16773,N_18467);
nand U24839 (N_24839,N_19361,N_16372);
or U24840 (N_24840,N_15000,N_18588);
xnor U24841 (N_24841,N_16552,N_18929);
and U24842 (N_24842,N_17154,N_15302);
xor U24843 (N_24843,N_17473,N_18393);
nor U24844 (N_24844,N_19869,N_18722);
or U24845 (N_24845,N_15635,N_17843);
or U24846 (N_24846,N_19044,N_15333);
and U24847 (N_24847,N_19891,N_15599);
or U24848 (N_24848,N_15301,N_19439);
nor U24849 (N_24849,N_19035,N_17339);
or U24850 (N_24850,N_18230,N_19506);
xnor U24851 (N_24851,N_19748,N_17029);
nand U24852 (N_24852,N_15280,N_18900);
nand U24853 (N_24853,N_18570,N_15166);
xnor U24854 (N_24854,N_18246,N_19887);
and U24855 (N_24855,N_19816,N_16202);
xnor U24856 (N_24856,N_16632,N_15992);
or U24857 (N_24857,N_19376,N_15883);
nand U24858 (N_24858,N_19717,N_16732);
and U24859 (N_24859,N_15492,N_15108);
nand U24860 (N_24860,N_18898,N_18080);
or U24861 (N_24861,N_16281,N_15484);
or U24862 (N_24862,N_18229,N_15949);
and U24863 (N_24863,N_17454,N_16373);
and U24864 (N_24864,N_16371,N_17961);
or U24865 (N_24865,N_15536,N_19799);
xnor U24866 (N_24866,N_15907,N_15595);
or U24867 (N_24867,N_17913,N_15159);
or U24868 (N_24868,N_16407,N_18630);
xnor U24869 (N_24869,N_15552,N_17553);
and U24870 (N_24870,N_15019,N_15589);
xnor U24871 (N_24871,N_15333,N_17867);
or U24872 (N_24872,N_19714,N_16549);
nand U24873 (N_24873,N_19063,N_19273);
and U24874 (N_24874,N_18380,N_15016);
nand U24875 (N_24875,N_15291,N_19367);
nand U24876 (N_24876,N_15207,N_15570);
and U24877 (N_24877,N_17414,N_15832);
or U24878 (N_24878,N_15582,N_18921);
nand U24879 (N_24879,N_16172,N_15791);
or U24880 (N_24880,N_18517,N_18850);
xnor U24881 (N_24881,N_18796,N_19339);
or U24882 (N_24882,N_17446,N_16129);
nand U24883 (N_24883,N_15502,N_17433);
and U24884 (N_24884,N_18827,N_19367);
nand U24885 (N_24885,N_19925,N_17953);
nand U24886 (N_24886,N_17899,N_15700);
or U24887 (N_24887,N_16531,N_16333);
nand U24888 (N_24888,N_15797,N_17604);
and U24889 (N_24889,N_16298,N_17677);
or U24890 (N_24890,N_18039,N_15395);
and U24891 (N_24891,N_19473,N_16907);
and U24892 (N_24892,N_18716,N_15291);
or U24893 (N_24893,N_19263,N_15822);
or U24894 (N_24894,N_19659,N_15677);
and U24895 (N_24895,N_19580,N_19501);
nor U24896 (N_24896,N_16146,N_17279);
and U24897 (N_24897,N_17536,N_15747);
or U24898 (N_24898,N_18491,N_19247);
or U24899 (N_24899,N_17477,N_19897);
or U24900 (N_24900,N_15100,N_15501);
or U24901 (N_24901,N_16705,N_15171);
or U24902 (N_24902,N_18677,N_15555);
nor U24903 (N_24903,N_17654,N_17243);
nor U24904 (N_24904,N_19372,N_17060);
nand U24905 (N_24905,N_16600,N_17239);
and U24906 (N_24906,N_15335,N_16589);
xor U24907 (N_24907,N_16003,N_18504);
and U24908 (N_24908,N_19096,N_17029);
and U24909 (N_24909,N_16861,N_17822);
nand U24910 (N_24910,N_16465,N_19128);
nand U24911 (N_24911,N_18279,N_15142);
and U24912 (N_24912,N_18199,N_16111);
nor U24913 (N_24913,N_15626,N_15654);
nand U24914 (N_24914,N_16628,N_16583);
nand U24915 (N_24915,N_17043,N_19736);
nand U24916 (N_24916,N_18887,N_19180);
xnor U24917 (N_24917,N_18334,N_16522);
or U24918 (N_24918,N_15637,N_18889);
or U24919 (N_24919,N_19496,N_18254);
xnor U24920 (N_24920,N_15354,N_15382);
xor U24921 (N_24921,N_17560,N_18104);
nand U24922 (N_24922,N_19589,N_15786);
and U24923 (N_24923,N_18248,N_15929);
and U24924 (N_24924,N_15158,N_15537);
nand U24925 (N_24925,N_18252,N_19296);
nand U24926 (N_24926,N_16154,N_17976);
or U24927 (N_24927,N_16965,N_16186);
nand U24928 (N_24928,N_18835,N_17882);
nand U24929 (N_24929,N_17761,N_17145);
nor U24930 (N_24930,N_16626,N_18117);
nand U24931 (N_24931,N_15936,N_16720);
nand U24932 (N_24932,N_15722,N_17190);
nand U24933 (N_24933,N_18898,N_19813);
xnor U24934 (N_24934,N_15605,N_15760);
or U24935 (N_24935,N_17401,N_15743);
or U24936 (N_24936,N_15710,N_18992);
and U24937 (N_24937,N_15590,N_16912);
and U24938 (N_24938,N_17806,N_18749);
and U24939 (N_24939,N_15278,N_17784);
xnor U24940 (N_24940,N_17703,N_16334);
nand U24941 (N_24941,N_17705,N_17993);
xnor U24942 (N_24942,N_15641,N_18882);
and U24943 (N_24943,N_17072,N_16839);
nor U24944 (N_24944,N_19863,N_16549);
and U24945 (N_24945,N_15232,N_16849);
xor U24946 (N_24946,N_17875,N_17920);
nor U24947 (N_24947,N_17715,N_15364);
and U24948 (N_24948,N_18177,N_15857);
and U24949 (N_24949,N_19575,N_15939);
nor U24950 (N_24950,N_16734,N_17147);
nor U24951 (N_24951,N_17457,N_16698);
nor U24952 (N_24952,N_17810,N_19368);
or U24953 (N_24953,N_19054,N_15928);
nor U24954 (N_24954,N_16816,N_19460);
xnor U24955 (N_24955,N_19853,N_19528);
and U24956 (N_24956,N_16904,N_16398);
or U24957 (N_24957,N_19219,N_17470);
or U24958 (N_24958,N_16602,N_17826);
and U24959 (N_24959,N_18916,N_17979);
or U24960 (N_24960,N_15955,N_17730);
and U24961 (N_24961,N_16550,N_19130);
nor U24962 (N_24962,N_19662,N_17805);
or U24963 (N_24963,N_19537,N_16747);
nand U24964 (N_24964,N_16271,N_17488);
nand U24965 (N_24965,N_16548,N_18335);
and U24966 (N_24966,N_15619,N_17751);
and U24967 (N_24967,N_16642,N_18905);
and U24968 (N_24968,N_18370,N_15422);
or U24969 (N_24969,N_15207,N_17428);
nand U24970 (N_24970,N_15100,N_16438);
and U24971 (N_24971,N_17277,N_16381);
or U24972 (N_24972,N_18195,N_19497);
nor U24973 (N_24973,N_17047,N_15744);
and U24974 (N_24974,N_17691,N_17910);
nand U24975 (N_24975,N_17813,N_15284);
and U24976 (N_24976,N_15836,N_19229);
nand U24977 (N_24977,N_19790,N_16299);
nand U24978 (N_24978,N_17221,N_17910);
nand U24979 (N_24979,N_19062,N_16850);
or U24980 (N_24980,N_18113,N_17944);
and U24981 (N_24981,N_15801,N_18957);
nor U24982 (N_24982,N_18527,N_19864);
or U24983 (N_24983,N_17438,N_17455);
and U24984 (N_24984,N_15715,N_16824);
nor U24985 (N_24985,N_19799,N_19689);
and U24986 (N_24986,N_19499,N_19366);
xor U24987 (N_24987,N_16545,N_19391);
nor U24988 (N_24988,N_17276,N_18671);
xnor U24989 (N_24989,N_15293,N_17356);
or U24990 (N_24990,N_16170,N_15379);
and U24991 (N_24991,N_16363,N_18409);
nand U24992 (N_24992,N_15788,N_15564);
or U24993 (N_24993,N_19639,N_16668);
nand U24994 (N_24994,N_19585,N_18446);
or U24995 (N_24995,N_15775,N_16199);
or U24996 (N_24996,N_15913,N_17972);
nand U24997 (N_24997,N_15669,N_15018);
nor U24998 (N_24998,N_16413,N_16982);
or U24999 (N_24999,N_18579,N_17306);
nor UO_0 (O_0,N_21199,N_23713);
or UO_1 (O_1,N_24537,N_24329);
nor UO_2 (O_2,N_24873,N_23246);
nand UO_3 (O_3,N_24415,N_20480);
nand UO_4 (O_4,N_22870,N_20094);
nor UO_5 (O_5,N_23849,N_22694);
and UO_6 (O_6,N_22071,N_21051);
xor UO_7 (O_7,N_24094,N_24503);
nor UO_8 (O_8,N_24919,N_23293);
xor UO_9 (O_9,N_22889,N_21813);
and UO_10 (O_10,N_20231,N_21423);
and UO_11 (O_11,N_23747,N_24476);
nor UO_12 (O_12,N_21574,N_23154);
nor UO_13 (O_13,N_21479,N_22545);
xnor UO_14 (O_14,N_22702,N_20404);
and UO_15 (O_15,N_24064,N_21755);
nand UO_16 (O_16,N_21925,N_20115);
nand UO_17 (O_17,N_23591,N_22407);
nor UO_18 (O_18,N_20758,N_21304);
xnor UO_19 (O_19,N_21689,N_21144);
nand UO_20 (O_20,N_20360,N_23541);
or UO_21 (O_21,N_22267,N_23385);
nand UO_22 (O_22,N_20046,N_20336);
xor UO_23 (O_23,N_21616,N_23182);
nand UO_24 (O_24,N_22945,N_24286);
and UO_25 (O_25,N_20259,N_24167);
or UO_26 (O_26,N_21712,N_21907);
xor UO_27 (O_27,N_23034,N_23181);
nand UO_28 (O_28,N_23267,N_22077);
nand UO_29 (O_29,N_20414,N_24275);
xnor UO_30 (O_30,N_20446,N_24558);
or UO_31 (O_31,N_23627,N_23798);
nor UO_32 (O_32,N_20813,N_23592);
xor UO_33 (O_33,N_24554,N_23758);
and UO_34 (O_34,N_24899,N_22848);
or UO_35 (O_35,N_21221,N_22719);
and UO_36 (O_36,N_23978,N_23765);
nor UO_37 (O_37,N_23669,N_20654);
nor UO_38 (O_38,N_24666,N_22661);
nor UO_39 (O_39,N_24788,N_20174);
nand UO_40 (O_40,N_20235,N_21254);
and UO_41 (O_41,N_22014,N_21873);
nor UO_42 (O_42,N_22191,N_20469);
nor UO_43 (O_43,N_20036,N_21333);
nor UO_44 (O_44,N_20303,N_22975);
and UO_45 (O_45,N_20605,N_23909);
or UO_46 (O_46,N_21128,N_20734);
nor UO_47 (O_47,N_24137,N_21795);
nor UO_48 (O_48,N_24359,N_21849);
nand UO_49 (O_49,N_22492,N_21044);
and UO_50 (O_50,N_20843,N_22557);
and UO_51 (O_51,N_23263,N_24341);
xor UO_52 (O_52,N_21968,N_20262);
xor UO_53 (O_53,N_20799,N_20375);
nand UO_54 (O_54,N_20715,N_22086);
nor UO_55 (O_55,N_23147,N_24163);
nand UO_56 (O_56,N_21883,N_23323);
nor UO_57 (O_57,N_24947,N_21361);
nor UO_58 (O_58,N_24598,N_24457);
xor UO_59 (O_59,N_23214,N_24791);
xor UO_60 (O_60,N_20114,N_22368);
xor UO_61 (O_61,N_20385,N_21776);
xnor UO_62 (O_62,N_21604,N_24195);
and UO_63 (O_63,N_21271,N_22477);
or UO_64 (O_64,N_20471,N_21154);
nor UO_65 (O_65,N_23762,N_22706);
nand UO_66 (O_66,N_24879,N_24378);
nor UO_67 (O_67,N_20570,N_22533);
and UO_68 (O_68,N_22094,N_23693);
or UO_69 (O_69,N_20678,N_23466);
xor UO_70 (O_70,N_21425,N_21259);
and UO_71 (O_71,N_23530,N_23371);
xor UO_72 (O_72,N_22644,N_20107);
or UO_73 (O_73,N_21684,N_20517);
nor UO_74 (O_74,N_22673,N_21270);
nand UO_75 (O_75,N_21920,N_21892);
xnor UO_76 (O_76,N_20428,N_22453);
and UO_77 (O_77,N_22118,N_20226);
or UO_78 (O_78,N_23170,N_21588);
or UO_79 (O_79,N_22339,N_20940);
xor UO_80 (O_80,N_23516,N_20892);
or UO_81 (O_81,N_20351,N_22507);
nor UO_82 (O_82,N_24015,N_20900);
nand UO_83 (O_83,N_24173,N_24135);
xnor UO_84 (O_84,N_24726,N_21420);
or UO_85 (O_85,N_23876,N_23949);
nand UO_86 (O_86,N_21295,N_23284);
xnor UO_87 (O_87,N_23957,N_21454);
nor UO_88 (O_88,N_23377,N_22396);
xor UO_89 (O_89,N_24449,N_24201);
or UO_90 (O_90,N_21785,N_23330);
and UO_91 (O_91,N_20111,N_22307);
and UO_92 (O_92,N_24865,N_20002);
nand UO_93 (O_93,N_20518,N_23690);
xor UO_94 (O_94,N_22567,N_21797);
nor UO_95 (O_95,N_24463,N_21758);
nor UO_96 (O_96,N_21284,N_23831);
nor UO_97 (O_97,N_23847,N_21382);
and UO_98 (O_98,N_20443,N_20688);
or UO_99 (O_99,N_21789,N_23917);
nand UO_100 (O_100,N_20060,N_24351);
nand UO_101 (O_101,N_20755,N_24908);
nand UO_102 (O_102,N_20902,N_24453);
nand UO_103 (O_103,N_22560,N_22050);
nor UO_104 (O_104,N_23929,N_23302);
xnor UO_105 (O_105,N_20301,N_23003);
xor UO_106 (O_106,N_20812,N_23961);
or UO_107 (O_107,N_24233,N_24701);
or UO_108 (O_108,N_23584,N_23059);
nor UO_109 (O_109,N_22640,N_20402);
and UO_110 (O_110,N_21083,N_21236);
nand UO_111 (O_111,N_22604,N_21895);
or UO_112 (O_112,N_22595,N_24176);
xor UO_113 (O_113,N_23103,N_21336);
xor UO_114 (O_114,N_20834,N_23020);
or UO_115 (O_115,N_24288,N_23763);
nand UO_116 (O_116,N_24221,N_21214);
xnor UO_117 (O_117,N_22419,N_22073);
nor UO_118 (O_118,N_24727,N_24323);
or UO_119 (O_119,N_22863,N_21028);
xor UO_120 (O_120,N_23060,N_23022);
or UO_121 (O_121,N_24047,N_21224);
or UO_122 (O_122,N_23805,N_24208);
xor UO_123 (O_123,N_22844,N_21519);
and UO_124 (O_124,N_24533,N_22357);
xnor UO_125 (O_125,N_23572,N_21134);
nor UO_126 (O_126,N_23688,N_21601);
nor UO_127 (O_127,N_24800,N_22808);
and UO_128 (O_128,N_24238,N_20559);
nor UO_129 (O_129,N_20269,N_21081);
nand UO_130 (O_130,N_21498,N_24615);
xnor UO_131 (O_131,N_23328,N_22196);
nor UO_132 (O_132,N_23485,N_22989);
nand UO_133 (O_133,N_24877,N_21411);
and UO_134 (O_134,N_21357,N_21025);
or UO_135 (O_135,N_23634,N_23667);
nor UO_136 (O_136,N_21335,N_21590);
nor UO_137 (O_137,N_23455,N_23185);
or UO_138 (O_138,N_24540,N_21978);
xnor UO_139 (O_139,N_23237,N_20791);
nand UO_140 (O_140,N_24355,N_23434);
or UO_141 (O_141,N_20736,N_24160);
xor UO_142 (O_142,N_24373,N_21235);
or UO_143 (O_143,N_23908,N_23474);
or UO_144 (O_144,N_24635,N_24215);
nor UO_145 (O_145,N_24369,N_23295);
nor UO_146 (O_146,N_23157,N_24515);
or UO_147 (O_147,N_22606,N_23991);
nand UO_148 (O_148,N_23934,N_24027);
nor UO_149 (O_149,N_20622,N_24979);
or UO_150 (O_150,N_24997,N_24781);
nand UO_151 (O_151,N_24614,N_20088);
xnor UO_152 (O_152,N_22963,N_22156);
or UO_153 (O_153,N_21072,N_21408);
nor UO_154 (O_154,N_22804,N_21084);
or UO_155 (O_155,N_23470,N_20143);
nand UO_156 (O_156,N_22360,N_20651);
nand UO_157 (O_157,N_24009,N_24092);
or UO_158 (O_158,N_24571,N_21954);
xor UO_159 (O_159,N_21359,N_21865);
or UO_160 (O_160,N_20390,N_24769);
nand UO_161 (O_161,N_20105,N_24721);
and UO_162 (O_162,N_20696,N_20358);
nand UO_163 (O_163,N_23821,N_23508);
nor UO_164 (O_164,N_22655,N_23895);
xor UO_165 (O_165,N_24446,N_20337);
xnor UO_166 (O_166,N_24656,N_23538);
and UO_167 (O_167,N_23160,N_22790);
nor UO_168 (O_168,N_20121,N_24146);
xor UO_169 (O_169,N_24921,N_21248);
nor UO_170 (O_170,N_23902,N_22389);
or UO_171 (O_171,N_22646,N_20242);
nand UO_172 (O_172,N_20458,N_22459);
or UO_173 (O_173,N_21662,N_22802);
nand UO_174 (O_174,N_20332,N_21265);
and UO_175 (O_175,N_21343,N_21063);
nor UO_176 (O_176,N_20648,N_22856);
xnor UO_177 (O_177,N_23412,N_23178);
or UO_178 (O_178,N_22705,N_24778);
nor UO_179 (O_179,N_21204,N_21914);
or UO_180 (O_180,N_22377,N_21033);
and UO_181 (O_181,N_23054,N_22809);
and UO_182 (O_182,N_22918,N_20700);
or UO_183 (O_183,N_24202,N_22337);
nand UO_184 (O_184,N_22229,N_20562);
or UO_185 (O_185,N_20815,N_20701);
nand UO_186 (O_186,N_21798,N_22596);
or UO_187 (O_187,N_22427,N_21419);
and UO_188 (O_188,N_24690,N_24290);
and UO_189 (O_189,N_24179,N_24093);
nand UO_190 (O_190,N_24466,N_21294);
or UO_191 (O_191,N_21185,N_22813);
nand UO_192 (O_192,N_23832,N_20667);
nand UO_193 (O_193,N_23623,N_20213);
xnor UO_194 (O_194,N_21181,N_21609);
xnor UO_195 (O_195,N_24244,N_20160);
and UO_196 (O_196,N_22738,N_20604);
xor UO_197 (O_197,N_23743,N_21014);
and UO_198 (O_198,N_20074,N_23979);
and UO_199 (O_199,N_20986,N_20705);
and UO_200 (O_200,N_22217,N_20629);
xnor UO_201 (O_201,N_24191,N_22394);
nor UO_202 (O_202,N_22944,N_21822);
and UO_203 (O_203,N_20208,N_23522);
and UO_204 (O_204,N_22031,N_24364);
and UO_205 (O_205,N_23988,N_22263);
or UO_206 (O_206,N_20221,N_21451);
nand UO_207 (O_207,N_24175,N_21661);
nor UO_208 (O_208,N_23777,N_22212);
xor UO_209 (O_209,N_20664,N_20322);
xor UO_210 (O_210,N_23676,N_22835);
or UO_211 (O_211,N_21735,N_22351);
nor UO_212 (O_212,N_20833,N_20917);
nor UO_213 (O_213,N_23685,N_24991);
nand UO_214 (O_214,N_24795,N_20253);
and UO_215 (O_215,N_23464,N_24810);
or UO_216 (O_216,N_21091,N_22950);
and UO_217 (O_217,N_23754,N_20906);
nor UO_218 (O_218,N_21583,N_23035);
and UO_219 (O_219,N_22795,N_20673);
and UO_220 (O_220,N_20426,N_21074);
xor UO_221 (O_221,N_21943,N_24524);
or UO_222 (O_222,N_24096,N_21473);
nor UO_223 (O_223,N_23752,N_21332);
and UO_224 (O_224,N_20842,N_22907);
nor UO_225 (O_225,N_21481,N_20445);
nand UO_226 (O_226,N_22296,N_23550);
or UO_227 (O_227,N_21017,N_23291);
nand UO_228 (O_228,N_24482,N_23131);
xor UO_229 (O_229,N_21029,N_21145);
xnor UO_230 (O_230,N_21971,N_21955);
or UO_231 (O_231,N_22214,N_23332);
and UO_232 (O_232,N_23290,N_24707);
nor UO_233 (O_233,N_21438,N_20492);
or UO_234 (O_234,N_21992,N_21956);
nand UO_235 (O_235,N_22826,N_22162);
nand UO_236 (O_236,N_23027,N_23531);
or UO_237 (O_237,N_20229,N_22842);
nand UO_238 (O_238,N_23241,N_24285);
nand UO_239 (O_239,N_20026,N_20432);
nor UO_240 (O_240,N_20788,N_20412);
nand UO_241 (O_241,N_22636,N_24081);
xnor UO_242 (O_242,N_20408,N_22805);
and UO_243 (O_243,N_21513,N_21200);
xnor UO_244 (O_244,N_24845,N_21685);
or UO_245 (O_245,N_23661,N_23966);
nor UO_246 (O_246,N_21514,N_23459);
nor UO_247 (O_247,N_22778,N_24336);
nand UO_248 (O_248,N_22704,N_22260);
nor UO_249 (O_249,N_24065,N_21958);
or UO_250 (O_250,N_21589,N_23543);
nand UO_251 (O_251,N_21984,N_20248);
and UO_252 (O_252,N_22986,N_24438);
and UO_253 (O_253,N_24264,N_21297);
xor UO_254 (O_254,N_21680,N_24621);
and UO_255 (O_255,N_20091,N_23800);
and UO_256 (O_256,N_21136,N_24079);
and UO_257 (O_257,N_20951,N_21375);
xor UO_258 (O_258,N_21036,N_21430);
and UO_259 (O_259,N_21174,N_23614);
nand UO_260 (O_260,N_21621,N_23827);
nor UO_261 (O_261,N_23318,N_23727);
xnor UO_262 (O_262,N_20218,N_21311);
xor UO_263 (O_263,N_24860,N_23636);
nor UO_264 (O_264,N_22581,N_22284);
xor UO_265 (O_265,N_24718,N_24145);
xor UO_266 (O_266,N_23447,N_21833);
xnor UO_267 (O_267,N_23233,N_24594);
or UO_268 (O_268,N_24266,N_22710);
xor UO_269 (O_269,N_22671,N_22448);
xnor UO_270 (O_270,N_21502,N_22592);
xnor UO_271 (O_271,N_20959,N_22574);
and UO_272 (O_272,N_20021,N_24862);
xnor UO_273 (O_273,N_22391,N_22350);
nand UO_274 (O_274,N_21002,N_22752);
nor UO_275 (O_275,N_20545,N_21846);
xor UO_276 (O_276,N_22811,N_24231);
xnor UO_277 (O_277,N_20746,N_21428);
nor UO_278 (O_278,N_23209,N_22353);
or UO_279 (O_279,N_21166,N_23803);
nor UO_280 (O_280,N_24222,N_21614);
or UO_281 (O_281,N_23392,N_22653);
and UO_282 (O_282,N_21815,N_24826);
and UO_283 (O_283,N_20627,N_23726);
and UO_284 (O_284,N_21731,N_21010);
nand UO_285 (O_285,N_22910,N_24715);
xnor UO_286 (O_286,N_20901,N_22895);
xnor UO_287 (O_287,N_21452,N_20274);
or UO_288 (O_288,N_21158,N_20437);
xor UO_289 (O_289,N_21360,N_21276);
xor UO_290 (O_290,N_20858,N_23311);
and UO_291 (O_291,N_22952,N_23383);
nand UO_292 (O_292,N_24057,N_22281);
nand UO_293 (O_293,N_22909,N_23360);
or UO_294 (O_294,N_21391,N_23225);
and UO_295 (O_295,N_22912,N_20095);
or UO_296 (O_296,N_22982,N_22893);
nand UO_297 (O_297,N_21178,N_24517);
xnor UO_298 (O_298,N_20591,N_23565);
or UO_299 (O_299,N_22106,N_23104);
nor UO_300 (O_300,N_23958,N_22046);
or UO_301 (O_301,N_21326,N_23768);
nand UO_302 (O_302,N_24172,N_20324);
or UO_303 (O_303,N_20884,N_24739);
nor UO_304 (O_304,N_20521,N_22248);
nor UO_305 (O_305,N_22463,N_20083);
or UO_306 (O_306,N_20693,N_24892);
xnor UO_307 (O_307,N_23331,N_21022);
xnor UO_308 (O_308,N_24067,N_23899);
nand UO_309 (O_309,N_22257,N_22745);
xnor UO_310 (O_310,N_20924,N_22528);
xnor UO_311 (O_311,N_21837,N_23269);
xnor UO_312 (O_312,N_24539,N_24317);
xor UO_313 (O_313,N_23808,N_20681);
nand UO_314 (O_314,N_23880,N_24210);
nand UO_315 (O_315,N_20044,N_23450);
nand UO_316 (O_316,N_21341,N_22981);
and UO_317 (O_317,N_24082,N_22499);
nand UO_318 (O_318,N_20581,N_23047);
xnor UO_319 (O_319,N_21031,N_24004);
and UO_320 (O_320,N_24780,N_23008);
or UO_321 (O_321,N_21635,N_20587);
and UO_322 (O_322,N_23396,N_20199);
xor UO_323 (O_323,N_20968,N_20668);
or UO_324 (O_324,N_20660,N_20930);
nor UO_325 (O_325,N_22019,N_24768);
nor UO_326 (O_326,N_21140,N_22529);
nand UO_327 (O_327,N_24294,N_24368);
and UO_328 (O_328,N_20364,N_20470);
xor UO_329 (O_329,N_22283,N_24812);
nor UO_330 (O_330,N_21413,N_23195);
nor UO_331 (O_331,N_22408,N_24471);
nand UO_332 (O_332,N_23132,N_20345);
xnor UO_333 (O_333,N_21750,N_20977);
nor UO_334 (O_334,N_22305,N_24134);
or UO_335 (O_335,N_23873,N_23879);
xnor UO_336 (O_336,N_24243,N_24034);
nand UO_337 (O_337,N_23426,N_24439);
nand UO_338 (O_338,N_21222,N_22992);
nor UO_339 (O_339,N_21272,N_23658);
and UO_340 (O_340,N_23981,N_20714);
or UO_341 (O_341,N_22278,N_21277);
and UO_342 (O_342,N_20703,N_21921);
or UO_343 (O_343,N_24646,N_23316);
nand UO_344 (O_344,N_22833,N_20058);
nor UO_345 (O_345,N_24218,N_23930);
nor UO_346 (O_346,N_20120,N_21996);
and UO_347 (O_347,N_23219,N_20739);
nand UO_348 (O_348,N_23493,N_23414);
or UO_349 (O_349,N_22697,N_20465);
nor UO_350 (O_350,N_20214,N_20781);
and UO_351 (O_351,N_23402,N_23420);
nor UO_352 (O_352,N_20707,N_22933);
nor UO_353 (O_353,N_20981,N_20420);
nand UO_354 (O_354,N_23792,N_21654);
nand UO_355 (O_355,N_23753,N_23424);
nor UO_356 (O_356,N_24031,N_23665);
or UO_357 (O_357,N_20975,N_21421);
or UO_358 (O_358,N_24502,N_21133);
or UO_359 (O_359,N_23845,N_23428);
nor UO_360 (O_360,N_21268,N_24050);
and UO_361 (O_361,N_21864,N_23514);
and UO_362 (O_362,N_23918,N_24929);
xor UO_363 (O_363,N_21538,N_20162);
and UO_364 (O_364,N_22227,N_22345);
and UO_365 (O_365,N_23629,N_20729);
nand UO_366 (O_366,N_22195,N_24808);
nor UO_367 (O_367,N_22166,N_23706);
or UO_368 (O_368,N_24869,N_23672);
nand UO_369 (O_369,N_22766,N_20989);
nor UO_370 (O_370,N_24629,N_22798);
xor UO_371 (O_371,N_23708,N_24616);
nor UO_372 (O_372,N_24078,N_24319);
or UO_373 (O_373,N_20575,N_22113);
nor UO_374 (O_374,N_20374,N_24687);
or UO_375 (O_375,N_21390,N_22875);
nand UO_376 (O_376,N_24054,N_23289);
or UO_377 (O_377,N_22017,N_23702);
or UO_378 (O_378,N_23595,N_24330);
or UO_379 (O_379,N_21664,N_20232);
nor UO_380 (O_380,N_20835,N_20383);
and UO_381 (O_381,N_21480,N_21392);
nor UO_382 (O_382,N_22759,N_24634);
or UO_383 (O_383,N_22139,N_24587);
nand UO_384 (O_384,N_22222,N_24550);
nor UO_385 (O_385,N_21827,N_23544);
nor UO_386 (O_386,N_23497,N_21179);
or UO_387 (O_387,N_22502,N_22371);
and UO_388 (O_388,N_20941,N_22615);
nand UO_389 (O_389,N_20683,N_20001);
or UO_390 (O_390,N_20777,N_20600);
nor UO_391 (O_391,N_23996,N_20102);
xnor UO_392 (O_392,N_24824,N_22347);
or UO_393 (O_393,N_20578,N_24933);
nand UO_394 (O_394,N_20376,N_24779);
nand UO_395 (O_395,N_24500,N_23163);
xnor UO_396 (O_396,N_21650,N_20343);
nand UO_397 (O_397,N_22243,N_22897);
nand UO_398 (O_398,N_22550,N_23098);
nor UO_399 (O_399,N_24032,N_24091);
nand UO_400 (O_400,N_23216,N_24362);
or UO_401 (O_401,N_24039,N_23787);
xnor UO_402 (O_402,N_21887,N_22318);
nand UO_403 (O_403,N_22445,N_21993);
or UO_404 (O_404,N_21592,N_24475);
xnor UO_405 (O_405,N_21894,N_24920);
and UO_406 (O_406,N_21637,N_20637);
and UO_407 (O_407,N_21830,N_24040);
nor UO_408 (O_408,N_24118,N_21156);
nor UO_409 (O_409,N_23609,N_23275);
or UO_410 (O_410,N_21879,N_24207);
or UO_411 (O_411,N_22796,N_24255);
nor UO_412 (O_412,N_20439,N_20506);
nand UO_413 (O_413,N_22877,N_20571);
and UO_414 (O_414,N_20104,N_20407);
nand UO_415 (O_415,N_24240,N_21505);
nor UO_416 (O_416,N_22469,N_23553);
xor UO_417 (O_417,N_24561,N_24966);
xnor UO_418 (O_418,N_24886,N_24254);
nor UO_419 (O_419,N_21545,N_22208);
and UO_420 (O_420,N_20388,N_22362);
nand UO_421 (O_421,N_24046,N_23306);
or UO_422 (O_422,N_22092,N_23074);
nor UO_423 (O_423,N_23339,N_23734);
and UO_424 (O_424,N_22979,N_20352);
nor UO_425 (O_425,N_20939,N_22059);
xor UO_426 (O_426,N_20574,N_20685);
and UO_427 (O_427,N_21310,N_22030);
nor UO_428 (O_428,N_20346,N_24949);
and UO_429 (O_429,N_20771,N_20396);
nand UO_430 (O_430,N_23061,N_24682);
nand UO_431 (O_431,N_21322,N_22664);
nand UO_432 (O_432,N_21003,N_22327);
nand UO_433 (O_433,N_22709,N_24575);
or UO_434 (O_434,N_24168,N_20418);
nor UO_435 (O_435,N_20152,N_20459);
or UO_436 (O_436,N_20020,N_20549);
nand UO_437 (O_437,N_24053,N_23458);
nand UO_438 (O_438,N_23631,N_23200);
or UO_439 (O_439,N_21032,N_22896);
xnor UO_440 (O_440,N_24511,N_24388);
and UO_441 (O_441,N_22878,N_20789);
nand UO_442 (O_442,N_22620,N_22652);
xnor UO_443 (O_443,N_24867,N_22876);
xnor UO_444 (O_444,N_21263,N_24427);
nand UO_445 (O_445,N_22633,N_21194);
nand UO_446 (O_446,N_22868,N_20988);
and UO_447 (O_447,N_20820,N_20141);
or UO_448 (O_448,N_24177,N_21959);
and UO_449 (O_449,N_22417,N_21399);
or UO_450 (O_450,N_20669,N_23203);
nand UO_451 (O_451,N_22503,N_22406);
nor UO_452 (O_452,N_24792,N_21707);
xnor UO_453 (O_453,N_20886,N_22899);
xnor UO_454 (O_454,N_24977,N_24102);
nand UO_455 (O_455,N_20960,N_20344);
and UO_456 (O_456,N_24674,N_23144);
xor UO_457 (O_457,N_20603,N_21824);
nand UO_458 (O_458,N_23611,N_22315);
and UO_459 (O_459,N_23612,N_21807);
nand UO_460 (O_460,N_23334,N_22591);
nor UO_461 (O_461,N_20686,N_20866);
xnor UO_462 (O_462,N_22900,N_21985);
and UO_463 (O_463,N_21195,N_21024);
or UO_464 (O_464,N_24596,N_20081);
xnor UO_465 (O_465,N_20034,N_20857);
nor UO_466 (O_466,N_21264,N_22270);
nand UO_467 (O_467,N_22570,N_22971);
nand UO_468 (O_468,N_21525,N_23893);
nor UO_469 (O_469,N_20453,N_22241);
nand UO_470 (O_470,N_20994,N_24352);
xor UO_471 (O_471,N_20010,N_21558);
nor UO_472 (O_472,N_21279,N_20150);
and UO_473 (O_473,N_24685,N_23770);
nor UO_474 (O_474,N_21274,N_24490);
xnor UO_475 (O_475,N_22756,N_20122);
nand UO_476 (O_476,N_22125,N_20524);
and UO_477 (O_477,N_21855,N_20539);
xor UO_478 (O_478,N_22983,N_22882);
and UO_479 (O_479,N_24435,N_24695);
nand UO_480 (O_480,N_24922,N_24915);
nand UO_481 (O_481,N_24732,N_21913);
or UO_482 (O_482,N_23265,N_20136);
xor UO_483 (O_483,N_24833,N_24619);
and UO_484 (O_484,N_23733,N_22236);
nor UO_485 (O_485,N_24220,N_20698);
and UO_486 (O_486,N_22621,N_20348);
nor UO_487 (O_487,N_20225,N_21368);
nand UO_488 (O_488,N_23956,N_22879);
nor UO_489 (O_489,N_22188,N_23348);
xor UO_490 (O_490,N_20185,N_23052);
xnor UO_491 (O_491,N_21871,N_22348);
nand UO_492 (O_492,N_22519,N_23325);
nor UO_493 (O_493,N_21205,N_24601);
nand UO_494 (O_494,N_24291,N_23193);
or UO_495 (O_495,N_20429,N_23883);
nor UO_496 (O_496,N_22980,N_24205);
nor UO_497 (O_497,N_23653,N_22524);
xor UO_498 (O_498,N_23812,N_24247);
xnor UO_499 (O_499,N_21492,N_22112);
nor UO_500 (O_500,N_24608,N_21120);
nand UO_501 (O_501,N_23083,N_22764);
nand UO_502 (O_502,N_24232,N_23578);
xor UO_503 (O_503,N_21292,N_24670);
or UO_504 (O_504,N_20012,N_23091);
or UO_505 (O_505,N_24532,N_20993);
and UO_506 (O_506,N_24104,N_20998);
nand UO_507 (O_507,N_24822,N_22429);
nor UO_508 (O_508,N_22940,N_21490);
or UO_509 (O_509,N_20464,N_21597);
and UO_510 (O_510,N_24954,N_22119);
and UO_511 (O_511,N_23344,N_21088);
or UO_512 (O_512,N_20188,N_21197);
or UO_513 (O_513,N_21692,N_22042);
xnor UO_514 (O_514,N_20792,N_20972);
xor UO_515 (O_515,N_23399,N_23249);
nand UO_516 (O_516,N_20838,N_21320);
nor UO_517 (O_517,N_24928,N_21546);
and UO_518 (O_518,N_22312,N_22388);
and UO_519 (O_519,N_24307,N_24496);
xor UO_520 (O_520,N_20145,N_22949);
or UO_521 (O_521,N_22669,N_20515);
and UO_522 (O_522,N_20742,N_21888);
nand UO_523 (O_523,N_20887,N_20171);
and UO_524 (O_524,N_21201,N_21239);
nor UO_525 (O_525,N_24553,N_24410);
xor UO_526 (O_526,N_24154,N_22128);
and UO_527 (O_527,N_23502,N_22052);
and UO_528 (O_528,N_22302,N_21867);
nor UO_529 (O_529,N_22022,N_23451);
nand UO_530 (O_530,N_21090,N_21157);
nand UO_531 (O_531,N_24497,N_23021);
and UO_532 (O_532,N_22380,N_23650);
or UO_533 (O_533,N_23581,N_23130);
and UO_534 (O_534,N_23382,N_24480);
nand UO_535 (O_535,N_23384,N_23985);
nor UO_536 (O_536,N_23971,N_23524);
xor UO_537 (O_537,N_20234,N_22043);
or UO_538 (O_538,N_24861,N_20065);
and UO_539 (O_539,N_20830,N_23745);
nand UO_540 (O_540,N_22551,N_21882);
nand UO_541 (O_541,N_24968,N_24406);
and UO_542 (O_542,N_22483,N_20825);
and UO_543 (O_543,N_23515,N_22735);
or UO_544 (O_544,N_22942,N_22485);
or UO_545 (O_545,N_23568,N_23475);
xnor UO_546 (O_546,N_21021,N_20455);
nor UO_547 (O_547,N_21551,N_21364);
xnor UO_548 (O_548,N_24133,N_24493);
nor UO_549 (O_549,N_20138,N_23867);
xnor UO_550 (O_550,N_21396,N_24262);
nand UO_551 (O_551,N_20384,N_21191);
and UO_552 (O_552,N_22714,N_23441);
or UO_553 (O_553,N_21436,N_21791);
and UO_554 (O_554,N_20116,N_24192);
nand UO_555 (O_555,N_21433,N_20211);
and UO_556 (O_556,N_21291,N_20661);
nand UO_557 (O_557,N_21644,N_21703);
nand UO_558 (O_558,N_20089,N_20580);
nor UO_559 (O_559,N_23076,N_21964);
nand UO_560 (O_560,N_22521,N_23887);
and UO_561 (O_561,N_22707,N_24890);
nand UO_562 (O_562,N_24999,N_22783);
or UO_563 (O_563,N_22775,N_24159);
xor UO_564 (O_564,N_22207,N_20617);
or UO_565 (O_565,N_24761,N_24110);
nand UO_566 (O_566,N_21889,N_24797);
nand UO_567 (O_567,N_20236,N_23327);
nand UO_568 (O_568,N_22987,N_22849);
nand UO_569 (O_569,N_20280,N_24782);
nand UO_570 (O_570,N_24277,N_21098);
xor UO_571 (O_571,N_23264,N_23287);
nor UO_572 (O_572,N_22497,N_22008);
nand UO_573 (O_573,N_23285,N_20377);
or UO_574 (O_574,N_23599,N_21249);
or UO_575 (O_575,N_23064,N_24253);
xnor UO_576 (O_576,N_20593,N_24857);
or UO_577 (O_577,N_21891,N_23546);
or UO_578 (O_578,N_20795,N_24297);
nor UO_579 (O_579,N_23579,N_22701);
nor UO_580 (O_580,N_20623,N_21973);
or UO_581 (O_581,N_23615,N_21234);
nand UO_582 (O_582,N_24250,N_24108);
xor UO_583 (O_583,N_24763,N_23610);
xor UO_584 (O_584,N_23699,N_23274);
nand UO_585 (O_585,N_20706,N_23442);
xnor UO_586 (O_586,N_24498,N_24750);
xor UO_587 (O_587,N_23602,N_22861);
xnor UO_588 (O_588,N_20353,N_24829);
xor UO_589 (O_589,N_22237,N_22943);
and UO_590 (O_590,N_23912,N_22153);
xor UO_591 (O_591,N_22925,N_22797);
xor UO_592 (O_592,N_20810,N_24736);
nand UO_593 (O_593,N_21919,N_24605);
or UO_594 (O_594,N_20646,N_21586);
nand UO_595 (O_595,N_20082,N_24944);
and UO_596 (O_596,N_24527,N_21575);
and UO_597 (O_597,N_24070,N_22970);
and UO_598 (O_598,N_21497,N_22698);
or UO_599 (O_599,N_24881,N_24432);
or UO_600 (O_600,N_24888,N_20447);
or UO_601 (O_601,N_24456,N_22097);
or UO_602 (O_602,N_20128,N_24296);
or UO_603 (O_603,N_24206,N_20255);
and UO_604 (O_604,N_24757,N_20929);
nor UO_605 (O_605,N_21303,N_21818);
nand UO_606 (O_606,N_22827,N_21220);
and UO_607 (O_607,N_21189,N_21602);
nand UO_608 (O_608,N_22763,N_21803);
nor UO_609 (O_609,N_23618,N_21666);
or UO_610 (O_610,N_22475,N_21345);
nand UO_611 (O_611,N_24508,N_21231);
nand UO_612 (O_612,N_23567,N_24798);
nor UO_613 (O_613,N_21135,N_24549);
nor UO_614 (O_614,N_21639,N_23095);
nor UO_615 (O_615,N_21915,N_24976);
or UO_616 (O_616,N_20572,N_20982);
and UO_617 (O_617,N_22845,N_20434);
or UO_618 (O_618,N_22807,N_23317);
and UO_619 (O_619,N_21811,N_21060);
nor UO_620 (O_620,N_20662,N_23102);
and UO_621 (O_621,N_21226,N_20849);
nor UO_622 (O_622,N_20913,N_21816);
nor UO_623 (O_623,N_23347,N_22006);
xnor UO_624 (O_624,N_22678,N_23660);
nand UO_625 (O_625,N_22904,N_23509);
and UO_626 (O_626,N_22231,N_22069);
nand UO_627 (O_627,N_20740,N_20357);
and UO_628 (O_628,N_22335,N_20076);
and UO_629 (O_629,N_22572,N_23722);
or UO_630 (O_630,N_23461,N_21064);
or UO_631 (O_631,N_20577,N_23129);
xor UO_632 (O_632,N_22325,N_22928);
nand UO_633 (O_633,N_24063,N_22741);
xor UO_634 (O_634,N_21605,N_20179);
nor UO_635 (O_635,N_24180,N_22150);
or UO_636 (O_636,N_24746,N_23046);
or UO_637 (O_637,N_24486,N_21407);
xnor UO_638 (O_638,N_24819,N_21071);
xor UO_639 (O_639,N_24917,N_20373);
nand UO_640 (O_640,N_22600,N_21431);
or UO_641 (O_641,N_23187,N_20264);
or UO_642 (O_642,N_21395,N_24424);
xor UO_643 (O_643,N_23279,N_21560);
xor UO_644 (O_644,N_23496,N_22654);
xor UO_645 (O_645,N_20797,N_21080);
xor UO_646 (O_646,N_23367,N_21289);
or UO_647 (O_647,N_22426,N_24593);
and UO_648 (O_648,N_22131,N_23589);
and UO_649 (O_649,N_23793,N_22254);
and UO_650 (O_650,N_23671,N_23418);
nand UO_651 (O_651,N_24401,N_22323);
nand UO_652 (O_652,N_20340,N_24030);
and UO_653 (O_653,N_21693,N_23149);
or UO_654 (O_654,N_24249,N_24940);
and UO_655 (O_655,N_23948,N_24038);
nand UO_656 (O_656,N_21584,N_21103);
nor UO_657 (O_657,N_22793,N_21011);
and UO_658 (O_658,N_23481,N_23683);
nand UO_659 (O_659,N_22068,N_23354);
or UO_660 (O_660,N_21773,N_23944);
and UO_661 (O_661,N_22005,N_21858);
nand UO_662 (O_662,N_20135,N_22657);
nor UO_663 (O_663,N_24741,N_23208);
nand UO_664 (O_664,N_20609,N_20085);
xor UO_665 (O_665,N_23309,N_21102);
xnor UO_666 (O_666,N_20008,N_20419);
nand UO_667 (O_667,N_23067,N_20992);
nand UO_668 (O_668,N_23229,N_24141);
and UO_669 (O_669,N_22820,N_22090);
nand UO_670 (O_670,N_24257,N_23959);
xor UO_671 (O_671,N_24209,N_21897);
xor UO_672 (O_672,N_23304,N_21893);
or UO_673 (O_673,N_21066,N_22361);
nor UO_674 (O_674,N_23633,N_20276);
nor UO_675 (O_675,N_21184,N_24204);
nor UO_676 (O_676,N_22095,N_24610);
xor UO_677 (O_677,N_20607,N_23086);
nand UO_678 (O_678,N_21255,N_24885);
nand UO_679 (O_679,N_20850,N_20327);
xor UO_680 (O_680,N_24584,N_21732);
and UO_681 (O_681,N_20477,N_22638);
nor UO_682 (O_682,N_20164,N_21108);
or UO_683 (O_683,N_22739,N_21093);
xnor UO_684 (O_684,N_22901,N_21376);
nand UO_685 (O_685,N_20508,N_21432);
nand UO_686 (O_686,N_23038,N_20087);
and UO_687 (O_687,N_21710,N_22048);
xnor UO_688 (O_688,N_22085,N_20938);
xor UO_689 (O_689,N_23528,N_24837);
or UO_690 (O_690,N_24491,N_23198);
and UO_691 (O_691,N_23169,N_21701);
or UO_692 (O_692,N_22384,N_21256);
xnor UO_693 (O_693,N_21192,N_21110);
and UO_694 (O_694,N_22319,N_21147);
nor UO_695 (O_695,N_23416,N_21125);
and UO_696 (O_696,N_21743,N_20769);
and UO_697 (O_697,N_20106,N_23397);
xor UO_698 (O_698,N_24567,N_21488);
nand UO_699 (O_699,N_23413,N_24265);
xnor UO_700 (O_700,N_22628,N_24305);
and UO_701 (O_701,N_24437,N_22806);
nor UO_702 (O_702,N_21491,N_23379);
and UO_703 (O_703,N_22369,N_22568);
and UO_704 (O_704,N_21061,N_22349);
nand UO_705 (O_705,N_24472,N_22286);
nor UO_706 (O_706,N_23010,N_22428);
xor UO_707 (O_707,N_20879,N_22712);
or UO_708 (O_708,N_23205,N_22765);
or UO_709 (O_709,N_21912,N_21878);
xnor UO_710 (O_710,N_22825,N_24753);
xnor UO_711 (O_711,N_22204,N_20209);
xor UO_712 (O_712,N_22198,N_23494);
or UO_713 (O_713,N_20594,N_21260);
and UO_714 (O_714,N_24194,N_22663);
nor UO_715 (O_715,N_21494,N_22951);
nand UO_716 (O_716,N_23588,N_23122);
and UO_717 (O_717,N_22383,N_21143);
nor UO_718 (O_718,N_22444,N_22740);
nor UO_719 (O_719,N_23718,N_21172);
nand UO_720 (O_720,N_20472,N_20704);
xor UO_721 (O_721,N_21160,N_20025);
xor UO_722 (O_722,N_24839,N_24412);
nor UO_723 (O_723,N_20759,N_22245);
and UO_724 (O_724,N_21977,N_22559);
xor UO_725 (O_725,N_22016,N_22421);
or UO_726 (O_726,N_23051,N_20865);
nor UO_727 (O_727,N_20063,N_24637);
xor UO_728 (O_728,N_20241,N_23679);
or UO_729 (O_729,N_21905,N_22699);
xnor UO_730 (O_730,N_22274,N_23863);
or UO_731 (O_731,N_21548,N_22787);
or UO_732 (O_732,N_24123,N_22496);
nor UO_733 (O_733,N_21046,N_22993);
nand UO_734 (O_734,N_21578,N_21922);
nor UO_735 (O_735,N_22974,N_21986);
nand UO_736 (O_736,N_22174,N_21372);
nor UO_737 (O_737,N_21966,N_22938);
nand UO_738 (O_738,N_21687,N_24374);
nor UO_739 (O_739,N_23482,N_24938);
or UO_740 (O_740,N_22478,N_24871);
nand UO_741 (O_741,N_21048,N_24478);
or UO_742 (O_742,N_23646,N_21266);
nand UO_743 (O_743,N_20598,N_24413);
nor UO_744 (O_744,N_20155,N_22405);
or UO_745 (O_745,N_20334,N_22732);
xor UO_746 (O_746,N_24676,N_24832);
or UO_747 (O_747,N_23161,N_23801);
xnor UO_748 (O_748,N_20394,N_20019);
nand UO_749 (O_749,N_22733,N_20168);
or UO_750 (O_750,N_24382,N_21718);
or UO_751 (O_751,N_20080,N_22098);
nor UO_752 (O_752,N_20800,N_20223);
nor UO_753 (O_753,N_20761,N_20247);
xnor UO_754 (O_754,N_22647,N_20809);
nor UO_755 (O_755,N_24327,N_22067);
and UO_756 (O_756,N_23123,N_24536);
and UO_757 (O_757,N_20778,N_21675);
xnor UO_758 (O_758,N_22033,N_20411);
nand UO_759 (O_759,N_20189,N_20069);
and UO_760 (O_760,N_21321,N_20124);
nor UO_761 (O_761,N_24119,N_20512);
nor UO_762 (O_762,N_21023,N_22919);
and UO_763 (O_763,N_24114,N_22536);
or UO_764 (O_764,N_23995,N_20882);
nand UO_765 (O_765,N_20793,N_21940);
xnor UO_766 (O_766,N_24083,N_20805);
and UO_767 (O_767,N_23963,N_22539);
xnor UO_768 (O_768,N_20984,N_22075);
xnor UO_769 (O_769,N_20329,N_23701);
xor UO_770 (O_770,N_21983,N_20196);
nand UO_771 (O_771,N_20183,N_21013);
and UO_772 (O_772,N_22382,N_21329);
nor UO_773 (O_773,N_21611,N_24136);
nor UO_774 (O_774,N_23704,N_21847);
nand UO_775 (O_775,N_24531,N_24821);
nand UO_776 (O_776,N_24452,N_22157);
nor UO_777 (O_777,N_20068,N_20505);
and UO_778 (O_778,N_20043,N_23997);
xor UO_779 (O_779,N_21386,N_23213);
xnor UO_780 (O_780,N_22481,N_22688);
xor UO_781 (O_781,N_21817,N_24251);
and UO_782 (O_782,N_23990,N_24772);
or UO_783 (O_783,N_24431,N_21472);
nor UO_784 (O_784,N_24357,N_20922);
and UO_785 (O_785,N_22392,N_24011);
nor UO_786 (O_786,N_21814,N_20967);
nand UO_787 (O_787,N_20413,N_23142);
nor UO_788 (O_788,N_24448,N_20057);
nand UO_789 (O_789,N_24153,N_22830);
nand UO_790 (O_790,N_21561,N_22931);
or UO_791 (O_791,N_24985,N_23664);
xor UO_792 (O_792,N_23651,N_21318);
and UO_793 (O_793,N_23480,N_20691);
nor UO_794 (O_794,N_24639,N_22401);
nor UO_795 (O_795,N_22573,N_22748);
nand UO_796 (O_796,N_21620,N_22309);
nor UO_797 (O_797,N_23946,N_22532);
xor UO_798 (O_798,N_20728,N_23359);
nand UO_799 (O_799,N_24675,N_21771);
or UO_800 (O_800,N_20955,N_23419);
and UO_801 (O_801,N_21799,N_21542);
nand UO_802 (O_802,N_22364,N_24606);
nand UO_803 (O_803,N_24187,N_22079);
nor UO_804 (O_804,N_20216,N_21496);
or UO_805 (O_805,N_22822,N_23582);
or UO_806 (O_806,N_21059,N_21945);
xor UO_807 (O_807,N_24495,N_24434);
nand UO_808 (O_808,N_22404,N_22965);
xnor UO_809 (O_809,N_22867,N_23391);
or UO_810 (O_810,N_23228,N_22635);
and UO_811 (O_811,N_24815,N_22101);
nand UO_812 (O_812,N_24563,N_23401);
or UO_813 (O_813,N_20468,N_24770);
or UO_814 (O_814,N_24542,N_21470);
and UO_815 (O_815,N_21705,N_24858);
or UO_816 (O_816,N_23974,N_22435);
and UO_817 (O_817,N_21981,N_24414);
nand UO_818 (O_818,N_22056,N_22012);
xnor UO_819 (O_819,N_23315,N_21465);
and UO_820 (O_820,N_24371,N_22385);
nor UO_821 (O_821,N_24139,N_22665);
and UO_822 (O_822,N_20460,N_22346);
xnor UO_823 (O_823,N_23152,N_24975);
nand UO_824 (O_824,N_23510,N_21449);
or UO_825 (O_825,N_22994,N_22437);
or UO_826 (O_826,N_21603,N_21587);
and UO_827 (O_827,N_24375,N_24530);
and UO_828 (O_828,N_22623,N_24538);
and UO_829 (O_829,N_22127,N_22409);
nor UO_830 (O_830,N_23542,N_20763);
nand UO_831 (O_831,N_23943,N_22894);
nor UO_832 (O_832,N_24577,N_20496);
nor UO_833 (O_833,N_24565,N_23040);
or UO_834 (O_834,N_24356,N_23986);
or UO_835 (O_835,N_24962,N_22637);
and UO_836 (O_836,N_21917,N_21450);
xnor UO_837 (O_837,N_23018,N_23093);
xnor UO_838 (O_838,N_20569,N_21327);
nand UO_839 (O_839,N_22363,N_20202);
or UO_840 (O_840,N_22141,N_20919);
and UO_841 (O_841,N_22137,N_23094);
and UO_842 (O_842,N_21012,N_24462);
nand UO_843 (O_843,N_22467,N_22768);
nor UO_844 (O_844,N_22556,N_23435);
nand UO_845 (O_845,N_21113,N_24699);
nor UO_846 (O_846,N_22252,N_23818);
and UO_847 (O_847,N_23532,N_20841);
nor UO_848 (O_848,N_22513,N_20430);
or UO_849 (O_849,N_23914,N_22929);
nor UO_850 (O_850,N_24308,N_22184);
and UO_851 (O_851,N_24636,N_20949);
nor UO_852 (O_852,N_22656,N_21338);
and UO_853 (O_853,N_21282,N_23019);
and UO_854 (O_854,N_21363,N_20735);
nor UO_855 (O_855,N_20952,N_23982);
nand UO_856 (O_856,N_23641,N_21043);
nor UO_857 (O_857,N_20448,N_20487);
nor UO_858 (O_858,N_21018,N_21749);
or UO_859 (O_859,N_22523,N_23117);
nor UO_860 (O_860,N_22181,N_20283);
xor UO_861 (O_861,N_24849,N_24591);
nor UO_862 (O_862,N_22905,N_22587);
and UO_863 (O_863,N_22594,N_20818);
or UO_864 (O_864,N_21939,N_21086);
nor UO_865 (O_865,N_21906,N_22358);
nand UO_866 (O_866,N_23409,N_21924);
nand UO_867 (O_867,N_23941,N_20220);
nor UO_868 (O_868,N_20647,N_23980);
or UO_869 (O_869,N_21961,N_22332);
xnor UO_870 (O_870,N_20245,N_23563);
nand UO_871 (O_871,N_20490,N_20393);
nand UO_872 (O_872,N_22934,N_24487);
and UO_873 (O_873,N_23276,N_21648);
nor UO_874 (O_874,N_21567,N_23896);
nand UO_875 (O_875,N_22015,N_20671);
and UO_876 (O_876,N_24510,N_21105);
nand UO_877 (O_877,N_21100,N_24229);
or UO_878 (O_878,N_23410,N_22218);
or UO_879 (O_879,N_23523,N_23924);
nor UO_880 (O_880,N_22365,N_20999);
and UO_881 (O_881,N_22911,N_23616);
and UO_882 (O_882,N_24345,N_22215);
and UO_883 (O_883,N_23159,N_24851);
and UO_884 (O_884,N_23240,N_20308);
xor UO_885 (O_885,N_24590,N_23113);
and UO_886 (O_886,N_21227,N_21132);
or UO_887 (O_887,N_23324,N_23207);
xor UO_888 (O_888,N_22221,N_22794);
nand UO_889 (O_889,N_20756,N_24704);
nor UO_890 (O_890,N_20205,N_20456);
or UO_891 (O_891,N_23190,N_20532);
and UO_892 (O_892,N_24989,N_20709);
nor UO_893 (O_893,N_21631,N_23574);
nor UO_894 (O_894,N_23262,N_21015);
xnor UO_895 (O_895,N_22799,N_20544);
xnor UO_896 (O_896,N_24631,N_23307);
or UO_897 (O_897,N_20366,N_20256);
or UO_898 (O_898,N_20062,N_20495);
nor UO_899 (O_899,N_21445,N_20554);
or UO_900 (O_900,N_22713,N_21872);
nand UO_901 (O_901,N_21169,N_24246);
nand UO_902 (O_902,N_24008,N_20452);
nand UO_903 (O_903,N_20804,N_22272);
nor UO_904 (O_904,N_24846,N_22874);
xor UO_905 (O_905,N_23141,N_23118);
nor UO_906 (O_906,N_24649,N_22727);
and UO_907 (O_907,N_22693,N_20557);
or UO_908 (O_908,N_21757,N_24394);
xor UO_909 (O_909,N_20870,N_24749);
nand UO_910 (O_910,N_22322,N_21840);
nor UO_911 (O_911,N_23903,N_23569);
nor UO_912 (O_912,N_24600,N_20212);
xnor UO_913 (O_913,N_21414,N_21862);
nand UO_914 (O_914,N_21461,N_20558);
and UO_915 (O_915,N_22990,N_21050);
xnor UO_916 (O_916,N_23846,N_23869);
xnor UO_917 (O_917,N_24714,N_22947);
xor UO_918 (O_918,N_20618,N_21659);
nand UO_919 (O_919,N_24706,N_23048);
nand UO_920 (O_920,N_24854,N_23146);
nand UO_921 (O_921,N_22966,N_23691);
nor UO_922 (O_922,N_21716,N_22142);
or UO_923 (O_923,N_21350,N_22815);
nor UO_924 (O_924,N_23861,N_23829);
nand UO_925 (O_925,N_21600,N_23521);
or UO_926 (O_926,N_21649,N_24751);
or UO_927 (O_927,N_23437,N_23711);
or UO_928 (O_928,N_20401,N_21005);
and UO_929 (O_929,N_23312,N_20392);
nand UO_930 (O_930,N_21275,N_22004);
nand UO_931 (O_931,N_22618,N_21418);
and UO_932 (O_932,N_21806,N_22381);
nor UO_933 (O_933,N_21107,N_21351);
or UO_934 (O_934,N_21290,N_20961);
or UO_935 (O_935,N_23029,N_22230);
nand UO_936 (O_936,N_22685,N_23603);
xnor UO_937 (O_937,N_21190,N_22643);
nor UO_938 (O_938,N_22412,N_21744);
or UO_939 (O_939,N_21804,N_20178);
xnor UO_940 (O_940,N_22490,N_23305);
nor UO_941 (O_941,N_21527,N_23199);
nand UO_942 (O_942,N_24223,N_21114);
and UO_943 (O_943,N_21175,N_21267);
xnor UO_944 (O_944,N_21258,N_24198);
or UO_945 (O_945,N_22178,N_20173);
or UO_946 (O_946,N_21020,N_20684);
nor UO_947 (O_947,N_23939,N_24103);
nand UO_948 (O_948,N_20310,N_23353);
or UO_949 (O_949,N_21671,N_21808);
xor UO_950 (O_950,N_20507,N_22531);
and UO_951 (O_951,N_20540,N_22750);
and UO_952 (O_952,N_20350,N_20197);
or UO_953 (O_953,N_22718,N_21507);
xnor UO_954 (O_954,N_23810,N_22730);
nand UO_955 (O_955,N_20314,N_21741);
xor UO_956 (O_956,N_20864,N_22542);
or UO_957 (O_957,N_22280,N_20258);
nor UO_958 (O_958,N_21899,N_20151);
nor UO_959 (O_959,N_23871,N_24679);
xnor UO_960 (O_960,N_23835,N_20500);
nand UO_961 (O_961,N_24731,N_20290);
nand UO_962 (O_962,N_23740,N_22906);
and UO_963 (O_963,N_20288,N_22864);
nor UO_964 (O_964,N_24399,N_20266);
and UO_965 (O_965,N_21835,N_23231);
xnor UO_966 (O_966,N_24391,N_21934);
or UO_967 (O_967,N_23491,N_20616);
nor UO_968 (O_968,N_23681,N_24354);
nand UO_969 (O_969,N_23970,N_23452);
and UO_970 (O_970,N_21936,N_23368);
nand UO_971 (O_971,N_23994,N_24937);
xor UO_972 (O_972,N_21041,N_23716);
nand UO_973 (O_973,N_20462,N_23492);
or UO_974 (O_974,N_23158,N_21729);
or UO_975 (O_975,N_20962,N_21403);
nor UO_976 (O_976,N_20597,N_22210);
nor UO_977 (O_977,N_22737,N_23687);
nand UO_978 (O_978,N_21860,N_20478);
nor UO_979 (O_979,N_20267,N_22114);
or UO_980 (O_980,N_23960,N_23955);
or UO_981 (O_981,N_24045,N_22650);
nand UO_982 (O_982,N_20286,N_24271);
and UO_983 (O_983,N_20638,N_23449);
nor UO_984 (O_984,N_23551,N_22482);
or UO_985 (O_985,N_22253,N_23662);
nor UO_986 (O_986,N_22675,N_24868);
and UO_987 (O_987,N_23031,N_23258);
nand UO_988 (O_988,N_20932,N_24331);
nor UO_989 (O_989,N_22968,N_24923);
and UO_990 (O_990,N_21826,N_24934);
and UO_991 (O_991,N_23280,N_22914);
and UO_992 (O_992,N_23242,N_24719);
or UO_993 (O_993,N_23292,N_21884);
xnor UO_994 (O_994,N_22791,N_20912);
or UO_995 (O_995,N_23968,N_24301);
xnor UO_996 (O_996,N_23465,N_21389);
nor UO_997 (O_997,N_20103,N_21424);
and UO_998 (O_998,N_22399,N_24887);
or UO_999 (O_999,N_21619,N_20282);
or UO_1000 (O_1000,N_20127,N_22356);
or UO_1001 (O_1001,N_23680,N_23273);
xnor UO_1002 (O_1002,N_21342,N_22213);
nand UO_1003 (O_1003,N_24292,N_21308);
or UO_1004 (O_1004,N_21821,N_21667);
or UO_1005 (O_1005,N_22062,N_21417);
nor UO_1006 (O_1006,N_22725,N_21096);
or UO_1007 (O_1007,N_22687,N_22575);
nand UO_1008 (O_1008,N_24411,N_20023);
nand UO_1009 (O_1009,N_23689,N_20092);
nor UO_1010 (O_1010,N_21746,N_20905);
nand UO_1011 (O_1011,N_21460,N_24625);
nand UO_1012 (O_1012,N_23405,N_23607);
or UO_1013 (O_1013,N_20125,N_21534);
nand UO_1014 (O_1014,N_22771,N_20299);
and UO_1015 (O_1015,N_22686,N_21448);
xor UO_1016 (O_1016,N_24442,N_20254);
and UO_1017 (O_1017,N_24258,N_21740);
and UO_1018 (O_1018,N_22537,N_23110);
or UO_1019 (O_1019,N_23741,N_22939);
nor UO_1020 (O_1020,N_21394,N_23746);
and UO_1021 (O_1021,N_22616,N_23760);
xnor UO_1022 (O_1022,N_22452,N_24948);
nor UO_1023 (O_1023,N_23001,N_21819);
xor UO_1024 (O_1024,N_23443,N_21346);
nor UO_1025 (O_1025,N_24003,N_20875);
xnor UO_1026 (O_1026,N_24525,N_21769);
nand UO_1027 (O_1027,N_24470,N_21262);
and UO_1028 (O_1028,N_21040,N_21730);
nand UO_1029 (O_1029,N_24874,N_21035);
or UO_1030 (O_1030,N_20222,N_21242);
xor UO_1031 (O_1031,N_20118,N_20894);
nor UO_1032 (O_1032,N_20154,N_24488);
xor UO_1033 (O_1033,N_20166,N_21153);
or UO_1034 (O_1034,N_21152,N_22423);
nor UO_1035 (O_1035,N_23604,N_21850);
xnor UO_1036 (O_1036,N_20801,N_24796);
nor UO_1037 (O_1037,N_24612,N_20354);
nor UO_1038 (O_1038,N_23423,N_21206);
and UO_1039 (O_1039,N_23571,N_24995);
and UO_1040 (O_1040,N_24642,N_21469);
nand UO_1041 (O_1041,N_22662,N_23462);
or UO_1042 (O_1042,N_22726,N_23253);
nand UO_1043 (O_1043,N_22977,N_24161);
or UO_1044 (O_1044,N_23761,N_21928);
nor UO_1045 (O_1045,N_21537,N_23172);
or UO_1046 (O_1046,N_22789,N_23684);
nor UO_1047 (O_1047,N_24384,N_21067);
nor UO_1048 (O_1048,N_24570,N_20817);
nand UO_1049 (O_1049,N_24855,N_20372);
or UO_1050 (O_1050,N_20854,N_23070);
nor UO_1051 (O_1051,N_23140,N_22852);
or UO_1052 (O_1052,N_24235,N_22070);
or UO_1053 (O_1053,N_21218,N_23039);
or UO_1054 (O_1054,N_21397,N_24302);
nand UO_1055 (O_1055,N_22530,N_20980);
nand UO_1056 (O_1056,N_23520,N_23457);
nand UO_1057 (O_1057,N_24655,N_20317);
and UO_1058 (O_1058,N_20665,N_23294);
and UO_1059 (O_1059,N_21529,N_21678);
and UO_1060 (O_1060,N_24820,N_21039);
xnor UO_1061 (O_1061,N_21141,N_23250);
xnor UO_1062 (O_1062,N_24310,N_23180);
xnor UO_1063 (O_1063,N_23940,N_22903);
or UO_1064 (O_1064,N_23100,N_22747);
nor UO_1065 (O_1065,N_24077,N_22088);
or UO_1066 (O_1066,N_21252,N_20666);
or UO_1067 (O_1067,N_20606,N_21466);
nor UO_1068 (O_1068,N_23310,N_20766);
nor UO_1069 (O_1069,N_21058,N_23725);
nand UO_1070 (O_1070,N_23972,N_22256);
xor UO_1071 (O_1071,N_24023,N_20956);
and UO_1072 (O_1072,N_24713,N_22287);
or UO_1073 (O_1073,N_24793,N_21938);
xor UO_1074 (O_1074,N_23270,N_21623);
nor UO_1075 (O_1075,N_24733,N_21579);
nor UO_1076 (O_1076,N_22108,N_20341);
and UO_1077 (O_1077,N_20548,N_23575);
xor UO_1078 (O_1078,N_22625,N_20583);
nor UO_1079 (O_1079,N_23900,N_24197);
xor UO_1080 (O_1080,N_21000,N_21503);
and UO_1081 (O_1081,N_20531,N_23719);
nand UO_1082 (O_1082,N_22742,N_20039);
or UO_1083 (O_1083,N_20931,N_20588);
and UO_1084 (O_1084,N_21929,N_23084);
nand UO_1085 (O_1085,N_23092,N_20614);
or UO_1086 (O_1086,N_23026,N_24020);
or UO_1087 (O_1087,N_24347,N_20421);
xor UO_1088 (O_1088,N_22753,N_22311);
xor UO_1089 (O_1089,N_21911,N_24380);
nor UO_1090 (O_1090,N_21443,N_22172);
or UO_1091 (O_1091,N_24492,N_21233);
nor UO_1092 (O_1092,N_22136,N_24479);
nor UO_1093 (O_1093,N_24927,N_20529);
or UO_1094 (O_1094,N_23013,N_20856);
xor UO_1095 (O_1095,N_21967,N_22244);
nand UO_1096 (O_1096,N_24853,N_24514);
nand UO_1097 (O_1097,N_20871,N_22890);
nand UO_1098 (O_1098,N_22767,N_24897);
nor UO_1099 (O_1099,N_23707,N_21047);
xor UO_1100 (O_1100,N_24033,N_20659);
nand UO_1101 (O_1101,N_21877,N_21612);
xor UO_1102 (O_1102,N_21111,N_23230);
and UO_1103 (O_1103,N_24035,N_22275);
and UO_1104 (O_1104,N_24807,N_21429);
or UO_1105 (O_1105,N_23888,N_22711);
nand UO_1106 (O_1106,N_22199,N_24069);
and UO_1107 (O_1107,N_20198,N_22223);
and UO_1108 (O_1108,N_21770,N_21406);
xor UO_1109 (O_1109,N_21844,N_23795);
xor UO_1110 (O_1110,N_23296,N_24474);
nor UO_1111 (O_1111,N_20802,N_21082);
and UO_1112 (O_1112,N_21240,N_22395);
nand UO_1113 (O_1113,N_22589,N_21323);
xnor UO_1114 (O_1114,N_22203,N_20679);
nor UO_1115 (O_1115,N_22259,N_23729);
nor UO_1116 (O_1116,N_24688,N_21285);
or UO_1117 (O_1117,N_23016,N_21657);
and UO_1118 (O_1118,N_23162,N_23606);
nand UO_1119 (O_1119,N_21694,N_22517);
nor UO_1120 (O_1120,N_21054,N_24386);
and UO_1121 (O_1121,N_24276,N_20915);
nand UO_1122 (O_1122,N_21306,N_21230);
or UO_1123 (O_1123,N_20386,N_21999);
nor UO_1124 (O_1124,N_23248,N_24450);
xnor UO_1125 (O_1125,N_24951,N_24633);
nand UO_1126 (O_1126,N_22476,N_23005);
nand UO_1127 (O_1127,N_23906,N_24072);
nor UO_1128 (O_1128,N_20853,N_21975);
nand UO_1129 (O_1129,N_24149,N_24528);
or UO_1130 (O_1130,N_22411,N_22578);
and UO_1131 (O_1131,N_21232,N_23698);
or UO_1132 (O_1132,N_23252,N_21640);
nand UO_1133 (O_1133,N_24526,N_20000);
nor UO_1134 (O_1134,N_21273,N_21008);
nor UO_1135 (O_1135,N_20292,N_23775);
and UO_1136 (O_1136,N_21019,N_20342);
nand UO_1137 (O_1137,N_22973,N_23548);
or UO_1138 (O_1138,N_22891,N_22340);
or UO_1139 (O_1139,N_22169,N_23737);
nor UO_1140 (O_1140,N_21880,N_20552);
nor UO_1141 (O_1141,N_24728,N_24010);
xnor UO_1142 (O_1142,N_21400,N_21440);
nor UO_1143 (O_1143,N_24980,N_21412);
nor UO_1144 (O_1144,N_23197,N_24409);
and UO_1145 (O_1145,N_24875,N_20649);
nand UO_1146 (O_1146,N_24196,N_23440);
nand UO_1147 (O_1147,N_21870,N_21780);
nor UO_1148 (O_1148,N_22233,N_24126);
nand UO_1149 (O_1149,N_22488,N_22462);
xnor UO_1150 (O_1150,N_24964,N_20592);
nor UO_1151 (O_1151,N_24552,N_22924);
xor UO_1152 (O_1152,N_21790,N_23872);
nand UO_1153 (O_1153,N_22538,N_21138);
or UO_1154 (O_1154,N_24018,N_20498);
nor UO_1155 (O_1155,N_23350,N_21533);
and UO_1156 (O_1156,N_20848,N_20006);
nor UO_1157 (O_1157,N_23023,N_21843);
and UO_1158 (O_1158,N_20181,N_21691);
xor UO_1159 (O_1159,N_24170,N_24397);
nor UO_1160 (O_1160,N_22130,N_24959);
and UO_1161 (O_1161,N_23017,N_22484);
nand UO_1162 (O_1162,N_23738,N_23490);
nand UO_1163 (O_1163,N_23951,N_20738);
or UO_1164 (O_1164,N_22326,N_23865);
nand UO_1165 (O_1165,N_23695,N_22932);
or UO_1166 (O_1166,N_22376,N_23714);
nand UO_1167 (O_1167,N_24840,N_22935);
nor UO_1168 (O_1168,N_22138,N_23259);
nand UO_1169 (O_1169,N_20934,N_21167);
nor UO_1170 (O_1170,N_24321,N_24381);
xnor UO_1171 (O_1171,N_20969,N_24464);
xor UO_1172 (O_1172,N_21665,N_22433);
and UO_1173 (O_1173,N_21385,N_23648);
nor UO_1174 (O_1174,N_21828,N_24901);
and UO_1175 (O_1175,N_23446,N_24700);
xnor UO_1176 (O_1176,N_23855,N_23365);
and UO_1177 (O_1177,N_22425,N_22465);
or UO_1178 (O_1178,N_24075,N_24076);
xnor UO_1179 (O_1179,N_20503,N_20261);
or UO_1180 (O_1180,N_23854,N_22553);
nand UO_1181 (O_1181,N_21997,N_24416);
xor UO_1182 (O_1182,N_22045,N_21596);
nand UO_1183 (O_1183,N_22187,N_20333);
or UO_1184 (O_1184,N_21148,N_20387);
or UO_1185 (O_1185,N_21334,N_24604);
xor UO_1186 (O_1186,N_20140,N_21365);
or UO_1187 (O_1187,N_21062,N_20860);
and UO_1188 (O_1188,N_21697,N_20371);
or UO_1189 (O_1189,N_22988,N_24315);
nand UO_1190 (O_1190,N_24002,N_21615);
xor UO_1191 (O_1191,N_24611,N_21916);
nor UO_1192 (O_1192,N_23366,N_21613);
xnor UO_1193 (O_1193,N_24971,N_21042);
and UO_1194 (O_1194,N_20716,N_22784);
or UO_1195 (O_1195,N_23965,N_24626);
nor UO_1196 (O_1196,N_20937,N_23945);
nor UO_1197 (O_1197,N_24755,N_21037);
nand UO_1198 (O_1198,N_22235,N_22689);
or UO_1199 (O_1199,N_20449,N_21876);
nand UO_1200 (O_1200,N_24256,N_22242);
nand UO_1201 (O_1201,N_20823,N_22061);
nor UO_1202 (O_1202,N_22018,N_24547);
and UO_1203 (O_1203,N_21753,N_20859);
nand UO_1204 (O_1204,N_24512,N_23321);
nand UO_1205 (O_1205,N_24212,N_24014);
and UO_1206 (O_1206,N_20936,N_23621);
nor UO_1207 (O_1207,N_21987,N_21377);
nand UO_1208 (O_1208,N_20485,N_24270);
or UO_1209 (O_1209,N_23739,N_24280);
xnor UO_1210 (O_1210,N_21706,N_20585);
and UO_1211 (O_1211,N_20306,N_24287);
or UO_1212 (O_1212,N_22468,N_20323);
nand UO_1213 (O_1213,N_21591,N_23227);
xor UO_1214 (O_1214,N_22152,N_21393);
xnor UO_1215 (O_1215,N_20175,N_22023);
nand UO_1216 (O_1216,N_20018,N_23594);
xor UO_1217 (O_1217,N_23183,N_23562);
nand UO_1218 (O_1218,N_23788,N_24467);
nor UO_1219 (O_1219,N_23381,N_23445);
nand UO_1220 (O_1220,N_20639,N_22997);
and UO_1221 (O_1221,N_24843,N_24930);
or UO_1222 (O_1222,N_22569,N_24764);
or UO_1223 (O_1223,N_23806,N_21796);
xor UO_1224 (O_1224,N_21087,N_21229);
xor UO_1225 (O_1225,N_21733,N_24426);
and UO_1226 (O_1226,N_21092,N_21187);
nand UO_1227 (O_1227,N_20207,N_23081);
and UO_1228 (O_1228,N_20645,N_24560);
and UO_1229 (O_1229,N_21544,N_21247);
and UO_1230 (O_1230,N_24366,N_24459);
xnor UO_1231 (O_1231,N_23121,N_21634);
and UO_1232 (O_1232,N_23479,N_22584);
xor UO_1233 (O_1233,N_20872,N_23853);
xnor UO_1234 (O_1234,N_22224,N_24363);
nand UO_1235 (O_1235,N_20457,N_21193);
xor UO_1236 (O_1236,N_21370,N_22320);
xor UO_1237 (O_1237,N_22455,N_21482);
xor UO_1238 (O_1238,N_23139,N_24926);
nand UO_1239 (O_1239,N_22370,N_22373);
nor UO_1240 (O_1240,N_24346,N_22458);
nand UO_1241 (O_1241,N_22978,N_23363);
nor UO_1242 (O_1242,N_21702,N_23682);
xnor UO_1243 (O_1243,N_21250,N_20307);
or UO_1244 (O_1244,N_23389,N_23109);
nor UO_1245 (O_1245,N_22565,N_22731);
nor UO_1246 (O_1246,N_23499,N_21555);
and UO_1247 (O_1247,N_20159,N_24105);
and UO_1248 (O_1248,N_23357,N_23151);
and UO_1249 (O_1249,N_24678,N_23932);
or UO_1250 (O_1250,N_20184,N_22579);
xnor UO_1251 (O_1251,N_20737,N_20829);
and UO_1252 (O_1252,N_22011,N_24863);
xnor UO_1253 (O_1253,N_20933,N_20033);
nand UO_1254 (O_1254,N_21636,N_23268);
or UO_1255 (O_1255,N_24758,N_20935);
and UO_1256 (O_1256,N_23313,N_24664);
nor UO_1257 (O_1257,N_23177,N_23272);
or UO_1258 (O_1258,N_22866,N_22431);
nor UO_1259 (O_1259,N_21782,N_21215);
nor UO_1260 (O_1260,N_20560,N_21119);
xnor UO_1261 (O_1261,N_23215,N_23923);
nor UO_1262 (O_1262,N_20911,N_22420);
or UO_1263 (O_1263,N_23785,N_20093);
nand UO_1264 (O_1264,N_21868,N_22660);
or UO_1265 (O_1265,N_21670,N_22956);
xnor UO_1266 (O_1266,N_23814,N_23580);
and UO_1267 (O_1267,N_24513,N_23620);
nor UO_1268 (O_1268,N_22814,N_23489);
or UO_1269 (O_1269,N_21520,N_21759);
xor UO_1270 (O_1270,N_23916,N_24760);
or UO_1271 (O_1271,N_21478,N_22603);
and UO_1272 (O_1272,N_20814,N_24916);
and UO_1273 (O_1273,N_20400,N_24661);
xor UO_1274 (O_1274,N_23484,N_23408);
or UO_1275 (O_1275,N_20807,N_24652);
or UO_1276 (O_1276,N_21738,N_23962);
nand UO_1277 (O_1277,N_21655,N_22703);
nor UO_1278 (O_1278,N_21056,N_24884);
nor UO_1279 (O_1279,N_23075,N_21927);
or UO_1280 (O_1280,N_21638,N_23501);
and UO_1281 (O_1281,N_20773,N_23352);
and UO_1282 (O_1282,N_24784,N_23476);
nor UO_1283 (O_1283,N_20101,N_22180);
xnor UO_1284 (O_1284,N_20765,N_24268);
and UO_1285 (O_1285,N_22457,N_21150);
and UO_1286 (O_1286,N_20945,N_24579);
and UO_1287 (O_1287,N_23429,N_24523);
nor UO_1288 (O_1288,N_20193,N_22617);
nand UO_1289 (O_1289,N_20845,N_21387);
nand UO_1290 (O_1290,N_20526,N_22102);
and UO_1291 (O_1291,N_23300,N_20909);
nand UO_1292 (O_1292,N_23600,N_22297);
nor UO_1293 (O_1293,N_23014,N_20753);
xor UO_1294 (O_1294,N_21522,N_24801);
nand UO_1295 (O_1295,N_24720,N_20380);
nor UO_1296 (O_1296,N_22872,N_22955);
or UO_1297 (O_1297,N_21339,N_23723);
xor UO_1298 (O_1298,N_22746,N_20440);
nor UO_1299 (O_1299,N_23799,N_23882);
nor UO_1300 (O_1300,N_21748,N_23513);
nor UO_1301 (O_1301,N_21646,N_20296);
nor UO_1302 (O_1302,N_21991,N_21543);
nor UO_1303 (O_1303,N_23471,N_20294);
or UO_1304 (O_1304,N_20287,N_22151);
nand UO_1305 (O_1305,N_24349,N_24454);
nor UO_1306 (O_1306,N_24468,N_20869);
nand UO_1307 (O_1307,N_21772,N_20615);
nand UO_1308 (O_1308,N_22074,N_20796);
nand UO_1309 (O_1309,N_22117,N_24499);
or UO_1310 (O_1310,N_22343,N_22504);
xnor UO_1311 (O_1311,N_24993,N_21793);
xnor UO_1312 (O_1312,N_24648,N_20896);
nand UO_1313 (O_1313,N_20997,N_24398);
nor UO_1314 (O_1314,N_22209,N_24402);
nor UO_1315 (O_1315,N_21832,N_24572);
nand UO_1316 (O_1316,N_22447,N_23069);
and UO_1317 (O_1317,N_20702,N_23834);
xor UO_1318 (O_1318,N_21030,N_21593);
or UO_1319 (O_1319,N_21535,N_24859);
and UO_1320 (O_1320,N_23066,N_24245);
nand UO_1321 (O_1321,N_21117,N_21775);
nand UO_1322 (O_1322,N_20878,N_24775);
and UO_1323 (O_1323,N_20476,N_21960);
or UO_1324 (O_1324,N_24494,N_24586);
and UO_1325 (O_1325,N_22487,N_20946);
or UO_1326 (O_1326,N_22786,N_24420);
or UO_1327 (O_1327,N_22418,N_20926);
and UO_1328 (O_1328,N_21287,N_21831);
nand UO_1329 (O_1329,N_21155,N_21007);
nand UO_1330 (O_1330,N_24085,N_22886);
nor UO_1331 (O_1331,N_21688,N_24735);
or UO_1332 (O_1332,N_21516,N_22124);
or UO_1333 (O_1333,N_24983,N_23898);
nor UO_1334 (O_1334,N_24698,N_24660);
nand UO_1335 (O_1335,N_20504,N_22761);
or UO_1336 (O_1336,N_24387,N_20533);
nor UO_1337 (O_1337,N_20249,N_22099);
xor UO_1338 (O_1338,N_24622,N_23744);
nor UO_1339 (O_1339,N_24982,N_22777);
or UO_1340 (O_1340,N_21366,N_24306);
xor UO_1341 (O_1341,N_23796,N_24613);
or UO_1342 (O_1342,N_23145,N_22116);
nor UO_1343 (O_1343,N_23105,N_21972);
xor UO_1344 (O_1344,N_20423,N_21952);
nand UO_1345 (O_1345,N_23202,N_21462);
or UO_1346 (O_1346,N_21681,N_24898);
xor UO_1347 (O_1347,N_22239,N_22430);
nor UO_1348 (O_1348,N_20642,N_23780);
nand UO_1349 (O_1349,N_24683,N_23372);
and UO_1350 (O_1350,N_24866,N_20454);
nor UO_1351 (O_1351,N_23422,N_21944);
or UO_1352 (O_1352,N_21577,N_23815);
nor UO_1353 (O_1353,N_20194,N_23101);
nor UO_1354 (O_1354,N_20978,N_22170);
or UO_1355 (O_1355,N_23025,N_24316);
nor UO_1356 (O_1356,N_23261,N_24748);
and UO_1357 (O_1357,N_23686,N_24961);
and UO_1358 (O_1358,N_22039,N_22946);
or UO_1359 (O_1359,N_24602,N_22415);
nor UO_1360 (O_1360,N_24668,N_24789);
or UO_1361 (O_1361,N_22708,N_21302);
or UO_1362 (O_1362,N_23720,N_21747);
xnor UO_1363 (O_1363,N_23340,N_21356);
xnor UO_1364 (O_1364,N_22436,N_22964);
or UO_1365 (O_1365,N_24028,N_20502);
xnor UO_1366 (O_1366,N_23226,N_21207);
nand UO_1367 (O_1367,N_24157,N_23043);
xor UO_1368 (O_1368,N_24936,N_22880);
or UO_1369 (O_1369,N_20098,N_20042);
xnor UO_1370 (O_1370,N_21918,N_20619);
nand UO_1371 (O_1371,N_22695,N_22610);
nor UO_1372 (O_1372,N_22053,N_22084);
xor UO_1373 (O_1373,N_24647,N_20643);
xnor UO_1374 (O_1374,N_21829,N_22144);
nand UO_1375 (O_1375,N_22386,N_20768);
or UO_1376 (O_1376,N_24939,N_20032);
or UO_1377 (O_1377,N_23314,N_20318);
nand UO_1378 (O_1378,N_24969,N_22920);
and UO_1379 (O_1379,N_20699,N_22821);
xnor UO_1380 (O_1380,N_22021,N_24747);
and UO_1381 (O_1381,N_23210,N_24059);
nand UO_1382 (O_1382,N_22205,N_24680);
xor UO_1383 (O_1383,N_20243,N_22352);
nor UO_1384 (O_1384,N_23478,N_20275);
nor UO_1385 (O_1385,N_23056,N_20743);
and UO_1386 (O_1386,N_24548,N_20436);
nand UO_1387 (O_1387,N_22605,N_22869);
nor UO_1388 (O_1388,N_23167,N_20289);
and UO_1389 (O_1389,N_22110,N_23937);
nor UO_1390 (O_1390,N_23333,N_20509);
or UO_1391 (O_1391,N_24100,N_23111);
nand UO_1392 (O_1392,N_23540,N_20260);
and UO_1393 (O_1393,N_20149,N_20215);
xor UO_1394 (O_1394,N_23778,N_23179);
nor UO_1395 (O_1395,N_20908,N_22439);
xor UO_1396 (O_1396,N_22122,N_22516);
nor UO_1397 (O_1397,N_21752,N_21781);
or UO_1398 (O_1398,N_21180,N_24216);
nand UO_1399 (O_1399,N_23088,N_24595);
nor UO_1400 (O_1400,N_21149,N_22510);
or UO_1401 (O_1401,N_23244,N_24902);
or UO_1402 (O_1402,N_20831,N_24506);
or UO_1403 (O_1403,N_23511,N_23393);
and UO_1404 (O_1404,N_24026,N_23886);
or UO_1405 (O_1405,N_24185,N_20943);
and UO_1406 (O_1406,N_20100,N_24348);
nand UO_1407 (O_1407,N_24095,N_21842);
or UO_1408 (O_1408,N_22471,N_24667);
and UO_1409 (O_1409,N_22937,N_20595);
and UO_1410 (O_1410,N_20230,N_21676);
nand UO_1411 (O_1411,N_20263,N_22200);
and UO_1412 (O_1412,N_21477,N_20086);
xor UO_1413 (O_1413,N_22626,N_23901);
or UO_1414 (O_1414,N_20599,N_21536);
nor UO_1415 (O_1415,N_20108,N_22622);
and UO_1416 (O_1416,N_22486,N_20861);
xnor UO_1417 (O_1417,N_20633,N_23759);
or UO_1418 (O_1418,N_24248,N_22040);
xor UO_1419 (O_1419,N_21509,N_22255);
and UO_1420 (O_1420,N_23586,N_24834);
xnor UO_1421 (O_1421,N_22840,N_23004);
nor UO_1422 (O_1422,N_21188,N_20059);
and UO_1423 (O_1423,N_23640,N_22220);
xnor UO_1424 (O_1424,N_22087,N_24169);
nand UO_1425 (O_1425,N_23255,N_20536);
xor UO_1426 (O_1426,N_23809,N_20573);
or UO_1427 (O_1427,N_21489,N_20365);
nand UO_1428 (O_1428,N_20099,N_23859);
nor UO_1429 (O_1429,N_23755,N_20602);
nand UO_1430 (O_1430,N_20991,N_20047);
and UO_1431 (O_1431,N_20653,N_22534);
xor UO_1432 (O_1432,N_20914,N_22508);
nor UO_1433 (O_1433,N_21212,N_23238);
or UO_1434 (O_1434,N_20491,N_23774);
nor UO_1435 (O_1435,N_23427,N_20191);
xnor UO_1436 (O_1436,N_20109,N_22562);
nor UO_1437 (O_1437,N_23301,N_20497);
nor UO_1438 (O_1438,N_21129,N_24436);
nor UO_1439 (O_1439,N_24389,N_23374);
nor UO_1440 (O_1440,N_22145,N_20576);
or UO_1441 (O_1441,N_23852,N_24794);
nand UO_1442 (O_1442,N_22851,N_20433);
nor UO_1443 (O_1443,N_24669,N_22692);
or UO_1444 (O_1444,N_24116,N_24269);
nor UO_1445 (O_1445,N_23370,N_24872);
or UO_1446 (O_1446,N_23534,N_20158);
nor UO_1447 (O_1447,N_24893,N_21439);
xnor UO_1448 (O_1448,N_20520,N_23133);
xnor UO_1449 (O_1449,N_24918,N_20007);
nand UO_1450 (O_1450,N_22959,N_24403);
nand UO_1451 (O_1451,N_21069,N_20655);
nor UO_1452 (O_1452,N_23721,N_22479);
and UO_1453 (O_1453,N_24469,N_20586);
or UO_1454 (O_1454,N_21288,N_20794);
or UO_1455 (O_1455,N_21768,N_24324);
and UO_1456 (O_1456,N_21787,N_21257);
nor UO_1457 (O_1457,N_24017,N_20048);
nand UO_1458 (O_1458,N_24787,N_21427);
xnor UO_1459 (O_1459,N_21562,N_23486);
or UO_1460 (O_1460,N_22216,N_24298);
or UO_1461 (O_1461,N_20129,N_23953);
xor UO_1462 (O_1462,N_21511,N_21183);
nand UO_1463 (O_1463,N_21352,N_24650);
nand UO_1464 (O_1464,N_22509,N_20186);
nor UO_1465 (O_1465,N_20790,N_24360);
and UO_1466 (O_1466,N_23642,N_24653);
or UO_1467 (O_1467,N_20511,N_23931);
nor UO_1468 (O_1468,N_21569,N_22262);
xnor UO_1469 (O_1469,N_20874,N_24708);
or UO_1470 (O_1470,N_23171,N_24358);
nand UO_1471 (O_1471,N_20953,N_22446);
xnor UO_1472 (O_1472,N_24994,N_23087);
or UO_1473 (O_1473,N_21727,N_24972);
nand UO_1474 (O_1474,N_21901,N_23055);
nand UO_1475 (O_1475,N_22800,N_24694);
and UO_1476 (O_1476,N_23403,N_23282);
xnor UO_1477 (O_1477,N_22251,N_24051);
and UO_1478 (O_1478,N_23730,N_23920);
and UO_1479 (O_1479,N_23769,N_21177);
xnor UO_1480 (O_1480,N_22576,N_22734);
nor UO_1481 (O_1481,N_20005,N_23647);
nand UO_1482 (O_1482,N_20783,N_22586);
nand UO_1483 (O_1483,N_24101,N_20824);
and UO_1484 (O_1484,N_24880,N_22310);
xor UO_1485 (O_1485,N_20051,N_24048);
nor UO_1486 (O_1486,N_20564,N_23976);
nor UO_1487 (O_1487,N_20004,N_21709);
nand UO_1488 (O_1488,N_22063,N_21647);
nor UO_1489 (O_1489,N_24407,N_24024);
xnor UO_1490 (O_1490,N_24709,N_21890);
nand UO_1491 (O_1491,N_22400,N_20525);
xor UO_1492 (O_1492,N_20551,N_23336);
nor UO_1493 (O_1493,N_21415,N_22013);
or UO_1494 (O_1494,N_22175,N_21594);
or UO_1495 (O_1495,N_24564,N_20641);
or UO_1496 (O_1496,N_23235,N_21182);
and UO_1497 (O_1497,N_21401,N_21723);
nor UO_1498 (O_1498,N_24127,N_24765);
nand UO_1499 (O_1499,N_23406,N_22480);
nor UO_1500 (O_1500,N_20689,N_22972);
nor UO_1501 (O_1501,N_23283,N_21931);
nor UO_1502 (O_1502,N_22024,N_24762);
nand UO_1503 (O_1503,N_20240,N_22577);
nor UO_1504 (O_1504,N_23525,N_21283);
xor UO_1505 (O_1505,N_23790,N_22683);
and UO_1506 (O_1506,N_20527,N_20486);
nand UO_1507 (O_1507,N_21315,N_24996);
nand UO_1508 (O_1508,N_20730,N_24361);
or UO_1509 (O_1509,N_22854,N_24507);
nor UO_1510 (O_1510,N_20139,N_22025);
xnor UO_1511 (O_1511,N_20711,N_23791);
and UO_1512 (O_1512,N_24627,N_23184);
and UO_1513 (O_1513,N_20251,N_21057);
xnor UO_1514 (O_1514,N_24062,N_21269);
or UO_1515 (O_1515,N_20204,N_21745);
xnor UO_1516 (O_1516,N_24460,N_22549);
nand UO_1517 (O_1517,N_23211,N_24681);
nand UO_1518 (O_1518,N_23731,N_23830);
xor UO_1519 (O_1519,N_22201,N_22202);
nand UO_1520 (O_1520,N_22953,N_23349);
or UO_1521 (O_1521,N_20037,N_20601);
nor UO_1522 (O_1522,N_22736,N_24541);
nand UO_1523 (O_1523,N_22941,N_20071);
nor UO_1524 (O_1524,N_23266,N_23894);
or UO_1525 (O_1525,N_23824,N_23369);
or UO_1526 (O_1526,N_22330,N_22146);
xor UO_1527 (O_1527,N_24242,N_23536);
nor UO_1528 (O_1528,N_21325,N_21794);
nor UO_1529 (O_1529,N_22855,N_20990);
nand UO_1530 (O_1530,N_21990,N_23041);
nor UO_1531 (O_1531,N_22674,N_24841);
nor UO_1532 (O_1532,N_23050,N_23138);
nand UO_1533 (O_1533,N_21896,N_23969);
or UO_1534 (O_1534,N_23925,N_24019);
nand UO_1535 (O_1535,N_24725,N_24903);
or UO_1536 (O_1536,N_24219,N_24581);
nor UO_1537 (O_1537,N_23000,N_20732);
nand UO_1538 (O_1538,N_20320,N_23559);
and UO_1539 (O_1539,N_24589,N_22372);
and UO_1540 (O_1540,N_23196,N_24521);
nand UO_1541 (O_1541,N_20009,N_24013);
xnor UO_1542 (O_1542,N_23058,N_20201);
xor UO_1543 (O_1543,N_24909,N_24827);
xnor UO_1544 (O_1544,N_20851,N_23545);
nand UO_1545 (O_1545,N_23247,N_22160);
nand UO_1546 (O_1546,N_23251,N_20250);
and UO_1547 (O_1547,N_22828,N_22792);
xnor UO_1548 (O_1548,N_20163,N_20822);
and UO_1549 (O_1549,N_22057,N_24744);
or UO_1550 (O_1550,N_21458,N_24335);
or UO_1551 (O_1551,N_20724,N_24074);
nand UO_1552 (O_1552,N_24314,N_21714);
nor UO_1553 (O_1553,N_23668,N_22629);
nor UO_1554 (O_1554,N_20339,N_23856);
nand UO_1555 (O_1555,N_23870,N_21243);
nand UO_1556 (O_1556,N_23644,N_24037);
and UO_1557 (O_1557,N_22183,N_24343);
nor UO_1558 (O_1558,N_24289,N_23217);
xnor UO_1559 (O_1559,N_23011,N_20708);
nand UO_1560 (O_1560,N_22027,N_20713);
nand UO_1561 (O_1561,N_22601,N_20921);
and UO_1562 (O_1562,N_23705,N_20522);
or UO_1563 (O_1563,N_24743,N_24461);
and UO_1564 (O_1564,N_20273,N_21980);
xnor UO_1565 (O_1565,N_21974,N_22066);
nand UO_1566 (O_1566,N_21875,N_23842);
nand UO_1567 (O_1567,N_21663,N_22246);
nor UO_1568 (O_1568,N_24907,N_23624);
nand UO_1569 (O_1569,N_20131,N_21524);
or UO_1570 (O_1570,N_20501,N_20903);
xor UO_1571 (O_1571,N_21006,N_24672);
and UO_1572 (O_1572,N_23378,N_23764);
or UO_1573 (O_1573,N_21838,N_22375);
nor UO_1574 (O_1574,N_23878,N_22922);
nand UO_1575 (O_1575,N_21841,N_23220);
nor UO_1576 (O_1576,N_21378,N_20628);
xnor UO_1577 (O_1577,N_22858,N_24894);
nor UO_1578 (O_1578,N_23537,N_21053);
or UO_1579 (O_1579,N_20640,N_21908);
xor UO_1580 (O_1580,N_24576,N_23983);
xnor UO_1581 (O_1581,N_21065,N_20877);
nand UO_1582 (O_1582,N_20450,N_23840);
and UO_1583 (O_1583,N_23411,N_23984);
xor UO_1584 (O_1584,N_22010,N_20228);
or UO_1585 (O_1585,N_20925,N_23288);
and UO_1586 (O_1586,N_24585,N_24376);
or UO_1587 (O_1587,N_21950,N_22720);
nor UO_1588 (O_1588,N_23833,N_24686);
and UO_1589 (O_1589,N_20787,N_24419);
nor UO_1590 (O_1590,N_23816,N_20844);
and UO_1591 (O_1591,N_24870,N_20885);
nand UO_1592 (O_1592,N_23089,N_24717);
nand UO_1593 (O_1593,N_22096,N_20482);
xor UO_1594 (O_1594,N_21101,N_24423);
nor UO_1595 (O_1595,N_24088,N_20717);
or UO_1596 (O_1596,N_24623,N_23577);
nand UO_1597 (O_1597,N_20024,N_20077);
xnor UO_1598 (O_1598,N_22232,N_22785);
and UO_1599 (O_1599,N_24737,N_22020);
nor UO_1600 (O_1600,N_24000,N_23860);
nor UO_1601 (O_1601,N_24665,N_23964);
nand UO_1602 (O_1602,N_22442,N_20475);
or UO_1603 (O_1603,N_21856,N_22917);
xnor UO_1604 (O_1604,N_21696,N_22996);
nand UO_1605 (O_1605,N_21196,N_20233);
and UO_1606 (O_1606,N_20553,N_23935);
nand UO_1607 (O_1607,N_22841,N_20053);
nand UO_1608 (O_1608,N_24444,N_20467);
or UO_1609 (O_1609,N_20976,N_24759);
and UO_1610 (O_1610,N_23062,N_24178);
nand UO_1611 (O_1611,N_20720,N_23448);
xor UO_1612 (O_1612,N_21495,N_21097);
xor UO_1613 (O_1613,N_21521,N_20762);
nand UO_1614 (O_1614,N_24813,N_20635);
xnor UO_1615 (O_1615,N_21564,N_20313);
nand UO_1616 (O_1616,N_21556,N_23375);
nor UO_1617 (O_1617,N_24817,N_23012);
nand UO_1618 (O_1618,N_24428,N_24313);
or UO_1619 (O_1619,N_20238,N_21900);
and UO_1620 (O_1620,N_23398,N_24941);
and UO_1621 (O_1621,N_22812,N_23335);
xnor UO_1622 (O_1622,N_20369,N_21568);
xnor UO_1623 (O_1623,N_23561,N_22960);
or UO_1624 (O_1624,N_24805,N_24773);
nand UO_1625 (O_1625,N_23977,N_22721);
and UO_1626 (O_1626,N_20680,N_24300);
or UO_1627 (O_1627,N_22680,N_24850);
xnor UO_1628 (O_1628,N_21300,N_23942);
nand UO_1629 (O_1629,N_21026,N_20534);
xor UO_1630 (O_1630,N_23436,N_23858);
nor UO_1631 (O_1631,N_20050,N_20898);
and UO_1632 (O_1632,N_23387,N_24673);
nor UO_1633 (O_1633,N_24913,N_22611);
nand UO_1634 (O_1634,N_23281,N_20624);
nand UO_1635 (O_1635,N_20156,N_20948);
nor UO_1636 (O_1636,N_24404,N_22898);
nand UO_1637 (O_1637,N_23175,N_23772);
nor UO_1638 (O_1638,N_21734,N_24188);
and UO_1639 (O_1639,N_21606,N_20479);
nor UO_1640 (O_1640,N_22219,N_22810);
or UO_1641 (O_1641,N_24162,N_20493);
xnor UO_1642 (O_1642,N_22378,N_21416);
xor UO_1643 (O_1643,N_20950,N_21383);
or UO_1644 (O_1644,N_20590,N_24501);
nand UO_1645 (O_1645,N_22498,N_20663);
xor UO_1646 (O_1646,N_20284,N_22091);
xnor UO_1647 (O_1647,N_24876,N_24150);
and UO_1648 (O_1648,N_22607,N_21902);
nand UO_1649 (O_1649,N_23533,N_21658);
nand UO_1650 (O_1650,N_24239,N_22774);
and UO_1651 (O_1651,N_21571,N_20442);
xor UO_1652 (O_1652,N_20049,N_20148);
nand UO_1653 (O_1653,N_21347,N_23933);
and UO_1654 (O_1654,N_22250,N_22044);
nor UO_1655 (O_1655,N_21281,N_21632);
and UO_1656 (O_1656,N_21839,N_24333);
or UO_1657 (O_1657,N_21089,N_20563);
or UO_1658 (O_1658,N_24809,N_21095);
nand UO_1659 (O_1659,N_23068,N_20803);
and UO_1660 (O_1660,N_20760,N_21965);
nand UO_1661 (O_1661,N_20890,N_24484);
nand UO_1662 (O_1662,N_22342,N_20078);
and UO_1663 (O_1663,N_21552,N_20126);
nor UO_1664 (O_1664,N_21052,N_21683);
and UO_1665 (O_1665,N_20674,N_23362);
xnor UO_1666 (O_1666,N_24651,N_24143);
xnor UO_1667 (O_1667,N_24186,N_24214);
nor UO_1668 (O_1668,N_24379,N_22338);
or UO_1669 (O_1669,N_20855,N_20888);
nor UO_1670 (O_1670,N_22291,N_20523);
and UO_1671 (O_1671,N_20427,N_22354);
nor UO_1672 (O_1672,N_22716,N_20285);
or UO_1673 (O_1673,N_23037,N_23529);
and UO_1674 (O_1674,N_23710,N_20725);
or UO_1675 (O_1675,N_22547,N_21314);
nor UO_1676 (O_1676,N_23526,N_22225);
nand UO_1677 (O_1677,N_20359,N_22770);
or UO_1678 (O_1678,N_24429,N_24856);
and UO_1679 (O_1679,N_20003,N_22197);
and UO_1680 (O_1680,N_20695,N_24831);
xnor UO_1681 (O_1681,N_22313,N_21549);
nand UO_1682 (O_1682,N_23007,N_23107);
and UO_1683 (O_1683,N_23877,N_23554);
and UO_1684 (O_1684,N_20029,N_24142);
nand UO_1685 (O_1685,N_23319,N_20546);
nor UO_1686 (O_1686,N_22543,N_20438);
and UO_1687 (O_1687,N_22608,N_20754);
nor UO_1688 (O_1688,N_22314,N_22072);
or UO_1689 (O_1689,N_24273,N_23696);
nand UO_1690 (O_1690,N_20582,N_21317);
nor UO_1691 (O_1691,N_22051,N_23779);
nand UO_1692 (O_1692,N_24299,N_24156);
xnor UO_1693 (O_1693,N_22065,N_20692);
or UO_1694 (O_1694,N_23789,N_23848);
xor UO_1695 (O_1695,N_21724,N_24697);
nor UO_1696 (O_1696,N_23390,N_22036);
nand UO_1697 (O_1697,N_21122,N_20305);
xor UO_1698 (O_1698,N_22000,N_22722);
or UO_1699 (O_1699,N_22520,N_24988);
xor UO_1700 (O_1700,N_24974,N_22865);
nor UO_1701 (O_1701,N_21173,N_21353);
or UO_1702 (O_1702,N_21045,N_24911);
or UO_1703 (O_1703,N_21547,N_22466);
xor UO_1704 (O_1704,N_20920,N_23657);
or UO_1705 (O_1705,N_23919,N_23601);
nor UO_1706 (O_1706,N_22054,N_24400);
nand UO_1707 (O_1707,N_20070,N_20064);
and UO_1708 (O_1708,N_24891,N_24990);
nand UO_1709 (O_1709,N_23320,N_22238);
and UO_1710 (O_1710,N_20723,N_24702);
nand UO_1711 (O_1711,N_21651,N_22723);
and UO_1712 (O_1712,N_24036,N_24211);
and UO_1713 (O_1713,N_22838,N_22461);
nor UO_1714 (O_1714,N_20550,N_21453);
xnor UO_1715 (O_1715,N_22414,N_23921);
xnor UO_1716 (O_1716,N_23692,N_20110);
nand UO_1717 (O_1717,N_24181,N_22438);
xnor UO_1718 (O_1718,N_23875,N_24705);
and UO_1719 (O_1719,N_20481,N_20474);
nand UO_1720 (O_1720,N_23337,N_24165);
nand UO_1721 (O_1721,N_22193,N_23841);
nor UO_1722 (O_1722,N_24228,N_23767);
xnor UO_1723 (O_1723,N_24806,N_21523);
and UO_1724 (O_1724,N_21532,N_23361);
xnor UO_1725 (O_1725,N_24711,N_20311);
or UO_1726 (O_1726,N_22133,N_23666);
nand UO_1727 (O_1727,N_20846,N_22161);
or UO_1728 (O_1728,N_24803,N_22450);
xnor UO_1729 (O_1729,N_23364,N_24106);
xnor UO_1730 (O_1730,N_24535,N_22029);
xor UO_1731 (O_1731,N_20061,N_24684);
or UO_1732 (O_1732,N_20038,N_21726);
xnor UO_1733 (O_1733,N_22916,N_20410);
xnor UO_1734 (O_1734,N_23206,N_21751);
nor UO_1735 (O_1735,N_21319,N_22277);
nor UO_1736 (O_1736,N_20170,N_21656);
or UO_1737 (O_1737,N_21409,N_21068);
and UO_1738 (O_1738,N_24925,N_24607);
nor UO_1739 (O_1739,N_22171,N_23724);
nand UO_1740 (O_1740,N_21713,N_20073);
xor UO_1741 (O_1741,N_23165,N_21164);
nand UO_1742 (O_1742,N_20381,N_21075);
xor UO_1743 (O_1743,N_23278,N_22676);
or UO_1744 (O_1744,N_22651,N_24950);
and UO_1745 (O_1745,N_23802,N_20368);
or UO_1746 (O_1746,N_21354,N_22760);
nand UO_1747 (O_1747,N_21976,N_21238);
nand UO_1748 (O_1748,N_24337,N_24723);
or UO_1749 (O_1749,N_21677,N_24303);
nand UO_1750 (O_1750,N_22908,N_20530);
nand UO_1751 (O_1751,N_22179,N_22402);
nand UO_1752 (O_1752,N_24117,N_22843);
and UO_1753 (O_1753,N_20528,N_23134);
nor UO_1754 (O_1754,N_24099,N_21778);
or UO_1755 (O_1755,N_23155,N_21373);
xor UO_1756 (O_1756,N_20772,N_24582);
or UO_1757 (O_1757,N_22265,N_22558);
xor UO_1758 (O_1758,N_22060,N_22515);
nand UO_1759 (O_1759,N_24001,N_21340);
and UO_1760 (O_1760,N_20161,N_23673);
nand UO_1761 (O_1761,N_23807,N_20489);
nand UO_1762 (O_1762,N_23063,N_20979);
nor UO_1763 (O_1763,N_21402,N_21624);
or UO_1764 (O_1764,N_24122,N_23742);
nand UO_1765 (O_1765,N_24970,N_20444);
nor UO_1766 (O_1766,N_23549,N_23728);
xnor UO_1767 (O_1767,N_21299,N_23356);
nor UO_1768 (O_1768,N_21027,N_21608);
and UO_1769 (O_1769,N_21585,N_23342);
and UO_1770 (O_1770,N_20963,N_23874);
nor UO_1771 (O_1771,N_20927,N_23425);
nor UO_1772 (O_1772,N_20422,N_20719);
xnor UO_1773 (O_1773,N_20827,N_23922);
or UO_1774 (O_1774,N_24007,N_21679);
or UO_1775 (O_1775,N_24830,N_22776);
nor UO_1776 (O_1776,N_21540,N_20672);
nand UO_1777 (O_1777,N_21923,N_24628);
and UO_1778 (O_1778,N_23341,N_20389);
or UO_1779 (O_1779,N_23002,N_22999);
nand UO_1780 (O_1780,N_24421,N_21800);
or UO_1781 (O_1781,N_23015,N_24545);
or UO_1782 (O_1782,N_23415,N_24477);
xnor UO_1783 (O_1783,N_20041,N_20741);
and UO_1784 (O_1784,N_24955,N_24574);
or UO_1785 (O_1785,N_21115,N_22540);
nor UO_1786 (O_1786,N_22926,N_22333);
or UO_1787 (O_1787,N_21645,N_23552);
nand UO_1788 (O_1788,N_23119,N_24225);
nand UO_1789 (O_1789,N_22081,N_21686);
nand UO_1790 (O_1790,N_23825,N_20297);
and UO_1791 (O_1791,N_23079,N_23608);
nor UO_1792 (O_1792,N_20779,N_20330);
and UO_1793 (O_1793,N_20579,N_23164);
and UO_1794 (O_1794,N_21162,N_20499);
xor UO_1795 (O_1795,N_23557,N_20319);
xor UO_1796 (O_1796,N_20634,N_21625);
nand UO_1797 (O_1797,N_20244,N_20881);
xnor UO_1798 (O_1798,N_24213,N_23938);
and UO_1799 (O_1799,N_21642,N_21809);
xnor UO_1800 (O_1800,N_22630,N_20355);
nor UO_1801 (O_1801,N_23519,N_20974);
or UO_1802 (O_1802,N_24987,N_22451);
xnor UO_1803 (O_1803,N_23204,N_23952);
nand UO_1804 (O_1804,N_20066,N_20612);
xor UO_1805 (O_1805,N_20697,N_22829);
xnor UO_1806 (O_1806,N_23114,N_24012);
and UO_1807 (O_1807,N_23495,N_22818);
and UO_1808 (O_1808,N_22334,N_20035);
nor UO_1809 (O_1809,N_23115,N_24043);
xor UO_1810 (O_1810,N_23456,N_24155);
or UO_1811 (O_1811,N_21246,N_23598);
nor UO_1812 (O_1812,N_23168,N_20895);
and UO_1813 (O_1813,N_20565,N_21404);
or UO_1814 (O_1814,N_20883,N_24543);
xor UO_1815 (O_1815,N_23239,N_24068);
nand UO_1816 (O_1816,N_24158,N_24318);
or UO_1817 (O_1817,N_22336,N_20441);
or UO_1818 (O_1818,N_22268,N_20718);
or UO_1819 (O_1819,N_23473,N_23837);
nor UO_1820 (O_1820,N_23176,N_22173);
nor UO_1821 (O_1821,N_20224,N_21953);
nand UO_1822 (O_1822,N_22552,N_23009);
nor UO_1823 (O_1823,N_23128,N_22434);
xnor UO_1824 (O_1824,N_22884,N_21937);
or UO_1825 (O_1825,N_21309,N_21457);
xor UO_1826 (O_1826,N_22249,N_20657);
nor UO_1827 (O_1827,N_21531,N_24630);
or UO_1828 (O_1828,N_24583,N_21209);
xnor UO_1829 (O_1829,N_20636,N_21788);
nor UO_1830 (O_1830,N_23593,N_20726);
nor UO_1831 (O_1831,N_20650,N_23322);
nand UO_1832 (O_1832,N_22915,N_22493);
nand UO_1833 (O_1833,N_22631,N_24148);
and UO_1834 (O_1834,N_23286,N_23358);
nor UO_1835 (O_1835,N_22505,N_21216);
xor UO_1836 (O_1836,N_20731,N_20473);
nor UO_1837 (O_1837,N_23926,N_21123);
nand UO_1838 (O_1838,N_21298,N_23622);
nor UO_1839 (O_1839,N_21358,N_20770);
and UO_1840 (O_1840,N_23596,N_24320);
nor UO_1841 (O_1841,N_22206,N_20620);
nor UO_1842 (O_1842,N_23864,N_22432);
or UO_1843 (O_1843,N_24417,N_21626);
nor UO_1844 (O_1844,N_24905,N_20177);
and UO_1845 (O_1845,N_20985,N_21501);
nor UO_1846 (O_1846,N_21118,N_21211);
nand UO_1847 (O_1847,N_21784,N_23078);
nand UO_1848 (O_1848,N_21767,N_23351);
or UO_1849 (O_1849,N_21848,N_22788);
xnor UO_1850 (O_1850,N_20075,N_23655);
nand UO_1851 (O_1851,N_20302,N_20958);
nor UO_1852 (O_1852,N_22624,N_23044);
nor UO_1853 (O_1853,N_22927,N_21699);
nor UO_1854 (O_1854,N_24021,N_24152);
or UO_1855 (O_1855,N_22294,N_20157);
xor UO_1856 (O_1856,N_22264,N_20298);
xor UO_1857 (O_1857,N_22316,N_23135);
nor UO_1858 (O_1858,N_21337,N_21244);
and UO_1859 (O_1859,N_20904,N_22599);
and UO_1860 (O_1860,N_22273,N_20774);
or UO_1861 (O_1861,N_22696,N_24080);
and UO_1862 (O_1862,N_22440,N_21344);
or UO_1863 (O_1863,N_23573,N_21165);
and UO_1864 (O_1864,N_21633,N_22413);
or UO_1865 (O_1865,N_24662,N_24073);
or UO_1866 (O_1866,N_21823,N_20084);
xnor UO_1867 (O_1867,N_23346,N_24566);
xnor UO_1868 (O_1868,N_24393,N_23150);
and UO_1869 (O_1869,N_21077,N_20610);
nand UO_1870 (O_1870,N_23467,N_24534);
xnor UO_1871 (O_1871,N_22715,N_21073);
nor UO_1872 (O_1872,N_21510,N_20367);
xnor UO_1873 (O_1873,N_20265,N_23073);
nand UO_1874 (O_1874,N_23345,N_24638);
and UO_1875 (O_1875,N_21444,N_22276);
nand UO_1876 (O_1876,N_22126,N_22182);
nor UO_1877 (O_1877,N_20670,N_22308);
xnor UO_1878 (O_1878,N_24730,N_22234);
nor UO_1879 (O_1879,N_20745,N_21582);
or UO_1880 (O_1880,N_22991,N_24125);
or UO_1881 (O_1881,N_21094,N_22582);
xnor UO_1882 (O_1882,N_20625,N_22831);
nand UO_1883 (O_1883,N_22460,N_23194);
or UO_1884 (O_1884,N_23570,N_21762);
xor UO_1885 (O_1885,N_22105,N_22757);
or UO_1886 (O_1886,N_22837,N_20712);
or UO_1887 (O_1887,N_21186,N_23843);
nor UO_1888 (O_1888,N_21630,N_24804);
and UO_1889 (O_1889,N_23477,N_23897);
or UO_1890 (O_1890,N_22470,N_24878);
and UO_1891 (O_1891,N_24963,N_23071);
nor UO_1892 (O_1892,N_23715,N_24377);
nand UO_1893 (O_1893,N_20767,N_24599);
xnor UO_1894 (O_1894,N_24071,N_20863);
nand UO_1895 (O_1895,N_23804,N_21774);
xor UO_1896 (O_1896,N_23053,N_22080);
or UO_1897 (O_1897,N_21293,N_23421);
xor UO_1898 (O_1898,N_24060,N_21009);
nand UO_1899 (O_1899,N_22563,N_23173);
xor UO_1900 (O_1900,N_24203,N_21737);
nor UO_1901 (O_1901,N_22832,N_23817);
nand UO_1902 (O_1902,N_20811,N_24910);
or UO_1903 (O_1903,N_21225,N_23257);
nor UO_1904 (O_1904,N_20119,N_20309);
nand UO_1905 (O_1905,N_20391,N_22155);
nand UO_1906 (O_1906,N_21853,N_21435);
xnor UO_1907 (O_1907,N_24592,N_24978);
nand UO_1908 (O_1908,N_24906,N_22103);
nor UO_1909 (O_1909,N_22324,N_23045);
and UO_1910 (O_1910,N_21126,N_24282);
and UO_1911 (O_1911,N_21660,N_24061);
xnor UO_1912 (O_1912,N_20466,N_21629);
nand UO_1913 (O_1913,N_22672,N_24942);
or UO_1914 (O_1914,N_23663,N_23866);
nor UO_1915 (O_1915,N_20897,N_22681);
or UO_1916 (O_1916,N_22387,N_23277);
or UO_1917 (O_1917,N_20190,N_22123);
or UO_1918 (O_1918,N_24447,N_24350);
nor UO_1919 (O_1919,N_21761,N_21554);
and UO_1920 (O_1920,N_21618,N_21085);
nand UO_1921 (O_1921,N_22506,N_23518);
or UO_1922 (O_1922,N_20918,N_22677);
nand UO_1923 (O_1923,N_20142,N_22003);
or UO_1924 (O_1924,N_20847,N_22744);
or UO_1925 (O_1925,N_21708,N_23717);
nor UO_1926 (O_1926,N_24802,N_22839);
and UO_1927 (O_1927,N_20519,N_21076);
or UO_1928 (O_1928,N_21756,N_23148);
or UO_1929 (O_1929,N_24657,N_20011);
nand UO_1930 (O_1930,N_23487,N_21374);
and UO_1931 (O_1931,N_24109,N_22659);
or UO_1932 (O_1932,N_23892,N_21330);
and UO_1933 (O_1933,N_22724,N_20278);
or UO_1934 (O_1934,N_23750,N_24617);
and UO_1935 (O_1935,N_24838,N_22041);
nand UO_1936 (O_1936,N_23998,N_23987);
nor UO_1937 (O_1937,N_22641,N_21857);
and UO_1938 (O_1938,N_24767,N_20356);
nand UO_1939 (O_1939,N_23127,N_22240);
or UO_1940 (O_1940,N_20608,N_21116);
or UO_1941 (O_1941,N_21099,N_21471);
nor UO_1942 (O_1942,N_24130,N_20832);
nand UO_1943 (O_1943,N_23783,N_22690);
and UO_1944 (O_1944,N_21557,N_20316);
xnor UO_1945 (O_1945,N_23297,N_21764);
or UO_1946 (O_1946,N_23700,N_20658);
nand UO_1947 (O_1947,N_22303,N_23097);
and UO_1948 (O_1948,N_21881,N_21570);
xnor UO_1949 (O_1949,N_21957,N_23675);
and UO_1950 (O_1950,N_24716,N_22749);
or UO_1951 (O_1951,N_23656,N_20424);
or UO_1952 (O_1952,N_24889,N_23432);
or UO_1953 (O_1953,N_20483,N_20013);
nor UO_1954 (O_1954,N_20246,N_24973);
nor UO_1955 (O_1955,N_22597,N_21673);
xnor UO_1956 (O_1956,N_24786,N_24946);
xor UO_1957 (O_1957,N_20694,N_23566);
or UO_1958 (O_1958,N_24620,N_20561);
nor UO_1959 (O_1959,N_24935,N_20300);
nor UO_1960 (O_1960,N_24392,N_24689);
nor UO_1961 (O_1961,N_21324,N_21786);
or UO_1962 (O_1962,N_24140,N_20054);
or UO_1963 (O_1963,N_22190,N_24261);
nand UO_1964 (O_1964,N_20370,N_24111);
xor UO_1965 (O_1965,N_21301,N_24113);
and UO_1966 (O_1966,N_22598,N_20206);
xnor UO_1967 (O_1967,N_22143,N_23654);
xor UO_1968 (O_1968,N_22836,N_20510);
and UO_1969 (O_1969,N_20942,N_24823);
or UO_1970 (O_1970,N_20630,N_24738);
xnor UO_1971 (O_1971,N_21168,N_21719);
and UO_1972 (O_1972,N_23260,N_23857);
nor UO_1973 (O_1973,N_21508,N_23085);
and UO_1974 (O_1974,N_20764,N_24234);
xnor UO_1975 (O_1975,N_22961,N_24084);
or UO_1976 (O_1976,N_23973,N_20113);
nand UO_1977 (O_1977,N_23703,N_23308);
nand UO_1978 (O_1978,N_23254,N_20964);
or UO_1979 (O_1979,N_20397,N_21580);
xnor UO_1980 (O_1980,N_21998,N_24293);
nor UO_1981 (O_1981,N_24056,N_22185);
or UO_1982 (O_1982,N_23080,N_24659);
nand UO_1983 (O_1983,N_23954,N_24774);
and UO_1984 (O_1984,N_23404,N_20123);
nor UO_1985 (O_1985,N_20589,N_22780);
nand UO_1986 (O_1986,N_24967,N_24904);
nor UO_1987 (O_1987,N_20484,N_22134);
nor UO_1988 (O_1988,N_23186,N_22329);
or UO_1989 (O_1989,N_23188,N_23192);
nand UO_1990 (O_1990,N_20786,N_24440);
nor UO_1991 (O_1991,N_23430,N_21704);
and UO_1992 (O_1992,N_22782,N_20733);
nor UO_1993 (O_1993,N_20052,N_23560);
xnor UO_1994 (O_1994,N_20027,N_23619);
and UO_1995 (O_1995,N_20415,N_23106);
nor UO_1996 (O_1996,N_21217,N_23433);
nor UO_1997 (O_1997,N_24952,N_20965);
nor UO_1998 (O_1998,N_20826,N_21866);
nor UO_1999 (O_1999,N_24953,N_21898);
and UO_2000 (O_2000,N_23460,N_24259);
nor UO_2001 (O_2001,N_24272,N_22627);
nor UO_2002 (O_2002,N_21903,N_20867);
nor UO_2003 (O_2003,N_24164,N_23756);
and UO_2004 (O_2004,N_24183,N_23555);
and UO_2005 (O_2005,N_20690,N_24334);
xor UO_2006 (O_2006,N_24281,N_22266);
or UO_2007 (O_2007,N_21739,N_21765);
and UO_2008 (O_2008,N_22379,N_23868);
nand UO_2009 (O_2009,N_22527,N_20361);
nand UO_2010 (O_2010,N_21994,N_20568);
nor UO_2011 (O_2011,N_22317,N_21442);
nand UO_2012 (O_2012,N_22292,N_22258);
nand UO_2013 (O_2013,N_22758,N_22211);
and UO_2014 (O_2014,N_21369,N_22717);
or UO_2015 (O_2015,N_22271,N_20399);
nand UO_2016 (O_2016,N_22583,N_23911);
nor UO_2017 (O_2017,N_20567,N_20406);
or UO_2018 (O_2018,N_21951,N_20750);
or UO_2019 (O_2019,N_23782,N_20880);
or UO_2020 (O_2020,N_21909,N_21437);
nor UO_2021 (O_2021,N_21280,N_23975);
nand UO_2022 (O_2022,N_24058,N_24932);
nor UO_2023 (O_2023,N_24556,N_24131);
and UO_2024 (O_2024,N_24644,N_24663);
nor UO_2025 (O_2025,N_22089,N_23355);
or UO_2026 (O_2026,N_22306,N_23828);
or UO_2027 (O_2027,N_20806,N_22700);
or UO_2028 (O_2028,N_21312,N_23488);
nand UO_2029 (O_2029,N_24353,N_20644);
nor UO_2030 (O_2030,N_23967,N_22100);
nor UO_2031 (O_2031,N_22135,N_21349);
nor UO_2032 (O_2032,N_20398,N_22962);
and UO_2033 (O_2033,N_24960,N_22398);
and UO_2034 (O_2034,N_24671,N_23373);
nand UO_2035 (O_2035,N_20137,N_23839);
nand UO_2036 (O_2036,N_20916,N_20626);
and UO_2037 (O_2037,N_20852,N_21034);
xnor UO_2038 (O_2038,N_21208,N_23635);
xnor UO_2039 (O_2039,N_20016,N_20328);
nor UO_2040 (O_2040,N_23590,N_24632);
nand UO_2041 (O_2041,N_24519,N_24129);
and UO_2042 (O_2042,N_20722,N_24847);
and UO_2043 (O_2043,N_22666,N_20611);
nor UO_2044 (O_2044,N_24529,N_23517);
nor UO_2045 (O_2045,N_20403,N_22148);
xnor UO_2046 (O_2046,N_22887,N_20710);
or UO_2047 (O_2047,N_21641,N_23993);
xnor UO_2048 (O_2048,N_21617,N_21512);
or UO_2049 (O_2049,N_22645,N_21969);
nor UO_2050 (O_2050,N_20808,N_22755);
or UO_2051 (O_2051,N_22985,N_21486);
nand UO_2052 (O_2052,N_20379,N_20417);
or UO_2053 (O_2053,N_24568,N_23630);
or UO_2054 (O_2054,N_23862,N_21820);
or UO_2055 (O_2055,N_23915,N_22298);
nand UO_2056 (O_2056,N_20014,N_23992);
or UO_2057 (O_2057,N_21219,N_23890);
or UO_2058 (O_2058,N_24914,N_24505);
nand UO_2059 (O_2059,N_21468,N_24151);
and UO_2060 (O_2060,N_24312,N_22424);
and UO_2061 (O_2061,N_24557,N_22366);
xnor UO_2062 (O_2062,N_22593,N_23400);
or UO_2063 (O_2063,N_20015,N_22001);
nand UO_2064 (O_2064,N_21989,N_22261);
xnor UO_2065 (O_2065,N_24692,N_24121);
or UO_2066 (O_2066,N_22518,N_24522);
and UO_2067 (O_2067,N_21367,N_21669);
and UO_2068 (O_2068,N_22192,N_24912);
nand UO_2069 (O_2069,N_24120,N_22321);
or UO_2070 (O_2070,N_20431,N_21463);
nand UO_2071 (O_2071,N_20112,N_21859);
xor UO_2072 (O_2072,N_24328,N_23735);
nand UO_2073 (O_2073,N_24489,N_24771);
or UO_2074 (O_2074,N_22416,N_21725);
nand UO_2075 (O_2075,N_20514,N_22779);
nand UO_2076 (O_2076,N_20435,N_20682);
and UO_2077 (O_2077,N_20631,N_23597);
nor UO_2078 (O_2078,N_20757,N_23587);
nand UO_2079 (O_2079,N_24555,N_21869);
nor UO_2080 (O_2080,N_20045,N_22168);
and UO_2081 (O_2081,N_20862,N_20325);
or UO_2082 (O_2082,N_22823,N_21805);
nor UO_2083 (O_2083,N_24089,N_21237);
xor UO_2084 (O_2084,N_20130,N_23613);
nor UO_2085 (O_2085,N_23736,N_22642);
and UO_2086 (O_2086,N_20219,N_24016);
or UO_2087 (O_2087,N_20584,N_24370);
and UO_2088 (O_2088,N_21935,N_20752);
nand UO_2089 (O_2089,N_22772,N_23694);
nor UO_2090 (O_2090,N_21131,N_22279);
or UO_2091 (O_2091,N_22514,N_23108);
nand UO_2092 (O_2092,N_20031,N_23732);
or UO_2093 (O_2093,N_23049,N_21722);
nand UO_2094 (O_2094,N_20555,N_21223);
or UO_2095 (O_2095,N_20954,N_22393);
and UO_2096 (O_2096,N_20543,N_20889);
nor UO_2097 (O_2097,N_23386,N_22817);
xnor UO_2098 (O_2098,N_23838,N_22441);
nor UO_2099 (O_2099,N_22819,N_24931);
xor UO_2100 (O_2100,N_21456,N_21203);
nor UO_2101 (O_2101,N_22454,N_22410);
and UO_2102 (O_2102,N_24691,N_23036);
and UO_2103 (O_2103,N_20335,N_21055);
or UO_2104 (O_2104,N_21142,N_21109);
and UO_2105 (O_2105,N_23794,N_20079);
or UO_2106 (O_2106,N_24742,N_24138);
nand UO_2107 (O_2107,N_24981,N_20613);
xor UO_2108 (O_2108,N_23678,N_23234);
or UO_2109 (O_2109,N_23712,N_20277);
xnor UO_2110 (O_2110,N_20416,N_24049);
xor UO_2111 (O_2111,N_20195,N_22093);
nor UO_2112 (O_2112,N_20819,N_21825);
nor UO_2113 (O_2113,N_23303,N_20270);
and UO_2114 (O_2114,N_21581,N_21016);
nor UO_2115 (O_2115,N_21078,N_24311);
nor UO_2116 (O_2116,N_21163,N_23166);
and UO_2117 (O_2117,N_22474,N_24573);
xor UO_2118 (O_2118,N_23947,N_23836);
nand UO_2119 (O_2119,N_23907,N_21979);
or UO_2120 (O_2120,N_20144,N_24603);
or UO_2121 (O_2121,N_21668,N_22154);
nor UO_2122 (O_2122,N_20656,N_22967);
xnor UO_2123 (O_2123,N_21381,N_20782);
nand UO_2124 (O_2124,N_24445,N_23236);
nand UO_2125 (O_2125,N_22120,N_24128);
nor UO_2126 (O_2126,N_22512,N_20744);
and UO_2127 (O_2127,N_23120,N_23652);
or UO_2128 (O_2128,N_21672,N_21124);
or UO_2129 (O_2129,N_20923,N_24260);
nor UO_2130 (O_2130,N_23558,N_23583);
nor UO_2131 (O_2131,N_20146,N_23201);
xnor UO_2132 (O_2132,N_22846,N_23453);
xor UO_2133 (O_2133,N_21783,N_20172);
nor UO_2134 (O_2134,N_20279,N_22083);
xor UO_2135 (O_2135,N_23472,N_24283);
and UO_2136 (O_2136,N_24451,N_24516);
and UO_2137 (O_2137,N_22403,N_21228);
or UO_2138 (O_2138,N_23605,N_23535);
nor UO_2139 (O_2139,N_20237,N_22670);
xnor UO_2140 (O_2140,N_21384,N_22743);
nor UO_2141 (O_2141,N_24365,N_21854);
nor UO_2142 (O_2142,N_23112,N_20349);
or UO_2143 (O_2143,N_24097,N_24776);
nand UO_2144 (O_2144,N_23082,N_22491);
xor UO_2145 (O_2145,N_22682,N_21610);
and UO_2146 (O_2146,N_20072,N_22226);
xor UO_2147 (O_2147,N_24559,N_23674);
and UO_2148 (O_2148,N_21812,N_20971);
or UO_2149 (O_2149,N_20378,N_21500);
or UO_2150 (O_2150,N_22801,N_24848);
and UO_2151 (O_2151,N_21171,N_21331);
or UO_2152 (O_2152,N_21861,N_21802);
or UO_2153 (O_2153,N_21559,N_20227);
nand UO_2154 (O_2154,N_24783,N_23823);
xor UO_2155 (O_2155,N_20747,N_21653);
xnor UO_2156 (O_2156,N_24408,N_22850);
or UO_2157 (O_2157,N_23156,N_20751);
and UO_2158 (O_2158,N_21518,N_23189);
xor UO_2159 (O_2159,N_24828,N_22803);
or UO_2160 (O_2160,N_20488,N_24852);
xor UO_2161 (O_2161,N_21982,N_20187);
xnor UO_2162 (O_2162,N_22554,N_23639);
nor UO_2163 (O_2163,N_21715,N_24943);
or UO_2164 (O_2164,N_21398,N_24465);
xor UO_2165 (O_2165,N_20957,N_23153);
or UO_2166 (O_2166,N_23748,N_22588);
nor UO_2167 (O_2167,N_22728,N_21553);
nor UO_2168 (O_2168,N_22473,N_21566);
or UO_2169 (O_2169,N_21483,N_23506);
xor UO_2170 (O_2170,N_22289,N_20494);
or UO_2171 (O_2171,N_22847,N_21410);
or UO_2172 (O_2172,N_23813,N_21278);
nand UO_2173 (O_2173,N_24640,N_22522);
nor UO_2174 (O_2174,N_21130,N_24481);
nand UO_2175 (O_2175,N_21863,N_21760);
xnor UO_2176 (O_2176,N_20987,N_22998);
nor UO_2177 (O_2177,N_21845,N_23245);
nor UO_2178 (O_2178,N_20566,N_22104);
nor UO_2179 (O_2179,N_24518,N_22564);
and UO_2180 (O_2180,N_22290,N_23243);
xor UO_2181 (O_2181,N_22026,N_22269);
nand UO_2182 (O_2182,N_20821,N_24799);
nor UO_2183 (O_2183,N_22754,N_24455);
nand UO_2184 (O_2184,N_24624,N_20995);
xnor UO_2185 (O_2185,N_23271,N_20117);
xnor UO_2186 (O_2186,N_21711,N_21763);
nand UO_2187 (O_2187,N_24693,N_21127);
and UO_2188 (O_2188,N_20947,N_22367);
or UO_2189 (O_2189,N_24044,N_22954);
xnor UO_2190 (O_2190,N_21933,N_24189);
xnor UO_2191 (O_2191,N_21506,N_22049);
nand UO_2192 (O_2192,N_23999,N_21241);
or UO_2193 (O_2193,N_22873,N_24041);
nand UO_2194 (O_2194,N_24325,N_24182);
nor UO_2195 (O_2195,N_23822,N_22525);
or UO_2196 (O_2196,N_20910,N_21995);
or UO_2197 (O_2197,N_22159,N_24226);
nand UO_2198 (O_2198,N_24115,N_22648);
nor UO_2199 (O_2199,N_24326,N_20096);
and UO_2200 (O_2200,N_24055,N_20281);
xnor UO_2201 (O_2201,N_21139,N_21176);
nor UO_2202 (O_2202,N_21499,N_21526);
or UO_2203 (O_2203,N_23329,N_20409);
and UO_2204 (O_2204,N_24641,N_23223);
and UO_2205 (O_2205,N_20382,N_23222);
nand UO_2206 (O_2206,N_21742,N_22489);
or UO_2207 (O_2207,N_23174,N_21159);
and UO_2208 (O_2208,N_22293,N_21910);
and UO_2209 (O_2209,N_22619,N_22449);
or UO_2210 (O_2210,N_23659,N_20017);
nor UO_2211 (O_2211,N_22544,N_23512);
or UO_2212 (O_2212,N_23077,N_22614);
and UO_2213 (O_2213,N_21484,N_22149);
nor UO_2214 (O_2214,N_22859,N_21720);
or UO_2215 (O_2215,N_20721,N_24147);
nor UO_2216 (O_2216,N_24132,N_21947);
xnor UO_2217 (O_2217,N_24956,N_23395);
nand UO_2218 (O_2218,N_22034,N_20516);
nor UO_2219 (O_2219,N_24544,N_21137);
xor UO_2220 (O_2220,N_24190,N_22300);
xnor UO_2221 (O_2221,N_20840,N_21674);
xnor UO_2222 (O_2222,N_23539,N_23504);
nand UO_2223 (O_2223,N_22769,N_24754);
and UO_2224 (O_2224,N_24274,N_22032);
and UO_2225 (O_2225,N_22494,N_24864);
and UO_2226 (O_2226,N_21355,N_21628);
and UO_2227 (O_2227,N_24171,N_24458);
or UO_2228 (O_2228,N_22857,N_20395);
nand UO_2229 (O_2229,N_24090,N_21700);
or UO_2230 (O_2230,N_24578,N_23885);
or UO_2231 (O_2231,N_24818,N_22923);
nor UO_2232 (O_2232,N_23891,N_23505);
nand UO_2233 (O_2233,N_21885,N_23585);
and UO_2234 (O_2234,N_20727,N_22464);
or UO_2235 (O_2235,N_21852,N_24618);
nand UO_2236 (O_2236,N_22984,N_22888);
nor UO_2237 (O_2237,N_22344,N_23376);
and UO_2238 (O_2238,N_21038,N_20363);
or UO_2239 (O_2239,N_20153,N_20547);
and UO_2240 (O_2240,N_21963,N_23784);
nand UO_2241 (O_2241,N_20538,N_23749);
nor UO_2242 (O_2242,N_21962,N_24367);
nand UO_2243 (O_2243,N_22109,N_24483);
and UO_2244 (O_2244,N_22751,N_24279);
and UO_2245 (O_2245,N_21652,N_23394);
nor UO_2246 (O_2246,N_24703,N_23438);
nor UO_2247 (O_2247,N_23072,N_24509);
nor UO_2248 (O_2248,N_20056,N_22328);
and UO_2249 (O_2249,N_21202,N_24900);
or UO_2250 (O_2250,N_20134,N_22649);
nor UO_2251 (O_2251,N_24433,N_22228);
nand UO_2252 (O_2252,N_24562,N_22076);
nor UO_2253 (O_2253,N_22177,N_21717);
nand UO_2254 (O_2254,N_24504,N_21607);
nor UO_2255 (O_2255,N_22107,N_22612);
xor UO_2256 (O_2256,N_20272,N_21539);
and UO_2257 (O_2257,N_23820,N_23626);
nand UO_2258 (O_2258,N_20837,N_22331);
nor UO_2259 (O_2259,N_21286,N_23576);
nand UO_2260 (O_2260,N_24304,N_24965);
nor UO_2261 (O_2261,N_24546,N_24025);
or UO_2262 (O_2262,N_24710,N_20868);
and UO_2263 (O_2263,N_23116,N_20996);
nor UO_2264 (O_2264,N_24342,N_21851);
nand UO_2265 (O_2265,N_21446,N_23645);
xnor UO_2266 (O_2266,N_23851,N_22500);
and UO_2267 (O_2267,N_22541,N_20239);
nor UO_2268 (O_2268,N_22555,N_20090);
or UO_2269 (O_2269,N_24551,N_23498);
or UO_2270 (O_2270,N_22781,N_24267);
or UO_2271 (O_2271,N_24372,N_20632);
nor UO_2272 (O_2272,N_22132,N_21517);
xor UO_2273 (O_2273,N_23126,N_22295);
or UO_2274 (O_2274,N_20326,N_21949);
or UO_2275 (O_2275,N_23483,N_20780);
nand UO_2276 (O_2276,N_21464,N_20028);
and UO_2277 (O_2277,N_21836,N_23927);
and UO_2278 (O_2278,N_24383,N_21487);
or UO_2279 (O_2279,N_23380,N_24107);
nor UO_2280 (O_2280,N_21834,N_23221);
and UO_2281 (O_2281,N_22078,N_24766);
or UO_2282 (O_2282,N_24785,N_21198);
or UO_2283 (O_2283,N_23439,N_24237);
xnor UO_2284 (O_2284,N_24895,N_21305);
xor UO_2285 (O_2285,N_24882,N_20828);
or UO_2286 (O_2286,N_23950,N_20097);
xnor UO_2287 (O_2287,N_24654,N_21380);
nor UO_2288 (O_2288,N_21515,N_20147);
or UO_2289 (O_2289,N_21504,N_21530);
xor UO_2290 (O_2290,N_24569,N_22058);
or UO_2291 (O_2291,N_23191,N_23811);
nor UO_2292 (O_2292,N_23556,N_21595);
or UO_2293 (O_2293,N_22679,N_20776);
nor UO_2294 (O_2294,N_24790,N_22691);
nand UO_2295 (O_2295,N_24835,N_21941);
nand UO_2296 (O_2296,N_22247,N_21766);
and UO_2297 (O_2297,N_20182,N_21528);
xor UO_2298 (O_2298,N_24052,N_22189);
or UO_2299 (O_2299,N_23905,N_24712);
xnor UO_2300 (O_2300,N_23751,N_22035);
nand UO_2301 (O_2301,N_24958,N_24677);
nor UO_2302 (O_2302,N_21926,N_23904);
and UO_2303 (O_2303,N_20338,N_22609);
nand UO_2304 (O_2304,N_24816,N_22355);
and UO_2305 (O_2305,N_23417,N_22121);
nor UO_2306 (O_2306,N_22958,N_21379);
nand UO_2307 (O_2307,N_23564,N_22082);
nor UO_2308 (O_2308,N_23771,N_22064);
or UO_2309 (O_2309,N_22007,N_20966);
and UO_2310 (O_2310,N_24984,N_23136);
nor UO_2311 (O_2311,N_22729,N_24199);
nor UO_2312 (O_2312,N_22038,N_21434);
and UO_2313 (O_2313,N_20676,N_23124);
and UO_2314 (O_2314,N_23256,N_21810);
or UO_2315 (O_2315,N_21474,N_20542);
nor UO_2316 (O_2316,N_23677,N_23547);
xnor UO_2317 (O_2317,N_24224,N_21721);
nand UO_2318 (O_2318,N_23936,N_20677);
or UO_2319 (O_2319,N_22883,N_21801);
or UO_2320 (O_2320,N_24588,N_21475);
nand UO_2321 (O_2321,N_24252,N_21942);
nor UO_2322 (O_2322,N_21261,N_23757);
nor UO_2323 (O_2323,N_20748,N_21598);
nor UO_2324 (O_2324,N_22613,N_22957);
nand UO_2325 (O_2325,N_22501,N_23643);
and UO_2326 (O_2326,N_22374,N_23507);
nand UO_2327 (O_2327,N_20257,N_23090);
or UO_2328 (O_2328,N_21467,N_23881);
nand UO_2329 (O_2329,N_22304,N_24395);
or UO_2330 (O_2330,N_24945,N_24184);
xor UO_2331 (O_2331,N_20180,N_23469);
nor UO_2332 (O_2332,N_22028,N_20836);
nand UO_2333 (O_2333,N_24166,N_22526);
nand UO_2334 (O_2334,N_22115,N_23819);
nor UO_2335 (O_2335,N_21426,N_24998);
xor UO_2336 (O_2336,N_23388,N_21441);
xor UO_2337 (O_2337,N_21736,N_20030);
nand UO_2338 (O_2338,N_20944,N_21572);
and UO_2339 (O_2339,N_23343,N_21121);
nand UO_2340 (O_2340,N_22892,N_24098);
or UO_2341 (O_2341,N_22511,N_21690);
xnor UO_2342 (O_2342,N_24756,N_23781);
or UO_2343 (O_2343,N_20200,N_21447);
and UO_2344 (O_2344,N_24729,N_21161);
or UO_2345 (O_2345,N_23527,N_23649);
nor UO_2346 (O_2346,N_24193,N_24724);
and UO_2347 (O_2347,N_24217,N_22969);
nor UO_2348 (O_2348,N_24473,N_20816);
xnor UO_2349 (O_2349,N_20315,N_20022);
xnor UO_2350 (O_2350,N_21792,N_24896);
and UO_2351 (O_2351,N_22341,N_20133);
nor UO_2352 (O_2352,N_24396,N_24174);
nor UO_2353 (O_2353,N_23889,N_23637);
nor UO_2354 (O_2354,N_22580,N_21049);
and UO_2355 (O_2355,N_24825,N_22976);
nand UO_2356 (O_2356,N_21932,N_23989);
nor UO_2357 (O_2357,N_20210,N_22881);
and UO_2358 (O_2358,N_20785,N_23212);
nand UO_2359 (O_2359,N_20891,N_20271);
nand UO_2360 (O_2360,N_22634,N_21251);
xor UO_2361 (O_2361,N_24200,N_24284);
nand UO_2362 (O_2362,N_23065,N_22147);
and UO_2363 (O_2363,N_23143,N_23030);
or UO_2364 (O_2364,N_22165,N_24112);
and UO_2365 (O_2365,N_22176,N_22773);
xnor UO_2366 (O_2366,N_23042,N_24278);
xor UO_2367 (O_2367,N_24777,N_24443);
nand UO_2368 (O_2368,N_22948,N_21316);
nand UO_2369 (O_2369,N_24957,N_24339);
or UO_2370 (O_2370,N_20040,N_21728);
nor UO_2371 (O_2371,N_24597,N_21563);
or UO_2372 (O_2372,N_22285,N_20873);
nand UO_2373 (O_2373,N_21455,N_23500);
nor UO_2374 (O_2374,N_24643,N_22535);
xor UO_2375 (O_2375,N_23910,N_22834);
and UO_2376 (O_2376,N_21405,N_22288);
and UO_2377 (O_2377,N_22047,N_22561);
xnor UO_2378 (O_2378,N_20556,N_21296);
nand UO_2379 (O_2379,N_21946,N_23125);
nor UO_2380 (O_2380,N_20970,N_24322);
nor UO_2381 (O_2381,N_20876,N_20907);
nor UO_2382 (O_2382,N_23826,N_22163);
xnor UO_2383 (O_2383,N_23913,N_21245);
or UO_2384 (O_2384,N_24418,N_23444);
or UO_2385 (O_2385,N_23298,N_22194);
or UO_2386 (O_2386,N_23928,N_24425);
nor UO_2387 (O_2387,N_20535,N_22443);
xnor UO_2388 (O_2388,N_23407,N_20055);
or UO_2389 (O_2389,N_21573,N_24422);
xor UO_2390 (O_2390,N_20217,N_24811);
and UO_2391 (O_2391,N_22129,N_21112);
or UO_2392 (O_2392,N_23697,N_24087);
or UO_2393 (O_2393,N_21970,N_23096);
xnor UO_2394 (O_2394,N_20775,N_21362);
or UO_2395 (O_2395,N_20347,N_23670);
or UO_2396 (O_2396,N_23503,N_21079);
xnor UO_2397 (O_2397,N_20169,N_23033);
and UO_2398 (O_2398,N_22658,N_21550);
and UO_2399 (O_2399,N_24441,N_20687);
nor UO_2400 (O_2400,N_21146,N_20513);
nor UO_2401 (O_2401,N_24645,N_21328);
xnor UO_2402 (O_2402,N_24609,N_22158);
or UO_2403 (O_2403,N_21682,N_22853);
and UO_2404 (O_2404,N_23463,N_24042);
and UO_2405 (O_2405,N_20798,N_24986);
nor UO_2406 (O_2406,N_21476,N_20893);
nand UO_2407 (O_2407,N_21576,N_20973);
or UO_2408 (O_2408,N_22397,N_24022);
or UO_2409 (O_2409,N_21070,N_20928);
and UO_2410 (O_2410,N_22571,N_22456);
nor UO_2411 (O_2411,N_22632,N_23632);
xor UO_2412 (O_2412,N_21388,N_21307);
nor UO_2413 (O_2413,N_20362,N_20463);
nand UO_2414 (O_2414,N_24309,N_23628);
xor UO_2415 (O_2415,N_21004,N_20192);
or UO_2416 (O_2416,N_24340,N_23766);
nor UO_2417 (O_2417,N_24722,N_22037);
or UO_2418 (O_2418,N_22422,N_20331);
nand UO_2419 (O_2419,N_22140,N_23024);
nor UO_2420 (O_2420,N_24344,N_23468);
or UO_2421 (O_2421,N_24740,N_20425);
and UO_2422 (O_2422,N_23028,N_22359);
nor UO_2423 (O_2423,N_21904,N_22390);
and UO_2424 (O_2424,N_21988,N_20839);
or UO_2425 (O_2425,N_22282,N_22602);
xor UO_2426 (O_2426,N_22590,N_24006);
nand UO_2427 (O_2427,N_22816,N_21886);
xor UO_2428 (O_2428,N_20295,N_22995);
nor UO_2429 (O_2429,N_20291,N_23218);
and UO_2430 (O_2430,N_20293,N_21643);
or UO_2431 (O_2431,N_23797,N_24745);
and UO_2432 (O_2432,N_24844,N_20268);
or UO_2433 (O_2433,N_24405,N_24124);
nand UO_2434 (O_2434,N_20067,N_21599);
xnor UO_2435 (O_2435,N_22871,N_23844);
nand UO_2436 (O_2436,N_23617,N_22762);
nor UO_2437 (O_2437,N_21948,N_22495);
or UO_2438 (O_2438,N_22862,N_22301);
nand UO_2439 (O_2439,N_24842,N_24029);
nor UO_2440 (O_2440,N_21106,N_24144);
or UO_2441 (O_2441,N_22055,N_24752);
nand UO_2442 (O_2442,N_23006,N_22936);
nor UO_2443 (O_2443,N_24992,N_23709);
nand UO_2444 (O_2444,N_23338,N_24814);
xor UO_2445 (O_2445,N_22186,N_22913);
xor UO_2446 (O_2446,N_24338,N_24430);
and UO_2447 (O_2447,N_24230,N_21779);
or UO_2448 (O_2448,N_21253,N_23786);
nand UO_2449 (O_2449,N_21210,N_22002);
nand UO_2450 (O_2450,N_23773,N_21371);
and UO_2451 (O_2451,N_24332,N_20451);
xor UO_2452 (O_2452,N_23057,N_22824);
or UO_2453 (O_2453,N_23431,N_20252);
xnor UO_2454 (O_2454,N_24734,N_24005);
and UO_2455 (O_2455,N_22684,N_24883);
xnor UO_2456 (O_2456,N_20784,N_21698);
nand UO_2457 (O_2457,N_22585,N_23454);
xnor UO_2458 (O_2458,N_22885,N_20537);
nand UO_2459 (O_2459,N_20203,N_21313);
nor UO_2460 (O_2460,N_21485,N_20405);
or UO_2461 (O_2461,N_21459,N_21874);
xor UO_2462 (O_2462,N_23099,N_22902);
nand UO_2463 (O_2463,N_20167,N_20899);
and UO_2464 (O_2464,N_23232,N_24520);
nand UO_2465 (O_2465,N_24658,N_21754);
or UO_2466 (O_2466,N_21541,N_24227);
xnor UO_2467 (O_2467,N_21493,N_20304);
nor UO_2468 (O_2468,N_21170,N_21565);
xor UO_2469 (O_2469,N_23299,N_21001);
nand UO_2470 (O_2470,N_20541,N_24390);
or UO_2471 (O_2471,N_24241,N_21213);
nand UO_2472 (O_2472,N_23638,N_24086);
nor UO_2473 (O_2473,N_22299,N_23850);
nand UO_2474 (O_2474,N_20461,N_22566);
or UO_2475 (O_2475,N_22009,N_20165);
and UO_2476 (O_2476,N_22668,N_23224);
xnor UO_2477 (O_2477,N_22472,N_23137);
nor UO_2478 (O_2478,N_20621,N_24924);
and UO_2479 (O_2479,N_24263,N_24696);
or UO_2480 (O_2480,N_20176,N_21777);
and UO_2481 (O_2481,N_21627,N_22111);
and UO_2482 (O_2482,N_20132,N_24236);
nand UO_2483 (O_2483,N_21695,N_22639);
nor UO_2484 (O_2484,N_21348,N_23326);
nor UO_2485 (O_2485,N_20652,N_21622);
nand UO_2486 (O_2486,N_22548,N_22164);
nand UO_2487 (O_2487,N_21422,N_23032);
nor UO_2488 (O_2488,N_20596,N_23625);
or UO_2489 (O_2489,N_24836,N_20749);
nand UO_2490 (O_2490,N_24485,N_24580);
xnor UO_2491 (O_2491,N_22921,N_22546);
nor UO_2492 (O_2492,N_20675,N_24385);
or UO_2493 (O_2493,N_22167,N_20983);
xor UO_2494 (O_2494,N_22930,N_20312);
xor UO_2495 (O_2495,N_24066,N_21151);
xor UO_2496 (O_2496,N_24295,N_23776);
nand UO_2497 (O_2497,N_22667,N_20321);
or UO_2498 (O_2498,N_23884,N_21930);
and UO_2499 (O_2499,N_21104,N_22860);
nor UO_2500 (O_2500,N_23111,N_20893);
nor UO_2501 (O_2501,N_23223,N_20381);
and UO_2502 (O_2502,N_23300,N_23547);
and UO_2503 (O_2503,N_22936,N_20813);
xnor UO_2504 (O_2504,N_20573,N_24168);
or UO_2505 (O_2505,N_21305,N_21861);
nand UO_2506 (O_2506,N_24590,N_21392);
xnor UO_2507 (O_2507,N_20730,N_20533);
or UO_2508 (O_2508,N_21958,N_22137);
nand UO_2509 (O_2509,N_21335,N_22932);
nand UO_2510 (O_2510,N_24691,N_22220);
nand UO_2511 (O_2511,N_20262,N_20385);
and UO_2512 (O_2512,N_22509,N_23124);
xnor UO_2513 (O_2513,N_20669,N_24159);
and UO_2514 (O_2514,N_24813,N_23423);
xor UO_2515 (O_2515,N_21928,N_22427);
nand UO_2516 (O_2516,N_23973,N_22060);
xnor UO_2517 (O_2517,N_21561,N_21133);
and UO_2518 (O_2518,N_24464,N_21170);
or UO_2519 (O_2519,N_23968,N_23138);
and UO_2520 (O_2520,N_20743,N_22119);
and UO_2521 (O_2521,N_24591,N_21944);
xor UO_2522 (O_2522,N_24159,N_22229);
or UO_2523 (O_2523,N_24630,N_22979);
and UO_2524 (O_2524,N_22503,N_24134);
or UO_2525 (O_2525,N_24328,N_23240);
and UO_2526 (O_2526,N_21361,N_24016);
and UO_2527 (O_2527,N_21709,N_20375);
xor UO_2528 (O_2528,N_20091,N_22538);
and UO_2529 (O_2529,N_24522,N_22457);
and UO_2530 (O_2530,N_23079,N_23516);
or UO_2531 (O_2531,N_20163,N_22397);
nor UO_2532 (O_2532,N_24809,N_22053);
and UO_2533 (O_2533,N_24511,N_22905);
and UO_2534 (O_2534,N_21350,N_24273);
and UO_2535 (O_2535,N_22041,N_20588);
and UO_2536 (O_2536,N_24768,N_23385);
xnor UO_2537 (O_2537,N_22044,N_24116);
xor UO_2538 (O_2538,N_23606,N_20006);
or UO_2539 (O_2539,N_21147,N_20304);
nand UO_2540 (O_2540,N_22056,N_21738);
or UO_2541 (O_2541,N_21745,N_20539);
and UO_2542 (O_2542,N_21006,N_22141);
xor UO_2543 (O_2543,N_20092,N_21493);
xor UO_2544 (O_2544,N_23470,N_22048);
nand UO_2545 (O_2545,N_22431,N_21993);
nor UO_2546 (O_2546,N_22905,N_23374);
xor UO_2547 (O_2547,N_22301,N_24894);
and UO_2548 (O_2548,N_20986,N_22864);
or UO_2549 (O_2549,N_22686,N_24111);
nor UO_2550 (O_2550,N_23243,N_20545);
xnor UO_2551 (O_2551,N_21034,N_22365);
or UO_2552 (O_2552,N_24874,N_22540);
nor UO_2553 (O_2553,N_23894,N_22677);
xor UO_2554 (O_2554,N_24267,N_24472);
and UO_2555 (O_2555,N_23420,N_21783);
nor UO_2556 (O_2556,N_23537,N_22251);
and UO_2557 (O_2557,N_21936,N_20030);
nand UO_2558 (O_2558,N_21119,N_21675);
nand UO_2559 (O_2559,N_21440,N_23970);
nand UO_2560 (O_2560,N_20825,N_21628);
xor UO_2561 (O_2561,N_24532,N_21595);
xor UO_2562 (O_2562,N_22343,N_22358);
and UO_2563 (O_2563,N_21690,N_23381);
nor UO_2564 (O_2564,N_21246,N_22841);
and UO_2565 (O_2565,N_20924,N_23625);
and UO_2566 (O_2566,N_20318,N_23537);
and UO_2567 (O_2567,N_21066,N_23219);
xnor UO_2568 (O_2568,N_20291,N_20678);
nor UO_2569 (O_2569,N_24622,N_23888);
nand UO_2570 (O_2570,N_24525,N_21432);
xnor UO_2571 (O_2571,N_21721,N_22250);
and UO_2572 (O_2572,N_22525,N_23666);
or UO_2573 (O_2573,N_24122,N_21268);
nand UO_2574 (O_2574,N_23818,N_20142);
nand UO_2575 (O_2575,N_20188,N_21370);
nor UO_2576 (O_2576,N_20489,N_23973);
and UO_2577 (O_2577,N_23932,N_21618);
nand UO_2578 (O_2578,N_23096,N_23587);
xor UO_2579 (O_2579,N_21487,N_22481);
nor UO_2580 (O_2580,N_22244,N_21001);
or UO_2581 (O_2581,N_20310,N_22584);
nand UO_2582 (O_2582,N_24249,N_22747);
and UO_2583 (O_2583,N_23262,N_21341);
nor UO_2584 (O_2584,N_20530,N_22752);
nand UO_2585 (O_2585,N_22413,N_20320);
nand UO_2586 (O_2586,N_24887,N_20915);
or UO_2587 (O_2587,N_24834,N_21361);
xor UO_2588 (O_2588,N_21485,N_21661);
nor UO_2589 (O_2589,N_22490,N_23972);
xor UO_2590 (O_2590,N_23302,N_23938);
and UO_2591 (O_2591,N_22864,N_22521);
or UO_2592 (O_2592,N_21883,N_22454);
and UO_2593 (O_2593,N_22361,N_24488);
nor UO_2594 (O_2594,N_22083,N_23536);
xor UO_2595 (O_2595,N_22941,N_22891);
nand UO_2596 (O_2596,N_23557,N_21066);
or UO_2597 (O_2597,N_24194,N_24881);
nor UO_2598 (O_2598,N_24061,N_20586);
and UO_2599 (O_2599,N_21119,N_20290);
or UO_2600 (O_2600,N_21133,N_20780);
nor UO_2601 (O_2601,N_21012,N_22778);
nand UO_2602 (O_2602,N_20256,N_24234);
and UO_2603 (O_2603,N_21477,N_20519);
nor UO_2604 (O_2604,N_22154,N_20426);
xor UO_2605 (O_2605,N_22757,N_22290);
nand UO_2606 (O_2606,N_24140,N_23068);
and UO_2607 (O_2607,N_20731,N_22431);
or UO_2608 (O_2608,N_20495,N_20665);
or UO_2609 (O_2609,N_21542,N_23623);
xor UO_2610 (O_2610,N_21204,N_20485);
or UO_2611 (O_2611,N_21088,N_20231);
xnor UO_2612 (O_2612,N_21419,N_24306);
and UO_2613 (O_2613,N_24979,N_22163);
nand UO_2614 (O_2614,N_24819,N_21525);
or UO_2615 (O_2615,N_23681,N_20748);
xor UO_2616 (O_2616,N_23490,N_24678);
xnor UO_2617 (O_2617,N_24558,N_21267);
xnor UO_2618 (O_2618,N_21302,N_20135);
nor UO_2619 (O_2619,N_21909,N_20645);
xor UO_2620 (O_2620,N_24400,N_24654);
and UO_2621 (O_2621,N_22017,N_21220);
and UO_2622 (O_2622,N_21866,N_21246);
nand UO_2623 (O_2623,N_23917,N_24665);
or UO_2624 (O_2624,N_22789,N_23297);
and UO_2625 (O_2625,N_24753,N_21702);
nand UO_2626 (O_2626,N_21636,N_20539);
or UO_2627 (O_2627,N_23866,N_24476);
nor UO_2628 (O_2628,N_22980,N_23004);
nand UO_2629 (O_2629,N_23920,N_24234);
xnor UO_2630 (O_2630,N_24309,N_22974);
and UO_2631 (O_2631,N_20818,N_24515);
nor UO_2632 (O_2632,N_22985,N_24871);
xnor UO_2633 (O_2633,N_20650,N_22449);
and UO_2634 (O_2634,N_22425,N_24194);
or UO_2635 (O_2635,N_21545,N_24192);
or UO_2636 (O_2636,N_23476,N_22883);
and UO_2637 (O_2637,N_23856,N_22019);
nand UO_2638 (O_2638,N_24165,N_23693);
and UO_2639 (O_2639,N_20406,N_23832);
nand UO_2640 (O_2640,N_22191,N_21336);
xor UO_2641 (O_2641,N_24872,N_24495);
and UO_2642 (O_2642,N_24392,N_20990);
nor UO_2643 (O_2643,N_24550,N_20664);
xnor UO_2644 (O_2644,N_24067,N_21661);
nor UO_2645 (O_2645,N_21513,N_22225);
nand UO_2646 (O_2646,N_24323,N_20389);
nor UO_2647 (O_2647,N_23694,N_22008);
or UO_2648 (O_2648,N_22488,N_20369);
nand UO_2649 (O_2649,N_23435,N_22099);
xnor UO_2650 (O_2650,N_21879,N_21148);
xor UO_2651 (O_2651,N_21204,N_21790);
nand UO_2652 (O_2652,N_21877,N_23710);
nand UO_2653 (O_2653,N_20062,N_20648);
nor UO_2654 (O_2654,N_23879,N_21492);
nand UO_2655 (O_2655,N_23064,N_22254);
and UO_2656 (O_2656,N_24840,N_21588);
nor UO_2657 (O_2657,N_20146,N_21022);
nor UO_2658 (O_2658,N_21290,N_20160);
nand UO_2659 (O_2659,N_23851,N_22858);
and UO_2660 (O_2660,N_23473,N_20304);
nor UO_2661 (O_2661,N_22743,N_24452);
nand UO_2662 (O_2662,N_23676,N_20342);
or UO_2663 (O_2663,N_21084,N_20881);
nor UO_2664 (O_2664,N_21805,N_20871);
and UO_2665 (O_2665,N_22758,N_21228);
nor UO_2666 (O_2666,N_21418,N_22581);
and UO_2667 (O_2667,N_20483,N_23701);
nand UO_2668 (O_2668,N_24194,N_23247);
nor UO_2669 (O_2669,N_21573,N_22915);
and UO_2670 (O_2670,N_24613,N_24869);
or UO_2671 (O_2671,N_22631,N_22539);
nand UO_2672 (O_2672,N_23292,N_20585);
nor UO_2673 (O_2673,N_24718,N_20904);
xor UO_2674 (O_2674,N_21469,N_22653);
nor UO_2675 (O_2675,N_23554,N_20759);
or UO_2676 (O_2676,N_20260,N_22157);
nor UO_2677 (O_2677,N_24583,N_21378);
and UO_2678 (O_2678,N_24640,N_23803);
nand UO_2679 (O_2679,N_22341,N_22498);
nor UO_2680 (O_2680,N_20782,N_24358);
and UO_2681 (O_2681,N_23998,N_24528);
nand UO_2682 (O_2682,N_24473,N_21695);
nand UO_2683 (O_2683,N_21104,N_24585);
nand UO_2684 (O_2684,N_23424,N_24700);
and UO_2685 (O_2685,N_23240,N_22477);
xnor UO_2686 (O_2686,N_24223,N_24169);
xnor UO_2687 (O_2687,N_22517,N_23041);
or UO_2688 (O_2688,N_23890,N_21849);
or UO_2689 (O_2689,N_23289,N_21243);
and UO_2690 (O_2690,N_24660,N_22181);
nand UO_2691 (O_2691,N_22983,N_21414);
and UO_2692 (O_2692,N_20650,N_24728);
and UO_2693 (O_2693,N_22967,N_22213);
and UO_2694 (O_2694,N_20401,N_21690);
or UO_2695 (O_2695,N_23459,N_20192);
or UO_2696 (O_2696,N_20863,N_20496);
nor UO_2697 (O_2697,N_21494,N_22005);
and UO_2698 (O_2698,N_20107,N_23568);
and UO_2699 (O_2699,N_24464,N_23661);
or UO_2700 (O_2700,N_23091,N_24104);
or UO_2701 (O_2701,N_24512,N_24853);
or UO_2702 (O_2702,N_21792,N_23321);
nor UO_2703 (O_2703,N_23917,N_22220);
or UO_2704 (O_2704,N_21358,N_21597);
nand UO_2705 (O_2705,N_20932,N_20828);
or UO_2706 (O_2706,N_20580,N_24238);
xnor UO_2707 (O_2707,N_21708,N_21382);
nand UO_2708 (O_2708,N_23452,N_24044);
nand UO_2709 (O_2709,N_20883,N_24766);
and UO_2710 (O_2710,N_20062,N_24293);
nor UO_2711 (O_2711,N_24496,N_21121);
or UO_2712 (O_2712,N_20340,N_23047);
or UO_2713 (O_2713,N_20236,N_24463);
xor UO_2714 (O_2714,N_24341,N_21766);
xor UO_2715 (O_2715,N_23852,N_24304);
xor UO_2716 (O_2716,N_22044,N_22142);
nand UO_2717 (O_2717,N_20183,N_23831);
xor UO_2718 (O_2718,N_21080,N_20893);
nand UO_2719 (O_2719,N_21438,N_24228);
and UO_2720 (O_2720,N_20820,N_21852);
nand UO_2721 (O_2721,N_23350,N_20201);
nor UO_2722 (O_2722,N_21640,N_24395);
nand UO_2723 (O_2723,N_24935,N_22448);
xor UO_2724 (O_2724,N_23408,N_22447);
nor UO_2725 (O_2725,N_23945,N_22679);
or UO_2726 (O_2726,N_23983,N_21045);
and UO_2727 (O_2727,N_20187,N_22118);
and UO_2728 (O_2728,N_22138,N_20573);
xnor UO_2729 (O_2729,N_20161,N_21415);
or UO_2730 (O_2730,N_21417,N_23201);
and UO_2731 (O_2731,N_20152,N_24078);
nand UO_2732 (O_2732,N_20666,N_24489);
and UO_2733 (O_2733,N_21727,N_22197);
or UO_2734 (O_2734,N_20867,N_21112);
nor UO_2735 (O_2735,N_22891,N_21700);
or UO_2736 (O_2736,N_23597,N_21960);
nand UO_2737 (O_2737,N_22337,N_20217);
nor UO_2738 (O_2738,N_24693,N_22664);
and UO_2739 (O_2739,N_21897,N_23828);
and UO_2740 (O_2740,N_23625,N_23576);
or UO_2741 (O_2741,N_22147,N_24501);
nor UO_2742 (O_2742,N_22530,N_21956);
xor UO_2743 (O_2743,N_21165,N_23467);
nor UO_2744 (O_2744,N_23826,N_24482);
nor UO_2745 (O_2745,N_20980,N_23623);
or UO_2746 (O_2746,N_23456,N_21605);
xnor UO_2747 (O_2747,N_21250,N_24698);
nand UO_2748 (O_2748,N_22657,N_24221);
or UO_2749 (O_2749,N_21322,N_20621);
nor UO_2750 (O_2750,N_22406,N_24876);
nor UO_2751 (O_2751,N_22391,N_21034);
and UO_2752 (O_2752,N_23782,N_20239);
or UO_2753 (O_2753,N_21880,N_24494);
and UO_2754 (O_2754,N_23927,N_22967);
xnor UO_2755 (O_2755,N_22015,N_23896);
or UO_2756 (O_2756,N_21195,N_22144);
xnor UO_2757 (O_2757,N_23650,N_23745);
nand UO_2758 (O_2758,N_20087,N_23093);
or UO_2759 (O_2759,N_24086,N_21534);
or UO_2760 (O_2760,N_24065,N_24531);
or UO_2761 (O_2761,N_21747,N_21796);
or UO_2762 (O_2762,N_20265,N_20958);
nor UO_2763 (O_2763,N_23860,N_22254);
xnor UO_2764 (O_2764,N_22518,N_20230);
nand UO_2765 (O_2765,N_22637,N_23470);
xnor UO_2766 (O_2766,N_22288,N_24239);
nand UO_2767 (O_2767,N_22820,N_22197);
or UO_2768 (O_2768,N_24520,N_21155);
or UO_2769 (O_2769,N_22049,N_21560);
xnor UO_2770 (O_2770,N_23522,N_21638);
and UO_2771 (O_2771,N_20579,N_22422);
nor UO_2772 (O_2772,N_21391,N_20621);
xor UO_2773 (O_2773,N_23626,N_20799);
or UO_2774 (O_2774,N_23510,N_22760);
nor UO_2775 (O_2775,N_22171,N_21346);
and UO_2776 (O_2776,N_20562,N_20418);
or UO_2777 (O_2777,N_21552,N_22286);
or UO_2778 (O_2778,N_24472,N_20194);
or UO_2779 (O_2779,N_21476,N_23899);
nand UO_2780 (O_2780,N_22073,N_20904);
or UO_2781 (O_2781,N_22323,N_21827);
nor UO_2782 (O_2782,N_23140,N_22582);
xor UO_2783 (O_2783,N_23366,N_23370);
nand UO_2784 (O_2784,N_23041,N_24165);
or UO_2785 (O_2785,N_22579,N_22764);
xnor UO_2786 (O_2786,N_20321,N_23510);
nand UO_2787 (O_2787,N_23189,N_22736);
nor UO_2788 (O_2788,N_23867,N_24417);
nor UO_2789 (O_2789,N_22370,N_24406);
and UO_2790 (O_2790,N_23878,N_24288);
or UO_2791 (O_2791,N_23092,N_24127);
or UO_2792 (O_2792,N_20903,N_23696);
nand UO_2793 (O_2793,N_21891,N_20672);
or UO_2794 (O_2794,N_20504,N_22182);
or UO_2795 (O_2795,N_23559,N_21616);
nand UO_2796 (O_2796,N_23813,N_24035);
or UO_2797 (O_2797,N_20315,N_20753);
nand UO_2798 (O_2798,N_24834,N_22521);
xor UO_2799 (O_2799,N_23721,N_23700);
xnor UO_2800 (O_2800,N_22386,N_20127);
nand UO_2801 (O_2801,N_21140,N_24536);
or UO_2802 (O_2802,N_22147,N_21309);
and UO_2803 (O_2803,N_24825,N_24011);
xor UO_2804 (O_2804,N_24503,N_24996);
nand UO_2805 (O_2805,N_23855,N_23028);
nor UO_2806 (O_2806,N_22386,N_24864);
xor UO_2807 (O_2807,N_20963,N_21664);
or UO_2808 (O_2808,N_21849,N_23150);
and UO_2809 (O_2809,N_24957,N_23589);
nor UO_2810 (O_2810,N_23720,N_23042);
or UO_2811 (O_2811,N_20701,N_20207);
nor UO_2812 (O_2812,N_22952,N_21483);
nand UO_2813 (O_2813,N_21934,N_23124);
nand UO_2814 (O_2814,N_23138,N_23472);
nor UO_2815 (O_2815,N_23995,N_24406);
or UO_2816 (O_2816,N_20916,N_23545);
nor UO_2817 (O_2817,N_20807,N_21736);
and UO_2818 (O_2818,N_23007,N_22352);
or UO_2819 (O_2819,N_23787,N_23551);
and UO_2820 (O_2820,N_22271,N_21443);
and UO_2821 (O_2821,N_24282,N_22639);
xnor UO_2822 (O_2822,N_23202,N_22951);
nor UO_2823 (O_2823,N_22022,N_24909);
and UO_2824 (O_2824,N_24200,N_23063);
nor UO_2825 (O_2825,N_22479,N_23768);
and UO_2826 (O_2826,N_24660,N_23648);
nor UO_2827 (O_2827,N_21363,N_20293);
nand UO_2828 (O_2828,N_24735,N_21546);
xnor UO_2829 (O_2829,N_20178,N_21270);
and UO_2830 (O_2830,N_23563,N_23725);
nand UO_2831 (O_2831,N_22935,N_23774);
nand UO_2832 (O_2832,N_23586,N_21260);
or UO_2833 (O_2833,N_20904,N_24312);
nor UO_2834 (O_2834,N_24895,N_21171);
nand UO_2835 (O_2835,N_22014,N_20942);
or UO_2836 (O_2836,N_22651,N_22100);
xor UO_2837 (O_2837,N_20946,N_24386);
nor UO_2838 (O_2838,N_20404,N_24629);
nand UO_2839 (O_2839,N_20432,N_21562);
nor UO_2840 (O_2840,N_24057,N_20680);
or UO_2841 (O_2841,N_20384,N_20219);
nand UO_2842 (O_2842,N_23721,N_23442);
or UO_2843 (O_2843,N_21773,N_24924);
nand UO_2844 (O_2844,N_22882,N_21164);
and UO_2845 (O_2845,N_23180,N_22961);
nor UO_2846 (O_2846,N_21199,N_22049);
and UO_2847 (O_2847,N_21646,N_24424);
xor UO_2848 (O_2848,N_22794,N_22085);
and UO_2849 (O_2849,N_21108,N_21991);
nor UO_2850 (O_2850,N_24462,N_23846);
and UO_2851 (O_2851,N_23123,N_21663);
nand UO_2852 (O_2852,N_21677,N_20691);
nor UO_2853 (O_2853,N_21636,N_21172);
nand UO_2854 (O_2854,N_22908,N_24861);
and UO_2855 (O_2855,N_20891,N_24805);
nor UO_2856 (O_2856,N_21158,N_24333);
or UO_2857 (O_2857,N_21470,N_24421);
or UO_2858 (O_2858,N_24895,N_22032);
nand UO_2859 (O_2859,N_21510,N_24613);
nand UO_2860 (O_2860,N_22011,N_21040);
nand UO_2861 (O_2861,N_23197,N_20963);
or UO_2862 (O_2862,N_21576,N_23659);
nand UO_2863 (O_2863,N_22077,N_24434);
or UO_2864 (O_2864,N_20755,N_21513);
and UO_2865 (O_2865,N_20045,N_23997);
nand UO_2866 (O_2866,N_22711,N_24053);
and UO_2867 (O_2867,N_21001,N_20814);
and UO_2868 (O_2868,N_22401,N_22455);
or UO_2869 (O_2869,N_23649,N_20502);
or UO_2870 (O_2870,N_21793,N_22524);
xnor UO_2871 (O_2871,N_23568,N_20289);
nand UO_2872 (O_2872,N_24821,N_22766);
or UO_2873 (O_2873,N_24732,N_24639);
and UO_2874 (O_2874,N_23678,N_21231);
nor UO_2875 (O_2875,N_24166,N_23433);
nand UO_2876 (O_2876,N_20614,N_20644);
or UO_2877 (O_2877,N_24666,N_22746);
xor UO_2878 (O_2878,N_23741,N_22887);
nand UO_2879 (O_2879,N_22072,N_23787);
nand UO_2880 (O_2880,N_22434,N_23573);
xor UO_2881 (O_2881,N_23104,N_21626);
or UO_2882 (O_2882,N_23962,N_24591);
nand UO_2883 (O_2883,N_21830,N_21617);
or UO_2884 (O_2884,N_20481,N_20011);
nand UO_2885 (O_2885,N_22168,N_24175);
nor UO_2886 (O_2886,N_20553,N_20988);
and UO_2887 (O_2887,N_24950,N_21034);
nor UO_2888 (O_2888,N_20179,N_24471);
xor UO_2889 (O_2889,N_22224,N_22387);
nand UO_2890 (O_2890,N_20904,N_24752);
xnor UO_2891 (O_2891,N_24854,N_22787);
nand UO_2892 (O_2892,N_21624,N_20871);
xor UO_2893 (O_2893,N_21070,N_23349);
nor UO_2894 (O_2894,N_22549,N_23901);
xor UO_2895 (O_2895,N_23116,N_22716);
nand UO_2896 (O_2896,N_24437,N_23275);
xor UO_2897 (O_2897,N_21959,N_23522);
xor UO_2898 (O_2898,N_22311,N_21559);
nand UO_2899 (O_2899,N_22650,N_24146);
nor UO_2900 (O_2900,N_24452,N_23648);
nand UO_2901 (O_2901,N_23648,N_24231);
nand UO_2902 (O_2902,N_22695,N_23037);
nand UO_2903 (O_2903,N_23601,N_24973);
nor UO_2904 (O_2904,N_22543,N_24883);
or UO_2905 (O_2905,N_24222,N_21253);
nand UO_2906 (O_2906,N_20977,N_24971);
and UO_2907 (O_2907,N_22904,N_22151);
or UO_2908 (O_2908,N_20066,N_20242);
xor UO_2909 (O_2909,N_22185,N_21286);
nand UO_2910 (O_2910,N_20759,N_22475);
nor UO_2911 (O_2911,N_22996,N_20333);
or UO_2912 (O_2912,N_20640,N_21098);
nand UO_2913 (O_2913,N_22445,N_24371);
and UO_2914 (O_2914,N_23234,N_24650);
or UO_2915 (O_2915,N_20427,N_22897);
and UO_2916 (O_2916,N_24734,N_21413);
xnor UO_2917 (O_2917,N_24718,N_20933);
or UO_2918 (O_2918,N_20552,N_22502);
nand UO_2919 (O_2919,N_20022,N_24594);
nand UO_2920 (O_2920,N_23574,N_21235);
and UO_2921 (O_2921,N_23814,N_20381);
xor UO_2922 (O_2922,N_20537,N_21631);
nor UO_2923 (O_2923,N_24085,N_20637);
and UO_2924 (O_2924,N_21083,N_23975);
or UO_2925 (O_2925,N_22081,N_20296);
nor UO_2926 (O_2926,N_20785,N_24413);
or UO_2927 (O_2927,N_21098,N_21173);
nor UO_2928 (O_2928,N_24585,N_20369);
and UO_2929 (O_2929,N_20463,N_20442);
and UO_2930 (O_2930,N_20413,N_24912);
nand UO_2931 (O_2931,N_21854,N_22535);
xnor UO_2932 (O_2932,N_22899,N_21159);
nor UO_2933 (O_2933,N_21818,N_24474);
nand UO_2934 (O_2934,N_24065,N_23812);
and UO_2935 (O_2935,N_21327,N_21809);
nand UO_2936 (O_2936,N_24520,N_24805);
or UO_2937 (O_2937,N_22673,N_23211);
and UO_2938 (O_2938,N_24138,N_24440);
or UO_2939 (O_2939,N_22282,N_21791);
or UO_2940 (O_2940,N_22173,N_22533);
or UO_2941 (O_2941,N_24961,N_21264);
nor UO_2942 (O_2942,N_22683,N_24116);
nand UO_2943 (O_2943,N_23864,N_20723);
or UO_2944 (O_2944,N_23342,N_24311);
and UO_2945 (O_2945,N_22932,N_22632);
xor UO_2946 (O_2946,N_22211,N_20732);
nor UO_2947 (O_2947,N_22166,N_24189);
nand UO_2948 (O_2948,N_22308,N_23939);
nand UO_2949 (O_2949,N_21566,N_20236);
nor UO_2950 (O_2950,N_24360,N_20385);
and UO_2951 (O_2951,N_21986,N_21744);
nand UO_2952 (O_2952,N_23948,N_23251);
xor UO_2953 (O_2953,N_22761,N_24048);
and UO_2954 (O_2954,N_23142,N_20015);
nand UO_2955 (O_2955,N_24970,N_21588);
and UO_2956 (O_2956,N_22988,N_24823);
xnor UO_2957 (O_2957,N_22978,N_23001);
and UO_2958 (O_2958,N_22563,N_24225);
or UO_2959 (O_2959,N_22395,N_24605);
nand UO_2960 (O_2960,N_21093,N_23965);
or UO_2961 (O_2961,N_24875,N_23797);
and UO_2962 (O_2962,N_23814,N_23086);
nand UO_2963 (O_2963,N_22409,N_24557);
xor UO_2964 (O_2964,N_20681,N_20740);
or UO_2965 (O_2965,N_20873,N_22385);
xnor UO_2966 (O_2966,N_24366,N_22430);
nand UO_2967 (O_2967,N_20529,N_23753);
and UO_2968 (O_2968,N_22441,N_24846);
xnor UO_2969 (O_2969,N_22370,N_24703);
and UO_2970 (O_2970,N_20564,N_22774);
xnor UO_2971 (O_2971,N_20430,N_23372);
nor UO_2972 (O_2972,N_24264,N_23779);
nand UO_2973 (O_2973,N_22078,N_22702);
or UO_2974 (O_2974,N_21987,N_23222);
xor UO_2975 (O_2975,N_20977,N_24578);
or UO_2976 (O_2976,N_21947,N_20897);
and UO_2977 (O_2977,N_23719,N_24951);
nor UO_2978 (O_2978,N_24296,N_20052);
xnor UO_2979 (O_2979,N_21660,N_24224);
nand UO_2980 (O_2980,N_24000,N_21990);
xnor UO_2981 (O_2981,N_20773,N_20435);
xnor UO_2982 (O_2982,N_20634,N_22942);
nor UO_2983 (O_2983,N_20463,N_20229);
and UO_2984 (O_2984,N_20111,N_22845);
nor UO_2985 (O_2985,N_24902,N_23378);
nand UO_2986 (O_2986,N_20636,N_24061);
or UO_2987 (O_2987,N_22281,N_21023);
nor UO_2988 (O_2988,N_20436,N_23749);
and UO_2989 (O_2989,N_22178,N_22343);
nand UO_2990 (O_2990,N_24344,N_20575);
and UO_2991 (O_2991,N_22932,N_21526);
and UO_2992 (O_2992,N_21000,N_21983);
nand UO_2993 (O_2993,N_23553,N_24034);
xor UO_2994 (O_2994,N_22272,N_23488);
and UO_2995 (O_2995,N_24610,N_24869);
nand UO_2996 (O_2996,N_23338,N_23264);
or UO_2997 (O_2997,N_20461,N_21458);
nand UO_2998 (O_2998,N_23847,N_22650);
xnor UO_2999 (O_2999,N_20556,N_21776);
endmodule