module basic_750_5000_1000_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_158,In_87);
or U1 (N_1,In_653,In_678);
or U2 (N_2,In_530,In_580);
nor U3 (N_3,In_371,In_14);
nand U4 (N_4,In_132,In_350);
or U5 (N_5,In_322,In_232);
nand U6 (N_6,In_298,In_253);
nor U7 (N_7,In_695,In_306);
and U8 (N_8,In_712,In_53);
or U9 (N_9,In_157,In_370);
nor U10 (N_10,In_6,In_195);
nand U11 (N_11,In_134,In_10);
xor U12 (N_12,In_86,In_403);
or U13 (N_13,In_553,In_171);
nor U14 (N_14,In_428,In_409);
and U15 (N_15,In_739,In_286);
and U16 (N_16,In_681,In_209);
xor U17 (N_17,In_542,In_565);
or U18 (N_18,In_235,In_315);
xnor U19 (N_19,In_360,In_1);
nor U20 (N_20,In_183,In_198);
xor U21 (N_21,In_321,In_36);
nand U22 (N_22,In_163,In_303);
nor U23 (N_23,In_486,In_213);
nor U24 (N_24,In_261,In_52);
nor U25 (N_25,In_452,In_622);
and U26 (N_26,In_71,In_7);
xor U27 (N_27,In_265,In_337);
xor U28 (N_28,In_494,In_423);
or U29 (N_29,In_586,In_335);
nand U30 (N_30,In_118,In_400);
and U31 (N_31,In_109,In_462);
xor U32 (N_32,In_473,In_546);
nand U33 (N_33,In_281,In_573);
nor U34 (N_34,In_351,In_356);
xor U35 (N_35,In_46,In_741);
xor U36 (N_36,In_187,In_254);
and U37 (N_37,In_567,In_655);
and U38 (N_38,In_675,In_59);
nor U39 (N_39,In_266,In_419);
nor U40 (N_40,In_644,In_556);
xnor U41 (N_41,In_463,In_51);
nand U42 (N_42,In_693,In_67);
nor U43 (N_43,In_152,In_402);
nor U44 (N_44,In_203,In_683);
and U45 (N_45,In_455,In_141);
or U46 (N_46,In_0,In_294);
or U47 (N_47,In_363,In_173);
or U48 (N_48,In_318,In_628);
or U49 (N_49,In_40,In_606);
and U50 (N_50,In_420,In_483);
nand U51 (N_51,In_398,In_588);
xnor U52 (N_52,In_456,In_305);
or U53 (N_53,In_710,In_373);
xnor U54 (N_54,In_296,In_627);
xnor U55 (N_55,In_507,In_746);
and U56 (N_56,In_139,In_295);
nor U57 (N_57,In_642,In_312);
nand U58 (N_58,In_110,In_93);
or U59 (N_59,In_368,In_285);
xor U60 (N_60,In_633,In_529);
or U61 (N_61,In_526,In_668);
nand U62 (N_62,In_416,In_411);
or U63 (N_63,In_242,In_449);
nor U64 (N_64,In_524,In_90);
and U65 (N_65,In_430,In_276);
and U66 (N_66,In_537,In_649);
nor U67 (N_67,In_278,In_592);
nand U68 (N_68,In_601,In_220);
and U69 (N_69,In_367,In_170);
nand U70 (N_70,In_11,In_98);
nand U71 (N_71,In_17,In_178);
nor U72 (N_72,In_260,In_585);
xnor U73 (N_73,In_311,In_397);
or U74 (N_74,In_83,In_582);
nand U75 (N_75,In_650,In_421);
xor U76 (N_76,In_221,In_167);
nand U77 (N_77,In_172,In_735);
nor U78 (N_78,In_268,In_418);
nor U79 (N_79,In_20,In_366);
or U80 (N_80,In_690,In_636);
nor U81 (N_81,In_129,In_2);
or U82 (N_82,In_682,In_116);
and U83 (N_83,In_37,In_89);
or U84 (N_84,In_245,In_273);
nand U85 (N_85,In_702,In_747);
nand U86 (N_86,In_234,In_517);
and U87 (N_87,In_694,In_262);
or U88 (N_88,In_660,In_279);
or U89 (N_89,In_16,In_503);
xor U90 (N_90,In_280,In_113);
nor U91 (N_91,In_436,In_344);
nand U92 (N_92,In_443,In_307);
and U93 (N_93,In_9,In_659);
xnor U94 (N_94,In_414,In_560);
nand U95 (N_95,In_640,In_676);
or U96 (N_96,In_346,In_597);
or U97 (N_97,In_404,In_239);
xor U98 (N_98,In_127,In_70);
nand U99 (N_99,In_26,In_251);
nand U100 (N_100,In_643,In_388);
nand U101 (N_101,In_248,In_444);
xor U102 (N_102,In_202,In_658);
or U103 (N_103,In_32,In_97);
nor U104 (N_104,N_58,In_680);
nor U105 (N_105,In_533,In_447);
xor U106 (N_106,In_50,In_527);
nand U107 (N_107,In_484,In_108);
or U108 (N_108,In_323,In_563);
and U109 (N_109,N_43,N_96);
or U110 (N_110,In_618,In_457);
and U111 (N_111,In_629,In_184);
nand U112 (N_112,N_15,In_107);
xnor U113 (N_113,In_561,In_258);
or U114 (N_114,In_128,In_723);
xnor U115 (N_115,In_410,In_392);
nor U116 (N_116,In_684,In_75);
and U117 (N_117,In_464,In_200);
nor U118 (N_118,In_39,In_510);
or U119 (N_119,In_282,In_631);
xor U120 (N_120,In_379,In_44);
and U121 (N_121,In_393,In_619);
or U122 (N_122,In_230,In_748);
xnor U123 (N_123,In_413,N_52);
xor U124 (N_124,In_308,In_732);
xor U125 (N_125,In_144,In_64);
xor U126 (N_126,N_11,N_90);
nand U127 (N_127,In_730,In_309);
or U128 (N_128,In_362,In_233);
nor U129 (N_129,In_38,In_332);
xnor U130 (N_130,In_646,In_709);
xnor U131 (N_131,In_607,N_74);
or U132 (N_132,In_255,In_632);
nand U133 (N_133,In_274,In_155);
nor U134 (N_134,In_704,In_28);
nand U135 (N_135,In_523,In_181);
nand U136 (N_136,N_9,N_67);
and U137 (N_137,In_288,In_13);
xnor U138 (N_138,In_243,In_249);
or U139 (N_139,N_79,In_283);
or U140 (N_140,In_117,In_737);
and U141 (N_141,In_501,In_445);
xor U142 (N_142,In_609,In_571);
nor U143 (N_143,In_626,In_199);
xor U144 (N_144,In_513,In_499);
and U145 (N_145,In_734,In_551);
xor U146 (N_146,In_478,In_347);
nand U147 (N_147,In_426,N_72);
nand U148 (N_148,N_17,In_505);
or U149 (N_149,N_23,In_512);
xor U150 (N_150,In_91,In_314);
and U151 (N_151,In_106,In_8);
and U152 (N_152,In_204,In_453);
and U153 (N_153,In_733,N_34);
nand U154 (N_154,In_361,N_95);
xnor U155 (N_155,In_349,In_461);
nor U156 (N_156,In_685,In_381);
or U157 (N_157,In_591,In_480);
and U158 (N_158,In_621,In_558);
and U159 (N_159,In_256,In_319);
or U160 (N_160,In_99,N_83);
and U161 (N_161,In_96,In_692);
xnor U162 (N_162,In_49,In_131);
or U163 (N_163,N_77,N_30);
nand U164 (N_164,In_688,In_497);
xor U165 (N_165,In_339,In_728);
or U166 (N_166,In_435,N_61);
xnor U167 (N_167,N_63,In_674);
nand U168 (N_168,In_481,In_603);
nor U169 (N_169,In_544,In_566);
xor U170 (N_170,N_80,In_667);
nor U171 (N_171,In_670,N_62);
and U172 (N_172,In_55,In_612);
nor U173 (N_173,In_577,In_531);
nand U174 (N_174,In_196,In_661);
nand U175 (N_175,In_749,In_472);
or U176 (N_176,In_162,In_210);
nor U177 (N_177,In_433,In_697);
nor U178 (N_178,In_405,N_55);
xor U179 (N_179,In_317,In_550);
xor U180 (N_180,N_47,N_88);
nand U181 (N_181,In_743,In_334);
xnor U182 (N_182,In_652,N_35);
or U183 (N_183,In_500,In_687);
xor U184 (N_184,N_40,In_143);
nor U185 (N_185,In_175,In_384);
nand U186 (N_186,In_431,In_665);
or U187 (N_187,In_194,N_68);
and U188 (N_188,In_145,In_263);
nand U189 (N_189,In_138,In_744);
or U190 (N_190,In_219,In_600);
or U191 (N_191,In_570,In_166);
and U192 (N_192,In_114,In_425);
or U193 (N_193,In_482,In_729);
and U194 (N_194,In_638,In_60);
xor U195 (N_195,In_545,In_630);
nand U196 (N_196,In_564,In_595);
nand U197 (N_197,In_569,In_536);
xnor U198 (N_198,In_345,In_721);
or U199 (N_199,In_460,In_62);
or U200 (N_200,N_183,In_590);
nor U201 (N_201,In_427,N_94);
nand U202 (N_202,N_4,In_669);
or U203 (N_203,In_713,In_76);
xor U204 (N_204,N_166,In_401);
xnor U205 (N_205,In_406,In_31);
and U206 (N_206,In_205,In_519);
xnor U207 (N_207,In_442,In_666);
nor U208 (N_208,N_177,In_664);
xnor U209 (N_209,N_131,In_641);
nand U210 (N_210,N_59,N_7);
xor U211 (N_211,N_110,In_333);
or U212 (N_212,In_58,N_159);
nand U213 (N_213,In_88,In_396);
and U214 (N_214,In_257,In_466);
xnor U215 (N_215,In_727,In_412);
and U216 (N_216,N_101,In_151);
nor U217 (N_217,In_156,In_718);
and U218 (N_218,N_194,N_78);
nor U219 (N_219,In_133,In_583);
nor U220 (N_220,In_73,In_575);
xor U221 (N_221,N_8,N_103);
xnor U222 (N_222,In_725,In_654);
nand U223 (N_223,In_555,N_115);
xor U224 (N_224,In_711,N_13);
nand U225 (N_225,N_36,N_132);
and U226 (N_226,In_57,In_68);
and U227 (N_227,In_521,N_107);
or U228 (N_228,N_111,N_190);
nand U229 (N_229,In_80,In_21);
or U230 (N_230,In_287,In_407);
xnor U231 (N_231,N_117,In_446);
nand U232 (N_232,N_25,In_341);
nand U233 (N_233,In_5,In_61);
or U234 (N_234,In_493,In_532);
xor U235 (N_235,N_152,In_391);
and U236 (N_236,In_515,In_559);
nor U237 (N_237,In_705,In_454);
nor U238 (N_238,N_118,In_225);
or U239 (N_239,In_549,In_95);
xor U240 (N_240,In_415,In_587);
nand U241 (N_241,N_102,In_161);
or U242 (N_242,N_142,N_56);
xor U243 (N_243,N_105,N_6);
nor U244 (N_244,In_543,In_422);
nand U245 (N_245,In_576,In_217);
and U246 (N_246,In_514,In_623);
nand U247 (N_247,In_535,In_488);
xnor U248 (N_248,In_441,In_140);
nor U249 (N_249,N_145,In_700);
xor U250 (N_250,In_635,In_142);
and U251 (N_251,In_338,In_689);
xnor U252 (N_252,N_139,N_185);
nor U253 (N_253,In_706,In_518);
nor U254 (N_254,N_157,N_60);
nor U255 (N_255,N_85,In_19);
xor U256 (N_256,In_496,In_238);
nand U257 (N_257,N_116,In_115);
or U258 (N_258,In_226,N_27);
or U259 (N_259,In_611,N_48);
nor U260 (N_260,In_126,In_111);
and U261 (N_261,In_369,In_105);
xor U262 (N_262,In_364,In_378);
xor U263 (N_263,In_620,In_651);
nor U264 (N_264,N_20,In_72);
nor U265 (N_265,In_374,In_495);
nand U266 (N_266,In_458,N_16);
nor U267 (N_267,In_477,In_214);
nor U268 (N_268,In_672,N_69);
nor U269 (N_269,In_179,In_182);
nor U270 (N_270,In_190,In_291);
xor U271 (N_271,In_568,N_87);
nor U272 (N_272,In_679,In_485);
or U273 (N_273,In_130,In_77);
nor U274 (N_274,In_35,N_189);
or U275 (N_275,N_129,N_89);
xor U276 (N_276,N_192,N_181);
nand U277 (N_277,N_22,N_2);
or U278 (N_278,In_284,In_584);
or U279 (N_279,In_252,In_720);
or U280 (N_280,In_699,N_98);
nor U281 (N_281,In_354,In_336);
xnor U282 (N_282,In_123,In_714);
and U283 (N_283,In_189,N_136);
nor U284 (N_284,In_608,In_185);
nand U285 (N_285,N_184,In_119);
xnor U286 (N_286,In_574,N_76);
xor U287 (N_287,In_313,In_228);
nand U288 (N_288,N_104,In_736);
and U289 (N_289,In_376,In_112);
nand U290 (N_290,In_240,In_717);
nand U291 (N_291,In_662,N_151);
nor U292 (N_292,In_100,N_65);
xor U293 (N_293,In_673,N_156);
and U294 (N_294,In_617,In_432);
or U295 (N_295,In_269,In_293);
xor U296 (N_296,N_46,N_188);
xnor U297 (N_297,N_44,In_65);
nor U298 (N_298,In_353,N_146);
or U299 (N_299,In_491,In_206);
nand U300 (N_300,In_125,In_557);
nand U301 (N_301,In_380,N_71);
xor U302 (N_302,N_242,In_511);
or U303 (N_303,N_70,In_297);
nor U304 (N_304,N_270,In_165);
or U305 (N_305,In_208,N_195);
xor U306 (N_306,N_256,N_128);
nor U307 (N_307,N_263,In_201);
nor U308 (N_308,In_614,In_552);
nand U309 (N_309,N_187,N_237);
and U310 (N_310,In_520,N_285);
or U311 (N_311,N_247,N_209);
nor U312 (N_312,In_48,In_489);
nor U313 (N_313,In_289,In_476);
or U314 (N_314,N_261,In_352);
nor U315 (N_315,N_121,N_228);
nor U316 (N_316,In_325,In_599);
or U317 (N_317,In_277,In_439);
nor U318 (N_318,N_205,N_172);
xor U319 (N_319,N_106,In_434);
or U320 (N_320,In_504,In_541);
xnor U321 (N_321,In_487,N_293);
or U322 (N_322,N_144,In_355);
xnor U323 (N_323,N_229,N_255);
nor U324 (N_324,In_417,In_387);
xor U325 (N_325,N_84,In_372);
and U326 (N_326,In_390,In_18);
nand U327 (N_327,N_119,N_239);
nand U328 (N_328,In_691,N_203);
xor U329 (N_329,In_3,N_86);
and U330 (N_330,N_279,In_331);
nor U331 (N_331,In_191,In_448);
nor U332 (N_332,In_12,N_134);
and U333 (N_333,In_137,N_206);
nor U334 (N_334,In_135,In_327);
nor U335 (N_335,N_26,N_73);
nor U336 (N_336,In_719,In_42);
nand U337 (N_337,In_290,N_100);
or U338 (N_338,In_197,In_740);
xnor U339 (N_339,N_31,In_386);
nand U340 (N_340,N_257,In_85);
or U341 (N_341,In_634,In_54);
nand U342 (N_342,In_359,In_696);
nor U343 (N_343,In_738,In_4);
or U344 (N_344,N_153,In_147);
or U345 (N_345,N_97,N_212);
nor U346 (N_346,In_69,In_176);
or U347 (N_347,N_292,N_141);
or U348 (N_348,N_260,In_304);
xor U349 (N_349,In_223,N_99);
nand U350 (N_350,In_43,N_213);
and U351 (N_351,In_229,N_168);
xor U352 (N_352,In_383,In_159);
or U353 (N_353,N_45,In_731);
nand U354 (N_354,N_114,In_385);
nor U355 (N_355,In_657,N_180);
or U356 (N_356,N_137,N_182);
or U357 (N_357,N_113,In_120);
xor U358 (N_358,N_37,N_286);
or U359 (N_359,N_173,In_222);
and U360 (N_360,N_240,In_365);
nor U361 (N_361,In_465,N_254);
xnor U362 (N_362,In_424,N_224);
or U363 (N_363,N_271,N_296);
nand U364 (N_364,N_92,N_193);
and U365 (N_365,N_29,In_528);
nand U366 (N_366,N_258,N_241);
xnor U367 (N_367,N_186,In_578);
nor U368 (N_368,N_167,N_0);
or U369 (N_369,In_707,In_136);
nor U370 (N_370,N_178,N_298);
nand U371 (N_371,N_171,In_343);
xnor U372 (N_372,In_389,N_273);
and U373 (N_373,In_330,N_295);
nor U374 (N_374,In_701,N_32);
xor U375 (N_375,N_276,In_742);
nor U376 (N_376,N_10,In_146);
or U377 (N_377,In_246,N_266);
xor U378 (N_378,N_109,In_522);
nand U379 (N_379,In_539,In_102);
or U380 (N_380,In_492,In_160);
xor U381 (N_381,In_180,N_154);
xnor U382 (N_382,In_177,In_438);
nor U383 (N_383,In_270,In_272);
and U384 (N_384,In_224,In_437);
xor U385 (N_385,In_540,In_328);
nand U386 (N_386,N_91,In_215);
or U387 (N_387,N_5,N_169);
nor U388 (N_388,N_126,N_75);
and U389 (N_389,N_252,N_28);
xnor U390 (N_390,N_18,N_42);
nand U391 (N_391,N_265,N_112);
nor U392 (N_392,N_197,N_272);
nor U393 (N_393,N_41,N_64);
or U394 (N_394,In_15,In_101);
or U395 (N_395,N_225,In_506);
nand U396 (N_396,In_467,In_148);
xor U397 (N_397,N_290,In_27);
nor U398 (N_398,In_236,N_51);
nor U399 (N_399,N_155,N_289);
nor U400 (N_400,N_356,N_19);
or U401 (N_401,In_340,In_342);
and U402 (N_402,In_244,N_352);
or U403 (N_403,In_192,In_22);
xnor U404 (N_404,In_216,In_218);
xor U405 (N_405,N_367,In_29);
nor U406 (N_406,In_663,N_288);
or U407 (N_407,N_338,In_186);
nand U408 (N_408,In_45,In_698);
and U409 (N_409,N_299,N_323);
or U410 (N_410,In_259,In_598);
xnor U411 (N_411,N_329,N_341);
and U412 (N_412,N_227,N_315);
nor U413 (N_413,In_724,In_271);
xor U414 (N_414,N_311,N_331);
xnor U415 (N_415,In_534,N_396);
nor U416 (N_416,N_327,N_373);
xor U417 (N_417,In_538,In_124);
xnor U418 (N_418,In_648,N_221);
nand U419 (N_419,In_47,N_202);
xnor U420 (N_420,N_243,N_316);
and U421 (N_421,N_303,N_349);
and U422 (N_422,N_382,In_227);
nor U423 (N_423,N_82,In_645);
and U424 (N_424,In_498,In_613);
or U425 (N_425,N_320,N_54);
nor U426 (N_426,N_322,In_329);
nor U427 (N_427,N_222,In_324);
and U428 (N_428,N_380,In_562);
and U429 (N_429,N_370,In_92);
nor U430 (N_430,In_677,In_469);
nor U431 (N_431,N_399,N_278);
nor U432 (N_432,In_84,In_326);
or U433 (N_433,In_479,In_726);
xor U434 (N_434,N_389,In_212);
nand U435 (N_435,N_333,N_210);
nor U436 (N_436,N_371,N_148);
nand U437 (N_437,N_138,In_716);
nand U438 (N_438,In_320,N_302);
nor U439 (N_439,N_305,N_386);
nand U440 (N_440,N_14,N_398);
and U441 (N_441,In_395,In_451);
and U442 (N_442,In_604,N_384);
xor U443 (N_443,N_211,N_281);
or U444 (N_444,N_306,N_348);
or U445 (N_445,In_267,N_163);
xnor U446 (N_446,N_130,In_34);
nand U447 (N_447,N_368,N_334);
or U448 (N_448,N_233,N_140);
nand U449 (N_449,N_264,N_365);
nand U450 (N_450,N_378,In_250);
and U451 (N_451,N_280,N_343);
nand U452 (N_452,N_358,N_223);
or U453 (N_453,N_218,N_354);
xor U454 (N_454,N_108,N_359);
nor U455 (N_455,N_339,N_304);
nor U456 (N_456,N_313,N_360);
xor U457 (N_457,N_385,In_722);
xor U458 (N_458,In_348,N_201);
or U459 (N_459,In_247,N_324);
xor U460 (N_460,N_283,In_399);
nand U461 (N_461,In_122,In_637);
xor U462 (N_462,In_302,In_554);
or U463 (N_463,In_300,In_164);
and U464 (N_464,N_49,In_450);
nor U465 (N_465,In_174,N_309);
nand U466 (N_466,In_375,N_287);
or U467 (N_467,N_149,N_390);
nand U468 (N_468,N_344,In_525);
or U469 (N_469,N_232,In_581);
nor U470 (N_470,N_332,N_238);
nor U471 (N_471,In_94,N_176);
xor U472 (N_472,In_516,N_357);
xnor U473 (N_473,N_214,In_490);
xnor U474 (N_474,N_362,In_188);
nor U475 (N_475,N_387,In_624);
xnor U476 (N_476,N_321,In_616);
or U477 (N_477,N_274,N_207);
or U478 (N_478,In_82,N_196);
and U479 (N_479,N_268,N_124);
and U480 (N_480,N_133,In_316);
and U481 (N_481,N_123,N_248);
nand U482 (N_482,In_193,N_179);
xnor U483 (N_483,In_241,N_164);
nor U484 (N_484,N_250,N_381);
or U485 (N_485,N_24,N_3);
xor U486 (N_486,N_282,In_81);
xnor U487 (N_487,In_231,In_23);
nor U488 (N_488,N_199,N_346);
xnor U489 (N_489,N_395,In_594);
and U490 (N_490,N_200,In_502);
nor U491 (N_491,N_253,In_671);
xnor U492 (N_492,N_297,In_275);
and U493 (N_493,N_291,In_429);
nand U494 (N_494,N_353,N_204);
and U495 (N_495,In_602,N_351);
nor U496 (N_496,In_169,In_74);
or U497 (N_497,N_342,In_647);
nand U498 (N_498,N_317,In_33);
nand U499 (N_499,N_215,N_364);
nand U500 (N_500,N_485,N_337);
xnor U501 (N_501,N_219,N_158);
nand U502 (N_502,N_347,N_127);
or U503 (N_503,In_104,N_463);
or U504 (N_504,N_496,N_401);
xor U505 (N_505,N_444,N_244);
or U506 (N_506,N_477,In_625);
nand U507 (N_507,N_445,In_103);
and U508 (N_508,N_147,In_149);
nor U509 (N_509,N_420,N_405);
nor U510 (N_510,In_56,N_461);
or U511 (N_511,N_437,N_208);
nor U512 (N_512,N_160,In_615);
nand U513 (N_513,N_383,N_165);
nand U514 (N_514,N_234,N_428);
xor U515 (N_515,N_464,N_495);
and U516 (N_516,N_406,N_39);
nand U517 (N_517,In_121,N_361);
xor U518 (N_518,N_415,N_439);
and U519 (N_519,In_686,N_236);
xor U520 (N_520,N_38,N_470);
nor U521 (N_521,N_408,N_220);
or U522 (N_522,N_314,In_41);
and U523 (N_523,N_328,In_656);
nor U524 (N_524,N_424,N_376);
or U525 (N_525,N_394,In_703);
and U526 (N_526,N_269,N_120);
nor U527 (N_527,In_66,N_455);
xor U528 (N_528,N_66,N_436);
nand U529 (N_529,N_404,In_292);
or U530 (N_530,N_475,N_473);
nor U531 (N_531,N_300,N_397);
nand U532 (N_532,In_745,N_417);
nand U533 (N_533,In_593,N_432);
nand U534 (N_534,N_465,N_479);
nand U535 (N_535,In_24,In_79);
nand U536 (N_536,N_478,In_471);
nand U537 (N_537,N_472,N_350);
and U538 (N_538,N_162,N_340);
or U539 (N_539,N_246,In_377);
and U540 (N_540,In_572,In_154);
or U541 (N_541,N_277,N_457);
xor U542 (N_542,N_326,In_264);
or U543 (N_543,In_30,N_427);
nor U544 (N_544,N_57,N_486);
nor U545 (N_545,In_150,In_358);
nand U546 (N_546,N_442,N_499);
and U547 (N_547,N_388,N_458);
xor U548 (N_548,N_336,N_456);
xor U549 (N_549,N_143,In_605);
nand U550 (N_550,N_426,N_391);
nor U551 (N_551,N_369,N_245);
nand U552 (N_552,N_307,N_216);
nor U553 (N_553,In_508,In_299);
or U554 (N_554,In_237,N_122);
and U555 (N_555,N_161,In_715);
nand U556 (N_556,N_423,In_610);
nor U557 (N_557,N_174,In_548);
nor U558 (N_558,In_310,N_251);
nand U559 (N_559,N_355,In_168);
nand U560 (N_560,N_482,N_443);
or U561 (N_561,N_191,N_308);
xnor U562 (N_562,N_462,N_488);
xnor U563 (N_563,In_301,N_446);
nor U564 (N_564,N_217,In_382);
nor U565 (N_565,N_363,N_435);
nor U566 (N_566,N_434,N_431);
or U567 (N_567,In_153,N_325);
and U568 (N_568,N_490,N_440);
xnor U569 (N_569,N_125,N_474);
and U570 (N_570,N_393,N_379);
nand U571 (N_571,N_310,In_579);
nor U572 (N_572,N_480,N_175);
and U573 (N_573,N_447,N_235);
xor U574 (N_574,In_25,N_400);
or U575 (N_575,N_377,N_471);
xor U576 (N_576,N_422,N_469);
nand U577 (N_577,N_452,N_198);
nor U578 (N_578,N_476,N_407);
nand U579 (N_579,N_438,In_596);
nand U580 (N_580,N_21,In_357);
or U581 (N_581,In_207,N_429);
and U582 (N_582,N_453,N_33);
nor U583 (N_583,N_53,N_81);
xor U584 (N_584,N_484,N_319);
nor U585 (N_585,N_284,N_275);
nand U586 (N_586,N_93,In_474);
or U587 (N_587,N_493,N_262);
nor U588 (N_588,N_491,N_409);
nor U589 (N_589,In_78,N_402);
nor U590 (N_590,N_335,N_413);
nand U591 (N_591,N_170,N_441);
nor U592 (N_592,N_454,N_450);
xor U593 (N_593,N_411,In_708);
nor U594 (N_594,N_430,N_318);
or U595 (N_595,N_481,N_412);
nor U596 (N_596,In_509,N_345);
xnor U597 (N_597,In_468,N_249);
nand U598 (N_598,N_135,In_211);
and U599 (N_599,N_451,N_12);
nor U600 (N_600,N_414,N_556);
nand U601 (N_601,N_570,N_585);
xnor U602 (N_602,N_545,N_595);
xor U603 (N_603,N_518,N_567);
or U604 (N_604,N_591,N_392);
or U605 (N_605,N_259,N_460);
or U606 (N_606,N_301,N_433);
and U607 (N_607,N_555,N_231);
xor U608 (N_608,N_468,N_563);
or U609 (N_609,N_593,N_559);
nand U610 (N_610,N_583,N_538);
xnor U611 (N_611,In_639,N_487);
xor U612 (N_612,N_521,N_226);
nand U613 (N_613,N_501,N_230);
nand U614 (N_614,N_554,N_526);
nand U615 (N_615,N_547,N_520);
nand U616 (N_616,N_573,N_528);
nor U617 (N_617,N_535,N_1);
and U618 (N_618,N_543,N_590);
nor U619 (N_619,N_516,N_561);
or U620 (N_620,N_586,N_588);
or U621 (N_621,In_408,N_448);
xnor U622 (N_622,N_574,N_410);
nor U623 (N_623,N_511,N_403);
xnor U624 (N_624,In_589,N_494);
nor U625 (N_625,N_587,N_489);
and U626 (N_626,N_425,N_504);
and U627 (N_627,N_374,N_544);
xnor U628 (N_628,N_421,N_366);
xnor U629 (N_629,N_416,N_575);
nand U630 (N_630,N_571,N_533);
nand U631 (N_631,N_312,N_502);
or U632 (N_632,N_527,In_63);
nand U633 (N_633,N_515,N_580);
nand U634 (N_634,N_550,N_517);
nand U635 (N_635,N_579,N_483);
or U636 (N_636,N_542,N_530);
nor U637 (N_637,N_582,In_440);
or U638 (N_638,N_566,N_534);
nor U639 (N_639,N_507,N_548);
nand U640 (N_640,N_524,N_506);
xor U641 (N_641,In_470,N_597);
nor U642 (N_642,N_525,N_562);
nand U643 (N_643,N_552,N_419);
and U644 (N_644,N_459,N_500);
nand U645 (N_645,In_547,N_565);
nor U646 (N_646,N_514,N_294);
or U647 (N_647,N_449,N_599);
or U648 (N_648,In_394,N_584);
nor U649 (N_649,N_564,N_498);
xnor U650 (N_650,N_513,N_577);
or U651 (N_651,N_569,N_558);
nand U652 (N_652,N_531,N_537);
and U653 (N_653,N_529,In_459);
and U654 (N_654,N_551,N_372);
and U655 (N_655,N_596,N_522);
or U656 (N_656,N_505,N_578);
nor U657 (N_657,N_492,N_467);
xnor U658 (N_658,N_540,N_330);
nor U659 (N_659,N_510,N_572);
and U660 (N_660,In_475,N_267);
and U661 (N_661,N_594,N_509);
or U662 (N_662,N_50,N_576);
and U663 (N_663,N_598,N_546);
and U664 (N_664,N_541,N_418);
nand U665 (N_665,N_549,N_523);
and U666 (N_666,N_375,N_581);
or U667 (N_667,N_560,N_553);
and U668 (N_668,N_592,N_557);
nand U669 (N_669,N_512,N_589);
or U670 (N_670,N_503,N_536);
or U671 (N_671,N_466,N_497);
and U672 (N_672,N_519,N_508);
or U673 (N_673,N_532,N_568);
nor U674 (N_674,N_539,N_150);
xor U675 (N_675,In_470,N_564);
and U676 (N_676,N_503,N_507);
nand U677 (N_677,N_529,N_556);
xor U678 (N_678,N_579,N_150);
nand U679 (N_679,In_470,N_549);
nand U680 (N_680,N_533,N_598);
or U681 (N_681,N_569,N_571);
xnor U682 (N_682,N_519,N_375);
or U683 (N_683,N_583,N_510);
or U684 (N_684,N_538,In_475);
and U685 (N_685,N_392,N_536);
nand U686 (N_686,N_598,N_421);
nor U687 (N_687,N_558,N_575);
nand U688 (N_688,N_513,N_508);
and U689 (N_689,N_559,N_267);
and U690 (N_690,N_414,N_410);
xor U691 (N_691,N_487,N_583);
nor U692 (N_692,N_503,N_526);
nor U693 (N_693,N_526,N_543);
and U694 (N_694,N_468,N_374);
nor U695 (N_695,N_467,N_525);
and U696 (N_696,N_449,N_528);
nor U697 (N_697,N_372,N_532);
and U698 (N_698,N_537,In_470);
and U699 (N_699,N_519,N_448);
or U700 (N_700,N_643,N_647);
xor U701 (N_701,N_686,N_670);
or U702 (N_702,N_622,N_629);
nor U703 (N_703,N_639,N_677);
and U704 (N_704,N_682,N_605);
and U705 (N_705,N_681,N_664);
xnor U706 (N_706,N_633,N_650);
xnor U707 (N_707,N_673,N_691);
xor U708 (N_708,N_678,N_679);
nor U709 (N_709,N_601,N_615);
or U710 (N_710,N_618,N_689);
nor U711 (N_711,N_614,N_602);
xor U712 (N_712,N_687,N_672);
or U713 (N_713,N_646,N_688);
or U714 (N_714,N_669,N_626);
or U715 (N_715,N_655,N_600);
nor U716 (N_716,N_627,N_685);
and U717 (N_717,N_628,N_698);
nand U718 (N_718,N_690,N_607);
nor U719 (N_719,N_638,N_663);
xnor U720 (N_720,N_652,N_620);
nand U721 (N_721,N_699,N_683);
xor U722 (N_722,N_634,N_611);
or U723 (N_723,N_657,N_693);
or U724 (N_724,N_665,N_616);
or U725 (N_725,N_642,N_649);
xnor U726 (N_726,N_624,N_623);
nand U727 (N_727,N_603,N_659);
and U728 (N_728,N_661,N_680);
nand U729 (N_729,N_609,N_658);
nand U730 (N_730,N_676,N_604);
xnor U731 (N_731,N_632,N_625);
xnor U732 (N_732,N_610,N_694);
and U733 (N_733,N_668,N_692);
and U734 (N_734,N_613,N_667);
or U735 (N_735,N_630,N_696);
nor U736 (N_736,N_662,N_641);
and U737 (N_737,N_654,N_644);
and U738 (N_738,N_631,N_645);
or U739 (N_739,N_675,N_635);
xnor U740 (N_740,N_656,N_619);
or U741 (N_741,N_660,N_653);
or U742 (N_742,N_640,N_695);
nor U743 (N_743,N_621,N_606);
or U744 (N_744,N_697,N_617);
and U745 (N_745,N_636,N_637);
and U746 (N_746,N_684,N_648);
xnor U747 (N_747,N_651,N_671);
nor U748 (N_748,N_612,N_666);
nand U749 (N_749,N_608,N_674);
and U750 (N_750,N_659,N_643);
or U751 (N_751,N_622,N_681);
and U752 (N_752,N_697,N_685);
and U753 (N_753,N_651,N_623);
or U754 (N_754,N_683,N_601);
xnor U755 (N_755,N_614,N_656);
nor U756 (N_756,N_613,N_601);
xor U757 (N_757,N_620,N_683);
xnor U758 (N_758,N_695,N_636);
or U759 (N_759,N_679,N_683);
nor U760 (N_760,N_687,N_629);
nand U761 (N_761,N_689,N_608);
and U762 (N_762,N_689,N_657);
nand U763 (N_763,N_603,N_664);
nor U764 (N_764,N_619,N_613);
and U765 (N_765,N_696,N_661);
nor U766 (N_766,N_646,N_698);
and U767 (N_767,N_692,N_664);
or U768 (N_768,N_622,N_633);
and U769 (N_769,N_615,N_659);
or U770 (N_770,N_654,N_602);
and U771 (N_771,N_687,N_694);
or U772 (N_772,N_648,N_697);
nand U773 (N_773,N_608,N_603);
nor U774 (N_774,N_641,N_685);
xnor U775 (N_775,N_667,N_647);
or U776 (N_776,N_647,N_637);
nand U777 (N_777,N_650,N_639);
nand U778 (N_778,N_662,N_646);
and U779 (N_779,N_621,N_628);
or U780 (N_780,N_697,N_627);
xnor U781 (N_781,N_641,N_686);
nor U782 (N_782,N_630,N_607);
and U783 (N_783,N_691,N_681);
nor U784 (N_784,N_699,N_691);
and U785 (N_785,N_669,N_642);
xor U786 (N_786,N_680,N_642);
and U787 (N_787,N_675,N_632);
nand U788 (N_788,N_668,N_600);
or U789 (N_789,N_641,N_665);
xnor U790 (N_790,N_621,N_676);
nor U791 (N_791,N_653,N_672);
and U792 (N_792,N_653,N_604);
and U793 (N_793,N_608,N_622);
nor U794 (N_794,N_620,N_639);
nor U795 (N_795,N_602,N_674);
or U796 (N_796,N_647,N_692);
nor U797 (N_797,N_668,N_662);
or U798 (N_798,N_645,N_640);
nor U799 (N_799,N_637,N_664);
or U800 (N_800,N_701,N_717);
and U801 (N_801,N_779,N_703);
nand U802 (N_802,N_712,N_790);
nand U803 (N_803,N_766,N_764);
and U804 (N_804,N_776,N_762);
nand U805 (N_805,N_714,N_722);
nand U806 (N_806,N_739,N_700);
nor U807 (N_807,N_768,N_741);
nand U808 (N_808,N_752,N_763);
nor U809 (N_809,N_743,N_785);
xnor U810 (N_810,N_760,N_798);
and U811 (N_811,N_729,N_702);
nor U812 (N_812,N_767,N_753);
nand U813 (N_813,N_799,N_783);
nand U814 (N_814,N_796,N_725);
xor U815 (N_815,N_737,N_784);
nand U816 (N_816,N_708,N_727);
nand U817 (N_817,N_733,N_755);
nand U818 (N_818,N_706,N_793);
nand U819 (N_819,N_787,N_786);
nor U820 (N_820,N_746,N_724);
or U821 (N_821,N_740,N_719);
xor U822 (N_822,N_769,N_720);
xor U823 (N_823,N_718,N_774);
or U824 (N_824,N_736,N_704);
and U825 (N_825,N_738,N_742);
and U826 (N_826,N_748,N_756);
nand U827 (N_827,N_773,N_709);
xnor U828 (N_828,N_795,N_735);
and U829 (N_829,N_734,N_751);
and U830 (N_830,N_758,N_771);
and U831 (N_831,N_726,N_745);
or U832 (N_832,N_797,N_723);
or U833 (N_833,N_705,N_791);
or U834 (N_834,N_759,N_707);
and U835 (N_835,N_761,N_780);
or U836 (N_836,N_713,N_754);
or U837 (N_837,N_731,N_775);
nand U838 (N_838,N_747,N_789);
nand U839 (N_839,N_772,N_728);
xor U840 (N_840,N_777,N_792);
and U841 (N_841,N_794,N_778);
and U842 (N_842,N_715,N_750);
or U843 (N_843,N_749,N_781);
xor U844 (N_844,N_711,N_765);
or U845 (N_845,N_716,N_757);
and U846 (N_846,N_730,N_744);
or U847 (N_847,N_721,N_770);
nor U848 (N_848,N_782,N_732);
xnor U849 (N_849,N_710,N_788);
and U850 (N_850,N_789,N_728);
and U851 (N_851,N_762,N_755);
and U852 (N_852,N_753,N_713);
nor U853 (N_853,N_713,N_780);
or U854 (N_854,N_760,N_774);
xor U855 (N_855,N_793,N_781);
xor U856 (N_856,N_792,N_755);
nor U857 (N_857,N_747,N_753);
and U858 (N_858,N_761,N_728);
or U859 (N_859,N_747,N_742);
or U860 (N_860,N_774,N_706);
xor U861 (N_861,N_717,N_760);
xnor U862 (N_862,N_776,N_741);
nand U863 (N_863,N_792,N_770);
and U864 (N_864,N_718,N_762);
and U865 (N_865,N_787,N_749);
or U866 (N_866,N_741,N_769);
nor U867 (N_867,N_792,N_723);
nor U868 (N_868,N_790,N_701);
and U869 (N_869,N_772,N_788);
xor U870 (N_870,N_737,N_741);
or U871 (N_871,N_773,N_725);
or U872 (N_872,N_731,N_716);
nor U873 (N_873,N_761,N_773);
or U874 (N_874,N_716,N_747);
and U875 (N_875,N_707,N_772);
and U876 (N_876,N_793,N_722);
xnor U877 (N_877,N_701,N_785);
or U878 (N_878,N_762,N_721);
xnor U879 (N_879,N_784,N_769);
xor U880 (N_880,N_726,N_743);
nor U881 (N_881,N_780,N_730);
nand U882 (N_882,N_766,N_740);
xor U883 (N_883,N_708,N_700);
nor U884 (N_884,N_747,N_723);
nand U885 (N_885,N_781,N_722);
xor U886 (N_886,N_747,N_718);
nor U887 (N_887,N_711,N_775);
nand U888 (N_888,N_790,N_747);
nor U889 (N_889,N_744,N_718);
or U890 (N_890,N_799,N_701);
and U891 (N_891,N_784,N_782);
or U892 (N_892,N_776,N_742);
or U893 (N_893,N_711,N_708);
xnor U894 (N_894,N_730,N_796);
or U895 (N_895,N_781,N_760);
and U896 (N_896,N_757,N_768);
or U897 (N_897,N_764,N_733);
or U898 (N_898,N_798,N_783);
nor U899 (N_899,N_772,N_765);
and U900 (N_900,N_870,N_830);
nand U901 (N_901,N_885,N_886);
xor U902 (N_902,N_881,N_883);
and U903 (N_903,N_801,N_836);
nor U904 (N_904,N_852,N_818);
nor U905 (N_905,N_897,N_887);
xor U906 (N_906,N_857,N_820);
or U907 (N_907,N_808,N_888);
xnor U908 (N_908,N_876,N_802);
and U909 (N_909,N_891,N_856);
nor U910 (N_910,N_865,N_833);
or U911 (N_911,N_828,N_827);
xor U912 (N_912,N_882,N_859);
or U913 (N_913,N_890,N_855);
xor U914 (N_914,N_806,N_893);
nand U915 (N_915,N_814,N_879);
or U916 (N_916,N_838,N_848);
or U917 (N_917,N_840,N_810);
nor U918 (N_918,N_869,N_804);
nor U919 (N_919,N_845,N_816);
or U920 (N_920,N_894,N_875);
nor U921 (N_921,N_825,N_867);
xor U922 (N_922,N_831,N_826);
or U923 (N_923,N_846,N_844);
or U924 (N_924,N_850,N_862);
xnor U925 (N_925,N_805,N_815);
nor U926 (N_926,N_842,N_800);
and U927 (N_927,N_877,N_878);
nand U928 (N_928,N_872,N_809);
and U929 (N_929,N_898,N_884);
nand U930 (N_930,N_861,N_839);
or U931 (N_931,N_854,N_863);
nor U932 (N_932,N_880,N_813);
and U933 (N_933,N_847,N_860);
nor U934 (N_934,N_821,N_823);
and U935 (N_935,N_832,N_851);
nand U936 (N_936,N_871,N_858);
and U937 (N_937,N_807,N_819);
and U938 (N_938,N_896,N_873);
or U939 (N_939,N_824,N_899);
nand U940 (N_940,N_834,N_835);
xnor U941 (N_941,N_811,N_864);
nor U942 (N_942,N_849,N_853);
nand U943 (N_943,N_868,N_866);
and U944 (N_944,N_822,N_829);
xor U945 (N_945,N_874,N_843);
or U946 (N_946,N_889,N_837);
nand U947 (N_947,N_895,N_841);
nand U948 (N_948,N_803,N_817);
or U949 (N_949,N_892,N_812);
nand U950 (N_950,N_819,N_808);
nor U951 (N_951,N_888,N_882);
nand U952 (N_952,N_864,N_871);
or U953 (N_953,N_811,N_878);
xnor U954 (N_954,N_824,N_858);
xnor U955 (N_955,N_820,N_833);
and U956 (N_956,N_882,N_884);
xnor U957 (N_957,N_832,N_891);
and U958 (N_958,N_802,N_862);
and U959 (N_959,N_848,N_821);
nand U960 (N_960,N_811,N_855);
nor U961 (N_961,N_858,N_893);
nor U962 (N_962,N_861,N_810);
and U963 (N_963,N_856,N_802);
xor U964 (N_964,N_888,N_823);
and U965 (N_965,N_893,N_884);
nor U966 (N_966,N_829,N_823);
and U967 (N_967,N_871,N_803);
xnor U968 (N_968,N_895,N_810);
nand U969 (N_969,N_896,N_831);
nor U970 (N_970,N_824,N_843);
and U971 (N_971,N_829,N_887);
nand U972 (N_972,N_872,N_846);
xor U973 (N_973,N_845,N_852);
or U974 (N_974,N_841,N_890);
xnor U975 (N_975,N_852,N_889);
or U976 (N_976,N_869,N_863);
and U977 (N_977,N_810,N_837);
nand U978 (N_978,N_888,N_871);
nand U979 (N_979,N_868,N_876);
nor U980 (N_980,N_876,N_844);
nor U981 (N_981,N_858,N_856);
nor U982 (N_982,N_880,N_834);
or U983 (N_983,N_876,N_803);
nand U984 (N_984,N_874,N_896);
xnor U985 (N_985,N_856,N_845);
or U986 (N_986,N_867,N_875);
xnor U987 (N_987,N_887,N_846);
nor U988 (N_988,N_874,N_873);
nor U989 (N_989,N_801,N_810);
and U990 (N_990,N_853,N_894);
nand U991 (N_991,N_866,N_848);
and U992 (N_992,N_826,N_834);
nand U993 (N_993,N_858,N_812);
nor U994 (N_994,N_844,N_823);
nor U995 (N_995,N_875,N_898);
or U996 (N_996,N_885,N_835);
xnor U997 (N_997,N_844,N_820);
and U998 (N_998,N_877,N_888);
nor U999 (N_999,N_854,N_831);
or U1000 (N_1000,N_955,N_919);
or U1001 (N_1001,N_970,N_949);
and U1002 (N_1002,N_910,N_929);
and U1003 (N_1003,N_962,N_920);
nand U1004 (N_1004,N_964,N_966);
and U1005 (N_1005,N_913,N_925);
xnor U1006 (N_1006,N_996,N_967);
nor U1007 (N_1007,N_911,N_994);
xor U1008 (N_1008,N_935,N_992);
and U1009 (N_1009,N_976,N_952);
or U1010 (N_1010,N_948,N_978);
or U1011 (N_1011,N_905,N_931);
nand U1012 (N_1012,N_977,N_960);
nor U1013 (N_1013,N_953,N_981);
nor U1014 (N_1014,N_941,N_938);
and U1015 (N_1015,N_969,N_984);
nand U1016 (N_1016,N_915,N_943);
nand U1017 (N_1017,N_958,N_940);
nor U1018 (N_1018,N_983,N_917);
and U1019 (N_1019,N_995,N_937);
xnor U1020 (N_1020,N_980,N_923);
xnor U1021 (N_1021,N_973,N_901);
nor U1022 (N_1022,N_971,N_999);
nor U1023 (N_1023,N_932,N_902);
or U1024 (N_1024,N_975,N_963);
and U1025 (N_1025,N_989,N_974);
nand U1026 (N_1026,N_934,N_908);
or U1027 (N_1027,N_986,N_936);
or U1028 (N_1028,N_924,N_909);
nand U1029 (N_1029,N_954,N_991);
nor U1030 (N_1030,N_945,N_930);
or U1031 (N_1031,N_979,N_903);
nand U1032 (N_1032,N_993,N_972);
or U1033 (N_1033,N_985,N_907);
nor U1034 (N_1034,N_946,N_912);
or U1035 (N_1035,N_957,N_918);
and U1036 (N_1036,N_922,N_968);
and U1037 (N_1037,N_950,N_921);
or U1038 (N_1038,N_988,N_900);
xnor U1039 (N_1039,N_961,N_956);
nand U1040 (N_1040,N_916,N_933);
or U1041 (N_1041,N_927,N_947);
and U1042 (N_1042,N_990,N_959);
and U1043 (N_1043,N_914,N_998);
nor U1044 (N_1044,N_942,N_951);
or U1045 (N_1045,N_904,N_928);
nand U1046 (N_1046,N_939,N_965);
xor U1047 (N_1047,N_944,N_997);
nand U1048 (N_1048,N_906,N_987);
nor U1049 (N_1049,N_982,N_926);
or U1050 (N_1050,N_942,N_972);
xnor U1051 (N_1051,N_995,N_998);
xor U1052 (N_1052,N_937,N_958);
and U1053 (N_1053,N_938,N_930);
nand U1054 (N_1054,N_946,N_966);
nand U1055 (N_1055,N_955,N_949);
and U1056 (N_1056,N_944,N_965);
or U1057 (N_1057,N_910,N_990);
nand U1058 (N_1058,N_963,N_914);
or U1059 (N_1059,N_959,N_993);
xor U1060 (N_1060,N_909,N_921);
nand U1061 (N_1061,N_969,N_917);
xnor U1062 (N_1062,N_901,N_924);
xnor U1063 (N_1063,N_913,N_911);
nand U1064 (N_1064,N_996,N_998);
or U1065 (N_1065,N_930,N_922);
and U1066 (N_1066,N_978,N_994);
or U1067 (N_1067,N_921,N_919);
nand U1068 (N_1068,N_948,N_975);
xnor U1069 (N_1069,N_937,N_916);
and U1070 (N_1070,N_981,N_926);
nor U1071 (N_1071,N_946,N_942);
and U1072 (N_1072,N_952,N_997);
nor U1073 (N_1073,N_980,N_919);
and U1074 (N_1074,N_919,N_927);
or U1075 (N_1075,N_959,N_998);
xnor U1076 (N_1076,N_937,N_941);
and U1077 (N_1077,N_919,N_965);
and U1078 (N_1078,N_920,N_947);
nand U1079 (N_1079,N_964,N_962);
and U1080 (N_1080,N_948,N_928);
and U1081 (N_1081,N_957,N_978);
or U1082 (N_1082,N_954,N_957);
xor U1083 (N_1083,N_993,N_961);
and U1084 (N_1084,N_938,N_923);
xnor U1085 (N_1085,N_970,N_923);
nor U1086 (N_1086,N_941,N_946);
nor U1087 (N_1087,N_959,N_963);
and U1088 (N_1088,N_916,N_980);
and U1089 (N_1089,N_936,N_957);
nor U1090 (N_1090,N_975,N_996);
and U1091 (N_1091,N_928,N_907);
xnor U1092 (N_1092,N_914,N_989);
xor U1093 (N_1093,N_925,N_956);
and U1094 (N_1094,N_956,N_970);
nor U1095 (N_1095,N_996,N_989);
and U1096 (N_1096,N_962,N_985);
nor U1097 (N_1097,N_919,N_901);
and U1098 (N_1098,N_910,N_978);
or U1099 (N_1099,N_976,N_954);
and U1100 (N_1100,N_1089,N_1019);
and U1101 (N_1101,N_1063,N_1056);
and U1102 (N_1102,N_1016,N_1006);
nand U1103 (N_1103,N_1042,N_1061);
nand U1104 (N_1104,N_1008,N_1012);
or U1105 (N_1105,N_1040,N_1034);
or U1106 (N_1106,N_1027,N_1064);
nor U1107 (N_1107,N_1041,N_1009);
and U1108 (N_1108,N_1033,N_1078);
nor U1109 (N_1109,N_1071,N_1075);
or U1110 (N_1110,N_1047,N_1059);
xnor U1111 (N_1111,N_1007,N_1085);
xnor U1112 (N_1112,N_1095,N_1050);
nand U1113 (N_1113,N_1076,N_1044);
xnor U1114 (N_1114,N_1024,N_1010);
or U1115 (N_1115,N_1096,N_1086);
and U1116 (N_1116,N_1066,N_1088);
nand U1117 (N_1117,N_1060,N_1022);
or U1118 (N_1118,N_1030,N_1026);
xnor U1119 (N_1119,N_1048,N_1020);
nor U1120 (N_1120,N_1094,N_1068);
or U1121 (N_1121,N_1082,N_1072);
and U1122 (N_1122,N_1097,N_1004);
nor U1123 (N_1123,N_1028,N_1081);
or U1124 (N_1124,N_1083,N_1053);
xor U1125 (N_1125,N_1052,N_1031);
or U1126 (N_1126,N_1002,N_1015);
or U1127 (N_1127,N_1036,N_1090);
nand U1128 (N_1128,N_1023,N_1039);
and U1129 (N_1129,N_1062,N_1003);
and U1130 (N_1130,N_1067,N_1054);
nand U1131 (N_1131,N_1073,N_1043);
nor U1132 (N_1132,N_1098,N_1057);
or U1133 (N_1133,N_1092,N_1087);
nand U1134 (N_1134,N_1070,N_1049);
xor U1135 (N_1135,N_1005,N_1065);
nand U1136 (N_1136,N_1046,N_1000);
nand U1137 (N_1137,N_1045,N_1084);
and U1138 (N_1138,N_1055,N_1032);
nor U1139 (N_1139,N_1080,N_1018);
xnor U1140 (N_1140,N_1079,N_1029);
nand U1141 (N_1141,N_1069,N_1077);
or U1142 (N_1142,N_1011,N_1093);
nor U1143 (N_1143,N_1091,N_1038);
nand U1144 (N_1144,N_1051,N_1001);
or U1145 (N_1145,N_1037,N_1017);
xnor U1146 (N_1146,N_1021,N_1074);
and U1147 (N_1147,N_1013,N_1014);
xor U1148 (N_1148,N_1099,N_1035);
xor U1149 (N_1149,N_1058,N_1025);
or U1150 (N_1150,N_1032,N_1041);
and U1151 (N_1151,N_1037,N_1030);
xnor U1152 (N_1152,N_1073,N_1049);
xnor U1153 (N_1153,N_1090,N_1094);
nor U1154 (N_1154,N_1020,N_1073);
nand U1155 (N_1155,N_1073,N_1010);
xor U1156 (N_1156,N_1032,N_1024);
and U1157 (N_1157,N_1095,N_1014);
xnor U1158 (N_1158,N_1092,N_1025);
or U1159 (N_1159,N_1026,N_1094);
nor U1160 (N_1160,N_1050,N_1055);
and U1161 (N_1161,N_1047,N_1098);
or U1162 (N_1162,N_1038,N_1007);
or U1163 (N_1163,N_1036,N_1063);
and U1164 (N_1164,N_1043,N_1094);
nand U1165 (N_1165,N_1043,N_1038);
or U1166 (N_1166,N_1029,N_1005);
and U1167 (N_1167,N_1088,N_1014);
or U1168 (N_1168,N_1096,N_1089);
nor U1169 (N_1169,N_1071,N_1099);
nand U1170 (N_1170,N_1038,N_1014);
and U1171 (N_1171,N_1090,N_1047);
nand U1172 (N_1172,N_1074,N_1080);
or U1173 (N_1173,N_1058,N_1007);
xor U1174 (N_1174,N_1058,N_1043);
nand U1175 (N_1175,N_1079,N_1073);
or U1176 (N_1176,N_1088,N_1019);
xnor U1177 (N_1177,N_1042,N_1017);
nand U1178 (N_1178,N_1016,N_1000);
and U1179 (N_1179,N_1064,N_1017);
or U1180 (N_1180,N_1085,N_1070);
nand U1181 (N_1181,N_1013,N_1038);
or U1182 (N_1182,N_1083,N_1030);
and U1183 (N_1183,N_1003,N_1048);
and U1184 (N_1184,N_1001,N_1088);
or U1185 (N_1185,N_1099,N_1059);
or U1186 (N_1186,N_1077,N_1017);
xnor U1187 (N_1187,N_1022,N_1064);
and U1188 (N_1188,N_1060,N_1026);
xnor U1189 (N_1189,N_1098,N_1076);
nor U1190 (N_1190,N_1023,N_1071);
and U1191 (N_1191,N_1066,N_1077);
nor U1192 (N_1192,N_1085,N_1082);
and U1193 (N_1193,N_1092,N_1049);
nor U1194 (N_1194,N_1034,N_1088);
or U1195 (N_1195,N_1098,N_1030);
and U1196 (N_1196,N_1015,N_1094);
or U1197 (N_1197,N_1015,N_1067);
nor U1198 (N_1198,N_1008,N_1030);
and U1199 (N_1199,N_1016,N_1032);
xnor U1200 (N_1200,N_1125,N_1143);
nor U1201 (N_1201,N_1176,N_1131);
xor U1202 (N_1202,N_1186,N_1115);
nand U1203 (N_1203,N_1105,N_1149);
xor U1204 (N_1204,N_1155,N_1193);
nand U1205 (N_1205,N_1194,N_1137);
xor U1206 (N_1206,N_1195,N_1122);
or U1207 (N_1207,N_1140,N_1180);
or U1208 (N_1208,N_1102,N_1162);
xor U1209 (N_1209,N_1185,N_1158);
nand U1210 (N_1210,N_1164,N_1111);
nor U1211 (N_1211,N_1116,N_1178);
and U1212 (N_1212,N_1146,N_1101);
and U1213 (N_1213,N_1129,N_1139);
or U1214 (N_1214,N_1174,N_1165);
or U1215 (N_1215,N_1189,N_1117);
and U1216 (N_1216,N_1190,N_1130);
or U1217 (N_1217,N_1151,N_1133);
and U1218 (N_1218,N_1150,N_1170);
xor U1219 (N_1219,N_1119,N_1153);
or U1220 (N_1220,N_1141,N_1166);
nor U1221 (N_1221,N_1144,N_1175);
nor U1222 (N_1222,N_1161,N_1159);
nor U1223 (N_1223,N_1160,N_1107);
nand U1224 (N_1224,N_1187,N_1181);
and U1225 (N_1225,N_1145,N_1114);
xnor U1226 (N_1226,N_1163,N_1192);
and U1227 (N_1227,N_1173,N_1157);
xnor U1228 (N_1228,N_1152,N_1169);
nand U1229 (N_1229,N_1132,N_1171);
xnor U1230 (N_1230,N_1103,N_1191);
nand U1231 (N_1231,N_1188,N_1127);
or U1232 (N_1232,N_1142,N_1108);
and U1233 (N_1233,N_1128,N_1124);
or U1234 (N_1234,N_1100,N_1182);
nand U1235 (N_1235,N_1134,N_1198);
nand U1236 (N_1236,N_1197,N_1136);
and U1237 (N_1237,N_1112,N_1147);
and U1238 (N_1238,N_1167,N_1148);
xor U1239 (N_1239,N_1113,N_1123);
xnor U1240 (N_1240,N_1199,N_1179);
and U1241 (N_1241,N_1126,N_1183);
nor U1242 (N_1242,N_1104,N_1120);
xnor U1243 (N_1243,N_1109,N_1184);
and U1244 (N_1244,N_1106,N_1138);
xor U1245 (N_1245,N_1196,N_1121);
nor U1246 (N_1246,N_1110,N_1177);
and U1247 (N_1247,N_1154,N_1118);
xor U1248 (N_1248,N_1156,N_1135);
nand U1249 (N_1249,N_1168,N_1172);
or U1250 (N_1250,N_1134,N_1185);
nand U1251 (N_1251,N_1158,N_1153);
nor U1252 (N_1252,N_1160,N_1152);
nand U1253 (N_1253,N_1171,N_1106);
xor U1254 (N_1254,N_1161,N_1102);
xor U1255 (N_1255,N_1145,N_1103);
nand U1256 (N_1256,N_1190,N_1177);
or U1257 (N_1257,N_1116,N_1177);
or U1258 (N_1258,N_1109,N_1120);
xnor U1259 (N_1259,N_1198,N_1152);
nand U1260 (N_1260,N_1133,N_1103);
xor U1261 (N_1261,N_1112,N_1104);
nor U1262 (N_1262,N_1143,N_1135);
and U1263 (N_1263,N_1117,N_1120);
and U1264 (N_1264,N_1153,N_1136);
nor U1265 (N_1265,N_1193,N_1139);
xnor U1266 (N_1266,N_1147,N_1196);
xnor U1267 (N_1267,N_1197,N_1138);
xnor U1268 (N_1268,N_1148,N_1144);
and U1269 (N_1269,N_1191,N_1189);
and U1270 (N_1270,N_1113,N_1171);
or U1271 (N_1271,N_1159,N_1169);
nor U1272 (N_1272,N_1186,N_1175);
xnor U1273 (N_1273,N_1106,N_1137);
nand U1274 (N_1274,N_1117,N_1141);
nand U1275 (N_1275,N_1151,N_1116);
and U1276 (N_1276,N_1182,N_1102);
xnor U1277 (N_1277,N_1136,N_1129);
or U1278 (N_1278,N_1178,N_1144);
or U1279 (N_1279,N_1141,N_1154);
nor U1280 (N_1280,N_1197,N_1153);
and U1281 (N_1281,N_1188,N_1100);
xor U1282 (N_1282,N_1106,N_1100);
and U1283 (N_1283,N_1100,N_1137);
or U1284 (N_1284,N_1199,N_1145);
and U1285 (N_1285,N_1118,N_1136);
nand U1286 (N_1286,N_1105,N_1181);
xor U1287 (N_1287,N_1100,N_1117);
nand U1288 (N_1288,N_1138,N_1119);
and U1289 (N_1289,N_1145,N_1152);
and U1290 (N_1290,N_1132,N_1130);
or U1291 (N_1291,N_1192,N_1165);
nand U1292 (N_1292,N_1189,N_1159);
or U1293 (N_1293,N_1162,N_1161);
nor U1294 (N_1294,N_1136,N_1182);
nand U1295 (N_1295,N_1114,N_1158);
nand U1296 (N_1296,N_1193,N_1179);
and U1297 (N_1297,N_1107,N_1114);
and U1298 (N_1298,N_1179,N_1105);
nor U1299 (N_1299,N_1155,N_1195);
and U1300 (N_1300,N_1290,N_1287);
and U1301 (N_1301,N_1244,N_1200);
or U1302 (N_1302,N_1204,N_1237);
nor U1303 (N_1303,N_1206,N_1221);
nor U1304 (N_1304,N_1214,N_1292);
or U1305 (N_1305,N_1230,N_1263);
nand U1306 (N_1306,N_1286,N_1291);
and U1307 (N_1307,N_1278,N_1267);
or U1308 (N_1308,N_1220,N_1295);
nand U1309 (N_1309,N_1213,N_1215);
and U1310 (N_1310,N_1251,N_1289);
nand U1311 (N_1311,N_1233,N_1275);
nor U1312 (N_1312,N_1285,N_1280);
nor U1313 (N_1313,N_1223,N_1205);
nand U1314 (N_1314,N_1265,N_1246);
nor U1315 (N_1315,N_1227,N_1226);
and U1316 (N_1316,N_1229,N_1299);
nand U1317 (N_1317,N_1212,N_1261);
nor U1318 (N_1318,N_1264,N_1234);
and U1319 (N_1319,N_1279,N_1236);
and U1320 (N_1320,N_1296,N_1259);
or U1321 (N_1321,N_1211,N_1274);
nand U1322 (N_1322,N_1268,N_1218);
or U1323 (N_1323,N_1248,N_1271);
and U1324 (N_1324,N_1238,N_1231);
nor U1325 (N_1325,N_1266,N_1262);
and U1326 (N_1326,N_1209,N_1272);
and U1327 (N_1327,N_1258,N_1216);
nand U1328 (N_1328,N_1201,N_1288);
nor U1329 (N_1329,N_1240,N_1239);
nand U1330 (N_1330,N_1222,N_1210);
nand U1331 (N_1331,N_1242,N_1297);
or U1332 (N_1332,N_1250,N_1273);
or U1333 (N_1333,N_1228,N_1235);
or U1334 (N_1334,N_1253,N_1241);
or U1335 (N_1335,N_1294,N_1219);
and U1336 (N_1336,N_1208,N_1202);
and U1337 (N_1337,N_1203,N_1260);
nand U1338 (N_1338,N_1293,N_1256);
nor U1339 (N_1339,N_1284,N_1298);
or U1340 (N_1340,N_1252,N_1254);
and U1341 (N_1341,N_1217,N_1225);
and U1342 (N_1342,N_1281,N_1224);
xnor U1343 (N_1343,N_1245,N_1270);
or U1344 (N_1344,N_1269,N_1232);
and U1345 (N_1345,N_1282,N_1249);
xnor U1346 (N_1346,N_1255,N_1257);
xor U1347 (N_1347,N_1283,N_1247);
nand U1348 (N_1348,N_1207,N_1276);
or U1349 (N_1349,N_1277,N_1243);
xnor U1350 (N_1350,N_1296,N_1243);
or U1351 (N_1351,N_1213,N_1280);
xor U1352 (N_1352,N_1221,N_1255);
nand U1353 (N_1353,N_1229,N_1241);
nor U1354 (N_1354,N_1296,N_1260);
nand U1355 (N_1355,N_1226,N_1243);
xnor U1356 (N_1356,N_1248,N_1215);
xor U1357 (N_1357,N_1296,N_1245);
and U1358 (N_1358,N_1239,N_1266);
nor U1359 (N_1359,N_1240,N_1261);
nand U1360 (N_1360,N_1206,N_1288);
or U1361 (N_1361,N_1270,N_1201);
and U1362 (N_1362,N_1278,N_1247);
nand U1363 (N_1363,N_1280,N_1239);
xnor U1364 (N_1364,N_1212,N_1272);
xnor U1365 (N_1365,N_1263,N_1280);
and U1366 (N_1366,N_1279,N_1298);
xor U1367 (N_1367,N_1208,N_1255);
and U1368 (N_1368,N_1263,N_1218);
and U1369 (N_1369,N_1211,N_1255);
and U1370 (N_1370,N_1297,N_1279);
xnor U1371 (N_1371,N_1265,N_1260);
nor U1372 (N_1372,N_1281,N_1207);
and U1373 (N_1373,N_1236,N_1237);
nor U1374 (N_1374,N_1220,N_1218);
or U1375 (N_1375,N_1273,N_1221);
and U1376 (N_1376,N_1223,N_1256);
or U1377 (N_1377,N_1242,N_1276);
nor U1378 (N_1378,N_1233,N_1209);
nor U1379 (N_1379,N_1233,N_1263);
or U1380 (N_1380,N_1227,N_1208);
nor U1381 (N_1381,N_1276,N_1269);
nor U1382 (N_1382,N_1242,N_1236);
and U1383 (N_1383,N_1255,N_1207);
nand U1384 (N_1384,N_1273,N_1256);
or U1385 (N_1385,N_1253,N_1270);
xnor U1386 (N_1386,N_1281,N_1204);
nor U1387 (N_1387,N_1208,N_1240);
xnor U1388 (N_1388,N_1266,N_1268);
xnor U1389 (N_1389,N_1240,N_1216);
xor U1390 (N_1390,N_1263,N_1294);
nand U1391 (N_1391,N_1247,N_1205);
or U1392 (N_1392,N_1272,N_1222);
nor U1393 (N_1393,N_1206,N_1210);
nor U1394 (N_1394,N_1214,N_1202);
or U1395 (N_1395,N_1204,N_1272);
nor U1396 (N_1396,N_1212,N_1276);
nand U1397 (N_1397,N_1259,N_1284);
and U1398 (N_1398,N_1279,N_1268);
nand U1399 (N_1399,N_1205,N_1245);
and U1400 (N_1400,N_1347,N_1353);
xor U1401 (N_1401,N_1319,N_1343);
and U1402 (N_1402,N_1389,N_1307);
nor U1403 (N_1403,N_1301,N_1312);
nor U1404 (N_1404,N_1327,N_1332);
and U1405 (N_1405,N_1352,N_1398);
nand U1406 (N_1406,N_1363,N_1323);
and U1407 (N_1407,N_1378,N_1390);
xor U1408 (N_1408,N_1383,N_1348);
nand U1409 (N_1409,N_1364,N_1349);
and U1410 (N_1410,N_1354,N_1385);
nor U1411 (N_1411,N_1310,N_1372);
or U1412 (N_1412,N_1380,N_1377);
xor U1413 (N_1413,N_1341,N_1340);
nand U1414 (N_1414,N_1395,N_1386);
xnor U1415 (N_1415,N_1333,N_1382);
nand U1416 (N_1416,N_1397,N_1350);
xnor U1417 (N_1417,N_1396,N_1342);
nand U1418 (N_1418,N_1315,N_1322);
and U1419 (N_1419,N_1374,N_1376);
nand U1420 (N_1420,N_1337,N_1367);
and U1421 (N_1421,N_1373,N_1392);
or U1422 (N_1422,N_1338,N_1318);
nor U1423 (N_1423,N_1399,N_1339);
nor U1424 (N_1424,N_1314,N_1303);
and U1425 (N_1425,N_1300,N_1311);
nor U1426 (N_1426,N_1324,N_1351);
xnor U1427 (N_1427,N_1391,N_1346);
nand U1428 (N_1428,N_1358,N_1330);
and U1429 (N_1429,N_1345,N_1362);
xor U1430 (N_1430,N_1335,N_1375);
or U1431 (N_1431,N_1344,N_1331);
nand U1432 (N_1432,N_1302,N_1365);
nor U1433 (N_1433,N_1394,N_1313);
nand U1434 (N_1434,N_1305,N_1321);
or U1435 (N_1435,N_1326,N_1309);
nand U1436 (N_1436,N_1379,N_1384);
xnor U1437 (N_1437,N_1369,N_1336);
or U1438 (N_1438,N_1355,N_1306);
nor U1439 (N_1439,N_1388,N_1359);
nand U1440 (N_1440,N_1317,N_1308);
nand U1441 (N_1441,N_1366,N_1316);
or U1442 (N_1442,N_1357,N_1370);
nor U1443 (N_1443,N_1368,N_1381);
nand U1444 (N_1444,N_1325,N_1304);
nand U1445 (N_1445,N_1356,N_1334);
and U1446 (N_1446,N_1360,N_1387);
and U1447 (N_1447,N_1329,N_1320);
or U1448 (N_1448,N_1393,N_1361);
or U1449 (N_1449,N_1328,N_1371);
nor U1450 (N_1450,N_1351,N_1388);
or U1451 (N_1451,N_1304,N_1307);
nor U1452 (N_1452,N_1315,N_1364);
or U1453 (N_1453,N_1373,N_1345);
xor U1454 (N_1454,N_1387,N_1319);
xor U1455 (N_1455,N_1323,N_1370);
xor U1456 (N_1456,N_1332,N_1314);
nand U1457 (N_1457,N_1361,N_1373);
and U1458 (N_1458,N_1367,N_1361);
nand U1459 (N_1459,N_1309,N_1347);
nor U1460 (N_1460,N_1330,N_1362);
nand U1461 (N_1461,N_1342,N_1352);
and U1462 (N_1462,N_1367,N_1336);
nand U1463 (N_1463,N_1371,N_1305);
nor U1464 (N_1464,N_1333,N_1370);
and U1465 (N_1465,N_1337,N_1355);
nand U1466 (N_1466,N_1385,N_1300);
nand U1467 (N_1467,N_1316,N_1375);
or U1468 (N_1468,N_1350,N_1324);
and U1469 (N_1469,N_1333,N_1371);
xnor U1470 (N_1470,N_1389,N_1371);
or U1471 (N_1471,N_1398,N_1307);
nor U1472 (N_1472,N_1344,N_1395);
nor U1473 (N_1473,N_1361,N_1300);
nor U1474 (N_1474,N_1322,N_1320);
and U1475 (N_1475,N_1346,N_1366);
or U1476 (N_1476,N_1363,N_1330);
nand U1477 (N_1477,N_1397,N_1316);
or U1478 (N_1478,N_1331,N_1396);
xnor U1479 (N_1479,N_1335,N_1304);
nand U1480 (N_1480,N_1365,N_1394);
or U1481 (N_1481,N_1384,N_1360);
nor U1482 (N_1482,N_1372,N_1392);
nand U1483 (N_1483,N_1323,N_1336);
or U1484 (N_1484,N_1350,N_1318);
xnor U1485 (N_1485,N_1314,N_1399);
xor U1486 (N_1486,N_1375,N_1348);
nand U1487 (N_1487,N_1325,N_1347);
and U1488 (N_1488,N_1324,N_1355);
xnor U1489 (N_1489,N_1358,N_1367);
xnor U1490 (N_1490,N_1340,N_1365);
xnor U1491 (N_1491,N_1307,N_1363);
xor U1492 (N_1492,N_1349,N_1336);
and U1493 (N_1493,N_1362,N_1318);
nand U1494 (N_1494,N_1346,N_1350);
nor U1495 (N_1495,N_1349,N_1334);
nand U1496 (N_1496,N_1399,N_1335);
xor U1497 (N_1497,N_1381,N_1318);
xnor U1498 (N_1498,N_1374,N_1377);
or U1499 (N_1499,N_1382,N_1367);
xor U1500 (N_1500,N_1462,N_1436);
nor U1501 (N_1501,N_1405,N_1433);
nand U1502 (N_1502,N_1411,N_1488);
and U1503 (N_1503,N_1406,N_1443);
xor U1504 (N_1504,N_1426,N_1463);
and U1505 (N_1505,N_1495,N_1490);
xnor U1506 (N_1506,N_1413,N_1438);
xnor U1507 (N_1507,N_1494,N_1469);
xor U1508 (N_1508,N_1479,N_1447);
or U1509 (N_1509,N_1415,N_1460);
or U1510 (N_1510,N_1465,N_1441);
and U1511 (N_1511,N_1427,N_1440);
and U1512 (N_1512,N_1412,N_1409);
nand U1513 (N_1513,N_1454,N_1464);
nand U1514 (N_1514,N_1492,N_1439);
and U1515 (N_1515,N_1467,N_1482);
xor U1516 (N_1516,N_1444,N_1486);
and U1517 (N_1517,N_1446,N_1472);
nor U1518 (N_1518,N_1407,N_1425);
and U1519 (N_1519,N_1496,N_1419);
nor U1520 (N_1520,N_1484,N_1455);
and U1521 (N_1521,N_1442,N_1481);
and U1522 (N_1522,N_1420,N_1487);
nand U1523 (N_1523,N_1498,N_1448);
and U1524 (N_1524,N_1416,N_1408);
nor U1525 (N_1525,N_1402,N_1445);
xnor U1526 (N_1526,N_1424,N_1431);
or U1527 (N_1527,N_1453,N_1475);
nor U1528 (N_1528,N_1421,N_1429);
nor U1529 (N_1529,N_1423,N_1458);
nor U1530 (N_1530,N_1477,N_1456);
and U1531 (N_1531,N_1478,N_1434);
or U1532 (N_1532,N_1450,N_1468);
nand U1533 (N_1533,N_1404,N_1474);
nor U1534 (N_1534,N_1432,N_1491);
xnor U1535 (N_1535,N_1461,N_1485);
nand U1536 (N_1536,N_1401,N_1493);
nor U1537 (N_1537,N_1403,N_1422);
nor U1538 (N_1538,N_1489,N_1497);
or U1539 (N_1539,N_1449,N_1466);
xor U1540 (N_1540,N_1410,N_1480);
nand U1541 (N_1541,N_1417,N_1418);
nor U1542 (N_1542,N_1435,N_1430);
nand U1543 (N_1543,N_1459,N_1471);
xor U1544 (N_1544,N_1476,N_1437);
and U1545 (N_1545,N_1428,N_1400);
or U1546 (N_1546,N_1483,N_1470);
nand U1547 (N_1547,N_1499,N_1457);
nor U1548 (N_1548,N_1451,N_1473);
or U1549 (N_1549,N_1452,N_1414);
nor U1550 (N_1550,N_1401,N_1427);
nor U1551 (N_1551,N_1498,N_1455);
xnor U1552 (N_1552,N_1401,N_1466);
and U1553 (N_1553,N_1448,N_1473);
xnor U1554 (N_1554,N_1456,N_1470);
nand U1555 (N_1555,N_1416,N_1425);
nand U1556 (N_1556,N_1453,N_1425);
or U1557 (N_1557,N_1419,N_1423);
nand U1558 (N_1558,N_1483,N_1463);
and U1559 (N_1559,N_1490,N_1474);
nor U1560 (N_1560,N_1461,N_1446);
nand U1561 (N_1561,N_1483,N_1446);
xor U1562 (N_1562,N_1444,N_1448);
and U1563 (N_1563,N_1478,N_1444);
xnor U1564 (N_1564,N_1459,N_1473);
and U1565 (N_1565,N_1480,N_1452);
xnor U1566 (N_1566,N_1485,N_1463);
and U1567 (N_1567,N_1472,N_1451);
nand U1568 (N_1568,N_1486,N_1464);
or U1569 (N_1569,N_1430,N_1485);
xnor U1570 (N_1570,N_1405,N_1465);
nor U1571 (N_1571,N_1421,N_1455);
nor U1572 (N_1572,N_1487,N_1431);
xor U1573 (N_1573,N_1463,N_1442);
and U1574 (N_1574,N_1444,N_1443);
and U1575 (N_1575,N_1424,N_1484);
nor U1576 (N_1576,N_1414,N_1400);
nor U1577 (N_1577,N_1400,N_1445);
or U1578 (N_1578,N_1438,N_1477);
or U1579 (N_1579,N_1419,N_1420);
nand U1580 (N_1580,N_1435,N_1461);
nand U1581 (N_1581,N_1490,N_1471);
nor U1582 (N_1582,N_1450,N_1480);
or U1583 (N_1583,N_1402,N_1418);
nor U1584 (N_1584,N_1429,N_1420);
nor U1585 (N_1585,N_1494,N_1415);
and U1586 (N_1586,N_1408,N_1468);
and U1587 (N_1587,N_1464,N_1440);
xnor U1588 (N_1588,N_1401,N_1408);
and U1589 (N_1589,N_1406,N_1430);
xnor U1590 (N_1590,N_1417,N_1430);
and U1591 (N_1591,N_1401,N_1467);
nor U1592 (N_1592,N_1402,N_1498);
or U1593 (N_1593,N_1486,N_1499);
xnor U1594 (N_1594,N_1412,N_1492);
nor U1595 (N_1595,N_1405,N_1455);
nor U1596 (N_1596,N_1461,N_1488);
or U1597 (N_1597,N_1452,N_1497);
nand U1598 (N_1598,N_1486,N_1434);
and U1599 (N_1599,N_1411,N_1486);
nand U1600 (N_1600,N_1539,N_1576);
or U1601 (N_1601,N_1568,N_1528);
nand U1602 (N_1602,N_1518,N_1561);
nor U1603 (N_1603,N_1574,N_1517);
nand U1604 (N_1604,N_1536,N_1534);
nand U1605 (N_1605,N_1549,N_1542);
and U1606 (N_1606,N_1594,N_1502);
and U1607 (N_1607,N_1564,N_1590);
and U1608 (N_1608,N_1543,N_1507);
and U1609 (N_1609,N_1533,N_1538);
and U1610 (N_1610,N_1521,N_1537);
xor U1611 (N_1611,N_1541,N_1560);
and U1612 (N_1612,N_1530,N_1524);
xor U1613 (N_1613,N_1555,N_1596);
xnor U1614 (N_1614,N_1579,N_1529);
nand U1615 (N_1615,N_1575,N_1565);
xnor U1616 (N_1616,N_1501,N_1514);
and U1617 (N_1617,N_1532,N_1588);
and U1618 (N_1618,N_1527,N_1525);
or U1619 (N_1619,N_1587,N_1552);
nor U1620 (N_1620,N_1523,N_1597);
or U1621 (N_1621,N_1520,N_1513);
or U1622 (N_1622,N_1506,N_1510);
and U1623 (N_1623,N_1591,N_1504);
xnor U1624 (N_1624,N_1546,N_1540);
xnor U1625 (N_1625,N_1547,N_1585);
and U1626 (N_1626,N_1572,N_1598);
xnor U1627 (N_1627,N_1551,N_1526);
or U1628 (N_1628,N_1595,N_1582);
or U1629 (N_1629,N_1592,N_1566);
and U1630 (N_1630,N_1578,N_1558);
nor U1631 (N_1631,N_1569,N_1505);
and U1632 (N_1632,N_1544,N_1556);
or U1633 (N_1633,N_1545,N_1509);
nor U1634 (N_1634,N_1531,N_1570);
xnor U1635 (N_1635,N_1573,N_1571);
xnor U1636 (N_1636,N_1508,N_1511);
nand U1637 (N_1637,N_1515,N_1554);
nor U1638 (N_1638,N_1593,N_1586);
or U1639 (N_1639,N_1500,N_1580);
xor U1640 (N_1640,N_1535,N_1562);
xor U1641 (N_1641,N_1519,N_1599);
xor U1642 (N_1642,N_1516,N_1557);
nand U1643 (N_1643,N_1512,N_1567);
nor U1644 (N_1644,N_1584,N_1548);
and U1645 (N_1645,N_1583,N_1522);
nand U1646 (N_1646,N_1577,N_1589);
or U1647 (N_1647,N_1559,N_1563);
nor U1648 (N_1648,N_1503,N_1553);
xnor U1649 (N_1649,N_1550,N_1581);
nor U1650 (N_1650,N_1500,N_1595);
xor U1651 (N_1651,N_1540,N_1579);
nor U1652 (N_1652,N_1509,N_1585);
or U1653 (N_1653,N_1580,N_1584);
nand U1654 (N_1654,N_1514,N_1594);
xnor U1655 (N_1655,N_1503,N_1534);
or U1656 (N_1656,N_1570,N_1577);
xnor U1657 (N_1657,N_1541,N_1514);
nand U1658 (N_1658,N_1517,N_1508);
and U1659 (N_1659,N_1533,N_1554);
nand U1660 (N_1660,N_1532,N_1597);
xnor U1661 (N_1661,N_1534,N_1541);
xor U1662 (N_1662,N_1520,N_1575);
nand U1663 (N_1663,N_1587,N_1577);
or U1664 (N_1664,N_1544,N_1550);
and U1665 (N_1665,N_1558,N_1555);
and U1666 (N_1666,N_1578,N_1555);
and U1667 (N_1667,N_1539,N_1598);
and U1668 (N_1668,N_1542,N_1548);
xor U1669 (N_1669,N_1560,N_1595);
nor U1670 (N_1670,N_1519,N_1509);
and U1671 (N_1671,N_1543,N_1506);
or U1672 (N_1672,N_1549,N_1560);
and U1673 (N_1673,N_1569,N_1564);
or U1674 (N_1674,N_1512,N_1540);
nand U1675 (N_1675,N_1589,N_1527);
nand U1676 (N_1676,N_1526,N_1516);
nor U1677 (N_1677,N_1525,N_1564);
and U1678 (N_1678,N_1556,N_1590);
and U1679 (N_1679,N_1558,N_1545);
or U1680 (N_1680,N_1529,N_1591);
and U1681 (N_1681,N_1560,N_1548);
xnor U1682 (N_1682,N_1547,N_1590);
and U1683 (N_1683,N_1587,N_1506);
or U1684 (N_1684,N_1531,N_1521);
nor U1685 (N_1685,N_1520,N_1596);
or U1686 (N_1686,N_1505,N_1520);
or U1687 (N_1687,N_1556,N_1574);
nand U1688 (N_1688,N_1541,N_1543);
and U1689 (N_1689,N_1544,N_1512);
nor U1690 (N_1690,N_1593,N_1504);
xor U1691 (N_1691,N_1580,N_1520);
and U1692 (N_1692,N_1589,N_1506);
xor U1693 (N_1693,N_1513,N_1511);
xnor U1694 (N_1694,N_1555,N_1510);
or U1695 (N_1695,N_1589,N_1501);
xor U1696 (N_1696,N_1525,N_1587);
and U1697 (N_1697,N_1500,N_1530);
and U1698 (N_1698,N_1501,N_1594);
nor U1699 (N_1699,N_1512,N_1536);
nand U1700 (N_1700,N_1623,N_1686);
or U1701 (N_1701,N_1695,N_1611);
and U1702 (N_1702,N_1618,N_1658);
nor U1703 (N_1703,N_1619,N_1661);
nand U1704 (N_1704,N_1601,N_1634);
xnor U1705 (N_1705,N_1622,N_1698);
nor U1706 (N_1706,N_1650,N_1620);
nand U1707 (N_1707,N_1668,N_1617);
nor U1708 (N_1708,N_1688,N_1645);
or U1709 (N_1709,N_1649,N_1672);
and U1710 (N_1710,N_1642,N_1607);
nand U1711 (N_1711,N_1643,N_1604);
nand U1712 (N_1712,N_1676,N_1696);
nor U1713 (N_1713,N_1651,N_1674);
nand U1714 (N_1714,N_1671,N_1662);
xor U1715 (N_1715,N_1614,N_1659);
nand U1716 (N_1716,N_1663,N_1664);
and U1717 (N_1717,N_1692,N_1630);
and U1718 (N_1718,N_1616,N_1641);
or U1719 (N_1719,N_1699,N_1631);
xor U1720 (N_1720,N_1646,N_1667);
and U1721 (N_1721,N_1687,N_1613);
nor U1722 (N_1722,N_1653,N_1605);
and U1723 (N_1723,N_1689,N_1632);
and U1724 (N_1724,N_1639,N_1656);
or U1725 (N_1725,N_1647,N_1638);
xnor U1726 (N_1726,N_1682,N_1683);
or U1727 (N_1727,N_1629,N_1657);
or U1728 (N_1728,N_1626,N_1625);
nor U1729 (N_1729,N_1606,N_1677);
nand U1730 (N_1730,N_1608,N_1691);
xnor U1731 (N_1731,N_1621,N_1600);
xor U1732 (N_1732,N_1654,N_1648);
and U1733 (N_1733,N_1681,N_1690);
and U1734 (N_1734,N_1678,N_1660);
xnor U1735 (N_1735,N_1652,N_1636);
nor U1736 (N_1736,N_1685,N_1612);
nand U1737 (N_1737,N_1615,N_1628);
or U1738 (N_1738,N_1669,N_1609);
xnor U1739 (N_1739,N_1694,N_1684);
or U1740 (N_1740,N_1644,N_1602);
nor U1741 (N_1741,N_1675,N_1697);
and U1742 (N_1742,N_1666,N_1670);
and U1743 (N_1743,N_1680,N_1627);
xor U1744 (N_1744,N_1693,N_1640);
nand U1745 (N_1745,N_1637,N_1610);
and U1746 (N_1746,N_1603,N_1679);
nor U1747 (N_1747,N_1624,N_1665);
nor U1748 (N_1748,N_1673,N_1635);
nor U1749 (N_1749,N_1633,N_1655);
or U1750 (N_1750,N_1646,N_1641);
or U1751 (N_1751,N_1696,N_1687);
or U1752 (N_1752,N_1685,N_1652);
nor U1753 (N_1753,N_1658,N_1611);
xnor U1754 (N_1754,N_1608,N_1658);
and U1755 (N_1755,N_1617,N_1621);
nand U1756 (N_1756,N_1689,N_1640);
and U1757 (N_1757,N_1676,N_1697);
and U1758 (N_1758,N_1695,N_1612);
nand U1759 (N_1759,N_1618,N_1687);
or U1760 (N_1760,N_1690,N_1636);
and U1761 (N_1761,N_1693,N_1657);
and U1762 (N_1762,N_1603,N_1645);
nand U1763 (N_1763,N_1652,N_1637);
nor U1764 (N_1764,N_1664,N_1699);
and U1765 (N_1765,N_1637,N_1648);
or U1766 (N_1766,N_1627,N_1653);
and U1767 (N_1767,N_1640,N_1623);
nor U1768 (N_1768,N_1641,N_1650);
xor U1769 (N_1769,N_1630,N_1681);
xnor U1770 (N_1770,N_1676,N_1698);
xnor U1771 (N_1771,N_1659,N_1693);
and U1772 (N_1772,N_1627,N_1681);
nor U1773 (N_1773,N_1650,N_1637);
or U1774 (N_1774,N_1668,N_1643);
xnor U1775 (N_1775,N_1636,N_1614);
xnor U1776 (N_1776,N_1633,N_1669);
or U1777 (N_1777,N_1620,N_1639);
or U1778 (N_1778,N_1666,N_1629);
nand U1779 (N_1779,N_1663,N_1611);
or U1780 (N_1780,N_1641,N_1664);
or U1781 (N_1781,N_1620,N_1631);
nor U1782 (N_1782,N_1679,N_1610);
or U1783 (N_1783,N_1660,N_1683);
nand U1784 (N_1784,N_1651,N_1645);
nor U1785 (N_1785,N_1685,N_1609);
xnor U1786 (N_1786,N_1692,N_1667);
or U1787 (N_1787,N_1657,N_1601);
nor U1788 (N_1788,N_1604,N_1686);
nor U1789 (N_1789,N_1678,N_1601);
nand U1790 (N_1790,N_1602,N_1607);
nand U1791 (N_1791,N_1644,N_1697);
or U1792 (N_1792,N_1679,N_1650);
or U1793 (N_1793,N_1662,N_1605);
nand U1794 (N_1794,N_1601,N_1682);
nor U1795 (N_1795,N_1671,N_1687);
nand U1796 (N_1796,N_1635,N_1609);
nand U1797 (N_1797,N_1613,N_1653);
xor U1798 (N_1798,N_1616,N_1661);
nand U1799 (N_1799,N_1680,N_1661);
nor U1800 (N_1800,N_1742,N_1791);
nor U1801 (N_1801,N_1726,N_1749);
or U1802 (N_1802,N_1799,N_1715);
or U1803 (N_1803,N_1720,N_1712);
nor U1804 (N_1804,N_1782,N_1705);
xnor U1805 (N_1805,N_1728,N_1797);
and U1806 (N_1806,N_1719,N_1716);
nor U1807 (N_1807,N_1713,N_1729);
xnor U1808 (N_1808,N_1745,N_1784);
nand U1809 (N_1809,N_1770,N_1798);
nor U1810 (N_1810,N_1732,N_1754);
and U1811 (N_1811,N_1706,N_1766);
and U1812 (N_1812,N_1738,N_1747);
nor U1813 (N_1813,N_1760,N_1762);
nor U1814 (N_1814,N_1739,N_1736);
and U1815 (N_1815,N_1750,N_1777);
xor U1816 (N_1816,N_1727,N_1744);
or U1817 (N_1817,N_1748,N_1700);
and U1818 (N_1818,N_1708,N_1788);
or U1819 (N_1819,N_1787,N_1772);
nor U1820 (N_1820,N_1761,N_1752);
and U1821 (N_1821,N_1711,N_1737);
and U1822 (N_1822,N_1725,N_1753);
nor U1823 (N_1823,N_1786,N_1769);
nand U1824 (N_1824,N_1743,N_1783);
and U1825 (N_1825,N_1794,N_1763);
or U1826 (N_1826,N_1768,N_1703);
nor U1827 (N_1827,N_1741,N_1723);
and U1828 (N_1828,N_1785,N_1709);
xor U1829 (N_1829,N_1775,N_1731);
and U1830 (N_1830,N_1710,N_1778);
xor U1831 (N_1831,N_1780,N_1702);
and U1832 (N_1832,N_1773,N_1756);
or U1833 (N_1833,N_1759,N_1740);
and U1834 (N_1834,N_1774,N_1722);
nor U1835 (N_1835,N_1792,N_1735);
and U1836 (N_1836,N_1796,N_1776);
nand U1837 (N_1837,N_1765,N_1790);
and U1838 (N_1838,N_1755,N_1734);
or U1839 (N_1839,N_1717,N_1771);
nand U1840 (N_1840,N_1789,N_1746);
and U1841 (N_1841,N_1751,N_1767);
nor U1842 (N_1842,N_1707,N_1779);
and U1843 (N_1843,N_1781,N_1724);
nand U1844 (N_1844,N_1758,N_1795);
and U1845 (N_1845,N_1701,N_1733);
xnor U1846 (N_1846,N_1730,N_1704);
nand U1847 (N_1847,N_1714,N_1793);
nand U1848 (N_1848,N_1757,N_1721);
and U1849 (N_1849,N_1764,N_1718);
and U1850 (N_1850,N_1777,N_1758);
xnor U1851 (N_1851,N_1710,N_1715);
or U1852 (N_1852,N_1735,N_1745);
xor U1853 (N_1853,N_1735,N_1701);
nand U1854 (N_1854,N_1786,N_1753);
xnor U1855 (N_1855,N_1766,N_1765);
nand U1856 (N_1856,N_1776,N_1778);
xnor U1857 (N_1857,N_1701,N_1795);
or U1858 (N_1858,N_1780,N_1782);
xnor U1859 (N_1859,N_1728,N_1736);
xnor U1860 (N_1860,N_1702,N_1733);
nor U1861 (N_1861,N_1720,N_1732);
or U1862 (N_1862,N_1780,N_1748);
nand U1863 (N_1863,N_1798,N_1750);
or U1864 (N_1864,N_1762,N_1730);
or U1865 (N_1865,N_1789,N_1732);
and U1866 (N_1866,N_1731,N_1780);
nor U1867 (N_1867,N_1787,N_1754);
and U1868 (N_1868,N_1796,N_1719);
nor U1869 (N_1869,N_1758,N_1737);
nor U1870 (N_1870,N_1704,N_1761);
nor U1871 (N_1871,N_1758,N_1711);
nand U1872 (N_1872,N_1716,N_1733);
and U1873 (N_1873,N_1781,N_1706);
xor U1874 (N_1874,N_1703,N_1702);
nand U1875 (N_1875,N_1791,N_1799);
xnor U1876 (N_1876,N_1793,N_1718);
xor U1877 (N_1877,N_1744,N_1785);
or U1878 (N_1878,N_1706,N_1762);
or U1879 (N_1879,N_1736,N_1721);
nor U1880 (N_1880,N_1776,N_1746);
or U1881 (N_1881,N_1749,N_1714);
nand U1882 (N_1882,N_1722,N_1753);
nor U1883 (N_1883,N_1741,N_1776);
and U1884 (N_1884,N_1747,N_1757);
xnor U1885 (N_1885,N_1728,N_1762);
xor U1886 (N_1886,N_1764,N_1779);
xor U1887 (N_1887,N_1795,N_1792);
xnor U1888 (N_1888,N_1779,N_1709);
xor U1889 (N_1889,N_1798,N_1776);
nand U1890 (N_1890,N_1739,N_1722);
nor U1891 (N_1891,N_1728,N_1709);
and U1892 (N_1892,N_1766,N_1725);
and U1893 (N_1893,N_1736,N_1767);
or U1894 (N_1894,N_1700,N_1711);
xor U1895 (N_1895,N_1772,N_1779);
nand U1896 (N_1896,N_1792,N_1744);
nor U1897 (N_1897,N_1702,N_1770);
and U1898 (N_1898,N_1730,N_1779);
or U1899 (N_1899,N_1787,N_1748);
or U1900 (N_1900,N_1879,N_1882);
xor U1901 (N_1901,N_1852,N_1886);
xor U1902 (N_1902,N_1851,N_1816);
xor U1903 (N_1903,N_1855,N_1895);
or U1904 (N_1904,N_1875,N_1831);
or U1905 (N_1905,N_1862,N_1848);
nor U1906 (N_1906,N_1865,N_1894);
and U1907 (N_1907,N_1802,N_1833);
xnor U1908 (N_1908,N_1843,N_1892);
nand U1909 (N_1909,N_1806,N_1844);
or U1910 (N_1910,N_1889,N_1869);
nor U1911 (N_1911,N_1840,N_1896);
nor U1912 (N_1912,N_1871,N_1813);
or U1913 (N_1913,N_1822,N_1881);
and U1914 (N_1914,N_1811,N_1846);
or U1915 (N_1915,N_1837,N_1810);
nand U1916 (N_1916,N_1899,N_1838);
nand U1917 (N_1917,N_1860,N_1803);
nor U1918 (N_1918,N_1842,N_1807);
and U1919 (N_1919,N_1870,N_1867);
or U1920 (N_1920,N_1821,N_1849);
or U1921 (N_1921,N_1858,N_1873);
and U1922 (N_1922,N_1830,N_1859);
and U1923 (N_1923,N_1808,N_1841);
nor U1924 (N_1924,N_1861,N_1839);
nand U1925 (N_1925,N_1887,N_1890);
or U1926 (N_1926,N_1850,N_1819);
and U1927 (N_1927,N_1868,N_1836);
nand U1928 (N_1928,N_1880,N_1888);
nor U1929 (N_1929,N_1872,N_1898);
xor U1930 (N_1930,N_1823,N_1829);
nor U1931 (N_1931,N_1812,N_1834);
xnor U1932 (N_1932,N_1883,N_1853);
xnor U1933 (N_1933,N_1826,N_1801);
xnor U1934 (N_1934,N_1815,N_1877);
nor U1935 (N_1935,N_1891,N_1863);
xor U1936 (N_1936,N_1827,N_1857);
nand U1937 (N_1937,N_1876,N_1828);
xor U1938 (N_1938,N_1884,N_1820);
xnor U1939 (N_1939,N_1835,N_1809);
or U1940 (N_1940,N_1885,N_1866);
nand U1941 (N_1941,N_1818,N_1893);
nor U1942 (N_1942,N_1854,N_1804);
xnor U1943 (N_1943,N_1878,N_1825);
nor U1944 (N_1944,N_1824,N_1874);
and U1945 (N_1945,N_1814,N_1832);
xor U1946 (N_1946,N_1856,N_1845);
or U1947 (N_1947,N_1805,N_1847);
nand U1948 (N_1948,N_1864,N_1817);
nand U1949 (N_1949,N_1897,N_1800);
xnor U1950 (N_1950,N_1809,N_1868);
or U1951 (N_1951,N_1803,N_1884);
nand U1952 (N_1952,N_1843,N_1874);
xnor U1953 (N_1953,N_1898,N_1887);
and U1954 (N_1954,N_1891,N_1819);
nor U1955 (N_1955,N_1829,N_1820);
or U1956 (N_1956,N_1890,N_1884);
xor U1957 (N_1957,N_1858,N_1887);
xnor U1958 (N_1958,N_1893,N_1839);
nor U1959 (N_1959,N_1897,N_1894);
nor U1960 (N_1960,N_1825,N_1803);
nor U1961 (N_1961,N_1809,N_1899);
nor U1962 (N_1962,N_1876,N_1820);
or U1963 (N_1963,N_1813,N_1834);
and U1964 (N_1964,N_1818,N_1806);
nand U1965 (N_1965,N_1843,N_1887);
nor U1966 (N_1966,N_1824,N_1827);
nor U1967 (N_1967,N_1824,N_1836);
or U1968 (N_1968,N_1831,N_1844);
nand U1969 (N_1969,N_1867,N_1872);
nor U1970 (N_1970,N_1867,N_1853);
and U1971 (N_1971,N_1882,N_1844);
and U1972 (N_1972,N_1899,N_1813);
nor U1973 (N_1973,N_1828,N_1806);
nand U1974 (N_1974,N_1897,N_1898);
xnor U1975 (N_1975,N_1884,N_1856);
or U1976 (N_1976,N_1835,N_1890);
nand U1977 (N_1977,N_1835,N_1807);
nand U1978 (N_1978,N_1833,N_1811);
or U1979 (N_1979,N_1805,N_1867);
and U1980 (N_1980,N_1818,N_1876);
nand U1981 (N_1981,N_1868,N_1860);
and U1982 (N_1982,N_1812,N_1849);
nor U1983 (N_1983,N_1883,N_1804);
or U1984 (N_1984,N_1848,N_1821);
and U1985 (N_1985,N_1806,N_1819);
nand U1986 (N_1986,N_1837,N_1881);
or U1987 (N_1987,N_1825,N_1894);
xor U1988 (N_1988,N_1859,N_1873);
and U1989 (N_1989,N_1837,N_1862);
and U1990 (N_1990,N_1831,N_1881);
xor U1991 (N_1991,N_1809,N_1858);
and U1992 (N_1992,N_1892,N_1890);
xor U1993 (N_1993,N_1869,N_1825);
nor U1994 (N_1994,N_1866,N_1820);
and U1995 (N_1995,N_1873,N_1895);
nand U1996 (N_1996,N_1805,N_1800);
nand U1997 (N_1997,N_1833,N_1894);
and U1998 (N_1998,N_1888,N_1803);
xnor U1999 (N_1999,N_1889,N_1853);
nor U2000 (N_2000,N_1940,N_1997);
nor U2001 (N_2001,N_1919,N_1956);
xor U2002 (N_2002,N_1907,N_1986);
nand U2003 (N_2003,N_1903,N_1924);
and U2004 (N_2004,N_1941,N_1916);
or U2005 (N_2005,N_1966,N_1948);
nor U2006 (N_2006,N_1909,N_1943);
nand U2007 (N_2007,N_1979,N_1954);
or U2008 (N_2008,N_1947,N_1944);
and U2009 (N_2009,N_1960,N_1958);
nor U2010 (N_2010,N_1901,N_1980);
nor U2011 (N_2011,N_1929,N_1964);
xor U2012 (N_2012,N_1982,N_1969);
and U2013 (N_2013,N_1923,N_1957);
and U2014 (N_2014,N_1955,N_1910);
nand U2015 (N_2015,N_1921,N_1928);
and U2016 (N_2016,N_1918,N_1987);
xnor U2017 (N_2017,N_1911,N_1912);
nand U2018 (N_2018,N_1936,N_1949);
or U2019 (N_2019,N_1959,N_1953);
or U2020 (N_2020,N_1968,N_1996);
nand U2021 (N_2021,N_1905,N_1937);
or U2022 (N_2022,N_1914,N_1970);
and U2023 (N_2023,N_1988,N_1971);
or U2024 (N_2024,N_1965,N_1917);
nor U2025 (N_2025,N_1934,N_1930);
or U2026 (N_2026,N_1961,N_1975);
or U2027 (N_2027,N_1981,N_1926);
nand U2028 (N_2028,N_1913,N_1974);
nor U2029 (N_2029,N_1922,N_1993);
nor U2030 (N_2030,N_1925,N_1927);
nor U2031 (N_2031,N_1994,N_1946);
nand U2032 (N_2032,N_1962,N_1963);
nand U2033 (N_2033,N_1931,N_1950);
xor U2034 (N_2034,N_1915,N_1977);
and U2035 (N_2035,N_1984,N_1952);
xnor U2036 (N_2036,N_1995,N_1933);
nor U2037 (N_2037,N_1989,N_1976);
xor U2038 (N_2038,N_1942,N_1932);
or U2039 (N_2039,N_1906,N_1990);
nand U2040 (N_2040,N_1983,N_1978);
xor U2041 (N_2041,N_1920,N_1998);
and U2042 (N_2042,N_1972,N_1902);
and U2043 (N_2043,N_1967,N_1939);
xnor U2044 (N_2044,N_1945,N_1908);
or U2045 (N_2045,N_1999,N_1985);
xor U2046 (N_2046,N_1991,N_1938);
nand U2047 (N_2047,N_1951,N_1973);
xnor U2048 (N_2048,N_1935,N_1900);
xnor U2049 (N_2049,N_1904,N_1992);
nand U2050 (N_2050,N_1916,N_1974);
and U2051 (N_2051,N_1934,N_1999);
or U2052 (N_2052,N_1940,N_1969);
and U2053 (N_2053,N_1939,N_1982);
or U2054 (N_2054,N_1907,N_1995);
or U2055 (N_2055,N_1987,N_1904);
or U2056 (N_2056,N_1992,N_1901);
xnor U2057 (N_2057,N_1991,N_1943);
nor U2058 (N_2058,N_1932,N_1988);
xnor U2059 (N_2059,N_1900,N_1964);
and U2060 (N_2060,N_1918,N_1952);
or U2061 (N_2061,N_1996,N_1961);
or U2062 (N_2062,N_1933,N_1966);
nand U2063 (N_2063,N_1961,N_1948);
nand U2064 (N_2064,N_1940,N_1929);
nor U2065 (N_2065,N_1955,N_1984);
nand U2066 (N_2066,N_1945,N_1900);
or U2067 (N_2067,N_1930,N_1955);
nand U2068 (N_2068,N_1959,N_1919);
nand U2069 (N_2069,N_1933,N_1929);
and U2070 (N_2070,N_1990,N_1983);
or U2071 (N_2071,N_1960,N_1954);
and U2072 (N_2072,N_1958,N_1920);
nor U2073 (N_2073,N_1977,N_1982);
and U2074 (N_2074,N_1990,N_1924);
nand U2075 (N_2075,N_1926,N_1921);
and U2076 (N_2076,N_1954,N_1984);
xor U2077 (N_2077,N_1945,N_1992);
nand U2078 (N_2078,N_1992,N_1962);
nor U2079 (N_2079,N_1937,N_1967);
and U2080 (N_2080,N_1982,N_1901);
and U2081 (N_2081,N_1950,N_1955);
xnor U2082 (N_2082,N_1941,N_1920);
or U2083 (N_2083,N_1997,N_1933);
nand U2084 (N_2084,N_1961,N_1954);
nor U2085 (N_2085,N_1980,N_1955);
nor U2086 (N_2086,N_1966,N_1975);
or U2087 (N_2087,N_1921,N_1948);
nand U2088 (N_2088,N_1904,N_1967);
nor U2089 (N_2089,N_1940,N_1982);
or U2090 (N_2090,N_1937,N_1914);
xor U2091 (N_2091,N_1935,N_1904);
xnor U2092 (N_2092,N_1900,N_1972);
nand U2093 (N_2093,N_1974,N_1971);
xor U2094 (N_2094,N_1976,N_1921);
nor U2095 (N_2095,N_1988,N_1916);
nor U2096 (N_2096,N_1921,N_1982);
nand U2097 (N_2097,N_1971,N_1986);
xnor U2098 (N_2098,N_1911,N_1925);
nor U2099 (N_2099,N_1957,N_1982);
xnor U2100 (N_2100,N_2042,N_2061);
or U2101 (N_2101,N_2076,N_2040);
or U2102 (N_2102,N_2086,N_2019);
nand U2103 (N_2103,N_2013,N_2082);
and U2104 (N_2104,N_2092,N_2056);
nor U2105 (N_2105,N_2090,N_2032);
nor U2106 (N_2106,N_2006,N_2023);
or U2107 (N_2107,N_2095,N_2059);
or U2108 (N_2108,N_2026,N_2087);
and U2109 (N_2109,N_2062,N_2081);
and U2110 (N_2110,N_2057,N_2080);
and U2111 (N_2111,N_2001,N_2065);
and U2112 (N_2112,N_2009,N_2016);
xnor U2113 (N_2113,N_2098,N_2071);
xor U2114 (N_2114,N_2067,N_2020);
and U2115 (N_2115,N_2091,N_2072);
and U2116 (N_2116,N_2097,N_2022);
nor U2117 (N_2117,N_2066,N_2075);
and U2118 (N_2118,N_2079,N_2003);
and U2119 (N_2119,N_2014,N_2054);
or U2120 (N_2120,N_2036,N_2045);
nand U2121 (N_2121,N_2039,N_2005);
and U2122 (N_2122,N_2094,N_2008);
nor U2123 (N_2123,N_2017,N_2063);
nor U2124 (N_2124,N_2078,N_2029);
and U2125 (N_2125,N_2046,N_2084);
and U2126 (N_2126,N_2038,N_2043);
xor U2127 (N_2127,N_2024,N_2033);
nor U2128 (N_2128,N_2050,N_2010);
xnor U2129 (N_2129,N_2030,N_2088);
or U2130 (N_2130,N_2047,N_2089);
xor U2131 (N_2131,N_2002,N_2053);
nor U2132 (N_2132,N_2069,N_2070);
and U2133 (N_2133,N_2015,N_2096);
nand U2134 (N_2134,N_2064,N_2041);
nand U2135 (N_2135,N_2048,N_2035);
and U2136 (N_2136,N_2044,N_2000);
xnor U2137 (N_2137,N_2074,N_2083);
nor U2138 (N_2138,N_2028,N_2012);
xor U2139 (N_2139,N_2049,N_2007);
or U2140 (N_2140,N_2055,N_2060);
and U2141 (N_2141,N_2034,N_2058);
xnor U2142 (N_2142,N_2011,N_2052);
or U2143 (N_2143,N_2037,N_2018);
and U2144 (N_2144,N_2021,N_2004);
xor U2145 (N_2145,N_2099,N_2093);
nand U2146 (N_2146,N_2073,N_2077);
xnor U2147 (N_2147,N_2085,N_2027);
xnor U2148 (N_2148,N_2031,N_2025);
nand U2149 (N_2149,N_2068,N_2051);
and U2150 (N_2150,N_2038,N_2073);
and U2151 (N_2151,N_2081,N_2044);
or U2152 (N_2152,N_2035,N_2062);
nor U2153 (N_2153,N_2009,N_2001);
xnor U2154 (N_2154,N_2035,N_2082);
and U2155 (N_2155,N_2061,N_2047);
nor U2156 (N_2156,N_2041,N_2047);
nand U2157 (N_2157,N_2014,N_2033);
nor U2158 (N_2158,N_2089,N_2002);
and U2159 (N_2159,N_2058,N_2060);
and U2160 (N_2160,N_2082,N_2000);
and U2161 (N_2161,N_2093,N_2085);
xnor U2162 (N_2162,N_2063,N_2099);
xnor U2163 (N_2163,N_2038,N_2034);
nand U2164 (N_2164,N_2054,N_2004);
and U2165 (N_2165,N_2036,N_2082);
and U2166 (N_2166,N_2029,N_2053);
nand U2167 (N_2167,N_2022,N_2079);
or U2168 (N_2168,N_2047,N_2052);
and U2169 (N_2169,N_2040,N_2033);
nor U2170 (N_2170,N_2026,N_2062);
or U2171 (N_2171,N_2033,N_2006);
xor U2172 (N_2172,N_2028,N_2029);
and U2173 (N_2173,N_2028,N_2067);
or U2174 (N_2174,N_2071,N_2053);
xnor U2175 (N_2175,N_2013,N_2092);
nor U2176 (N_2176,N_2069,N_2083);
nor U2177 (N_2177,N_2062,N_2096);
nand U2178 (N_2178,N_2084,N_2062);
and U2179 (N_2179,N_2083,N_2051);
or U2180 (N_2180,N_2020,N_2031);
or U2181 (N_2181,N_2072,N_2046);
and U2182 (N_2182,N_2007,N_2035);
or U2183 (N_2183,N_2032,N_2044);
nand U2184 (N_2184,N_2005,N_2019);
nand U2185 (N_2185,N_2092,N_2016);
or U2186 (N_2186,N_2048,N_2034);
xor U2187 (N_2187,N_2049,N_2068);
nand U2188 (N_2188,N_2014,N_2031);
or U2189 (N_2189,N_2081,N_2087);
xnor U2190 (N_2190,N_2041,N_2053);
and U2191 (N_2191,N_2096,N_2039);
xor U2192 (N_2192,N_2092,N_2063);
nor U2193 (N_2193,N_2063,N_2029);
nand U2194 (N_2194,N_2008,N_2061);
nand U2195 (N_2195,N_2071,N_2078);
or U2196 (N_2196,N_2086,N_2085);
or U2197 (N_2197,N_2050,N_2048);
xnor U2198 (N_2198,N_2048,N_2053);
and U2199 (N_2199,N_2071,N_2099);
xor U2200 (N_2200,N_2165,N_2149);
or U2201 (N_2201,N_2114,N_2137);
and U2202 (N_2202,N_2158,N_2167);
nand U2203 (N_2203,N_2124,N_2198);
and U2204 (N_2204,N_2142,N_2121);
nor U2205 (N_2205,N_2182,N_2104);
or U2206 (N_2206,N_2156,N_2177);
xnor U2207 (N_2207,N_2190,N_2191);
or U2208 (N_2208,N_2153,N_2196);
nor U2209 (N_2209,N_2123,N_2100);
and U2210 (N_2210,N_2143,N_2129);
or U2211 (N_2211,N_2157,N_2145);
nand U2212 (N_2212,N_2175,N_2146);
nand U2213 (N_2213,N_2172,N_2115);
and U2214 (N_2214,N_2128,N_2164);
or U2215 (N_2215,N_2116,N_2103);
nor U2216 (N_2216,N_2152,N_2132);
and U2217 (N_2217,N_2151,N_2102);
or U2218 (N_2218,N_2184,N_2193);
or U2219 (N_2219,N_2179,N_2140);
or U2220 (N_2220,N_2178,N_2147);
nand U2221 (N_2221,N_2195,N_2105);
nor U2222 (N_2222,N_2118,N_2117);
or U2223 (N_2223,N_2141,N_2136);
and U2224 (N_2224,N_2106,N_2181);
or U2225 (N_2225,N_2162,N_2159);
nor U2226 (N_2226,N_2180,N_2134);
nor U2227 (N_2227,N_2168,N_2107);
nor U2228 (N_2228,N_2160,N_2185);
nor U2229 (N_2229,N_2188,N_2108);
xnor U2230 (N_2230,N_2183,N_2148);
and U2231 (N_2231,N_2173,N_2144);
nand U2232 (N_2232,N_2186,N_2131);
nor U2233 (N_2233,N_2138,N_2176);
or U2234 (N_2234,N_2150,N_2154);
or U2235 (N_2235,N_2169,N_2199);
nand U2236 (N_2236,N_2187,N_2189);
nand U2237 (N_2237,N_2133,N_2126);
and U2238 (N_2238,N_2171,N_2110);
nand U2239 (N_2239,N_2166,N_2101);
nand U2240 (N_2240,N_2112,N_2135);
nand U2241 (N_2241,N_2120,N_2163);
and U2242 (N_2242,N_2170,N_2125);
xor U2243 (N_2243,N_2194,N_2155);
nor U2244 (N_2244,N_2174,N_2161);
nand U2245 (N_2245,N_2139,N_2192);
nor U2246 (N_2246,N_2119,N_2109);
nor U2247 (N_2247,N_2130,N_2111);
nand U2248 (N_2248,N_2113,N_2197);
nand U2249 (N_2249,N_2122,N_2127);
nand U2250 (N_2250,N_2142,N_2151);
nand U2251 (N_2251,N_2171,N_2132);
or U2252 (N_2252,N_2151,N_2125);
nor U2253 (N_2253,N_2168,N_2127);
nor U2254 (N_2254,N_2135,N_2106);
xnor U2255 (N_2255,N_2194,N_2135);
nor U2256 (N_2256,N_2181,N_2116);
nor U2257 (N_2257,N_2137,N_2199);
and U2258 (N_2258,N_2115,N_2125);
or U2259 (N_2259,N_2166,N_2183);
or U2260 (N_2260,N_2159,N_2118);
xnor U2261 (N_2261,N_2199,N_2138);
nand U2262 (N_2262,N_2153,N_2114);
xnor U2263 (N_2263,N_2191,N_2116);
nand U2264 (N_2264,N_2112,N_2158);
and U2265 (N_2265,N_2105,N_2126);
and U2266 (N_2266,N_2199,N_2102);
nand U2267 (N_2267,N_2153,N_2143);
nor U2268 (N_2268,N_2161,N_2168);
nor U2269 (N_2269,N_2157,N_2155);
xor U2270 (N_2270,N_2130,N_2155);
nand U2271 (N_2271,N_2173,N_2151);
and U2272 (N_2272,N_2178,N_2199);
xor U2273 (N_2273,N_2162,N_2127);
nor U2274 (N_2274,N_2162,N_2143);
nand U2275 (N_2275,N_2110,N_2140);
or U2276 (N_2276,N_2134,N_2160);
or U2277 (N_2277,N_2119,N_2147);
nand U2278 (N_2278,N_2180,N_2112);
or U2279 (N_2279,N_2184,N_2180);
xor U2280 (N_2280,N_2136,N_2194);
and U2281 (N_2281,N_2146,N_2154);
nand U2282 (N_2282,N_2101,N_2195);
or U2283 (N_2283,N_2168,N_2165);
and U2284 (N_2284,N_2183,N_2175);
and U2285 (N_2285,N_2172,N_2147);
nor U2286 (N_2286,N_2171,N_2119);
and U2287 (N_2287,N_2184,N_2125);
and U2288 (N_2288,N_2141,N_2146);
xor U2289 (N_2289,N_2184,N_2143);
xor U2290 (N_2290,N_2125,N_2196);
nand U2291 (N_2291,N_2115,N_2157);
nor U2292 (N_2292,N_2149,N_2146);
nand U2293 (N_2293,N_2132,N_2164);
xnor U2294 (N_2294,N_2141,N_2176);
xor U2295 (N_2295,N_2183,N_2117);
nand U2296 (N_2296,N_2103,N_2126);
and U2297 (N_2297,N_2198,N_2166);
and U2298 (N_2298,N_2102,N_2136);
nand U2299 (N_2299,N_2114,N_2185);
or U2300 (N_2300,N_2220,N_2201);
or U2301 (N_2301,N_2232,N_2217);
xor U2302 (N_2302,N_2277,N_2209);
xor U2303 (N_2303,N_2257,N_2250);
nand U2304 (N_2304,N_2278,N_2276);
and U2305 (N_2305,N_2244,N_2283);
and U2306 (N_2306,N_2290,N_2282);
and U2307 (N_2307,N_2236,N_2251);
and U2308 (N_2308,N_2242,N_2245);
nor U2309 (N_2309,N_2269,N_2254);
or U2310 (N_2310,N_2279,N_2203);
and U2311 (N_2311,N_2206,N_2240);
nand U2312 (N_2312,N_2284,N_2252);
and U2313 (N_2313,N_2299,N_2208);
or U2314 (N_2314,N_2261,N_2272);
xor U2315 (N_2315,N_2291,N_2259);
or U2316 (N_2316,N_2210,N_2298);
and U2317 (N_2317,N_2204,N_2215);
xor U2318 (N_2318,N_2213,N_2295);
nor U2319 (N_2319,N_2293,N_2268);
xor U2320 (N_2320,N_2207,N_2256);
nor U2321 (N_2321,N_2239,N_2292);
nand U2322 (N_2322,N_2285,N_2273);
nand U2323 (N_2323,N_2200,N_2267);
and U2324 (N_2324,N_2294,N_2297);
xor U2325 (N_2325,N_2264,N_2202);
or U2326 (N_2326,N_2255,N_2270);
xor U2327 (N_2327,N_2234,N_2262);
or U2328 (N_2328,N_2265,N_2289);
nand U2329 (N_2329,N_2275,N_2288);
nor U2330 (N_2330,N_2243,N_2235);
xnor U2331 (N_2331,N_2266,N_2260);
and U2332 (N_2332,N_2253,N_2230);
and U2333 (N_2333,N_2224,N_2246);
nor U2334 (N_2334,N_2271,N_2248);
nor U2335 (N_2335,N_2238,N_2222);
nor U2336 (N_2336,N_2263,N_2227);
and U2337 (N_2337,N_2214,N_2205);
nor U2338 (N_2338,N_2247,N_2218);
nor U2339 (N_2339,N_2223,N_2221);
nand U2340 (N_2340,N_2219,N_2280);
nor U2341 (N_2341,N_2286,N_2229);
or U2342 (N_2342,N_2237,N_2228);
or U2343 (N_2343,N_2231,N_2296);
xor U2344 (N_2344,N_2226,N_2216);
nor U2345 (N_2345,N_2249,N_2233);
nor U2346 (N_2346,N_2281,N_2212);
nor U2347 (N_2347,N_2211,N_2274);
and U2348 (N_2348,N_2258,N_2287);
nand U2349 (N_2349,N_2241,N_2225);
xnor U2350 (N_2350,N_2210,N_2235);
xor U2351 (N_2351,N_2270,N_2294);
nor U2352 (N_2352,N_2266,N_2209);
xnor U2353 (N_2353,N_2212,N_2223);
or U2354 (N_2354,N_2234,N_2287);
or U2355 (N_2355,N_2253,N_2276);
and U2356 (N_2356,N_2210,N_2232);
or U2357 (N_2357,N_2277,N_2272);
nor U2358 (N_2358,N_2285,N_2205);
and U2359 (N_2359,N_2273,N_2252);
nor U2360 (N_2360,N_2215,N_2202);
or U2361 (N_2361,N_2203,N_2204);
nand U2362 (N_2362,N_2266,N_2263);
xnor U2363 (N_2363,N_2256,N_2280);
nand U2364 (N_2364,N_2205,N_2280);
xnor U2365 (N_2365,N_2211,N_2293);
nand U2366 (N_2366,N_2284,N_2272);
nand U2367 (N_2367,N_2225,N_2243);
or U2368 (N_2368,N_2233,N_2242);
nor U2369 (N_2369,N_2220,N_2258);
nand U2370 (N_2370,N_2234,N_2267);
and U2371 (N_2371,N_2279,N_2270);
or U2372 (N_2372,N_2217,N_2292);
nand U2373 (N_2373,N_2286,N_2270);
and U2374 (N_2374,N_2298,N_2206);
and U2375 (N_2375,N_2280,N_2224);
nor U2376 (N_2376,N_2221,N_2290);
and U2377 (N_2377,N_2282,N_2278);
or U2378 (N_2378,N_2259,N_2220);
or U2379 (N_2379,N_2241,N_2283);
nand U2380 (N_2380,N_2242,N_2228);
xnor U2381 (N_2381,N_2205,N_2274);
nand U2382 (N_2382,N_2220,N_2206);
nor U2383 (N_2383,N_2264,N_2214);
nor U2384 (N_2384,N_2247,N_2225);
xor U2385 (N_2385,N_2245,N_2232);
nand U2386 (N_2386,N_2278,N_2224);
nor U2387 (N_2387,N_2215,N_2292);
nor U2388 (N_2388,N_2232,N_2273);
xor U2389 (N_2389,N_2223,N_2211);
and U2390 (N_2390,N_2277,N_2207);
and U2391 (N_2391,N_2275,N_2249);
xnor U2392 (N_2392,N_2282,N_2271);
nor U2393 (N_2393,N_2295,N_2243);
nor U2394 (N_2394,N_2285,N_2268);
xor U2395 (N_2395,N_2234,N_2296);
xnor U2396 (N_2396,N_2234,N_2283);
and U2397 (N_2397,N_2279,N_2242);
xnor U2398 (N_2398,N_2297,N_2279);
xnor U2399 (N_2399,N_2289,N_2204);
and U2400 (N_2400,N_2306,N_2308);
nor U2401 (N_2401,N_2390,N_2329);
nand U2402 (N_2402,N_2330,N_2394);
xor U2403 (N_2403,N_2303,N_2319);
or U2404 (N_2404,N_2346,N_2348);
nand U2405 (N_2405,N_2354,N_2388);
or U2406 (N_2406,N_2322,N_2324);
nand U2407 (N_2407,N_2326,N_2312);
nor U2408 (N_2408,N_2341,N_2344);
nor U2409 (N_2409,N_2379,N_2301);
or U2410 (N_2410,N_2321,N_2364);
nand U2411 (N_2411,N_2313,N_2389);
nand U2412 (N_2412,N_2356,N_2315);
nor U2413 (N_2413,N_2358,N_2304);
nand U2414 (N_2414,N_2333,N_2382);
and U2415 (N_2415,N_2342,N_2355);
xor U2416 (N_2416,N_2369,N_2334);
xnor U2417 (N_2417,N_2328,N_2373);
nor U2418 (N_2418,N_2338,N_2353);
or U2419 (N_2419,N_2383,N_2300);
and U2420 (N_2420,N_2366,N_2398);
nand U2421 (N_2421,N_2397,N_2316);
and U2422 (N_2422,N_2349,N_2370);
and U2423 (N_2423,N_2395,N_2331);
and U2424 (N_2424,N_2336,N_2343);
xnor U2425 (N_2425,N_2361,N_2302);
nand U2426 (N_2426,N_2337,N_2332);
or U2427 (N_2427,N_2362,N_2384);
or U2428 (N_2428,N_2386,N_2325);
nor U2429 (N_2429,N_2339,N_2335);
xor U2430 (N_2430,N_2352,N_2305);
xor U2431 (N_2431,N_2327,N_2314);
nand U2432 (N_2432,N_2323,N_2310);
xor U2433 (N_2433,N_2345,N_2318);
nand U2434 (N_2434,N_2385,N_2309);
nand U2435 (N_2435,N_2377,N_2376);
and U2436 (N_2436,N_2387,N_2378);
xor U2437 (N_2437,N_2367,N_2347);
nor U2438 (N_2438,N_2375,N_2359);
and U2439 (N_2439,N_2372,N_2311);
nor U2440 (N_2440,N_2360,N_2391);
and U2441 (N_2441,N_2357,N_2340);
nor U2442 (N_2442,N_2392,N_2363);
and U2443 (N_2443,N_2365,N_2374);
xnor U2444 (N_2444,N_2350,N_2351);
nor U2445 (N_2445,N_2317,N_2381);
and U2446 (N_2446,N_2368,N_2320);
and U2447 (N_2447,N_2393,N_2307);
nand U2448 (N_2448,N_2399,N_2371);
or U2449 (N_2449,N_2396,N_2380);
and U2450 (N_2450,N_2390,N_2368);
nand U2451 (N_2451,N_2369,N_2317);
nor U2452 (N_2452,N_2325,N_2363);
nor U2453 (N_2453,N_2393,N_2389);
and U2454 (N_2454,N_2320,N_2307);
or U2455 (N_2455,N_2378,N_2399);
nand U2456 (N_2456,N_2374,N_2318);
xor U2457 (N_2457,N_2331,N_2373);
xor U2458 (N_2458,N_2313,N_2329);
nand U2459 (N_2459,N_2306,N_2334);
and U2460 (N_2460,N_2310,N_2379);
nand U2461 (N_2461,N_2383,N_2367);
nand U2462 (N_2462,N_2322,N_2308);
nor U2463 (N_2463,N_2331,N_2398);
nand U2464 (N_2464,N_2301,N_2399);
and U2465 (N_2465,N_2392,N_2328);
nand U2466 (N_2466,N_2382,N_2308);
and U2467 (N_2467,N_2378,N_2312);
nor U2468 (N_2468,N_2320,N_2328);
or U2469 (N_2469,N_2334,N_2316);
nor U2470 (N_2470,N_2371,N_2316);
or U2471 (N_2471,N_2353,N_2301);
xnor U2472 (N_2472,N_2319,N_2316);
or U2473 (N_2473,N_2352,N_2362);
xnor U2474 (N_2474,N_2376,N_2321);
nor U2475 (N_2475,N_2303,N_2326);
and U2476 (N_2476,N_2375,N_2387);
or U2477 (N_2477,N_2399,N_2339);
nand U2478 (N_2478,N_2322,N_2384);
nand U2479 (N_2479,N_2376,N_2352);
nor U2480 (N_2480,N_2383,N_2376);
nor U2481 (N_2481,N_2306,N_2322);
or U2482 (N_2482,N_2352,N_2328);
and U2483 (N_2483,N_2352,N_2319);
nand U2484 (N_2484,N_2367,N_2304);
xnor U2485 (N_2485,N_2325,N_2337);
xnor U2486 (N_2486,N_2373,N_2308);
nor U2487 (N_2487,N_2302,N_2307);
and U2488 (N_2488,N_2364,N_2344);
xor U2489 (N_2489,N_2354,N_2306);
xor U2490 (N_2490,N_2378,N_2345);
nand U2491 (N_2491,N_2308,N_2366);
nor U2492 (N_2492,N_2390,N_2359);
nand U2493 (N_2493,N_2301,N_2320);
nor U2494 (N_2494,N_2319,N_2385);
xor U2495 (N_2495,N_2361,N_2325);
nor U2496 (N_2496,N_2323,N_2307);
xnor U2497 (N_2497,N_2332,N_2302);
and U2498 (N_2498,N_2382,N_2378);
nor U2499 (N_2499,N_2378,N_2367);
or U2500 (N_2500,N_2400,N_2479);
xnor U2501 (N_2501,N_2412,N_2495);
nor U2502 (N_2502,N_2474,N_2469);
xor U2503 (N_2503,N_2451,N_2409);
nand U2504 (N_2504,N_2423,N_2422);
nor U2505 (N_2505,N_2421,N_2468);
or U2506 (N_2506,N_2498,N_2406);
nor U2507 (N_2507,N_2436,N_2490);
xor U2508 (N_2508,N_2420,N_2488);
nand U2509 (N_2509,N_2411,N_2448);
nand U2510 (N_2510,N_2454,N_2483);
and U2511 (N_2511,N_2491,N_2418);
and U2512 (N_2512,N_2433,N_2492);
nor U2513 (N_2513,N_2416,N_2478);
or U2514 (N_2514,N_2489,N_2464);
and U2515 (N_2515,N_2494,N_2486);
nor U2516 (N_2516,N_2430,N_2467);
or U2517 (N_2517,N_2426,N_2499);
xnor U2518 (N_2518,N_2480,N_2481);
nand U2519 (N_2519,N_2405,N_2460);
nor U2520 (N_2520,N_2401,N_2424);
and U2521 (N_2521,N_2415,N_2475);
nor U2522 (N_2522,N_2459,N_2442);
nand U2523 (N_2523,N_2487,N_2439);
and U2524 (N_2524,N_2482,N_2404);
or U2525 (N_2525,N_2477,N_2493);
or U2526 (N_2526,N_2452,N_2458);
nand U2527 (N_2527,N_2413,N_2443);
or U2528 (N_2528,N_2461,N_2438);
and U2529 (N_2529,N_2435,N_2425);
nor U2530 (N_2530,N_2496,N_2408);
and U2531 (N_2531,N_2462,N_2437);
and U2532 (N_2532,N_2410,N_2497);
and U2533 (N_2533,N_2434,N_2402);
or U2534 (N_2534,N_2476,N_2466);
and U2535 (N_2535,N_2414,N_2419);
and U2536 (N_2536,N_2455,N_2463);
or U2537 (N_2537,N_2447,N_2450);
and U2538 (N_2538,N_2444,N_2471);
and U2539 (N_2539,N_2446,N_2457);
or U2540 (N_2540,N_2427,N_2453);
or U2541 (N_2541,N_2445,N_2449);
nor U2542 (N_2542,N_2417,N_2431);
and U2543 (N_2543,N_2472,N_2485);
and U2544 (N_2544,N_2441,N_2465);
nand U2545 (N_2545,N_2484,N_2432);
nor U2546 (N_2546,N_2428,N_2440);
nor U2547 (N_2547,N_2473,N_2429);
or U2548 (N_2548,N_2470,N_2456);
nor U2549 (N_2549,N_2403,N_2407);
and U2550 (N_2550,N_2466,N_2463);
and U2551 (N_2551,N_2484,N_2490);
nand U2552 (N_2552,N_2415,N_2484);
nand U2553 (N_2553,N_2434,N_2446);
xor U2554 (N_2554,N_2471,N_2448);
and U2555 (N_2555,N_2458,N_2429);
xnor U2556 (N_2556,N_2496,N_2448);
nand U2557 (N_2557,N_2451,N_2473);
or U2558 (N_2558,N_2470,N_2440);
and U2559 (N_2559,N_2418,N_2431);
and U2560 (N_2560,N_2498,N_2488);
or U2561 (N_2561,N_2471,N_2413);
nor U2562 (N_2562,N_2420,N_2427);
xor U2563 (N_2563,N_2444,N_2498);
xnor U2564 (N_2564,N_2452,N_2433);
nand U2565 (N_2565,N_2412,N_2491);
and U2566 (N_2566,N_2488,N_2452);
or U2567 (N_2567,N_2452,N_2446);
and U2568 (N_2568,N_2422,N_2479);
nand U2569 (N_2569,N_2403,N_2496);
and U2570 (N_2570,N_2495,N_2497);
xnor U2571 (N_2571,N_2407,N_2406);
nand U2572 (N_2572,N_2442,N_2447);
xnor U2573 (N_2573,N_2429,N_2490);
and U2574 (N_2574,N_2471,N_2406);
nand U2575 (N_2575,N_2462,N_2488);
xnor U2576 (N_2576,N_2487,N_2438);
or U2577 (N_2577,N_2452,N_2496);
nor U2578 (N_2578,N_2464,N_2409);
nand U2579 (N_2579,N_2455,N_2416);
xnor U2580 (N_2580,N_2443,N_2427);
xor U2581 (N_2581,N_2466,N_2470);
nand U2582 (N_2582,N_2437,N_2412);
and U2583 (N_2583,N_2462,N_2421);
xnor U2584 (N_2584,N_2488,N_2444);
nand U2585 (N_2585,N_2464,N_2402);
and U2586 (N_2586,N_2493,N_2478);
xnor U2587 (N_2587,N_2437,N_2467);
nand U2588 (N_2588,N_2418,N_2498);
or U2589 (N_2589,N_2457,N_2403);
nor U2590 (N_2590,N_2481,N_2464);
nor U2591 (N_2591,N_2471,N_2458);
nand U2592 (N_2592,N_2457,N_2451);
and U2593 (N_2593,N_2453,N_2424);
nor U2594 (N_2594,N_2466,N_2448);
nor U2595 (N_2595,N_2437,N_2423);
nand U2596 (N_2596,N_2418,N_2447);
xnor U2597 (N_2597,N_2484,N_2402);
xnor U2598 (N_2598,N_2416,N_2418);
and U2599 (N_2599,N_2435,N_2480);
or U2600 (N_2600,N_2595,N_2513);
or U2601 (N_2601,N_2549,N_2547);
nor U2602 (N_2602,N_2556,N_2531);
and U2603 (N_2603,N_2581,N_2582);
nor U2604 (N_2604,N_2597,N_2544);
nor U2605 (N_2605,N_2598,N_2553);
xor U2606 (N_2606,N_2555,N_2593);
nor U2607 (N_2607,N_2523,N_2580);
nor U2608 (N_2608,N_2563,N_2583);
and U2609 (N_2609,N_2514,N_2548);
nand U2610 (N_2610,N_2565,N_2503);
nand U2611 (N_2611,N_2517,N_2594);
xnor U2612 (N_2612,N_2568,N_2530);
nor U2613 (N_2613,N_2520,N_2518);
or U2614 (N_2614,N_2509,N_2529);
xnor U2615 (N_2615,N_2552,N_2561);
nand U2616 (N_2616,N_2502,N_2510);
and U2617 (N_2617,N_2500,N_2579);
xor U2618 (N_2618,N_2526,N_2539);
or U2619 (N_2619,N_2507,N_2542);
xnor U2620 (N_2620,N_2586,N_2540);
or U2621 (N_2621,N_2576,N_2562);
or U2622 (N_2622,N_2559,N_2537);
nor U2623 (N_2623,N_2578,N_2599);
and U2624 (N_2624,N_2541,N_2588);
and U2625 (N_2625,N_2558,N_2525);
xor U2626 (N_2626,N_2546,N_2560);
xnor U2627 (N_2627,N_2590,N_2564);
nand U2628 (N_2628,N_2521,N_2522);
xor U2629 (N_2629,N_2527,N_2516);
nand U2630 (N_2630,N_2575,N_2591);
xnor U2631 (N_2631,N_2534,N_2596);
and U2632 (N_2632,N_2524,N_2567);
xor U2633 (N_2633,N_2554,N_2566);
and U2634 (N_2634,N_2573,N_2589);
or U2635 (N_2635,N_2501,N_2587);
nor U2636 (N_2636,N_2528,N_2569);
nor U2637 (N_2637,N_2515,N_2572);
xnor U2638 (N_2638,N_2543,N_2574);
nand U2639 (N_2639,N_2519,N_2506);
or U2640 (N_2640,N_2508,N_2557);
and U2641 (N_2641,N_2536,N_2571);
nand U2642 (N_2642,N_2533,N_2584);
nand U2643 (N_2643,N_2505,N_2532);
or U2644 (N_2644,N_2511,N_2577);
nand U2645 (N_2645,N_2512,N_2535);
nand U2646 (N_2646,N_2551,N_2570);
nand U2647 (N_2647,N_2538,N_2504);
nand U2648 (N_2648,N_2545,N_2585);
and U2649 (N_2649,N_2592,N_2550);
nand U2650 (N_2650,N_2513,N_2551);
xor U2651 (N_2651,N_2547,N_2529);
nor U2652 (N_2652,N_2570,N_2592);
xnor U2653 (N_2653,N_2554,N_2543);
xor U2654 (N_2654,N_2597,N_2545);
or U2655 (N_2655,N_2522,N_2529);
and U2656 (N_2656,N_2531,N_2595);
nor U2657 (N_2657,N_2532,N_2588);
and U2658 (N_2658,N_2585,N_2566);
nand U2659 (N_2659,N_2563,N_2537);
nor U2660 (N_2660,N_2541,N_2567);
and U2661 (N_2661,N_2563,N_2596);
nor U2662 (N_2662,N_2515,N_2540);
and U2663 (N_2663,N_2557,N_2510);
xnor U2664 (N_2664,N_2575,N_2535);
and U2665 (N_2665,N_2513,N_2520);
xor U2666 (N_2666,N_2513,N_2501);
or U2667 (N_2667,N_2504,N_2505);
and U2668 (N_2668,N_2548,N_2565);
nor U2669 (N_2669,N_2571,N_2555);
or U2670 (N_2670,N_2519,N_2527);
or U2671 (N_2671,N_2538,N_2566);
xnor U2672 (N_2672,N_2545,N_2522);
nand U2673 (N_2673,N_2571,N_2520);
nand U2674 (N_2674,N_2586,N_2526);
nor U2675 (N_2675,N_2580,N_2520);
and U2676 (N_2676,N_2518,N_2553);
nand U2677 (N_2677,N_2502,N_2565);
xor U2678 (N_2678,N_2556,N_2551);
or U2679 (N_2679,N_2520,N_2548);
or U2680 (N_2680,N_2504,N_2541);
and U2681 (N_2681,N_2593,N_2578);
or U2682 (N_2682,N_2534,N_2519);
nand U2683 (N_2683,N_2589,N_2531);
xnor U2684 (N_2684,N_2567,N_2543);
or U2685 (N_2685,N_2533,N_2554);
nor U2686 (N_2686,N_2598,N_2508);
nand U2687 (N_2687,N_2517,N_2533);
nand U2688 (N_2688,N_2532,N_2581);
nand U2689 (N_2689,N_2528,N_2526);
or U2690 (N_2690,N_2514,N_2596);
nand U2691 (N_2691,N_2586,N_2511);
nor U2692 (N_2692,N_2542,N_2559);
nor U2693 (N_2693,N_2576,N_2587);
or U2694 (N_2694,N_2539,N_2596);
and U2695 (N_2695,N_2545,N_2534);
nor U2696 (N_2696,N_2573,N_2540);
nand U2697 (N_2697,N_2504,N_2560);
nor U2698 (N_2698,N_2581,N_2556);
and U2699 (N_2699,N_2546,N_2509);
xnor U2700 (N_2700,N_2606,N_2653);
xor U2701 (N_2701,N_2646,N_2608);
xnor U2702 (N_2702,N_2613,N_2654);
and U2703 (N_2703,N_2655,N_2677);
xnor U2704 (N_2704,N_2679,N_2621);
xnor U2705 (N_2705,N_2672,N_2673);
nand U2706 (N_2706,N_2604,N_2636);
nand U2707 (N_2707,N_2625,N_2682);
or U2708 (N_2708,N_2647,N_2684);
or U2709 (N_2709,N_2631,N_2670);
nand U2710 (N_2710,N_2652,N_2609);
xor U2711 (N_2711,N_2618,N_2615);
and U2712 (N_2712,N_2664,N_2602);
nor U2713 (N_2713,N_2690,N_2661);
nand U2714 (N_2714,N_2641,N_2614);
nor U2715 (N_2715,N_2603,N_2628);
nor U2716 (N_2716,N_2619,N_2666);
nor U2717 (N_2717,N_2697,N_2627);
xnor U2718 (N_2718,N_2637,N_2688);
xor U2719 (N_2719,N_2650,N_2651);
or U2720 (N_2720,N_2639,N_2668);
and U2721 (N_2721,N_2695,N_2676);
or U2722 (N_2722,N_2671,N_2674);
nor U2723 (N_2723,N_2638,N_2605);
nand U2724 (N_2724,N_2642,N_2691);
nor U2725 (N_2725,N_2665,N_2622);
and U2726 (N_2726,N_2626,N_2610);
nor U2727 (N_2727,N_2683,N_2623);
nand U2728 (N_2728,N_2669,N_2624);
nand U2729 (N_2729,N_2660,N_2675);
and U2730 (N_2730,N_2698,N_2630);
or U2731 (N_2731,N_2617,N_2645);
or U2732 (N_2732,N_2632,N_2680);
nor U2733 (N_2733,N_2640,N_2696);
nand U2734 (N_2734,N_2667,N_2633);
xnor U2735 (N_2735,N_2687,N_2612);
nand U2736 (N_2736,N_2678,N_2620);
nor U2737 (N_2737,N_2649,N_2635);
xnor U2738 (N_2738,N_2611,N_2658);
or U2739 (N_2739,N_2659,N_2600);
xor U2740 (N_2740,N_2656,N_2681);
xor U2741 (N_2741,N_2648,N_2663);
or U2742 (N_2742,N_2685,N_2686);
nand U2743 (N_2743,N_2644,N_2692);
nand U2744 (N_2744,N_2657,N_2699);
and U2745 (N_2745,N_2662,N_2616);
or U2746 (N_2746,N_2634,N_2693);
xnor U2747 (N_2747,N_2601,N_2694);
and U2748 (N_2748,N_2629,N_2607);
and U2749 (N_2749,N_2689,N_2643);
nand U2750 (N_2750,N_2608,N_2616);
and U2751 (N_2751,N_2613,N_2617);
xor U2752 (N_2752,N_2628,N_2600);
nor U2753 (N_2753,N_2654,N_2691);
nand U2754 (N_2754,N_2666,N_2651);
xor U2755 (N_2755,N_2661,N_2695);
nor U2756 (N_2756,N_2613,N_2606);
nand U2757 (N_2757,N_2629,N_2646);
and U2758 (N_2758,N_2645,N_2649);
or U2759 (N_2759,N_2699,N_2674);
xor U2760 (N_2760,N_2668,N_2633);
or U2761 (N_2761,N_2659,N_2637);
xor U2762 (N_2762,N_2688,N_2693);
nor U2763 (N_2763,N_2609,N_2658);
and U2764 (N_2764,N_2663,N_2696);
or U2765 (N_2765,N_2691,N_2639);
and U2766 (N_2766,N_2612,N_2670);
nor U2767 (N_2767,N_2628,N_2648);
xor U2768 (N_2768,N_2631,N_2676);
nor U2769 (N_2769,N_2605,N_2690);
nor U2770 (N_2770,N_2698,N_2674);
xor U2771 (N_2771,N_2618,N_2691);
or U2772 (N_2772,N_2679,N_2672);
nor U2773 (N_2773,N_2673,N_2633);
nor U2774 (N_2774,N_2649,N_2692);
and U2775 (N_2775,N_2653,N_2675);
and U2776 (N_2776,N_2676,N_2681);
nor U2777 (N_2777,N_2606,N_2649);
or U2778 (N_2778,N_2673,N_2631);
nand U2779 (N_2779,N_2690,N_2682);
nand U2780 (N_2780,N_2670,N_2682);
nor U2781 (N_2781,N_2609,N_2622);
nand U2782 (N_2782,N_2646,N_2667);
nand U2783 (N_2783,N_2697,N_2681);
nand U2784 (N_2784,N_2685,N_2695);
nand U2785 (N_2785,N_2609,N_2621);
nor U2786 (N_2786,N_2640,N_2658);
xnor U2787 (N_2787,N_2609,N_2690);
nor U2788 (N_2788,N_2663,N_2608);
and U2789 (N_2789,N_2638,N_2603);
or U2790 (N_2790,N_2620,N_2675);
and U2791 (N_2791,N_2666,N_2664);
xor U2792 (N_2792,N_2699,N_2652);
nand U2793 (N_2793,N_2621,N_2690);
nand U2794 (N_2794,N_2683,N_2603);
and U2795 (N_2795,N_2644,N_2613);
or U2796 (N_2796,N_2635,N_2604);
xnor U2797 (N_2797,N_2645,N_2606);
xnor U2798 (N_2798,N_2663,N_2619);
nand U2799 (N_2799,N_2631,N_2634);
nand U2800 (N_2800,N_2761,N_2748);
and U2801 (N_2801,N_2733,N_2792);
nand U2802 (N_2802,N_2723,N_2711);
or U2803 (N_2803,N_2778,N_2726);
or U2804 (N_2804,N_2776,N_2734);
and U2805 (N_2805,N_2714,N_2762);
nand U2806 (N_2806,N_2757,N_2750);
nand U2807 (N_2807,N_2797,N_2755);
xor U2808 (N_2808,N_2764,N_2717);
nand U2809 (N_2809,N_2704,N_2788);
and U2810 (N_2810,N_2721,N_2722);
or U2811 (N_2811,N_2708,N_2705);
and U2812 (N_2812,N_2775,N_2703);
nand U2813 (N_2813,N_2732,N_2765);
nor U2814 (N_2814,N_2749,N_2707);
nand U2815 (N_2815,N_2766,N_2742);
xnor U2816 (N_2816,N_2740,N_2796);
or U2817 (N_2817,N_2741,N_2710);
or U2818 (N_2818,N_2728,N_2798);
or U2819 (N_2819,N_2747,N_2702);
and U2820 (N_2820,N_2771,N_2712);
xnor U2821 (N_2821,N_2727,N_2752);
nand U2822 (N_2822,N_2791,N_2706);
nor U2823 (N_2823,N_2774,N_2751);
xor U2824 (N_2824,N_2730,N_2782);
xor U2825 (N_2825,N_2767,N_2737);
or U2826 (N_2826,N_2746,N_2719);
xor U2827 (N_2827,N_2779,N_2738);
nand U2828 (N_2828,N_2786,N_2799);
or U2829 (N_2829,N_2773,N_2787);
nor U2830 (N_2830,N_2718,N_2790);
or U2831 (N_2831,N_2735,N_2743);
xnor U2832 (N_2832,N_2729,N_2758);
or U2833 (N_2833,N_2793,N_2772);
nand U2834 (N_2834,N_2731,N_2716);
nand U2835 (N_2835,N_2744,N_2725);
xor U2836 (N_2836,N_2763,N_2724);
or U2837 (N_2837,N_2769,N_2736);
nor U2838 (N_2838,N_2760,N_2754);
or U2839 (N_2839,N_2720,N_2781);
nand U2840 (N_2840,N_2700,N_2795);
nand U2841 (N_2841,N_2745,N_2739);
and U2842 (N_2842,N_2770,N_2753);
and U2843 (N_2843,N_2794,N_2785);
xnor U2844 (N_2844,N_2715,N_2768);
xor U2845 (N_2845,N_2759,N_2713);
or U2846 (N_2846,N_2701,N_2756);
or U2847 (N_2847,N_2784,N_2780);
or U2848 (N_2848,N_2783,N_2777);
and U2849 (N_2849,N_2789,N_2709);
nand U2850 (N_2850,N_2779,N_2725);
or U2851 (N_2851,N_2754,N_2755);
nand U2852 (N_2852,N_2750,N_2778);
xnor U2853 (N_2853,N_2748,N_2774);
xor U2854 (N_2854,N_2788,N_2702);
nor U2855 (N_2855,N_2720,N_2729);
xnor U2856 (N_2856,N_2716,N_2762);
xor U2857 (N_2857,N_2770,N_2760);
xnor U2858 (N_2858,N_2741,N_2732);
and U2859 (N_2859,N_2723,N_2746);
xor U2860 (N_2860,N_2720,N_2700);
or U2861 (N_2861,N_2761,N_2794);
xor U2862 (N_2862,N_2777,N_2769);
nand U2863 (N_2863,N_2788,N_2739);
nor U2864 (N_2864,N_2749,N_2734);
xnor U2865 (N_2865,N_2738,N_2736);
nand U2866 (N_2866,N_2775,N_2779);
nand U2867 (N_2867,N_2763,N_2768);
and U2868 (N_2868,N_2785,N_2727);
and U2869 (N_2869,N_2767,N_2721);
and U2870 (N_2870,N_2783,N_2706);
and U2871 (N_2871,N_2772,N_2702);
and U2872 (N_2872,N_2798,N_2714);
and U2873 (N_2873,N_2726,N_2701);
nor U2874 (N_2874,N_2704,N_2731);
nor U2875 (N_2875,N_2745,N_2768);
xor U2876 (N_2876,N_2748,N_2710);
xnor U2877 (N_2877,N_2786,N_2782);
nand U2878 (N_2878,N_2787,N_2768);
xor U2879 (N_2879,N_2752,N_2751);
and U2880 (N_2880,N_2762,N_2731);
and U2881 (N_2881,N_2765,N_2749);
nand U2882 (N_2882,N_2761,N_2730);
or U2883 (N_2883,N_2703,N_2734);
nand U2884 (N_2884,N_2738,N_2718);
nor U2885 (N_2885,N_2735,N_2755);
or U2886 (N_2886,N_2709,N_2776);
nand U2887 (N_2887,N_2754,N_2784);
xor U2888 (N_2888,N_2728,N_2783);
nor U2889 (N_2889,N_2747,N_2796);
nand U2890 (N_2890,N_2704,N_2750);
nand U2891 (N_2891,N_2785,N_2751);
nand U2892 (N_2892,N_2741,N_2797);
nor U2893 (N_2893,N_2736,N_2722);
nand U2894 (N_2894,N_2706,N_2705);
nor U2895 (N_2895,N_2705,N_2799);
or U2896 (N_2896,N_2789,N_2724);
and U2897 (N_2897,N_2787,N_2742);
or U2898 (N_2898,N_2774,N_2764);
xnor U2899 (N_2899,N_2775,N_2776);
nand U2900 (N_2900,N_2816,N_2810);
and U2901 (N_2901,N_2883,N_2880);
nand U2902 (N_2902,N_2875,N_2856);
and U2903 (N_2903,N_2825,N_2867);
or U2904 (N_2904,N_2819,N_2863);
xor U2905 (N_2905,N_2820,N_2812);
nor U2906 (N_2906,N_2841,N_2852);
or U2907 (N_2907,N_2865,N_2824);
xnor U2908 (N_2908,N_2871,N_2803);
nand U2909 (N_2909,N_2831,N_2848);
nor U2910 (N_2910,N_2832,N_2872);
or U2911 (N_2911,N_2813,N_2862);
nor U2912 (N_2912,N_2879,N_2817);
or U2913 (N_2913,N_2853,N_2881);
and U2914 (N_2914,N_2894,N_2833);
nand U2915 (N_2915,N_2839,N_2829);
nand U2916 (N_2916,N_2847,N_2830);
or U2917 (N_2917,N_2844,N_2861);
nand U2918 (N_2918,N_2842,N_2873);
nor U2919 (N_2919,N_2874,N_2887);
xor U2920 (N_2920,N_2850,N_2814);
nor U2921 (N_2921,N_2869,N_2870);
nor U2922 (N_2922,N_2866,N_2818);
or U2923 (N_2923,N_2892,N_2860);
or U2924 (N_2924,N_2800,N_2859);
nand U2925 (N_2925,N_2849,N_2827);
xnor U2926 (N_2926,N_2806,N_2837);
and U2927 (N_2927,N_2890,N_2885);
nor U2928 (N_2928,N_2822,N_2882);
and U2929 (N_2929,N_2835,N_2828);
and U2930 (N_2930,N_2807,N_2899);
nor U2931 (N_2931,N_2815,N_2895);
nand U2932 (N_2932,N_2896,N_2889);
nand U2933 (N_2933,N_2811,N_2878);
and U2934 (N_2934,N_2834,N_2851);
nand U2935 (N_2935,N_2821,N_2838);
or U2936 (N_2936,N_2802,N_2840);
xor U2937 (N_2937,N_2804,N_2876);
or U2938 (N_2938,N_2893,N_2843);
and U2939 (N_2939,N_2855,N_2809);
and U2940 (N_2940,N_2801,N_2898);
nand U2941 (N_2941,N_2877,N_2891);
nor U2942 (N_2942,N_2805,N_2858);
xnor U2943 (N_2943,N_2864,N_2854);
xor U2944 (N_2944,N_2857,N_2845);
xnor U2945 (N_2945,N_2846,N_2884);
nor U2946 (N_2946,N_2826,N_2886);
and U2947 (N_2947,N_2836,N_2888);
or U2948 (N_2948,N_2868,N_2823);
xnor U2949 (N_2949,N_2897,N_2808);
xnor U2950 (N_2950,N_2881,N_2806);
nor U2951 (N_2951,N_2898,N_2840);
or U2952 (N_2952,N_2892,N_2885);
nor U2953 (N_2953,N_2872,N_2830);
or U2954 (N_2954,N_2817,N_2885);
nor U2955 (N_2955,N_2800,N_2867);
xor U2956 (N_2956,N_2873,N_2867);
or U2957 (N_2957,N_2803,N_2884);
and U2958 (N_2958,N_2860,N_2893);
nand U2959 (N_2959,N_2850,N_2857);
nand U2960 (N_2960,N_2869,N_2813);
nor U2961 (N_2961,N_2897,N_2894);
xnor U2962 (N_2962,N_2809,N_2863);
and U2963 (N_2963,N_2856,N_2849);
and U2964 (N_2964,N_2895,N_2854);
nand U2965 (N_2965,N_2833,N_2818);
and U2966 (N_2966,N_2861,N_2830);
xnor U2967 (N_2967,N_2804,N_2802);
or U2968 (N_2968,N_2849,N_2870);
and U2969 (N_2969,N_2817,N_2867);
xor U2970 (N_2970,N_2897,N_2874);
xnor U2971 (N_2971,N_2866,N_2857);
xor U2972 (N_2972,N_2840,N_2844);
and U2973 (N_2973,N_2888,N_2806);
and U2974 (N_2974,N_2877,N_2811);
and U2975 (N_2975,N_2830,N_2891);
nor U2976 (N_2976,N_2864,N_2800);
and U2977 (N_2977,N_2885,N_2888);
nor U2978 (N_2978,N_2855,N_2822);
and U2979 (N_2979,N_2870,N_2817);
nor U2980 (N_2980,N_2887,N_2846);
xor U2981 (N_2981,N_2802,N_2868);
or U2982 (N_2982,N_2855,N_2817);
nor U2983 (N_2983,N_2889,N_2817);
and U2984 (N_2984,N_2845,N_2876);
nand U2985 (N_2985,N_2805,N_2832);
and U2986 (N_2986,N_2808,N_2833);
and U2987 (N_2987,N_2898,N_2848);
xor U2988 (N_2988,N_2811,N_2808);
nand U2989 (N_2989,N_2893,N_2856);
xor U2990 (N_2990,N_2876,N_2869);
nor U2991 (N_2991,N_2830,N_2892);
or U2992 (N_2992,N_2868,N_2833);
nor U2993 (N_2993,N_2856,N_2861);
and U2994 (N_2994,N_2802,N_2849);
nor U2995 (N_2995,N_2842,N_2808);
and U2996 (N_2996,N_2836,N_2857);
xor U2997 (N_2997,N_2809,N_2880);
xor U2998 (N_2998,N_2868,N_2803);
nand U2999 (N_2999,N_2856,N_2848);
nor U3000 (N_3000,N_2976,N_2925);
and U3001 (N_3001,N_2965,N_2908);
nand U3002 (N_3002,N_2955,N_2972);
nand U3003 (N_3003,N_2924,N_2941);
nor U3004 (N_3004,N_2985,N_2979);
nand U3005 (N_3005,N_2969,N_2993);
xnor U3006 (N_3006,N_2942,N_2905);
nand U3007 (N_3007,N_2921,N_2975);
nor U3008 (N_3008,N_2920,N_2981);
and U3009 (N_3009,N_2961,N_2947);
or U3010 (N_3010,N_2938,N_2919);
or U3011 (N_3011,N_2923,N_2903);
nor U3012 (N_3012,N_2967,N_2987);
or U3013 (N_3013,N_2915,N_2988);
nor U3014 (N_3014,N_2926,N_2999);
and U3015 (N_3015,N_2962,N_2940);
and U3016 (N_3016,N_2964,N_2950);
or U3017 (N_3017,N_2902,N_2968);
nor U3018 (N_3018,N_2939,N_2970);
or U3019 (N_3019,N_2907,N_2954);
and U3020 (N_3020,N_2945,N_2960);
nand U3021 (N_3021,N_2997,N_2912);
xnor U3022 (N_3022,N_2918,N_2971);
or U3023 (N_3023,N_2934,N_2930);
nor U3024 (N_3024,N_2906,N_2909);
or U3025 (N_3025,N_2914,N_2978);
or U3026 (N_3026,N_2913,N_2910);
and U3027 (N_3027,N_2929,N_2928);
nand U3028 (N_3028,N_2935,N_2984);
nor U3029 (N_3029,N_2952,N_2901);
and U3030 (N_3030,N_2922,N_2957);
xnor U3031 (N_3031,N_2958,N_2904);
or U3032 (N_3032,N_2900,N_2990);
xor U3033 (N_3033,N_2973,N_2977);
nor U3034 (N_3034,N_2949,N_2916);
nor U3035 (N_3035,N_2998,N_2994);
or U3036 (N_3036,N_2948,N_2959);
and U3037 (N_3037,N_2937,N_2992);
or U3038 (N_3038,N_2917,N_2932);
xor U3039 (N_3039,N_2982,N_2936);
and U3040 (N_3040,N_2963,N_2989);
and U3041 (N_3041,N_2996,N_2943);
and U3042 (N_3042,N_2983,N_2995);
nand U3043 (N_3043,N_2927,N_2980);
nor U3044 (N_3044,N_2966,N_2931);
nor U3045 (N_3045,N_2944,N_2953);
or U3046 (N_3046,N_2951,N_2946);
and U3047 (N_3047,N_2956,N_2974);
or U3048 (N_3048,N_2986,N_2933);
or U3049 (N_3049,N_2991,N_2911);
nand U3050 (N_3050,N_2991,N_2946);
xor U3051 (N_3051,N_2962,N_2900);
or U3052 (N_3052,N_2953,N_2917);
nor U3053 (N_3053,N_2943,N_2954);
and U3054 (N_3054,N_2949,N_2939);
and U3055 (N_3055,N_2965,N_2987);
and U3056 (N_3056,N_2982,N_2922);
xnor U3057 (N_3057,N_2997,N_2963);
xnor U3058 (N_3058,N_2988,N_2972);
nand U3059 (N_3059,N_2959,N_2924);
or U3060 (N_3060,N_2911,N_2958);
xor U3061 (N_3061,N_2979,N_2986);
nand U3062 (N_3062,N_2918,N_2985);
and U3063 (N_3063,N_2973,N_2955);
and U3064 (N_3064,N_2953,N_2904);
nand U3065 (N_3065,N_2940,N_2976);
nand U3066 (N_3066,N_2931,N_2900);
xor U3067 (N_3067,N_2994,N_2966);
nor U3068 (N_3068,N_2993,N_2979);
xnor U3069 (N_3069,N_2930,N_2967);
nand U3070 (N_3070,N_2908,N_2929);
or U3071 (N_3071,N_2910,N_2917);
xor U3072 (N_3072,N_2933,N_2957);
and U3073 (N_3073,N_2935,N_2921);
nor U3074 (N_3074,N_2963,N_2987);
and U3075 (N_3075,N_2994,N_2952);
xnor U3076 (N_3076,N_2981,N_2996);
nor U3077 (N_3077,N_2997,N_2941);
and U3078 (N_3078,N_2909,N_2963);
nand U3079 (N_3079,N_2947,N_2942);
or U3080 (N_3080,N_2967,N_2915);
xnor U3081 (N_3081,N_2980,N_2934);
nor U3082 (N_3082,N_2963,N_2901);
nand U3083 (N_3083,N_2951,N_2913);
nor U3084 (N_3084,N_2983,N_2958);
or U3085 (N_3085,N_2928,N_2963);
xnor U3086 (N_3086,N_2936,N_2914);
nor U3087 (N_3087,N_2957,N_2949);
nand U3088 (N_3088,N_2935,N_2916);
xnor U3089 (N_3089,N_2970,N_2911);
nand U3090 (N_3090,N_2980,N_2999);
nor U3091 (N_3091,N_2977,N_2908);
nand U3092 (N_3092,N_2993,N_2906);
and U3093 (N_3093,N_2920,N_2954);
or U3094 (N_3094,N_2931,N_2934);
xnor U3095 (N_3095,N_2964,N_2999);
xnor U3096 (N_3096,N_2998,N_2957);
and U3097 (N_3097,N_2934,N_2951);
and U3098 (N_3098,N_2993,N_2926);
xor U3099 (N_3099,N_2936,N_2951);
nand U3100 (N_3100,N_3069,N_3013);
xnor U3101 (N_3101,N_3031,N_3059);
nand U3102 (N_3102,N_3004,N_3075);
xnor U3103 (N_3103,N_3006,N_3020);
nor U3104 (N_3104,N_3012,N_3081);
xor U3105 (N_3105,N_3024,N_3052);
nor U3106 (N_3106,N_3021,N_3068);
nor U3107 (N_3107,N_3089,N_3077);
nand U3108 (N_3108,N_3027,N_3061);
or U3109 (N_3109,N_3040,N_3057);
nor U3110 (N_3110,N_3017,N_3063);
and U3111 (N_3111,N_3084,N_3051);
nand U3112 (N_3112,N_3030,N_3009);
or U3113 (N_3113,N_3073,N_3053);
xor U3114 (N_3114,N_3048,N_3007);
xor U3115 (N_3115,N_3092,N_3085);
and U3116 (N_3116,N_3083,N_3082);
and U3117 (N_3117,N_3072,N_3045);
xor U3118 (N_3118,N_3026,N_3039);
and U3119 (N_3119,N_3042,N_3003);
or U3120 (N_3120,N_3023,N_3094);
nor U3121 (N_3121,N_3091,N_3014);
nand U3122 (N_3122,N_3034,N_3001);
xnor U3123 (N_3123,N_3038,N_3055);
and U3124 (N_3124,N_3071,N_3022);
xor U3125 (N_3125,N_3065,N_3025);
xor U3126 (N_3126,N_3043,N_3044);
nand U3127 (N_3127,N_3010,N_3016);
nor U3128 (N_3128,N_3000,N_3032);
nor U3129 (N_3129,N_3097,N_3090);
and U3130 (N_3130,N_3033,N_3066);
xor U3131 (N_3131,N_3058,N_3049);
nor U3132 (N_3132,N_3060,N_3098);
nor U3133 (N_3133,N_3064,N_3087);
and U3134 (N_3134,N_3056,N_3093);
nand U3135 (N_3135,N_3079,N_3037);
xor U3136 (N_3136,N_3008,N_3076);
xor U3137 (N_3137,N_3005,N_3054);
nand U3138 (N_3138,N_3019,N_3080);
and U3139 (N_3139,N_3011,N_3074);
nor U3140 (N_3140,N_3028,N_3088);
nand U3141 (N_3141,N_3041,N_3035);
nand U3142 (N_3142,N_3029,N_3002);
and U3143 (N_3143,N_3062,N_3078);
or U3144 (N_3144,N_3046,N_3015);
nor U3145 (N_3145,N_3086,N_3099);
xor U3146 (N_3146,N_3067,N_3096);
nand U3147 (N_3147,N_3047,N_3095);
nor U3148 (N_3148,N_3050,N_3036);
or U3149 (N_3149,N_3070,N_3018);
or U3150 (N_3150,N_3098,N_3028);
xnor U3151 (N_3151,N_3001,N_3011);
xor U3152 (N_3152,N_3096,N_3047);
and U3153 (N_3153,N_3082,N_3086);
or U3154 (N_3154,N_3068,N_3078);
xnor U3155 (N_3155,N_3047,N_3053);
nand U3156 (N_3156,N_3070,N_3060);
and U3157 (N_3157,N_3051,N_3044);
nand U3158 (N_3158,N_3052,N_3038);
and U3159 (N_3159,N_3091,N_3074);
or U3160 (N_3160,N_3068,N_3081);
and U3161 (N_3161,N_3075,N_3025);
and U3162 (N_3162,N_3034,N_3083);
xnor U3163 (N_3163,N_3063,N_3053);
nand U3164 (N_3164,N_3035,N_3095);
or U3165 (N_3165,N_3050,N_3071);
nand U3166 (N_3166,N_3007,N_3059);
and U3167 (N_3167,N_3059,N_3050);
or U3168 (N_3168,N_3082,N_3044);
nor U3169 (N_3169,N_3097,N_3051);
and U3170 (N_3170,N_3034,N_3066);
xnor U3171 (N_3171,N_3017,N_3081);
or U3172 (N_3172,N_3085,N_3047);
nand U3173 (N_3173,N_3041,N_3083);
nand U3174 (N_3174,N_3060,N_3048);
or U3175 (N_3175,N_3045,N_3023);
or U3176 (N_3176,N_3036,N_3073);
nand U3177 (N_3177,N_3005,N_3043);
nor U3178 (N_3178,N_3024,N_3028);
nor U3179 (N_3179,N_3054,N_3034);
nor U3180 (N_3180,N_3005,N_3060);
nand U3181 (N_3181,N_3067,N_3033);
nand U3182 (N_3182,N_3003,N_3038);
nand U3183 (N_3183,N_3092,N_3069);
and U3184 (N_3184,N_3070,N_3085);
or U3185 (N_3185,N_3051,N_3080);
and U3186 (N_3186,N_3028,N_3006);
nand U3187 (N_3187,N_3096,N_3001);
xnor U3188 (N_3188,N_3034,N_3051);
and U3189 (N_3189,N_3021,N_3074);
or U3190 (N_3190,N_3028,N_3081);
nand U3191 (N_3191,N_3011,N_3070);
or U3192 (N_3192,N_3067,N_3079);
or U3193 (N_3193,N_3062,N_3025);
xor U3194 (N_3194,N_3032,N_3025);
and U3195 (N_3195,N_3090,N_3043);
and U3196 (N_3196,N_3067,N_3003);
and U3197 (N_3197,N_3013,N_3006);
nor U3198 (N_3198,N_3060,N_3045);
and U3199 (N_3199,N_3052,N_3045);
and U3200 (N_3200,N_3192,N_3182);
xnor U3201 (N_3201,N_3137,N_3184);
nor U3202 (N_3202,N_3166,N_3138);
and U3203 (N_3203,N_3171,N_3126);
or U3204 (N_3204,N_3157,N_3136);
nor U3205 (N_3205,N_3140,N_3156);
and U3206 (N_3206,N_3180,N_3188);
nor U3207 (N_3207,N_3141,N_3119);
xor U3208 (N_3208,N_3111,N_3146);
and U3209 (N_3209,N_3128,N_3115);
nor U3210 (N_3210,N_3186,N_3101);
xor U3211 (N_3211,N_3187,N_3104);
nor U3212 (N_3212,N_3160,N_3132);
and U3213 (N_3213,N_3143,N_3190);
xnor U3214 (N_3214,N_3118,N_3189);
nor U3215 (N_3215,N_3183,N_3103);
nor U3216 (N_3216,N_3169,N_3114);
or U3217 (N_3217,N_3127,N_3170);
and U3218 (N_3218,N_3196,N_3122);
and U3219 (N_3219,N_3154,N_3155);
nand U3220 (N_3220,N_3113,N_3194);
nor U3221 (N_3221,N_3130,N_3106);
or U3222 (N_3222,N_3147,N_3150);
and U3223 (N_3223,N_3159,N_3198);
xor U3224 (N_3224,N_3109,N_3123);
and U3225 (N_3225,N_3125,N_3185);
nor U3226 (N_3226,N_3135,N_3149);
and U3227 (N_3227,N_3151,N_3131);
xor U3228 (N_3228,N_3108,N_3139);
xnor U3229 (N_3229,N_3176,N_3134);
nand U3230 (N_3230,N_3177,N_3178);
nand U3231 (N_3231,N_3102,N_3129);
or U3232 (N_3232,N_3153,N_3173);
or U3233 (N_3233,N_3164,N_3144);
nand U3234 (N_3234,N_3116,N_3167);
nor U3235 (N_3235,N_3162,N_3191);
or U3236 (N_3236,N_3181,N_3120);
nand U3237 (N_3237,N_3121,N_3174);
nand U3238 (N_3238,N_3110,N_3195);
xnor U3239 (N_3239,N_3133,N_3168);
and U3240 (N_3240,N_3165,N_3172);
or U3241 (N_3241,N_3107,N_3142);
nor U3242 (N_3242,N_3163,N_3161);
nand U3243 (N_3243,N_3145,N_3179);
xnor U3244 (N_3244,N_3152,N_3158);
or U3245 (N_3245,N_3105,N_3100);
or U3246 (N_3246,N_3112,N_3117);
nor U3247 (N_3247,N_3193,N_3148);
nand U3248 (N_3248,N_3124,N_3175);
nand U3249 (N_3249,N_3197,N_3199);
xnor U3250 (N_3250,N_3139,N_3120);
or U3251 (N_3251,N_3163,N_3116);
xor U3252 (N_3252,N_3166,N_3148);
and U3253 (N_3253,N_3106,N_3139);
and U3254 (N_3254,N_3166,N_3134);
nand U3255 (N_3255,N_3108,N_3186);
nand U3256 (N_3256,N_3128,N_3114);
nor U3257 (N_3257,N_3168,N_3196);
and U3258 (N_3258,N_3148,N_3128);
xor U3259 (N_3259,N_3143,N_3142);
xor U3260 (N_3260,N_3129,N_3124);
or U3261 (N_3261,N_3149,N_3166);
and U3262 (N_3262,N_3191,N_3110);
nand U3263 (N_3263,N_3191,N_3125);
nand U3264 (N_3264,N_3177,N_3135);
xor U3265 (N_3265,N_3158,N_3110);
xor U3266 (N_3266,N_3120,N_3171);
or U3267 (N_3267,N_3182,N_3119);
xnor U3268 (N_3268,N_3122,N_3121);
nor U3269 (N_3269,N_3174,N_3127);
xnor U3270 (N_3270,N_3196,N_3185);
nand U3271 (N_3271,N_3103,N_3173);
and U3272 (N_3272,N_3148,N_3154);
nor U3273 (N_3273,N_3183,N_3116);
nor U3274 (N_3274,N_3111,N_3154);
xor U3275 (N_3275,N_3125,N_3113);
nand U3276 (N_3276,N_3197,N_3123);
xnor U3277 (N_3277,N_3106,N_3152);
nand U3278 (N_3278,N_3140,N_3130);
xor U3279 (N_3279,N_3166,N_3136);
or U3280 (N_3280,N_3197,N_3134);
xor U3281 (N_3281,N_3119,N_3156);
or U3282 (N_3282,N_3160,N_3167);
xor U3283 (N_3283,N_3198,N_3132);
or U3284 (N_3284,N_3111,N_3130);
nor U3285 (N_3285,N_3131,N_3107);
and U3286 (N_3286,N_3157,N_3146);
nor U3287 (N_3287,N_3161,N_3189);
nor U3288 (N_3288,N_3154,N_3133);
xor U3289 (N_3289,N_3101,N_3173);
nor U3290 (N_3290,N_3139,N_3156);
and U3291 (N_3291,N_3188,N_3181);
xor U3292 (N_3292,N_3148,N_3169);
nor U3293 (N_3293,N_3135,N_3166);
xnor U3294 (N_3294,N_3137,N_3176);
or U3295 (N_3295,N_3151,N_3176);
xor U3296 (N_3296,N_3179,N_3133);
and U3297 (N_3297,N_3141,N_3193);
and U3298 (N_3298,N_3179,N_3184);
xnor U3299 (N_3299,N_3170,N_3182);
nor U3300 (N_3300,N_3237,N_3287);
xor U3301 (N_3301,N_3214,N_3261);
nor U3302 (N_3302,N_3294,N_3216);
xnor U3303 (N_3303,N_3242,N_3297);
nand U3304 (N_3304,N_3263,N_3262);
nand U3305 (N_3305,N_3243,N_3212);
nor U3306 (N_3306,N_3202,N_3293);
nor U3307 (N_3307,N_3267,N_3217);
xor U3308 (N_3308,N_3296,N_3285);
xnor U3309 (N_3309,N_3247,N_3288);
or U3310 (N_3310,N_3249,N_3256);
or U3311 (N_3311,N_3221,N_3281);
xnor U3312 (N_3312,N_3225,N_3265);
xor U3313 (N_3313,N_3222,N_3269);
nand U3314 (N_3314,N_3250,N_3205);
nor U3315 (N_3315,N_3259,N_3207);
xnor U3316 (N_3316,N_3226,N_3224);
xnor U3317 (N_3317,N_3213,N_3264);
nor U3318 (N_3318,N_3273,N_3280);
nand U3319 (N_3319,N_3291,N_3209);
and U3320 (N_3320,N_3268,N_3282);
xor U3321 (N_3321,N_3274,N_3206);
nand U3322 (N_3322,N_3277,N_3246);
nand U3323 (N_3323,N_3292,N_3276);
xnor U3324 (N_3324,N_3231,N_3234);
xnor U3325 (N_3325,N_3215,N_3283);
nor U3326 (N_3326,N_3245,N_3255);
xor U3327 (N_3327,N_3232,N_3229);
xnor U3328 (N_3328,N_3244,N_3275);
nand U3329 (N_3329,N_3295,N_3236);
xor U3330 (N_3330,N_3235,N_3211);
nor U3331 (N_3331,N_3272,N_3270);
and U3332 (N_3332,N_3223,N_3258);
xnor U3333 (N_3333,N_3278,N_3290);
or U3334 (N_3334,N_3254,N_3218);
nor U3335 (N_3335,N_3253,N_3220);
nor U3336 (N_3336,N_3299,N_3279);
nand U3337 (N_3337,N_3289,N_3238);
nor U3338 (N_3338,N_3228,N_3271);
nand U3339 (N_3339,N_3257,N_3204);
nor U3340 (N_3340,N_3266,N_3298);
xor U3341 (N_3341,N_3201,N_3233);
nor U3342 (N_3342,N_3248,N_3260);
xor U3343 (N_3343,N_3240,N_3252);
xor U3344 (N_3344,N_3203,N_3284);
or U3345 (N_3345,N_3227,N_3239);
nand U3346 (N_3346,N_3200,N_3219);
nor U3347 (N_3347,N_3230,N_3208);
nor U3348 (N_3348,N_3251,N_3210);
xnor U3349 (N_3349,N_3286,N_3241);
xor U3350 (N_3350,N_3251,N_3219);
and U3351 (N_3351,N_3231,N_3293);
nor U3352 (N_3352,N_3271,N_3277);
xnor U3353 (N_3353,N_3266,N_3250);
xnor U3354 (N_3354,N_3213,N_3221);
xor U3355 (N_3355,N_3201,N_3276);
nand U3356 (N_3356,N_3233,N_3295);
or U3357 (N_3357,N_3210,N_3232);
or U3358 (N_3358,N_3255,N_3251);
or U3359 (N_3359,N_3253,N_3283);
xnor U3360 (N_3360,N_3237,N_3254);
and U3361 (N_3361,N_3265,N_3291);
or U3362 (N_3362,N_3238,N_3210);
and U3363 (N_3363,N_3235,N_3207);
nor U3364 (N_3364,N_3286,N_3271);
nand U3365 (N_3365,N_3221,N_3283);
xnor U3366 (N_3366,N_3210,N_3296);
nor U3367 (N_3367,N_3226,N_3204);
nand U3368 (N_3368,N_3282,N_3257);
and U3369 (N_3369,N_3237,N_3247);
and U3370 (N_3370,N_3268,N_3297);
and U3371 (N_3371,N_3282,N_3285);
nor U3372 (N_3372,N_3268,N_3276);
xor U3373 (N_3373,N_3222,N_3276);
nor U3374 (N_3374,N_3262,N_3208);
nand U3375 (N_3375,N_3211,N_3291);
xor U3376 (N_3376,N_3246,N_3233);
or U3377 (N_3377,N_3284,N_3280);
or U3378 (N_3378,N_3222,N_3246);
or U3379 (N_3379,N_3281,N_3212);
nor U3380 (N_3380,N_3266,N_3226);
nand U3381 (N_3381,N_3219,N_3298);
nor U3382 (N_3382,N_3280,N_3203);
or U3383 (N_3383,N_3269,N_3209);
nor U3384 (N_3384,N_3258,N_3253);
or U3385 (N_3385,N_3265,N_3224);
nand U3386 (N_3386,N_3252,N_3294);
or U3387 (N_3387,N_3275,N_3267);
nand U3388 (N_3388,N_3251,N_3274);
or U3389 (N_3389,N_3254,N_3248);
and U3390 (N_3390,N_3257,N_3201);
xor U3391 (N_3391,N_3203,N_3221);
nand U3392 (N_3392,N_3235,N_3299);
xor U3393 (N_3393,N_3222,N_3245);
nand U3394 (N_3394,N_3226,N_3203);
xor U3395 (N_3395,N_3278,N_3228);
and U3396 (N_3396,N_3268,N_3208);
nor U3397 (N_3397,N_3289,N_3246);
nand U3398 (N_3398,N_3272,N_3283);
xor U3399 (N_3399,N_3227,N_3249);
nor U3400 (N_3400,N_3315,N_3387);
nand U3401 (N_3401,N_3352,N_3357);
or U3402 (N_3402,N_3308,N_3375);
or U3403 (N_3403,N_3351,N_3322);
or U3404 (N_3404,N_3377,N_3341);
xor U3405 (N_3405,N_3390,N_3355);
xor U3406 (N_3406,N_3339,N_3321);
nor U3407 (N_3407,N_3381,N_3396);
xor U3408 (N_3408,N_3394,N_3371);
xnor U3409 (N_3409,N_3342,N_3338);
or U3410 (N_3410,N_3316,N_3327);
and U3411 (N_3411,N_3376,N_3320);
or U3412 (N_3412,N_3325,N_3319);
or U3413 (N_3413,N_3361,N_3368);
xor U3414 (N_3414,N_3305,N_3388);
nand U3415 (N_3415,N_3374,N_3380);
nand U3416 (N_3416,N_3310,N_3335);
nand U3417 (N_3417,N_3306,N_3329);
or U3418 (N_3418,N_3349,N_3372);
and U3419 (N_3419,N_3370,N_3331);
nor U3420 (N_3420,N_3345,N_3399);
and U3421 (N_3421,N_3328,N_3397);
xor U3422 (N_3422,N_3389,N_3369);
xor U3423 (N_3423,N_3363,N_3340);
or U3424 (N_3424,N_3364,N_3354);
or U3425 (N_3425,N_3343,N_3353);
nand U3426 (N_3426,N_3303,N_3382);
xor U3427 (N_3427,N_3356,N_3350);
and U3428 (N_3428,N_3366,N_3337);
xor U3429 (N_3429,N_3398,N_3348);
nor U3430 (N_3430,N_3314,N_3367);
or U3431 (N_3431,N_3307,N_3323);
xnor U3432 (N_3432,N_3334,N_3362);
nand U3433 (N_3433,N_3365,N_3378);
nand U3434 (N_3434,N_3309,N_3373);
nor U3435 (N_3435,N_3330,N_3391);
or U3436 (N_3436,N_3379,N_3385);
or U3437 (N_3437,N_3317,N_3301);
or U3438 (N_3438,N_3318,N_3336);
or U3439 (N_3439,N_3384,N_3312);
nor U3440 (N_3440,N_3313,N_3383);
or U3441 (N_3441,N_3360,N_3300);
and U3442 (N_3442,N_3311,N_3393);
nand U3443 (N_3443,N_3324,N_3359);
nor U3444 (N_3444,N_3333,N_3358);
xnor U3445 (N_3445,N_3332,N_3344);
or U3446 (N_3446,N_3392,N_3302);
nor U3447 (N_3447,N_3347,N_3346);
or U3448 (N_3448,N_3326,N_3395);
or U3449 (N_3449,N_3386,N_3304);
nand U3450 (N_3450,N_3390,N_3337);
nor U3451 (N_3451,N_3336,N_3302);
xor U3452 (N_3452,N_3327,N_3351);
nand U3453 (N_3453,N_3349,N_3313);
nor U3454 (N_3454,N_3326,N_3311);
and U3455 (N_3455,N_3388,N_3397);
and U3456 (N_3456,N_3378,N_3300);
or U3457 (N_3457,N_3367,N_3393);
xnor U3458 (N_3458,N_3304,N_3317);
nor U3459 (N_3459,N_3353,N_3316);
xor U3460 (N_3460,N_3317,N_3369);
or U3461 (N_3461,N_3328,N_3368);
or U3462 (N_3462,N_3394,N_3365);
and U3463 (N_3463,N_3397,N_3391);
and U3464 (N_3464,N_3302,N_3395);
and U3465 (N_3465,N_3345,N_3367);
nand U3466 (N_3466,N_3393,N_3378);
nor U3467 (N_3467,N_3355,N_3358);
or U3468 (N_3468,N_3353,N_3304);
or U3469 (N_3469,N_3358,N_3390);
nor U3470 (N_3470,N_3384,N_3310);
xnor U3471 (N_3471,N_3375,N_3312);
nand U3472 (N_3472,N_3333,N_3334);
xnor U3473 (N_3473,N_3324,N_3372);
nor U3474 (N_3474,N_3343,N_3320);
and U3475 (N_3475,N_3361,N_3327);
or U3476 (N_3476,N_3319,N_3367);
xor U3477 (N_3477,N_3357,N_3343);
nand U3478 (N_3478,N_3313,N_3305);
xnor U3479 (N_3479,N_3393,N_3301);
xor U3480 (N_3480,N_3371,N_3363);
nor U3481 (N_3481,N_3392,N_3367);
and U3482 (N_3482,N_3392,N_3300);
nand U3483 (N_3483,N_3384,N_3338);
nand U3484 (N_3484,N_3378,N_3316);
nand U3485 (N_3485,N_3341,N_3333);
nand U3486 (N_3486,N_3313,N_3318);
and U3487 (N_3487,N_3398,N_3386);
nor U3488 (N_3488,N_3309,N_3319);
xor U3489 (N_3489,N_3306,N_3383);
nand U3490 (N_3490,N_3360,N_3395);
or U3491 (N_3491,N_3392,N_3342);
nand U3492 (N_3492,N_3309,N_3387);
nor U3493 (N_3493,N_3335,N_3387);
or U3494 (N_3494,N_3393,N_3375);
or U3495 (N_3495,N_3334,N_3318);
nor U3496 (N_3496,N_3304,N_3366);
nand U3497 (N_3497,N_3302,N_3378);
xnor U3498 (N_3498,N_3376,N_3307);
or U3499 (N_3499,N_3300,N_3342);
or U3500 (N_3500,N_3457,N_3460);
nor U3501 (N_3501,N_3476,N_3495);
nor U3502 (N_3502,N_3435,N_3430);
nand U3503 (N_3503,N_3409,N_3454);
and U3504 (N_3504,N_3446,N_3470);
or U3505 (N_3505,N_3425,N_3483);
nand U3506 (N_3506,N_3444,N_3485);
and U3507 (N_3507,N_3453,N_3471);
xor U3508 (N_3508,N_3486,N_3438);
and U3509 (N_3509,N_3431,N_3490);
and U3510 (N_3510,N_3449,N_3404);
or U3511 (N_3511,N_3488,N_3480);
and U3512 (N_3512,N_3473,N_3417);
xor U3513 (N_3513,N_3456,N_3419);
nand U3514 (N_3514,N_3434,N_3422);
xor U3515 (N_3515,N_3415,N_3478);
and U3516 (N_3516,N_3439,N_3464);
nor U3517 (N_3517,N_3463,N_3436);
nor U3518 (N_3518,N_3429,N_3465);
or U3519 (N_3519,N_3420,N_3493);
or U3520 (N_3520,N_3479,N_3400);
nand U3521 (N_3521,N_3452,N_3487);
and U3522 (N_3522,N_3402,N_3491);
or U3523 (N_3523,N_3401,N_3426);
xnor U3524 (N_3524,N_3461,N_3459);
nor U3525 (N_3525,N_3418,N_3462);
xor U3526 (N_3526,N_3428,N_3497);
or U3527 (N_3527,N_3472,N_3403);
nand U3528 (N_3528,N_3443,N_3416);
and U3529 (N_3529,N_3482,N_3477);
xor U3530 (N_3530,N_3437,N_3407);
nor U3531 (N_3531,N_3467,N_3408);
xnor U3532 (N_3532,N_3498,N_3412);
xor U3533 (N_3533,N_3423,N_3499);
nor U3534 (N_3534,N_3458,N_3448);
xor U3535 (N_3535,N_3455,N_3410);
xnor U3536 (N_3536,N_3447,N_3468);
or U3537 (N_3537,N_3474,N_3451);
and U3538 (N_3538,N_3445,N_3494);
or U3539 (N_3539,N_3414,N_3432);
xnor U3540 (N_3540,N_3440,N_3489);
xor U3541 (N_3541,N_3475,N_3466);
nand U3542 (N_3542,N_3433,N_3421);
xor U3543 (N_3543,N_3406,N_3492);
and U3544 (N_3544,N_3450,N_3442);
nor U3545 (N_3545,N_3413,N_3441);
xor U3546 (N_3546,N_3496,N_3481);
xor U3547 (N_3547,N_3405,N_3427);
nand U3548 (N_3548,N_3424,N_3411);
xnor U3549 (N_3549,N_3484,N_3469);
nand U3550 (N_3550,N_3430,N_3412);
or U3551 (N_3551,N_3475,N_3491);
and U3552 (N_3552,N_3421,N_3418);
and U3553 (N_3553,N_3458,N_3439);
or U3554 (N_3554,N_3450,N_3422);
nor U3555 (N_3555,N_3446,N_3412);
nand U3556 (N_3556,N_3485,N_3424);
and U3557 (N_3557,N_3418,N_3403);
xor U3558 (N_3558,N_3445,N_3449);
nand U3559 (N_3559,N_3460,N_3469);
xor U3560 (N_3560,N_3446,N_3411);
nand U3561 (N_3561,N_3423,N_3480);
nor U3562 (N_3562,N_3440,N_3405);
nor U3563 (N_3563,N_3438,N_3495);
nand U3564 (N_3564,N_3447,N_3454);
nand U3565 (N_3565,N_3406,N_3469);
nand U3566 (N_3566,N_3497,N_3445);
nand U3567 (N_3567,N_3473,N_3419);
nor U3568 (N_3568,N_3465,N_3408);
nand U3569 (N_3569,N_3440,N_3427);
nand U3570 (N_3570,N_3494,N_3437);
and U3571 (N_3571,N_3444,N_3464);
nand U3572 (N_3572,N_3464,N_3428);
xnor U3573 (N_3573,N_3439,N_3440);
xor U3574 (N_3574,N_3414,N_3495);
nand U3575 (N_3575,N_3438,N_3426);
or U3576 (N_3576,N_3439,N_3478);
or U3577 (N_3577,N_3441,N_3450);
xnor U3578 (N_3578,N_3496,N_3485);
or U3579 (N_3579,N_3443,N_3412);
nand U3580 (N_3580,N_3409,N_3440);
xnor U3581 (N_3581,N_3438,N_3409);
xnor U3582 (N_3582,N_3430,N_3495);
nand U3583 (N_3583,N_3434,N_3495);
or U3584 (N_3584,N_3406,N_3404);
xor U3585 (N_3585,N_3435,N_3409);
and U3586 (N_3586,N_3423,N_3425);
xor U3587 (N_3587,N_3451,N_3419);
nor U3588 (N_3588,N_3423,N_3400);
and U3589 (N_3589,N_3485,N_3497);
xor U3590 (N_3590,N_3490,N_3496);
or U3591 (N_3591,N_3467,N_3453);
and U3592 (N_3592,N_3480,N_3454);
xnor U3593 (N_3593,N_3415,N_3418);
nor U3594 (N_3594,N_3484,N_3473);
nor U3595 (N_3595,N_3412,N_3415);
or U3596 (N_3596,N_3468,N_3420);
and U3597 (N_3597,N_3442,N_3464);
and U3598 (N_3598,N_3410,N_3494);
and U3599 (N_3599,N_3440,N_3491);
nand U3600 (N_3600,N_3538,N_3599);
nor U3601 (N_3601,N_3584,N_3573);
and U3602 (N_3602,N_3564,N_3582);
nor U3603 (N_3603,N_3569,N_3567);
and U3604 (N_3604,N_3596,N_3513);
or U3605 (N_3605,N_3592,N_3525);
xor U3606 (N_3606,N_3536,N_3557);
nand U3607 (N_3607,N_3574,N_3549);
xnor U3608 (N_3608,N_3529,N_3591);
nand U3609 (N_3609,N_3581,N_3516);
or U3610 (N_3610,N_3590,N_3539);
nand U3611 (N_3611,N_3544,N_3527);
xor U3612 (N_3612,N_3506,N_3555);
nor U3613 (N_3613,N_3552,N_3585);
nand U3614 (N_3614,N_3563,N_3597);
and U3615 (N_3615,N_3534,N_3562);
and U3616 (N_3616,N_3508,N_3532);
nor U3617 (N_3617,N_3505,N_3509);
nor U3618 (N_3618,N_3512,N_3519);
xor U3619 (N_3619,N_3528,N_3551);
nor U3620 (N_3620,N_3500,N_3570);
nor U3621 (N_3621,N_3543,N_3514);
xnor U3622 (N_3622,N_3580,N_3504);
and U3623 (N_3623,N_3571,N_3542);
or U3624 (N_3624,N_3583,N_3541);
xor U3625 (N_3625,N_3598,N_3507);
xor U3626 (N_3626,N_3588,N_3537);
nor U3627 (N_3627,N_3548,N_3595);
or U3628 (N_3628,N_3550,N_3587);
or U3629 (N_3629,N_3530,N_3578);
or U3630 (N_3630,N_3502,N_3511);
and U3631 (N_3631,N_3560,N_3503);
and U3632 (N_3632,N_3510,N_3554);
nor U3633 (N_3633,N_3579,N_3566);
and U3634 (N_3634,N_3546,N_3593);
or U3635 (N_3635,N_3565,N_3577);
or U3636 (N_3636,N_3576,N_3545);
and U3637 (N_3637,N_3526,N_3524);
nor U3638 (N_3638,N_3522,N_3553);
and U3639 (N_3639,N_3594,N_3575);
nand U3640 (N_3640,N_3523,N_3556);
nor U3641 (N_3641,N_3586,N_3520);
xor U3642 (N_3642,N_3572,N_3515);
or U3643 (N_3643,N_3518,N_3568);
or U3644 (N_3644,N_3521,N_3531);
xor U3645 (N_3645,N_3559,N_3517);
or U3646 (N_3646,N_3547,N_3535);
xor U3647 (N_3647,N_3501,N_3561);
nand U3648 (N_3648,N_3558,N_3533);
or U3649 (N_3649,N_3589,N_3540);
nand U3650 (N_3650,N_3543,N_3565);
xor U3651 (N_3651,N_3522,N_3584);
nor U3652 (N_3652,N_3545,N_3524);
nor U3653 (N_3653,N_3523,N_3522);
and U3654 (N_3654,N_3593,N_3553);
xor U3655 (N_3655,N_3517,N_3591);
and U3656 (N_3656,N_3596,N_3550);
nand U3657 (N_3657,N_3523,N_3562);
nand U3658 (N_3658,N_3588,N_3539);
nand U3659 (N_3659,N_3594,N_3513);
nor U3660 (N_3660,N_3581,N_3520);
and U3661 (N_3661,N_3565,N_3516);
nand U3662 (N_3662,N_3530,N_3500);
nand U3663 (N_3663,N_3533,N_3536);
xor U3664 (N_3664,N_3533,N_3508);
xor U3665 (N_3665,N_3531,N_3583);
nand U3666 (N_3666,N_3568,N_3546);
and U3667 (N_3667,N_3587,N_3523);
nor U3668 (N_3668,N_3552,N_3528);
or U3669 (N_3669,N_3542,N_3515);
and U3670 (N_3670,N_3564,N_3514);
or U3671 (N_3671,N_3513,N_3593);
or U3672 (N_3672,N_3502,N_3586);
xnor U3673 (N_3673,N_3581,N_3592);
nor U3674 (N_3674,N_3568,N_3596);
nand U3675 (N_3675,N_3559,N_3555);
nor U3676 (N_3676,N_3556,N_3582);
xor U3677 (N_3677,N_3520,N_3555);
or U3678 (N_3678,N_3568,N_3515);
or U3679 (N_3679,N_3568,N_3583);
and U3680 (N_3680,N_3598,N_3506);
xnor U3681 (N_3681,N_3588,N_3529);
or U3682 (N_3682,N_3500,N_3585);
nor U3683 (N_3683,N_3542,N_3547);
or U3684 (N_3684,N_3560,N_3587);
and U3685 (N_3685,N_3516,N_3540);
or U3686 (N_3686,N_3588,N_3570);
xnor U3687 (N_3687,N_3593,N_3575);
xor U3688 (N_3688,N_3570,N_3553);
nor U3689 (N_3689,N_3574,N_3585);
nor U3690 (N_3690,N_3560,N_3508);
and U3691 (N_3691,N_3554,N_3581);
xor U3692 (N_3692,N_3545,N_3591);
or U3693 (N_3693,N_3521,N_3548);
or U3694 (N_3694,N_3589,N_3529);
and U3695 (N_3695,N_3535,N_3553);
nand U3696 (N_3696,N_3550,N_3593);
nand U3697 (N_3697,N_3579,N_3557);
nor U3698 (N_3698,N_3535,N_3551);
and U3699 (N_3699,N_3514,N_3594);
nand U3700 (N_3700,N_3682,N_3625);
and U3701 (N_3701,N_3671,N_3628);
or U3702 (N_3702,N_3640,N_3618);
nor U3703 (N_3703,N_3624,N_3637);
xor U3704 (N_3704,N_3600,N_3663);
nor U3705 (N_3705,N_3673,N_3680);
xor U3706 (N_3706,N_3643,N_3614);
xnor U3707 (N_3707,N_3642,N_3659);
nand U3708 (N_3708,N_3690,N_3626);
nor U3709 (N_3709,N_3620,N_3647);
and U3710 (N_3710,N_3653,N_3603);
or U3711 (N_3711,N_3660,N_3612);
xor U3712 (N_3712,N_3662,N_3652);
and U3713 (N_3713,N_3692,N_3687);
and U3714 (N_3714,N_3609,N_3633);
nand U3715 (N_3715,N_3613,N_3617);
or U3716 (N_3716,N_3666,N_3641);
or U3717 (N_3717,N_3693,N_3650);
and U3718 (N_3718,N_3689,N_3648);
nand U3719 (N_3719,N_3622,N_3669);
xnor U3720 (N_3720,N_3675,N_3646);
and U3721 (N_3721,N_3639,N_3661);
xnor U3722 (N_3722,N_3679,N_3615);
nand U3723 (N_3723,N_3676,N_3636);
xnor U3724 (N_3724,N_3657,N_3605);
xnor U3725 (N_3725,N_3645,N_3616);
and U3726 (N_3726,N_3697,N_3698);
nand U3727 (N_3727,N_3694,N_3601);
and U3728 (N_3728,N_3658,N_3607);
xor U3729 (N_3729,N_3649,N_3634);
and U3730 (N_3730,N_3677,N_3670);
nor U3731 (N_3731,N_3629,N_3638);
nand U3732 (N_3732,N_3683,N_3611);
or U3733 (N_3733,N_3656,N_3668);
or U3734 (N_3734,N_3674,N_3699);
and U3735 (N_3735,N_3602,N_3696);
nand U3736 (N_3736,N_3684,N_3621);
nand U3737 (N_3737,N_3608,N_3681);
or U3738 (N_3738,N_3655,N_3667);
and U3739 (N_3739,N_3631,N_3627);
nand U3740 (N_3740,N_3678,N_3665);
and U3741 (N_3741,N_3623,N_3606);
or U3742 (N_3742,N_3619,N_3610);
nor U3743 (N_3743,N_3654,N_3688);
xnor U3744 (N_3744,N_3632,N_3630);
xor U3745 (N_3745,N_3691,N_3635);
and U3746 (N_3746,N_3664,N_3686);
nor U3747 (N_3747,N_3672,N_3695);
and U3748 (N_3748,N_3685,N_3604);
nor U3749 (N_3749,N_3651,N_3644);
xor U3750 (N_3750,N_3674,N_3637);
xor U3751 (N_3751,N_3685,N_3616);
nand U3752 (N_3752,N_3678,N_3629);
nand U3753 (N_3753,N_3627,N_3623);
or U3754 (N_3754,N_3667,N_3625);
nand U3755 (N_3755,N_3626,N_3660);
and U3756 (N_3756,N_3689,N_3645);
or U3757 (N_3757,N_3695,N_3601);
xnor U3758 (N_3758,N_3638,N_3605);
or U3759 (N_3759,N_3639,N_3627);
xor U3760 (N_3760,N_3640,N_3644);
or U3761 (N_3761,N_3640,N_3672);
and U3762 (N_3762,N_3614,N_3662);
xnor U3763 (N_3763,N_3668,N_3655);
or U3764 (N_3764,N_3634,N_3624);
xor U3765 (N_3765,N_3672,N_3699);
and U3766 (N_3766,N_3675,N_3637);
xor U3767 (N_3767,N_3618,N_3685);
or U3768 (N_3768,N_3658,N_3696);
and U3769 (N_3769,N_3672,N_3696);
nor U3770 (N_3770,N_3628,N_3630);
nand U3771 (N_3771,N_3694,N_3622);
or U3772 (N_3772,N_3616,N_3641);
nand U3773 (N_3773,N_3668,N_3664);
nand U3774 (N_3774,N_3663,N_3641);
nor U3775 (N_3775,N_3667,N_3648);
nand U3776 (N_3776,N_3659,N_3681);
nor U3777 (N_3777,N_3664,N_3639);
or U3778 (N_3778,N_3670,N_3618);
or U3779 (N_3779,N_3625,N_3653);
nor U3780 (N_3780,N_3669,N_3604);
nand U3781 (N_3781,N_3663,N_3672);
nor U3782 (N_3782,N_3612,N_3668);
nand U3783 (N_3783,N_3673,N_3642);
nor U3784 (N_3784,N_3653,N_3615);
nor U3785 (N_3785,N_3627,N_3681);
and U3786 (N_3786,N_3688,N_3646);
nand U3787 (N_3787,N_3674,N_3684);
and U3788 (N_3788,N_3681,N_3657);
or U3789 (N_3789,N_3603,N_3649);
or U3790 (N_3790,N_3650,N_3627);
nor U3791 (N_3791,N_3671,N_3634);
or U3792 (N_3792,N_3678,N_3675);
or U3793 (N_3793,N_3690,N_3688);
nand U3794 (N_3794,N_3618,N_3696);
xnor U3795 (N_3795,N_3606,N_3672);
nor U3796 (N_3796,N_3695,N_3687);
and U3797 (N_3797,N_3649,N_3680);
nor U3798 (N_3798,N_3618,N_3686);
and U3799 (N_3799,N_3602,N_3657);
nor U3800 (N_3800,N_3722,N_3764);
xnor U3801 (N_3801,N_3761,N_3787);
or U3802 (N_3802,N_3745,N_3721);
or U3803 (N_3803,N_3748,N_3790);
xor U3804 (N_3804,N_3735,N_3799);
xnor U3805 (N_3805,N_3734,N_3792);
or U3806 (N_3806,N_3771,N_3736);
and U3807 (N_3807,N_3783,N_3767);
xnor U3808 (N_3808,N_3757,N_3714);
nand U3809 (N_3809,N_3754,N_3760);
nor U3810 (N_3810,N_3747,N_3766);
and U3811 (N_3811,N_3763,N_3780);
nand U3812 (N_3812,N_3795,N_3788);
or U3813 (N_3813,N_3708,N_3753);
nand U3814 (N_3814,N_3728,N_3774);
xor U3815 (N_3815,N_3785,N_3789);
nor U3816 (N_3816,N_3713,N_3777);
and U3817 (N_3817,N_3719,N_3733);
xor U3818 (N_3818,N_3773,N_3756);
xor U3819 (N_3819,N_3707,N_3731);
nand U3820 (N_3820,N_3749,N_3779);
xor U3821 (N_3821,N_3700,N_3702);
nor U3822 (N_3822,N_3770,N_3703);
xor U3823 (N_3823,N_3751,N_3744);
xor U3824 (N_3824,N_3704,N_3781);
xnor U3825 (N_3825,N_3759,N_3726);
nor U3826 (N_3826,N_3720,N_3794);
or U3827 (N_3827,N_3762,N_3709);
nand U3828 (N_3828,N_3725,N_3715);
nor U3829 (N_3829,N_3778,N_3739);
xnor U3830 (N_3830,N_3797,N_3758);
xor U3831 (N_3831,N_3717,N_3798);
nor U3832 (N_3832,N_3730,N_3738);
and U3833 (N_3833,N_3750,N_3723);
xor U3834 (N_3834,N_3712,N_3782);
nor U3835 (N_3835,N_3769,N_3765);
nand U3836 (N_3836,N_3791,N_3752);
nand U3837 (N_3837,N_3742,N_3716);
nand U3838 (N_3838,N_3701,N_3768);
nand U3839 (N_3839,N_3776,N_3746);
nor U3840 (N_3840,N_3718,N_3784);
nor U3841 (N_3841,N_3743,N_3793);
nor U3842 (N_3842,N_3706,N_3705);
nand U3843 (N_3843,N_3755,N_3740);
or U3844 (N_3844,N_3732,N_3796);
or U3845 (N_3845,N_3786,N_3727);
and U3846 (N_3846,N_3772,N_3737);
xnor U3847 (N_3847,N_3724,N_3710);
nand U3848 (N_3848,N_3711,N_3729);
nor U3849 (N_3849,N_3775,N_3741);
and U3850 (N_3850,N_3744,N_3736);
nand U3851 (N_3851,N_3756,N_3738);
nor U3852 (N_3852,N_3753,N_3704);
nor U3853 (N_3853,N_3731,N_3762);
nand U3854 (N_3854,N_3792,N_3726);
and U3855 (N_3855,N_3790,N_3789);
or U3856 (N_3856,N_3738,N_3715);
and U3857 (N_3857,N_3799,N_3755);
xor U3858 (N_3858,N_3737,N_3773);
or U3859 (N_3859,N_3714,N_3772);
xnor U3860 (N_3860,N_3782,N_3783);
or U3861 (N_3861,N_3746,N_3774);
nor U3862 (N_3862,N_3756,N_3743);
nand U3863 (N_3863,N_3780,N_3743);
and U3864 (N_3864,N_3755,N_3789);
or U3865 (N_3865,N_3721,N_3716);
xnor U3866 (N_3866,N_3733,N_3722);
and U3867 (N_3867,N_3764,N_3731);
and U3868 (N_3868,N_3765,N_3781);
xor U3869 (N_3869,N_3751,N_3745);
and U3870 (N_3870,N_3780,N_3744);
and U3871 (N_3871,N_3758,N_3771);
or U3872 (N_3872,N_3777,N_3705);
nor U3873 (N_3873,N_3797,N_3784);
nand U3874 (N_3874,N_3799,N_3743);
or U3875 (N_3875,N_3775,N_3759);
nand U3876 (N_3876,N_3738,N_3788);
or U3877 (N_3877,N_3746,N_3736);
and U3878 (N_3878,N_3749,N_3773);
and U3879 (N_3879,N_3751,N_3732);
xor U3880 (N_3880,N_3790,N_3778);
and U3881 (N_3881,N_3708,N_3774);
nand U3882 (N_3882,N_3762,N_3767);
nor U3883 (N_3883,N_3798,N_3719);
and U3884 (N_3884,N_3730,N_3760);
and U3885 (N_3885,N_3773,N_3706);
and U3886 (N_3886,N_3741,N_3736);
nand U3887 (N_3887,N_3750,N_3727);
nor U3888 (N_3888,N_3720,N_3746);
xnor U3889 (N_3889,N_3776,N_3757);
and U3890 (N_3890,N_3729,N_3791);
nor U3891 (N_3891,N_3741,N_3733);
or U3892 (N_3892,N_3753,N_3729);
xor U3893 (N_3893,N_3735,N_3719);
xor U3894 (N_3894,N_3730,N_3773);
xnor U3895 (N_3895,N_3766,N_3780);
and U3896 (N_3896,N_3770,N_3789);
xor U3897 (N_3897,N_3777,N_3755);
nand U3898 (N_3898,N_3755,N_3788);
nor U3899 (N_3899,N_3716,N_3771);
nand U3900 (N_3900,N_3899,N_3892);
nand U3901 (N_3901,N_3820,N_3816);
xnor U3902 (N_3902,N_3812,N_3876);
and U3903 (N_3903,N_3890,N_3839);
xor U3904 (N_3904,N_3888,N_3875);
xor U3905 (N_3905,N_3869,N_3857);
nand U3906 (N_3906,N_3872,N_3814);
and U3907 (N_3907,N_3884,N_3877);
and U3908 (N_3908,N_3878,N_3826);
and U3909 (N_3909,N_3880,N_3840);
and U3910 (N_3910,N_3803,N_3870);
nor U3911 (N_3911,N_3838,N_3883);
or U3912 (N_3912,N_3868,N_3879);
and U3913 (N_3913,N_3859,N_3801);
nor U3914 (N_3914,N_3889,N_3846);
or U3915 (N_3915,N_3860,N_3853);
nor U3916 (N_3916,N_3864,N_3849);
xnor U3917 (N_3917,N_3821,N_3873);
and U3918 (N_3918,N_3866,N_3871);
or U3919 (N_3919,N_3828,N_3894);
or U3920 (N_3920,N_3896,N_3844);
and U3921 (N_3921,N_3893,N_3855);
or U3922 (N_3922,N_3835,N_3810);
nor U3923 (N_3923,N_3848,N_3837);
and U3924 (N_3924,N_3819,N_3809);
xor U3925 (N_3925,N_3852,N_3858);
nor U3926 (N_3926,N_3845,N_3836);
xnor U3927 (N_3927,N_3811,N_3834);
nand U3928 (N_3928,N_3824,N_3813);
xnor U3929 (N_3929,N_3887,N_3818);
or U3930 (N_3930,N_3867,N_3808);
or U3931 (N_3931,N_3815,N_3850);
nor U3932 (N_3932,N_3805,N_3847);
or U3933 (N_3933,N_3863,N_3862);
or U3934 (N_3934,N_3802,N_3895);
nor U3935 (N_3935,N_3856,N_3817);
nor U3936 (N_3936,N_3822,N_3800);
or U3937 (N_3937,N_3885,N_3806);
and U3938 (N_3938,N_3881,N_3842);
nand U3939 (N_3939,N_3854,N_3874);
xnor U3940 (N_3940,N_3829,N_3807);
or U3941 (N_3941,N_3865,N_3886);
or U3942 (N_3942,N_3841,N_3827);
nand U3943 (N_3943,N_3825,N_3898);
or U3944 (N_3944,N_3897,N_3843);
nand U3945 (N_3945,N_3833,N_3830);
or U3946 (N_3946,N_3804,N_3823);
or U3947 (N_3947,N_3851,N_3831);
xnor U3948 (N_3948,N_3832,N_3882);
and U3949 (N_3949,N_3861,N_3891);
nand U3950 (N_3950,N_3844,N_3882);
nor U3951 (N_3951,N_3878,N_3825);
or U3952 (N_3952,N_3896,N_3856);
or U3953 (N_3953,N_3869,N_3875);
nand U3954 (N_3954,N_3832,N_3814);
xnor U3955 (N_3955,N_3812,N_3807);
nand U3956 (N_3956,N_3880,N_3831);
xor U3957 (N_3957,N_3810,N_3862);
and U3958 (N_3958,N_3839,N_3802);
nor U3959 (N_3959,N_3803,N_3846);
and U3960 (N_3960,N_3815,N_3813);
and U3961 (N_3961,N_3866,N_3818);
nand U3962 (N_3962,N_3866,N_3826);
nor U3963 (N_3963,N_3876,N_3832);
nor U3964 (N_3964,N_3892,N_3870);
or U3965 (N_3965,N_3890,N_3815);
and U3966 (N_3966,N_3882,N_3875);
xnor U3967 (N_3967,N_3876,N_3847);
and U3968 (N_3968,N_3821,N_3883);
nand U3969 (N_3969,N_3847,N_3884);
nand U3970 (N_3970,N_3878,N_3831);
or U3971 (N_3971,N_3824,N_3864);
nor U3972 (N_3972,N_3893,N_3849);
nand U3973 (N_3973,N_3806,N_3875);
nand U3974 (N_3974,N_3835,N_3871);
or U3975 (N_3975,N_3823,N_3849);
nor U3976 (N_3976,N_3894,N_3870);
nor U3977 (N_3977,N_3817,N_3846);
xor U3978 (N_3978,N_3869,N_3810);
or U3979 (N_3979,N_3887,N_3871);
or U3980 (N_3980,N_3835,N_3884);
nor U3981 (N_3981,N_3813,N_3854);
nand U3982 (N_3982,N_3899,N_3852);
or U3983 (N_3983,N_3834,N_3845);
or U3984 (N_3984,N_3848,N_3866);
xor U3985 (N_3985,N_3823,N_3841);
nand U3986 (N_3986,N_3827,N_3836);
nand U3987 (N_3987,N_3861,N_3832);
xnor U3988 (N_3988,N_3800,N_3890);
nor U3989 (N_3989,N_3801,N_3821);
nand U3990 (N_3990,N_3884,N_3870);
and U3991 (N_3991,N_3876,N_3862);
xnor U3992 (N_3992,N_3839,N_3887);
nor U3993 (N_3993,N_3800,N_3855);
nor U3994 (N_3994,N_3859,N_3848);
or U3995 (N_3995,N_3878,N_3810);
xor U3996 (N_3996,N_3898,N_3827);
nand U3997 (N_3997,N_3878,N_3898);
and U3998 (N_3998,N_3818,N_3894);
nor U3999 (N_3999,N_3830,N_3811);
nand U4000 (N_4000,N_3934,N_3909);
or U4001 (N_4001,N_3932,N_3935);
nor U4002 (N_4002,N_3978,N_3941);
nand U4003 (N_4003,N_3956,N_3971);
xnor U4004 (N_4004,N_3915,N_3949);
xnor U4005 (N_4005,N_3994,N_3986);
and U4006 (N_4006,N_3985,N_3925);
nor U4007 (N_4007,N_3951,N_3976);
or U4008 (N_4008,N_3902,N_3983);
nand U4009 (N_4009,N_3900,N_3953);
nor U4010 (N_4010,N_3995,N_3920);
or U4011 (N_4011,N_3905,N_3926);
nand U4012 (N_4012,N_3962,N_3943);
nand U4013 (N_4013,N_3945,N_3931);
and U4014 (N_4014,N_3910,N_3969);
xnor U4015 (N_4015,N_3992,N_3991);
nand U4016 (N_4016,N_3924,N_3997);
and U4017 (N_4017,N_3998,N_3947);
xor U4018 (N_4018,N_3963,N_3955);
nand U4019 (N_4019,N_3903,N_3946);
and U4020 (N_4020,N_3959,N_3929);
and U4021 (N_4021,N_3950,N_3993);
nor U4022 (N_4022,N_3906,N_3927);
and U4023 (N_4023,N_3936,N_3973);
or U4024 (N_4024,N_3921,N_3988);
or U4025 (N_4025,N_3967,N_3948);
or U4026 (N_4026,N_3960,N_3970);
or U4027 (N_4027,N_3979,N_3982);
xnor U4028 (N_4028,N_3972,N_3964);
nand U4029 (N_4029,N_3981,N_3965);
nand U4030 (N_4030,N_3954,N_3937);
or U4031 (N_4031,N_3919,N_3916);
xor U4032 (N_4032,N_3907,N_3975);
and U4033 (N_4033,N_3966,N_3958);
or U4034 (N_4034,N_3996,N_3928);
and U4035 (N_4035,N_3939,N_3904);
and U4036 (N_4036,N_3930,N_3974);
and U4037 (N_4037,N_3914,N_3908);
xnor U4038 (N_4038,N_3922,N_3913);
or U4039 (N_4039,N_3990,N_3999);
and U4040 (N_4040,N_3933,N_3957);
nand U4041 (N_4041,N_3912,N_3987);
nor U4042 (N_4042,N_3917,N_3901);
xnor U4043 (N_4043,N_3938,N_3989);
xor U4044 (N_4044,N_3940,N_3984);
xnor U4045 (N_4045,N_3952,N_3911);
nor U4046 (N_4046,N_3944,N_3968);
nor U4047 (N_4047,N_3977,N_3961);
xor U4048 (N_4048,N_3942,N_3918);
or U4049 (N_4049,N_3980,N_3923);
nor U4050 (N_4050,N_3975,N_3955);
nor U4051 (N_4051,N_3934,N_3936);
and U4052 (N_4052,N_3950,N_3970);
nand U4053 (N_4053,N_3953,N_3918);
nand U4054 (N_4054,N_3998,N_3927);
nand U4055 (N_4055,N_3971,N_3980);
or U4056 (N_4056,N_3970,N_3909);
and U4057 (N_4057,N_3911,N_3901);
nand U4058 (N_4058,N_3920,N_3975);
nor U4059 (N_4059,N_3957,N_3999);
nor U4060 (N_4060,N_3909,N_3994);
and U4061 (N_4061,N_3985,N_3969);
or U4062 (N_4062,N_3905,N_3963);
nor U4063 (N_4063,N_3924,N_3904);
or U4064 (N_4064,N_3997,N_3992);
and U4065 (N_4065,N_3939,N_3922);
nor U4066 (N_4066,N_3909,N_3953);
or U4067 (N_4067,N_3940,N_3935);
nand U4068 (N_4068,N_3977,N_3994);
or U4069 (N_4069,N_3997,N_3953);
and U4070 (N_4070,N_3918,N_3937);
or U4071 (N_4071,N_3993,N_3980);
nor U4072 (N_4072,N_3957,N_3911);
nand U4073 (N_4073,N_3904,N_3913);
nand U4074 (N_4074,N_3963,N_3935);
and U4075 (N_4075,N_3978,N_3913);
nor U4076 (N_4076,N_3989,N_3956);
nor U4077 (N_4077,N_3945,N_3980);
nand U4078 (N_4078,N_3964,N_3942);
nand U4079 (N_4079,N_3927,N_3946);
or U4080 (N_4080,N_3996,N_3940);
xnor U4081 (N_4081,N_3932,N_3976);
nor U4082 (N_4082,N_3988,N_3945);
or U4083 (N_4083,N_3993,N_3960);
or U4084 (N_4084,N_3937,N_3998);
xor U4085 (N_4085,N_3983,N_3904);
nand U4086 (N_4086,N_3922,N_3947);
xor U4087 (N_4087,N_3916,N_3973);
nand U4088 (N_4088,N_3956,N_3978);
nand U4089 (N_4089,N_3997,N_3929);
and U4090 (N_4090,N_3981,N_3946);
nor U4091 (N_4091,N_3969,N_3947);
or U4092 (N_4092,N_3964,N_3908);
and U4093 (N_4093,N_3988,N_3927);
xnor U4094 (N_4094,N_3980,N_3981);
xnor U4095 (N_4095,N_3964,N_3975);
or U4096 (N_4096,N_3907,N_3940);
and U4097 (N_4097,N_3904,N_3982);
nand U4098 (N_4098,N_3922,N_3954);
xor U4099 (N_4099,N_3907,N_3954);
or U4100 (N_4100,N_4025,N_4014);
nand U4101 (N_4101,N_4022,N_4080);
or U4102 (N_4102,N_4030,N_4090);
nand U4103 (N_4103,N_4049,N_4086);
and U4104 (N_4104,N_4092,N_4037);
xnor U4105 (N_4105,N_4088,N_4012);
nor U4106 (N_4106,N_4020,N_4028);
xnor U4107 (N_4107,N_4074,N_4091);
and U4108 (N_4108,N_4076,N_4057);
nor U4109 (N_4109,N_4003,N_4061);
nor U4110 (N_4110,N_4045,N_4042);
nand U4111 (N_4111,N_4089,N_4084);
or U4112 (N_4112,N_4078,N_4079);
and U4113 (N_4113,N_4032,N_4008);
xor U4114 (N_4114,N_4058,N_4070);
and U4115 (N_4115,N_4072,N_4063);
nor U4116 (N_4116,N_4095,N_4098);
nand U4117 (N_4117,N_4009,N_4011);
or U4118 (N_4118,N_4067,N_4062);
and U4119 (N_4119,N_4016,N_4059);
or U4120 (N_4120,N_4017,N_4006);
xnor U4121 (N_4121,N_4060,N_4043);
and U4122 (N_4122,N_4015,N_4064);
and U4123 (N_4123,N_4066,N_4093);
nor U4124 (N_4124,N_4035,N_4085);
or U4125 (N_4125,N_4082,N_4010);
and U4126 (N_4126,N_4018,N_4021);
or U4127 (N_4127,N_4039,N_4099);
or U4128 (N_4128,N_4046,N_4094);
nand U4129 (N_4129,N_4002,N_4096);
and U4130 (N_4130,N_4050,N_4068);
xor U4131 (N_4131,N_4024,N_4007);
nor U4132 (N_4132,N_4054,N_4081);
nand U4133 (N_4133,N_4077,N_4097);
xor U4134 (N_4134,N_4029,N_4033);
nor U4135 (N_4135,N_4026,N_4052);
nand U4136 (N_4136,N_4056,N_4065);
nor U4137 (N_4137,N_4027,N_4040);
xnor U4138 (N_4138,N_4053,N_4004);
xor U4139 (N_4139,N_4005,N_4048);
xor U4140 (N_4140,N_4038,N_4031);
xnor U4141 (N_4141,N_4023,N_4044);
and U4142 (N_4142,N_4000,N_4055);
nand U4143 (N_4143,N_4047,N_4041);
nand U4144 (N_4144,N_4071,N_4013);
nand U4145 (N_4145,N_4069,N_4075);
and U4146 (N_4146,N_4034,N_4036);
nand U4147 (N_4147,N_4083,N_4001);
xnor U4148 (N_4148,N_4087,N_4019);
xnor U4149 (N_4149,N_4073,N_4051);
nor U4150 (N_4150,N_4030,N_4088);
or U4151 (N_4151,N_4062,N_4068);
or U4152 (N_4152,N_4047,N_4061);
or U4153 (N_4153,N_4020,N_4006);
or U4154 (N_4154,N_4027,N_4029);
nor U4155 (N_4155,N_4000,N_4097);
or U4156 (N_4156,N_4098,N_4062);
nand U4157 (N_4157,N_4025,N_4009);
and U4158 (N_4158,N_4090,N_4041);
xor U4159 (N_4159,N_4098,N_4084);
nor U4160 (N_4160,N_4092,N_4084);
nor U4161 (N_4161,N_4082,N_4078);
nor U4162 (N_4162,N_4038,N_4047);
nand U4163 (N_4163,N_4012,N_4089);
xnor U4164 (N_4164,N_4052,N_4060);
xor U4165 (N_4165,N_4062,N_4038);
nand U4166 (N_4166,N_4032,N_4099);
and U4167 (N_4167,N_4060,N_4054);
or U4168 (N_4168,N_4062,N_4053);
or U4169 (N_4169,N_4099,N_4037);
nor U4170 (N_4170,N_4033,N_4098);
nor U4171 (N_4171,N_4034,N_4064);
nand U4172 (N_4172,N_4080,N_4098);
or U4173 (N_4173,N_4084,N_4028);
xnor U4174 (N_4174,N_4014,N_4058);
and U4175 (N_4175,N_4042,N_4047);
and U4176 (N_4176,N_4042,N_4009);
xor U4177 (N_4177,N_4029,N_4071);
and U4178 (N_4178,N_4057,N_4025);
nand U4179 (N_4179,N_4018,N_4089);
nand U4180 (N_4180,N_4008,N_4039);
xnor U4181 (N_4181,N_4091,N_4060);
nor U4182 (N_4182,N_4095,N_4094);
nor U4183 (N_4183,N_4037,N_4086);
or U4184 (N_4184,N_4087,N_4064);
or U4185 (N_4185,N_4094,N_4048);
nand U4186 (N_4186,N_4039,N_4010);
and U4187 (N_4187,N_4018,N_4004);
xor U4188 (N_4188,N_4082,N_4028);
nand U4189 (N_4189,N_4083,N_4070);
nand U4190 (N_4190,N_4035,N_4060);
xnor U4191 (N_4191,N_4058,N_4081);
nand U4192 (N_4192,N_4063,N_4096);
or U4193 (N_4193,N_4075,N_4073);
xor U4194 (N_4194,N_4056,N_4055);
nand U4195 (N_4195,N_4015,N_4083);
nor U4196 (N_4196,N_4068,N_4009);
or U4197 (N_4197,N_4099,N_4033);
nor U4198 (N_4198,N_4081,N_4021);
xor U4199 (N_4199,N_4054,N_4011);
or U4200 (N_4200,N_4124,N_4113);
nor U4201 (N_4201,N_4197,N_4118);
xnor U4202 (N_4202,N_4138,N_4162);
nor U4203 (N_4203,N_4192,N_4125);
and U4204 (N_4204,N_4190,N_4189);
nor U4205 (N_4205,N_4196,N_4149);
or U4206 (N_4206,N_4155,N_4115);
nor U4207 (N_4207,N_4116,N_4133);
xor U4208 (N_4208,N_4156,N_4121);
and U4209 (N_4209,N_4104,N_4117);
or U4210 (N_4210,N_4161,N_4164);
or U4211 (N_4211,N_4131,N_4129);
xor U4212 (N_4212,N_4168,N_4195);
nand U4213 (N_4213,N_4109,N_4150);
xnor U4214 (N_4214,N_4185,N_4144);
and U4215 (N_4215,N_4176,N_4140);
nor U4216 (N_4216,N_4169,N_4148);
and U4217 (N_4217,N_4163,N_4100);
xor U4218 (N_4218,N_4101,N_4122);
nand U4219 (N_4219,N_4105,N_4154);
xnor U4220 (N_4220,N_4183,N_4191);
and U4221 (N_4221,N_4132,N_4119);
and U4222 (N_4222,N_4174,N_4160);
or U4223 (N_4223,N_4120,N_4199);
or U4224 (N_4224,N_4186,N_4159);
or U4225 (N_4225,N_4193,N_4142);
and U4226 (N_4226,N_4108,N_4103);
or U4227 (N_4227,N_4146,N_4110);
or U4228 (N_4228,N_4127,N_4166);
and U4229 (N_4229,N_4145,N_4187);
or U4230 (N_4230,N_4143,N_4152);
or U4231 (N_4231,N_4111,N_4181);
nand U4232 (N_4232,N_4123,N_4158);
nand U4233 (N_4233,N_4128,N_4171);
and U4234 (N_4234,N_4165,N_4112);
nand U4235 (N_4235,N_4141,N_4114);
xor U4236 (N_4236,N_4182,N_4175);
xnor U4237 (N_4237,N_4135,N_4177);
nor U4238 (N_4238,N_4151,N_4106);
and U4239 (N_4239,N_4172,N_4107);
nand U4240 (N_4240,N_4170,N_4147);
xor U4241 (N_4241,N_4194,N_4184);
nor U4242 (N_4242,N_4198,N_4178);
or U4243 (N_4243,N_4157,N_4134);
or U4244 (N_4244,N_4180,N_4188);
and U4245 (N_4245,N_4173,N_4167);
or U4246 (N_4246,N_4126,N_4136);
nor U4247 (N_4247,N_4130,N_4153);
xor U4248 (N_4248,N_4137,N_4139);
xor U4249 (N_4249,N_4102,N_4179);
xor U4250 (N_4250,N_4126,N_4158);
or U4251 (N_4251,N_4155,N_4146);
and U4252 (N_4252,N_4161,N_4131);
nor U4253 (N_4253,N_4169,N_4179);
and U4254 (N_4254,N_4103,N_4173);
and U4255 (N_4255,N_4174,N_4129);
xnor U4256 (N_4256,N_4192,N_4106);
nor U4257 (N_4257,N_4115,N_4136);
and U4258 (N_4258,N_4130,N_4113);
and U4259 (N_4259,N_4168,N_4186);
and U4260 (N_4260,N_4181,N_4109);
or U4261 (N_4261,N_4174,N_4100);
nor U4262 (N_4262,N_4140,N_4117);
nand U4263 (N_4263,N_4164,N_4181);
nand U4264 (N_4264,N_4176,N_4149);
or U4265 (N_4265,N_4161,N_4193);
nor U4266 (N_4266,N_4124,N_4172);
and U4267 (N_4267,N_4169,N_4156);
or U4268 (N_4268,N_4138,N_4158);
nor U4269 (N_4269,N_4124,N_4126);
xor U4270 (N_4270,N_4147,N_4129);
or U4271 (N_4271,N_4119,N_4138);
xnor U4272 (N_4272,N_4192,N_4145);
nand U4273 (N_4273,N_4175,N_4126);
and U4274 (N_4274,N_4105,N_4182);
nand U4275 (N_4275,N_4161,N_4187);
or U4276 (N_4276,N_4178,N_4126);
or U4277 (N_4277,N_4198,N_4148);
nor U4278 (N_4278,N_4196,N_4136);
nor U4279 (N_4279,N_4104,N_4169);
nand U4280 (N_4280,N_4144,N_4128);
or U4281 (N_4281,N_4102,N_4174);
or U4282 (N_4282,N_4186,N_4135);
xnor U4283 (N_4283,N_4113,N_4155);
nor U4284 (N_4284,N_4197,N_4131);
nor U4285 (N_4285,N_4134,N_4114);
xor U4286 (N_4286,N_4136,N_4122);
xor U4287 (N_4287,N_4124,N_4102);
nor U4288 (N_4288,N_4111,N_4110);
nor U4289 (N_4289,N_4119,N_4108);
xnor U4290 (N_4290,N_4184,N_4103);
or U4291 (N_4291,N_4187,N_4192);
and U4292 (N_4292,N_4109,N_4166);
nand U4293 (N_4293,N_4119,N_4131);
nand U4294 (N_4294,N_4130,N_4185);
and U4295 (N_4295,N_4107,N_4180);
or U4296 (N_4296,N_4176,N_4133);
and U4297 (N_4297,N_4162,N_4159);
nand U4298 (N_4298,N_4166,N_4141);
nand U4299 (N_4299,N_4129,N_4171);
or U4300 (N_4300,N_4235,N_4276);
xor U4301 (N_4301,N_4206,N_4217);
or U4302 (N_4302,N_4254,N_4292);
or U4303 (N_4303,N_4277,N_4234);
and U4304 (N_4304,N_4255,N_4211);
nand U4305 (N_4305,N_4257,N_4222);
nand U4306 (N_4306,N_4230,N_4214);
xor U4307 (N_4307,N_4262,N_4231);
or U4308 (N_4308,N_4295,N_4224);
nand U4309 (N_4309,N_4250,N_4291);
nand U4310 (N_4310,N_4202,N_4243);
or U4311 (N_4311,N_4218,N_4248);
nor U4312 (N_4312,N_4278,N_4282);
or U4313 (N_4313,N_4239,N_4207);
or U4314 (N_4314,N_4273,N_4251);
or U4315 (N_4315,N_4256,N_4299);
xor U4316 (N_4316,N_4237,N_4279);
and U4317 (N_4317,N_4280,N_4210);
or U4318 (N_4318,N_4260,N_4221);
nand U4319 (N_4319,N_4200,N_4223);
nand U4320 (N_4320,N_4227,N_4212);
nand U4321 (N_4321,N_4269,N_4252);
and U4322 (N_4322,N_4209,N_4268);
nor U4323 (N_4323,N_4274,N_4245);
or U4324 (N_4324,N_4275,N_4205);
nor U4325 (N_4325,N_4242,N_4265);
and U4326 (N_4326,N_4246,N_4287);
xor U4327 (N_4327,N_4232,N_4293);
or U4328 (N_4328,N_4238,N_4288);
or U4329 (N_4329,N_4215,N_4261);
and U4330 (N_4330,N_4247,N_4226);
nand U4331 (N_4331,N_4270,N_4263);
or U4332 (N_4332,N_4281,N_4219);
xnor U4333 (N_4333,N_4297,N_4208);
xor U4334 (N_4334,N_4290,N_4244);
or U4335 (N_4335,N_4272,N_4284);
nand U4336 (N_4336,N_4298,N_4220);
nor U4337 (N_4337,N_4286,N_4225);
or U4338 (N_4338,N_4229,N_4259);
or U4339 (N_4339,N_4285,N_4264);
xnor U4340 (N_4340,N_4267,N_4271);
nor U4341 (N_4341,N_4294,N_4258);
or U4342 (N_4342,N_4283,N_4216);
nor U4343 (N_4343,N_4241,N_4289);
or U4344 (N_4344,N_4204,N_4240);
nand U4345 (N_4345,N_4249,N_4296);
or U4346 (N_4346,N_4213,N_4236);
nor U4347 (N_4347,N_4266,N_4201);
xnor U4348 (N_4348,N_4253,N_4233);
nor U4349 (N_4349,N_4203,N_4228);
nand U4350 (N_4350,N_4257,N_4215);
nor U4351 (N_4351,N_4255,N_4213);
xor U4352 (N_4352,N_4295,N_4251);
and U4353 (N_4353,N_4208,N_4222);
nand U4354 (N_4354,N_4260,N_4258);
nand U4355 (N_4355,N_4251,N_4269);
nand U4356 (N_4356,N_4262,N_4200);
and U4357 (N_4357,N_4277,N_4275);
nor U4358 (N_4358,N_4242,N_4251);
xor U4359 (N_4359,N_4289,N_4226);
nand U4360 (N_4360,N_4234,N_4223);
nor U4361 (N_4361,N_4278,N_4296);
nand U4362 (N_4362,N_4262,N_4263);
nand U4363 (N_4363,N_4218,N_4288);
or U4364 (N_4364,N_4237,N_4229);
nor U4365 (N_4365,N_4254,N_4203);
or U4366 (N_4366,N_4298,N_4275);
or U4367 (N_4367,N_4292,N_4229);
xor U4368 (N_4368,N_4224,N_4297);
and U4369 (N_4369,N_4297,N_4251);
nand U4370 (N_4370,N_4240,N_4262);
xnor U4371 (N_4371,N_4290,N_4242);
nor U4372 (N_4372,N_4224,N_4245);
or U4373 (N_4373,N_4272,N_4250);
nor U4374 (N_4374,N_4216,N_4237);
xnor U4375 (N_4375,N_4249,N_4230);
nor U4376 (N_4376,N_4222,N_4202);
nand U4377 (N_4377,N_4254,N_4264);
nand U4378 (N_4378,N_4286,N_4224);
nand U4379 (N_4379,N_4264,N_4225);
or U4380 (N_4380,N_4290,N_4243);
or U4381 (N_4381,N_4280,N_4291);
nor U4382 (N_4382,N_4263,N_4298);
nand U4383 (N_4383,N_4283,N_4264);
and U4384 (N_4384,N_4283,N_4277);
and U4385 (N_4385,N_4286,N_4269);
nand U4386 (N_4386,N_4216,N_4289);
nor U4387 (N_4387,N_4253,N_4285);
nor U4388 (N_4388,N_4258,N_4259);
nor U4389 (N_4389,N_4271,N_4236);
xnor U4390 (N_4390,N_4289,N_4234);
nand U4391 (N_4391,N_4288,N_4226);
nand U4392 (N_4392,N_4298,N_4294);
xor U4393 (N_4393,N_4263,N_4249);
nor U4394 (N_4394,N_4251,N_4267);
nor U4395 (N_4395,N_4241,N_4263);
nand U4396 (N_4396,N_4264,N_4293);
or U4397 (N_4397,N_4299,N_4279);
nand U4398 (N_4398,N_4296,N_4235);
and U4399 (N_4399,N_4283,N_4227);
xor U4400 (N_4400,N_4396,N_4328);
nor U4401 (N_4401,N_4378,N_4361);
xor U4402 (N_4402,N_4379,N_4332);
xor U4403 (N_4403,N_4301,N_4367);
nor U4404 (N_4404,N_4347,N_4334);
and U4405 (N_4405,N_4393,N_4356);
nand U4406 (N_4406,N_4380,N_4304);
nor U4407 (N_4407,N_4398,N_4300);
nor U4408 (N_4408,N_4302,N_4359);
nor U4409 (N_4409,N_4349,N_4331);
nand U4410 (N_4410,N_4314,N_4366);
xnor U4411 (N_4411,N_4386,N_4310);
nand U4412 (N_4412,N_4390,N_4374);
and U4413 (N_4413,N_4348,N_4344);
nor U4414 (N_4414,N_4355,N_4372);
nand U4415 (N_4415,N_4337,N_4336);
nand U4416 (N_4416,N_4354,N_4353);
and U4417 (N_4417,N_4381,N_4322);
xor U4418 (N_4418,N_4341,N_4320);
nand U4419 (N_4419,N_4307,N_4329);
nor U4420 (N_4420,N_4382,N_4357);
xor U4421 (N_4421,N_4313,N_4387);
and U4422 (N_4422,N_4338,N_4309);
xnor U4423 (N_4423,N_4364,N_4317);
nand U4424 (N_4424,N_4391,N_4335);
nor U4425 (N_4425,N_4345,N_4315);
xor U4426 (N_4426,N_4318,N_4326);
xnor U4427 (N_4427,N_4308,N_4389);
or U4428 (N_4428,N_4360,N_4312);
nor U4429 (N_4429,N_4333,N_4395);
or U4430 (N_4430,N_4316,N_4394);
nor U4431 (N_4431,N_4384,N_4365);
nand U4432 (N_4432,N_4311,N_4397);
nand U4433 (N_4433,N_4392,N_4376);
or U4434 (N_4434,N_4305,N_4399);
xnor U4435 (N_4435,N_4369,N_4385);
nor U4436 (N_4436,N_4321,N_4383);
or U4437 (N_4437,N_4375,N_4330);
and U4438 (N_4438,N_4368,N_4371);
xnor U4439 (N_4439,N_4388,N_4358);
and U4440 (N_4440,N_4363,N_4325);
and U4441 (N_4441,N_4352,N_4373);
nor U4442 (N_4442,N_4346,N_4343);
and U4443 (N_4443,N_4339,N_4350);
nor U4444 (N_4444,N_4351,N_4327);
nand U4445 (N_4445,N_4370,N_4342);
or U4446 (N_4446,N_4340,N_4324);
nor U4447 (N_4447,N_4377,N_4319);
and U4448 (N_4448,N_4323,N_4303);
nor U4449 (N_4449,N_4306,N_4362);
and U4450 (N_4450,N_4333,N_4386);
or U4451 (N_4451,N_4323,N_4368);
xor U4452 (N_4452,N_4396,N_4390);
xnor U4453 (N_4453,N_4331,N_4303);
and U4454 (N_4454,N_4350,N_4305);
or U4455 (N_4455,N_4359,N_4313);
nand U4456 (N_4456,N_4369,N_4329);
or U4457 (N_4457,N_4374,N_4398);
nand U4458 (N_4458,N_4333,N_4370);
nand U4459 (N_4459,N_4305,N_4336);
or U4460 (N_4460,N_4383,N_4305);
xnor U4461 (N_4461,N_4345,N_4312);
or U4462 (N_4462,N_4338,N_4399);
nand U4463 (N_4463,N_4387,N_4330);
and U4464 (N_4464,N_4342,N_4375);
nor U4465 (N_4465,N_4339,N_4360);
nor U4466 (N_4466,N_4387,N_4376);
and U4467 (N_4467,N_4331,N_4383);
nand U4468 (N_4468,N_4311,N_4307);
nor U4469 (N_4469,N_4323,N_4356);
and U4470 (N_4470,N_4300,N_4399);
nor U4471 (N_4471,N_4346,N_4327);
or U4472 (N_4472,N_4328,N_4379);
and U4473 (N_4473,N_4385,N_4381);
or U4474 (N_4474,N_4346,N_4360);
and U4475 (N_4475,N_4354,N_4314);
nand U4476 (N_4476,N_4390,N_4337);
nand U4477 (N_4477,N_4303,N_4344);
nor U4478 (N_4478,N_4386,N_4330);
nand U4479 (N_4479,N_4334,N_4397);
nor U4480 (N_4480,N_4395,N_4343);
or U4481 (N_4481,N_4342,N_4318);
and U4482 (N_4482,N_4334,N_4354);
xnor U4483 (N_4483,N_4396,N_4368);
nor U4484 (N_4484,N_4399,N_4371);
xor U4485 (N_4485,N_4325,N_4331);
and U4486 (N_4486,N_4397,N_4345);
and U4487 (N_4487,N_4371,N_4324);
nand U4488 (N_4488,N_4324,N_4374);
nand U4489 (N_4489,N_4340,N_4390);
xor U4490 (N_4490,N_4330,N_4389);
and U4491 (N_4491,N_4326,N_4367);
or U4492 (N_4492,N_4361,N_4399);
nand U4493 (N_4493,N_4364,N_4386);
nor U4494 (N_4494,N_4300,N_4394);
and U4495 (N_4495,N_4303,N_4320);
and U4496 (N_4496,N_4362,N_4308);
nor U4497 (N_4497,N_4362,N_4395);
nor U4498 (N_4498,N_4304,N_4384);
and U4499 (N_4499,N_4366,N_4363);
and U4500 (N_4500,N_4434,N_4466);
nand U4501 (N_4501,N_4482,N_4453);
and U4502 (N_4502,N_4454,N_4435);
or U4503 (N_4503,N_4418,N_4451);
nand U4504 (N_4504,N_4440,N_4415);
and U4505 (N_4505,N_4468,N_4413);
and U4506 (N_4506,N_4472,N_4423);
and U4507 (N_4507,N_4474,N_4449);
xor U4508 (N_4508,N_4467,N_4444);
nand U4509 (N_4509,N_4441,N_4475);
xor U4510 (N_4510,N_4490,N_4484);
nand U4511 (N_4511,N_4462,N_4430);
nor U4512 (N_4512,N_4405,N_4414);
nand U4513 (N_4513,N_4412,N_4450);
xor U4514 (N_4514,N_4429,N_4498);
nand U4515 (N_4515,N_4446,N_4481);
or U4516 (N_4516,N_4406,N_4464);
xor U4517 (N_4517,N_4404,N_4433);
and U4518 (N_4518,N_4438,N_4443);
xor U4519 (N_4519,N_4420,N_4458);
and U4520 (N_4520,N_4419,N_4447);
nand U4521 (N_4521,N_4428,N_4456);
nand U4522 (N_4522,N_4410,N_4496);
or U4523 (N_4523,N_4457,N_4480);
nand U4524 (N_4524,N_4465,N_4460);
nand U4525 (N_4525,N_4494,N_4495);
or U4526 (N_4526,N_4424,N_4479);
nand U4527 (N_4527,N_4483,N_4452);
nand U4528 (N_4528,N_4499,N_4455);
nor U4529 (N_4529,N_4432,N_4470);
or U4530 (N_4530,N_4476,N_4477);
and U4531 (N_4531,N_4426,N_4488);
or U4532 (N_4532,N_4437,N_4448);
nand U4533 (N_4533,N_4493,N_4497);
nand U4534 (N_4534,N_4411,N_4469);
nand U4535 (N_4535,N_4409,N_4459);
and U4536 (N_4536,N_4485,N_4436);
or U4537 (N_4537,N_4463,N_4402);
nand U4538 (N_4538,N_4416,N_4417);
xor U4539 (N_4539,N_4471,N_4407);
nor U4540 (N_4540,N_4492,N_4478);
nand U4541 (N_4541,N_4461,N_4491);
xnor U4542 (N_4542,N_4425,N_4427);
xor U4543 (N_4543,N_4442,N_4431);
and U4544 (N_4544,N_4486,N_4489);
or U4545 (N_4545,N_4401,N_4408);
nor U4546 (N_4546,N_4445,N_4422);
nor U4547 (N_4547,N_4421,N_4400);
xor U4548 (N_4548,N_4487,N_4403);
and U4549 (N_4549,N_4473,N_4439);
xor U4550 (N_4550,N_4456,N_4429);
xnor U4551 (N_4551,N_4415,N_4418);
nand U4552 (N_4552,N_4440,N_4485);
and U4553 (N_4553,N_4400,N_4431);
nor U4554 (N_4554,N_4416,N_4444);
or U4555 (N_4555,N_4403,N_4469);
or U4556 (N_4556,N_4491,N_4453);
nor U4557 (N_4557,N_4427,N_4430);
or U4558 (N_4558,N_4439,N_4470);
and U4559 (N_4559,N_4403,N_4443);
or U4560 (N_4560,N_4497,N_4473);
or U4561 (N_4561,N_4402,N_4496);
xnor U4562 (N_4562,N_4424,N_4427);
xnor U4563 (N_4563,N_4422,N_4440);
nand U4564 (N_4564,N_4482,N_4404);
and U4565 (N_4565,N_4400,N_4488);
nor U4566 (N_4566,N_4459,N_4463);
and U4567 (N_4567,N_4449,N_4402);
xnor U4568 (N_4568,N_4452,N_4446);
nand U4569 (N_4569,N_4408,N_4476);
xnor U4570 (N_4570,N_4447,N_4442);
nor U4571 (N_4571,N_4430,N_4481);
nand U4572 (N_4572,N_4405,N_4443);
nor U4573 (N_4573,N_4428,N_4411);
or U4574 (N_4574,N_4417,N_4406);
xnor U4575 (N_4575,N_4438,N_4426);
nand U4576 (N_4576,N_4447,N_4472);
and U4577 (N_4577,N_4469,N_4444);
xnor U4578 (N_4578,N_4401,N_4472);
and U4579 (N_4579,N_4424,N_4477);
and U4580 (N_4580,N_4461,N_4459);
or U4581 (N_4581,N_4422,N_4467);
and U4582 (N_4582,N_4453,N_4493);
nor U4583 (N_4583,N_4471,N_4497);
xnor U4584 (N_4584,N_4493,N_4475);
xor U4585 (N_4585,N_4458,N_4481);
or U4586 (N_4586,N_4469,N_4423);
xnor U4587 (N_4587,N_4491,N_4464);
and U4588 (N_4588,N_4449,N_4425);
nand U4589 (N_4589,N_4413,N_4478);
nand U4590 (N_4590,N_4471,N_4448);
xor U4591 (N_4591,N_4486,N_4429);
xor U4592 (N_4592,N_4481,N_4489);
nor U4593 (N_4593,N_4420,N_4405);
nor U4594 (N_4594,N_4429,N_4463);
and U4595 (N_4595,N_4411,N_4402);
and U4596 (N_4596,N_4491,N_4404);
and U4597 (N_4597,N_4450,N_4492);
nand U4598 (N_4598,N_4458,N_4423);
nor U4599 (N_4599,N_4484,N_4405);
and U4600 (N_4600,N_4519,N_4552);
nor U4601 (N_4601,N_4580,N_4558);
and U4602 (N_4602,N_4557,N_4527);
nor U4603 (N_4603,N_4595,N_4537);
nor U4604 (N_4604,N_4512,N_4530);
nand U4605 (N_4605,N_4506,N_4590);
and U4606 (N_4606,N_4539,N_4501);
and U4607 (N_4607,N_4518,N_4500);
or U4608 (N_4608,N_4520,N_4572);
xnor U4609 (N_4609,N_4589,N_4591);
and U4610 (N_4610,N_4560,N_4551);
and U4611 (N_4611,N_4599,N_4581);
nor U4612 (N_4612,N_4575,N_4579);
and U4613 (N_4613,N_4505,N_4542);
nor U4614 (N_4614,N_4521,N_4561);
and U4615 (N_4615,N_4574,N_4514);
or U4616 (N_4616,N_4546,N_4577);
nor U4617 (N_4617,N_4503,N_4523);
and U4618 (N_4618,N_4508,N_4531);
nor U4619 (N_4619,N_4532,N_4540);
xor U4620 (N_4620,N_4550,N_4536);
nor U4621 (N_4621,N_4522,N_4555);
nor U4622 (N_4622,N_4568,N_4563);
or U4623 (N_4623,N_4596,N_4524);
or U4624 (N_4624,N_4588,N_4593);
nor U4625 (N_4625,N_4544,N_4587);
or U4626 (N_4626,N_4571,N_4516);
nand U4627 (N_4627,N_4556,N_4549);
xor U4628 (N_4628,N_4598,N_4597);
xor U4629 (N_4629,N_4517,N_4559);
xnor U4630 (N_4630,N_4528,N_4566);
and U4631 (N_4631,N_4535,N_4534);
xnor U4632 (N_4632,N_4576,N_4529);
nand U4633 (N_4633,N_4504,N_4510);
nor U4634 (N_4634,N_4569,N_4509);
nor U4635 (N_4635,N_4573,N_4570);
and U4636 (N_4636,N_4592,N_4565);
or U4637 (N_4637,N_4533,N_4511);
nor U4638 (N_4638,N_4526,N_4564);
and U4639 (N_4639,N_4525,N_4562);
nand U4640 (N_4640,N_4507,N_4578);
nand U4641 (N_4641,N_4554,N_4584);
or U4642 (N_4642,N_4541,N_4543);
and U4643 (N_4643,N_4553,N_4547);
or U4644 (N_4644,N_4515,N_4585);
and U4645 (N_4645,N_4545,N_4567);
and U4646 (N_4646,N_4582,N_4513);
nand U4647 (N_4647,N_4586,N_4594);
nor U4648 (N_4648,N_4583,N_4538);
or U4649 (N_4649,N_4502,N_4548);
xor U4650 (N_4650,N_4502,N_4537);
and U4651 (N_4651,N_4563,N_4573);
nand U4652 (N_4652,N_4570,N_4562);
xor U4653 (N_4653,N_4550,N_4583);
and U4654 (N_4654,N_4509,N_4500);
or U4655 (N_4655,N_4537,N_4572);
and U4656 (N_4656,N_4596,N_4541);
and U4657 (N_4657,N_4526,N_4561);
xnor U4658 (N_4658,N_4570,N_4517);
and U4659 (N_4659,N_4546,N_4518);
xnor U4660 (N_4660,N_4583,N_4532);
or U4661 (N_4661,N_4514,N_4544);
and U4662 (N_4662,N_4519,N_4563);
and U4663 (N_4663,N_4514,N_4520);
xnor U4664 (N_4664,N_4517,N_4592);
nor U4665 (N_4665,N_4570,N_4540);
and U4666 (N_4666,N_4589,N_4560);
nor U4667 (N_4667,N_4550,N_4594);
xnor U4668 (N_4668,N_4573,N_4502);
xor U4669 (N_4669,N_4598,N_4584);
or U4670 (N_4670,N_4580,N_4541);
or U4671 (N_4671,N_4561,N_4588);
nand U4672 (N_4672,N_4563,N_4548);
nor U4673 (N_4673,N_4509,N_4523);
nor U4674 (N_4674,N_4599,N_4554);
or U4675 (N_4675,N_4576,N_4571);
or U4676 (N_4676,N_4591,N_4542);
and U4677 (N_4677,N_4520,N_4578);
nor U4678 (N_4678,N_4587,N_4592);
xor U4679 (N_4679,N_4504,N_4549);
or U4680 (N_4680,N_4573,N_4516);
and U4681 (N_4681,N_4539,N_4541);
xnor U4682 (N_4682,N_4525,N_4526);
and U4683 (N_4683,N_4564,N_4569);
nand U4684 (N_4684,N_4547,N_4592);
or U4685 (N_4685,N_4546,N_4563);
xnor U4686 (N_4686,N_4535,N_4500);
nor U4687 (N_4687,N_4519,N_4520);
xnor U4688 (N_4688,N_4532,N_4578);
or U4689 (N_4689,N_4599,N_4579);
xor U4690 (N_4690,N_4539,N_4585);
and U4691 (N_4691,N_4596,N_4558);
nor U4692 (N_4692,N_4507,N_4511);
nor U4693 (N_4693,N_4552,N_4558);
nand U4694 (N_4694,N_4588,N_4547);
and U4695 (N_4695,N_4544,N_4513);
nor U4696 (N_4696,N_4516,N_4546);
or U4697 (N_4697,N_4557,N_4582);
or U4698 (N_4698,N_4562,N_4545);
xor U4699 (N_4699,N_4597,N_4517);
or U4700 (N_4700,N_4624,N_4692);
xnor U4701 (N_4701,N_4601,N_4631);
xor U4702 (N_4702,N_4609,N_4616);
or U4703 (N_4703,N_4694,N_4612);
and U4704 (N_4704,N_4604,N_4614);
nor U4705 (N_4705,N_4625,N_4648);
nand U4706 (N_4706,N_4677,N_4646);
xor U4707 (N_4707,N_4608,N_4618);
xnor U4708 (N_4708,N_4663,N_4666);
and U4709 (N_4709,N_4688,N_4623);
nand U4710 (N_4710,N_4647,N_4684);
or U4711 (N_4711,N_4602,N_4665);
nor U4712 (N_4712,N_4613,N_4699);
nor U4713 (N_4713,N_4657,N_4641);
nor U4714 (N_4714,N_4653,N_4680);
nor U4715 (N_4715,N_4644,N_4645);
nor U4716 (N_4716,N_4621,N_4696);
nand U4717 (N_4717,N_4679,N_4635);
nand U4718 (N_4718,N_4670,N_4629);
and U4719 (N_4719,N_4634,N_4676);
and U4720 (N_4720,N_4654,N_4638);
xnor U4721 (N_4721,N_4667,N_4606);
nand U4722 (N_4722,N_4627,N_4697);
nand U4723 (N_4723,N_4682,N_4642);
nand U4724 (N_4724,N_4620,N_4600);
or U4725 (N_4725,N_4632,N_4685);
and U4726 (N_4726,N_4674,N_4690);
nand U4727 (N_4727,N_4649,N_4658);
or U4728 (N_4728,N_4659,N_4671);
or U4729 (N_4729,N_4630,N_4689);
nor U4730 (N_4730,N_4643,N_4622);
and U4731 (N_4731,N_4617,N_4664);
nand U4732 (N_4732,N_4628,N_4675);
and U4733 (N_4733,N_4603,N_4673);
nor U4734 (N_4734,N_4672,N_4611);
nor U4735 (N_4735,N_4637,N_4687);
and U4736 (N_4736,N_4640,N_4691);
or U4737 (N_4737,N_4619,N_4698);
nor U4738 (N_4738,N_4655,N_4660);
or U4739 (N_4739,N_4678,N_4615);
or U4740 (N_4740,N_4650,N_4661);
xnor U4741 (N_4741,N_4633,N_4607);
and U4742 (N_4742,N_4605,N_4681);
or U4743 (N_4743,N_4662,N_4652);
and U4744 (N_4744,N_4651,N_4683);
and U4745 (N_4745,N_4668,N_4695);
or U4746 (N_4746,N_4626,N_4610);
and U4747 (N_4747,N_4693,N_4639);
or U4748 (N_4748,N_4656,N_4686);
or U4749 (N_4749,N_4669,N_4636);
nand U4750 (N_4750,N_4662,N_4640);
or U4751 (N_4751,N_4680,N_4609);
xnor U4752 (N_4752,N_4673,N_4671);
xor U4753 (N_4753,N_4620,N_4662);
or U4754 (N_4754,N_4687,N_4609);
nand U4755 (N_4755,N_4628,N_4656);
nand U4756 (N_4756,N_4646,N_4606);
nand U4757 (N_4757,N_4636,N_4670);
and U4758 (N_4758,N_4688,N_4639);
or U4759 (N_4759,N_4671,N_4656);
nor U4760 (N_4760,N_4640,N_4619);
and U4761 (N_4761,N_4652,N_4670);
nand U4762 (N_4762,N_4683,N_4637);
and U4763 (N_4763,N_4650,N_4652);
and U4764 (N_4764,N_4659,N_4608);
xor U4765 (N_4765,N_4676,N_4602);
or U4766 (N_4766,N_4606,N_4698);
or U4767 (N_4767,N_4606,N_4623);
nand U4768 (N_4768,N_4688,N_4681);
nand U4769 (N_4769,N_4678,N_4632);
and U4770 (N_4770,N_4642,N_4670);
nand U4771 (N_4771,N_4657,N_4684);
and U4772 (N_4772,N_4695,N_4652);
nand U4773 (N_4773,N_4690,N_4675);
or U4774 (N_4774,N_4640,N_4631);
nand U4775 (N_4775,N_4609,N_4602);
and U4776 (N_4776,N_4612,N_4659);
nor U4777 (N_4777,N_4621,N_4644);
nor U4778 (N_4778,N_4673,N_4688);
xnor U4779 (N_4779,N_4677,N_4640);
or U4780 (N_4780,N_4682,N_4635);
nand U4781 (N_4781,N_4682,N_4669);
nand U4782 (N_4782,N_4640,N_4605);
nor U4783 (N_4783,N_4621,N_4601);
xor U4784 (N_4784,N_4686,N_4692);
or U4785 (N_4785,N_4650,N_4618);
nor U4786 (N_4786,N_4649,N_4637);
xnor U4787 (N_4787,N_4688,N_4618);
nand U4788 (N_4788,N_4684,N_4683);
and U4789 (N_4789,N_4681,N_4612);
or U4790 (N_4790,N_4604,N_4644);
or U4791 (N_4791,N_4655,N_4671);
nand U4792 (N_4792,N_4695,N_4686);
xnor U4793 (N_4793,N_4643,N_4682);
and U4794 (N_4794,N_4609,N_4653);
xnor U4795 (N_4795,N_4690,N_4678);
nand U4796 (N_4796,N_4611,N_4643);
xnor U4797 (N_4797,N_4652,N_4677);
nand U4798 (N_4798,N_4635,N_4626);
xnor U4799 (N_4799,N_4689,N_4656);
xnor U4800 (N_4800,N_4766,N_4765);
nor U4801 (N_4801,N_4762,N_4767);
nor U4802 (N_4802,N_4711,N_4764);
nand U4803 (N_4803,N_4744,N_4797);
xor U4804 (N_4804,N_4717,N_4709);
and U4805 (N_4805,N_4719,N_4780);
or U4806 (N_4806,N_4723,N_4735);
or U4807 (N_4807,N_4726,N_4712);
nor U4808 (N_4808,N_4720,N_4704);
xnor U4809 (N_4809,N_4763,N_4787);
or U4810 (N_4810,N_4757,N_4792);
nand U4811 (N_4811,N_4722,N_4736);
nor U4812 (N_4812,N_4786,N_4734);
nor U4813 (N_4813,N_4713,N_4776);
or U4814 (N_4814,N_4741,N_4783);
xnor U4815 (N_4815,N_4739,N_4759);
xnor U4816 (N_4816,N_4707,N_4756);
and U4817 (N_4817,N_4721,N_4751);
and U4818 (N_4818,N_4742,N_4710);
or U4819 (N_4819,N_4724,N_4799);
or U4820 (N_4820,N_4788,N_4702);
xor U4821 (N_4821,N_4705,N_4729);
nand U4822 (N_4822,N_4761,N_4714);
nand U4823 (N_4823,N_4773,N_4774);
nor U4824 (N_4824,N_4778,N_4725);
or U4825 (N_4825,N_4790,N_4769);
and U4826 (N_4826,N_4755,N_4747);
or U4827 (N_4827,N_4775,N_4795);
xnor U4828 (N_4828,N_4701,N_4781);
and U4829 (N_4829,N_4745,N_4703);
and U4830 (N_4830,N_4708,N_4700);
xor U4831 (N_4831,N_4749,N_4748);
nand U4832 (N_4832,N_4754,N_4743);
or U4833 (N_4833,N_4794,N_4715);
xor U4834 (N_4834,N_4737,N_4716);
or U4835 (N_4835,N_4728,N_4784);
or U4836 (N_4836,N_4771,N_4730);
xor U4837 (N_4837,N_4732,N_4777);
nor U4838 (N_4838,N_4758,N_4798);
nand U4839 (N_4839,N_4768,N_4740);
and U4840 (N_4840,N_4793,N_4785);
nor U4841 (N_4841,N_4738,N_4752);
xnor U4842 (N_4842,N_4750,N_4746);
nor U4843 (N_4843,N_4731,N_4789);
or U4844 (N_4844,N_4753,N_4760);
nand U4845 (N_4845,N_4727,N_4706);
and U4846 (N_4846,N_4796,N_4791);
nor U4847 (N_4847,N_4772,N_4718);
xnor U4848 (N_4848,N_4733,N_4779);
nor U4849 (N_4849,N_4782,N_4770);
xnor U4850 (N_4850,N_4779,N_4768);
xnor U4851 (N_4851,N_4792,N_4730);
xor U4852 (N_4852,N_4708,N_4715);
xnor U4853 (N_4853,N_4709,N_4764);
nand U4854 (N_4854,N_4741,N_4749);
nand U4855 (N_4855,N_4794,N_4768);
nand U4856 (N_4856,N_4741,N_4745);
and U4857 (N_4857,N_4794,N_4772);
and U4858 (N_4858,N_4791,N_4767);
nor U4859 (N_4859,N_4764,N_4722);
nor U4860 (N_4860,N_4700,N_4748);
nor U4861 (N_4861,N_4729,N_4734);
nand U4862 (N_4862,N_4790,N_4778);
or U4863 (N_4863,N_4749,N_4792);
or U4864 (N_4864,N_4790,N_4717);
xor U4865 (N_4865,N_4796,N_4782);
or U4866 (N_4866,N_4716,N_4784);
nor U4867 (N_4867,N_4736,N_4743);
and U4868 (N_4868,N_4732,N_4729);
nand U4869 (N_4869,N_4723,N_4700);
xnor U4870 (N_4870,N_4785,N_4736);
or U4871 (N_4871,N_4723,N_4740);
nand U4872 (N_4872,N_4785,N_4777);
and U4873 (N_4873,N_4749,N_4729);
and U4874 (N_4874,N_4732,N_4704);
or U4875 (N_4875,N_4760,N_4721);
or U4876 (N_4876,N_4778,N_4799);
and U4877 (N_4877,N_4779,N_4780);
xor U4878 (N_4878,N_4733,N_4748);
nor U4879 (N_4879,N_4731,N_4705);
nor U4880 (N_4880,N_4720,N_4782);
xor U4881 (N_4881,N_4783,N_4785);
and U4882 (N_4882,N_4738,N_4709);
and U4883 (N_4883,N_4782,N_4768);
and U4884 (N_4884,N_4778,N_4709);
nand U4885 (N_4885,N_4708,N_4749);
nand U4886 (N_4886,N_4725,N_4727);
and U4887 (N_4887,N_4765,N_4705);
nand U4888 (N_4888,N_4739,N_4732);
xnor U4889 (N_4889,N_4742,N_4763);
xnor U4890 (N_4890,N_4737,N_4787);
or U4891 (N_4891,N_4759,N_4723);
nor U4892 (N_4892,N_4779,N_4757);
or U4893 (N_4893,N_4740,N_4792);
xor U4894 (N_4894,N_4725,N_4724);
or U4895 (N_4895,N_4742,N_4729);
xor U4896 (N_4896,N_4732,N_4780);
and U4897 (N_4897,N_4767,N_4774);
and U4898 (N_4898,N_4774,N_4719);
xor U4899 (N_4899,N_4730,N_4779);
nor U4900 (N_4900,N_4890,N_4873);
nor U4901 (N_4901,N_4819,N_4814);
xor U4902 (N_4902,N_4813,N_4855);
and U4903 (N_4903,N_4823,N_4889);
xnor U4904 (N_4904,N_4883,N_4816);
nor U4905 (N_4905,N_4820,N_4830);
or U4906 (N_4906,N_4805,N_4863);
and U4907 (N_4907,N_4858,N_4853);
nor U4908 (N_4908,N_4899,N_4870);
and U4909 (N_4909,N_4840,N_4839);
xor U4910 (N_4910,N_4831,N_4868);
or U4911 (N_4911,N_4829,N_4821);
or U4912 (N_4912,N_4812,N_4886);
and U4913 (N_4913,N_4884,N_4854);
xnor U4914 (N_4914,N_4895,N_4859);
xor U4915 (N_4915,N_4869,N_4826);
xnor U4916 (N_4916,N_4843,N_4896);
and U4917 (N_4917,N_4803,N_4865);
or U4918 (N_4918,N_4887,N_4862);
xor U4919 (N_4919,N_4804,N_4818);
and U4920 (N_4920,N_4898,N_4802);
and U4921 (N_4921,N_4892,N_4817);
nor U4922 (N_4922,N_4842,N_4837);
xor U4923 (N_4923,N_4838,N_4841);
xor U4924 (N_4924,N_4864,N_4801);
xnor U4925 (N_4925,N_4894,N_4891);
xnor U4926 (N_4926,N_4860,N_4893);
or U4927 (N_4927,N_4827,N_4881);
xnor U4928 (N_4928,N_4815,N_4822);
nor U4929 (N_4929,N_4861,N_4879);
nand U4930 (N_4930,N_4825,N_4828);
nor U4931 (N_4931,N_4852,N_4888);
or U4932 (N_4932,N_4836,N_4848);
or U4933 (N_4933,N_4846,N_4844);
nand U4934 (N_4934,N_4800,N_4847);
nor U4935 (N_4935,N_4857,N_4850);
nor U4936 (N_4936,N_4810,N_4834);
or U4937 (N_4937,N_4807,N_4876);
nor U4938 (N_4938,N_4809,N_4845);
and U4939 (N_4939,N_4811,N_4877);
or U4940 (N_4940,N_4866,N_4856);
and U4941 (N_4941,N_4851,N_4867);
or U4942 (N_4942,N_4875,N_4878);
nand U4943 (N_4943,N_4880,N_4885);
and U4944 (N_4944,N_4824,N_4897);
xnor U4945 (N_4945,N_4874,N_4871);
nor U4946 (N_4946,N_4849,N_4835);
nor U4947 (N_4947,N_4882,N_4808);
or U4948 (N_4948,N_4832,N_4872);
nand U4949 (N_4949,N_4806,N_4833);
and U4950 (N_4950,N_4811,N_4844);
or U4951 (N_4951,N_4888,N_4881);
and U4952 (N_4952,N_4862,N_4846);
xnor U4953 (N_4953,N_4828,N_4899);
nand U4954 (N_4954,N_4865,N_4813);
or U4955 (N_4955,N_4807,N_4812);
xor U4956 (N_4956,N_4854,N_4881);
or U4957 (N_4957,N_4874,N_4895);
or U4958 (N_4958,N_4846,N_4819);
or U4959 (N_4959,N_4858,N_4887);
xnor U4960 (N_4960,N_4824,N_4822);
and U4961 (N_4961,N_4843,N_4852);
nand U4962 (N_4962,N_4860,N_4809);
and U4963 (N_4963,N_4865,N_4831);
xor U4964 (N_4964,N_4803,N_4845);
xnor U4965 (N_4965,N_4847,N_4801);
nor U4966 (N_4966,N_4853,N_4800);
nor U4967 (N_4967,N_4874,N_4896);
or U4968 (N_4968,N_4838,N_4876);
and U4969 (N_4969,N_4843,N_4848);
xor U4970 (N_4970,N_4817,N_4849);
xor U4971 (N_4971,N_4822,N_4804);
xor U4972 (N_4972,N_4842,N_4800);
nand U4973 (N_4973,N_4805,N_4830);
or U4974 (N_4974,N_4853,N_4870);
or U4975 (N_4975,N_4860,N_4827);
nor U4976 (N_4976,N_4832,N_4889);
or U4977 (N_4977,N_4825,N_4831);
nand U4978 (N_4978,N_4847,N_4806);
nor U4979 (N_4979,N_4852,N_4868);
nor U4980 (N_4980,N_4892,N_4858);
nand U4981 (N_4981,N_4884,N_4836);
nand U4982 (N_4982,N_4835,N_4833);
nand U4983 (N_4983,N_4870,N_4875);
xor U4984 (N_4984,N_4852,N_4829);
or U4985 (N_4985,N_4861,N_4833);
nor U4986 (N_4986,N_4887,N_4876);
xor U4987 (N_4987,N_4893,N_4870);
xor U4988 (N_4988,N_4867,N_4845);
nor U4989 (N_4989,N_4812,N_4802);
or U4990 (N_4990,N_4825,N_4870);
xor U4991 (N_4991,N_4811,N_4881);
and U4992 (N_4992,N_4832,N_4883);
nor U4993 (N_4993,N_4842,N_4851);
xor U4994 (N_4994,N_4837,N_4857);
nor U4995 (N_4995,N_4820,N_4897);
nand U4996 (N_4996,N_4808,N_4828);
nand U4997 (N_4997,N_4811,N_4866);
nor U4998 (N_4998,N_4884,N_4880);
or U4999 (N_4999,N_4880,N_4849);
and UO_0 (O_0,N_4907,N_4917);
nand UO_1 (O_1,N_4989,N_4938);
or UO_2 (O_2,N_4957,N_4979);
nor UO_3 (O_3,N_4974,N_4918);
xnor UO_4 (O_4,N_4995,N_4975);
nand UO_5 (O_5,N_4943,N_4992);
nor UO_6 (O_6,N_4971,N_4984);
xor UO_7 (O_7,N_4961,N_4988);
xnor UO_8 (O_8,N_4922,N_4948);
and UO_9 (O_9,N_4967,N_4919);
and UO_10 (O_10,N_4966,N_4930);
and UO_11 (O_11,N_4977,N_4923);
or UO_12 (O_12,N_4900,N_4913);
and UO_13 (O_13,N_4910,N_4991);
xor UO_14 (O_14,N_4973,N_4963);
xnor UO_15 (O_15,N_4920,N_4903);
nor UO_16 (O_16,N_4928,N_4987);
nand UO_17 (O_17,N_4906,N_4924);
or UO_18 (O_18,N_4914,N_4908);
or UO_19 (O_19,N_4932,N_4921);
nor UO_20 (O_20,N_4901,N_4981);
xnor UO_21 (O_21,N_4999,N_4986);
nor UO_22 (O_22,N_4952,N_4965);
xnor UO_23 (O_23,N_4985,N_4941);
xnor UO_24 (O_24,N_4994,N_4997);
xor UO_25 (O_25,N_4946,N_4970);
xor UO_26 (O_26,N_4935,N_4976);
or UO_27 (O_27,N_4990,N_4936);
or UO_28 (O_28,N_4912,N_4944);
nor UO_29 (O_29,N_4951,N_4939);
nand UO_30 (O_30,N_4955,N_4933);
or UO_31 (O_31,N_4956,N_4940);
nand UO_32 (O_32,N_4998,N_4926);
xnor UO_33 (O_33,N_4925,N_4969);
and UO_34 (O_34,N_4949,N_4959);
nand UO_35 (O_35,N_4947,N_4958);
and UO_36 (O_36,N_4945,N_4904);
and UO_37 (O_37,N_4942,N_4931);
nand UO_38 (O_38,N_4916,N_4911);
xor UO_39 (O_39,N_4902,N_4960);
nor UO_40 (O_40,N_4980,N_4953);
or UO_41 (O_41,N_4964,N_4929);
nand UO_42 (O_42,N_4909,N_4927);
or UO_43 (O_43,N_4937,N_4983);
nand UO_44 (O_44,N_4950,N_4996);
nand UO_45 (O_45,N_4978,N_4993);
nor UO_46 (O_46,N_4905,N_4962);
xor UO_47 (O_47,N_4915,N_4982);
nor UO_48 (O_48,N_4972,N_4954);
nand UO_49 (O_49,N_4968,N_4934);
nor UO_50 (O_50,N_4963,N_4929);
nor UO_51 (O_51,N_4965,N_4967);
or UO_52 (O_52,N_4957,N_4927);
nand UO_53 (O_53,N_4951,N_4986);
nand UO_54 (O_54,N_4938,N_4930);
nand UO_55 (O_55,N_4958,N_4985);
xor UO_56 (O_56,N_4976,N_4983);
nor UO_57 (O_57,N_4915,N_4910);
or UO_58 (O_58,N_4920,N_4990);
and UO_59 (O_59,N_4976,N_4907);
and UO_60 (O_60,N_4916,N_4998);
xor UO_61 (O_61,N_4929,N_4957);
nand UO_62 (O_62,N_4949,N_4922);
xor UO_63 (O_63,N_4975,N_4932);
nand UO_64 (O_64,N_4966,N_4919);
or UO_65 (O_65,N_4906,N_4989);
or UO_66 (O_66,N_4952,N_4988);
nand UO_67 (O_67,N_4993,N_4942);
xnor UO_68 (O_68,N_4932,N_4947);
nand UO_69 (O_69,N_4985,N_4953);
or UO_70 (O_70,N_4984,N_4912);
xor UO_71 (O_71,N_4971,N_4926);
nand UO_72 (O_72,N_4945,N_4946);
and UO_73 (O_73,N_4999,N_4966);
and UO_74 (O_74,N_4962,N_4966);
and UO_75 (O_75,N_4992,N_4980);
or UO_76 (O_76,N_4920,N_4952);
and UO_77 (O_77,N_4973,N_4918);
and UO_78 (O_78,N_4915,N_4983);
or UO_79 (O_79,N_4901,N_4999);
nor UO_80 (O_80,N_4989,N_4990);
nand UO_81 (O_81,N_4982,N_4922);
nor UO_82 (O_82,N_4965,N_4904);
nand UO_83 (O_83,N_4991,N_4923);
nand UO_84 (O_84,N_4964,N_4915);
nor UO_85 (O_85,N_4947,N_4981);
or UO_86 (O_86,N_4976,N_4932);
nor UO_87 (O_87,N_4919,N_4972);
and UO_88 (O_88,N_4924,N_4903);
and UO_89 (O_89,N_4978,N_4934);
nor UO_90 (O_90,N_4957,N_4904);
and UO_91 (O_91,N_4999,N_4989);
nor UO_92 (O_92,N_4988,N_4971);
nor UO_93 (O_93,N_4955,N_4999);
and UO_94 (O_94,N_4997,N_4925);
nand UO_95 (O_95,N_4996,N_4948);
xnor UO_96 (O_96,N_4980,N_4935);
nand UO_97 (O_97,N_4955,N_4927);
xnor UO_98 (O_98,N_4990,N_4921);
xnor UO_99 (O_99,N_4935,N_4987);
and UO_100 (O_100,N_4991,N_4924);
nand UO_101 (O_101,N_4900,N_4914);
nor UO_102 (O_102,N_4966,N_4950);
xor UO_103 (O_103,N_4930,N_4980);
xnor UO_104 (O_104,N_4949,N_4992);
nor UO_105 (O_105,N_4910,N_4946);
and UO_106 (O_106,N_4979,N_4960);
nand UO_107 (O_107,N_4904,N_4961);
and UO_108 (O_108,N_4980,N_4919);
nor UO_109 (O_109,N_4957,N_4975);
xnor UO_110 (O_110,N_4922,N_4967);
or UO_111 (O_111,N_4975,N_4983);
nand UO_112 (O_112,N_4957,N_4949);
or UO_113 (O_113,N_4941,N_4909);
nand UO_114 (O_114,N_4931,N_4925);
nor UO_115 (O_115,N_4985,N_4986);
and UO_116 (O_116,N_4943,N_4928);
nand UO_117 (O_117,N_4984,N_4904);
and UO_118 (O_118,N_4949,N_4921);
xor UO_119 (O_119,N_4945,N_4908);
xnor UO_120 (O_120,N_4924,N_4922);
nand UO_121 (O_121,N_4975,N_4922);
xor UO_122 (O_122,N_4941,N_4934);
nor UO_123 (O_123,N_4919,N_4903);
xnor UO_124 (O_124,N_4914,N_4930);
or UO_125 (O_125,N_4911,N_4956);
and UO_126 (O_126,N_4912,N_4953);
nor UO_127 (O_127,N_4931,N_4991);
xor UO_128 (O_128,N_4984,N_4972);
and UO_129 (O_129,N_4913,N_4966);
xnor UO_130 (O_130,N_4983,N_4968);
nand UO_131 (O_131,N_4969,N_4914);
or UO_132 (O_132,N_4945,N_4988);
or UO_133 (O_133,N_4918,N_4995);
xor UO_134 (O_134,N_4961,N_4912);
and UO_135 (O_135,N_4981,N_4970);
xnor UO_136 (O_136,N_4981,N_4935);
or UO_137 (O_137,N_4915,N_4981);
nand UO_138 (O_138,N_4923,N_4934);
nand UO_139 (O_139,N_4904,N_4947);
nand UO_140 (O_140,N_4902,N_4938);
or UO_141 (O_141,N_4908,N_4962);
nor UO_142 (O_142,N_4926,N_4960);
nand UO_143 (O_143,N_4961,N_4986);
xnor UO_144 (O_144,N_4917,N_4962);
and UO_145 (O_145,N_4958,N_4957);
nand UO_146 (O_146,N_4931,N_4977);
nand UO_147 (O_147,N_4914,N_4918);
nand UO_148 (O_148,N_4915,N_4951);
and UO_149 (O_149,N_4982,N_4950);
nand UO_150 (O_150,N_4950,N_4975);
nand UO_151 (O_151,N_4965,N_4936);
and UO_152 (O_152,N_4931,N_4967);
or UO_153 (O_153,N_4909,N_4925);
nand UO_154 (O_154,N_4919,N_4994);
and UO_155 (O_155,N_4984,N_4915);
xnor UO_156 (O_156,N_4916,N_4913);
nand UO_157 (O_157,N_4986,N_4910);
and UO_158 (O_158,N_4921,N_4991);
or UO_159 (O_159,N_4923,N_4907);
and UO_160 (O_160,N_4973,N_4972);
nor UO_161 (O_161,N_4935,N_4999);
nor UO_162 (O_162,N_4919,N_4974);
nor UO_163 (O_163,N_4908,N_4913);
or UO_164 (O_164,N_4962,N_4980);
nor UO_165 (O_165,N_4931,N_4970);
and UO_166 (O_166,N_4920,N_4940);
nor UO_167 (O_167,N_4948,N_4981);
xor UO_168 (O_168,N_4968,N_4931);
nor UO_169 (O_169,N_4951,N_4911);
xnor UO_170 (O_170,N_4978,N_4919);
xnor UO_171 (O_171,N_4931,N_4957);
and UO_172 (O_172,N_4947,N_4927);
or UO_173 (O_173,N_4915,N_4978);
or UO_174 (O_174,N_4911,N_4972);
xnor UO_175 (O_175,N_4992,N_4977);
nor UO_176 (O_176,N_4989,N_4982);
nor UO_177 (O_177,N_4922,N_4904);
nor UO_178 (O_178,N_4968,N_4989);
xor UO_179 (O_179,N_4954,N_4941);
nand UO_180 (O_180,N_4940,N_4951);
and UO_181 (O_181,N_4908,N_4900);
xor UO_182 (O_182,N_4906,N_4973);
xnor UO_183 (O_183,N_4908,N_4932);
and UO_184 (O_184,N_4948,N_4906);
or UO_185 (O_185,N_4920,N_4971);
xnor UO_186 (O_186,N_4902,N_4904);
nand UO_187 (O_187,N_4996,N_4940);
nand UO_188 (O_188,N_4926,N_4964);
nor UO_189 (O_189,N_4901,N_4937);
nand UO_190 (O_190,N_4906,N_4964);
nor UO_191 (O_191,N_4953,N_4964);
or UO_192 (O_192,N_4940,N_4974);
nor UO_193 (O_193,N_4913,N_4934);
nor UO_194 (O_194,N_4900,N_4973);
nand UO_195 (O_195,N_4909,N_4987);
xor UO_196 (O_196,N_4919,N_4924);
and UO_197 (O_197,N_4962,N_4914);
and UO_198 (O_198,N_4915,N_4959);
or UO_199 (O_199,N_4913,N_4939);
or UO_200 (O_200,N_4964,N_4902);
nor UO_201 (O_201,N_4966,N_4973);
xor UO_202 (O_202,N_4967,N_4937);
nand UO_203 (O_203,N_4926,N_4992);
nand UO_204 (O_204,N_4935,N_4979);
nor UO_205 (O_205,N_4915,N_4973);
and UO_206 (O_206,N_4973,N_4976);
xor UO_207 (O_207,N_4988,N_4922);
or UO_208 (O_208,N_4904,N_4920);
xor UO_209 (O_209,N_4928,N_4929);
nor UO_210 (O_210,N_4905,N_4913);
nor UO_211 (O_211,N_4962,N_4919);
nand UO_212 (O_212,N_4994,N_4905);
nand UO_213 (O_213,N_4939,N_4966);
nand UO_214 (O_214,N_4924,N_4987);
nor UO_215 (O_215,N_4901,N_4942);
nor UO_216 (O_216,N_4953,N_4906);
nand UO_217 (O_217,N_4998,N_4913);
and UO_218 (O_218,N_4990,N_4966);
or UO_219 (O_219,N_4903,N_4911);
and UO_220 (O_220,N_4907,N_4912);
or UO_221 (O_221,N_4987,N_4950);
and UO_222 (O_222,N_4912,N_4914);
and UO_223 (O_223,N_4990,N_4993);
nor UO_224 (O_224,N_4919,N_4986);
and UO_225 (O_225,N_4981,N_4900);
nand UO_226 (O_226,N_4900,N_4994);
or UO_227 (O_227,N_4901,N_4923);
and UO_228 (O_228,N_4907,N_4966);
nor UO_229 (O_229,N_4964,N_4996);
or UO_230 (O_230,N_4901,N_4972);
or UO_231 (O_231,N_4978,N_4961);
or UO_232 (O_232,N_4930,N_4917);
nand UO_233 (O_233,N_4972,N_4912);
nor UO_234 (O_234,N_4965,N_4919);
xor UO_235 (O_235,N_4959,N_4916);
and UO_236 (O_236,N_4914,N_4949);
or UO_237 (O_237,N_4975,N_4920);
and UO_238 (O_238,N_4945,N_4900);
nand UO_239 (O_239,N_4948,N_4974);
nor UO_240 (O_240,N_4955,N_4973);
nand UO_241 (O_241,N_4953,N_4999);
and UO_242 (O_242,N_4941,N_4924);
and UO_243 (O_243,N_4982,N_4966);
or UO_244 (O_244,N_4924,N_4960);
and UO_245 (O_245,N_4956,N_4948);
nand UO_246 (O_246,N_4951,N_4977);
or UO_247 (O_247,N_4916,N_4955);
xor UO_248 (O_248,N_4908,N_4930);
nand UO_249 (O_249,N_4958,N_4979);
and UO_250 (O_250,N_4942,N_4969);
xnor UO_251 (O_251,N_4935,N_4940);
nor UO_252 (O_252,N_4958,N_4934);
nand UO_253 (O_253,N_4928,N_4918);
or UO_254 (O_254,N_4958,N_4900);
or UO_255 (O_255,N_4946,N_4999);
xnor UO_256 (O_256,N_4914,N_4973);
nor UO_257 (O_257,N_4929,N_4981);
nand UO_258 (O_258,N_4967,N_4995);
nand UO_259 (O_259,N_4979,N_4923);
and UO_260 (O_260,N_4957,N_4948);
nand UO_261 (O_261,N_4915,N_4942);
xnor UO_262 (O_262,N_4988,N_4949);
or UO_263 (O_263,N_4992,N_4914);
nand UO_264 (O_264,N_4975,N_4939);
xnor UO_265 (O_265,N_4933,N_4980);
or UO_266 (O_266,N_4968,N_4922);
nand UO_267 (O_267,N_4937,N_4924);
and UO_268 (O_268,N_4987,N_4915);
xnor UO_269 (O_269,N_4930,N_4945);
and UO_270 (O_270,N_4942,N_4972);
xor UO_271 (O_271,N_4972,N_4933);
nand UO_272 (O_272,N_4951,N_4950);
nand UO_273 (O_273,N_4944,N_4999);
nand UO_274 (O_274,N_4938,N_4914);
nor UO_275 (O_275,N_4963,N_4931);
and UO_276 (O_276,N_4918,N_4930);
and UO_277 (O_277,N_4963,N_4978);
and UO_278 (O_278,N_4922,N_4921);
or UO_279 (O_279,N_4938,N_4910);
nand UO_280 (O_280,N_4934,N_4925);
nand UO_281 (O_281,N_4937,N_4935);
nor UO_282 (O_282,N_4960,N_4980);
xor UO_283 (O_283,N_4977,N_4995);
or UO_284 (O_284,N_4948,N_4913);
nor UO_285 (O_285,N_4983,N_4922);
and UO_286 (O_286,N_4922,N_4918);
or UO_287 (O_287,N_4974,N_4902);
nand UO_288 (O_288,N_4926,N_4974);
nor UO_289 (O_289,N_4963,N_4928);
nor UO_290 (O_290,N_4931,N_4975);
xor UO_291 (O_291,N_4921,N_4965);
or UO_292 (O_292,N_4986,N_4913);
xnor UO_293 (O_293,N_4995,N_4998);
nor UO_294 (O_294,N_4982,N_4975);
xnor UO_295 (O_295,N_4948,N_4937);
and UO_296 (O_296,N_4958,N_4949);
and UO_297 (O_297,N_4937,N_4959);
and UO_298 (O_298,N_4949,N_4967);
or UO_299 (O_299,N_4953,N_4955);
and UO_300 (O_300,N_4907,N_4927);
nand UO_301 (O_301,N_4998,N_4955);
xnor UO_302 (O_302,N_4946,N_4995);
and UO_303 (O_303,N_4962,N_4901);
nand UO_304 (O_304,N_4902,N_4958);
and UO_305 (O_305,N_4988,N_4986);
xor UO_306 (O_306,N_4966,N_4924);
nand UO_307 (O_307,N_4901,N_4963);
nor UO_308 (O_308,N_4924,N_4930);
nor UO_309 (O_309,N_4990,N_4994);
nand UO_310 (O_310,N_4987,N_4911);
or UO_311 (O_311,N_4943,N_4914);
xnor UO_312 (O_312,N_4927,N_4992);
and UO_313 (O_313,N_4944,N_4907);
nand UO_314 (O_314,N_4951,N_4902);
xnor UO_315 (O_315,N_4972,N_4925);
or UO_316 (O_316,N_4992,N_4915);
and UO_317 (O_317,N_4988,N_4977);
or UO_318 (O_318,N_4949,N_4916);
nand UO_319 (O_319,N_4951,N_4925);
or UO_320 (O_320,N_4909,N_4993);
or UO_321 (O_321,N_4973,N_4964);
or UO_322 (O_322,N_4958,N_4905);
and UO_323 (O_323,N_4925,N_4968);
and UO_324 (O_324,N_4958,N_4992);
and UO_325 (O_325,N_4926,N_4945);
or UO_326 (O_326,N_4925,N_4905);
nor UO_327 (O_327,N_4916,N_4961);
or UO_328 (O_328,N_4924,N_4913);
and UO_329 (O_329,N_4986,N_4940);
nor UO_330 (O_330,N_4966,N_4952);
nor UO_331 (O_331,N_4929,N_4942);
nand UO_332 (O_332,N_4906,N_4961);
or UO_333 (O_333,N_4981,N_4932);
and UO_334 (O_334,N_4901,N_4950);
and UO_335 (O_335,N_4989,N_4965);
nand UO_336 (O_336,N_4954,N_4969);
and UO_337 (O_337,N_4928,N_4952);
nor UO_338 (O_338,N_4906,N_4922);
and UO_339 (O_339,N_4904,N_4962);
nor UO_340 (O_340,N_4967,N_4961);
or UO_341 (O_341,N_4927,N_4921);
and UO_342 (O_342,N_4998,N_4942);
and UO_343 (O_343,N_4931,N_4989);
nand UO_344 (O_344,N_4995,N_4996);
and UO_345 (O_345,N_4932,N_4900);
and UO_346 (O_346,N_4993,N_4947);
nor UO_347 (O_347,N_4905,N_4967);
and UO_348 (O_348,N_4927,N_4914);
and UO_349 (O_349,N_4949,N_4938);
or UO_350 (O_350,N_4936,N_4939);
xor UO_351 (O_351,N_4995,N_4974);
and UO_352 (O_352,N_4916,N_4968);
nor UO_353 (O_353,N_4907,N_4942);
xnor UO_354 (O_354,N_4975,N_4916);
nand UO_355 (O_355,N_4937,N_4956);
nand UO_356 (O_356,N_4924,N_4929);
and UO_357 (O_357,N_4904,N_4907);
nor UO_358 (O_358,N_4904,N_4935);
and UO_359 (O_359,N_4925,N_4989);
nand UO_360 (O_360,N_4995,N_4900);
nor UO_361 (O_361,N_4998,N_4966);
or UO_362 (O_362,N_4980,N_4977);
or UO_363 (O_363,N_4953,N_4919);
nor UO_364 (O_364,N_4931,N_4918);
xor UO_365 (O_365,N_4947,N_4900);
nand UO_366 (O_366,N_4970,N_4953);
xnor UO_367 (O_367,N_4944,N_4909);
or UO_368 (O_368,N_4996,N_4986);
nor UO_369 (O_369,N_4940,N_4909);
and UO_370 (O_370,N_4974,N_4956);
and UO_371 (O_371,N_4976,N_4999);
and UO_372 (O_372,N_4911,N_4929);
nand UO_373 (O_373,N_4965,N_4910);
nor UO_374 (O_374,N_4975,N_4917);
or UO_375 (O_375,N_4909,N_4992);
xnor UO_376 (O_376,N_4915,N_4995);
nand UO_377 (O_377,N_4904,N_4964);
xnor UO_378 (O_378,N_4944,N_4916);
xor UO_379 (O_379,N_4957,N_4995);
and UO_380 (O_380,N_4931,N_4956);
nor UO_381 (O_381,N_4982,N_4916);
xnor UO_382 (O_382,N_4927,N_4912);
or UO_383 (O_383,N_4986,N_4962);
nor UO_384 (O_384,N_4988,N_4981);
nor UO_385 (O_385,N_4917,N_4974);
nor UO_386 (O_386,N_4917,N_4992);
xor UO_387 (O_387,N_4974,N_4905);
nand UO_388 (O_388,N_4989,N_4934);
or UO_389 (O_389,N_4932,N_4986);
nor UO_390 (O_390,N_4921,N_4924);
nor UO_391 (O_391,N_4991,N_4950);
xor UO_392 (O_392,N_4951,N_4944);
or UO_393 (O_393,N_4982,N_4952);
xor UO_394 (O_394,N_4973,N_4962);
nor UO_395 (O_395,N_4995,N_4958);
nand UO_396 (O_396,N_4978,N_4937);
xnor UO_397 (O_397,N_4996,N_4987);
and UO_398 (O_398,N_4936,N_4988);
and UO_399 (O_399,N_4924,N_4952);
nor UO_400 (O_400,N_4900,N_4910);
nor UO_401 (O_401,N_4910,N_4905);
xnor UO_402 (O_402,N_4971,N_4927);
or UO_403 (O_403,N_4965,N_4962);
nor UO_404 (O_404,N_4957,N_4988);
or UO_405 (O_405,N_4973,N_4952);
and UO_406 (O_406,N_4970,N_4979);
or UO_407 (O_407,N_4983,N_4989);
or UO_408 (O_408,N_4920,N_4989);
and UO_409 (O_409,N_4931,N_4927);
or UO_410 (O_410,N_4941,N_4914);
and UO_411 (O_411,N_4935,N_4920);
xor UO_412 (O_412,N_4985,N_4979);
or UO_413 (O_413,N_4957,N_4959);
nor UO_414 (O_414,N_4931,N_4952);
xor UO_415 (O_415,N_4961,N_4937);
nor UO_416 (O_416,N_4923,N_4935);
and UO_417 (O_417,N_4960,N_4927);
nand UO_418 (O_418,N_4939,N_4935);
xnor UO_419 (O_419,N_4932,N_4901);
nor UO_420 (O_420,N_4976,N_4954);
xnor UO_421 (O_421,N_4947,N_4984);
nor UO_422 (O_422,N_4988,N_4925);
nand UO_423 (O_423,N_4965,N_4948);
or UO_424 (O_424,N_4997,N_4948);
and UO_425 (O_425,N_4997,N_4981);
and UO_426 (O_426,N_4972,N_4928);
nor UO_427 (O_427,N_4993,N_4917);
nor UO_428 (O_428,N_4939,N_4908);
nor UO_429 (O_429,N_4977,N_4985);
and UO_430 (O_430,N_4967,N_4975);
and UO_431 (O_431,N_4954,N_4930);
xor UO_432 (O_432,N_4963,N_4940);
xor UO_433 (O_433,N_4912,N_4911);
and UO_434 (O_434,N_4932,N_4909);
and UO_435 (O_435,N_4914,N_4942);
and UO_436 (O_436,N_4986,N_4903);
or UO_437 (O_437,N_4912,N_4977);
nor UO_438 (O_438,N_4960,N_4978);
xor UO_439 (O_439,N_4936,N_4999);
xor UO_440 (O_440,N_4954,N_4902);
nand UO_441 (O_441,N_4900,N_4983);
nand UO_442 (O_442,N_4953,N_4922);
nand UO_443 (O_443,N_4937,N_4990);
or UO_444 (O_444,N_4990,N_4982);
xnor UO_445 (O_445,N_4966,N_4960);
nand UO_446 (O_446,N_4923,N_4914);
xnor UO_447 (O_447,N_4926,N_4928);
nor UO_448 (O_448,N_4965,N_4925);
and UO_449 (O_449,N_4929,N_4933);
or UO_450 (O_450,N_4904,N_4968);
nand UO_451 (O_451,N_4935,N_4996);
and UO_452 (O_452,N_4954,N_4992);
or UO_453 (O_453,N_4914,N_4944);
xnor UO_454 (O_454,N_4920,N_4900);
nand UO_455 (O_455,N_4948,N_4966);
nand UO_456 (O_456,N_4924,N_4984);
nor UO_457 (O_457,N_4976,N_4977);
xor UO_458 (O_458,N_4911,N_4908);
or UO_459 (O_459,N_4936,N_4935);
nand UO_460 (O_460,N_4949,N_4999);
and UO_461 (O_461,N_4917,N_4998);
nor UO_462 (O_462,N_4923,N_4944);
nand UO_463 (O_463,N_4951,N_4994);
nand UO_464 (O_464,N_4976,N_4913);
nand UO_465 (O_465,N_4958,N_4912);
nor UO_466 (O_466,N_4903,N_4990);
nor UO_467 (O_467,N_4919,N_4945);
or UO_468 (O_468,N_4995,N_4930);
xnor UO_469 (O_469,N_4985,N_4993);
or UO_470 (O_470,N_4962,N_4935);
and UO_471 (O_471,N_4968,N_4903);
and UO_472 (O_472,N_4918,N_4985);
and UO_473 (O_473,N_4956,N_4932);
xnor UO_474 (O_474,N_4969,N_4982);
and UO_475 (O_475,N_4918,N_4950);
and UO_476 (O_476,N_4910,N_4922);
nand UO_477 (O_477,N_4978,N_4944);
nor UO_478 (O_478,N_4946,N_4900);
nand UO_479 (O_479,N_4918,N_4904);
nor UO_480 (O_480,N_4918,N_4963);
nor UO_481 (O_481,N_4932,N_4993);
xnor UO_482 (O_482,N_4934,N_4986);
xor UO_483 (O_483,N_4972,N_4921);
and UO_484 (O_484,N_4930,N_4900);
nand UO_485 (O_485,N_4922,N_4965);
nor UO_486 (O_486,N_4992,N_4902);
xor UO_487 (O_487,N_4957,N_4955);
or UO_488 (O_488,N_4943,N_4915);
or UO_489 (O_489,N_4904,N_4901);
and UO_490 (O_490,N_4919,N_4993);
nor UO_491 (O_491,N_4953,N_4929);
nor UO_492 (O_492,N_4904,N_4999);
or UO_493 (O_493,N_4988,N_4929);
nand UO_494 (O_494,N_4925,N_4936);
xor UO_495 (O_495,N_4983,N_4988);
nand UO_496 (O_496,N_4969,N_4902);
nand UO_497 (O_497,N_4976,N_4924);
nand UO_498 (O_498,N_4901,N_4987);
nor UO_499 (O_499,N_4981,N_4940);
or UO_500 (O_500,N_4937,N_4984);
nand UO_501 (O_501,N_4938,N_4970);
and UO_502 (O_502,N_4944,N_4901);
nand UO_503 (O_503,N_4967,N_4940);
xnor UO_504 (O_504,N_4983,N_4950);
or UO_505 (O_505,N_4969,N_4936);
or UO_506 (O_506,N_4913,N_4978);
xnor UO_507 (O_507,N_4935,N_4958);
xor UO_508 (O_508,N_4993,N_4927);
or UO_509 (O_509,N_4994,N_4914);
nand UO_510 (O_510,N_4992,N_4984);
and UO_511 (O_511,N_4990,N_4963);
or UO_512 (O_512,N_4960,N_4964);
nor UO_513 (O_513,N_4981,N_4975);
nor UO_514 (O_514,N_4940,N_4952);
xor UO_515 (O_515,N_4973,N_4942);
or UO_516 (O_516,N_4994,N_4928);
nand UO_517 (O_517,N_4948,N_4935);
xnor UO_518 (O_518,N_4954,N_4919);
and UO_519 (O_519,N_4909,N_4931);
nand UO_520 (O_520,N_4971,N_4932);
nor UO_521 (O_521,N_4975,N_4928);
nand UO_522 (O_522,N_4907,N_4931);
nor UO_523 (O_523,N_4954,N_4942);
xor UO_524 (O_524,N_4925,N_4901);
nor UO_525 (O_525,N_4906,N_4968);
or UO_526 (O_526,N_4985,N_4930);
or UO_527 (O_527,N_4980,N_4955);
xnor UO_528 (O_528,N_4992,N_4939);
nand UO_529 (O_529,N_4947,N_4998);
nor UO_530 (O_530,N_4912,N_4945);
xor UO_531 (O_531,N_4970,N_4937);
and UO_532 (O_532,N_4973,N_4943);
nand UO_533 (O_533,N_4969,N_4966);
xnor UO_534 (O_534,N_4952,N_4945);
nand UO_535 (O_535,N_4900,N_4915);
and UO_536 (O_536,N_4956,N_4939);
nand UO_537 (O_537,N_4963,N_4911);
nor UO_538 (O_538,N_4906,N_4913);
xnor UO_539 (O_539,N_4962,N_4927);
nand UO_540 (O_540,N_4953,N_4995);
xor UO_541 (O_541,N_4917,N_4935);
xor UO_542 (O_542,N_4934,N_4995);
and UO_543 (O_543,N_4923,N_4940);
nor UO_544 (O_544,N_4952,N_4983);
xor UO_545 (O_545,N_4925,N_4947);
or UO_546 (O_546,N_4942,N_4905);
or UO_547 (O_547,N_4939,N_4902);
nand UO_548 (O_548,N_4907,N_4980);
nor UO_549 (O_549,N_4971,N_4914);
or UO_550 (O_550,N_4937,N_4931);
xor UO_551 (O_551,N_4959,N_4964);
or UO_552 (O_552,N_4973,N_4957);
or UO_553 (O_553,N_4941,N_4937);
nand UO_554 (O_554,N_4953,N_4936);
nor UO_555 (O_555,N_4971,N_4900);
or UO_556 (O_556,N_4929,N_4956);
or UO_557 (O_557,N_4963,N_4938);
nand UO_558 (O_558,N_4965,N_4956);
and UO_559 (O_559,N_4959,N_4958);
nor UO_560 (O_560,N_4927,N_4948);
or UO_561 (O_561,N_4986,N_4989);
or UO_562 (O_562,N_4976,N_4948);
nand UO_563 (O_563,N_4980,N_4947);
or UO_564 (O_564,N_4936,N_4951);
nor UO_565 (O_565,N_4963,N_4900);
xnor UO_566 (O_566,N_4912,N_4993);
nand UO_567 (O_567,N_4951,N_4941);
or UO_568 (O_568,N_4958,N_4937);
xor UO_569 (O_569,N_4999,N_4930);
or UO_570 (O_570,N_4909,N_4915);
and UO_571 (O_571,N_4923,N_4946);
nor UO_572 (O_572,N_4962,N_4931);
nand UO_573 (O_573,N_4968,N_4990);
nor UO_574 (O_574,N_4972,N_4918);
xor UO_575 (O_575,N_4941,N_4989);
nor UO_576 (O_576,N_4945,N_4903);
and UO_577 (O_577,N_4958,N_4981);
or UO_578 (O_578,N_4945,N_4942);
nand UO_579 (O_579,N_4920,N_4955);
xor UO_580 (O_580,N_4952,N_4979);
nor UO_581 (O_581,N_4918,N_4967);
xor UO_582 (O_582,N_4949,N_4908);
and UO_583 (O_583,N_4956,N_4924);
nand UO_584 (O_584,N_4991,N_4989);
nand UO_585 (O_585,N_4904,N_4975);
nand UO_586 (O_586,N_4922,N_4996);
and UO_587 (O_587,N_4911,N_4970);
or UO_588 (O_588,N_4975,N_4903);
and UO_589 (O_589,N_4937,N_4997);
or UO_590 (O_590,N_4910,N_4902);
and UO_591 (O_591,N_4945,N_4971);
xnor UO_592 (O_592,N_4952,N_4975);
nand UO_593 (O_593,N_4997,N_4921);
nor UO_594 (O_594,N_4968,N_4966);
and UO_595 (O_595,N_4956,N_4985);
or UO_596 (O_596,N_4926,N_4953);
or UO_597 (O_597,N_4972,N_4931);
or UO_598 (O_598,N_4994,N_4956);
and UO_599 (O_599,N_4954,N_4920);
nand UO_600 (O_600,N_4918,N_4997);
xnor UO_601 (O_601,N_4989,N_4949);
xor UO_602 (O_602,N_4916,N_4900);
and UO_603 (O_603,N_4996,N_4980);
xor UO_604 (O_604,N_4929,N_4976);
or UO_605 (O_605,N_4974,N_4936);
nor UO_606 (O_606,N_4911,N_4964);
nand UO_607 (O_607,N_4946,N_4975);
and UO_608 (O_608,N_4993,N_4938);
and UO_609 (O_609,N_4992,N_4918);
nor UO_610 (O_610,N_4986,N_4933);
nand UO_611 (O_611,N_4956,N_4993);
nor UO_612 (O_612,N_4926,N_4901);
and UO_613 (O_613,N_4976,N_4982);
and UO_614 (O_614,N_4962,N_4944);
xnor UO_615 (O_615,N_4986,N_4954);
nor UO_616 (O_616,N_4945,N_4924);
xor UO_617 (O_617,N_4988,N_4963);
nand UO_618 (O_618,N_4995,N_4938);
and UO_619 (O_619,N_4900,N_4989);
or UO_620 (O_620,N_4973,N_4924);
nor UO_621 (O_621,N_4929,N_4973);
xor UO_622 (O_622,N_4940,N_4914);
or UO_623 (O_623,N_4931,N_4930);
and UO_624 (O_624,N_4909,N_4956);
or UO_625 (O_625,N_4943,N_4913);
or UO_626 (O_626,N_4932,N_4945);
nor UO_627 (O_627,N_4910,N_4941);
nand UO_628 (O_628,N_4973,N_4903);
xor UO_629 (O_629,N_4991,N_4966);
nor UO_630 (O_630,N_4988,N_4933);
and UO_631 (O_631,N_4999,N_4921);
nand UO_632 (O_632,N_4918,N_4941);
xor UO_633 (O_633,N_4971,N_4964);
xnor UO_634 (O_634,N_4981,N_4971);
xor UO_635 (O_635,N_4945,N_4986);
and UO_636 (O_636,N_4923,N_4974);
or UO_637 (O_637,N_4971,N_4911);
or UO_638 (O_638,N_4980,N_4981);
nand UO_639 (O_639,N_4902,N_4911);
and UO_640 (O_640,N_4967,N_4936);
nor UO_641 (O_641,N_4992,N_4930);
xnor UO_642 (O_642,N_4954,N_4978);
nand UO_643 (O_643,N_4922,N_4941);
xnor UO_644 (O_644,N_4987,N_4902);
nor UO_645 (O_645,N_4977,N_4952);
and UO_646 (O_646,N_4916,N_4931);
nand UO_647 (O_647,N_4999,N_4948);
and UO_648 (O_648,N_4903,N_4925);
nand UO_649 (O_649,N_4977,N_4969);
nor UO_650 (O_650,N_4935,N_4930);
and UO_651 (O_651,N_4945,N_4955);
nor UO_652 (O_652,N_4981,N_4927);
xnor UO_653 (O_653,N_4917,N_4966);
nand UO_654 (O_654,N_4935,N_4941);
nor UO_655 (O_655,N_4908,N_4961);
xnor UO_656 (O_656,N_4966,N_4996);
nor UO_657 (O_657,N_4997,N_4914);
and UO_658 (O_658,N_4996,N_4982);
nand UO_659 (O_659,N_4936,N_4966);
and UO_660 (O_660,N_4992,N_4993);
xor UO_661 (O_661,N_4941,N_4977);
and UO_662 (O_662,N_4931,N_4969);
nand UO_663 (O_663,N_4925,N_4996);
nor UO_664 (O_664,N_4958,N_4954);
or UO_665 (O_665,N_4923,N_4931);
and UO_666 (O_666,N_4923,N_4915);
nor UO_667 (O_667,N_4928,N_4944);
nand UO_668 (O_668,N_4965,N_4926);
nand UO_669 (O_669,N_4901,N_4927);
nand UO_670 (O_670,N_4937,N_4954);
xnor UO_671 (O_671,N_4993,N_4984);
xor UO_672 (O_672,N_4933,N_4906);
nor UO_673 (O_673,N_4916,N_4951);
and UO_674 (O_674,N_4926,N_4994);
and UO_675 (O_675,N_4923,N_4951);
nor UO_676 (O_676,N_4960,N_4945);
nor UO_677 (O_677,N_4989,N_4996);
and UO_678 (O_678,N_4995,N_4952);
and UO_679 (O_679,N_4959,N_4987);
nor UO_680 (O_680,N_4937,N_4942);
and UO_681 (O_681,N_4936,N_4957);
nand UO_682 (O_682,N_4971,N_4948);
nor UO_683 (O_683,N_4944,N_4983);
nand UO_684 (O_684,N_4916,N_4954);
or UO_685 (O_685,N_4918,N_4905);
and UO_686 (O_686,N_4943,N_4920);
or UO_687 (O_687,N_4956,N_4997);
nand UO_688 (O_688,N_4906,N_4939);
nand UO_689 (O_689,N_4941,N_4998);
nor UO_690 (O_690,N_4933,N_4935);
xnor UO_691 (O_691,N_4991,N_4917);
xor UO_692 (O_692,N_4933,N_4999);
nand UO_693 (O_693,N_4991,N_4981);
nand UO_694 (O_694,N_4951,N_4988);
xnor UO_695 (O_695,N_4982,N_4913);
nand UO_696 (O_696,N_4947,N_4955);
nor UO_697 (O_697,N_4958,N_4996);
or UO_698 (O_698,N_4977,N_4935);
nor UO_699 (O_699,N_4981,N_4979);
and UO_700 (O_700,N_4910,N_4945);
xor UO_701 (O_701,N_4916,N_4981);
xor UO_702 (O_702,N_4980,N_4926);
nand UO_703 (O_703,N_4933,N_4949);
or UO_704 (O_704,N_4903,N_4917);
nand UO_705 (O_705,N_4915,N_4994);
and UO_706 (O_706,N_4964,N_4925);
nor UO_707 (O_707,N_4963,N_4955);
nand UO_708 (O_708,N_4967,N_4935);
nor UO_709 (O_709,N_4968,N_4911);
nand UO_710 (O_710,N_4943,N_4958);
nor UO_711 (O_711,N_4988,N_4970);
nand UO_712 (O_712,N_4948,N_4998);
nor UO_713 (O_713,N_4934,N_4964);
and UO_714 (O_714,N_4931,N_4911);
xnor UO_715 (O_715,N_4959,N_4984);
nor UO_716 (O_716,N_4924,N_4909);
or UO_717 (O_717,N_4983,N_4959);
nor UO_718 (O_718,N_4923,N_4900);
xor UO_719 (O_719,N_4995,N_4987);
nor UO_720 (O_720,N_4941,N_4923);
or UO_721 (O_721,N_4913,N_4985);
nor UO_722 (O_722,N_4986,N_4979);
or UO_723 (O_723,N_4933,N_4961);
and UO_724 (O_724,N_4917,N_4910);
nand UO_725 (O_725,N_4944,N_4904);
nor UO_726 (O_726,N_4901,N_4977);
and UO_727 (O_727,N_4985,N_4900);
nand UO_728 (O_728,N_4905,N_4914);
or UO_729 (O_729,N_4974,N_4966);
nor UO_730 (O_730,N_4989,N_4950);
or UO_731 (O_731,N_4961,N_4934);
xnor UO_732 (O_732,N_4987,N_4964);
nor UO_733 (O_733,N_4950,N_4908);
xor UO_734 (O_734,N_4905,N_4930);
and UO_735 (O_735,N_4958,N_4946);
or UO_736 (O_736,N_4972,N_4937);
and UO_737 (O_737,N_4988,N_4948);
nor UO_738 (O_738,N_4985,N_4945);
nand UO_739 (O_739,N_4941,N_4903);
nand UO_740 (O_740,N_4927,N_4920);
xor UO_741 (O_741,N_4939,N_4960);
nor UO_742 (O_742,N_4990,N_4967);
nand UO_743 (O_743,N_4915,N_4966);
nor UO_744 (O_744,N_4985,N_4950);
or UO_745 (O_745,N_4986,N_4950);
nand UO_746 (O_746,N_4932,N_4997);
nor UO_747 (O_747,N_4933,N_4912);
nor UO_748 (O_748,N_4969,N_4934);
or UO_749 (O_749,N_4988,N_4984);
xnor UO_750 (O_750,N_4997,N_4922);
or UO_751 (O_751,N_4929,N_4934);
and UO_752 (O_752,N_4909,N_4950);
nand UO_753 (O_753,N_4955,N_4986);
and UO_754 (O_754,N_4907,N_4991);
nand UO_755 (O_755,N_4950,N_4926);
nand UO_756 (O_756,N_4995,N_4947);
nor UO_757 (O_757,N_4935,N_4968);
nor UO_758 (O_758,N_4908,N_4969);
nand UO_759 (O_759,N_4955,N_4942);
nand UO_760 (O_760,N_4956,N_4984);
nand UO_761 (O_761,N_4974,N_4927);
nor UO_762 (O_762,N_4905,N_4988);
nor UO_763 (O_763,N_4956,N_4959);
xor UO_764 (O_764,N_4973,N_4938);
or UO_765 (O_765,N_4979,N_4971);
nand UO_766 (O_766,N_4958,N_4975);
nor UO_767 (O_767,N_4936,N_4955);
and UO_768 (O_768,N_4956,N_4964);
xor UO_769 (O_769,N_4974,N_4958);
and UO_770 (O_770,N_4958,N_4910);
nor UO_771 (O_771,N_4918,N_4913);
xnor UO_772 (O_772,N_4945,N_4966);
nor UO_773 (O_773,N_4975,N_4979);
nand UO_774 (O_774,N_4957,N_4952);
or UO_775 (O_775,N_4943,N_4976);
xor UO_776 (O_776,N_4967,N_4903);
xor UO_777 (O_777,N_4992,N_4935);
nor UO_778 (O_778,N_4933,N_4907);
and UO_779 (O_779,N_4910,N_4962);
xor UO_780 (O_780,N_4984,N_4926);
nand UO_781 (O_781,N_4988,N_4926);
xor UO_782 (O_782,N_4971,N_4939);
nor UO_783 (O_783,N_4925,N_4977);
or UO_784 (O_784,N_4909,N_4985);
and UO_785 (O_785,N_4914,N_4910);
xnor UO_786 (O_786,N_4945,N_4958);
or UO_787 (O_787,N_4951,N_4918);
or UO_788 (O_788,N_4970,N_4978);
xor UO_789 (O_789,N_4947,N_4905);
xnor UO_790 (O_790,N_4921,N_4946);
nand UO_791 (O_791,N_4942,N_4987);
xnor UO_792 (O_792,N_4937,N_4911);
nand UO_793 (O_793,N_4945,N_4906);
or UO_794 (O_794,N_4970,N_4960);
nor UO_795 (O_795,N_4986,N_4915);
or UO_796 (O_796,N_4963,N_4982);
or UO_797 (O_797,N_4933,N_4953);
nor UO_798 (O_798,N_4932,N_4950);
nor UO_799 (O_799,N_4986,N_4998);
nand UO_800 (O_800,N_4916,N_4953);
and UO_801 (O_801,N_4954,N_4948);
or UO_802 (O_802,N_4964,N_4945);
and UO_803 (O_803,N_4922,N_4999);
nand UO_804 (O_804,N_4915,N_4920);
nor UO_805 (O_805,N_4972,N_4908);
nand UO_806 (O_806,N_4928,N_4932);
xor UO_807 (O_807,N_4924,N_4989);
nor UO_808 (O_808,N_4984,N_4952);
or UO_809 (O_809,N_4930,N_4946);
or UO_810 (O_810,N_4939,N_4930);
or UO_811 (O_811,N_4916,N_4923);
or UO_812 (O_812,N_4977,N_4944);
nand UO_813 (O_813,N_4909,N_4935);
or UO_814 (O_814,N_4926,N_4997);
xor UO_815 (O_815,N_4919,N_4937);
and UO_816 (O_816,N_4903,N_4909);
nor UO_817 (O_817,N_4999,N_4902);
xnor UO_818 (O_818,N_4945,N_4941);
or UO_819 (O_819,N_4942,N_4966);
nand UO_820 (O_820,N_4947,N_4930);
nand UO_821 (O_821,N_4927,N_4963);
nand UO_822 (O_822,N_4905,N_4961);
nand UO_823 (O_823,N_4944,N_4945);
and UO_824 (O_824,N_4988,N_4968);
and UO_825 (O_825,N_4962,N_4909);
and UO_826 (O_826,N_4931,N_4974);
and UO_827 (O_827,N_4906,N_4936);
and UO_828 (O_828,N_4921,N_4962);
nor UO_829 (O_829,N_4955,N_4994);
nor UO_830 (O_830,N_4957,N_4944);
and UO_831 (O_831,N_4933,N_4971);
xnor UO_832 (O_832,N_4980,N_4987);
xnor UO_833 (O_833,N_4989,N_4979);
nor UO_834 (O_834,N_4986,N_4908);
nand UO_835 (O_835,N_4967,N_4978);
nand UO_836 (O_836,N_4971,N_4930);
nand UO_837 (O_837,N_4977,N_4942);
nand UO_838 (O_838,N_4947,N_4902);
nand UO_839 (O_839,N_4911,N_4981);
xor UO_840 (O_840,N_4970,N_4903);
or UO_841 (O_841,N_4937,N_4940);
and UO_842 (O_842,N_4987,N_4933);
nand UO_843 (O_843,N_4974,N_4997);
nor UO_844 (O_844,N_4929,N_4989);
or UO_845 (O_845,N_4996,N_4930);
or UO_846 (O_846,N_4975,N_4960);
xnor UO_847 (O_847,N_4931,N_4933);
or UO_848 (O_848,N_4998,N_4945);
xnor UO_849 (O_849,N_4998,N_4956);
nand UO_850 (O_850,N_4991,N_4941);
nand UO_851 (O_851,N_4977,N_4959);
nor UO_852 (O_852,N_4936,N_4973);
nor UO_853 (O_853,N_4917,N_4982);
or UO_854 (O_854,N_4942,N_4983);
and UO_855 (O_855,N_4911,N_4942);
or UO_856 (O_856,N_4998,N_4912);
and UO_857 (O_857,N_4948,N_4915);
nand UO_858 (O_858,N_4928,N_4938);
nor UO_859 (O_859,N_4993,N_4988);
nor UO_860 (O_860,N_4970,N_4962);
and UO_861 (O_861,N_4997,N_4917);
nand UO_862 (O_862,N_4949,N_4976);
xor UO_863 (O_863,N_4946,N_4942);
nor UO_864 (O_864,N_4947,N_4907);
nor UO_865 (O_865,N_4926,N_4918);
nor UO_866 (O_866,N_4935,N_4995);
nand UO_867 (O_867,N_4933,N_4928);
xnor UO_868 (O_868,N_4906,N_4949);
and UO_869 (O_869,N_4921,N_4984);
xnor UO_870 (O_870,N_4947,N_4944);
nor UO_871 (O_871,N_4954,N_4906);
nor UO_872 (O_872,N_4957,N_4918);
and UO_873 (O_873,N_4974,N_4934);
xor UO_874 (O_874,N_4990,N_4957);
and UO_875 (O_875,N_4928,N_4922);
nand UO_876 (O_876,N_4903,N_4946);
and UO_877 (O_877,N_4967,N_4966);
nand UO_878 (O_878,N_4929,N_4902);
nand UO_879 (O_879,N_4903,N_4961);
and UO_880 (O_880,N_4951,N_4914);
nor UO_881 (O_881,N_4916,N_4993);
nor UO_882 (O_882,N_4971,N_4936);
nor UO_883 (O_883,N_4994,N_4907);
and UO_884 (O_884,N_4919,N_4992);
or UO_885 (O_885,N_4939,N_4932);
or UO_886 (O_886,N_4900,N_4978);
or UO_887 (O_887,N_4903,N_4930);
nand UO_888 (O_888,N_4979,N_4918);
nand UO_889 (O_889,N_4963,N_4949);
nor UO_890 (O_890,N_4928,N_4945);
or UO_891 (O_891,N_4969,N_4974);
xor UO_892 (O_892,N_4949,N_4929);
nor UO_893 (O_893,N_4909,N_4914);
nor UO_894 (O_894,N_4943,N_4969);
nor UO_895 (O_895,N_4900,N_4948);
xor UO_896 (O_896,N_4989,N_4948);
and UO_897 (O_897,N_4955,N_4902);
nor UO_898 (O_898,N_4943,N_4931);
and UO_899 (O_899,N_4926,N_4961);
xnor UO_900 (O_900,N_4937,N_4930);
or UO_901 (O_901,N_4969,N_4951);
and UO_902 (O_902,N_4977,N_4913);
xor UO_903 (O_903,N_4916,N_4935);
nand UO_904 (O_904,N_4981,N_4908);
and UO_905 (O_905,N_4942,N_4910);
nand UO_906 (O_906,N_4953,N_4945);
nand UO_907 (O_907,N_4947,N_4969);
and UO_908 (O_908,N_4970,N_4993);
or UO_909 (O_909,N_4962,N_4938);
nor UO_910 (O_910,N_4934,N_4926);
and UO_911 (O_911,N_4953,N_4960);
xor UO_912 (O_912,N_4929,N_4909);
or UO_913 (O_913,N_4981,N_4985);
nand UO_914 (O_914,N_4915,N_4929);
or UO_915 (O_915,N_4922,N_4984);
and UO_916 (O_916,N_4911,N_4939);
nand UO_917 (O_917,N_4976,N_4994);
and UO_918 (O_918,N_4948,N_4921);
nand UO_919 (O_919,N_4970,N_4921);
xnor UO_920 (O_920,N_4962,N_4902);
and UO_921 (O_921,N_4979,N_4914);
nand UO_922 (O_922,N_4910,N_4997);
xnor UO_923 (O_923,N_4951,N_4931);
xor UO_924 (O_924,N_4909,N_4988);
xor UO_925 (O_925,N_4942,N_4992);
or UO_926 (O_926,N_4908,N_4984);
xnor UO_927 (O_927,N_4938,N_4936);
or UO_928 (O_928,N_4933,N_4948);
nor UO_929 (O_929,N_4902,N_4925);
nor UO_930 (O_930,N_4915,N_4946);
or UO_931 (O_931,N_4998,N_4901);
nand UO_932 (O_932,N_4925,N_4976);
nor UO_933 (O_933,N_4925,N_4952);
xor UO_934 (O_934,N_4936,N_4933);
or UO_935 (O_935,N_4908,N_4943);
and UO_936 (O_936,N_4922,N_4969);
nand UO_937 (O_937,N_4938,N_4960);
nand UO_938 (O_938,N_4937,N_4985);
and UO_939 (O_939,N_4969,N_4915);
xor UO_940 (O_940,N_4971,N_4906);
or UO_941 (O_941,N_4970,N_4965);
nor UO_942 (O_942,N_4974,N_4928);
or UO_943 (O_943,N_4981,N_4952);
xor UO_944 (O_944,N_4909,N_4999);
nor UO_945 (O_945,N_4995,N_4932);
nor UO_946 (O_946,N_4908,N_4915);
nand UO_947 (O_947,N_4988,N_4982);
xnor UO_948 (O_948,N_4919,N_4977);
nand UO_949 (O_949,N_4989,N_4922);
nand UO_950 (O_950,N_4917,N_4994);
nand UO_951 (O_951,N_4908,N_4929);
xor UO_952 (O_952,N_4969,N_4944);
nor UO_953 (O_953,N_4914,N_4925);
xor UO_954 (O_954,N_4985,N_4970);
or UO_955 (O_955,N_4906,N_4974);
and UO_956 (O_956,N_4999,N_4969);
and UO_957 (O_957,N_4973,N_4980);
and UO_958 (O_958,N_4938,N_4974);
xnor UO_959 (O_959,N_4947,N_4921);
or UO_960 (O_960,N_4943,N_4998);
xor UO_961 (O_961,N_4990,N_4922);
nor UO_962 (O_962,N_4976,N_4947);
xnor UO_963 (O_963,N_4969,N_4941);
nor UO_964 (O_964,N_4934,N_4902);
and UO_965 (O_965,N_4948,N_4987);
xor UO_966 (O_966,N_4979,N_4905);
and UO_967 (O_967,N_4968,N_4981);
xnor UO_968 (O_968,N_4943,N_4903);
nand UO_969 (O_969,N_4973,N_4981);
xor UO_970 (O_970,N_4920,N_4991);
nand UO_971 (O_971,N_4965,N_4939);
and UO_972 (O_972,N_4940,N_4916);
xor UO_973 (O_973,N_4926,N_4976);
or UO_974 (O_974,N_4973,N_4937);
and UO_975 (O_975,N_4918,N_4916);
xnor UO_976 (O_976,N_4932,N_4946);
or UO_977 (O_977,N_4997,N_4933);
or UO_978 (O_978,N_4928,N_4911);
nand UO_979 (O_979,N_4937,N_4902);
xor UO_980 (O_980,N_4933,N_4916);
and UO_981 (O_981,N_4991,N_4914);
and UO_982 (O_982,N_4964,N_4966);
nand UO_983 (O_983,N_4945,N_4968);
nor UO_984 (O_984,N_4958,N_4993);
nor UO_985 (O_985,N_4989,N_4966);
or UO_986 (O_986,N_4965,N_4908);
nand UO_987 (O_987,N_4919,N_4943);
nor UO_988 (O_988,N_4926,N_4941);
nand UO_989 (O_989,N_4936,N_4989);
nand UO_990 (O_990,N_4912,N_4991);
or UO_991 (O_991,N_4936,N_4993);
xnor UO_992 (O_992,N_4927,N_4982);
or UO_993 (O_993,N_4969,N_4952);
xnor UO_994 (O_994,N_4992,N_4986);
and UO_995 (O_995,N_4905,N_4986);
and UO_996 (O_996,N_4936,N_4998);
nand UO_997 (O_997,N_4947,N_4901);
and UO_998 (O_998,N_4905,N_4903);
nand UO_999 (O_999,N_4954,N_4912);
endmodule