module basic_500_3000_500_50_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_487,In_250);
nand U1 (N_1,In_273,In_245);
nor U2 (N_2,In_341,In_422);
nand U3 (N_3,In_134,In_52);
nor U4 (N_4,In_121,In_50);
and U5 (N_5,In_164,In_254);
xor U6 (N_6,In_329,In_198);
or U7 (N_7,In_381,In_491);
or U8 (N_8,In_349,In_103);
nor U9 (N_9,In_377,In_217);
nand U10 (N_10,In_396,In_367);
nor U11 (N_11,In_441,In_335);
and U12 (N_12,In_306,In_202);
nor U13 (N_13,In_383,In_236);
and U14 (N_14,In_168,In_462);
or U15 (N_15,In_379,In_19);
nor U16 (N_16,In_151,In_117);
nand U17 (N_17,In_291,In_498);
nor U18 (N_18,In_384,In_222);
and U19 (N_19,In_21,In_209);
nor U20 (N_20,In_17,In_97);
nand U21 (N_21,In_106,In_118);
nand U22 (N_22,In_392,In_373);
nor U23 (N_23,In_0,In_128);
or U24 (N_24,In_249,In_44);
nor U25 (N_25,In_166,In_137);
or U26 (N_26,In_444,In_193);
nand U27 (N_27,In_362,In_9);
nand U28 (N_28,In_451,In_154);
or U29 (N_29,In_16,In_140);
or U30 (N_30,In_276,In_264);
and U31 (N_31,In_472,In_442);
and U32 (N_32,In_400,In_350);
or U33 (N_33,In_330,In_471);
or U34 (N_34,In_94,In_234);
nand U35 (N_35,In_275,In_135);
nand U36 (N_36,In_30,In_191);
nor U37 (N_37,In_211,In_443);
nand U38 (N_38,In_409,In_175);
nor U39 (N_39,In_78,In_160);
nor U40 (N_40,In_65,In_169);
or U41 (N_41,In_390,In_456);
and U42 (N_42,In_71,In_252);
and U43 (N_43,In_382,In_120);
or U44 (N_44,In_33,In_55);
nor U45 (N_45,In_133,In_369);
nand U46 (N_46,In_486,In_4);
or U47 (N_47,In_149,In_40);
nand U48 (N_48,In_380,In_453);
and U49 (N_49,In_60,In_212);
nor U50 (N_50,In_270,In_282);
and U51 (N_51,In_189,In_26);
and U52 (N_52,In_385,In_351);
nor U53 (N_53,In_87,In_468);
or U54 (N_54,In_455,In_267);
and U55 (N_55,In_296,In_495);
or U56 (N_56,In_263,In_63);
nand U57 (N_57,In_326,In_96);
xnor U58 (N_58,In_277,In_39);
and U59 (N_59,In_257,In_424);
nand U60 (N_60,In_307,N_41);
nor U61 (N_61,N_32,In_49);
or U62 (N_62,In_337,In_450);
nor U63 (N_63,In_51,In_14);
nand U64 (N_64,N_24,In_53);
or U65 (N_65,In_315,In_430);
nand U66 (N_66,In_253,In_186);
nor U67 (N_67,In_170,In_311);
nor U68 (N_68,In_32,In_100);
and U69 (N_69,In_181,N_2);
nand U70 (N_70,In_232,N_16);
nand U71 (N_71,In_320,In_338);
xnor U72 (N_72,In_62,In_79);
nor U73 (N_73,In_332,In_167);
and U74 (N_74,In_246,In_2);
nand U75 (N_75,In_425,In_23);
or U76 (N_76,In_297,In_477);
and U77 (N_77,In_475,In_298);
nor U78 (N_78,In_45,N_48);
nor U79 (N_79,In_397,N_27);
nor U80 (N_80,N_15,In_208);
or U81 (N_81,In_386,In_428);
nor U82 (N_82,In_493,In_7);
or U83 (N_83,In_204,In_439);
and U84 (N_84,In_159,In_139);
and U85 (N_85,In_287,In_301);
xor U86 (N_86,In_334,In_378);
and U87 (N_87,In_354,N_36);
nand U88 (N_88,In_346,In_247);
and U89 (N_89,In_288,In_388);
or U90 (N_90,In_131,In_344);
and U91 (N_91,N_20,In_130);
nand U92 (N_92,In_156,In_129);
nand U93 (N_93,In_454,In_331);
nand U94 (N_94,In_242,In_15);
nand U95 (N_95,In_153,In_283);
and U96 (N_96,In_469,In_219);
nand U97 (N_97,In_115,In_8);
and U98 (N_98,In_436,In_438);
and U99 (N_99,In_461,In_99);
nand U100 (N_100,In_229,In_426);
nor U101 (N_101,In_465,In_418);
and U102 (N_102,In_196,In_147);
and U103 (N_103,In_324,In_278);
nand U104 (N_104,In_101,In_490);
nor U105 (N_105,In_13,N_42);
or U106 (N_106,In_172,In_340);
or U107 (N_107,In_412,In_228);
nor U108 (N_108,In_41,In_81);
or U109 (N_109,N_46,In_31);
or U110 (N_110,In_104,In_393);
or U111 (N_111,In_448,In_132);
nor U112 (N_112,In_323,In_398);
nor U113 (N_113,In_110,In_358);
and U114 (N_114,In_423,In_59);
or U115 (N_115,In_479,In_427);
nand U116 (N_116,In_47,In_178);
or U117 (N_117,In_368,In_70);
and U118 (N_118,In_224,In_176);
or U119 (N_119,In_42,In_35);
and U120 (N_120,N_56,In_113);
and U121 (N_121,In_304,In_309);
or U122 (N_122,In_310,In_119);
or U123 (N_123,In_437,In_464);
nor U124 (N_124,In_74,In_294);
and U125 (N_125,In_312,In_6);
or U126 (N_126,N_60,In_12);
xnor U127 (N_127,In_333,In_43);
or U128 (N_128,N_66,In_109);
and U129 (N_129,N_22,N_104);
and U130 (N_130,In_480,In_405);
or U131 (N_131,In_210,In_321);
or U132 (N_132,N_12,N_89);
nand U133 (N_133,In_407,N_37);
nor U134 (N_134,In_457,In_286);
nand U135 (N_135,In_90,In_238);
nand U136 (N_136,N_57,In_459);
and U137 (N_137,In_36,N_10);
and U138 (N_138,N_82,N_119);
or U139 (N_139,In_492,In_375);
nor U140 (N_140,In_243,In_395);
nand U141 (N_141,In_230,In_325);
or U142 (N_142,In_201,In_488);
xnor U143 (N_143,In_419,In_187);
or U144 (N_144,In_80,N_105);
and U145 (N_145,In_458,In_163);
xor U146 (N_146,In_445,In_410);
xor U147 (N_147,In_225,In_279);
nand U148 (N_148,N_21,N_88);
nor U149 (N_149,N_77,In_145);
nor U150 (N_150,N_92,In_227);
nand U151 (N_151,In_190,N_49);
or U152 (N_152,In_83,In_484);
or U153 (N_153,In_162,In_370);
nor U154 (N_154,N_5,In_173);
nand U155 (N_155,In_299,In_274);
or U156 (N_156,In_417,In_372);
or U157 (N_157,In_481,In_497);
and U158 (N_158,N_58,In_218);
and U159 (N_159,N_81,In_75);
nor U160 (N_160,In_353,N_53);
or U161 (N_161,In_239,N_91);
and U162 (N_162,N_78,In_72);
nor U163 (N_163,In_256,In_446);
or U164 (N_164,N_102,In_293);
or U165 (N_165,N_50,In_387);
nand U166 (N_166,In_406,In_220);
nand U167 (N_167,In_91,In_214);
nor U168 (N_168,In_179,In_108);
nand U169 (N_169,In_322,In_197);
or U170 (N_170,In_295,In_415);
nand U171 (N_171,In_272,In_308);
and U172 (N_172,In_411,In_64);
nand U173 (N_173,N_67,In_391);
nor U174 (N_174,N_117,In_258);
or U175 (N_175,N_87,N_7);
xnor U176 (N_176,In_434,In_18);
nor U177 (N_177,In_376,In_404);
nand U178 (N_178,In_319,N_61);
nand U179 (N_179,N_26,In_356);
and U180 (N_180,In_98,In_474);
nand U181 (N_181,In_213,N_43);
or U182 (N_182,In_399,N_14);
xor U183 (N_183,N_151,In_216);
or U184 (N_184,In_192,In_374);
nor U185 (N_185,In_478,N_80);
or U186 (N_186,N_148,N_55);
and U187 (N_187,In_56,N_68);
or U188 (N_188,In_467,N_123);
or U189 (N_189,N_94,In_207);
and U190 (N_190,In_269,In_261);
nor U191 (N_191,In_182,In_327);
nor U192 (N_192,In_66,N_171);
nand U193 (N_193,In_313,In_460);
and U194 (N_194,In_260,In_174);
nand U195 (N_195,In_482,N_96);
and U196 (N_196,In_318,In_221);
nor U197 (N_197,N_110,In_73);
and U198 (N_198,In_302,In_116);
or U199 (N_199,In_266,In_69);
or U200 (N_200,N_133,In_150);
nand U201 (N_201,In_251,In_343);
and U202 (N_202,In_328,N_150);
nor U203 (N_203,N_116,N_31);
and U204 (N_204,N_44,N_152);
and U205 (N_205,N_164,In_280);
nor U206 (N_206,N_11,N_4);
or U207 (N_207,In_171,In_124);
and U208 (N_208,N_84,In_185);
nor U209 (N_209,N_172,N_69);
nand U210 (N_210,In_111,N_141);
and U211 (N_211,N_155,In_226);
and U212 (N_212,N_40,N_8);
or U213 (N_213,N_139,N_126);
or U214 (N_214,In_303,N_134);
nor U215 (N_215,N_85,In_57);
or U216 (N_216,In_177,In_352);
nor U217 (N_217,N_158,N_19);
and U218 (N_218,N_109,In_403);
and U219 (N_219,In_401,N_153);
and U220 (N_220,N_18,N_0);
or U221 (N_221,In_355,N_173);
nor U222 (N_222,In_494,In_24);
nor U223 (N_223,N_86,In_366);
or U224 (N_224,In_360,In_155);
or U225 (N_225,N_140,In_284);
or U226 (N_226,N_115,In_152);
nor U227 (N_227,N_179,N_17);
or U228 (N_228,In_433,In_416);
or U229 (N_229,In_414,In_84);
and U230 (N_230,In_194,In_144);
and U231 (N_231,In_314,In_499);
nor U232 (N_232,In_183,N_165);
nor U233 (N_233,In_3,In_180);
nand U234 (N_234,In_483,N_136);
nand U235 (N_235,In_489,In_339);
and U236 (N_236,In_496,In_259);
nand U237 (N_237,In_88,In_285);
and U238 (N_238,In_447,N_28);
nor U239 (N_239,In_364,In_289);
nor U240 (N_240,N_220,In_281);
or U241 (N_241,N_224,N_65);
and U242 (N_242,N_183,In_89);
and U243 (N_243,N_121,N_194);
nor U244 (N_244,In_271,In_54);
and U245 (N_245,N_62,In_27);
or U246 (N_246,In_205,In_233);
and U247 (N_247,N_120,In_10);
nand U248 (N_248,In_107,In_5);
xnor U249 (N_249,In_58,In_161);
and U250 (N_250,In_25,N_122);
nand U251 (N_251,In_206,In_429);
nand U252 (N_252,In_265,N_13);
or U253 (N_253,N_127,N_113);
nand U254 (N_254,In_348,N_191);
xor U255 (N_255,N_132,N_30);
nand U256 (N_256,In_143,In_215);
nand U257 (N_257,N_25,In_82);
nand U258 (N_258,N_1,N_149);
and U259 (N_259,In_449,N_231);
nor U260 (N_260,N_198,In_262);
or U261 (N_261,In_290,N_29);
nor U262 (N_262,N_235,In_141);
nand U263 (N_263,N_226,In_11);
nor U264 (N_264,N_76,In_61);
nor U265 (N_265,In_359,In_466);
xnor U266 (N_266,N_214,In_114);
and U267 (N_267,In_68,N_176);
nor U268 (N_268,N_9,N_73);
nand U269 (N_269,N_156,N_168);
or U270 (N_270,N_147,N_97);
or U271 (N_271,N_169,N_202);
xnor U272 (N_272,In_248,N_210);
or U273 (N_273,N_129,In_292);
nand U274 (N_274,N_200,N_72);
and U275 (N_275,N_237,In_200);
nor U276 (N_276,In_77,In_29);
nor U277 (N_277,N_54,In_300);
and U278 (N_278,In_138,N_112);
nand U279 (N_279,N_34,In_476);
or U280 (N_280,N_6,In_127);
nand U281 (N_281,N_209,N_114);
nand U282 (N_282,In_361,In_421);
and U283 (N_283,In_402,In_37);
or U284 (N_284,In_1,N_130);
nand U285 (N_285,N_182,N_192);
and U286 (N_286,N_203,In_158);
or U287 (N_287,N_197,N_145);
and U288 (N_288,N_181,N_228);
nor U289 (N_289,In_389,In_432);
nor U290 (N_290,N_186,In_420);
and U291 (N_291,N_144,N_51);
nor U292 (N_292,N_229,In_345);
or U293 (N_293,N_63,N_79);
nor U294 (N_294,N_178,N_195);
and U295 (N_295,N_207,In_244);
nor U296 (N_296,N_95,N_99);
or U297 (N_297,In_95,N_234);
or U298 (N_298,N_154,In_241);
or U299 (N_299,In_371,N_64);
xor U300 (N_300,N_242,N_283);
or U301 (N_301,N_268,N_90);
xor U302 (N_302,N_189,N_135);
and U303 (N_303,In_188,N_143);
xnor U304 (N_304,In_85,In_102);
or U305 (N_305,N_272,In_473);
and U306 (N_306,In_223,N_170);
and U307 (N_307,N_47,N_59);
nor U308 (N_308,N_247,In_255);
and U309 (N_309,In_485,N_240);
nand U310 (N_310,N_74,In_76);
and U311 (N_311,N_244,N_248);
or U312 (N_312,N_52,In_336);
xnor U313 (N_313,N_251,N_296);
nand U314 (N_314,N_124,N_193);
nor U315 (N_315,In_92,N_75);
nor U316 (N_316,N_245,N_142);
xor U317 (N_317,N_223,In_235);
nand U318 (N_318,In_148,N_280);
nand U319 (N_319,N_269,In_46);
nand U320 (N_320,In_165,N_295);
nor U321 (N_321,N_222,N_218);
or U322 (N_322,N_157,N_83);
nor U323 (N_323,In_408,In_452);
or U324 (N_324,In_125,N_190);
nor U325 (N_325,N_264,N_282);
nand U326 (N_326,N_299,N_286);
nor U327 (N_327,N_232,N_125);
and U328 (N_328,N_162,N_215);
and U329 (N_329,N_262,N_294);
and U330 (N_330,In_28,N_257);
nor U331 (N_331,N_225,N_45);
and U332 (N_332,N_177,N_111);
and U333 (N_333,N_35,In_122);
and U334 (N_334,N_106,N_216);
or U335 (N_335,N_199,N_188);
nor U336 (N_336,N_230,In_463);
and U337 (N_337,In_38,N_250);
or U338 (N_338,In_240,N_233);
nor U339 (N_339,N_39,N_258);
nor U340 (N_340,N_281,N_298);
nand U341 (N_341,In_435,N_270);
and U342 (N_342,N_175,N_276);
nand U343 (N_343,N_180,N_118);
and U344 (N_344,N_128,N_212);
nor U345 (N_345,N_289,N_261);
and U346 (N_346,In_268,N_208);
nand U347 (N_347,N_206,N_187);
nand U348 (N_348,N_108,N_267);
nor U349 (N_349,N_217,N_273);
or U350 (N_350,In_184,N_213);
and U351 (N_351,In_67,In_305);
or U352 (N_352,N_101,N_271);
nor U353 (N_353,N_205,N_288);
or U354 (N_354,N_239,In_105);
and U355 (N_355,In_48,N_23);
or U356 (N_356,N_146,N_293);
nor U357 (N_357,N_278,N_204);
or U358 (N_358,N_98,N_236);
nand U359 (N_359,In_126,N_211);
nor U360 (N_360,N_318,N_312);
nor U361 (N_361,N_354,N_323);
nor U362 (N_362,In_357,N_185);
nor U363 (N_363,N_315,N_329);
nor U364 (N_364,N_351,N_305);
or U365 (N_365,N_291,N_343);
nand U366 (N_366,N_227,In_440);
and U367 (N_367,In_413,N_266);
nor U368 (N_368,N_334,N_238);
nand U369 (N_369,N_246,In_231);
nor U370 (N_370,N_330,N_322);
and U371 (N_371,N_353,N_260);
or U372 (N_372,N_292,N_253);
nand U373 (N_373,N_357,N_160);
or U374 (N_374,In_237,N_319);
nand U375 (N_375,N_302,In_316);
nand U376 (N_376,In_470,N_317);
and U377 (N_377,N_355,N_196);
nor U378 (N_378,N_303,In_431);
or U379 (N_379,N_252,In_394);
or U380 (N_380,N_174,N_314);
nor U381 (N_381,In_34,N_359);
or U382 (N_382,N_321,N_100);
or U383 (N_383,N_326,N_332);
or U384 (N_384,In_342,N_255);
nand U385 (N_385,N_103,N_308);
nand U386 (N_386,In_199,N_304);
nor U387 (N_387,In_142,In_365);
nand U388 (N_388,In_195,N_279);
nor U389 (N_389,In_203,N_137);
nand U390 (N_390,In_20,N_325);
nor U391 (N_391,N_320,N_290);
nor U392 (N_392,N_341,N_301);
nor U393 (N_393,N_306,In_347);
and U394 (N_394,N_346,N_316);
nand U395 (N_395,N_336,N_311);
nor U396 (N_396,N_167,N_33);
or U397 (N_397,N_331,In_317);
or U398 (N_398,N_241,N_159);
nand U399 (N_399,N_166,N_284);
and U400 (N_400,N_259,N_71);
nand U401 (N_401,N_348,N_70);
nor U402 (N_402,N_256,N_352);
and U403 (N_403,N_356,N_327);
nor U404 (N_404,N_38,In_136);
and U405 (N_405,In_22,N_243);
and U406 (N_406,N_131,N_307);
and U407 (N_407,In_86,N_93);
or U408 (N_408,N_339,N_249);
nor U409 (N_409,In_93,N_324);
and U410 (N_410,N_287,N_285);
nand U411 (N_411,N_221,N_340);
or U412 (N_412,N_274,In_146);
nand U413 (N_413,In_157,N_338);
and U414 (N_414,N_342,N_3);
nor U415 (N_415,N_358,N_138);
nor U416 (N_416,N_335,N_350);
nor U417 (N_417,N_163,N_328);
or U418 (N_418,N_344,N_349);
or U419 (N_419,N_265,In_123);
nand U420 (N_420,N_107,N_309);
and U421 (N_421,N_370,N_360);
nor U422 (N_422,N_384,N_400);
and U423 (N_423,N_406,N_219);
nand U424 (N_424,N_380,N_378);
nand U425 (N_425,N_161,In_112);
nor U426 (N_426,N_409,N_381);
and U427 (N_427,N_390,N_414);
or U428 (N_428,N_399,N_391);
or U429 (N_429,N_333,N_394);
or U430 (N_430,N_410,N_382);
or U431 (N_431,N_337,N_397);
xor U432 (N_432,N_413,N_368);
or U433 (N_433,N_416,N_411);
nand U434 (N_434,N_263,N_407);
and U435 (N_435,N_345,N_395);
and U436 (N_436,N_365,N_377);
nor U437 (N_437,N_387,N_389);
nor U438 (N_438,N_402,N_310);
nor U439 (N_439,N_363,N_419);
and U440 (N_440,N_375,N_386);
nor U441 (N_441,N_277,N_376);
and U442 (N_442,N_371,N_404);
nor U443 (N_443,N_364,N_254);
and U444 (N_444,N_361,N_418);
nor U445 (N_445,N_313,In_363);
and U446 (N_446,N_275,N_417);
nor U447 (N_447,N_396,N_388);
or U448 (N_448,N_405,N_369);
nor U449 (N_449,N_383,N_367);
or U450 (N_450,N_201,N_300);
nand U451 (N_451,N_403,N_379);
and U452 (N_452,N_297,N_373);
or U453 (N_453,N_392,N_366);
or U454 (N_454,N_408,N_362);
nand U455 (N_455,N_385,N_415);
and U456 (N_456,N_347,N_412);
and U457 (N_457,N_372,N_184);
or U458 (N_458,N_401,N_374);
and U459 (N_459,N_398,N_393);
nor U460 (N_460,N_300,N_297);
nor U461 (N_461,In_112,N_309);
nand U462 (N_462,N_361,N_380);
or U463 (N_463,N_313,N_415);
nand U464 (N_464,N_376,N_387);
or U465 (N_465,N_297,N_368);
and U466 (N_466,N_201,N_107);
and U467 (N_467,N_219,N_390);
nand U468 (N_468,N_365,N_161);
nand U469 (N_469,N_418,N_161);
and U470 (N_470,N_362,N_364);
or U471 (N_471,N_361,N_390);
and U472 (N_472,N_402,N_366);
nand U473 (N_473,N_297,N_408);
nand U474 (N_474,N_372,N_371);
nor U475 (N_475,N_376,N_345);
or U476 (N_476,N_377,N_390);
and U477 (N_477,In_112,N_380);
and U478 (N_478,N_378,N_366);
or U479 (N_479,N_380,N_387);
nand U480 (N_480,N_475,N_455);
nand U481 (N_481,N_468,N_442);
and U482 (N_482,N_461,N_453);
nor U483 (N_483,N_423,N_430);
or U484 (N_484,N_433,N_431);
and U485 (N_485,N_459,N_474);
nor U486 (N_486,N_471,N_470);
and U487 (N_487,N_448,N_456);
nor U488 (N_488,N_472,N_449);
nand U489 (N_489,N_477,N_447);
nand U490 (N_490,N_422,N_432);
nor U491 (N_491,N_439,N_421);
nor U492 (N_492,N_464,N_444);
or U493 (N_493,N_450,N_463);
nand U494 (N_494,N_425,N_427);
or U495 (N_495,N_462,N_435);
nand U496 (N_496,N_437,N_476);
or U497 (N_497,N_445,N_428);
nand U498 (N_498,N_443,N_454);
nand U499 (N_499,N_465,N_446);
and U500 (N_500,N_473,N_434);
nand U501 (N_501,N_466,N_441);
or U502 (N_502,N_424,N_452);
or U503 (N_503,N_438,N_420);
and U504 (N_504,N_467,N_458);
nor U505 (N_505,N_479,N_426);
nor U506 (N_506,N_429,N_436);
nor U507 (N_507,N_451,N_478);
nand U508 (N_508,N_460,N_440);
nand U509 (N_509,N_469,N_457);
and U510 (N_510,N_461,N_424);
and U511 (N_511,N_420,N_434);
or U512 (N_512,N_457,N_470);
or U513 (N_513,N_436,N_469);
and U514 (N_514,N_430,N_442);
nor U515 (N_515,N_443,N_426);
or U516 (N_516,N_468,N_463);
or U517 (N_517,N_436,N_430);
or U518 (N_518,N_473,N_437);
nand U519 (N_519,N_479,N_427);
and U520 (N_520,N_459,N_430);
nor U521 (N_521,N_432,N_445);
nor U522 (N_522,N_445,N_446);
and U523 (N_523,N_432,N_472);
nand U524 (N_524,N_421,N_424);
or U525 (N_525,N_463,N_470);
nand U526 (N_526,N_473,N_430);
nor U527 (N_527,N_441,N_478);
or U528 (N_528,N_432,N_459);
and U529 (N_529,N_455,N_421);
and U530 (N_530,N_449,N_443);
or U531 (N_531,N_445,N_452);
nand U532 (N_532,N_421,N_476);
or U533 (N_533,N_430,N_443);
nor U534 (N_534,N_445,N_437);
nand U535 (N_535,N_433,N_477);
and U536 (N_536,N_475,N_478);
and U537 (N_537,N_468,N_479);
and U538 (N_538,N_462,N_427);
nor U539 (N_539,N_440,N_451);
or U540 (N_540,N_491,N_539);
nor U541 (N_541,N_529,N_521);
nand U542 (N_542,N_536,N_534);
nor U543 (N_543,N_489,N_530);
and U544 (N_544,N_496,N_525);
or U545 (N_545,N_483,N_493);
and U546 (N_546,N_533,N_497);
or U547 (N_547,N_486,N_517);
nor U548 (N_548,N_537,N_526);
and U549 (N_549,N_490,N_507);
or U550 (N_550,N_538,N_516);
nand U551 (N_551,N_528,N_492);
nand U552 (N_552,N_501,N_495);
nand U553 (N_553,N_494,N_512);
nand U554 (N_554,N_488,N_535);
nand U555 (N_555,N_509,N_482);
and U556 (N_556,N_518,N_531);
nand U557 (N_557,N_520,N_485);
nor U558 (N_558,N_508,N_487);
and U559 (N_559,N_524,N_499);
and U560 (N_560,N_532,N_505);
nor U561 (N_561,N_506,N_523);
or U562 (N_562,N_502,N_510);
nand U563 (N_563,N_504,N_498);
or U564 (N_564,N_515,N_519);
nor U565 (N_565,N_522,N_481);
nand U566 (N_566,N_500,N_514);
nand U567 (N_567,N_511,N_480);
nor U568 (N_568,N_527,N_513);
and U569 (N_569,N_484,N_503);
or U570 (N_570,N_515,N_501);
nor U571 (N_571,N_523,N_492);
or U572 (N_572,N_534,N_528);
or U573 (N_573,N_528,N_486);
nand U574 (N_574,N_506,N_486);
or U575 (N_575,N_490,N_501);
or U576 (N_576,N_481,N_520);
nand U577 (N_577,N_499,N_532);
and U578 (N_578,N_519,N_494);
or U579 (N_579,N_485,N_528);
nand U580 (N_580,N_528,N_515);
nor U581 (N_581,N_524,N_490);
or U582 (N_582,N_504,N_486);
nand U583 (N_583,N_481,N_514);
nand U584 (N_584,N_495,N_538);
nand U585 (N_585,N_529,N_484);
and U586 (N_586,N_490,N_526);
nor U587 (N_587,N_532,N_513);
nor U588 (N_588,N_514,N_493);
and U589 (N_589,N_538,N_492);
nor U590 (N_590,N_533,N_495);
or U591 (N_591,N_499,N_529);
nor U592 (N_592,N_513,N_489);
nand U593 (N_593,N_507,N_485);
nor U594 (N_594,N_492,N_537);
or U595 (N_595,N_507,N_531);
or U596 (N_596,N_500,N_504);
and U597 (N_597,N_525,N_522);
or U598 (N_598,N_531,N_516);
nand U599 (N_599,N_506,N_484);
or U600 (N_600,N_575,N_578);
nor U601 (N_601,N_596,N_592);
nand U602 (N_602,N_571,N_544);
nor U603 (N_603,N_565,N_552);
or U604 (N_604,N_559,N_597);
or U605 (N_605,N_593,N_581);
nand U606 (N_606,N_567,N_572);
and U607 (N_607,N_594,N_598);
and U608 (N_608,N_568,N_557);
nand U609 (N_609,N_550,N_573);
nor U610 (N_610,N_579,N_558);
nand U611 (N_611,N_547,N_560);
nor U612 (N_612,N_545,N_564);
or U613 (N_613,N_577,N_555);
or U614 (N_614,N_586,N_570);
and U615 (N_615,N_556,N_588);
and U616 (N_616,N_548,N_549);
or U617 (N_617,N_584,N_554);
and U618 (N_618,N_553,N_540);
nand U619 (N_619,N_561,N_595);
and U620 (N_620,N_587,N_541);
nor U621 (N_621,N_582,N_569);
nand U622 (N_622,N_542,N_562);
nor U623 (N_623,N_551,N_563);
nand U624 (N_624,N_590,N_543);
or U625 (N_625,N_574,N_599);
nor U626 (N_626,N_583,N_591);
and U627 (N_627,N_566,N_585);
nand U628 (N_628,N_546,N_580);
xor U629 (N_629,N_576,N_589);
nor U630 (N_630,N_585,N_558);
and U631 (N_631,N_598,N_542);
nand U632 (N_632,N_566,N_590);
nor U633 (N_633,N_597,N_564);
and U634 (N_634,N_577,N_544);
nor U635 (N_635,N_578,N_548);
xnor U636 (N_636,N_561,N_598);
or U637 (N_637,N_543,N_552);
nand U638 (N_638,N_546,N_599);
nor U639 (N_639,N_568,N_558);
nor U640 (N_640,N_575,N_598);
nor U641 (N_641,N_599,N_584);
nor U642 (N_642,N_595,N_590);
and U643 (N_643,N_572,N_582);
and U644 (N_644,N_575,N_585);
nor U645 (N_645,N_561,N_583);
and U646 (N_646,N_595,N_570);
nor U647 (N_647,N_582,N_573);
or U648 (N_648,N_574,N_542);
nand U649 (N_649,N_563,N_582);
and U650 (N_650,N_547,N_551);
nor U651 (N_651,N_587,N_542);
and U652 (N_652,N_555,N_587);
or U653 (N_653,N_562,N_570);
nor U654 (N_654,N_557,N_543);
and U655 (N_655,N_585,N_542);
nor U656 (N_656,N_580,N_569);
and U657 (N_657,N_594,N_576);
nand U658 (N_658,N_591,N_542);
or U659 (N_659,N_563,N_592);
and U660 (N_660,N_649,N_618);
or U661 (N_661,N_652,N_634);
nor U662 (N_662,N_651,N_609);
or U663 (N_663,N_607,N_625);
nor U664 (N_664,N_639,N_624);
and U665 (N_665,N_600,N_659);
nand U666 (N_666,N_611,N_627);
nand U667 (N_667,N_613,N_605);
and U668 (N_668,N_604,N_628);
nor U669 (N_669,N_644,N_612);
or U670 (N_670,N_619,N_633);
nor U671 (N_671,N_635,N_626);
nand U672 (N_672,N_647,N_614);
or U673 (N_673,N_658,N_630);
or U674 (N_674,N_620,N_657);
and U675 (N_675,N_641,N_643);
nor U676 (N_676,N_617,N_610);
nand U677 (N_677,N_616,N_602);
or U678 (N_678,N_650,N_623);
or U679 (N_679,N_603,N_632);
nor U680 (N_680,N_606,N_640);
or U681 (N_681,N_655,N_621);
or U682 (N_682,N_638,N_646);
and U683 (N_683,N_653,N_629);
or U684 (N_684,N_656,N_648);
nand U685 (N_685,N_631,N_636);
or U686 (N_686,N_645,N_654);
nor U687 (N_687,N_642,N_601);
nand U688 (N_688,N_637,N_615);
xnor U689 (N_689,N_608,N_622);
and U690 (N_690,N_601,N_613);
or U691 (N_691,N_647,N_649);
nand U692 (N_692,N_619,N_627);
and U693 (N_693,N_656,N_606);
nand U694 (N_694,N_653,N_633);
xnor U695 (N_695,N_605,N_655);
and U696 (N_696,N_604,N_655);
nor U697 (N_697,N_646,N_645);
nand U698 (N_698,N_617,N_639);
and U699 (N_699,N_648,N_624);
and U700 (N_700,N_651,N_603);
or U701 (N_701,N_611,N_626);
nor U702 (N_702,N_606,N_643);
or U703 (N_703,N_604,N_605);
and U704 (N_704,N_618,N_640);
nand U705 (N_705,N_615,N_613);
nand U706 (N_706,N_644,N_642);
nand U707 (N_707,N_642,N_624);
nand U708 (N_708,N_627,N_604);
nand U709 (N_709,N_628,N_653);
nand U710 (N_710,N_638,N_611);
and U711 (N_711,N_648,N_626);
nand U712 (N_712,N_622,N_600);
nand U713 (N_713,N_636,N_656);
or U714 (N_714,N_645,N_644);
and U715 (N_715,N_618,N_628);
and U716 (N_716,N_620,N_605);
nor U717 (N_717,N_628,N_643);
nand U718 (N_718,N_607,N_648);
nor U719 (N_719,N_644,N_625);
and U720 (N_720,N_692,N_703);
and U721 (N_721,N_718,N_674);
nor U722 (N_722,N_663,N_708);
and U723 (N_723,N_662,N_695);
or U724 (N_724,N_672,N_668);
nor U725 (N_725,N_661,N_697);
or U726 (N_726,N_706,N_677);
or U727 (N_727,N_682,N_685);
nor U728 (N_728,N_689,N_716);
nor U729 (N_729,N_701,N_669);
nand U730 (N_730,N_714,N_704);
and U731 (N_731,N_671,N_681);
and U732 (N_732,N_675,N_717);
or U733 (N_733,N_688,N_711);
nor U734 (N_734,N_699,N_710);
nand U735 (N_735,N_684,N_683);
and U736 (N_736,N_690,N_694);
or U737 (N_737,N_691,N_715);
xor U738 (N_738,N_687,N_693);
and U739 (N_739,N_667,N_664);
or U740 (N_740,N_698,N_680);
and U741 (N_741,N_660,N_678);
xnor U742 (N_742,N_673,N_665);
or U743 (N_743,N_709,N_707);
or U744 (N_744,N_713,N_679);
nor U745 (N_745,N_666,N_712);
nand U746 (N_746,N_670,N_700);
nand U747 (N_747,N_719,N_686);
and U748 (N_748,N_705,N_696);
or U749 (N_749,N_702,N_676);
and U750 (N_750,N_675,N_698);
and U751 (N_751,N_690,N_674);
and U752 (N_752,N_684,N_662);
or U753 (N_753,N_670,N_681);
nor U754 (N_754,N_692,N_675);
or U755 (N_755,N_700,N_719);
nand U756 (N_756,N_700,N_699);
or U757 (N_757,N_676,N_670);
nor U758 (N_758,N_715,N_663);
nand U759 (N_759,N_689,N_671);
nand U760 (N_760,N_689,N_713);
xnor U761 (N_761,N_670,N_677);
or U762 (N_762,N_719,N_712);
nor U763 (N_763,N_677,N_688);
nand U764 (N_764,N_712,N_698);
nor U765 (N_765,N_670,N_698);
nand U766 (N_766,N_693,N_703);
nand U767 (N_767,N_716,N_678);
or U768 (N_768,N_703,N_702);
and U769 (N_769,N_712,N_660);
nand U770 (N_770,N_685,N_719);
nand U771 (N_771,N_673,N_705);
or U772 (N_772,N_685,N_690);
and U773 (N_773,N_664,N_712);
and U774 (N_774,N_673,N_718);
xnor U775 (N_775,N_686,N_707);
and U776 (N_776,N_696,N_665);
nand U777 (N_777,N_707,N_711);
and U778 (N_778,N_700,N_662);
nand U779 (N_779,N_717,N_676);
and U780 (N_780,N_760,N_722);
nor U781 (N_781,N_739,N_721);
nand U782 (N_782,N_764,N_771);
and U783 (N_783,N_731,N_756);
nor U784 (N_784,N_769,N_736);
nand U785 (N_785,N_754,N_751);
or U786 (N_786,N_765,N_767);
or U787 (N_787,N_758,N_747);
nand U788 (N_788,N_777,N_729);
and U789 (N_789,N_757,N_761);
or U790 (N_790,N_743,N_772);
or U791 (N_791,N_779,N_773);
nor U792 (N_792,N_774,N_766);
or U793 (N_793,N_724,N_735);
or U794 (N_794,N_753,N_759);
nor U795 (N_795,N_726,N_727);
and U796 (N_796,N_768,N_770);
nand U797 (N_797,N_748,N_738);
nand U798 (N_798,N_741,N_740);
nor U799 (N_799,N_732,N_763);
nor U800 (N_800,N_733,N_720);
or U801 (N_801,N_750,N_776);
and U802 (N_802,N_728,N_737);
and U803 (N_803,N_775,N_742);
and U804 (N_804,N_745,N_734);
or U805 (N_805,N_778,N_755);
nand U806 (N_806,N_746,N_749);
and U807 (N_807,N_762,N_723);
or U808 (N_808,N_725,N_752);
and U809 (N_809,N_730,N_744);
nand U810 (N_810,N_734,N_757);
and U811 (N_811,N_757,N_770);
and U812 (N_812,N_771,N_740);
and U813 (N_813,N_738,N_759);
or U814 (N_814,N_750,N_774);
or U815 (N_815,N_762,N_748);
and U816 (N_816,N_720,N_739);
or U817 (N_817,N_720,N_736);
or U818 (N_818,N_745,N_757);
and U819 (N_819,N_734,N_749);
nor U820 (N_820,N_724,N_748);
and U821 (N_821,N_740,N_736);
or U822 (N_822,N_729,N_721);
and U823 (N_823,N_724,N_728);
nor U824 (N_824,N_732,N_738);
or U825 (N_825,N_727,N_748);
xor U826 (N_826,N_759,N_768);
nor U827 (N_827,N_738,N_739);
xnor U828 (N_828,N_727,N_752);
nand U829 (N_829,N_763,N_759);
xor U830 (N_830,N_766,N_739);
nor U831 (N_831,N_778,N_735);
nor U832 (N_832,N_764,N_747);
nor U833 (N_833,N_762,N_749);
nand U834 (N_834,N_743,N_734);
or U835 (N_835,N_720,N_778);
nor U836 (N_836,N_759,N_746);
and U837 (N_837,N_732,N_730);
or U838 (N_838,N_766,N_731);
and U839 (N_839,N_739,N_764);
or U840 (N_840,N_797,N_794);
and U841 (N_841,N_800,N_801);
xor U842 (N_842,N_822,N_839);
or U843 (N_843,N_834,N_807);
nand U844 (N_844,N_829,N_826);
or U845 (N_845,N_833,N_817);
nand U846 (N_846,N_790,N_836);
and U847 (N_847,N_802,N_835);
nand U848 (N_848,N_820,N_806);
nor U849 (N_849,N_785,N_808);
and U850 (N_850,N_798,N_821);
nor U851 (N_851,N_791,N_799);
nand U852 (N_852,N_792,N_832);
or U853 (N_853,N_823,N_819);
nor U854 (N_854,N_818,N_787);
and U855 (N_855,N_796,N_812);
nand U856 (N_856,N_816,N_824);
nor U857 (N_857,N_804,N_830);
and U858 (N_858,N_828,N_782);
nand U859 (N_859,N_803,N_838);
and U860 (N_860,N_811,N_825);
and U861 (N_861,N_810,N_781);
or U862 (N_862,N_793,N_815);
and U863 (N_863,N_814,N_795);
nand U864 (N_864,N_837,N_789);
nor U865 (N_865,N_783,N_827);
nand U866 (N_866,N_788,N_784);
nor U867 (N_867,N_786,N_813);
or U868 (N_868,N_805,N_809);
or U869 (N_869,N_780,N_831);
nor U870 (N_870,N_829,N_832);
and U871 (N_871,N_794,N_781);
or U872 (N_872,N_816,N_820);
or U873 (N_873,N_784,N_822);
nor U874 (N_874,N_829,N_793);
nand U875 (N_875,N_792,N_788);
and U876 (N_876,N_797,N_821);
nand U877 (N_877,N_787,N_795);
nor U878 (N_878,N_818,N_813);
nand U879 (N_879,N_830,N_838);
or U880 (N_880,N_806,N_814);
and U881 (N_881,N_788,N_828);
or U882 (N_882,N_788,N_824);
nand U883 (N_883,N_828,N_829);
nor U884 (N_884,N_822,N_786);
or U885 (N_885,N_824,N_802);
or U886 (N_886,N_786,N_789);
nand U887 (N_887,N_785,N_828);
nor U888 (N_888,N_807,N_789);
nor U889 (N_889,N_833,N_813);
nor U890 (N_890,N_785,N_812);
or U891 (N_891,N_798,N_781);
xor U892 (N_892,N_839,N_788);
or U893 (N_893,N_830,N_839);
or U894 (N_894,N_800,N_836);
nor U895 (N_895,N_789,N_825);
nor U896 (N_896,N_813,N_836);
xor U897 (N_897,N_782,N_795);
and U898 (N_898,N_783,N_826);
or U899 (N_899,N_816,N_828);
nor U900 (N_900,N_852,N_853);
xor U901 (N_901,N_894,N_898);
and U902 (N_902,N_883,N_865);
and U903 (N_903,N_868,N_846);
nand U904 (N_904,N_870,N_848);
and U905 (N_905,N_866,N_863);
and U906 (N_906,N_871,N_874);
and U907 (N_907,N_878,N_860);
or U908 (N_908,N_877,N_844);
or U909 (N_909,N_882,N_845);
nand U910 (N_910,N_876,N_847);
and U911 (N_911,N_892,N_859);
xor U912 (N_912,N_890,N_889);
or U913 (N_913,N_857,N_841);
nand U914 (N_914,N_862,N_886);
nor U915 (N_915,N_879,N_884);
nor U916 (N_916,N_875,N_867);
nor U917 (N_917,N_849,N_897);
and U918 (N_918,N_864,N_885);
and U919 (N_919,N_896,N_858);
nand U920 (N_920,N_895,N_887);
or U921 (N_921,N_880,N_855);
nor U922 (N_922,N_843,N_873);
or U923 (N_923,N_840,N_842);
nor U924 (N_924,N_891,N_861);
and U925 (N_925,N_872,N_899);
or U926 (N_926,N_888,N_869);
nand U927 (N_927,N_854,N_851);
nor U928 (N_928,N_850,N_881);
and U929 (N_929,N_856,N_893);
nand U930 (N_930,N_880,N_877);
or U931 (N_931,N_889,N_858);
nor U932 (N_932,N_849,N_840);
or U933 (N_933,N_893,N_879);
and U934 (N_934,N_876,N_851);
and U935 (N_935,N_882,N_858);
or U936 (N_936,N_899,N_862);
nand U937 (N_937,N_877,N_873);
xor U938 (N_938,N_859,N_895);
and U939 (N_939,N_864,N_840);
and U940 (N_940,N_855,N_886);
or U941 (N_941,N_870,N_879);
nor U942 (N_942,N_850,N_878);
nand U943 (N_943,N_875,N_878);
nand U944 (N_944,N_868,N_850);
and U945 (N_945,N_880,N_851);
nand U946 (N_946,N_865,N_880);
and U947 (N_947,N_844,N_859);
nand U948 (N_948,N_880,N_858);
nand U949 (N_949,N_878,N_862);
and U950 (N_950,N_854,N_862);
and U951 (N_951,N_889,N_887);
nand U952 (N_952,N_897,N_894);
nand U953 (N_953,N_856,N_855);
or U954 (N_954,N_891,N_862);
or U955 (N_955,N_859,N_879);
and U956 (N_956,N_869,N_854);
nor U957 (N_957,N_896,N_881);
or U958 (N_958,N_848,N_854);
nor U959 (N_959,N_858,N_867);
nor U960 (N_960,N_904,N_922);
and U961 (N_961,N_920,N_919);
and U962 (N_962,N_957,N_915);
or U963 (N_963,N_911,N_954);
and U964 (N_964,N_901,N_959);
nor U965 (N_965,N_929,N_905);
nor U966 (N_966,N_914,N_917);
nor U967 (N_967,N_948,N_908);
nor U968 (N_968,N_938,N_925);
nor U969 (N_969,N_928,N_932);
or U970 (N_970,N_909,N_937);
xnor U971 (N_971,N_907,N_931);
nand U972 (N_972,N_947,N_944);
and U973 (N_973,N_955,N_918);
xnor U974 (N_974,N_933,N_953);
xor U975 (N_975,N_913,N_934);
or U976 (N_976,N_949,N_923);
nand U977 (N_977,N_902,N_916);
nand U978 (N_978,N_945,N_900);
nand U979 (N_979,N_935,N_940);
and U980 (N_980,N_941,N_958);
and U981 (N_981,N_939,N_952);
nor U982 (N_982,N_910,N_950);
nand U983 (N_983,N_956,N_930);
and U984 (N_984,N_926,N_924);
nor U985 (N_985,N_946,N_903);
nand U986 (N_986,N_951,N_927);
nor U987 (N_987,N_921,N_912);
or U988 (N_988,N_943,N_936);
nor U989 (N_989,N_906,N_942);
nor U990 (N_990,N_941,N_949);
or U991 (N_991,N_927,N_926);
and U992 (N_992,N_947,N_939);
nor U993 (N_993,N_938,N_917);
or U994 (N_994,N_958,N_915);
nor U995 (N_995,N_947,N_913);
xnor U996 (N_996,N_949,N_905);
or U997 (N_997,N_906,N_944);
nor U998 (N_998,N_951,N_935);
and U999 (N_999,N_906,N_953);
and U1000 (N_1000,N_921,N_958);
or U1001 (N_1001,N_900,N_943);
nor U1002 (N_1002,N_957,N_931);
nor U1003 (N_1003,N_913,N_950);
nor U1004 (N_1004,N_950,N_920);
nor U1005 (N_1005,N_942,N_919);
or U1006 (N_1006,N_949,N_933);
xnor U1007 (N_1007,N_914,N_923);
nand U1008 (N_1008,N_935,N_945);
xnor U1009 (N_1009,N_925,N_922);
nor U1010 (N_1010,N_923,N_946);
or U1011 (N_1011,N_936,N_928);
xor U1012 (N_1012,N_902,N_901);
xnor U1013 (N_1013,N_927,N_928);
or U1014 (N_1014,N_929,N_904);
nor U1015 (N_1015,N_920,N_907);
or U1016 (N_1016,N_929,N_933);
nor U1017 (N_1017,N_928,N_952);
and U1018 (N_1018,N_925,N_945);
nand U1019 (N_1019,N_907,N_954);
xnor U1020 (N_1020,N_997,N_991);
nand U1021 (N_1021,N_1019,N_985);
nand U1022 (N_1022,N_1008,N_965);
or U1023 (N_1023,N_969,N_1000);
or U1024 (N_1024,N_1015,N_1013);
nand U1025 (N_1025,N_992,N_1001);
or U1026 (N_1026,N_979,N_1014);
or U1027 (N_1027,N_999,N_962);
nor U1028 (N_1028,N_1012,N_994);
nor U1029 (N_1029,N_1002,N_1018);
and U1030 (N_1030,N_1009,N_1006);
or U1031 (N_1031,N_998,N_981);
nand U1032 (N_1032,N_975,N_989);
nor U1033 (N_1033,N_1010,N_986);
and U1034 (N_1034,N_976,N_967);
and U1035 (N_1035,N_961,N_978);
xnor U1036 (N_1036,N_995,N_970);
nand U1037 (N_1037,N_968,N_977);
and U1038 (N_1038,N_980,N_1007);
or U1039 (N_1039,N_1005,N_966);
nand U1040 (N_1040,N_973,N_964);
and U1041 (N_1041,N_1016,N_1004);
nor U1042 (N_1042,N_983,N_963);
and U1043 (N_1043,N_996,N_982);
nor U1044 (N_1044,N_972,N_974);
nand U1045 (N_1045,N_984,N_1003);
and U1046 (N_1046,N_971,N_960);
nand U1047 (N_1047,N_990,N_1017);
or U1048 (N_1048,N_1011,N_987);
nor U1049 (N_1049,N_988,N_993);
and U1050 (N_1050,N_1016,N_965);
and U1051 (N_1051,N_1005,N_1011);
nor U1052 (N_1052,N_960,N_1004);
or U1053 (N_1053,N_977,N_1002);
nor U1054 (N_1054,N_976,N_989);
nor U1055 (N_1055,N_1005,N_991);
and U1056 (N_1056,N_1014,N_1002);
nand U1057 (N_1057,N_973,N_962);
or U1058 (N_1058,N_969,N_1007);
nand U1059 (N_1059,N_985,N_983);
and U1060 (N_1060,N_980,N_965);
and U1061 (N_1061,N_963,N_969);
nor U1062 (N_1062,N_1011,N_964);
nand U1063 (N_1063,N_982,N_991);
and U1064 (N_1064,N_969,N_989);
and U1065 (N_1065,N_985,N_1009);
or U1066 (N_1066,N_1013,N_966);
and U1067 (N_1067,N_1018,N_993);
nand U1068 (N_1068,N_1011,N_988);
and U1069 (N_1069,N_993,N_991);
or U1070 (N_1070,N_1019,N_988);
nand U1071 (N_1071,N_970,N_1013);
and U1072 (N_1072,N_988,N_967);
and U1073 (N_1073,N_967,N_968);
nor U1074 (N_1074,N_974,N_992);
and U1075 (N_1075,N_961,N_989);
and U1076 (N_1076,N_981,N_986);
nand U1077 (N_1077,N_990,N_972);
and U1078 (N_1078,N_971,N_996);
and U1079 (N_1079,N_962,N_993);
and U1080 (N_1080,N_1061,N_1064);
nor U1081 (N_1081,N_1058,N_1068);
nand U1082 (N_1082,N_1028,N_1070);
nor U1083 (N_1083,N_1037,N_1026);
nor U1084 (N_1084,N_1073,N_1056);
nand U1085 (N_1085,N_1044,N_1054);
nor U1086 (N_1086,N_1074,N_1060);
nand U1087 (N_1087,N_1065,N_1035);
nor U1088 (N_1088,N_1050,N_1071);
nor U1089 (N_1089,N_1055,N_1034);
nand U1090 (N_1090,N_1043,N_1039);
and U1091 (N_1091,N_1048,N_1041);
and U1092 (N_1092,N_1076,N_1072);
or U1093 (N_1093,N_1022,N_1052);
nor U1094 (N_1094,N_1063,N_1046);
and U1095 (N_1095,N_1042,N_1067);
nor U1096 (N_1096,N_1059,N_1051);
nand U1097 (N_1097,N_1078,N_1027);
nor U1098 (N_1098,N_1047,N_1031);
and U1099 (N_1099,N_1075,N_1077);
nor U1100 (N_1100,N_1069,N_1040);
nand U1101 (N_1101,N_1025,N_1023);
or U1102 (N_1102,N_1030,N_1036);
or U1103 (N_1103,N_1057,N_1038);
or U1104 (N_1104,N_1062,N_1045);
nand U1105 (N_1105,N_1024,N_1020);
nor U1106 (N_1106,N_1032,N_1033);
or U1107 (N_1107,N_1079,N_1021);
or U1108 (N_1108,N_1053,N_1029);
and U1109 (N_1109,N_1049,N_1066);
and U1110 (N_1110,N_1027,N_1020);
or U1111 (N_1111,N_1075,N_1057);
or U1112 (N_1112,N_1063,N_1027);
and U1113 (N_1113,N_1066,N_1075);
or U1114 (N_1114,N_1026,N_1079);
nand U1115 (N_1115,N_1061,N_1066);
nor U1116 (N_1116,N_1021,N_1029);
nor U1117 (N_1117,N_1028,N_1058);
and U1118 (N_1118,N_1041,N_1045);
and U1119 (N_1119,N_1026,N_1043);
and U1120 (N_1120,N_1037,N_1064);
and U1121 (N_1121,N_1051,N_1064);
or U1122 (N_1122,N_1021,N_1068);
and U1123 (N_1123,N_1036,N_1056);
nor U1124 (N_1124,N_1077,N_1079);
and U1125 (N_1125,N_1035,N_1078);
nor U1126 (N_1126,N_1055,N_1030);
and U1127 (N_1127,N_1053,N_1043);
nor U1128 (N_1128,N_1056,N_1058);
nor U1129 (N_1129,N_1061,N_1024);
nand U1130 (N_1130,N_1052,N_1037);
nor U1131 (N_1131,N_1038,N_1051);
or U1132 (N_1132,N_1037,N_1049);
or U1133 (N_1133,N_1062,N_1059);
nand U1134 (N_1134,N_1035,N_1049);
xnor U1135 (N_1135,N_1020,N_1032);
nor U1136 (N_1136,N_1078,N_1020);
nor U1137 (N_1137,N_1060,N_1044);
and U1138 (N_1138,N_1059,N_1022);
or U1139 (N_1139,N_1049,N_1045);
nor U1140 (N_1140,N_1128,N_1102);
nor U1141 (N_1141,N_1090,N_1104);
nand U1142 (N_1142,N_1121,N_1127);
and U1143 (N_1143,N_1089,N_1101);
and U1144 (N_1144,N_1080,N_1135);
nor U1145 (N_1145,N_1130,N_1137);
and U1146 (N_1146,N_1126,N_1098);
nand U1147 (N_1147,N_1113,N_1087);
and U1148 (N_1148,N_1118,N_1133);
nor U1149 (N_1149,N_1112,N_1129);
nand U1150 (N_1150,N_1115,N_1086);
and U1151 (N_1151,N_1119,N_1081);
nor U1152 (N_1152,N_1100,N_1103);
nand U1153 (N_1153,N_1120,N_1094);
or U1154 (N_1154,N_1106,N_1093);
nor U1155 (N_1155,N_1131,N_1116);
nand U1156 (N_1156,N_1107,N_1095);
and U1157 (N_1157,N_1139,N_1123);
nand U1158 (N_1158,N_1136,N_1138);
and U1159 (N_1159,N_1109,N_1134);
nand U1160 (N_1160,N_1117,N_1082);
and U1161 (N_1161,N_1132,N_1110);
or U1162 (N_1162,N_1122,N_1085);
or U1163 (N_1163,N_1097,N_1096);
and U1164 (N_1164,N_1124,N_1092);
nand U1165 (N_1165,N_1088,N_1083);
nor U1166 (N_1166,N_1114,N_1105);
nand U1167 (N_1167,N_1125,N_1099);
or U1168 (N_1168,N_1084,N_1108);
nand U1169 (N_1169,N_1091,N_1111);
nor U1170 (N_1170,N_1123,N_1128);
nand U1171 (N_1171,N_1118,N_1120);
and U1172 (N_1172,N_1103,N_1106);
nand U1173 (N_1173,N_1083,N_1100);
or U1174 (N_1174,N_1105,N_1093);
or U1175 (N_1175,N_1113,N_1101);
or U1176 (N_1176,N_1118,N_1100);
and U1177 (N_1177,N_1110,N_1111);
nor U1178 (N_1178,N_1098,N_1119);
or U1179 (N_1179,N_1134,N_1139);
and U1180 (N_1180,N_1121,N_1108);
and U1181 (N_1181,N_1095,N_1115);
or U1182 (N_1182,N_1090,N_1086);
and U1183 (N_1183,N_1136,N_1131);
or U1184 (N_1184,N_1135,N_1090);
and U1185 (N_1185,N_1117,N_1083);
or U1186 (N_1186,N_1086,N_1111);
nor U1187 (N_1187,N_1095,N_1111);
nand U1188 (N_1188,N_1118,N_1080);
nor U1189 (N_1189,N_1128,N_1089);
and U1190 (N_1190,N_1093,N_1101);
or U1191 (N_1191,N_1125,N_1096);
and U1192 (N_1192,N_1138,N_1097);
and U1193 (N_1193,N_1114,N_1122);
nand U1194 (N_1194,N_1134,N_1138);
nor U1195 (N_1195,N_1094,N_1101);
nand U1196 (N_1196,N_1108,N_1114);
or U1197 (N_1197,N_1125,N_1094);
and U1198 (N_1198,N_1137,N_1122);
nand U1199 (N_1199,N_1126,N_1132);
nor U1200 (N_1200,N_1197,N_1172);
nor U1201 (N_1201,N_1161,N_1191);
xnor U1202 (N_1202,N_1145,N_1152);
nor U1203 (N_1203,N_1144,N_1182);
or U1204 (N_1204,N_1175,N_1187);
nor U1205 (N_1205,N_1190,N_1167);
and U1206 (N_1206,N_1194,N_1165);
nand U1207 (N_1207,N_1147,N_1150);
nor U1208 (N_1208,N_1183,N_1146);
and U1209 (N_1209,N_1174,N_1148);
or U1210 (N_1210,N_1157,N_1184);
nand U1211 (N_1211,N_1192,N_1163);
nor U1212 (N_1212,N_1140,N_1180);
or U1213 (N_1213,N_1160,N_1141);
and U1214 (N_1214,N_1195,N_1189);
nor U1215 (N_1215,N_1171,N_1178);
nor U1216 (N_1216,N_1154,N_1176);
or U1217 (N_1217,N_1158,N_1166);
or U1218 (N_1218,N_1149,N_1181);
nand U1219 (N_1219,N_1155,N_1173);
nand U1220 (N_1220,N_1164,N_1162);
nor U1221 (N_1221,N_1143,N_1170);
xnor U1222 (N_1222,N_1159,N_1142);
or U1223 (N_1223,N_1185,N_1196);
and U1224 (N_1224,N_1193,N_1179);
nand U1225 (N_1225,N_1186,N_1156);
nand U1226 (N_1226,N_1177,N_1199);
or U1227 (N_1227,N_1198,N_1151);
nand U1228 (N_1228,N_1168,N_1169);
nand U1229 (N_1229,N_1188,N_1153);
nand U1230 (N_1230,N_1168,N_1156);
nor U1231 (N_1231,N_1166,N_1177);
and U1232 (N_1232,N_1163,N_1141);
or U1233 (N_1233,N_1162,N_1199);
nand U1234 (N_1234,N_1148,N_1157);
nor U1235 (N_1235,N_1181,N_1182);
nand U1236 (N_1236,N_1180,N_1156);
and U1237 (N_1237,N_1193,N_1199);
nor U1238 (N_1238,N_1185,N_1148);
or U1239 (N_1239,N_1177,N_1167);
and U1240 (N_1240,N_1169,N_1162);
or U1241 (N_1241,N_1154,N_1164);
nand U1242 (N_1242,N_1197,N_1198);
nand U1243 (N_1243,N_1157,N_1155);
or U1244 (N_1244,N_1150,N_1185);
nand U1245 (N_1245,N_1162,N_1180);
and U1246 (N_1246,N_1167,N_1152);
nor U1247 (N_1247,N_1148,N_1159);
nand U1248 (N_1248,N_1169,N_1144);
and U1249 (N_1249,N_1154,N_1196);
or U1250 (N_1250,N_1196,N_1178);
or U1251 (N_1251,N_1171,N_1144);
and U1252 (N_1252,N_1183,N_1177);
nor U1253 (N_1253,N_1199,N_1142);
or U1254 (N_1254,N_1145,N_1149);
nor U1255 (N_1255,N_1183,N_1142);
nor U1256 (N_1256,N_1183,N_1149);
and U1257 (N_1257,N_1167,N_1151);
and U1258 (N_1258,N_1152,N_1162);
nor U1259 (N_1259,N_1195,N_1166);
nor U1260 (N_1260,N_1211,N_1206);
nor U1261 (N_1261,N_1234,N_1201);
and U1262 (N_1262,N_1225,N_1228);
nor U1263 (N_1263,N_1253,N_1243);
nor U1264 (N_1264,N_1241,N_1249);
nor U1265 (N_1265,N_1257,N_1212);
or U1266 (N_1266,N_1240,N_1209);
nand U1267 (N_1267,N_1251,N_1245);
or U1268 (N_1268,N_1219,N_1258);
and U1269 (N_1269,N_1255,N_1256);
or U1270 (N_1270,N_1223,N_1214);
nand U1271 (N_1271,N_1254,N_1230);
and U1272 (N_1272,N_1250,N_1242);
or U1273 (N_1273,N_1218,N_1247);
or U1274 (N_1274,N_1252,N_1221);
or U1275 (N_1275,N_1205,N_1217);
or U1276 (N_1276,N_1244,N_1220);
or U1277 (N_1277,N_1227,N_1213);
nand U1278 (N_1278,N_1235,N_1232);
nand U1279 (N_1279,N_1246,N_1210);
and U1280 (N_1280,N_1204,N_1259);
or U1281 (N_1281,N_1207,N_1215);
or U1282 (N_1282,N_1233,N_1216);
or U1283 (N_1283,N_1229,N_1237);
xor U1284 (N_1284,N_1238,N_1231);
and U1285 (N_1285,N_1203,N_1224);
or U1286 (N_1286,N_1222,N_1248);
nor U1287 (N_1287,N_1202,N_1226);
or U1288 (N_1288,N_1239,N_1200);
nor U1289 (N_1289,N_1208,N_1236);
or U1290 (N_1290,N_1247,N_1237);
nor U1291 (N_1291,N_1256,N_1223);
xnor U1292 (N_1292,N_1213,N_1246);
or U1293 (N_1293,N_1257,N_1224);
or U1294 (N_1294,N_1203,N_1231);
nor U1295 (N_1295,N_1204,N_1200);
nand U1296 (N_1296,N_1226,N_1209);
or U1297 (N_1297,N_1241,N_1245);
and U1298 (N_1298,N_1207,N_1212);
xnor U1299 (N_1299,N_1232,N_1224);
xnor U1300 (N_1300,N_1236,N_1219);
nor U1301 (N_1301,N_1252,N_1219);
nand U1302 (N_1302,N_1252,N_1248);
or U1303 (N_1303,N_1243,N_1216);
nand U1304 (N_1304,N_1244,N_1201);
nor U1305 (N_1305,N_1252,N_1250);
xnor U1306 (N_1306,N_1212,N_1240);
nor U1307 (N_1307,N_1232,N_1208);
nor U1308 (N_1308,N_1255,N_1206);
nand U1309 (N_1309,N_1213,N_1235);
xnor U1310 (N_1310,N_1254,N_1243);
nand U1311 (N_1311,N_1240,N_1224);
nor U1312 (N_1312,N_1206,N_1252);
and U1313 (N_1313,N_1255,N_1240);
nor U1314 (N_1314,N_1250,N_1241);
nand U1315 (N_1315,N_1202,N_1206);
nand U1316 (N_1316,N_1253,N_1223);
or U1317 (N_1317,N_1209,N_1202);
or U1318 (N_1318,N_1222,N_1216);
or U1319 (N_1319,N_1226,N_1215);
and U1320 (N_1320,N_1284,N_1264);
nor U1321 (N_1321,N_1280,N_1265);
or U1322 (N_1322,N_1267,N_1304);
or U1323 (N_1323,N_1281,N_1303);
nor U1324 (N_1324,N_1286,N_1319);
nor U1325 (N_1325,N_1288,N_1294);
and U1326 (N_1326,N_1262,N_1273);
nand U1327 (N_1327,N_1309,N_1275);
and U1328 (N_1328,N_1314,N_1301);
and U1329 (N_1329,N_1299,N_1297);
xnor U1330 (N_1330,N_1261,N_1298);
or U1331 (N_1331,N_1285,N_1306);
nand U1332 (N_1332,N_1310,N_1305);
nor U1333 (N_1333,N_1268,N_1300);
or U1334 (N_1334,N_1276,N_1293);
nor U1335 (N_1335,N_1316,N_1272);
and U1336 (N_1336,N_1274,N_1307);
or U1337 (N_1337,N_1270,N_1308);
or U1338 (N_1338,N_1317,N_1313);
and U1339 (N_1339,N_1269,N_1260);
or U1340 (N_1340,N_1289,N_1291);
xor U1341 (N_1341,N_1266,N_1315);
and U1342 (N_1342,N_1287,N_1312);
nor U1343 (N_1343,N_1283,N_1292);
nor U1344 (N_1344,N_1290,N_1271);
nor U1345 (N_1345,N_1302,N_1318);
and U1346 (N_1346,N_1279,N_1263);
or U1347 (N_1347,N_1277,N_1295);
or U1348 (N_1348,N_1296,N_1278);
xor U1349 (N_1349,N_1282,N_1311);
nor U1350 (N_1350,N_1312,N_1277);
nor U1351 (N_1351,N_1297,N_1276);
and U1352 (N_1352,N_1267,N_1302);
nand U1353 (N_1353,N_1315,N_1276);
nand U1354 (N_1354,N_1299,N_1300);
or U1355 (N_1355,N_1305,N_1307);
nor U1356 (N_1356,N_1317,N_1297);
nand U1357 (N_1357,N_1278,N_1309);
or U1358 (N_1358,N_1298,N_1309);
and U1359 (N_1359,N_1310,N_1276);
nand U1360 (N_1360,N_1285,N_1288);
or U1361 (N_1361,N_1267,N_1300);
nand U1362 (N_1362,N_1291,N_1279);
nor U1363 (N_1363,N_1292,N_1276);
xor U1364 (N_1364,N_1287,N_1267);
and U1365 (N_1365,N_1270,N_1295);
and U1366 (N_1366,N_1265,N_1287);
nand U1367 (N_1367,N_1260,N_1313);
and U1368 (N_1368,N_1293,N_1265);
nor U1369 (N_1369,N_1303,N_1279);
or U1370 (N_1370,N_1264,N_1276);
and U1371 (N_1371,N_1314,N_1268);
nor U1372 (N_1372,N_1270,N_1286);
or U1373 (N_1373,N_1309,N_1285);
and U1374 (N_1374,N_1261,N_1275);
nor U1375 (N_1375,N_1282,N_1286);
and U1376 (N_1376,N_1266,N_1300);
nand U1377 (N_1377,N_1279,N_1315);
nand U1378 (N_1378,N_1295,N_1275);
nor U1379 (N_1379,N_1314,N_1307);
or U1380 (N_1380,N_1338,N_1340);
or U1381 (N_1381,N_1349,N_1333);
or U1382 (N_1382,N_1359,N_1323);
and U1383 (N_1383,N_1344,N_1324);
nand U1384 (N_1384,N_1366,N_1358);
nor U1385 (N_1385,N_1339,N_1336);
nor U1386 (N_1386,N_1357,N_1365);
nand U1387 (N_1387,N_1352,N_1362);
nor U1388 (N_1388,N_1320,N_1375);
and U1389 (N_1389,N_1364,N_1377);
nand U1390 (N_1390,N_1335,N_1343);
nand U1391 (N_1391,N_1329,N_1360);
and U1392 (N_1392,N_1345,N_1361);
and U1393 (N_1393,N_1356,N_1325);
nand U1394 (N_1394,N_1330,N_1371);
or U1395 (N_1395,N_1354,N_1334);
nand U1396 (N_1396,N_1327,N_1372);
or U1397 (N_1397,N_1326,N_1346);
or U1398 (N_1398,N_1348,N_1355);
nor U1399 (N_1399,N_1332,N_1347);
and U1400 (N_1400,N_1322,N_1337);
and U1401 (N_1401,N_1376,N_1321);
and U1402 (N_1402,N_1351,N_1367);
and U1403 (N_1403,N_1368,N_1373);
nor U1404 (N_1404,N_1350,N_1353);
nand U1405 (N_1405,N_1342,N_1331);
and U1406 (N_1406,N_1379,N_1378);
or U1407 (N_1407,N_1341,N_1363);
nor U1408 (N_1408,N_1374,N_1328);
nor U1409 (N_1409,N_1370,N_1369);
nand U1410 (N_1410,N_1371,N_1372);
nand U1411 (N_1411,N_1370,N_1332);
nand U1412 (N_1412,N_1372,N_1344);
nor U1413 (N_1413,N_1357,N_1329);
nor U1414 (N_1414,N_1378,N_1377);
or U1415 (N_1415,N_1334,N_1344);
nor U1416 (N_1416,N_1355,N_1376);
and U1417 (N_1417,N_1370,N_1338);
xnor U1418 (N_1418,N_1373,N_1320);
or U1419 (N_1419,N_1334,N_1374);
and U1420 (N_1420,N_1322,N_1335);
nor U1421 (N_1421,N_1330,N_1353);
nand U1422 (N_1422,N_1363,N_1355);
nand U1423 (N_1423,N_1368,N_1338);
or U1424 (N_1424,N_1367,N_1353);
and U1425 (N_1425,N_1349,N_1321);
nor U1426 (N_1426,N_1320,N_1374);
or U1427 (N_1427,N_1373,N_1362);
nor U1428 (N_1428,N_1321,N_1346);
nand U1429 (N_1429,N_1340,N_1337);
nand U1430 (N_1430,N_1326,N_1335);
nand U1431 (N_1431,N_1365,N_1353);
nor U1432 (N_1432,N_1331,N_1330);
or U1433 (N_1433,N_1325,N_1340);
or U1434 (N_1434,N_1365,N_1329);
nand U1435 (N_1435,N_1353,N_1374);
and U1436 (N_1436,N_1372,N_1347);
or U1437 (N_1437,N_1354,N_1366);
and U1438 (N_1438,N_1336,N_1371);
nor U1439 (N_1439,N_1350,N_1343);
xor U1440 (N_1440,N_1418,N_1419);
nor U1441 (N_1441,N_1411,N_1408);
or U1442 (N_1442,N_1429,N_1393);
or U1443 (N_1443,N_1413,N_1435);
nor U1444 (N_1444,N_1386,N_1415);
and U1445 (N_1445,N_1384,N_1428);
nor U1446 (N_1446,N_1433,N_1438);
nand U1447 (N_1447,N_1398,N_1432);
and U1448 (N_1448,N_1390,N_1405);
and U1449 (N_1449,N_1426,N_1391);
or U1450 (N_1450,N_1427,N_1407);
or U1451 (N_1451,N_1421,N_1431);
and U1452 (N_1452,N_1403,N_1385);
nor U1453 (N_1453,N_1397,N_1401);
or U1454 (N_1454,N_1439,N_1420);
and U1455 (N_1455,N_1388,N_1406);
or U1456 (N_1456,N_1394,N_1399);
nand U1457 (N_1457,N_1404,N_1417);
or U1458 (N_1458,N_1389,N_1412);
and U1459 (N_1459,N_1416,N_1402);
xor U1460 (N_1460,N_1380,N_1424);
or U1461 (N_1461,N_1400,N_1383);
and U1462 (N_1462,N_1382,N_1392);
nor U1463 (N_1463,N_1423,N_1422);
nand U1464 (N_1464,N_1387,N_1396);
nand U1465 (N_1465,N_1434,N_1381);
xor U1466 (N_1466,N_1425,N_1414);
and U1467 (N_1467,N_1409,N_1437);
nor U1468 (N_1468,N_1410,N_1430);
nand U1469 (N_1469,N_1436,N_1395);
or U1470 (N_1470,N_1406,N_1380);
nor U1471 (N_1471,N_1417,N_1380);
nand U1472 (N_1472,N_1408,N_1438);
nor U1473 (N_1473,N_1394,N_1422);
and U1474 (N_1474,N_1408,N_1434);
nand U1475 (N_1475,N_1439,N_1390);
nor U1476 (N_1476,N_1395,N_1432);
nand U1477 (N_1477,N_1413,N_1401);
and U1478 (N_1478,N_1390,N_1418);
or U1479 (N_1479,N_1411,N_1427);
and U1480 (N_1480,N_1389,N_1381);
and U1481 (N_1481,N_1429,N_1409);
nor U1482 (N_1482,N_1390,N_1381);
nor U1483 (N_1483,N_1437,N_1426);
nand U1484 (N_1484,N_1382,N_1399);
xnor U1485 (N_1485,N_1404,N_1386);
or U1486 (N_1486,N_1428,N_1396);
nand U1487 (N_1487,N_1425,N_1388);
nor U1488 (N_1488,N_1409,N_1413);
nand U1489 (N_1489,N_1423,N_1431);
nand U1490 (N_1490,N_1393,N_1416);
and U1491 (N_1491,N_1423,N_1396);
nand U1492 (N_1492,N_1418,N_1422);
nor U1493 (N_1493,N_1420,N_1412);
nor U1494 (N_1494,N_1409,N_1398);
nand U1495 (N_1495,N_1381,N_1416);
and U1496 (N_1496,N_1436,N_1390);
and U1497 (N_1497,N_1395,N_1435);
or U1498 (N_1498,N_1385,N_1422);
and U1499 (N_1499,N_1426,N_1418);
nor U1500 (N_1500,N_1476,N_1486);
or U1501 (N_1501,N_1472,N_1462);
or U1502 (N_1502,N_1453,N_1495);
nor U1503 (N_1503,N_1444,N_1478);
and U1504 (N_1504,N_1487,N_1491);
or U1505 (N_1505,N_1499,N_1442);
nor U1506 (N_1506,N_1443,N_1452);
and U1507 (N_1507,N_1460,N_1498);
or U1508 (N_1508,N_1490,N_1466);
and U1509 (N_1509,N_1441,N_1448);
or U1510 (N_1510,N_1492,N_1479);
nor U1511 (N_1511,N_1473,N_1485);
nor U1512 (N_1512,N_1480,N_1474);
and U1513 (N_1513,N_1481,N_1461);
and U1514 (N_1514,N_1477,N_1464);
and U1515 (N_1515,N_1497,N_1467);
or U1516 (N_1516,N_1446,N_1494);
and U1517 (N_1517,N_1459,N_1493);
or U1518 (N_1518,N_1445,N_1496);
nand U1519 (N_1519,N_1440,N_1468);
or U1520 (N_1520,N_1484,N_1456);
or U1521 (N_1521,N_1449,N_1455);
xor U1522 (N_1522,N_1451,N_1463);
or U1523 (N_1523,N_1471,N_1483);
and U1524 (N_1524,N_1489,N_1488);
nand U1525 (N_1525,N_1457,N_1454);
or U1526 (N_1526,N_1458,N_1469);
and U1527 (N_1527,N_1447,N_1475);
nand U1528 (N_1528,N_1482,N_1450);
and U1529 (N_1529,N_1470,N_1465);
nand U1530 (N_1530,N_1453,N_1496);
nor U1531 (N_1531,N_1468,N_1494);
nor U1532 (N_1532,N_1444,N_1457);
or U1533 (N_1533,N_1475,N_1463);
nor U1534 (N_1534,N_1475,N_1479);
and U1535 (N_1535,N_1449,N_1468);
nand U1536 (N_1536,N_1452,N_1497);
or U1537 (N_1537,N_1485,N_1458);
nand U1538 (N_1538,N_1447,N_1449);
or U1539 (N_1539,N_1456,N_1497);
and U1540 (N_1540,N_1463,N_1483);
nand U1541 (N_1541,N_1461,N_1483);
nand U1542 (N_1542,N_1481,N_1489);
and U1543 (N_1543,N_1471,N_1493);
nor U1544 (N_1544,N_1492,N_1494);
nand U1545 (N_1545,N_1499,N_1467);
nand U1546 (N_1546,N_1440,N_1486);
or U1547 (N_1547,N_1489,N_1445);
nand U1548 (N_1548,N_1459,N_1474);
or U1549 (N_1549,N_1496,N_1447);
nand U1550 (N_1550,N_1498,N_1468);
nor U1551 (N_1551,N_1462,N_1448);
nand U1552 (N_1552,N_1441,N_1494);
and U1553 (N_1553,N_1455,N_1470);
nand U1554 (N_1554,N_1498,N_1461);
or U1555 (N_1555,N_1469,N_1468);
nand U1556 (N_1556,N_1478,N_1497);
nor U1557 (N_1557,N_1482,N_1448);
nand U1558 (N_1558,N_1492,N_1481);
and U1559 (N_1559,N_1483,N_1458);
and U1560 (N_1560,N_1552,N_1533);
or U1561 (N_1561,N_1551,N_1525);
nor U1562 (N_1562,N_1534,N_1542);
nor U1563 (N_1563,N_1500,N_1502);
xnor U1564 (N_1564,N_1557,N_1523);
nor U1565 (N_1565,N_1514,N_1524);
and U1566 (N_1566,N_1540,N_1521);
nand U1567 (N_1567,N_1508,N_1518);
or U1568 (N_1568,N_1555,N_1503);
nand U1569 (N_1569,N_1559,N_1515);
or U1570 (N_1570,N_1535,N_1516);
nor U1571 (N_1571,N_1506,N_1528);
nand U1572 (N_1572,N_1548,N_1550);
or U1573 (N_1573,N_1546,N_1526);
nand U1574 (N_1574,N_1547,N_1544);
or U1575 (N_1575,N_1513,N_1501);
or U1576 (N_1576,N_1531,N_1509);
xnor U1577 (N_1577,N_1549,N_1553);
nor U1578 (N_1578,N_1537,N_1541);
nor U1579 (N_1579,N_1532,N_1527);
nor U1580 (N_1580,N_1530,N_1519);
nand U1581 (N_1581,N_1512,N_1538);
and U1582 (N_1582,N_1545,N_1505);
nor U1583 (N_1583,N_1558,N_1511);
or U1584 (N_1584,N_1543,N_1536);
nor U1585 (N_1585,N_1522,N_1520);
nand U1586 (N_1586,N_1517,N_1510);
and U1587 (N_1587,N_1554,N_1556);
or U1588 (N_1588,N_1539,N_1529);
nor U1589 (N_1589,N_1504,N_1507);
nand U1590 (N_1590,N_1526,N_1549);
or U1591 (N_1591,N_1547,N_1521);
and U1592 (N_1592,N_1542,N_1546);
or U1593 (N_1593,N_1533,N_1530);
nand U1594 (N_1594,N_1557,N_1528);
nor U1595 (N_1595,N_1523,N_1555);
and U1596 (N_1596,N_1502,N_1552);
and U1597 (N_1597,N_1526,N_1551);
nand U1598 (N_1598,N_1500,N_1508);
nor U1599 (N_1599,N_1543,N_1506);
nand U1600 (N_1600,N_1557,N_1522);
nand U1601 (N_1601,N_1525,N_1552);
nor U1602 (N_1602,N_1537,N_1521);
or U1603 (N_1603,N_1543,N_1520);
nor U1604 (N_1604,N_1518,N_1501);
nor U1605 (N_1605,N_1530,N_1507);
nand U1606 (N_1606,N_1543,N_1512);
or U1607 (N_1607,N_1518,N_1511);
nor U1608 (N_1608,N_1551,N_1531);
and U1609 (N_1609,N_1513,N_1539);
nor U1610 (N_1610,N_1531,N_1528);
and U1611 (N_1611,N_1509,N_1557);
or U1612 (N_1612,N_1511,N_1531);
and U1613 (N_1613,N_1506,N_1515);
xnor U1614 (N_1614,N_1511,N_1527);
or U1615 (N_1615,N_1556,N_1536);
nand U1616 (N_1616,N_1513,N_1519);
xnor U1617 (N_1617,N_1510,N_1557);
and U1618 (N_1618,N_1537,N_1553);
nor U1619 (N_1619,N_1510,N_1526);
nand U1620 (N_1620,N_1584,N_1593);
and U1621 (N_1621,N_1579,N_1569);
and U1622 (N_1622,N_1604,N_1608);
nand U1623 (N_1623,N_1601,N_1582);
nand U1624 (N_1624,N_1592,N_1561);
xor U1625 (N_1625,N_1607,N_1591);
nand U1626 (N_1626,N_1586,N_1560);
nor U1627 (N_1627,N_1567,N_1575);
nor U1628 (N_1628,N_1589,N_1619);
nand U1629 (N_1629,N_1603,N_1581);
nand U1630 (N_1630,N_1600,N_1590);
nor U1631 (N_1631,N_1580,N_1606);
and U1632 (N_1632,N_1574,N_1587);
nand U1633 (N_1633,N_1570,N_1596);
and U1634 (N_1634,N_1566,N_1615);
nor U1635 (N_1635,N_1618,N_1599);
or U1636 (N_1636,N_1602,N_1616);
nor U1637 (N_1637,N_1594,N_1598);
nor U1638 (N_1638,N_1585,N_1563);
nand U1639 (N_1639,N_1609,N_1605);
and U1640 (N_1640,N_1613,N_1565);
or U1641 (N_1641,N_1597,N_1583);
nor U1642 (N_1642,N_1562,N_1568);
nand U1643 (N_1643,N_1572,N_1578);
and U1644 (N_1644,N_1571,N_1564);
xor U1645 (N_1645,N_1573,N_1612);
or U1646 (N_1646,N_1577,N_1588);
nor U1647 (N_1647,N_1610,N_1617);
nor U1648 (N_1648,N_1595,N_1576);
nor U1649 (N_1649,N_1611,N_1614);
xor U1650 (N_1650,N_1597,N_1570);
or U1651 (N_1651,N_1598,N_1618);
nand U1652 (N_1652,N_1601,N_1614);
or U1653 (N_1653,N_1573,N_1611);
and U1654 (N_1654,N_1575,N_1618);
or U1655 (N_1655,N_1573,N_1577);
or U1656 (N_1656,N_1560,N_1577);
and U1657 (N_1657,N_1578,N_1580);
nor U1658 (N_1658,N_1602,N_1574);
and U1659 (N_1659,N_1611,N_1561);
or U1660 (N_1660,N_1565,N_1571);
xnor U1661 (N_1661,N_1594,N_1591);
nand U1662 (N_1662,N_1605,N_1579);
nand U1663 (N_1663,N_1619,N_1611);
nand U1664 (N_1664,N_1568,N_1600);
nor U1665 (N_1665,N_1578,N_1605);
nor U1666 (N_1666,N_1585,N_1578);
nor U1667 (N_1667,N_1611,N_1575);
nor U1668 (N_1668,N_1563,N_1613);
nor U1669 (N_1669,N_1606,N_1568);
nand U1670 (N_1670,N_1583,N_1571);
or U1671 (N_1671,N_1609,N_1598);
or U1672 (N_1672,N_1604,N_1598);
and U1673 (N_1673,N_1586,N_1585);
nor U1674 (N_1674,N_1562,N_1565);
and U1675 (N_1675,N_1571,N_1608);
and U1676 (N_1676,N_1599,N_1611);
nor U1677 (N_1677,N_1619,N_1614);
or U1678 (N_1678,N_1607,N_1614);
or U1679 (N_1679,N_1562,N_1614);
nand U1680 (N_1680,N_1633,N_1652);
and U1681 (N_1681,N_1677,N_1625);
nor U1682 (N_1682,N_1662,N_1620);
nand U1683 (N_1683,N_1665,N_1661);
nor U1684 (N_1684,N_1631,N_1657);
nor U1685 (N_1685,N_1674,N_1658);
or U1686 (N_1686,N_1637,N_1668);
nand U1687 (N_1687,N_1653,N_1670);
nor U1688 (N_1688,N_1621,N_1628);
nand U1689 (N_1689,N_1679,N_1654);
and U1690 (N_1690,N_1622,N_1623);
or U1691 (N_1691,N_1647,N_1646);
nand U1692 (N_1692,N_1626,N_1673);
or U1693 (N_1693,N_1663,N_1667);
nand U1694 (N_1694,N_1629,N_1660);
or U1695 (N_1695,N_1678,N_1644);
or U1696 (N_1696,N_1675,N_1635);
nand U1697 (N_1697,N_1638,N_1651);
or U1698 (N_1698,N_1641,N_1645);
nor U1699 (N_1699,N_1642,N_1639);
nor U1700 (N_1700,N_1650,N_1655);
nand U1701 (N_1701,N_1634,N_1636);
nor U1702 (N_1702,N_1649,N_1632);
nor U1703 (N_1703,N_1666,N_1656);
or U1704 (N_1704,N_1671,N_1627);
or U1705 (N_1705,N_1664,N_1630);
nand U1706 (N_1706,N_1643,N_1659);
or U1707 (N_1707,N_1672,N_1669);
nor U1708 (N_1708,N_1676,N_1624);
or U1709 (N_1709,N_1648,N_1640);
or U1710 (N_1710,N_1675,N_1664);
or U1711 (N_1711,N_1660,N_1669);
and U1712 (N_1712,N_1657,N_1665);
nand U1713 (N_1713,N_1622,N_1670);
or U1714 (N_1714,N_1666,N_1675);
nor U1715 (N_1715,N_1670,N_1621);
or U1716 (N_1716,N_1628,N_1659);
nor U1717 (N_1717,N_1654,N_1668);
nor U1718 (N_1718,N_1622,N_1646);
and U1719 (N_1719,N_1661,N_1645);
and U1720 (N_1720,N_1635,N_1666);
or U1721 (N_1721,N_1652,N_1667);
xor U1722 (N_1722,N_1642,N_1643);
and U1723 (N_1723,N_1665,N_1622);
or U1724 (N_1724,N_1632,N_1676);
or U1725 (N_1725,N_1645,N_1652);
and U1726 (N_1726,N_1674,N_1661);
nor U1727 (N_1727,N_1676,N_1645);
nand U1728 (N_1728,N_1637,N_1644);
nand U1729 (N_1729,N_1665,N_1621);
and U1730 (N_1730,N_1641,N_1670);
nand U1731 (N_1731,N_1673,N_1678);
nand U1732 (N_1732,N_1662,N_1675);
nand U1733 (N_1733,N_1638,N_1676);
and U1734 (N_1734,N_1671,N_1648);
nor U1735 (N_1735,N_1624,N_1636);
or U1736 (N_1736,N_1659,N_1663);
nand U1737 (N_1737,N_1654,N_1672);
or U1738 (N_1738,N_1641,N_1658);
nand U1739 (N_1739,N_1679,N_1665);
or U1740 (N_1740,N_1710,N_1706);
or U1741 (N_1741,N_1713,N_1725);
and U1742 (N_1742,N_1727,N_1690);
or U1743 (N_1743,N_1732,N_1693);
nor U1744 (N_1744,N_1684,N_1707);
nor U1745 (N_1745,N_1698,N_1683);
nor U1746 (N_1746,N_1739,N_1685);
nor U1747 (N_1747,N_1724,N_1712);
xnor U1748 (N_1748,N_1682,N_1705);
nand U1749 (N_1749,N_1720,N_1731);
nand U1750 (N_1750,N_1708,N_1704);
nor U1751 (N_1751,N_1715,N_1703);
and U1752 (N_1752,N_1717,N_1692);
nand U1753 (N_1753,N_1700,N_1699);
nand U1754 (N_1754,N_1686,N_1730);
and U1755 (N_1755,N_1733,N_1728);
nand U1756 (N_1756,N_1711,N_1736);
nand U1757 (N_1757,N_1722,N_1735);
or U1758 (N_1758,N_1687,N_1701);
nor U1759 (N_1759,N_1696,N_1695);
nor U1760 (N_1760,N_1737,N_1697);
nand U1761 (N_1761,N_1738,N_1691);
nor U1762 (N_1762,N_1688,N_1723);
nor U1763 (N_1763,N_1702,N_1689);
nor U1764 (N_1764,N_1718,N_1681);
nand U1765 (N_1765,N_1721,N_1716);
or U1766 (N_1766,N_1729,N_1726);
or U1767 (N_1767,N_1734,N_1719);
and U1768 (N_1768,N_1694,N_1714);
nand U1769 (N_1769,N_1709,N_1680);
nand U1770 (N_1770,N_1686,N_1738);
or U1771 (N_1771,N_1723,N_1680);
and U1772 (N_1772,N_1695,N_1702);
or U1773 (N_1773,N_1724,N_1719);
or U1774 (N_1774,N_1715,N_1720);
and U1775 (N_1775,N_1697,N_1693);
and U1776 (N_1776,N_1736,N_1707);
nand U1777 (N_1777,N_1682,N_1687);
nand U1778 (N_1778,N_1689,N_1688);
nand U1779 (N_1779,N_1718,N_1686);
or U1780 (N_1780,N_1688,N_1684);
nor U1781 (N_1781,N_1726,N_1699);
nor U1782 (N_1782,N_1697,N_1707);
and U1783 (N_1783,N_1695,N_1708);
or U1784 (N_1784,N_1706,N_1737);
xnor U1785 (N_1785,N_1716,N_1737);
nand U1786 (N_1786,N_1693,N_1717);
nor U1787 (N_1787,N_1680,N_1697);
or U1788 (N_1788,N_1681,N_1714);
and U1789 (N_1789,N_1707,N_1720);
nand U1790 (N_1790,N_1714,N_1690);
nand U1791 (N_1791,N_1701,N_1697);
and U1792 (N_1792,N_1699,N_1723);
and U1793 (N_1793,N_1705,N_1692);
and U1794 (N_1794,N_1687,N_1685);
or U1795 (N_1795,N_1698,N_1693);
and U1796 (N_1796,N_1705,N_1686);
and U1797 (N_1797,N_1704,N_1738);
nor U1798 (N_1798,N_1720,N_1710);
nand U1799 (N_1799,N_1722,N_1701);
nor U1800 (N_1800,N_1751,N_1765);
nor U1801 (N_1801,N_1757,N_1744);
nand U1802 (N_1802,N_1758,N_1780);
nand U1803 (N_1803,N_1774,N_1793);
nor U1804 (N_1804,N_1770,N_1776);
and U1805 (N_1805,N_1782,N_1768);
nor U1806 (N_1806,N_1779,N_1745);
nand U1807 (N_1807,N_1786,N_1798);
nor U1808 (N_1808,N_1746,N_1748);
or U1809 (N_1809,N_1755,N_1742);
nand U1810 (N_1810,N_1775,N_1781);
nand U1811 (N_1811,N_1771,N_1797);
xor U1812 (N_1812,N_1778,N_1741);
and U1813 (N_1813,N_1749,N_1740);
and U1814 (N_1814,N_1766,N_1762);
or U1815 (N_1815,N_1772,N_1785);
and U1816 (N_1816,N_1799,N_1767);
and U1817 (N_1817,N_1753,N_1752);
or U1818 (N_1818,N_1764,N_1790);
nor U1819 (N_1819,N_1773,N_1796);
nor U1820 (N_1820,N_1777,N_1794);
or U1821 (N_1821,N_1784,N_1792);
and U1822 (N_1822,N_1763,N_1747);
or U1823 (N_1823,N_1791,N_1788);
and U1824 (N_1824,N_1743,N_1750);
nand U1825 (N_1825,N_1756,N_1760);
nor U1826 (N_1826,N_1787,N_1795);
nor U1827 (N_1827,N_1769,N_1783);
and U1828 (N_1828,N_1789,N_1759);
nor U1829 (N_1829,N_1754,N_1761);
nand U1830 (N_1830,N_1742,N_1768);
nand U1831 (N_1831,N_1762,N_1752);
and U1832 (N_1832,N_1772,N_1753);
and U1833 (N_1833,N_1779,N_1751);
and U1834 (N_1834,N_1779,N_1784);
nand U1835 (N_1835,N_1752,N_1776);
or U1836 (N_1836,N_1797,N_1755);
and U1837 (N_1837,N_1752,N_1774);
and U1838 (N_1838,N_1784,N_1764);
nor U1839 (N_1839,N_1772,N_1740);
or U1840 (N_1840,N_1753,N_1776);
or U1841 (N_1841,N_1787,N_1768);
or U1842 (N_1842,N_1779,N_1787);
nor U1843 (N_1843,N_1784,N_1754);
or U1844 (N_1844,N_1783,N_1760);
nor U1845 (N_1845,N_1751,N_1773);
and U1846 (N_1846,N_1744,N_1792);
nor U1847 (N_1847,N_1749,N_1781);
nor U1848 (N_1848,N_1765,N_1766);
and U1849 (N_1849,N_1754,N_1787);
xnor U1850 (N_1850,N_1797,N_1782);
nor U1851 (N_1851,N_1756,N_1796);
or U1852 (N_1852,N_1789,N_1782);
nand U1853 (N_1853,N_1763,N_1797);
nand U1854 (N_1854,N_1769,N_1785);
nor U1855 (N_1855,N_1756,N_1767);
and U1856 (N_1856,N_1784,N_1765);
nor U1857 (N_1857,N_1762,N_1794);
or U1858 (N_1858,N_1792,N_1781);
and U1859 (N_1859,N_1751,N_1767);
or U1860 (N_1860,N_1839,N_1811);
nor U1861 (N_1861,N_1830,N_1804);
nand U1862 (N_1862,N_1803,N_1801);
and U1863 (N_1863,N_1844,N_1824);
and U1864 (N_1864,N_1828,N_1821);
and U1865 (N_1865,N_1826,N_1853);
nor U1866 (N_1866,N_1815,N_1849);
nand U1867 (N_1867,N_1846,N_1800);
nand U1868 (N_1868,N_1838,N_1848);
xor U1869 (N_1869,N_1859,N_1823);
nor U1870 (N_1870,N_1825,N_1837);
and U1871 (N_1871,N_1814,N_1847);
or U1872 (N_1872,N_1845,N_1832);
nor U1873 (N_1873,N_1843,N_1840);
or U1874 (N_1874,N_1808,N_1834);
or U1875 (N_1875,N_1831,N_1802);
and U1876 (N_1876,N_1807,N_1819);
or U1877 (N_1877,N_1851,N_1810);
nand U1878 (N_1878,N_1858,N_1827);
or U1879 (N_1879,N_1835,N_1841);
nand U1880 (N_1880,N_1842,N_1850);
or U1881 (N_1881,N_1820,N_1818);
nor U1882 (N_1882,N_1809,N_1822);
or U1883 (N_1883,N_1854,N_1817);
nor U1884 (N_1884,N_1857,N_1836);
and U1885 (N_1885,N_1852,N_1856);
nor U1886 (N_1886,N_1806,N_1816);
or U1887 (N_1887,N_1812,N_1855);
or U1888 (N_1888,N_1829,N_1805);
nor U1889 (N_1889,N_1833,N_1813);
nor U1890 (N_1890,N_1833,N_1817);
and U1891 (N_1891,N_1831,N_1815);
nand U1892 (N_1892,N_1809,N_1820);
nand U1893 (N_1893,N_1856,N_1807);
nand U1894 (N_1894,N_1859,N_1852);
and U1895 (N_1895,N_1805,N_1843);
and U1896 (N_1896,N_1816,N_1854);
nor U1897 (N_1897,N_1809,N_1856);
nor U1898 (N_1898,N_1844,N_1809);
nand U1899 (N_1899,N_1840,N_1833);
and U1900 (N_1900,N_1859,N_1834);
and U1901 (N_1901,N_1846,N_1815);
nor U1902 (N_1902,N_1845,N_1829);
nand U1903 (N_1903,N_1804,N_1838);
or U1904 (N_1904,N_1803,N_1829);
nor U1905 (N_1905,N_1832,N_1848);
or U1906 (N_1906,N_1841,N_1859);
and U1907 (N_1907,N_1818,N_1852);
nand U1908 (N_1908,N_1829,N_1853);
or U1909 (N_1909,N_1825,N_1854);
or U1910 (N_1910,N_1831,N_1855);
nor U1911 (N_1911,N_1804,N_1837);
nand U1912 (N_1912,N_1806,N_1817);
and U1913 (N_1913,N_1830,N_1827);
and U1914 (N_1914,N_1838,N_1806);
and U1915 (N_1915,N_1854,N_1827);
and U1916 (N_1916,N_1836,N_1849);
or U1917 (N_1917,N_1836,N_1811);
or U1918 (N_1918,N_1843,N_1831);
nor U1919 (N_1919,N_1806,N_1839);
or U1920 (N_1920,N_1881,N_1894);
and U1921 (N_1921,N_1890,N_1883);
nor U1922 (N_1922,N_1867,N_1866);
or U1923 (N_1923,N_1918,N_1860);
nor U1924 (N_1924,N_1863,N_1893);
or U1925 (N_1925,N_1865,N_1898);
nand U1926 (N_1926,N_1864,N_1904);
nand U1927 (N_1927,N_1911,N_1862);
or U1928 (N_1928,N_1875,N_1905);
nand U1929 (N_1929,N_1903,N_1884);
nor U1930 (N_1930,N_1886,N_1878);
nor U1931 (N_1931,N_1917,N_1870);
or U1932 (N_1932,N_1869,N_1914);
nand U1933 (N_1933,N_1888,N_1915);
nor U1934 (N_1934,N_1861,N_1901);
nor U1935 (N_1935,N_1891,N_1913);
and U1936 (N_1936,N_1882,N_1896);
nor U1937 (N_1937,N_1909,N_1907);
nand U1938 (N_1938,N_1895,N_1885);
or U1939 (N_1939,N_1877,N_1876);
and U1940 (N_1940,N_1872,N_1912);
or U1941 (N_1941,N_1889,N_1874);
and U1942 (N_1942,N_1879,N_1910);
nor U1943 (N_1943,N_1892,N_1871);
nand U1944 (N_1944,N_1916,N_1906);
nand U1945 (N_1945,N_1887,N_1873);
nor U1946 (N_1946,N_1880,N_1868);
and U1947 (N_1947,N_1908,N_1897);
and U1948 (N_1948,N_1919,N_1900);
xnor U1949 (N_1949,N_1899,N_1902);
or U1950 (N_1950,N_1863,N_1901);
nor U1951 (N_1951,N_1909,N_1879);
nand U1952 (N_1952,N_1880,N_1876);
or U1953 (N_1953,N_1907,N_1894);
or U1954 (N_1954,N_1911,N_1870);
nand U1955 (N_1955,N_1872,N_1911);
nor U1956 (N_1956,N_1877,N_1914);
or U1957 (N_1957,N_1867,N_1883);
and U1958 (N_1958,N_1902,N_1885);
nor U1959 (N_1959,N_1887,N_1882);
nor U1960 (N_1960,N_1880,N_1862);
nand U1961 (N_1961,N_1886,N_1868);
or U1962 (N_1962,N_1911,N_1892);
nor U1963 (N_1963,N_1878,N_1899);
and U1964 (N_1964,N_1870,N_1905);
or U1965 (N_1965,N_1879,N_1887);
nor U1966 (N_1966,N_1871,N_1867);
or U1967 (N_1967,N_1876,N_1862);
and U1968 (N_1968,N_1870,N_1909);
or U1969 (N_1969,N_1892,N_1917);
or U1970 (N_1970,N_1884,N_1885);
and U1971 (N_1971,N_1901,N_1912);
or U1972 (N_1972,N_1892,N_1909);
nand U1973 (N_1973,N_1883,N_1891);
nor U1974 (N_1974,N_1875,N_1898);
or U1975 (N_1975,N_1919,N_1863);
and U1976 (N_1976,N_1908,N_1909);
or U1977 (N_1977,N_1861,N_1881);
and U1978 (N_1978,N_1870,N_1899);
and U1979 (N_1979,N_1869,N_1880);
nor U1980 (N_1980,N_1979,N_1968);
nor U1981 (N_1981,N_1927,N_1957);
and U1982 (N_1982,N_1921,N_1936);
nand U1983 (N_1983,N_1955,N_1930);
xnor U1984 (N_1984,N_1967,N_1922);
or U1985 (N_1985,N_1975,N_1920);
or U1986 (N_1986,N_1951,N_1932);
or U1987 (N_1987,N_1952,N_1923);
and U1988 (N_1988,N_1933,N_1925);
or U1989 (N_1989,N_1959,N_1966);
or U1990 (N_1990,N_1943,N_1969);
nand U1991 (N_1991,N_1972,N_1953);
nor U1992 (N_1992,N_1940,N_1945);
nand U1993 (N_1993,N_1941,N_1960);
nor U1994 (N_1994,N_1964,N_1947);
nor U1995 (N_1995,N_1944,N_1937);
nor U1996 (N_1996,N_1973,N_1958);
nor U1997 (N_1997,N_1939,N_1946);
nand U1998 (N_1998,N_1950,N_1977);
nand U1999 (N_1999,N_1948,N_1949);
nand U2000 (N_2000,N_1931,N_1954);
nand U2001 (N_2001,N_1978,N_1965);
nand U2002 (N_2002,N_1976,N_1935);
nand U2003 (N_2003,N_1924,N_1942);
nand U2004 (N_2004,N_1962,N_1963);
nor U2005 (N_2005,N_1970,N_1956);
nor U2006 (N_2006,N_1934,N_1926);
nand U2007 (N_2007,N_1928,N_1961);
nor U2008 (N_2008,N_1971,N_1974);
and U2009 (N_2009,N_1938,N_1929);
nand U2010 (N_2010,N_1973,N_1956);
nand U2011 (N_2011,N_1924,N_1966);
nor U2012 (N_2012,N_1923,N_1931);
and U2013 (N_2013,N_1974,N_1934);
nor U2014 (N_2014,N_1951,N_1942);
and U2015 (N_2015,N_1948,N_1974);
and U2016 (N_2016,N_1959,N_1936);
nand U2017 (N_2017,N_1940,N_1972);
and U2018 (N_2018,N_1956,N_1924);
nor U2019 (N_2019,N_1978,N_1941);
or U2020 (N_2020,N_1972,N_1978);
and U2021 (N_2021,N_1978,N_1969);
nor U2022 (N_2022,N_1971,N_1933);
nor U2023 (N_2023,N_1941,N_1921);
nor U2024 (N_2024,N_1956,N_1930);
xnor U2025 (N_2025,N_1973,N_1929);
or U2026 (N_2026,N_1942,N_1948);
nand U2027 (N_2027,N_1956,N_1927);
nor U2028 (N_2028,N_1979,N_1931);
nand U2029 (N_2029,N_1920,N_1933);
and U2030 (N_2030,N_1944,N_1930);
nand U2031 (N_2031,N_1943,N_1933);
and U2032 (N_2032,N_1922,N_1955);
nand U2033 (N_2033,N_1951,N_1958);
or U2034 (N_2034,N_1970,N_1975);
or U2035 (N_2035,N_1960,N_1978);
nand U2036 (N_2036,N_1925,N_1936);
or U2037 (N_2037,N_1925,N_1951);
xor U2038 (N_2038,N_1943,N_1971);
nor U2039 (N_2039,N_1964,N_1965);
and U2040 (N_2040,N_1997,N_2032);
nand U2041 (N_2041,N_2003,N_2005);
and U2042 (N_2042,N_2017,N_1993);
nand U2043 (N_2043,N_2006,N_2038);
and U2044 (N_2044,N_1991,N_2000);
or U2045 (N_2045,N_2008,N_2009);
nor U2046 (N_2046,N_1985,N_2018);
nor U2047 (N_2047,N_2019,N_2015);
nor U2048 (N_2048,N_1992,N_1986);
nor U2049 (N_2049,N_2022,N_2011);
and U2050 (N_2050,N_2027,N_2025);
nand U2051 (N_2051,N_1980,N_1995);
or U2052 (N_2052,N_2035,N_1987);
nand U2053 (N_2053,N_1989,N_1996);
or U2054 (N_2054,N_2004,N_1983);
and U2055 (N_2055,N_2002,N_2016);
or U2056 (N_2056,N_2012,N_2007);
or U2057 (N_2057,N_2020,N_2030);
nor U2058 (N_2058,N_2028,N_2036);
and U2059 (N_2059,N_2033,N_2031);
nand U2060 (N_2060,N_2034,N_1994);
nand U2061 (N_2061,N_1984,N_2010);
or U2062 (N_2062,N_2024,N_2014);
nor U2063 (N_2063,N_1981,N_2001);
or U2064 (N_2064,N_2023,N_2037);
or U2065 (N_2065,N_1999,N_1990);
and U2066 (N_2066,N_1988,N_2013);
and U2067 (N_2067,N_1982,N_2039);
nor U2068 (N_2068,N_2021,N_2026);
or U2069 (N_2069,N_2029,N_1998);
nor U2070 (N_2070,N_2014,N_2005);
nand U2071 (N_2071,N_2027,N_1981);
and U2072 (N_2072,N_1982,N_1998);
nand U2073 (N_2073,N_2018,N_1986);
and U2074 (N_2074,N_2000,N_1992);
nand U2075 (N_2075,N_1989,N_2011);
nor U2076 (N_2076,N_2015,N_1998);
nand U2077 (N_2077,N_2025,N_1986);
nor U2078 (N_2078,N_2008,N_1996);
nor U2079 (N_2079,N_2018,N_2021);
or U2080 (N_2080,N_1999,N_2012);
or U2081 (N_2081,N_2007,N_1996);
and U2082 (N_2082,N_2013,N_2009);
nand U2083 (N_2083,N_2017,N_1996);
nand U2084 (N_2084,N_2029,N_2035);
nand U2085 (N_2085,N_2001,N_1988);
nor U2086 (N_2086,N_1999,N_1987);
nand U2087 (N_2087,N_1981,N_2015);
and U2088 (N_2088,N_2021,N_2031);
and U2089 (N_2089,N_2018,N_2031);
nor U2090 (N_2090,N_2013,N_2039);
nand U2091 (N_2091,N_1993,N_2009);
nand U2092 (N_2092,N_1989,N_2031);
nor U2093 (N_2093,N_1981,N_1995);
and U2094 (N_2094,N_2013,N_2022);
or U2095 (N_2095,N_2009,N_1984);
nand U2096 (N_2096,N_1981,N_1985);
nand U2097 (N_2097,N_2027,N_2037);
nand U2098 (N_2098,N_2000,N_2001);
nor U2099 (N_2099,N_2033,N_1997);
nand U2100 (N_2100,N_2068,N_2043);
and U2101 (N_2101,N_2044,N_2054);
nand U2102 (N_2102,N_2073,N_2098);
and U2103 (N_2103,N_2057,N_2086);
and U2104 (N_2104,N_2091,N_2041);
or U2105 (N_2105,N_2074,N_2046);
nand U2106 (N_2106,N_2081,N_2072);
nor U2107 (N_2107,N_2092,N_2050);
or U2108 (N_2108,N_2067,N_2080);
nor U2109 (N_2109,N_2042,N_2053);
nor U2110 (N_2110,N_2078,N_2052);
and U2111 (N_2111,N_2084,N_2045);
nor U2112 (N_2112,N_2090,N_2060);
nand U2113 (N_2113,N_2055,N_2099);
and U2114 (N_2114,N_2065,N_2096);
or U2115 (N_2115,N_2063,N_2059);
and U2116 (N_2116,N_2082,N_2070);
nand U2117 (N_2117,N_2075,N_2058);
nor U2118 (N_2118,N_2097,N_2089);
nor U2119 (N_2119,N_2069,N_2040);
and U2120 (N_2120,N_2056,N_2061);
nand U2121 (N_2121,N_2047,N_2095);
or U2122 (N_2122,N_2048,N_2093);
nand U2123 (N_2123,N_2066,N_2087);
xor U2124 (N_2124,N_2049,N_2064);
or U2125 (N_2125,N_2079,N_2062);
nand U2126 (N_2126,N_2076,N_2077);
nand U2127 (N_2127,N_2051,N_2083);
or U2128 (N_2128,N_2088,N_2094);
nor U2129 (N_2129,N_2071,N_2085);
and U2130 (N_2130,N_2041,N_2072);
nor U2131 (N_2131,N_2087,N_2060);
nand U2132 (N_2132,N_2081,N_2042);
nor U2133 (N_2133,N_2066,N_2099);
nor U2134 (N_2134,N_2077,N_2073);
and U2135 (N_2135,N_2067,N_2041);
or U2136 (N_2136,N_2042,N_2054);
nor U2137 (N_2137,N_2061,N_2046);
nand U2138 (N_2138,N_2045,N_2096);
and U2139 (N_2139,N_2075,N_2090);
and U2140 (N_2140,N_2093,N_2077);
nor U2141 (N_2141,N_2043,N_2055);
and U2142 (N_2142,N_2092,N_2058);
and U2143 (N_2143,N_2062,N_2042);
nor U2144 (N_2144,N_2084,N_2072);
nand U2145 (N_2145,N_2073,N_2043);
or U2146 (N_2146,N_2055,N_2077);
and U2147 (N_2147,N_2061,N_2047);
nand U2148 (N_2148,N_2096,N_2088);
or U2149 (N_2149,N_2054,N_2091);
and U2150 (N_2150,N_2067,N_2043);
nor U2151 (N_2151,N_2064,N_2092);
and U2152 (N_2152,N_2071,N_2045);
nor U2153 (N_2153,N_2087,N_2054);
and U2154 (N_2154,N_2046,N_2045);
or U2155 (N_2155,N_2083,N_2045);
and U2156 (N_2156,N_2090,N_2047);
xor U2157 (N_2157,N_2077,N_2075);
and U2158 (N_2158,N_2082,N_2099);
and U2159 (N_2159,N_2058,N_2088);
nand U2160 (N_2160,N_2102,N_2148);
or U2161 (N_2161,N_2133,N_2158);
and U2162 (N_2162,N_2104,N_2137);
or U2163 (N_2163,N_2108,N_2125);
nor U2164 (N_2164,N_2115,N_2155);
and U2165 (N_2165,N_2100,N_2149);
and U2166 (N_2166,N_2152,N_2157);
nand U2167 (N_2167,N_2136,N_2109);
and U2168 (N_2168,N_2146,N_2154);
nand U2169 (N_2169,N_2123,N_2121);
nand U2170 (N_2170,N_2111,N_2144);
nand U2171 (N_2171,N_2138,N_2129);
nand U2172 (N_2172,N_2120,N_2106);
xor U2173 (N_2173,N_2122,N_2107);
and U2174 (N_2174,N_2143,N_2110);
nand U2175 (N_2175,N_2130,N_2139);
and U2176 (N_2176,N_2145,N_2140);
and U2177 (N_2177,N_2103,N_2118);
or U2178 (N_2178,N_2142,N_2119);
nor U2179 (N_2179,N_2105,N_2135);
nor U2180 (N_2180,N_2114,N_2126);
nand U2181 (N_2181,N_2159,N_2131);
or U2182 (N_2182,N_2124,N_2132);
and U2183 (N_2183,N_2141,N_2127);
nand U2184 (N_2184,N_2156,N_2150);
or U2185 (N_2185,N_2116,N_2101);
nand U2186 (N_2186,N_2117,N_2128);
xnor U2187 (N_2187,N_2151,N_2134);
or U2188 (N_2188,N_2113,N_2112);
nand U2189 (N_2189,N_2153,N_2147);
nand U2190 (N_2190,N_2130,N_2137);
nand U2191 (N_2191,N_2119,N_2105);
nand U2192 (N_2192,N_2146,N_2151);
nor U2193 (N_2193,N_2124,N_2155);
or U2194 (N_2194,N_2153,N_2132);
nand U2195 (N_2195,N_2108,N_2157);
and U2196 (N_2196,N_2138,N_2134);
nand U2197 (N_2197,N_2144,N_2112);
or U2198 (N_2198,N_2132,N_2129);
nand U2199 (N_2199,N_2147,N_2152);
nand U2200 (N_2200,N_2114,N_2109);
or U2201 (N_2201,N_2121,N_2122);
and U2202 (N_2202,N_2152,N_2101);
nor U2203 (N_2203,N_2146,N_2141);
nand U2204 (N_2204,N_2105,N_2154);
or U2205 (N_2205,N_2148,N_2155);
nand U2206 (N_2206,N_2101,N_2151);
nor U2207 (N_2207,N_2158,N_2108);
nand U2208 (N_2208,N_2135,N_2119);
nor U2209 (N_2209,N_2102,N_2132);
nand U2210 (N_2210,N_2151,N_2133);
or U2211 (N_2211,N_2106,N_2158);
nor U2212 (N_2212,N_2154,N_2113);
nor U2213 (N_2213,N_2114,N_2156);
nand U2214 (N_2214,N_2158,N_2102);
and U2215 (N_2215,N_2104,N_2130);
nand U2216 (N_2216,N_2104,N_2124);
and U2217 (N_2217,N_2125,N_2134);
nand U2218 (N_2218,N_2107,N_2131);
or U2219 (N_2219,N_2125,N_2149);
and U2220 (N_2220,N_2169,N_2185);
and U2221 (N_2221,N_2196,N_2199);
nand U2222 (N_2222,N_2218,N_2174);
nor U2223 (N_2223,N_2160,N_2203);
or U2224 (N_2224,N_2165,N_2194);
or U2225 (N_2225,N_2187,N_2163);
nand U2226 (N_2226,N_2183,N_2167);
and U2227 (N_2227,N_2175,N_2193);
nand U2228 (N_2228,N_2180,N_2200);
and U2229 (N_2229,N_2166,N_2190);
nor U2230 (N_2230,N_2176,N_2164);
nand U2231 (N_2231,N_2195,N_2181);
xnor U2232 (N_2232,N_2209,N_2177);
nand U2233 (N_2233,N_2168,N_2208);
nor U2234 (N_2234,N_2178,N_2179);
nor U2235 (N_2235,N_2205,N_2162);
nand U2236 (N_2236,N_2170,N_2172);
and U2237 (N_2237,N_2219,N_2201);
nand U2238 (N_2238,N_2192,N_2161);
or U2239 (N_2239,N_2204,N_2173);
nand U2240 (N_2240,N_2215,N_2171);
nand U2241 (N_2241,N_2184,N_2214);
or U2242 (N_2242,N_2217,N_2197);
nand U2243 (N_2243,N_2216,N_2189);
and U2244 (N_2244,N_2188,N_2202);
or U2245 (N_2245,N_2213,N_2212);
or U2246 (N_2246,N_2198,N_2210);
nand U2247 (N_2247,N_2186,N_2182);
xnor U2248 (N_2248,N_2207,N_2191);
nor U2249 (N_2249,N_2211,N_2206);
or U2250 (N_2250,N_2201,N_2174);
or U2251 (N_2251,N_2165,N_2161);
nor U2252 (N_2252,N_2213,N_2218);
nor U2253 (N_2253,N_2214,N_2174);
nor U2254 (N_2254,N_2207,N_2215);
and U2255 (N_2255,N_2205,N_2176);
nand U2256 (N_2256,N_2194,N_2186);
or U2257 (N_2257,N_2193,N_2168);
or U2258 (N_2258,N_2191,N_2213);
nand U2259 (N_2259,N_2198,N_2184);
and U2260 (N_2260,N_2214,N_2192);
nor U2261 (N_2261,N_2186,N_2163);
or U2262 (N_2262,N_2183,N_2173);
or U2263 (N_2263,N_2168,N_2169);
nand U2264 (N_2264,N_2173,N_2198);
nand U2265 (N_2265,N_2164,N_2181);
nand U2266 (N_2266,N_2171,N_2217);
nand U2267 (N_2267,N_2219,N_2196);
and U2268 (N_2268,N_2197,N_2191);
or U2269 (N_2269,N_2174,N_2177);
or U2270 (N_2270,N_2193,N_2198);
and U2271 (N_2271,N_2203,N_2215);
or U2272 (N_2272,N_2176,N_2169);
and U2273 (N_2273,N_2169,N_2180);
or U2274 (N_2274,N_2192,N_2212);
or U2275 (N_2275,N_2189,N_2179);
nor U2276 (N_2276,N_2182,N_2207);
or U2277 (N_2277,N_2203,N_2180);
nor U2278 (N_2278,N_2184,N_2188);
nand U2279 (N_2279,N_2213,N_2208);
nor U2280 (N_2280,N_2246,N_2266);
or U2281 (N_2281,N_2254,N_2275);
nor U2282 (N_2282,N_2237,N_2274);
nor U2283 (N_2283,N_2245,N_2240);
or U2284 (N_2284,N_2265,N_2232);
or U2285 (N_2285,N_2220,N_2272);
or U2286 (N_2286,N_2277,N_2263);
and U2287 (N_2287,N_2270,N_2231);
nand U2288 (N_2288,N_2248,N_2269);
nand U2289 (N_2289,N_2271,N_2243);
and U2290 (N_2290,N_2257,N_2258);
nand U2291 (N_2291,N_2227,N_2255);
and U2292 (N_2292,N_2250,N_2236);
and U2293 (N_2293,N_2242,N_2268);
nor U2294 (N_2294,N_2259,N_2221);
and U2295 (N_2295,N_2224,N_2230);
or U2296 (N_2296,N_2226,N_2239);
or U2297 (N_2297,N_2238,N_2249);
nand U2298 (N_2298,N_2244,N_2234);
nand U2299 (N_2299,N_2273,N_2225);
or U2300 (N_2300,N_2247,N_2260);
nor U2301 (N_2301,N_2222,N_2262);
or U2302 (N_2302,N_2251,N_2229);
nand U2303 (N_2303,N_2223,N_2235);
nand U2304 (N_2304,N_2267,N_2233);
or U2305 (N_2305,N_2278,N_2276);
nand U2306 (N_2306,N_2241,N_2261);
nand U2307 (N_2307,N_2264,N_2256);
and U2308 (N_2308,N_2252,N_2253);
and U2309 (N_2309,N_2228,N_2279);
nor U2310 (N_2310,N_2242,N_2257);
and U2311 (N_2311,N_2258,N_2263);
nand U2312 (N_2312,N_2251,N_2224);
nand U2313 (N_2313,N_2230,N_2229);
and U2314 (N_2314,N_2251,N_2268);
and U2315 (N_2315,N_2258,N_2222);
or U2316 (N_2316,N_2249,N_2272);
nand U2317 (N_2317,N_2245,N_2264);
or U2318 (N_2318,N_2222,N_2247);
and U2319 (N_2319,N_2251,N_2232);
nand U2320 (N_2320,N_2264,N_2271);
nand U2321 (N_2321,N_2224,N_2276);
or U2322 (N_2322,N_2270,N_2242);
nor U2323 (N_2323,N_2230,N_2278);
or U2324 (N_2324,N_2221,N_2265);
or U2325 (N_2325,N_2229,N_2258);
and U2326 (N_2326,N_2245,N_2263);
and U2327 (N_2327,N_2276,N_2251);
and U2328 (N_2328,N_2233,N_2222);
or U2329 (N_2329,N_2252,N_2237);
nor U2330 (N_2330,N_2258,N_2244);
or U2331 (N_2331,N_2279,N_2271);
nand U2332 (N_2332,N_2256,N_2235);
or U2333 (N_2333,N_2238,N_2276);
or U2334 (N_2334,N_2253,N_2229);
and U2335 (N_2335,N_2242,N_2243);
nand U2336 (N_2336,N_2267,N_2222);
and U2337 (N_2337,N_2231,N_2239);
nand U2338 (N_2338,N_2274,N_2275);
nand U2339 (N_2339,N_2262,N_2234);
or U2340 (N_2340,N_2308,N_2320);
or U2341 (N_2341,N_2287,N_2292);
nor U2342 (N_2342,N_2326,N_2317);
and U2343 (N_2343,N_2296,N_2337);
nor U2344 (N_2344,N_2303,N_2289);
or U2345 (N_2345,N_2290,N_2325);
nand U2346 (N_2346,N_2305,N_2310);
nand U2347 (N_2347,N_2314,N_2284);
nand U2348 (N_2348,N_2313,N_2307);
nand U2349 (N_2349,N_2298,N_2283);
and U2350 (N_2350,N_2309,N_2286);
nand U2351 (N_2351,N_2329,N_2335);
nor U2352 (N_2352,N_2301,N_2333);
or U2353 (N_2353,N_2306,N_2280);
and U2354 (N_2354,N_2318,N_2316);
nand U2355 (N_2355,N_2281,N_2300);
and U2356 (N_2356,N_2299,N_2330);
nor U2357 (N_2357,N_2327,N_2338);
and U2358 (N_2358,N_2332,N_2288);
or U2359 (N_2359,N_2282,N_2323);
nand U2360 (N_2360,N_2294,N_2302);
nand U2361 (N_2361,N_2339,N_2334);
and U2362 (N_2362,N_2336,N_2319);
or U2363 (N_2363,N_2321,N_2324);
nor U2364 (N_2364,N_2293,N_2285);
nor U2365 (N_2365,N_2295,N_2311);
or U2366 (N_2366,N_2315,N_2291);
nor U2367 (N_2367,N_2297,N_2304);
nand U2368 (N_2368,N_2328,N_2312);
nor U2369 (N_2369,N_2322,N_2331);
or U2370 (N_2370,N_2310,N_2287);
nand U2371 (N_2371,N_2286,N_2308);
nor U2372 (N_2372,N_2299,N_2324);
and U2373 (N_2373,N_2292,N_2298);
nor U2374 (N_2374,N_2318,N_2281);
nand U2375 (N_2375,N_2313,N_2328);
and U2376 (N_2376,N_2320,N_2281);
nand U2377 (N_2377,N_2334,N_2282);
nor U2378 (N_2378,N_2319,N_2291);
and U2379 (N_2379,N_2304,N_2332);
nor U2380 (N_2380,N_2285,N_2333);
or U2381 (N_2381,N_2329,N_2309);
nor U2382 (N_2382,N_2286,N_2293);
nor U2383 (N_2383,N_2297,N_2329);
nor U2384 (N_2384,N_2330,N_2339);
and U2385 (N_2385,N_2310,N_2338);
nand U2386 (N_2386,N_2327,N_2318);
and U2387 (N_2387,N_2300,N_2298);
nand U2388 (N_2388,N_2336,N_2332);
nand U2389 (N_2389,N_2318,N_2284);
nor U2390 (N_2390,N_2300,N_2287);
nand U2391 (N_2391,N_2289,N_2290);
nor U2392 (N_2392,N_2325,N_2294);
and U2393 (N_2393,N_2325,N_2326);
xnor U2394 (N_2394,N_2323,N_2289);
or U2395 (N_2395,N_2337,N_2308);
or U2396 (N_2396,N_2307,N_2286);
or U2397 (N_2397,N_2280,N_2294);
nand U2398 (N_2398,N_2305,N_2295);
nand U2399 (N_2399,N_2330,N_2302);
or U2400 (N_2400,N_2342,N_2347);
nand U2401 (N_2401,N_2376,N_2393);
nand U2402 (N_2402,N_2389,N_2348);
or U2403 (N_2403,N_2354,N_2363);
nand U2404 (N_2404,N_2399,N_2367);
or U2405 (N_2405,N_2381,N_2359);
and U2406 (N_2406,N_2378,N_2371);
nand U2407 (N_2407,N_2386,N_2375);
and U2408 (N_2408,N_2358,N_2346);
nor U2409 (N_2409,N_2349,N_2361);
and U2410 (N_2410,N_2351,N_2385);
nand U2411 (N_2411,N_2341,N_2366);
nand U2412 (N_2412,N_2382,N_2365);
nand U2413 (N_2413,N_2340,N_2350);
nand U2414 (N_2414,N_2391,N_2395);
or U2415 (N_2415,N_2369,N_2352);
nor U2416 (N_2416,N_2380,N_2343);
or U2417 (N_2417,N_2357,N_2394);
nand U2418 (N_2418,N_2374,N_2383);
nor U2419 (N_2419,N_2390,N_2398);
nor U2420 (N_2420,N_2345,N_2373);
and U2421 (N_2421,N_2397,N_2387);
nand U2422 (N_2422,N_2379,N_2364);
and U2423 (N_2423,N_2356,N_2353);
and U2424 (N_2424,N_2372,N_2362);
and U2425 (N_2425,N_2368,N_2355);
or U2426 (N_2426,N_2388,N_2370);
or U2427 (N_2427,N_2377,N_2396);
nand U2428 (N_2428,N_2360,N_2392);
nor U2429 (N_2429,N_2384,N_2344);
or U2430 (N_2430,N_2392,N_2394);
and U2431 (N_2431,N_2394,N_2379);
nand U2432 (N_2432,N_2392,N_2370);
nor U2433 (N_2433,N_2386,N_2378);
or U2434 (N_2434,N_2374,N_2349);
and U2435 (N_2435,N_2390,N_2373);
or U2436 (N_2436,N_2391,N_2384);
nand U2437 (N_2437,N_2372,N_2384);
or U2438 (N_2438,N_2352,N_2373);
nor U2439 (N_2439,N_2396,N_2342);
or U2440 (N_2440,N_2359,N_2398);
and U2441 (N_2441,N_2384,N_2382);
or U2442 (N_2442,N_2357,N_2369);
and U2443 (N_2443,N_2370,N_2382);
nand U2444 (N_2444,N_2374,N_2360);
or U2445 (N_2445,N_2352,N_2368);
or U2446 (N_2446,N_2367,N_2371);
and U2447 (N_2447,N_2359,N_2345);
or U2448 (N_2448,N_2355,N_2386);
and U2449 (N_2449,N_2352,N_2340);
nand U2450 (N_2450,N_2381,N_2393);
nor U2451 (N_2451,N_2382,N_2352);
nand U2452 (N_2452,N_2371,N_2397);
nand U2453 (N_2453,N_2399,N_2358);
or U2454 (N_2454,N_2353,N_2347);
and U2455 (N_2455,N_2354,N_2392);
nor U2456 (N_2456,N_2377,N_2374);
nor U2457 (N_2457,N_2378,N_2388);
nor U2458 (N_2458,N_2389,N_2379);
nor U2459 (N_2459,N_2352,N_2342);
nand U2460 (N_2460,N_2416,N_2413);
and U2461 (N_2461,N_2425,N_2448);
or U2462 (N_2462,N_2419,N_2433);
xor U2463 (N_2463,N_2430,N_2451);
nor U2464 (N_2464,N_2410,N_2440);
nor U2465 (N_2465,N_2421,N_2459);
nor U2466 (N_2466,N_2449,N_2428);
nand U2467 (N_2467,N_2408,N_2434);
nor U2468 (N_2468,N_2450,N_2402);
nor U2469 (N_2469,N_2457,N_2422);
or U2470 (N_2470,N_2444,N_2417);
or U2471 (N_2471,N_2405,N_2426);
nand U2472 (N_2472,N_2435,N_2407);
nand U2473 (N_2473,N_2412,N_2438);
or U2474 (N_2474,N_2411,N_2420);
nor U2475 (N_2475,N_2453,N_2455);
nor U2476 (N_2476,N_2406,N_2404);
and U2477 (N_2477,N_2447,N_2403);
and U2478 (N_2478,N_2418,N_2414);
or U2479 (N_2479,N_2443,N_2401);
xor U2480 (N_2480,N_2442,N_2439);
or U2481 (N_2481,N_2454,N_2441);
nor U2482 (N_2482,N_2458,N_2432);
and U2483 (N_2483,N_2409,N_2431);
nor U2484 (N_2484,N_2445,N_2429);
and U2485 (N_2485,N_2437,N_2456);
or U2486 (N_2486,N_2415,N_2427);
nor U2487 (N_2487,N_2436,N_2452);
and U2488 (N_2488,N_2424,N_2446);
nor U2489 (N_2489,N_2400,N_2423);
and U2490 (N_2490,N_2439,N_2413);
nand U2491 (N_2491,N_2401,N_2432);
or U2492 (N_2492,N_2450,N_2438);
nor U2493 (N_2493,N_2411,N_2409);
or U2494 (N_2494,N_2451,N_2406);
or U2495 (N_2495,N_2418,N_2441);
nor U2496 (N_2496,N_2433,N_2440);
or U2497 (N_2497,N_2401,N_2415);
nor U2498 (N_2498,N_2432,N_2445);
or U2499 (N_2499,N_2447,N_2428);
nor U2500 (N_2500,N_2439,N_2424);
nor U2501 (N_2501,N_2446,N_2409);
nand U2502 (N_2502,N_2434,N_2420);
and U2503 (N_2503,N_2425,N_2410);
or U2504 (N_2504,N_2420,N_2446);
nand U2505 (N_2505,N_2441,N_2449);
nand U2506 (N_2506,N_2452,N_2426);
nand U2507 (N_2507,N_2431,N_2439);
or U2508 (N_2508,N_2419,N_2455);
nand U2509 (N_2509,N_2421,N_2415);
nand U2510 (N_2510,N_2436,N_2432);
or U2511 (N_2511,N_2448,N_2456);
and U2512 (N_2512,N_2421,N_2454);
or U2513 (N_2513,N_2444,N_2410);
nor U2514 (N_2514,N_2457,N_2400);
and U2515 (N_2515,N_2426,N_2413);
nand U2516 (N_2516,N_2410,N_2420);
nor U2517 (N_2517,N_2420,N_2432);
nand U2518 (N_2518,N_2430,N_2452);
nand U2519 (N_2519,N_2401,N_2404);
nor U2520 (N_2520,N_2482,N_2477);
or U2521 (N_2521,N_2476,N_2512);
nand U2522 (N_2522,N_2499,N_2465);
nand U2523 (N_2523,N_2508,N_2469);
nor U2524 (N_2524,N_2474,N_2488);
nor U2525 (N_2525,N_2489,N_2496);
nor U2526 (N_2526,N_2509,N_2467);
and U2527 (N_2527,N_2507,N_2494);
nor U2528 (N_2528,N_2514,N_2513);
nor U2529 (N_2529,N_2492,N_2478);
or U2530 (N_2530,N_2519,N_2511);
and U2531 (N_2531,N_2461,N_2466);
nor U2532 (N_2532,N_2485,N_2502);
nor U2533 (N_2533,N_2503,N_2515);
or U2534 (N_2534,N_2464,N_2497);
nand U2535 (N_2535,N_2475,N_2491);
nand U2536 (N_2536,N_2483,N_2463);
or U2537 (N_2537,N_2498,N_2479);
and U2538 (N_2538,N_2495,N_2470);
and U2539 (N_2539,N_2472,N_2501);
or U2540 (N_2540,N_2462,N_2517);
and U2541 (N_2541,N_2468,N_2471);
nand U2542 (N_2542,N_2487,N_2500);
nand U2543 (N_2543,N_2460,N_2486);
nor U2544 (N_2544,N_2504,N_2518);
and U2545 (N_2545,N_2481,N_2484);
nand U2546 (N_2546,N_2506,N_2516);
and U2547 (N_2547,N_2493,N_2473);
nor U2548 (N_2548,N_2490,N_2480);
or U2549 (N_2549,N_2505,N_2510);
nor U2550 (N_2550,N_2466,N_2479);
and U2551 (N_2551,N_2497,N_2482);
nor U2552 (N_2552,N_2517,N_2495);
nor U2553 (N_2553,N_2500,N_2472);
nor U2554 (N_2554,N_2509,N_2518);
or U2555 (N_2555,N_2516,N_2507);
or U2556 (N_2556,N_2509,N_2478);
and U2557 (N_2557,N_2501,N_2510);
or U2558 (N_2558,N_2508,N_2519);
nor U2559 (N_2559,N_2518,N_2516);
xnor U2560 (N_2560,N_2487,N_2513);
nand U2561 (N_2561,N_2484,N_2501);
nand U2562 (N_2562,N_2460,N_2477);
nand U2563 (N_2563,N_2493,N_2484);
and U2564 (N_2564,N_2518,N_2513);
and U2565 (N_2565,N_2488,N_2506);
and U2566 (N_2566,N_2489,N_2516);
and U2567 (N_2567,N_2474,N_2501);
and U2568 (N_2568,N_2481,N_2507);
nor U2569 (N_2569,N_2515,N_2471);
or U2570 (N_2570,N_2487,N_2480);
and U2571 (N_2571,N_2483,N_2502);
nor U2572 (N_2572,N_2473,N_2468);
nor U2573 (N_2573,N_2509,N_2490);
or U2574 (N_2574,N_2512,N_2518);
nand U2575 (N_2575,N_2511,N_2516);
and U2576 (N_2576,N_2461,N_2474);
or U2577 (N_2577,N_2467,N_2496);
nand U2578 (N_2578,N_2472,N_2510);
nor U2579 (N_2579,N_2511,N_2515);
nand U2580 (N_2580,N_2573,N_2570);
nand U2581 (N_2581,N_2553,N_2564);
or U2582 (N_2582,N_2537,N_2531);
nor U2583 (N_2583,N_2577,N_2526);
or U2584 (N_2584,N_2566,N_2550);
or U2585 (N_2585,N_2528,N_2532);
or U2586 (N_2586,N_2554,N_2574);
or U2587 (N_2587,N_2562,N_2540);
and U2588 (N_2588,N_2545,N_2567);
nand U2589 (N_2589,N_2552,N_2578);
or U2590 (N_2590,N_2558,N_2575);
nor U2591 (N_2591,N_2547,N_2521);
nor U2592 (N_2592,N_2534,N_2576);
and U2593 (N_2593,N_2565,N_2525);
or U2594 (N_2594,N_2546,N_2569);
nor U2595 (N_2595,N_2530,N_2563);
or U2596 (N_2596,N_2538,N_2559);
and U2597 (N_2597,N_2527,N_2541);
and U2598 (N_2598,N_2539,N_2542);
or U2599 (N_2599,N_2557,N_2522);
nand U2600 (N_2600,N_2520,N_2544);
or U2601 (N_2601,N_2549,N_2572);
nand U2602 (N_2602,N_2523,N_2579);
nand U2603 (N_2603,N_2533,N_2536);
nand U2604 (N_2604,N_2535,N_2555);
nand U2605 (N_2605,N_2529,N_2568);
and U2606 (N_2606,N_2543,N_2560);
nand U2607 (N_2607,N_2556,N_2571);
and U2608 (N_2608,N_2548,N_2551);
nor U2609 (N_2609,N_2524,N_2561);
nand U2610 (N_2610,N_2578,N_2542);
nand U2611 (N_2611,N_2538,N_2553);
nand U2612 (N_2612,N_2558,N_2549);
nand U2613 (N_2613,N_2532,N_2568);
or U2614 (N_2614,N_2551,N_2534);
and U2615 (N_2615,N_2570,N_2535);
nor U2616 (N_2616,N_2533,N_2527);
xnor U2617 (N_2617,N_2573,N_2575);
or U2618 (N_2618,N_2555,N_2576);
xor U2619 (N_2619,N_2578,N_2549);
or U2620 (N_2620,N_2546,N_2527);
nor U2621 (N_2621,N_2528,N_2559);
nor U2622 (N_2622,N_2531,N_2540);
or U2623 (N_2623,N_2571,N_2553);
or U2624 (N_2624,N_2542,N_2529);
nand U2625 (N_2625,N_2564,N_2558);
or U2626 (N_2626,N_2547,N_2573);
and U2627 (N_2627,N_2543,N_2555);
nand U2628 (N_2628,N_2562,N_2559);
nand U2629 (N_2629,N_2531,N_2534);
nor U2630 (N_2630,N_2569,N_2527);
nor U2631 (N_2631,N_2565,N_2548);
nand U2632 (N_2632,N_2559,N_2550);
nor U2633 (N_2633,N_2575,N_2523);
nor U2634 (N_2634,N_2552,N_2572);
and U2635 (N_2635,N_2521,N_2568);
nand U2636 (N_2636,N_2544,N_2526);
or U2637 (N_2637,N_2556,N_2566);
and U2638 (N_2638,N_2538,N_2562);
and U2639 (N_2639,N_2540,N_2573);
or U2640 (N_2640,N_2581,N_2599);
and U2641 (N_2641,N_2629,N_2625);
or U2642 (N_2642,N_2606,N_2594);
or U2643 (N_2643,N_2603,N_2591);
nand U2644 (N_2644,N_2628,N_2602);
and U2645 (N_2645,N_2635,N_2639);
and U2646 (N_2646,N_2612,N_2634);
nand U2647 (N_2647,N_2585,N_2632);
nand U2648 (N_2648,N_2589,N_2621);
or U2649 (N_2649,N_2609,N_2618);
nand U2650 (N_2650,N_2631,N_2611);
or U2651 (N_2651,N_2608,N_2584);
or U2652 (N_2652,N_2590,N_2601);
nor U2653 (N_2653,N_2583,N_2624);
and U2654 (N_2654,N_2595,N_2638);
nand U2655 (N_2655,N_2592,N_2613);
nor U2656 (N_2656,N_2622,N_2626);
nand U2657 (N_2657,N_2586,N_2614);
nand U2658 (N_2658,N_2620,N_2582);
and U2659 (N_2659,N_2616,N_2600);
nand U2660 (N_2660,N_2607,N_2637);
nand U2661 (N_2661,N_2617,N_2610);
nor U2662 (N_2662,N_2605,N_2587);
nor U2663 (N_2663,N_2580,N_2596);
and U2664 (N_2664,N_2627,N_2636);
and U2665 (N_2665,N_2615,N_2623);
and U2666 (N_2666,N_2598,N_2588);
nor U2667 (N_2667,N_2630,N_2593);
and U2668 (N_2668,N_2597,N_2604);
or U2669 (N_2669,N_2633,N_2619);
nor U2670 (N_2670,N_2619,N_2614);
or U2671 (N_2671,N_2639,N_2583);
nor U2672 (N_2672,N_2586,N_2602);
or U2673 (N_2673,N_2635,N_2627);
and U2674 (N_2674,N_2634,N_2630);
and U2675 (N_2675,N_2621,N_2618);
and U2676 (N_2676,N_2638,N_2587);
nor U2677 (N_2677,N_2621,N_2639);
or U2678 (N_2678,N_2625,N_2638);
and U2679 (N_2679,N_2623,N_2585);
xnor U2680 (N_2680,N_2639,N_2631);
nor U2681 (N_2681,N_2602,N_2634);
nor U2682 (N_2682,N_2602,N_2589);
or U2683 (N_2683,N_2614,N_2604);
nor U2684 (N_2684,N_2587,N_2597);
xnor U2685 (N_2685,N_2588,N_2613);
or U2686 (N_2686,N_2623,N_2606);
nor U2687 (N_2687,N_2596,N_2602);
nor U2688 (N_2688,N_2580,N_2612);
or U2689 (N_2689,N_2611,N_2581);
nor U2690 (N_2690,N_2616,N_2623);
and U2691 (N_2691,N_2611,N_2601);
or U2692 (N_2692,N_2611,N_2634);
or U2693 (N_2693,N_2637,N_2595);
nand U2694 (N_2694,N_2600,N_2597);
nor U2695 (N_2695,N_2607,N_2624);
and U2696 (N_2696,N_2637,N_2625);
nand U2697 (N_2697,N_2615,N_2605);
nand U2698 (N_2698,N_2596,N_2593);
and U2699 (N_2699,N_2611,N_2614);
nand U2700 (N_2700,N_2651,N_2666);
or U2701 (N_2701,N_2660,N_2691);
and U2702 (N_2702,N_2648,N_2679);
and U2703 (N_2703,N_2699,N_2680);
and U2704 (N_2704,N_2655,N_2658);
and U2705 (N_2705,N_2698,N_2692);
nand U2706 (N_2706,N_2675,N_2672);
or U2707 (N_2707,N_2656,N_2644);
and U2708 (N_2708,N_2650,N_2677);
or U2709 (N_2709,N_2682,N_2649);
nand U2710 (N_2710,N_2684,N_2678);
or U2711 (N_2711,N_2686,N_2657);
nand U2712 (N_2712,N_2654,N_2653);
nand U2713 (N_2713,N_2674,N_2667);
and U2714 (N_2714,N_2643,N_2670);
nand U2715 (N_2715,N_2673,N_2665);
and U2716 (N_2716,N_2695,N_2676);
nand U2717 (N_2717,N_2659,N_2669);
nor U2718 (N_2718,N_2652,N_2697);
nand U2719 (N_2719,N_2641,N_2640);
or U2720 (N_2720,N_2662,N_2646);
and U2721 (N_2721,N_2689,N_2664);
nor U2722 (N_2722,N_2668,N_2685);
nor U2723 (N_2723,N_2681,N_2688);
or U2724 (N_2724,N_2693,N_2647);
nor U2725 (N_2725,N_2694,N_2683);
and U2726 (N_2726,N_2663,N_2696);
or U2727 (N_2727,N_2642,N_2661);
nand U2728 (N_2728,N_2645,N_2687);
and U2729 (N_2729,N_2671,N_2690);
nor U2730 (N_2730,N_2681,N_2671);
and U2731 (N_2731,N_2655,N_2645);
or U2732 (N_2732,N_2660,N_2661);
nor U2733 (N_2733,N_2679,N_2678);
nor U2734 (N_2734,N_2680,N_2681);
or U2735 (N_2735,N_2657,N_2695);
or U2736 (N_2736,N_2685,N_2674);
nor U2737 (N_2737,N_2665,N_2651);
or U2738 (N_2738,N_2644,N_2669);
and U2739 (N_2739,N_2657,N_2673);
or U2740 (N_2740,N_2670,N_2695);
or U2741 (N_2741,N_2693,N_2644);
and U2742 (N_2742,N_2681,N_2664);
nand U2743 (N_2743,N_2662,N_2684);
xnor U2744 (N_2744,N_2647,N_2681);
or U2745 (N_2745,N_2698,N_2689);
nand U2746 (N_2746,N_2680,N_2696);
nand U2747 (N_2747,N_2695,N_2683);
or U2748 (N_2748,N_2677,N_2691);
and U2749 (N_2749,N_2676,N_2678);
nand U2750 (N_2750,N_2675,N_2679);
nand U2751 (N_2751,N_2663,N_2682);
or U2752 (N_2752,N_2679,N_2684);
and U2753 (N_2753,N_2657,N_2648);
nor U2754 (N_2754,N_2645,N_2665);
xnor U2755 (N_2755,N_2671,N_2655);
nand U2756 (N_2756,N_2680,N_2666);
or U2757 (N_2757,N_2658,N_2691);
nor U2758 (N_2758,N_2657,N_2693);
or U2759 (N_2759,N_2679,N_2685);
nor U2760 (N_2760,N_2752,N_2744);
or U2761 (N_2761,N_2726,N_2728);
or U2762 (N_2762,N_2754,N_2715);
and U2763 (N_2763,N_2722,N_2733);
or U2764 (N_2764,N_2741,N_2713);
nor U2765 (N_2765,N_2743,N_2756);
nand U2766 (N_2766,N_2706,N_2723);
nand U2767 (N_2767,N_2740,N_2748);
nor U2768 (N_2768,N_2700,N_2757);
nor U2769 (N_2769,N_2710,N_2711);
or U2770 (N_2770,N_2758,N_2735);
nor U2771 (N_2771,N_2750,N_2701);
and U2772 (N_2772,N_2705,N_2717);
nand U2773 (N_2773,N_2753,N_2719);
nor U2774 (N_2774,N_2747,N_2720);
or U2775 (N_2775,N_2751,N_2745);
nand U2776 (N_2776,N_2746,N_2725);
and U2777 (N_2777,N_2704,N_2724);
nand U2778 (N_2778,N_2739,N_2718);
nand U2779 (N_2779,N_2703,N_2731);
or U2780 (N_2780,N_2755,N_2707);
or U2781 (N_2781,N_2709,N_2759);
or U2782 (N_2782,N_2730,N_2712);
xnor U2783 (N_2783,N_2702,N_2714);
nand U2784 (N_2784,N_2736,N_2742);
nand U2785 (N_2785,N_2727,N_2734);
or U2786 (N_2786,N_2737,N_2729);
nand U2787 (N_2787,N_2738,N_2732);
nand U2788 (N_2788,N_2721,N_2749);
nor U2789 (N_2789,N_2708,N_2716);
and U2790 (N_2790,N_2738,N_2729);
nor U2791 (N_2791,N_2735,N_2717);
nand U2792 (N_2792,N_2711,N_2732);
nor U2793 (N_2793,N_2708,N_2756);
nor U2794 (N_2794,N_2750,N_2735);
or U2795 (N_2795,N_2727,N_2755);
or U2796 (N_2796,N_2720,N_2730);
and U2797 (N_2797,N_2737,N_2747);
and U2798 (N_2798,N_2746,N_2754);
and U2799 (N_2799,N_2754,N_2731);
nor U2800 (N_2800,N_2728,N_2737);
nand U2801 (N_2801,N_2757,N_2735);
nand U2802 (N_2802,N_2737,N_2756);
nor U2803 (N_2803,N_2752,N_2720);
or U2804 (N_2804,N_2741,N_2755);
or U2805 (N_2805,N_2716,N_2723);
nor U2806 (N_2806,N_2744,N_2738);
nand U2807 (N_2807,N_2734,N_2716);
nand U2808 (N_2808,N_2744,N_2721);
and U2809 (N_2809,N_2757,N_2738);
nor U2810 (N_2810,N_2719,N_2715);
or U2811 (N_2811,N_2743,N_2725);
nor U2812 (N_2812,N_2716,N_2707);
nor U2813 (N_2813,N_2725,N_2710);
or U2814 (N_2814,N_2730,N_2700);
nor U2815 (N_2815,N_2711,N_2756);
and U2816 (N_2816,N_2700,N_2758);
or U2817 (N_2817,N_2722,N_2730);
and U2818 (N_2818,N_2712,N_2736);
nand U2819 (N_2819,N_2711,N_2750);
and U2820 (N_2820,N_2810,N_2772);
nand U2821 (N_2821,N_2816,N_2796);
nor U2822 (N_2822,N_2793,N_2764);
nand U2823 (N_2823,N_2779,N_2763);
nand U2824 (N_2824,N_2802,N_2807);
nand U2825 (N_2825,N_2787,N_2790);
nand U2826 (N_2826,N_2804,N_2760);
nor U2827 (N_2827,N_2765,N_2791);
or U2828 (N_2828,N_2792,N_2770);
nor U2829 (N_2829,N_2812,N_2761);
nor U2830 (N_2830,N_2771,N_2769);
nand U2831 (N_2831,N_2811,N_2784);
nand U2832 (N_2832,N_2794,N_2776);
nor U2833 (N_2833,N_2798,N_2777);
or U2834 (N_2834,N_2782,N_2800);
nor U2835 (N_2835,N_2799,N_2775);
and U2836 (N_2836,N_2785,N_2795);
nand U2837 (N_2837,N_2783,N_2767);
or U2838 (N_2838,N_2801,N_2808);
xnor U2839 (N_2839,N_2766,N_2806);
or U2840 (N_2840,N_2819,N_2788);
or U2841 (N_2841,N_2809,N_2778);
or U2842 (N_2842,N_2813,N_2803);
and U2843 (N_2843,N_2805,N_2768);
nand U2844 (N_2844,N_2774,N_2780);
and U2845 (N_2845,N_2797,N_2773);
or U2846 (N_2846,N_2762,N_2781);
nand U2847 (N_2847,N_2818,N_2817);
or U2848 (N_2848,N_2786,N_2789);
and U2849 (N_2849,N_2815,N_2814);
nor U2850 (N_2850,N_2785,N_2793);
and U2851 (N_2851,N_2805,N_2815);
and U2852 (N_2852,N_2803,N_2779);
or U2853 (N_2853,N_2796,N_2772);
and U2854 (N_2854,N_2782,N_2783);
nand U2855 (N_2855,N_2767,N_2772);
nand U2856 (N_2856,N_2800,N_2803);
nor U2857 (N_2857,N_2778,N_2769);
nor U2858 (N_2858,N_2773,N_2793);
or U2859 (N_2859,N_2781,N_2776);
nor U2860 (N_2860,N_2761,N_2787);
or U2861 (N_2861,N_2816,N_2790);
nand U2862 (N_2862,N_2793,N_2809);
nor U2863 (N_2863,N_2793,N_2816);
nand U2864 (N_2864,N_2791,N_2784);
nand U2865 (N_2865,N_2800,N_2780);
and U2866 (N_2866,N_2806,N_2785);
and U2867 (N_2867,N_2779,N_2777);
and U2868 (N_2868,N_2796,N_2784);
nor U2869 (N_2869,N_2811,N_2797);
nor U2870 (N_2870,N_2813,N_2771);
and U2871 (N_2871,N_2772,N_2808);
or U2872 (N_2872,N_2775,N_2780);
nor U2873 (N_2873,N_2811,N_2782);
or U2874 (N_2874,N_2779,N_2762);
or U2875 (N_2875,N_2800,N_2802);
nand U2876 (N_2876,N_2809,N_2796);
nor U2877 (N_2877,N_2789,N_2768);
xor U2878 (N_2878,N_2790,N_2783);
or U2879 (N_2879,N_2805,N_2806);
or U2880 (N_2880,N_2821,N_2878);
nand U2881 (N_2881,N_2873,N_2870);
nor U2882 (N_2882,N_2866,N_2828);
and U2883 (N_2883,N_2829,N_2825);
and U2884 (N_2884,N_2846,N_2862);
nor U2885 (N_2885,N_2842,N_2848);
nor U2886 (N_2886,N_2852,N_2849);
or U2887 (N_2887,N_2853,N_2850);
nand U2888 (N_2888,N_2869,N_2864);
nand U2889 (N_2889,N_2841,N_2820);
and U2890 (N_2890,N_2868,N_2824);
or U2891 (N_2891,N_2856,N_2833);
and U2892 (N_2892,N_2877,N_2836);
and U2893 (N_2893,N_2871,N_2826);
or U2894 (N_2894,N_2844,N_2879);
nor U2895 (N_2895,N_2865,N_2835);
or U2896 (N_2896,N_2860,N_2867);
nand U2897 (N_2897,N_2861,N_2858);
nor U2898 (N_2898,N_2874,N_2831);
nand U2899 (N_2899,N_2827,N_2822);
and U2900 (N_2900,N_2851,N_2839);
and U2901 (N_2901,N_2832,N_2830);
nor U2902 (N_2902,N_2876,N_2847);
or U2903 (N_2903,N_2823,N_2872);
nand U2904 (N_2904,N_2834,N_2837);
nor U2905 (N_2905,N_2855,N_2838);
nand U2906 (N_2906,N_2857,N_2859);
and U2907 (N_2907,N_2863,N_2854);
or U2908 (N_2908,N_2843,N_2840);
nand U2909 (N_2909,N_2845,N_2875);
or U2910 (N_2910,N_2873,N_2841);
or U2911 (N_2911,N_2841,N_2864);
nand U2912 (N_2912,N_2879,N_2833);
nand U2913 (N_2913,N_2825,N_2827);
and U2914 (N_2914,N_2863,N_2851);
nand U2915 (N_2915,N_2849,N_2851);
nor U2916 (N_2916,N_2826,N_2868);
and U2917 (N_2917,N_2840,N_2855);
and U2918 (N_2918,N_2825,N_2877);
or U2919 (N_2919,N_2847,N_2845);
nor U2920 (N_2920,N_2848,N_2857);
and U2921 (N_2921,N_2828,N_2869);
and U2922 (N_2922,N_2877,N_2835);
nand U2923 (N_2923,N_2866,N_2841);
nor U2924 (N_2924,N_2844,N_2872);
nand U2925 (N_2925,N_2838,N_2823);
nand U2926 (N_2926,N_2820,N_2857);
nor U2927 (N_2927,N_2846,N_2857);
xnor U2928 (N_2928,N_2874,N_2846);
or U2929 (N_2929,N_2835,N_2845);
and U2930 (N_2930,N_2853,N_2824);
and U2931 (N_2931,N_2820,N_2872);
or U2932 (N_2932,N_2872,N_2861);
nor U2933 (N_2933,N_2838,N_2875);
and U2934 (N_2934,N_2844,N_2863);
nand U2935 (N_2935,N_2839,N_2842);
or U2936 (N_2936,N_2874,N_2866);
and U2937 (N_2937,N_2860,N_2879);
nand U2938 (N_2938,N_2856,N_2820);
nor U2939 (N_2939,N_2832,N_2849);
or U2940 (N_2940,N_2930,N_2928);
nand U2941 (N_2941,N_2901,N_2907);
or U2942 (N_2942,N_2886,N_2931);
and U2943 (N_2943,N_2917,N_2897);
nand U2944 (N_2944,N_2923,N_2922);
or U2945 (N_2945,N_2888,N_2937);
nor U2946 (N_2946,N_2889,N_2898);
nand U2947 (N_2947,N_2899,N_2925);
nand U2948 (N_2948,N_2903,N_2934);
and U2949 (N_2949,N_2906,N_2935);
or U2950 (N_2950,N_2924,N_2919);
and U2951 (N_2951,N_2914,N_2936);
nor U2952 (N_2952,N_2882,N_2920);
and U2953 (N_2953,N_2894,N_2926);
nand U2954 (N_2954,N_2938,N_2893);
or U2955 (N_2955,N_2916,N_2891);
nand U2956 (N_2956,N_2887,N_2910);
and U2957 (N_2957,N_2933,N_2881);
or U2958 (N_2958,N_2915,N_2927);
xnor U2959 (N_2959,N_2884,N_2918);
nand U2960 (N_2960,N_2932,N_2890);
and U2961 (N_2961,N_2905,N_2912);
nor U2962 (N_2962,N_2921,N_2929);
nor U2963 (N_2963,N_2908,N_2909);
nor U2964 (N_2964,N_2896,N_2892);
or U2965 (N_2965,N_2913,N_2885);
xnor U2966 (N_2966,N_2900,N_2911);
nor U2967 (N_2967,N_2904,N_2939);
or U2968 (N_2968,N_2902,N_2880);
and U2969 (N_2969,N_2895,N_2883);
and U2970 (N_2970,N_2938,N_2884);
nand U2971 (N_2971,N_2920,N_2909);
nor U2972 (N_2972,N_2903,N_2893);
nand U2973 (N_2973,N_2898,N_2890);
or U2974 (N_2974,N_2890,N_2928);
or U2975 (N_2975,N_2928,N_2916);
and U2976 (N_2976,N_2919,N_2908);
and U2977 (N_2977,N_2918,N_2888);
and U2978 (N_2978,N_2888,N_2933);
and U2979 (N_2979,N_2899,N_2912);
and U2980 (N_2980,N_2898,N_2901);
nor U2981 (N_2981,N_2880,N_2906);
or U2982 (N_2982,N_2920,N_2927);
nand U2983 (N_2983,N_2888,N_2917);
or U2984 (N_2984,N_2906,N_2902);
nand U2985 (N_2985,N_2880,N_2905);
or U2986 (N_2986,N_2883,N_2896);
nand U2987 (N_2987,N_2881,N_2920);
and U2988 (N_2988,N_2894,N_2920);
or U2989 (N_2989,N_2937,N_2881);
and U2990 (N_2990,N_2886,N_2937);
nor U2991 (N_2991,N_2891,N_2896);
or U2992 (N_2992,N_2922,N_2895);
nor U2993 (N_2993,N_2897,N_2881);
and U2994 (N_2994,N_2883,N_2925);
or U2995 (N_2995,N_2895,N_2889);
or U2996 (N_2996,N_2937,N_2917);
nand U2997 (N_2997,N_2881,N_2891);
nor U2998 (N_2998,N_2932,N_2904);
nor U2999 (N_2999,N_2896,N_2909);
nand UO_0 (O_0,N_2963,N_2942);
nand UO_1 (O_1,N_2982,N_2960);
and UO_2 (O_2,N_2983,N_2997);
nor UO_3 (O_3,N_2946,N_2940);
nor UO_4 (O_4,N_2992,N_2993);
and UO_5 (O_5,N_2944,N_2947);
nand UO_6 (O_6,N_2943,N_2956);
nand UO_7 (O_7,N_2959,N_2953);
xnor UO_8 (O_8,N_2998,N_2978);
nand UO_9 (O_9,N_2954,N_2969);
and UO_10 (O_10,N_2984,N_2968);
and UO_11 (O_11,N_2981,N_2964);
nor UO_12 (O_12,N_2941,N_2975);
or UO_13 (O_13,N_2961,N_2996);
xnor UO_14 (O_14,N_2977,N_2962);
nand UO_15 (O_15,N_2971,N_2986);
nand UO_16 (O_16,N_2987,N_2999);
nor UO_17 (O_17,N_2988,N_2958);
nor UO_18 (O_18,N_2967,N_2966);
or UO_19 (O_19,N_2991,N_2974);
nor UO_20 (O_20,N_2949,N_2972);
nor UO_21 (O_21,N_2990,N_2994);
nand UO_22 (O_22,N_2980,N_2995);
and UO_23 (O_23,N_2955,N_2957);
or UO_24 (O_24,N_2965,N_2985);
or UO_25 (O_25,N_2948,N_2989);
xnor UO_26 (O_26,N_2951,N_2976);
nor UO_27 (O_27,N_2979,N_2950);
or UO_28 (O_28,N_2952,N_2945);
and UO_29 (O_29,N_2973,N_2970);
nand UO_30 (O_30,N_2999,N_2975);
nand UO_31 (O_31,N_2970,N_2977);
and UO_32 (O_32,N_2952,N_2940);
nor UO_33 (O_33,N_2995,N_2958);
or UO_34 (O_34,N_2966,N_2973);
or UO_35 (O_35,N_2973,N_2978);
nor UO_36 (O_36,N_2996,N_2946);
or UO_37 (O_37,N_2956,N_2960);
nor UO_38 (O_38,N_2976,N_2949);
xor UO_39 (O_39,N_2942,N_2991);
nand UO_40 (O_40,N_2974,N_2949);
nor UO_41 (O_41,N_2947,N_2974);
or UO_42 (O_42,N_2987,N_2991);
and UO_43 (O_43,N_2950,N_2980);
and UO_44 (O_44,N_2993,N_2962);
nand UO_45 (O_45,N_2971,N_2956);
nor UO_46 (O_46,N_2953,N_2973);
and UO_47 (O_47,N_2998,N_2991);
and UO_48 (O_48,N_2979,N_2984);
nor UO_49 (O_49,N_2947,N_2960);
nor UO_50 (O_50,N_2959,N_2954);
and UO_51 (O_51,N_2991,N_2947);
and UO_52 (O_52,N_2947,N_2951);
nand UO_53 (O_53,N_2953,N_2944);
nor UO_54 (O_54,N_2983,N_2978);
or UO_55 (O_55,N_2973,N_2981);
nand UO_56 (O_56,N_2997,N_2993);
and UO_57 (O_57,N_2953,N_2992);
and UO_58 (O_58,N_2976,N_2992);
and UO_59 (O_59,N_2989,N_2998);
nand UO_60 (O_60,N_2952,N_2941);
nor UO_61 (O_61,N_2984,N_2961);
and UO_62 (O_62,N_2975,N_2973);
nor UO_63 (O_63,N_2985,N_2958);
and UO_64 (O_64,N_2960,N_2948);
nand UO_65 (O_65,N_2980,N_2983);
or UO_66 (O_66,N_2997,N_2990);
or UO_67 (O_67,N_2972,N_2942);
or UO_68 (O_68,N_2949,N_2946);
nor UO_69 (O_69,N_2976,N_2980);
nand UO_70 (O_70,N_2977,N_2999);
nand UO_71 (O_71,N_2948,N_2951);
nand UO_72 (O_72,N_2955,N_2986);
nor UO_73 (O_73,N_2956,N_2957);
and UO_74 (O_74,N_2982,N_2996);
and UO_75 (O_75,N_2955,N_2959);
nand UO_76 (O_76,N_2993,N_2998);
and UO_77 (O_77,N_2992,N_2998);
nand UO_78 (O_78,N_2954,N_2974);
nand UO_79 (O_79,N_2952,N_2996);
or UO_80 (O_80,N_2967,N_2985);
and UO_81 (O_81,N_2975,N_2951);
nor UO_82 (O_82,N_2943,N_2991);
nand UO_83 (O_83,N_2994,N_2953);
and UO_84 (O_84,N_2964,N_2971);
nor UO_85 (O_85,N_2967,N_2965);
or UO_86 (O_86,N_2949,N_2959);
nand UO_87 (O_87,N_2973,N_2948);
and UO_88 (O_88,N_2984,N_2974);
or UO_89 (O_89,N_2969,N_2987);
and UO_90 (O_90,N_2968,N_2967);
nand UO_91 (O_91,N_2963,N_2984);
xnor UO_92 (O_92,N_2941,N_2958);
or UO_93 (O_93,N_2995,N_2966);
or UO_94 (O_94,N_2982,N_2962);
and UO_95 (O_95,N_2980,N_2986);
or UO_96 (O_96,N_2956,N_2961);
nor UO_97 (O_97,N_2981,N_2971);
nor UO_98 (O_98,N_2974,N_2957);
nand UO_99 (O_99,N_2953,N_2999);
or UO_100 (O_100,N_2948,N_2976);
or UO_101 (O_101,N_2955,N_2940);
nor UO_102 (O_102,N_2966,N_2992);
nand UO_103 (O_103,N_2961,N_2982);
nand UO_104 (O_104,N_2958,N_2966);
and UO_105 (O_105,N_2999,N_2956);
or UO_106 (O_106,N_2978,N_2996);
nand UO_107 (O_107,N_2949,N_2997);
nor UO_108 (O_108,N_2942,N_2995);
or UO_109 (O_109,N_2956,N_2996);
or UO_110 (O_110,N_2993,N_2942);
or UO_111 (O_111,N_2955,N_2990);
nand UO_112 (O_112,N_2994,N_2989);
or UO_113 (O_113,N_2964,N_2966);
nor UO_114 (O_114,N_2997,N_2961);
and UO_115 (O_115,N_2992,N_2961);
and UO_116 (O_116,N_2955,N_2981);
or UO_117 (O_117,N_2967,N_2960);
xnor UO_118 (O_118,N_2966,N_2990);
and UO_119 (O_119,N_2958,N_2955);
or UO_120 (O_120,N_2962,N_2976);
or UO_121 (O_121,N_2941,N_2986);
nand UO_122 (O_122,N_2984,N_2980);
nand UO_123 (O_123,N_2958,N_2975);
and UO_124 (O_124,N_2990,N_2996);
or UO_125 (O_125,N_2949,N_2984);
nor UO_126 (O_126,N_2994,N_2968);
nor UO_127 (O_127,N_2979,N_2994);
nor UO_128 (O_128,N_2964,N_2985);
or UO_129 (O_129,N_2956,N_2972);
nor UO_130 (O_130,N_2993,N_2960);
or UO_131 (O_131,N_2974,N_2941);
nand UO_132 (O_132,N_2951,N_2985);
and UO_133 (O_133,N_2967,N_2970);
nand UO_134 (O_134,N_2963,N_2945);
and UO_135 (O_135,N_2984,N_2992);
nor UO_136 (O_136,N_2992,N_2962);
xnor UO_137 (O_137,N_2950,N_2984);
and UO_138 (O_138,N_2993,N_2971);
nand UO_139 (O_139,N_2996,N_2986);
nor UO_140 (O_140,N_2957,N_2971);
nor UO_141 (O_141,N_2982,N_2945);
and UO_142 (O_142,N_2967,N_2972);
or UO_143 (O_143,N_2957,N_2978);
or UO_144 (O_144,N_2949,N_2953);
or UO_145 (O_145,N_2995,N_2955);
and UO_146 (O_146,N_2985,N_2969);
and UO_147 (O_147,N_2981,N_2966);
or UO_148 (O_148,N_2989,N_2985);
nor UO_149 (O_149,N_2952,N_2983);
nand UO_150 (O_150,N_2974,N_2955);
nand UO_151 (O_151,N_2990,N_2984);
nand UO_152 (O_152,N_2949,N_2945);
nor UO_153 (O_153,N_2999,N_2996);
and UO_154 (O_154,N_2944,N_2945);
nor UO_155 (O_155,N_2959,N_2975);
nand UO_156 (O_156,N_2986,N_2958);
nor UO_157 (O_157,N_2960,N_2979);
nor UO_158 (O_158,N_2946,N_2950);
nand UO_159 (O_159,N_2959,N_2983);
nor UO_160 (O_160,N_2957,N_2985);
or UO_161 (O_161,N_2999,N_2989);
xnor UO_162 (O_162,N_2982,N_2943);
or UO_163 (O_163,N_2954,N_2999);
or UO_164 (O_164,N_2972,N_2947);
or UO_165 (O_165,N_2946,N_2973);
nand UO_166 (O_166,N_2965,N_2999);
nor UO_167 (O_167,N_2973,N_2965);
or UO_168 (O_168,N_2971,N_2946);
xnor UO_169 (O_169,N_2997,N_2941);
nor UO_170 (O_170,N_2977,N_2940);
nor UO_171 (O_171,N_2944,N_2971);
nand UO_172 (O_172,N_2966,N_2972);
nor UO_173 (O_173,N_2999,N_2971);
nor UO_174 (O_174,N_2956,N_2983);
nor UO_175 (O_175,N_2985,N_2986);
and UO_176 (O_176,N_2957,N_2989);
nand UO_177 (O_177,N_2992,N_2979);
or UO_178 (O_178,N_2993,N_2982);
and UO_179 (O_179,N_2973,N_2964);
and UO_180 (O_180,N_2977,N_2954);
or UO_181 (O_181,N_2970,N_2965);
nand UO_182 (O_182,N_2996,N_2980);
or UO_183 (O_183,N_2998,N_2951);
or UO_184 (O_184,N_2941,N_2960);
or UO_185 (O_185,N_2981,N_2976);
nand UO_186 (O_186,N_2967,N_2954);
nor UO_187 (O_187,N_2964,N_2979);
or UO_188 (O_188,N_2999,N_2969);
or UO_189 (O_189,N_2968,N_2942);
nand UO_190 (O_190,N_2948,N_2979);
or UO_191 (O_191,N_2988,N_2963);
nor UO_192 (O_192,N_2988,N_2948);
or UO_193 (O_193,N_2943,N_2955);
nand UO_194 (O_194,N_2998,N_2965);
or UO_195 (O_195,N_2985,N_2972);
and UO_196 (O_196,N_2957,N_2970);
and UO_197 (O_197,N_2982,N_2986);
nand UO_198 (O_198,N_2965,N_2990);
xor UO_199 (O_199,N_2994,N_2981);
nor UO_200 (O_200,N_2971,N_2968);
nand UO_201 (O_201,N_2940,N_2989);
nand UO_202 (O_202,N_2991,N_2950);
and UO_203 (O_203,N_2986,N_2943);
or UO_204 (O_204,N_2973,N_2990);
nand UO_205 (O_205,N_2990,N_2951);
nor UO_206 (O_206,N_2990,N_2970);
or UO_207 (O_207,N_2950,N_2997);
or UO_208 (O_208,N_2983,N_2999);
nand UO_209 (O_209,N_2946,N_2964);
nand UO_210 (O_210,N_2987,N_2941);
nor UO_211 (O_211,N_2953,N_2997);
nand UO_212 (O_212,N_2981,N_2977);
nor UO_213 (O_213,N_2959,N_2961);
and UO_214 (O_214,N_2947,N_2976);
or UO_215 (O_215,N_2979,N_2942);
nor UO_216 (O_216,N_2955,N_2991);
nor UO_217 (O_217,N_2969,N_2943);
or UO_218 (O_218,N_2963,N_2951);
nor UO_219 (O_219,N_2941,N_2948);
nor UO_220 (O_220,N_2951,N_2941);
and UO_221 (O_221,N_2976,N_2953);
or UO_222 (O_222,N_2945,N_2973);
or UO_223 (O_223,N_2990,N_2993);
nand UO_224 (O_224,N_2990,N_2988);
nor UO_225 (O_225,N_2966,N_2942);
nand UO_226 (O_226,N_2976,N_2960);
xnor UO_227 (O_227,N_2989,N_2975);
nor UO_228 (O_228,N_2956,N_2986);
or UO_229 (O_229,N_2961,N_2967);
or UO_230 (O_230,N_2945,N_2948);
and UO_231 (O_231,N_2987,N_2971);
or UO_232 (O_232,N_2980,N_2977);
or UO_233 (O_233,N_2974,N_2978);
or UO_234 (O_234,N_2952,N_2979);
nor UO_235 (O_235,N_2981,N_2982);
nor UO_236 (O_236,N_2964,N_2954);
or UO_237 (O_237,N_2971,N_2948);
nor UO_238 (O_238,N_2980,N_2941);
or UO_239 (O_239,N_2997,N_2985);
xnor UO_240 (O_240,N_2997,N_2957);
or UO_241 (O_241,N_2962,N_2960);
nand UO_242 (O_242,N_2997,N_2980);
nor UO_243 (O_243,N_2974,N_2979);
and UO_244 (O_244,N_2994,N_2976);
or UO_245 (O_245,N_2943,N_2948);
or UO_246 (O_246,N_2941,N_2992);
and UO_247 (O_247,N_2949,N_2998);
nand UO_248 (O_248,N_2963,N_2992);
nand UO_249 (O_249,N_2950,N_2981);
nand UO_250 (O_250,N_2994,N_2977);
and UO_251 (O_251,N_2959,N_2969);
nor UO_252 (O_252,N_2945,N_2965);
or UO_253 (O_253,N_2976,N_2943);
nor UO_254 (O_254,N_2943,N_2973);
xor UO_255 (O_255,N_2957,N_2962);
nand UO_256 (O_256,N_2980,N_2970);
or UO_257 (O_257,N_2986,N_2988);
nand UO_258 (O_258,N_2946,N_2954);
nor UO_259 (O_259,N_2957,N_2967);
nor UO_260 (O_260,N_2968,N_2953);
nand UO_261 (O_261,N_2972,N_2974);
nand UO_262 (O_262,N_2981,N_2956);
or UO_263 (O_263,N_2982,N_2955);
or UO_264 (O_264,N_2989,N_2949);
or UO_265 (O_265,N_2951,N_2981);
nor UO_266 (O_266,N_2964,N_2996);
nor UO_267 (O_267,N_2957,N_2964);
and UO_268 (O_268,N_2940,N_2981);
nor UO_269 (O_269,N_2948,N_2982);
and UO_270 (O_270,N_2963,N_2959);
and UO_271 (O_271,N_2975,N_2965);
nor UO_272 (O_272,N_2960,N_2959);
and UO_273 (O_273,N_2977,N_2988);
and UO_274 (O_274,N_2941,N_2981);
nor UO_275 (O_275,N_2977,N_2949);
and UO_276 (O_276,N_2972,N_2970);
nor UO_277 (O_277,N_2952,N_2997);
nand UO_278 (O_278,N_2984,N_2966);
and UO_279 (O_279,N_2981,N_2960);
and UO_280 (O_280,N_2988,N_2985);
and UO_281 (O_281,N_2955,N_2997);
or UO_282 (O_282,N_2983,N_2990);
xnor UO_283 (O_283,N_2998,N_2999);
nand UO_284 (O_284,N_2960,N_2953);
nand UO_285 (O_285,N_2969,N_2961);
or UO_286 (O_286,N_2977,N_2943);
and UO_287 (O_287,N_2989,N_2956);
nor UO_288 (O_288,N_2966,N_2983);
nand UO_289 (O_289,N_2961,N_2991);
nor UO_290 (O_290,N_2969,N_2990);
nor UO_291 (O_291,N_2989,N_2962);
and UO_292 (O_292,N_2974,N_2965);
and UO_293 (O_293,N_2980,N_2969);
nand UO_294 (O_294,N_2955,N_2998);
nor UO_295 (O_295,N_2973,N_2942);
nand UO_296 (O_296,N_2972,N_2965);
nand UO_297 (O_297,N_2984,N_2972);
or UO_298 (O_298,N_2988,N_2991);
or UO_299 (O_299,N_2947,N_2965);
or UO_300 (O_300,N_2999,N_2985);
nor UO_301 (O_301,N_2975,N_2964);
and UO_302 (O_302,N_2980,N_2992);
and UO_303 (O_303,N_2961,N_2952);
or UO_304 (O_304,N_2982,N_2968);
or UO_305 (O_305,N_2946,N_2960);
nor UO_306 (O_306,N_2961,N_2949);
and UO_307 (O_307,N_2995,N_2986);
and UO_308 (O_308,N_2953,N_2981);
nand UO_309 (O_309,N_2989,N_2986);
nand UO_310 (O_310,N_2949,N_2952);
xor UO_311 (O_311,N_2996,N_2968);
nand UO_312 (O_312,N_2942,N_2990);
nand UO_313 (O_313,N_2958,N_2980);
xor UO_314 (O_314,N_2984,N_2948);
nor UO_315 (O_315,N_2973,N_2986);
nor UO_316 (O_316,N_2966,N_2988);
nor UO_317 (O_317,N_2946,N_2988);
and UO_318 (O_318,N_2989,N_2973);
nand UO_319 (O_319,N_2958,N_2962);
or UO_320 (O_320,N_2942,N_2996);
and UO_321 (O_321,N_2948,N_2996);
nand UO_322 (O_322,N_2970,N_2993);
and UO_323 (O_323,N_2997,N_2954);
nor UO_324 (O_324,N_2975,N_2986);
xnor UO_325 (O_325,N_2955,N_2950);
or UO_326 (O_326,N_2998,N_2994);
and UO_327 (O_327,N_2985,N_2982);
nor UO_328 (O_328,N_2998,N_2945);
nor UO_329 (O_329,N_2957,N_2940);
and UO_330 (O_330,N_2960,N_2991);
and UO_331 (O_331,N_2985,N_2946);
and UO_332 (O_332,N_2984,N_2996);
nor UO_333 (O_333,N_2971,N_2980);
and UO_334 (O_334,N_2982,N_2952);
nor UO_335 (O_335,N_2952,N_2967);
nor UO_336 (O_336,N_2966,N_2943);
nand UO_337 (O_337,N_2966,N_2998);
nor UO_338 (O_338,N_2940,N_2944);
nor UO_339 (O_339,N_2961,N_2946);
and UO_340 (O_340,N_2948,N_2983);
nor UO_341 (O_341,N_2973,N_2963);
or UO_342 (O_342,N_2944,N_2992);
nor UO_343 (O_343,N_2942,N_2982);
or UO_344 (O_344,N_2972,N_2961);
nand UO_345 (O_345,N_2950,N_2964);
or UO_346 (O_346,N_2971,N_2974);
nand UO_347 (O_347,N_2990,N_2944);
or UO_348 (O_348,N_2945,N_2942);
nor UO_349 (O_349,N_2949,N_2985);
nand UO_350 (O_350,N_2950,N_2987);
nand UO_351 (O_351,N_2996,N_2995);
or UO_352 (O_352,N_2953,N_2941);
nand UO_353 (O_353,N_2999,N_2968);
nand UO_354 (O_354,N_2980,N_2966);
nand UO_355 (O_355,N_2959,N_2988);
and UO_356 (O_356,N_2992,N_2986);
nor UO_357 (O_357,N_2998,N_2985);
or UO_358 (O_358,N_2999,N_2941);
nor UO_359 (O_359,N_2995,N_2978);
or UO_360 (O_360,N_2946,N_2958);
nand UO_361 (O_361,N_2956,N_2975);
or UO_362 (O_362,N_2970,N_2996);
nor UO_363 (O_363,N_2942,N_2952);
nor UO_364 (O_364,N_2956,N_2976);
nand UO_365 (O_365,N_2985,N_2973);
nand UO_366 (O_366,N_2993,N_2940);
nand UO_367 (O_367,N_2948,N_2963);
nor UO_368 (O_368,N_2985,N_2978);
or UO_369 (O_369,N_2973,N_2974);
and UO_370 (O_370,N_2983,N_2987);
nand UO_371 (O_371,N_2970,N_2988);
nor UO_372 (O_372,N_2970,N_2945);
nand UO_373 (O_373,N_2975,N_2977);
nand UO_374 (O_374,N_2940,N_2951);
or UO_375 (O_375,N_2973,N_2952);
nand UO_376 (O_376,N_2992,N_2990);
nand UO_377 (O_377,N_2959,N_2940);
nand UO_378 (O_378,N_2960,N_2972);
or UO_379 (O_379,N_2968,N_2966);
and UO_380 (O_380,N_2958,N_2952);
or UO_381 (O_381,N_2979,N_2986);
nor UO_382 (O_382,N_2948,N_2998);
and UO_383 (O_383,N_2948,N_2956);
and UO_384 (O_384,N_2962,N_2973);
and UO_385 (O_385,N_2983,N_2965);
and UO_386 (O_386,N_2969,N_2975);
nand UO_387 (O_387,N_2975,N_2982);
and UO_388 (O_388,N_2959,N_2980);
nand UO_389 (O_389,N_2962,N_2979);
nand UO_390 (O_390,N_2959,N_2981);
nand UO_391 (O_391,N_2989,N_2968);
and UO_392 (O_392,N_2962,N_2963);
or UO_393 (O_393,N_2952,N_2980);
nor UO_394 (O_394,N_2972,N_2968);
and UO_395 (O_395,N_2972,N_2946);
or UO_396 (O_396,N_2997,N_2992);
nand UO_397 (O_397,N_2962,N_2996);
nor UO_398 (O_398,N_2993,N_2958);
nor UO_399 (O_399,N_2943,N_2974);
and UO_400 (O_400,N_2965,N_2994);
nor UO_401 (O_401,N_2986,N_2966);
or UO_402 (O_402,N_2991,N_2993);
nand UO_403 (O_403,N_2943,N_2988);
and UO_404 (O_404,N_2954,N_2980);
and UO_405 (O_405,N_2970,N_2952);
and UO_406 (O_406,N_2950,N_2953);
or UO_407 (O_407,N_2967,N_2984);
nand UO_408 (O_408,N_2955,N_2963);
nor UO_409 (O_409,N_2995,N_2976);
nor UO_410 (O_410,N_2995,N_2999);
nand UO_411 (O_411,N_2953,N_2972);
nor UO_412 (O_412,N_2940,N_2949);
nor UO_413 (O_413,N_2960,N_2952);
nor UO_414 (O_414,N_2973,N_2954);
or UO_415 (O_415,N_2974,N_2945);
nor UO_416 (O_416,N_2994,N_2958);
and UO_417 (O_417,N_2979,N_2958);
or UO_418 (O_418,N_2978,N_2965);
nand UO_419 (O_419,N_2945,N_2999);
nand UO_420 (O_420,N_2979,N_2965);
nand UO_421 (O_421,N_2987,N_2953);
nand UO_422 (O_422,N_2977,N_2979);
nor UO_423 (O_423,N_2995,N_2969);
nand UO_424 (O_424,N_2982,N_2963);
and UO_425 (O_425,N_2987,N_2996);
nor UO_426 (O_426,N_2945,N_2977);
or UO_427 (O_427,N_2994,N_2962);
or UO_428 (O_428,N_2983,N_2986);
and UO_429 (O_429,N_2993,N_2966);
and UO_430 (O_430,N_2985,N_2954);
or UO_431 (O_431,N_2981,N_2991);
nand UO_432 (O_432,N_2947,N_2959);
and UO_433 (O_433,N_2977,N_2953);
nand UO_434 (O_434,N_2968,N_2949);
and UO_435 (O_435,N_2960,N_2975);
and UO_436 (O_436,N_2950,N_2956);
or UO_437 (O_437,N_2953,N_2990);
nand UO_438 (O_438,N_2948,N_2978);
nor UO_439 (O_439,N_2997,N_2979);
xor UO_440 (O_440,N_2942,N_2959);
nor UO_441 (O_441,N_2986,N_2998);
and UO_442 (O_442,N_2957,N_2992);
or UO_443 (O_443,N_2976,N_2946);
or UO_444 (O_444,N_2958,N_2987);
and UO_445 (O_445,N_2983,N_2950);
or UO_446 (O_446,N_2941,N_2973);
nand UO_447 (O_447,N_2944,N_2974);
or UO_448 (O_448,N_2946,N_2947);
nand UO_449 (O_449,N_2967,N_2982);
nor UO_450 (O_450,N_2972,N_2988);
or UO_451 (O_451,N_2951,N_2983);
nor UO_452 (O_452,N_2967,N_2987);
nor UO_453 (O_453,N_2994,N_2948);
and UO_454 (O_454,N_2999,N_2981);
nor UO_455 (O_455,N_2987,N_2940);
nand UO_456 (O_456,N_2955,N_2969);
nand UO_457 (O_457,N_2971,N_2991);
nor UO_458 (O_458,N_2977,N_2957);
or UO_459 (O_459,N_2952,N_2950);
or UO_460 (O_460,N_2964,N_2994);
nor UO_461 (O_461,N_2948,N_2966);
or UO_462 (O_462,N_2963,N_2969);
and UO_463 (O_463,N_2993,N_2972);
and UO_464 (O_464,N_2965,N_2988);
or UO_465 (O_465,N_2981,N_2978);
or UO_466 (O_466,N_2959,N_2944);
nor UO_467 (O_467,N_2995,N_2965);
xnor UO_468 (O_468,N_2956,N_2970);
or UO_469 (O_469,N_2946,N_2986);
or UO_470 (O_470,N_2986,N_2977);
nor UO_471 (O_471,N_2960,N_2966);
and UO_472 (O_472,N_2945,N_2940);
or UO_473 (O_473,N_2997,N_2951);
and UO_474 (O_474,N_2992,N_2971);
nor UO_475 (O_475,N_2971,N_2952);
xnor UO_476 (O_476,N_2994,N_2946);
or UO_477 (O_477,N_2941,N_2949);
and UO_478 (O_478,N_2955,N_2941);
or UO_479 (O_479,N_2993,N_2957);
nor UO_480 (O_480,N_2987,N_2974);
or UO_481 (O_481,N_2946,N_2969);
and UO_482 (O_482,N_2984,N_2955);
and UO_483 (O_483,N_2992,N_2956);
nor UO_484 (O_484,N_2964,N_2944);
xor UO_485 (O_485,N_2988,N_2987);
nand UO_486 (O_486,N_2982,N_2995);
and UO_487 (O_487,N_2947,N_2986);
and UO_488 (O_488,N_2940,N_2956);
nand UO_489 (O_489,N_2985,N_2942);
or UO_490 (O_490,N_2949,N_2948);
nor UO_491 (O_491,N_2947,N_2955);
nor UO_492 (O_492,N_2985,N_2980);
nor UO_493 (O_493,N_2952,N_2956);
nor UO_494 (O_494,N_2967,N_2991);
nand UO_495 (O_495,N_2950,N_2940);
xnor UO_496 (O_496,N_2960,N_2942);
nor UO_497 (O_497,N_2954,N_2990);
or UO_498 (O_498,N_2953,N_2967);
nor UO_499 (O_499,N_2988,N_2951);
endmodule