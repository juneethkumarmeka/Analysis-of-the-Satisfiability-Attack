module basic_1500_15000_2000_75_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_458,In_991);
nor U1 (N_1,In_1495,In_423);
and U2 (N_2,In_692,In_1085);
xnor U3 (N_3,In_1365,In_941);
xnor U4 (N_4,In_6,In_608);
and U5 (N_5,In_647,In_1160);
xor U6 (N_6,In_709,In_751);
xor U7 (N_7,In_1334,In_1093);
and U8 (N_8,In_1161,In_1314);
or U9 (N_9,In_710,In_1186);
and U10 (N_10,In_65,In_939);
nor U11 (N_11,In_407,In_822);
nor U12 (N_12,In_1348,In_628);
nor U13 (N_13,In_209,In_1385);
or U14 (N_14,In_210,In_576);
and U15 (N_15,In_1122,In_1062);
xor U16 (N_16,In_800,In_323);
and U17 (N_17,In_777,In_203);
xor U18 (N_18,In_688,In_821);
nand U19 (N_19,In_656,In_24);
and U20 (N_20,In_781,In_1191);
or U21 (N_21,In_808,In_363);
and U22 (N_22,In_389,In_1281);
and U23 (N_23,In_181,In_326);
and U24 (N_24,In_55,In_318);
nand U25 (N_25,In_857,In_796);
or U26 (N_26,In_1342,In_330);
and U27 (N_27,In_737,In_1194);
and U28 (N_28,In_607,In_726);
nand U29 (N_29,In_75,In_695);
xor U30 (N_30,In_1114,In_1100);
nand U31 (N_31,In_1293,In_1286);
nor U32 (N_32,In_561,In_228);
nand U33 (N_33,In_1356,In_520);
and U34 (N_34,In_190,In_1136);
and U35 (N_35,In_759,In_1479);
nand U36 (N_36,In_570,In_1108);
xnor U37 (N_37,In_300,In_817);
xor U38 (N_38,In_527,In_1013);
and U39 (N_39,In_568,In_148);
nand U40 (N_40,In_590,In_1467);
or U41 (N_41,In_114,In_943);
or U42 (N_42,In_802,In_1390);
and U43 (N_43,In_866,In_658);
nor U44 (N_44,In_1192,In_31);
and U45 (N_45,In_1435,In_1273);
xnor U46 (N_46,In_672,In_522);
nor U47 (N_47,In_95,In_534);
and U48 (N_48,In_451,In_677);
and U49 (N_49,In_722,In_1204);
nand U50 (N_50,In_671,In_643);
or U51 (N_51,In_913,In_917);
or U52 (N_52,In_689,In_119);
nor U53 (N_53,In_305,In_401);
xor U54 (N_54,In_895,In_415);
nor U55 (N_55,In_724,In_1301);
and U56 (N_56,In_1229,In_627);
nor U57 (N_57,In_1035,In_188);
xnor U58 (N_58,In_135,In_34);
nand U59 (N_59,In_799,In_894);
or U60 (N_60,In_748,In_126);
or U61 (N_61,In_12,In_1140);
nand U62 (N_62,In_1487,In_680);
nor U63 (N_63,In_327,In_310);
xor U64 (N_64,In_20,In_771);
nand U65 (N_65,In_1378,In_1317);
xor U66 (N_66,In_954,In_521);
or U67 (N_67,In_984,In_195);
xor U68 (N_68,In_179,In_1185);
or U69 (N_69,In_388,In_1172);
or U70 (N_70,In_558,In_98);
xor U71 (N_71,In_809,In_452);
xor U72 (N_72,In_1022,In_366);
nor U73 (N_73,In_497,In_642);
and U74 (N_74,In_1488,In_812);
and U75 (N_75,In_1383,In_96);
nand U76 (N_76,In_1170,In_583);
and U77 (N_77,In_619,In_226);
nand U78 (N_78,In_43,In_836);
or U79 (N_79,In_436,In_1391);
xor U80 (N_80,In_1133,In_636);
and U81 (N_81,In_546,In_1368);
nor U82 (N_82,In_1375,In_1112);
and U83 (N_83,In_1327,In_1041);
and U84 (N_84,In_1296,In_1);
nor U85 (N_85,In_632,In_1490);
and U86 (N_86,In_1092,In_316);
or U87 (N_87,In_883,In_158);
xnor U88 (N_88,In_453,In_1277);
or U89 (N_89,In_1279,In_850);
xnor U90 (N_90,In_25,In_249);
xnor U91 (N_91,In_354,In_1451);
and U92 (N_92,In_871,In_942);
nand U93 (N_93,In_392,In_683);
xnor U94 (N_94,In_236,In_145);
and U95 (N_95,In_707,In_386);
nor U96 (N_96,In_912,In_693);
or U97 (N_97,In_1208,In_1266);
nor U98 (N_98,In_832,In_514);
nand U99 (N_99,In_506,In_1494);
and U100 (N_100,In_1312,In_1103);
nand U101 (N_101,In_294,In_1057);
nand U102 (N_102,In_845,In_640);
nand U103 (N_103,In_1267,In_1280);
nor U104 (N_104,In_633,In_1384);
nand U105 (N_105,In_1349,In_1351);
or U106 (N_106,In_1309,In_390);
nor U107 (N_107,In_69,In_512);
or U108 (N_108,In_1269,In_1037);
xor U109 (N_109,In_106,In_1329);
and U110 (N_110,In_189,In_509);
xnor U111 (N_111,In_807,In_923);
nand U112 (N_112,In_754,In_752);
nand U113 (N_113,In_56,In_1123);
or U114 (N_114,In_306,In_903);
and U115 (N_115,In_1463,In_296);
nor U116 (N_116,In_694,In_1496);
and U117 (N_117,In_581,In_345);
and U118 (N_118,In_1213,In_1178);
nand U119 (N_119,In_381,In_1295);
nand U120 (N_120,In_519,In_591);
nor U121 (N_121,In_595,In_1343);
nand U122 (N_122,In_770,In_52);
xnor U123 (N_123,In_1283,In_1104);
xor U124 (N_124,In_816,In_276);
nand U125 (N_125,In_379,In_610);
xnor U126 (N_126,In_1054,In_690);
nor U127 (N_127,In_1429,In_717);
and U128 (N_128,In_1012,In_612);
nor U129 (N_129,In_909,In_32);
nand U130 (N_130,In_140,In_8);
or U131 (N_131,In_653,In_284);
nand U132 (N_132,In_83,In_990);
xnor U133 (N_133,In_793,In_1302);
xnor U134 (N_134,In_960,In_47);
and U135 (N_135,In_412,In_670);
nor U136 (N_136,In_686,In_860);
xnor U137 (N_137,In_1124,In_938);
and U138 (N_138,In_1336,In_1203);
and U139 (N_139,In_668,In_964);
and U140 (N_140,In_71,In_1011);
xor U141 (N_141,In_347,In_955);
and U142 (N_142,In_1241,In_257);
nor U143 (N_143,In_852,In_1426);
nand U144 (N_144,In_993,In_729);
or U145 (N_145,In_1119,In_206);
nor U146 (N_146,In_250,In_1307);
xor U147 (N_147,In_1436,In_1238);
nor U148 (N_148,In_545,In_215);
xnor U149 (N_149,In_160,In_1313);
and U150 (N_150,In_108,In_157);
xnor U151 (N_151,In_1067,In_747);
or U152 (N_152,In_929,In_21);
nor U153 (N_153,In_1082,In_838);
or U154 (N_154,In_734,In_865);
nand U155 (N_155,In_1205,In_467);
and U156 (N_156,In_485,In_283);
nand U157 (N_157,In_1007,In_1315);
or U158 (N_158,In_1345,In_496);
xnor U159 (N_159,In_271,In_476);
xor U160 (N_160,In_1347,In_378);
and U161 (N_161,In_208,In_1405);
nand U162 (N_162,In_1472,In_718);
nand U163 (N_163,In_1017,In_1038);
nor U164 (N_164,In_996,In_1409);
xnor U165 (N_165,In_1246,In_1043);
and U166 (N_166,In_1476,In_471);
nor U167 (N_167,In_1094,In_785);
nor U168 (N_168,In_248,In_166);
or U169 (N_169,In_367,In_792);
nand U170 (N_170,In_932,In_535);
and U171 (N_171,In_1239,In_398);
nand U172 (N_172,In_1097,In_107);
nand U173 (N_173,In_635,In_40);
and U174 (N_174,In_1005,In_616);
xnor U175 (N_175,In_699,In_1392);
xnor U176 (N_176,In_580,In_1020);
nor U177 (N_177,In_1252,In_233);
and U178 (N_178,In_1287,In_118);
nand U179 (N_179,In_742,In_1319);
nand U180 (N_180,In_144,In_1394);
or U181 (N_181,In_7,In_1402);
xnor U182 (N_182,In_730,In_891);
xnor U183 (N_183,In_1053,In_925);
nand U184 (N_184,In_584,In_530);
nor U185 (N_185,In_30,In_665);
nor U186 (N_186,In_1395,In_1438);
or U187 (N_187,In_1481,In_893);
xor U188 (N_188,In_202,In_319);
or U189 (N_189,In_597,In_659);
or U190 (N_190,In_1200,In_46);
and U191 (N_191,In_1176,In_844);
nand U192 (N_192,In_1387,In_1175);
xnor U193 (N_193,In_151,In_432);
and U194 (N_194,In_370,In_1432);
nand U195 (N_195,In_1400,In_593);
nor U196 (N_196,In_1486,In_1498);
and U197 (N_197,In_1270,In_442);
xnor U198 (N_198,In_657,In_1066);
or U199 (N_199,In_337,In_981);
and U200 (N_200,N_95,In_1259);
nand U201 (N_201,In_59,N_134);
nor U202 (N_202,In_353,In_525);
nor U203 (N_203,In_1377,In_185);
nor U204 (N_204,In_1388,In_352);
and U205 (N_205,In_1121,In_1234);
nor U206 (N_206,In_192,N_196);
and U207 (N_207,In_557,In_1000);
nand U208 (N_208,In_502,In_1138);
or U209 (N_209,In_849,In_798);
and U210 (N_210,In_368,In_239);
xnor U211 (N_211,In_1499,In_1389);
xnor U212 (N_212,In_1397,In_908);
xor U213 (N_213,N_148,In_933);
nand U214 (N_214,N_8,In_28);
xnor U215 (N_215,N_75,In_1332);
nand U216 (N_216,N_55,In_505);
and U217 (N_217,In_872,N_86);
nand U218 (N_218,In_252,In_297);
and U219 (N_219,N_79,In_242);
or U220 (N_220,In_246,In_155);
nand U221 (N_221,In_961,In_380);
xor U222 (N_222,In_399,In_552);
nor U223 (N_223,In_1224,In_988);
nand U224 (N_224,In_1217,N_87);
and U225 (N_225,In_272,In_782);
and U226 (N_226,In_163,In_1257);
xor U227 (N_227,In_997,N_174);
or U228 (N_228,In_769,N_93);
and U229 (N_229,In_928,In_90);
nand U230 (N_230,N_115,In_18);
nor U231 (N_231,In_786,In_92);
nor U232 (N_232,In_1333,In_788);
nor U233 (N_233,In_1227,In_574);
nor U234 (N_234,In_1144,In_1320);
or U235 (N_235,In_1181,In_851);
nor U236 (N_236,In_1316,In_614);
and U237 (N_237,In_1148,In_281);
nand U238 (N_238,N_41,In_1360);
or U239 (N_239,In_182,In_419);
nand U240 (N_240,In_13,In_554);
or U241 (N_241,N_82,In_870);
nand U242 (N_242,In_1272,In_978);
xnor U243 (N_243,In_958,In_606);
nand U244 (N_244,In_231,In_1029);
or U245 (N_245,In_501,In_1271);
xnor U246 (N_246,In_644,In_1129);
nor U247 (N_247,In_445,In_803);
nor U248 (N_248,In_1090,In_667);
xor U249 (N_249,In_384,In_727);
nand U250 (N_250,In_806,N_162);
and U251 (N_251,In_930,N_72);
and U252 (N_252,In_868,In_555);
nand U253 (N_253,In_1457,In_475);
nor U254 (N_254,In_701,In_256);
and U255 (N_255,In_719,In_1081);
nand U256 (N_256,In_1045,In_1163);
nor U257 (N_257,N_27,In_1485);
nand U258 (N_258,In_507,In_712);
xnor U259 (N_259,In_1446,N_137);
and U260 (N_260,In_200,In_842);
or U261 (N_261,In_750,In_1105);
or U262 (N_262,In_481,N_121);
and U263 (N_263,In_130,N_163);
nand U264 (N_264,In_311,In_1423);
nand U265 (N_265,In_240,In_1084);
xnor U266 (N_266,In_1251,N_46);
and U267 (N_267,In_649,In_101);
and U268 (N_268,In_198,In_1417);
nand U269 (N_269,In_674,N_140);
nor U270 (N_270,In_819,In_1031);
nor U271 (N_271,In_324,In_1344);
nor U272 (N_272,In_23,In_1125);
nand U273 (N_273,In_890,In_758);
xnor U274 (N_274,In_251,In_1352);
nor U275 (N_275,N_71,In_936);
and U276 (N_276,In_333,In_457);
nor U277 (N_277,N_111,In_794);
nand U278 (N_278,In_431,In_149);
nand U279 (N_279,In_111,In_315);
and U280 (N_280,N_183,In_863);
nand U281 (N_281,In_1089,In_605);
nand U282 (N_282,In_914,In_499);
and U283 (N_283,In_818,In_312);
nor U284 (N_284,In_387,In_48);
nor U285 (N_285,In_599,In_847);
nand U286 (N_286,In_877,In_159);
and U287 (N_287,In_1132,N_130);
nand U288 (N_288,In_654,In_325);
or U289 (N_289,N_139,In_843);
xnor U290 (N_290,In_1294,In_575);
nor U291 (N_291,In_985,In_334);
xnor U292 (N_292,In_829,In_639);
xor U293 (N_293,In_1357,In_1036);
nand U294 (N_294,In_438,N_67);
nor U295 (N_295,In_298,In_110);
nor U296 (N_296,In_317,In_549);
nand U297 (N_297,In_238,In_1465);
nand U298 (N_298,In_214,In_886);
or U299 (N_299,N_173,In_704);
nand U300 (N_300,In_572,N_29);
and U301 (N_301,In_362,In_1300);
nand U302 (N_302,In_394,In_1049);
and U303 (N_303,In_1323,In_579);
xnor U304 (N_304,In_949,In_684);
and U305 (N_305,In_815,In_728);
and U306 (N_306,In_1080,In_732);
nand U307 (N_307,In_524,In_447);
nor U308 (N_308,In_217,In_1071);
and U309 (N_309,In_375,N_26);
nand U310 (N_310,In_146,In_259);
nand U311 (N_311,In_1372,In_772);
and U312 (N_312,N_84,In_1202);
nor U313 (N_313,In_503,In_889);
nand U314 (N_314,N_61,In_1308);
and U315 (N_315,In_918,N_195);
or U316 (N_316,In_1461,In_22);
xnor U317 (N_317,In_982,In_428);
xnor U318 (N_318,In_68,In_1127);
and U319 (N_319,In_1154,In_1077);
xnor U320 (N_320,In_1034,In_765);
xor U321 (N_321,In_651,In_1275);
or U322 (N_322,In_582,In_1219);
or U323 (N_323,In_1420,In_846);
nor U324 (N_324,N_132,N_192);
nand U325 (N_325,In_1015,In_420);
xnor U326 (N_326,In_377,In_129);
nor U327 (N_327,In_1276,In_966);
xnor U328 (N_328,N_151,In_813);
nor U329 (N_329,In_896,In_416);
nor U330 (N_330,In_1024,In_1424);
or U331 (N_331,In_980,In_735);
nand U332 (N_332,In_539,In_437);
nand U333 (N_333,In_935,In_1059);
xor U334 (N_334,In_213,In_897);
xor U335 (N_335,In_265,In_620);
nor U336 (N_336,In_725,In_738);
xor U337 (N_337,N_16,In_1450);
and U338 (N_338,In_1422,In_916);
nand U339 (N_339,In_624,In_790);
and U340 (N_340,In_266,In_1367);
xor U341 (N_341,In_666,N_22);
xor U342 (N_342,In_953,In_1381);
or U343 (N_343,In_791,In_1149);
or U344 (N_344,N_36,In_878);
nor U345 (N_345,In_355,In_253);
nand U346 (N_346,In_1455,In_1289);
xor U347 (N_347,In_461,In_876);
or U348 (N_348,In_926,In_1078);
nor U349 (N_349,In_127,In_542);
nand U350 (N_350,In_422,In_1413);
xnor U351 (N_351,In_102,N_4);
nand U352 (N_352,In_444,N_127);
xnor U353 (N_353,In_679,In_691);
and U354 (N_354,In_596,In_1142);
nor U355 (N_355,In_478,In_435);
nand U356 (N_356,In_1492,In_1070);
xnor U357 (N_357,In_1025,In_212);
or U358 (N_358,In_1366,In_99);
nand U359 (N_359,In_232,N_193);
xor U360 (N_360,N_96,In_267);
xor U361 (N_361,In_421,In_905);
nand U362 (N_362,In_856,In_439);
xnor U363 (N_363,N_145,In_1353);
nor U364 (N_364,In_810,In_466);
and U365 (N_365,N_40,In_559);
or U366 (N_366,In_1079,N_166);
or U367 (N_367,In_569,In_29);
xnor U368 (N_368,In_1173,In_901);
xnor U369 (N_369,N_182,In_950);
or U370 (N_370,In_180,In_1197);
nand U371 (N_371,In_811,In_641);
nand U372 (N_372,In_702,In_626);
and U373 (N_373,In_529,In_1134);
nand U374 (N_374,In_348,In_1087);
xor U375 (N_375,In_280,In_1177);
nor U376 (N_376,In_837,In_743);
nand U377 (N_377,In_540,In_0);
nor U378 (N_378,In_369,In_864);
xor U379 (N_379,In_1260,In_269);
or U380 (N_380,In_971,In_1354);
or U381 (N_381,In_646,In_38);
xnor U382 (N_382,In_1325,N_116);
nor U383 (N_383,In_840,In_125);
or U384 (N_384,N_33,In_650);
nand U385 (N_385,N_47,In_1456);
nand U386 (N_386,N_23,In_992);
and U387 (N_387,N_39,In_1139);
and U388 (N_388,In_621,In_1131);
or U389 (N_389,In_915,In_74);
nor U390 (N_390,In_678,N_106);
xnor U391 (N_391,In_587,In_516);
and U392 (N_392,In_1184,In_1477);
nand U393 (N_393,In_1410,In_1230);
and U394 (N_394,In_81,In_1051);
xnor U395 (N_395,In_264,In_35);
xor U396 (N_396,In_254,In_1180);
nor U397 (N_397,In_338,In_1050);
nor U398 (N_398,N_5,In_136);
nor U399 (N_399,N_6,In_94);
or U400 (N_400,N_164,In_495);
nor U401 (N_401,In_839,In_746);
or U402 (N_402,N_152,In_1117);
or U403 (N_403,In_655,N_398);
xor U404 (N_404,In_1158,In_1425);
nor U405 (N_405,N_279,In_426);
or U406 (N_406,N_49,N_161);
nor U407 (N_407,In_1466,In_304);
and U408 (N_408,In_773,In_273);
and U409 (N_409,N_56,In_1475);
nor U410 (N_410,In_413,In_731);
and U411 (N_411,N_198,In_875);
nand U412 (N_412,In_541,In_1374);
or U413 (N_413,N_147,N_153);
or U414 (N_414,In_417,N_209);
and U415 (N_415,In_1310,N_157);
xnor U416 (N_416,N_266,In_609);
nand U417 (N_417,N_158,In_1109);
or U418 (N_418,In_1399,In_430);
nor U419 (N_419,In_16,In_623);
xnor U420 (N_420,In_1428,In_613);
nand U421 (N_421,In_469,In_1253);
nand U422 (N_422,N_382,In_128);
xor U423 (N_423,N_108,N_262);
nor U424 (N_424,In_287,In_1222);
nand U425 (N_425,In_93,In_898);
or U426 (N_426,In_598,In_979);
nand U427 (N_427,N_114,In_1411);
xnor U428 (N_428,In_660,In_1376);
and U429 (N_429,N_112,N_83);
or U430 (N_430,N_270,N_248);
xor U431 (N_431,In_260,N_48);
and U432 (N_432,N_227,In_219);
or U433 (N_433,N_323,N_277);
or U434 (N_434,N_315,In_900);
and U435 (N_435,In_274,N_200);
and U436 (N_436,In_757,N_276);
or U437 (N_437,N_274,In_879);
nand U438 (N_438,In_974,In_1305);
nor U439 (N_439,In_617,In_1023);
or U440 (N_440,N_35,N_380);
nor U441 (N_441,N_230,In_1099);
or U442 (N_442,In_87,N_344);
or U443 (N_443,In_1221,In_1137);
and U444 (N_444,In_382,In_1198);
xor U445 (N_445,In_987,N_346);
nor U446 (N_446,N_288,In_1047);
and U447 (N_447,N_388,In_1183);
or U448 (N_448,In_313,In_427);
and U449 (N_449,In_594,N_189);
nor U450 (N_450,In_131,In_825);
xor U451 (N_451,In_622,In_1009);
xnor U452 (N_452,N_291,In_45);
xnor U453 (N_453,N_17,In_764);
and U454 (N_454,In_638,In_488);
nand U455 (N_455,In_329,In_328);
xnor U456 (N_456,In_784,In_681);
xor U457 (N_457,In_973,N_348);
nor U458 (N_458,In_1046,In_1240);
nor U459 (N_459,In_1497,In_880);
xor U460 (N_460,In_66,In_50);
xnor U461 (N_461,In_927,In_571);
xor U462 (N_462,N_303,In_295);
nor U463 (N_463,In_563,In_1225);
xor U464 (N_464,In_424,In_714);
nand U465 (N_465,In_1003,N_177);
or U466 (N_466,N_14,In_491);
or U467 (N_467,In_397,In_869);
or U468 (N_468,N_21,In_1261);
xnor U469 (N_469,In_207,In_1016);
xor U470 (N_470,In_1430,N_392);
xnor U471 (N_471,N_194,N_370);
nand U472 (N_472,N_15,N_30);
xor U473 (N_473,N_190,N_214);
and U474 (N_474,N_349,N_231);
xor U475 (N_475,In_162,In_711);
xor U476 (N_476,N_204,N_149);
or U477 (N_477,N_54,In_1040);
and U478 (N_478,N_13,N_18);
or U479 (N_479,In_1021,In_1006);
or U480 (N_480,In_1107,In_201);
and U481 (N_481,N_103,N_360);
or U482 (N_482,In_1361,In_1218);
nand U483 (N_483,In_1091,In_904);
or U484 (N_484,N_363,N_241);
xnor U485 (N_485,In_1118,In_945);
or U486 (N_486,In_855,N_311);
xnor U487 (N_487,In_286,N_356);
xnor U488 (N_488,N_142,In_592);
xnor U489 (N_489,In_1350,N_321);
and U490 (N_490,In_134,In_279);
and U491 (N_491,N_282,In_1339);
nand U492 (N_492,In_1268,N_373);
or U493 (N_493,In_986,In_1478);
or U494 (N_494,In_1026,N_38);
nor U495 (N_495,In_1207,In_1453);
nand U496 (N_496,N_271,N_237);
and U497 (N_497,In_972,In_346);
xnor U498 (N_498,N_299,In_448);
nand U499 (N_499,In_51,In_1076);
and U500 (N_500,In_1331,N_239);
and U501 (N_501,In_1433,In_396);
nand U502 (N_502,In_995,N_302);
xor U503 (N_503,In_761,In_72);
nor U504 (N_504,In_1454,In_685);
nand U505 (N_505,N_208,In_376);
or U506 (N_506,In_1115,In_511);
xor U507 (N_507,In_828,In_744);
nor U508 (N_508,In_994,In_335);
and U509 (N_509,In_1065,In_137);
nand U510 (N_510,N_244,In_139);
nand U511 (N_511,In_77,In_874);
or U512 (N_512,N_179,In_736);
or U513 (N_513,In_1074,N_375);
nor U514 (N_514,In_814,N_117);
nor U515 (N_515,In_1382,In_910);
or U516 (N_516,N_171,In_361);
or U517 (N_517,In_492,N_59);
nor U518 (N_518,N_333,In_175);
nor U519 (N_519,N_2,N_184);
xnor U520 (N_520,In_551,In_696);
nor U521 (N_521,In_703,In_1171);
xor U522 (N_522,In_1068,In_211);
nor U523 (N_523,In_460,In_86);
and U524 (N_524,N_272,In_1165);
nand U525 (N_525,N_281,N_10);
nor U526 (N_526,In_383,In_687);
nor U527 (N_527,In_400,N_19);
xnor U528 (N_528,In_153,In_795);
nor U529 (N_529,In_766,In_1042);
and U530 (N_530,In_1322,In_277);
and U531 (N_531,In_853,In_245);
and U532 (N_532,N_386,In_1462);
or U533 (N_533,In_1458,In_465);
xnor U534 (N_534,In_1075,N_207);
nand U535 (N_535,In_1328,N_252);
xnor U536 (N_536,N_135,N_31);
xnor U537 (N_537,In_156,In_823);
nand U538 (N_538,N_68,In_1156);
nor U539 (N_539,In_220,N_219);
nand U540 (N_540,In_454,N_70);
nand U541 (N_541,In_343,In_112);
and U542 (N_542,N_397,In_79);
nand U543 (N_543,In_538,In_1159);
and U544 (N_544,In_391,In_1233);
nand U545 (N_545,In_556,In_440);
nor U546 (N_546,In_1468,In_404);
and U547 (N_547,In_1414,In_1044);
xnor U548 (N_548,N_144,In_14);
and U549 (N_549,In_637,N_234);
and U550 (N_550,In_969,In_706);
or U551 (N_551,In_1027,In_648);
nand U552 (N_552,In_768,In_1146);
or U553 (N_553,In_1169,In_723);
xor U554 (N_554,In_441,In_115);
xor U555 (N_555,N_229,In_204);
or U556 (N_556,In_1439,In_498);
nand U557 (N_557,In_170,In_767);
nand U558 (N_558,In_1209,In_473);
nand U559 (N_559,In_241,In_116);
nor U560 (N_560,In_449,N_343);
and U561 (N_561,In_937,In_341);
and U562 (N_562,N_267,N_57);
and U563 (N_563,N_225,In_477);
xor U564 (N_564,N_328,In_268);
nor U565 (N_565,In_1004,N_294);
and U566 (N_566,In_716,In_531);
nor U567 (N_567,In_1482,In_340);
nand U568 (N_568,In_508,In_831);
nand U569 (N_569,In_120,N_352);
nand U570 (N_570,In_824,In_1232);
or U571 (N_571,N_42,In_199);
nand U572 (N_572,N_354,In_1471);
nor U573 (N_573,In_1063,In_255);
and U574 (N_574,N_203,N_283);
or U575 (N_575,In_924,In_1064);
nand U576 (N_576,In_247,In_1008);
xor U577 (N_577,In_906,In_775);
nand U578 (N_578,N_245,In_109);
xnor U579 (N_579,In_976,In_73);
nand U580 (N_580,In_15,In_1039);
nor U581 (N_581,In_600,In_54);
xnor U582 (N_582,In_1048,In_862);
nor U583 (N_583,In_1358,In_1110);
or U584 (N_584,In_167,In_1069);
nand U585 (N_585,In_536,In_84);
nor U586 (N_586,N_202,In_873);
xor U587 (N_587,In_487,In_1179);
and U588 (N_588,In_3,In_1437);
or U589 (N_589,In_164,In_1404);
or U590 (N_590,N_92,In_360);
and U591 (N_591,In_1126,In_1228);
xor U592 (N_592,In_10,N_60);
xnor U593 (N_593,N_76,In_303);
nor U594 (N_594,In_1459,In_1206);
xor U595 (N_595,N_371,In_395);
xnor U596 (N_596,In_1265,In_564);
nor U597 (N_597,In_1396,In_523);
xor U598 (N_598,N_289,In_500);
nand U599 (N_599,N_307,N_205);
xnor U600 (N_600,In_957,In_920);
or U601 (N_601,In_243,In_1106);
nor U602 (N_602,In_698,In_434);
and U603 (N_603,N_471,N_421);
xnor U604 (N_604,N_104,In_1056);
xnor U605 (N_605,In_493,N_486);
or U606 (N_606,N_541,In_1442);
nand U607 (N_607,In_975,In_602);
nand U608 (N_608,N_9,N_320);
xnor U609 (N_609,N_133,N_107);
xor U610 (N_610,N_206,N_540);
or U611 (N_611,N_359,In_26);
and U612 (N_612,N_150,In_762);
nand U613 (N_613,In_763,N_374);
or U614 (N_614,In_244,In_174);
or U615 (N_615,In_224,In_1483);
nor U616 (N_616,N_263,In_1335);
or U617 (N_617,In_588,In_85);
nor U618 (N_618,In_36,In_374);
nand U619 (N_619,N_85,In_510);
xor U620 (N_620,N_400,N_453);
nand U621 (N_621,N_460,N_293);
or U622 (N_622,N_589,In_700);
nand U623 (N_623,N_1,N_261);
or U624 (N_624,N_362,In_1406);
and U625 (N_625,In_1058,In_161);
nand U626 (N_626,In_372,In_947);
nor U627 (N_627,In_1096,In_143);
or U628 (N_628,In_1263,N_378);
or U629 (N_629,In_1452,N_32);
nand U630 (N_630,In_526,N_548);
and U631 (N_631,N_390,In_1448);
xor U632 (N_632,N_520,In_789);
or U633 (N_633,In_154,N_488);
and U634 (N_634,N_594,N_466);
nor U635 (N_635,N_576,N_3);
xor U636 (N_636,N_90,N_45);
and U637 (N_637,N_236,In_1306);
nor U638 (N_638,In_1445,In_783);
xor U639 (N_639,In_446,N_91);
nor U640 (N_640,In_1278,N_395);
or U641 (N_641,N_191,In_411);
xor U642 (N_642,N_213,In_537);
and U643 (N_643,In_715,N_569);
or U644 (N_644,N_470,In_1248);
or U645 (N_645,In_922,N_50);
or U646 (N_646,In_1311,N_243);
or U647 (N_647,In_804,In_1018);
xnor U648 (N_648,In_631,N_165);
xor U649 (N_649,In_176,N_479);
nor U650 (N_650,N_287,N_585);
and U651 (N_651,N_559,In_60);
nor U652 (N_652,In_1220,In_58);
or U653 (N_653,In_899,In_117);
nor U654 (N_654,N_537,In_963);
nor U655 (N_655,N_431,In_835);
nor U656 (N_656,N_167,In_336);
or U657 (N_657,In_1464,N_210);
nand U658 (N_658,In_1086,N_572);
and U659 (N_659,In_39,N_74);
nand U660 (N_660,In_652,N_278);
nand U661 (N_661,N_458,N_259);
and U662 (N_662,In_1371,N_98);
and U663 (N_663,N_357,N_226);
and U664 (N_664,In_1355,In_867);
and U665 (N_665,In_708,N_393);
nand U666 (N_666,In_408,N_405);
nand U667 (N_667,N_467,In_755);
and U668 (N_668,In_1285,In_1190);
nor U669 (N_669,N_181,N_457);
nor U670 (N_670,N_563,In_349);
and U671 (N_671,In_61,N_310);
xnor U672 (N_672,N_368,N_20);
or U673 (N_673,N_436,N_461);
nor U674 (N_674,N_564,In_547);
or U675 (N_675,N_146,N_529);
and U676 (N_676,N_215,In_1447);
or U677 (N_677,In_1282,In_713);
nand U678 (N_678,In_308,In_1489);
nor U679 (N_679,In_1151,N_577);
nor U680 (N_680,In_406,N_560);
nor U681 (N_681,N_358,N_440);
or U682 (N_682,In_172,N_442);
or U683 (N_683,N_480,In_892);
and U684 (N_684,In_1244,N_543);
and U685 (N_685,In_258,N_450);
xnor U686 (N_686,In_911,N_176);
and U687 (N_687,In_1237,In_578);
nor U688 (N_688,In_1258,In_409);
xor U689 (N_689,N_325,In_1288);
and U690 (N_690,In_1098,In_948);
xor U691 (N_691,In_49,In_1421);
and U692 (N_692,N_175,In_970);
xnor U693 (N_693,N_250,In_482);
or U694 (N_694,N_37,In_567);
nand U695 (N_695,N_62,N_355);
xnor U696 (N_696,N_387,N_493);
nand U697 (N_697,N_329,In_1250);
and U698 (N_698,In_1166,In_1236);
nor U699 (N_699,N_305,N_481);
and U700 (N_700,In_1150,N_553);
or U701 (N_701,In_1182,In_1440);
and U702 (N_702,In_967,In_1195);
nor U703 (N_703,In_88,In_1284);
or U704 (N_704,N_550,N_273);
and U705 (N_705,N_69,In_841);
nor U706 (N_706,N_517,N_126);
and U707 (N_707,N_224,In_797);
nand U708 (N_708,N_597,In_1162);
nand U709 (N_709,In_1324,N_268);
xnor U710 (N_710,In_53,N_437);
or U711 (N_711,In_235,N_413);
and U712 (N_712,In_468,In_601);
nor U713 (N_713,In_1255,N_332);
and U714 (N_714,N_155,In_1393);
xor U715 (N_715,In_1187,N_170);
or U716 (N_716,In_19,In_733);
or U717 (N_717,In_740,In_741);
and U718 (N_718,N_506,N_419);
and U719 (N_719,N_519,In_634);
or U720 (N_720,N_218,N_596);
and U721 (N_721,N_223,In_1341);
nor U722 (N_722,In_1174,In_630);
or U723 (N_723,In_615,N_212);
nand U724 (N_724,N_172,In_625);
and U725 (N_725,N_455,N_504);
or U726 (N_726,In_1214,In_225);
nand U727 (N_727,N_159,N_547);
and U728 (N_728,In_721,N_510);
xnor U729 (N_729,In_1441,In_881);
or U730 (N_730,In_1291,In_589);
and U731 (N_731,N_284,N_415);
or U732 (N_732,In_1243,In_1135);
xnor U733 (N_733,N_396,In_302);
or U734 (N_734,In_262,N_416);
nand U735 (N_735,In_1431,N_385);
nand U736 (N_736,In_1330,In_462);
xor U737 (N_737,N_383,In_618);
and U738 (N_738,In_494,In_956);
or U739 (N_739,In_952,In_339);
xnor U740 (N_740,In_774,N_592);
or U741 (N_741,In_104,In_293);
nor U742 (N_742,In_483,N_446);
nand U743 (N_743,In_193,N_327);
nor U744 (N_744,N_249,N_505);
nand U745 (N_745,In_749,In_357);
or U746 (N_746,In_165,In_504);
nor U747 (N_747,N_290,N_465);
xnor U748 (N_748,In_309,N_468);
or U749 (N_749,In_885,N_314);
xnor U750 (N_750,N_136,In_1427);
or U751 (N_751,N_430,N_337);
or U752 (N_752,N_485,N_306);
xor U753 (N_753,N_435,In_1363);
nor U754 (N_754,N_242,In_1088);
or U755 (N_755,In_27,N_34);
and U756 (N_756,N_591,In_70);
nor U757 (N_757,N_424,N_526);
xor U758 (N_758,In_977,N_570);
nand U759 (N_759,N_80,In_403);
nand U760 (N_760,N_102,In_1380);
xor U761 (N_761,In_787,N_318);
nand U762 (N_762,In_1299,N_562);
and U763 (N_763,In_221,N_401);
or U764 (N_764,In_351,In_1412);
xnor U765 (N_765,In_1130,N_491);
and U766 (N_766,N_507,N_571);
nand U767 (N_767,N_509,In_301);
xnor U768 (N_768,N_459,In_290);
xnor U769 (N_769,In_968,In_1010);
and U770 (N_770,N_501,N_301);
and U771 (N_771,N_469,In_470);
nor U772 (N_772,In_278,N_521);
or U773 (N_773,In_227,N_530);
xor U774 (N_774,N_97,N_285);
or U775 (N_775,In_1073,In_1157);
nor U776 (N_776,N_326,In_289);
xor U777 (N_777,N_366,N_118);
or U778 (N_778,N_351,In_1398);
nand U779 (N_779,In_332,N_418);
or U780 (N_780,In_801,In_834);
nor U781 (N_781,N_316,N_556);
xor U782 (N_782,In_940,In_100);
nor U783 (N_783,In_902,In_1101);
nand U784 (N_784,In_1321,In_124);
and U785 (N_785,N_77,N_511);
nor U786 (N_786,In_1480,N_347);
nor U787 (N_787,N_240,N_257);
nand U788 (N_788,N_180,N_260);
and U789 (N_789,N_404,N_534);
nand U790 (N_790,In_320,In_756);
or U791 (N_791,N_89,In_1223);
xnor U792 (N_792,N_296,N_384);
nand U793 (N_793,In_57,In_780);
xnor U794 (N_794,In_67,In_42);
nand U795 (N_795,In_934,In_1337);
nand U796 (N_796,N_211,In_611);
or U797 (N_797,In_528,N_28);
nand U798 (N_798,In_474,N_12);
or U799 (N_799,In_661,N_531);
nor U800 (N_800,N_699,In_888);
nor U801 (N_801,N_647,In_147);
and U802 (N_802,In_669,In_1147);
xnor U803 (N_803,N_81,N_409);
xor U804 (N_804,In_560,N_747);
nand U805 (N_805,N_376,N_621);
nand U806 (N_806,In_662,N_717);
nand U807 (N_807,N_732,In_344);
nand U808 (N_808,N_715,N_721);
nor U809 (N_809,N_755,N_587);
nor U810 (N_810,N_702,In_9);
nand U811 (N_811,N_496,N_643);
xnor U812 (N_812,In_138,N_489);
and U813 (N_813,In_645,N_113);
and U814 (N_814,N_632,N_779);
xnor U815 (N_815,N_532,N_625);
xnor U816 (N_816,In_270,N_762);
and U817 (N_817,N_546,In_169);
or U818 (N_818,In_887,N_353);
nor U819 (N_819,N_317,In_550);
xor U820 (N_820,N_319,N_123);
nor U821 (N_821,In_833,N_331);
and U822 (N_822,N_775,In_11);
nor U823 (N_823,In_1061,N_300);
or U824 (N_824,N_777,In_1152);
xor U825 (N_825,In_105,In_858);
nor U826 (N_826,N_528,N_513);
or U827 (N_827,N_628,In_517);
nor U828 (N_828,N_372,N_188);
xor U829 (N_829,In_5,N_737);
nor U830 (N_830,In_848,N_653);
xor U831 (N_831,N_369,N_538);
nor U832 (N_832,N_593,In_456);
nand U833 (N_833,N_629,N_238);
xor U834 (N_834,In_229,N_656);
xor U835 (N_835,N_710,In_425);
nor U836 (N_836,N_718,N_739);
xnor U837 (N_837,N_601,In_1052);
nor U838 (N_838,N_429,N_246);
nor U839 (N_839,N_565,N_655);
nor U840 (N_840,In_1167,In_1111);
and U841 (N_841,N_535,In_184);
or U842 (N_842,N_539,N_586);
nor U843 (N_843,N_609,N_462);
and U844 (N_844,N_472,N_120);
and U845 (N_845,N_487,N_708);
xnor U846 (N_846,N_549,In_544);
and U847 (N_847,N_233,In_322);
or U848 (N_848,N_402,In_1373);
nand U849 (N_849,N_668,In_97);
nor U850 (N_850,In_82,N_131);
and U851 (N_851,In_999,N_661);
nand U852 (N_852,N_707,N_686);
nand U853 (N_853,N_361,N_687);
and U854 (N_854,N_663,N_449);
and U855 (N_855,N_473,In_1469);
or U856 (N_856,N_697,N_367);
xnor U857 (N_857,N_566,In_113);
and U858 (N_858,N_638,In_1434);
nand U859 (N_859,N_769,In_205);
and U860 (N_860,In_356,In_921);
nor U861 (N_861,N_125,N_0);
or U862 (N_862,N_714,In_285);
or U863 (N_863,N_654,N_492);
and U864 (N_864,N_474,In_358);
and U865 (N_865,N_247,In_402);
nand U866 (N_866,In_548,In_1113);
or U867 (N_867,N_784,N_610);
nor U868 (N_868,In_123,N_729);
and U869 (N_869,In_586,N_607);
or U870 (N_870,In_103,In_1196);
and U871 (N_871,In_1292,In_33);
xnor U872 (N_872,In_359,In_745);
or U873 (N_873,N_408,In_373);
or U874 (N_874,In_884,N_216);
or U875 (N_875,In_951,In_983);
nand U876 (N_876,In_1303,N_154);
xnor U877 (N_877,In_1155,N_53);
nor U878 (N_878,In_1095,N_99);
xnor U879 (N_879,N_426,In_573);
or U880 (N_880,N_64,N_156);
nor U881 (N_881,N_744,N_24);
and U882 (N_882,N_66,In_1083);
xnor U883 (N_883,N_308,In_577);
xor U884 (N_884,N_787,In_275);
nand U885 (N_885,N_723,In_1369);
xor U886 (N_886,In_861,In_486);
or U887 (N_887,N_776,N_536);
nor U888 (N_888,N_619,N_434);
or U889 (N_889,N_313,N_551);
nand U890 (N_890,N_731,N_799);
nand U891 (N_891,N_603,N_324);
nand U892 (N_892,N_605,N_379);
nand U893 (N_893,In_261,N_758);
nor U894 (N_894,N_753,N_767);
nor U895 (N_895,In_1443,N_399);
or U896 (N_896,N_286,N_693);
or U897 (N_897,N_88,In_543);
and U898 (N_898,N_584,In_959);
nor U899 (N_899,In_371,N_341);
nand U900 (N_900,N_783,In_2);
or U901 (N_901,In_1449,N_574);
xor U902 (N_902,In_321,In_664);
and U903 (N_903,In_826,N_187);
nor U904 (N_904,N_512,N_641);
nor U905 (N_905,N_598,In_4);
nor U906 (N_906,In_63,In_944);
or U907 (N_907,N_667,N_669);
and U908 (N_908,N_676,In_1304);
nand U909 (N_909,In_1408,N_7);
xor U910 (N_910,N_339,In_1235);
nor U911 (N_911,In_1143,N_78);
nor U912 (N_912,N_774,N_620);
or U913 (N_913,N_498,N_524);
nor U914 (N_914,In_859,In_1254);
and U915 (N_915,In_1460,N_626);
nand U916 (N_916,N_691,N_414);
xor U917 (N_917,N_454,N_527);
or U918 (N_918,N_269,N_350);
or U919 (N_919,In_675,In_1474);
nor U920 (N_920,N_642,N_627);
nand U921 (N_921,N_722,N_738);
nor U922 (N_922,N_477,In_282);
nor U923 (N_923,N_750,In_121);
and U924 (N_924,In_1028,N_796);
nand U925 (N_925,In_1364,In_414);
and U926 (N_926,In_1264,N_502);
xnor U927 (N_927,In_778,N_757);
xnor U928 (N_928,N_518,In_1060);
xor U929 (N_929,N_336,In_472);
or U930 (N_930,In_1491,N_433);
nand U931 (N_931,N_407,N_345);
or U932 (N_932,N_611,N_258);
xnor U933 (N_933,N_25,In_222);
xor U934 (N_934,N_599,N_770);
or U935 (N_935,In_1216,N_220);
or U936 (N_936,In_1201,In_1245);
nand U937 (N_937,N_312,In_484);
xnor U938 (N_938,N_636,N_256);
nand U939 (N_939,N_322,In_429);
nand U940 (N_940,In_882,In_17);
nor U941 (N_941,In_171,N_746);
nor U942 (N_942,N_612,N_644);
and U943 (N_943,N_11,N_682);
nand U944 (N_944,N_709,In_604);
nand U945 (N_945,N_748,N_110);
xor U946 (N_946,In_183,N_701);
xor U947 (N_947,N_772,N_795);
and U948 (N_948,N_542,In_532);
and U949 (N_949,In_1386,N_377);
nor U950 (N_950,N_417,N_766);
nand U951 (N_951,N_445,N_595);
and U952 (N_952,N_334,In_1153);
and U953 (N_953,In_1141,N_651);
xor U954 (N_954,N_232,In_230);
and U955 (N_955,In_150,In_1338);
or U956 (N_956,N_143,N_664);
nand U957 (N_957,In_133,N_394);
nor U958 (N_958,N_475,N_615);
nor U959 (N_959,In_1032,N_652);
xnor U960 (N_960,N_786,N_365);
nand U961 (N_961,N_456,N_515);
xnor U962 (N_962,N_782,N_659);
xor U963 (N_963,In_64,In_1014);
and U964 (N_964,In_463,N_160);
xor U965 (N_965,N_742,N_614);
or U966 (N_966,In_178,N_635);
nand U967 (N_967,N_255,N_555);
xor U968 (N_968,N_703,N_391);
or U969 (N_969,N_444,In_44);
and U970 (N_970,N_275,In_1001);
xor U971 (N_971,In_805,In_673);
nand U972 (N_972,N_412,In_490);
nor U973 (N_973,N_484,N_447);
or U974 (N_974,In_1415,In_565);
or U975 (N_975,In_1002,In_1403);
and U976 (N_976,N_792,In_1033);
nor U977 (N_977,N_790,N_734);
or U978 (N_978,In_433,N_427);
nor U979 (N_979,In_307,In_80);
or U980 (N_980,In_603,In_676);
or U981 (N_981,N_428,In_173);
and U982 (N_982,In_776,N_773);
xnor U983 (N_983,In_1262,In_237);
or U984 (N_984,N_670,In_89);
xnor U985 (N_985,N_756,N_389);
and U986 (N_986,In_464,N_558);
xor U987 (N_987,In_562,N_743);
nand U988 (N_988,N_700,N_490);
or U989 (N_989,N_448,N_441);
xor U990 (N_990,N_228,N_43);
xor U991 (N_991,N_705,N_690);
and U992 (N_992,In_1359,N_580);
nor U993 (N_993,N_735,In_585);
and U994 (N_994,N_295,In_1199);
nand U995 (N_995,N_622,In_1210);
and U996 (N_996,N_613,N_335);
xor U997 (N_997,In_1274,In_141);
and U998 (N_998,N_483,N_788);
nor U999 (N_999,In_1120,N_780);
and U1000 (N_1000,N_990,N_124);
or U1001 (N_1001,In_515,N_514);
xor U1002 (N_1002,N_695,N_842);
xor U1003 (N_1003,N_561,N_808);
or U1004 (N_1004,N_898,N_798);
or U1005 (N_1005,N_950,In_1362);
and U1006 (N_1006,In_1484,In_1072);
nand U1007 (N_1007,In_350,N_821);
nand U1008 (N_1008,N_423,N_789);
and U1009 (N_1009,N_494,N_778);
nand U1010 (N_1010,N_646,In_218);
nand U1011 (N_1011,In_1055,N_832);
and U1012 (N_1012,In_1346,In_450);
nand U1013 (N_1013,N_94,In_291);
and U1014 (N_1014,N_829,In_919);
and U1015 (N_1015,N_982,N_552);
and U1016 (N_1016,N_438,N_716);
xor U1017 (N_1017,N_822,N_971);
xnor U1018 (N_1018,N_880,N_73);
nand U1019 (N_1019,In_1444,N_733);
or U1020 (N_1020,N_840,N_523);
or U1021 (N_1021,In_479,N_745);
nor U1022 (N_1022,N_836,N_940);
or U1023 (N_1023,N_724,N_930);
nand U1024 (N_1024,In_753,In_1231);
xnor U1025 (N_1025,N_895,N_955);
xor U1026 (N_1026,N_122,N_874);
xnor U1027 (N_1027,N_711,N_837);
and U1028 (N_1028,In_410,In_405);
nand U1029 (N_1029,N_806,N_403);
and U1030 (N_1030,N_848,N_883);
nor U1031 (N_1031,N_338,N_921);
nor U1032 (N_1032,N_839,N_844);
nor U1033 (N_1033,N_928,N_452);
and U1034 (N_1034,N_973,In_518);
nor U1035 (N_1035,N_857,N_956);
nor U1036 (N_1036,N_740,In_1379);
nand U1037 (N_1037,N_650,N_827);
xnor U1038 (N_1038,N_820,N_533);
or U1039 (N_1039,N_280,N_941);
or U1040 (N_1040,In_682,N_926);
or U1041 (N_1041,N_816,N_925);
xor U1042 (N_1042,N_105,N_896);
or U1043 (N_1043,N_478,In_292);
nand U1044 (N_1044,In_1326,N_960);
and U1045 (N_1045,N_910,In_827);
nand U1046 (N_1046,N_841,N_963);
nand U1047 (N_1047,N_364,N_522);
xnor U1048 (N_1048,N_994,N_680);
nor U1049 (N_1049,In_393,In_705);
nand U1050 (N_1050,In_1019,In_41);
xnor U1051 (N_1051,In_459,In_418);
and U1052 (N_1052,In_1211,N_100);
or U1053 (N_1053,N_819,N_861);
and U1054 (N_1054,N_567,N_128);
xnor U1055 (N_1055,N_761,In_998);
xnor U1056 (N_1056,In_1145,In_720);
xor U1057 (N_1057,N_919,N_516);
and U1058 (N_1058,N_725,N_915);
or U1059 (N_1059,N_942,N_864);
nor U1060 (N_1060,N_791,N_894);
or U1061 (N_1061,N_503,N_649);
or U1062 (N_1062,In_1242,N_932);
and U1063 (N_1063,N_933,N_943);
nor U1064 (N_1064,In_1030,N_616);
nand U1065 (N_1065,In_191,N_913);
and U1066 (N_1066,N_588,In_78);
nor U1067 (N_1067,In_1188,N_917);
xnor U1068 (N_1068,N_859,N_44);
or U1069 (N_1069,N_849,In_197);
xnor U1070 (N_1070,N_58,N_499);
nand U1071 (N_1071,N_557,N_443);
or U1072 (N_1072,In_1290,N_909);
or U1073 (N_1073,N_815,N_858);
xnor U1074 (N_1074,In_288,N_648);
nand U1075 (N_1075,N_831,In_177);
nand U1076 (N_1076,N_508,N_671);
xnor U1077 (N_1077,In_854,N_685);
or U1078 (N_1078,N_949,N_825);
nand U1079 (N_1079,N_974,N_938);
and U1080 (N_1080,N_970,In_1226);
or U1081 (N_1081,In_342,In_1215);
or U1082 (N_1082,N_406,N_838);
nand U1083 (N_1083,N_637,N_771);
and U1084 (N_1084,N_264,In_1164);
xor U1085 (N_1085,N_886,N_119);
or U1086 (N_1086,N_727,In_566);
or U1087 (N_1087,N_579,In_132);
nand U1088 (N_1088,N_677,N_197);
and U1089 (N_1089,N_292,N_988);
nand U1090 (N_1090,N_634,N_869);
nand U1091 (N_1091,N_420,N_851);
xor U1092 (N_1092,N_726,N_807);
and U1093 (N_1093,N_604,N_882);
nor U1094 (N_1094,N_662,N_201);
and U1095 (N_1095,N_954,N_673);
nor U1096 (N_1096,N_482,N_425);
and U1097 (N_1097,N_951,N_168);
nand U1098 (N_1098,N_854,N_253);
xnor U1099 (N_1099,N_980,N_961);
nor U1100 (N_1100,In_1256,N_178);
and U1101 (N_1101,N_760,N_965);
or U1102 (N_1102,In_907,N_765);
nand U1103 (N_1103,In_513,N_763);
or U1104 (N_1104,N_976,N_683);
and U1105 (N_1105,N_730,In_168);
nand U1106 (N_1106,N_907,N_410);
and U1107 (N_1107,In_1318,N_828);
and U1108 (N_1108,N_698,In_1473);
nor U1109 (N_1109,N_814,N_781);
nor U1110 (N_1110,N_958,N_330);
nand U1111 (N_1111,N_794,N_924);
nor U1112 (N_1112,N_889,N_986);
nand U1113 (N_1113,N_65,N_340);
xor U1114 (N_1114,N_853,N_893);
or U1115 (N_1115,In_1370,In_455);
or U1116 (N_1116,N_879,N_871);
and U1117 (N_1117,N_675,N_63);
or U1118 (N_1118,N_997,In_62);
or U1119 (N_1119,N_631,N_860);
nor U1120 (N_1120,N_785,In_37);
xnor U1121 (N_1121,N_602,N_904);
nand U1122 (N_1122,N_749,N_923);
nand U1123 (N_1123,N_759,N_679);
or U1124 (N_1124,In_1297,N_251);
nor U1125 (N_1125,In_739,N_684);
xor U1126 (N_1126,In_1340,N_464);
and U1127 (N_1127,N_497,In_1470);
xor U1128 (N_1128,N_713,In_76);
xnor U1129 (N_1129,N_583,N_138);
and U1130 (N_1130,N_876,N_884);
xnor U1131 (N_1131,N_852,N_797);
nand U1132 (N_1132,N_704,In_1116);
xnor U1133 (N_1133,In_820,In_663);
nand U1134 (N_1134,N_969,N_606);
xnor U1135 (N_1135,N_947,N_983);
nand U1136 (N_1136,In_1419,In_830);
nand U1137 (N_1137,N_692,N_914);
or U1138 (N_1138,N_617,N_495);
nand U1139 (N_1139,In_186,N_500);
xor U1140 (N_1140,In_553,N_935);
xnor U1141 (N_1141,In_1128,N_525);
xnor U1142 (N_1142,N_141,N_900);
or U1143 (N_1143,N_812,N_891);
and U1144 (N_1144,N_169,N_899);
or U1145 (N_1145,In_1418,N_865);
nand U1146 (N_1146,N_934,N_639);
nor U1147 (N_1147,N_948,In_931);
xor U1148 (N_1148,In_1401,N_600);
xor U1149 (N_1149,N_897,N_575);
nor U1150 (N_1150,N_968,In_697);
xnor U1151 (N_1151,N_801,N_217);
xor U1152 (N_1152,N_830,N_811);
nand U1153 (N_1153,N_813,N_998);
nand U1154 (N_1154,N_222,N_186);
nand U1155 (N_1155,In_1189,N_846);
or U1156 (N_1156,N_903,N_902);
nor U1157 (N_1157,N_867,In_299);
nand U1158 (N_1158,N_728,N_981);
or U1159 (N_1159,In_365,N_826);
and U1160 (N_1160,N_411,N_665);
nand U1161 (N_1161,N_381,N_987);
or U1162 (N_1162,N_235,In_533);
and U1163 (N_1163,N_835,N_706);
xor U1164 (N_1164,N_764,In_946);
xnor U1165 (N_1165,In_263,N_922);
xor U1166 (N_1166,N_977,N_872);
and U1167 (N_1167,In_234,In_223);
nor U1168 (N_1168,N_953,N_967);
or U1169 (N_1169,In_1102,N_939);
or U1170 (N_1170,N_199,N_678);
xor U1171 (N_1171,N_254,N_833);
nor U1172 (N_1172,N_630,In_314);
nand U1173 (N_1173,In_1249,N_752);
or U1174 (N_1174,N_996,N_877);
or U1175 (N_1175,N_463,N_863);
nor U1176 (N_1176,N_952,N_696);
or U1177 (N_1177,N_995,In_962);
xor U1178 (N_1178,In_1407,N_937);
xnor U1179 (N_1179,N_875,N_694);
or U1180 (N_1180,In_629,In_443);
or U1181 (N_1181,N_101,N_309);
xor U1182 (N_1182,N_297,In_779);
xnor U1183 (N_1183,In_1212,N_608);
nor U1184 (N_1184,N_802,N_800);
nor U1185 (N_1185,N_422,N_432);
nand U1186 (N_1186,N_342,N_768);
nor U1187 (N_1187,N_972,In_194);
xnor U1188 (N_1188,N_870,N_885);
and U1189 (N_1189,N_658,N_451);
nand U1190 (N_1190,N_810,N_855);
nand U1191 (N_1191,N_873,In_965);
nor U1192 (N_1192,N_911,N_945);
and U1193 (N_1193,N_568,N_590);
and U1194 (N_1194,N_979,In_760);
xnor U1195 (N_1195,N_52,N_581);
nand U1196 (N_1196,N_984,N_736);
and U1197 (N_1197,N_304,In_91);
or U1198 (N_1198,N_298,N_666);
nor U1199 (N_1199,In_385,N_964);
nor U1200 (N_1200,N_1055,N_1033);
nor U1201 (N_1201,N_185,N_623);
or U1202 (N_1202,N_1086,In_1168);
or U1203 (N_1203,N_1198,N_1176);
nor U1204 (N_1204,N_1175,N_1101);
or U1205 (N_1205,N_1188,N_1156);
or U1206 (N_1206,N_1062,N_1074);
or U1207 (N_1207,N_1039,N_1158);
nor U1208 (N_1208,N_1006,N_754);
nand U1209 (N_1209,N_1001,N_975);
xnor U1210 (N_1210,N_1182,N_887);
nor U1211 (N_1211,N_751,N_823);
and U1212 (N_1212,In_187,N_1108);
or U1213 (N_1213,N_1093,N_1098);
and U1214 (N_1214,N_1183,N_1145);
and U1215 (N_1215,N_1149,N_1120);
and U1216 (N_1216,N_1085,In_1416);
or U1217 (N_1217,N_1121,N_862);
nand U1218 (N_1218,N_1030,N_993);
or U1219 (N_1219,N_1007,N_1073);
or U1220 (N_1220,N_1014,N_1009);
or U1221 (N_1221,N_817,N_1087);
or U1222 (N_1222,N_1169,N_1049);
nand U1223 (N_1223,In_489,N_1063);
nor U1224 (N_1224,N_957,N_1137);
nor U1225 (N_1225,N_1119,N_1037);
or U1226 (N_1226,In_1298,N_1047);
and U1227 (N_1227,N_1186,N_1140);
or U1228 (N_1228,N_1181,N_1163);
nand U1229 (N_1229,N_944,N_1032);
or U1230 (N_1230,N_1122,N_927);
or U1231 (N_1231,In_1493,N_809);
or U1232 (N_1232,N_1179,N_1022);
nor U1233 (N_1233,N_1027,N_265);
and U1234 (N_1234,N_1038,N_920);
nand U1235 (N_1235,N_1010,N_1069);
or U1236 (N_1236,N_1150,N_674);
and U1237 (N_1237,In_331,N_1123);
nand U1238 (N_1238,N_1133,N_1003);
xor U1239 (N_1239,N_1161,N_908);
nor U1240 (N_1240,N_1005,N_962);
nor U1241 (N_1241,N_1109,N_1154);
or U1242 (N_1242,N_1167,N_573);
xnor U1243 (N_1243,N_890,N_1065);
and U1244 (N_1244,N_931,N_657);
or U1245 (N_1245,N_1084,N_1050);
or U1246 (N_1246,N_1095,N_1178);
nor U1247 (N_1247,In_1193,In_216);
nor U1248 (N_1248,N_1042,N_929);
nand U1249 (N_1249,N_1015,N_741);
or U1250 (N_1250,N_1185,N_1075);
or U1251 (N_1251,N_1083,N_633);
xor U1252 (N_1252,N_1076,N_834);
or U1253 (N_1253,N_554,N_1096);
or U1254 (N_1254,N_1056,N_1131);
and U1255 (N_1255,N_1000,N_1172);
nand U1256 (N_1256,N_582,N_1193);
and U1257 (N_1257,N_1170,N_1192);
and U1258 (N_1258,N_1045,N_966);
and U1259 (N_1259,N_1148,N_1152);
xnor U1260 (N_1260,In_989,N_1124);
xnor U1261 (N_1261,N_1008,N_1160);
nor U1262 (N_1262,N_850,N_720);
xor U1263 (N_1263,N_1012,In_152);
nand U1264 (N_1264,N_545,N_1088);
xor U1265 (N_1265,N_618,N_1103);
xor U1266 (N_1266,N_892,N_1144);
and U1267 (N_1267,N_1031,N_1190);
or U1268 (N_1268,N_645,N_1051);
or U1269 (N_1269,N_1196,N_805);
and U1270 (N_1270,N_1164,N_991);
nand U1271 (N_1271,N_1147,In_122);
or U1272 (N_1272,N_1128,N_1082);
or U1273 (N_1273,N_689,N_818);
xor U1274 (N_1274,N_1125,N_1048);
nand U1275 (N_1275,N_803,N_901);
and U1276 (N_1276,In_196,N_1028);
nand U1277 (N_1277,N_1094,N_1174);
nor U1278 (N_1278,N_1070,N_1110);
nand U1279 (N_1279,N_1146,N_578);
or U1280 (N_1280,N_1024,N_1004);
and U1281 (N_1281,N_1171,N_1112);
or U1282 (N_1282,N_1080,N_1023);
or U1283 (N_1283,N_1187,N_906);
nor U1284 (N_1284,N_688,N_1113);
nand U1285 (N_1285,N_1043,N_1081);
xnor U1286 (N_1286,N_1162,N_1177);
xnor U1287 (N_1287,N_1115,N_1130);
or U1288 (N_1288,N_1077,N_1194);
xnor U1289 (N_1289,N_1066,N_1138);
nand U1290 (N_1290,N_1016,N_1002);
nand U1291 (N_1291,N_1180,N_221);
and U1292 (N_1292,N_916,N_1114);
nor U1293 (N_1293,N_992,N_1060);
nand U1294 (N_1294,N_999,N_1117);
nor U1295 (N_1295,N_1097,In_142);
xnor U1296 (N_1296,N_1054,N_1091);
nand U1297 (N_1297,N_1199,N_1107);
nor U1298 (N_1298,N_978,N_1026);
nand U1299 (N_1299,N_1139,N_712);
xnor U1300 (N_1300,N_624,N_719);
nand U1301 (N_1301,N_1034,N_51);
xor U1302 (N_1302,N_672,N_1035);
nor U1303 (N_1303,N_1126,N_1078);
and U1304 (N_1304,N_856,N_1025);
and U1305 (N_1305,N_793,In_364);
nor U1306 (N_1306,N_1041,N_1153);
and U1307 (N_1307,N_1099,N_1197);
nand U1308 (N_1308,N_1155,N_1105);
nand U1309 (N_1309,N_1159,N_985);
nand U1310 (N_1310,N_1020,N_129);
nand U1311 (N_1311,N_476,N_1036);
and U1312 (N_1312,N_918,N_1021);
and U1313 (N_1313,N_878,N_1104);
or U1314 (N_1314,N_544,N_1143);
nand U1315 (N_1315,N_959,N_1090);
and U1316 (N_1316,N_1029,N_1151);
xor U1317 (N_1317,N_905,N_1079);
nand U1318 (N_1318,N_1011,N_1071);
nor U1319 (N_1319,N_1013,N_946);
nand U1320 (N_1320,N_1017,N_1106);
or U1321 (N_1321,N_881,N_1195);
or U1322 (N_1322,N_1061,N_1040);
or U1323 (N_1323,N_1165,N_1092);
and U1324 (N_1324,In_1247,N_1132);
nand U1325 (N_1325,N_1191,N_1118);
nor U1326 (N_1326,N_866,N_1184);
nand U1327 (N_1327,In_480,N_1052);
nor U1328 (N_1328,N_1018,N_1019);
nand U1329 (N_1329,N_1134,N_1100);
nand U1330 (N_1330,N_1135,N_439);
nand U1331 (N_1331,N_1072,N_989);
nor U1332 (N_1332,N_804,N_1157);
nor U1333 (N_1333,N_888,N_1116);
nand U1334 (N_1334,N_868,N_1046);
or U1335 (N_1335,N_845,N_1142);
xnor U1336 (N_1336,N_1166,N_936);
or U1337 (N_1337,N_847,N_824);
and U1338 (N_1338,N_1111,N_1136);
or U1339 (N_1339,N_1067,N_843);
xor U1340 (N_1340,N_660,N_1089);
xor U1341 (N_1341,N_1053,N_640);
and U1342 (N_1342,N_1064,N_1189);
or U1343 (N_1343,N_1068,N_681);
and U1344 (N_1344,N_1102,N_1059);
and U1345 (N_1345,N_1129,N_1173);
or U1346 (N_1346,N_1044,N_1168);
nand U1347 (N_1347,N_912,N_1058);
and U1348 (N_1348,N_109,N_1141);
nand U1349 (N_1349,N_1057,N_1127);
nand U1350 (N_1350,N_901,In_489);
or U1351 (N_1351,N_1073,N_918);
xor U1352 (N_1352,N_712,N_1087);
nor U1353 (N_1353,N_1097,N_1196);
nor U1354 (N_1354,N_1081,N_1060);
and U1355 (N_1355,N_1095,N_660);
and U1356 (N_1356,N_936,N_805);
and U1357 (N_1357,N_905,N_1192);
and U1358 (N_1358,N_887,N_1103);
xnor U1359 (N_1359,N_1126,N_1024);
and U1360 (N_1360,N_992,N_1070);
nor U1361 (N_1361,N_578,N_689);
nor U1362 (N_1362,N_1029,N_881);
and U1363 (N_1363,N_1150,N_741);
nand U1364 (N_1364,N_1057,N_1119);
nor U1365 (N_1365,N_1002,N_1174);
and U1366 (N_1366,N_1195,In_364);
nand U1367 (N_1367,N_1185,N_1122);
nand U1368 (N_1368,N_1086,N_803);
nor U1369 (N_1369,N_1013,N_1136);
nor U1370 (N_1370,N_962,N_1117);
xnor U1371 (N_1371,N_823,N_1052);
or U1372 (N_1372,N_751,N_929);
nand U1373 (N_1373,N_845,N_1176);
or U1374 (N_1374,N_544,N_1179);
nand U1375 (N_1375,N_439,N_1011);
nor U1376 (N_1376,N_1075,N_887);
nand U1377 (N_1377,N_847,N_1075);
or U1378 (N_1378,N_1059,N_1029);
nand U1379 (N_1379,N_1160,N_1062);
nand U1380 (N_1380,N_1141,N_1139);
xnor U1381 (N_1381,N_1170,N_809);
or U1382 (N_1382,N_1120,N_843);
nand U1383 (N_1383,In_187,N_843);
nor U1384 (N_1384,N_1012,N_1098);
nor U1385 (N_1385,N_1082,N_1184);
nand U1386 (N_1386,In_989,N_936);
nor U1387 (N_1387,N_1015,N_1032);
or U1388 (N_1388,N_751,N_1075);
nand U1389 (N_1389,N_1080,N_809);
xor U1390 (N_1390,N_1162,N_1059);
and U1391 (N_1391,N_1128,N_51);
xnor U1392 (N_1392,N_862,N_1198);
or U1393 (N_1393,In_364,N_1165);
or U1394 (N_1394,In_152,N_1130);
and U1395 (N_1395,N_1161,In_480);
xor U1396 (N_1396,N_1057,N_1129);
or U1397 (N_1397,In_1247,N_545);
and U1398 (N_1398,N_966,N_1047);
xnor U1399 (N_1399,N_1098,N_1058);
or U1400 (N_1400,N_1354,N_1306);
xnor U1401 (N_1401,N_1372,N_1283);
nand U1402 (N_1402,N_1399,N_1208);
nand U1403 (N_1403,N_1371,N_1266);
and U1404 (N_1404,N_1298,N_1340);
nand U1405 (N_1405,N_1263,N_1308);
and U1406 (N_1406,N_1359,N_1320);
xor U1407 (N_1407,N_1318,N_1336);
or U1408 (N_1408,N_1322,N_1309);
nor U1409 (N_1409,N_1381,N_1316);
xor U1410 (N_1410,N_1343,N_1357);
or U1411 (N_1411,N_1330,N_1366);
and U1412 (N_1412,N_1230,N_1206);
or U1413 (N_1413,N_1284,N_1386);
and U1414 (N_1414,N_1291,N_1204);
and U1415 (N_1415,N_1240,N_1302);
xnor U1416 (N_1416,N_1334,N_1243);
nand U1417 (N_1417,N_1258,N_1325);
and U1418 (N_1418,N_1278,N_1224);
or U1419 (N_1419,N_1254,N_1235);
nor U1420 (N_1420,N_1247,N_1241);
nor U1421 (N_1421,N_1294,N_1317);
nor U1422 (N_1422,N_1290,N_1349);
nand U1423 (N_1423,N_1391,N_1388);
or U1424 (N_1424,N_1233,N_1213);
xor U1425 (N_1425,N_1314,N_1209);
nand U1426 (N_1426,N_1344,N_1389);
or U1427 (N_1427,N_1383,N_1397);
or U1428 (N_1428,N_1212,N_1288);
nand U1429 (N_1429,N_1211,N_1362);
nor U1430 (N_1430,N_1394,N_1356);
and U1431 (N_1431,N_1214,N_1238);
and U1432 (N_1432,N_1202,N_1382);
xor U1433 (N_1433,N_1257,N_1215);
xnor U1434 (N_1434,N_1210,N_1274);
nor U1435 (N_1435,N_1355,N_1228);
or U1436 (N_1436,N_1244,N_1255);
nand U1437 (N_1437,N_1220,N_1368);
xor U1438 (N_1438,N_1326,N_1364);
and U1439 (N_1439,N_1226,N_1269);
or U1440 (N_1440,N_1396,N_1286);
and U1441 (N_1441,N_1239,N_1345);
and U1442 (N_1442,N_1310,N_1221);
or U1443 (N_1443,N_1376,N_1268);
or U1444 (N_1444,N_1271,N_1387);
and U1445 (N_1445,N_1361,N_1207);
nor U1446 (N_1446,N_1232,N_1242);
nor U1447 (N_1447,N_1217,N_1385);
nand U1448 (N_1448,N_1281,N_1335);
and U1449 (N_1449,N_1229,N_1236);
and U1450 (N_1450,N_1327,N_1216);
or U1451 (N_1451,N_1300,N_1259);
nand U1452 (N_1452,N_1350,N_1201);
nor U1453 (N_1453,N_1348,N_1267);
nor U1454 (N_1454,N_1360,N_1223);
xor U1455 (N_1455,N_1313,N_1351);
nor U1456 (N_1456,N_1265,N_1358);
or U1457 (N_1457,N_1338,N_1295);
nand U1458 (N_1458,N_1253,N_1287);
xor U1459 (N_1459,N_1324,N_1378);
nor U1460 (N_1460,N_1252,N_1273);
xnor U1461 (N_1461,N_1332,N_1304);
xnor U1462 (N_1462,N_1393,N_1367);
nand U1463 (N_1463,N_1299,N_1303);
or U1464 (N_1464,N_1374,N_1337);
and U1465 (N_1465,N_1296,N_1363);
and U1466 (N_1466,N_1333,N_1395);
or U1467 (N_1467,N_1312,N_1231);
xor U1468 (N_1468,N_1219,N_1256);
and U1469 (N_1469,N_1237,N_1323);
and U1470 (N_1470,N_1365,N_1275);
and U1471 (N_1471,N_1276,N_1331);
and U1472 (N_1472,N_1342,N_1297);
and U1473 (N_1473,N_1260,N_1264);
and U1474 (N_1474,N_1369,N_1305);
and U1475 (N_1475,N_1321,N_1234);
nor U1476 (N_1476,N_1315,N_1262);
or U1477 (N_1477,N_1270,N_1319);
nor U1478 (N_1478,N_1339,N_1272);
xnor U1479 (N_1479,N_1289,N_1375);
or U1480 (N_1480,N_1329,N_1245);
nor U1481 (N_1481,N_1370,N_1249);
xnor U1482 (N_1482,N_1218,N_1246);
nor U1483 (N_1483,N_1248,N_1377);
or U1484 (N_1484,N_1341,N_1293);
nor U1485 (N_1485,N_1277,N_1353);
nand U1486 (N_1486,N_1301,N_1398);
and U1487 (N_1487,N_1282,N_1261);
nor U1488 (N_1488,N_1222,N_1380);
and U1489 (N_1489,N_1352,N_1205);
nor U1490 (N_1490,N_1251,N_1347);
or U1491 (N_1491,N_1292,N_1227);
and U1492 (N_1492,N_1250,N_1311);
and U1493 (N_1493,N_1225,N_1280);
nor U1494 (N_1494,N_1346,N_1307);
nand U1495 (N_1495,N_1203,N_1285);
xor U1496 (N_1496,N_1200,N_1390);
nor U1497 (N_1497,N_1373,N_1279);
xor U1498 (N_1498,N_1384,N_1379);
and U1499 (N_1499,N_1328,N_1392);
xor U1500 (N_1500,N_1236,N_1281);
xor U1501 (N_1501,N_1383,N_1250);
or U1502 (N_1502,N_1237,N_1216);
nand U1503 (N_1503,N_1349,N_1362);
xnor U1504 (N_1504,N_1305,N_1278);
nor U1505 (N_1505,N_1389,N_1367);
xor U1506 (N_1506,N_1276,N_1355);
xnor U1507 (N_1507,N_1286,N_1360);
and U1508 (N_1508,N_1230,N_1389);
and U1509 (N_1509,N_1388,N_1245);
and U1510 (N_1510,N_1277,N_1287);
nor U1511 (N_1511,N_1287,N_1371);
nand U1512 (N_1512,N_1256,N_1279);
nand U1513 (N_1513,N_1291,N_1237);
and U1514 (N_1514,N_1298,N_1399);
nand U1515 (N_1515,N_1237,N_1268);
xor U1516 (N_1516,N_1280,N_1327);
xnor U1517 (N_1517,N_1233,N_1273);
and U1518 (N_1518,N_1206,N_1323);
nand U1519 (N_1519,N_1276,N_1393);
nand U1520 (N_1520,N_1228,N_1378);
nor U1521 (N_1521,N_1340,N_1388);
and U1522 (N_1522,N_1322,N_1383);
nor U1523 (N_1523,N_1309,N_1272);
or U1524 (N_1524,N_1225,N_1330);
nand U1525 (N_1525,N_1396,N_1212);
or U1526 (N_1526,N_1335,N_1211);
nand U1527 (N_1527,N_1305,N_1274);
and U1528 (N_1528,N_1228,N_1247);
nor U1529 (N_1529,N_1339,N_1239);
xor U1530 (N_1530,N_1290,N_1326);
and U1531 (N_1531,N_1368,N_1337);
and U1532 (N_1532,N_1249,N_1254);
nor U1533 (N_1533,N_1256,N_1275);
nor U1534 (N_1534,N_1363,N_1217);
nor U1535 (N_1535,N_1381,N_1340);
and U1536 (N_1536,N_1339,N_1219);
nand U1537 (N_1537,N_1220,N_1291);
xor U1538 (N_1538,N_1371,N_1387);
and U1539 (N_1539,N_1263,N_1267);
xor U1540 (N_1540,N_1285,N_1213);
nor U1541 (N_1541,N_1214,N_1204);
xor U1542 (N_1542,N_1311,N_1377);
nor U1543 (N_1543,N_1324,N_1257);
and U1544 (N_1544,N_1357,N_1276);
xor U1545 (N_1545,N_1238,N_1360);
nand U1546 (N_1546,N_1213,N_1279);
or U1547 (N_1547,N_1245,N_1338);
xnor U1548 (N_1548,N_1239,N_1229);
xor U1549 (N_1549,N_1278,N_1284);
xnor U1550 (N_1550,N_1394,N_1213);
and U1551 (N_1551,N_1384,N_1269);
nand U1552 (N_1552,N_1335,N_1237);
xor U1553 (N_1553,N_1217,N_1252);
nand U1554 (N_1554,N_1229,N_1387);
nor U1555 (N_1555,N_1305,N_1261);
and U1556 (N_1556,N_1251,N_1393);
xor U1557 (N_1557,N_1259,N_1248);
nor U1558 (N_1558,N_1278,N_1354);
xnor U1559 (N_1559,N_1270,N_1217);
nor U1560 (N_1560,N_1385,N_1231);
xnor U1561 (N_1561,N_1301,N_1254);
or U1562 (N_1562,N_1345,N_1251);
xor U1563 (N_1563,N_1284,N_1291);
and U1564 (N_1564,N_1370,N_1208);
xor U1565 (N_1565,N_1340,N_1365);
nor U1566 (N_1566,N_1327,N_1390);
and U1567 (N_1567,N_1210,N_1287);
nand U1568 (N_1568,N_1399,N_1363);
nor U1569 (N_1569,N_1279,N_1226);
or U1570 (N_1570,N_1241,N_1211);
xor U1571 (N_1571,N_1253,N_1250);
nand U1572 (N_1572,N_1220,N_1261);
nor U1573 (N_1573,N_1204,N_1215);
nand U1574 (N_1574,N_1223,N_1257);
nor U1575 (N_1575,N_1348,N_1359);
nand U1576 (N_1576,N_1235,N_1261);
xor U1577 (N_1577,N_1221,N_1372);
nand U1578 (N_1578,N_1251,N_1255);
and U1579 (N_1579,N_1380,N_1356);
and U1580 (N_1580,N_1366,N_1206);
nand U1581 (N_1581,N_1354,N_1375);
and U1582 (N_1582,N_1339,N_1215);
xor U1583 (N_1583,N_1252,N_1390);
xnor U1584 (N_1584,N_1205,N_1277);
and U1585 (N_1585,N_1398,N_1352);
nor U1586 (N_1586,N_1222,N_1399);
and U1587 (N_1587,N_1309,N_1204);
and U1588 (N_1588,N_1240,N_1306);
and U1589 (N_1589,N_1399,N_1214);
and U1590 (N_1590,N_1327,N_1373);
and U1591 (N_1591,N_1368,N_1350);
nor U1592 (N_1592,N_1211,N_1238);
or U1593 (N_1593,N_1332,N_1278);
or U1594 (N_1594,N_1324,N_1276);
nor U1595 (N_1595,N_1388,N_1279);
nand U1596 (N_1596,N_1287,N_1351);
or U1597 (N_1597,N_1272,N_1266);
nor U1598 (N_1598,N_1272,N_1383);
nor U1599 (N_1599,N_1216,N_1382);
or U1600 (N_1600,N_1591,N_1455);
nand U1601 (N_1601,N_1446,N_1562);
xnor U1602 (N_1602,N_1467,N_1571);
xnor U1603 (N_1603,N_1484,N_1550);
xor U1604 (N_1604,N_1542,N_1423);
and U1605 (N_1605,N_1464,N_1470);
nand U1606 (N_1606,N_1449,N_1521);
xnor U1607 (N_1607,N_1556,N_1437);
xor U1608 (N_1608,N_1412,N_1445);
or U1609 (N_1609,N_1472,N_1414);
nor U1610 (N_1610,N_1428,N_1590);
or U1611 (N_1611,N_1430,N_1485);
and U1612 (N_1612,N_1543,N_1536);
xnor U1613 (N_1613,N_1429,N_1501);
nand U1614 (N_1614,N_1422,N_1535);
nor U1615 (N_1615,N_1481,N_1490);
nand U1616 (N_1616,N_1496,N_1400);
nand U1617 (N_1617,N_1581,N_1456);
or U1618 (N_1618,N_1506,N_1584);
or U1619 (N_1619,N_1463,N_1447);
nand U1620 (N_1620,N_1586,N_1576);
or U1621 (N_1621,N_1408,N_1596);
or U1622 (N_1622,N_1440,N_1554);
or U1623 (N_1623,N_1419,N_1523);
xor U1624 (N_1624,N_1413,N_1541);
nand U1625 (N_1625,N_1459,N_1431);
and U1626 (N_1626,N_1478,N_1540);
or U1627 (N_1627,N_1493,N_1451);
nor U1628 (N_1628,N_1469,N_1508);
nand U1629 (N_1629,N_1551,N_1417);
nand U1630 (N_1630,N_1516,N_1595);
or U1631 (N_1631,N_1533,N_1570);
or U1632 (N_1632,N_1473,N_1477);
xor U1633 (N_1633,N_1534,N_1424);
nand U1634 (N_1634,N_1404,N_1442);
or U1635 (N_1635,N_1439,N_1402);
and U1636 (N_1636,N_1486,N_1525);
xnor U1637 (N_1637,N_1582,N_1465);
nor U1638 (N_1638,N_1528,N_1436);
or U1639 (N_1639,N_1460,N_1583);
or U1640 (N_1640,N_1507,N_1409);
nand U1641 (N_1641,N_1432,N_1443);
xnor U1642 (N_1642,N_1433,N_1574);
xnor U1643 (N_1643,N_1580,N_1509);
or U1644 (N_1644,N_1549,N_1587);
nand U1645 (N_1645,N_1558,N_1572);
xnor U1646 (N_1646,N_1401,N_1559);
and U1647 (N_1647,N_1526,N_1524);
xnor U1648 (N_1648,N_1548,N_1598);
and U1649 (N_1649,N_1427,N_1519);
xnor U1650 (N_1650,N_1561,N_1483);
nand U1651 (N_1651,N_1421,N_1527);
and U1652 (N_1652,N_1530,N_1438);
nor U1653 (N_1653,N_1546,N_1539);
nand U1654 (N_1654,N_1471,N_1579);
nand U1655 (N_1655,N_1488,N_1515);
nor U1656 (N_1656,N_1480,N_1599);
or U1657 (N_1657,N_1563,N_1538);
or U1658 (N_1658,N_1499,N_1434);
xnor U1659 (N_1659,N_1479,N_1453);
xor U1660 (N_1660,N_1510,N_1594);
and U1661 (N_1661,N_1593,N_1537);
nor U1662 (N_1662,N_1411,N_1588);
and U1663 (N_1663,N_1466,N_1575);
or U1664 (N_1664,N_1457,N_1512);
nor U1665 (N_1665,N_1448,N_1529);
and U1666 (N_1666,N_1544,N_1518);
nand U1667 (N_1667,N_1491,N_1407);
and U1668 (N_1668,N_1415,N_1597);
nand U1669 (N_1669,N_1566,N_1435);
nand U1670 (N_1670,N_1452,N_1441);
and U1671 (N_1671,N_1405,N_1568);
and U1672 (N_1672,N_1592,N_1560);
nand U1673 (N_1673,N_1557,N_1418);
nand U1674 (N_1674,N_1450,N_1474);
or U1675 (N_1675,N_1578,N_1454);
nand U1676 (N_1676,N_1468,N_1520);
nand U1677 (N_1677,N_1564,N_1555);
xor U1678 (N_1678,N_1406,N_1545);
nor U1679 (N_1679,N_1553,N_1410);
nor U1680 (N_1680,N_1497,N_1502);
xnor U1681 (N_1681,N_1589,N_1476);
nand U1682 (N_1682,N_1416,N_1425);
or U1683 (N_1683,N_1492,N_1514);
nand U1684 (N_1684,N_1577,N_1503);
or U1685 (N_1685,N_1522,N_1585);
nand U1686 (N_1686,N_1495,N_1504);
or U1687 (N_1687,N_1482,N_1426);
xnor U1688 (N_1688,N_1444,N_1517);
or U1689 (N_1689,N_1500,N_1475);
xor U1690 (N_1690,N_1552,N_1487);
and U1691 (N_1691,N_1403,N_1573);
and U1692 (N_1692,N_1569,N_1567);
or U1693 (N_1693,N_1505,N_1420);
xnor U1694 (N_1694,N_1462,N_1498);
or U1695 (N_1695,N_1513,N_1489);
or U1696 (N_1696,N_1547,N_1461);
and U1697 (N_1697,N_1494,N_1565);
and U1698 (N_1698,N_1532,N_1511);
or U1699 (N_1699,N_1531,N_1458);
and U1700 (N_1700,N_1433,N_1577);
nor U1701 (N_1701,N_1429,N_1531);
and U1702 (N_1702,N_1509,N_1494);
nor U1703 (N_1703,N_1466,N_1464);
nor U1704 (N_1704,N_1592,N_1426);
or U1705 (N_1705,N_1424,N_1552);
nand U1706 (N_1706,N_1565,N_1558);
xor U1707 (N_1707,N_1508,N_1569);
xor U1708 (N_1708,N_1448,N_1482);
and U1709 (N_1709,N_1558,N_1440);
and U1710 (N_1710,N_1586,N_1439);
xor U1711 (N_1711,N_1599,N_1529);
nand U1712 (N_1712,N_1432,N_1533);
xnor U1713 (N_1713,N_1472,N_1526);
or U1714 (N_1714,N_1595,N_1472);
nand U1715 (N_1715,N_1551,N_1469);
nand U1716 (N_1716,N_1460,N_1512);
or U1717 (N_1717,N_1515,N_1421);
and U1718 (N_1718,N_1464,N_1489);
or U1719 (N_1719,N_1425,N_1423);
nor U1720 (N_1720,N_1494,N_1431);
nand U1721 (N_1721,N_1534,N_1423);
nor U1722 (N_1722,N_1458,N_1581);
or U1723 (N_1723,N_1570,N_1561);
or U1724 (N_1724,N_1461,N_1505);
and U1725 (N_1725,N_1456,N_1542);
xor U1726 (N_1726,N_1465,N_1572);
or U1727 (N_1727,N_1574,N_1427);
nor U1728 (N_1728,N_1452,N_1420);
nand U1729 (N_1729,N_1576,N_1578);
or U1730 (N_1730,N_1507,N_1476);
nor U1731 (N_1731,N_1437,N_1525);
xor U1732 (N_1732,N_1589,N_1424);
nor U1733 (N_1733,N_1477,N_1467);
xnor U1734 (N_1734,N_1461,N_1566);
nor U1735 (N_1735,N_1592,N_1528);
xor U1736 (N_1736,N_1584,N_1556);
xnor U1737 (N_1737,N_1500,N_1599);
nand U1738 (N_1738,N_1598,N_1448);
nor U1739 (N_1739,N_1504,N_1430);
or U1740 (N_1740,N_1536,N_1572);
nor U1741 (N_1741,N_1495,N_1568);
or U1742 (N_1742,N_1571,N_1586);
and U1743 (N_1743,N_1416,N_1522);
or U1744 (N_1744,N_1480,N_1455);
nor U1745 (N_1745,N_1535,N_1556);
nor U1746 (N_1746,N_1412,N_1557);
nand U1747 (N_1747,N_1546,N_1564);
xor U1748 (N_1748,N_1504,N_1507);
or U1749 (N_1749,N_1565,N_1495);
xor U1750 (N_1750,N_1561,N_1592);
xor U1751 (N_1751,N_1573,N_1425);
nor U1752 (N_1752,N_1512,N_1569);
or U1753 (N_1753,N_1515,N_1445);
xor U1754 (N_1754,N_1419,N_1437);
nor U1755 (N_1755,N_1571,N_1431);
nand U1756 (N_1756,N_1455,N_1599);
and U1757 (N_1757,N_1554,N_1583);
and U1758 (N_1758,N_1413,N_1457);
and U1759 (N_1759,N_1524,N_1406);
nor U1760 (N_1760,N_1475,N_1430);
or U1761 (N_1761,N_1457,N_1542);
or U1762 (N_1762,N_1575,N_1461);
xor U1763 (N_1763,N_1572,N_1555);
xor U1764 (N_1764,N_1551,N_1463);
and U1765 (N_1765,N_1591,N_1450);
or U1766 (N_1766,N_1549,N_1533);
xnor U1767 (N_1767,N_1415,N_1479);
nor U1768 (N_1768,N_1561,N_1544);
or U1769 (N_1769,N_1457,N_1543);
and U1770 (N_1770,N_1451,N_1446);
xnor U1771 (N_1771,N_1553,N_1520);
and U1772 (N_1772,N_1550,N_1449);
or U1773 (N_1773,N_1539,N_1433);
nor U1774 (N_1774,N_1484,N_1402);
nor U1775 (N_1775,N_1525,N_1401);
or U1776 (N_1776,N_1525,N_1447);
nand U1777 (N_1777,N_1434,N_1521);
xor U1778 (N_1778,N_1555,N_1583);
and U1779 (N_1779,N_1411,N_1427);
nand U1780 (N_1780,N_1462,N_1583);
and U1781 (N_1781,N_1556,N_1447);
xor U1782 (N_1782,N_1431,N_1456);
and U1783 (N_1783,N_1536,N_1595);
and U1784 (N_1784,N_1425,N_1527);
nand U1785 (N_1785,N_1518,N_1439);
xnor U1786 (N_1786,N_1445,N_1534);
and U1787 (N_1787,N_1448,N_1545);
and U1788 (N_1788,N_1582,N_1477);
xnor U1789 (N_1789,N_1464,N_1408);
or U1790 (N_1790,N_1488,N_1587);
nor U1791 (N_1791,N_1528,N_1456);
or U1792 (N_1792,N_1490,N_1498);
nor U1793 (N_1793,N_1558,N_1447);
nor U1794 (N_1794,N_1493,N_1498);
or U1795 (N_1795,N_1413,N_1588);
nand U1796 (N_1796,N_1539,N_1543);
nor U1797 (N_1797,N_1447,N_1533);
and U1798 (N_1798,N_1407,N_1580);
nor U1799 (N_1799,N_1572,N_1442);
and U1800 (N_1800,N_1672,N_1678);
xnor U1801 (N_1801,N_1706,N_1743);
nor U1802 (N_1802,N_1606,N_1659);
nor U1803 (N_1803,N_1708,N_1753);
nand U1804 (N_1804,N_1602,N_1693);
nor U1805 (N_1805,N_1728,N_1699);
nand U1806 (N_1806,N_1795,N_1788);
nor U1807 (N_1807,N_1636,N_1700);
or U1808 (N_1808,N_1628,N_1662);
xor U1809 (N_1809,N_1610,N_1658);
and U1810 (N_1810,N_1644,N_1749);
nor U1811 (N_1811,N_1718,N_1710);
nand U1812 (N_1812,N_1782,N_1769);
or U1813 (N_1813,N_1637,N_1676);
nand U1814 (N_1814,N_1740,N_1737);
xnor U1815 (N_1815,N_1721,N_1746);
nand U1816 (N_1816,N_1609,N_1686);
nand U1817 (N_1817,N_1777,N_1695);
nand U1818 (N_1818,N_1652,N_1622);
or U1819 (N_1819,N_1705,N_1729);
xnor U1820 (N_1820,N_1698,N_1771);
and U1821 (N_1821,N_1768,N_1781);
nor U1822 (N_1822,N_1685,N_1641);
or U1823 (N_1823,N_1717,N_1601);
xor U1824 (N_1824,N_1635,N_1785);
or U1825 (N_1825,N_1611,N_1660);
and U1826 (N_1826,N_1664,N_1724);
or U1827 (N_1827,N_1701,N_1713);
nor U1828 (N_1828,N_1666,N_1655);
and U1829 (N_1829,N_1793,N_1742);
nand U1830 (N_1830,N_1689,N_1703);
xnor U1831 (N_1831,N_1677,N_1603);
nand U1832 (N_1832,N_1744,N_1670);
and U1833 (N_1833,N_1620,N_1779);
nor U1834 (N_1834,N_1735,N_1646);
nand U1835 (N_1835,N_1605,N_1764);
nand U1836 (N_1836,N_1702,N_1684);
nor U1837 (N_1837,N_1600,N_1680);
or U1838 (N_1838,N_1778,N_1661);
or U1839 (N_1839,N_1757,N_1725);
and U1840 (N_1840,N_1648,N_1651);
and U1841 (N_1841,N_1714,N_1668);
xnor U1842 (N_1842,N_1681,N_1691);
nor U1843 (N_1843,N_1650,N_1607);
or U1844 (N_1844,N_1712,N_1615);
nand U1845 (N_1845,N_1716,N_1747);
xnor U1846 (N_1846,N_1707,N_1623);
nor U1847 (N_1847,N_1687,N_1625);
xor U1848 (N_1848,N_1791,N_1745);
or U1849 (N_1849,N_1783,N_1673);
and U1850 (N_1850,N_1794,N_1624);
nor U1851 (N_1851,N_1629,N_1604);
nand U1852 (N_1852,N_1682,N_1733);
nor U1853 (N_1853,N_1762,N_1739);
nand U1854 (N_1854,N_1734,N_1690);
and U1855 (N_1855,N_1760,N_1797);
nand U1856 (N_1856,N_1627,N_1649);
and U1857 (N_1857,N_1674,N_1723);
and U1858 (N_1858,N_1616,N_1633);
nand U1859 (N_1859,N_1763,N_1715);
nand U1860 (N_1860,N_1752,N_1748);
nor U1861 (N_1861,N_1639,N_1799);
nand U1862 (N_1862,N_1730,N_1675);
nand U1863 (N_1863,N_1770,N_1772);
and U1864 (N_1864,N_1653,N_1726);
nor U1865 (N_1865,N_1694,N_1786);
and U1866 (N_1866,N_1640,N_1741);
xnor U1867 (N_1867,N_1732,N_1767);
or U1868 (N_1868,N_1711,N_1665);
and U1869 (N_1869,N_1618,N_1631);
and U1870 (N_1870,N_1679,N_1758);
nand U1871 (N_1871,N_1789,N_1643);
xnor U1872 (N_1872,N_1619,N_1796);
xnor U1873 (N_1873,N_1780,N_1663);
or U1874 (N_1874,N_1671,N_1765);
nor U1875 (N_1875,N_1634,N_1656);
or U1876 (N_1876,N_1642,N_1654);
nor U1877 (N_1877,N_1759,N_1755);
xor U1878 (N_1878,N_1683,N_1614);
nor U1879 (N_1879,N_1696,N_1756);
xnor U1880 (N_1880,N_1657,N_1688);
and U1881 (N_1881,N_1638,N_1784);
xnor U1882 (N_1882,N_1612,N_1632);
nor U1883 (N_1883,N_1754,N_1751);
or U1884 (N_1884,N_1738,N_1719);
xor U1885 (N_1885,N_1761,N_1626);
nor U1886 (N_1886,N_1630,N_1720);
xnor U1887 (N_1887,N_1667,N_1775);
or U1888 (N_1888,N_1645,N_1727);
nand U1889 (N_1889,N_1647,N_1776);
nor U1890 (N_1890,N_1669,N_1704);
or U1891 (N_1891,N_1621,N_1697);
xor U1892 (N_1892,N_1617,N_1731);
nor U1893 (N_1893,N_1766,N_1787);
and U1894 (N_1894,N_1773,N_1790);
nand U1895 (N_1895,N_1792,N_1722);
xnor U1896 (N_1896,N_1692,N_1798);
and U1897 (N_1897,N_1613,N_1709);
xnor U1898 (N_1898,N_1774,N_1750);
nand U1899 (N_1899,N_1736,N_1608);
and U1900 (N_1900,N_1628,N_1631);
xnor U1901 (N_1901,N_1787,N_1622);
nand U1902 (N_1902,N_1745,N_1624);
and U1903 (N_1903,N_1793,N_1711);
xnor U1904 (N_1904,N_1689,N_1604);
or U1905 (N_1905,N_1649,N_1689);
nand U1906 (N_1906,N_1751,N_1623);
and U1907 (N_1907,N_1740,N_1728);
and U1908 (N_1908,N_1754,N_1702);
nand U1909 (N_1909,N_1644,N_1759);
xnor U1910 (N_1910,N_1739,N_1661);
or U1911 (N_1911,N_1665,N_1602);
nand U1912 (N_1912,N_1711,N_1619);
nand U1913 (N_1913,N_1608,N_1664);
nor U1914 (N_1914,N_1706,N_1737);
and U1915 (N_1915,N_1640,N_1632);
xor U1916 (N_1916,N_1654,N_1748);
xor U1917 (N_1917,N_1662,N_1706);
xnor U1918 (N_1918,N_1741,N_1674);
nand U1919 (N_1919,N_1742,N_1772);
nand U1920 (N_1920,N_1693,N_1798);
nor U1921 (N_1921,N_1728,N_1628);
nand U1922 (N_1922,N_1735,N_1607);
xor U1923 (N_1923,N_1611,N_1694);
nand U1924 (N_1924,N_1773,N_1764);
nor U1925 (N_1925,N_1629,N_1650);
xnor U1926 (N_1926,N_1609,N_1794);
xor U1927 (N_1927,N_1721,N_1781);
xnor U1928 (N_1928,N_1760,N_1733);
xor U1929 (N_1929,N_1636,N_1742);
nor U1930 (N_1930,N_1667,N_1702);
and U1931 (N_1931,N_1649,N_1673);
nor U1932 (N_1932,N_1628,N_1743);
nor U1933 (N_1933,N_1673,N_1661);
and U1934 (N_1934,N_1628,N_1685);
nor U1935 (N_1935,N_1769,N_1707);
nor U1936 (N_1936,N_1645,N_1785);
nand U1937 (N_1937,N_1794,N_1647);
xor U1938 (N_1938,N_1689,N_1738);
and U1939 (N_1939,N_1735,N_1672);
nor U1940 (N_1940,N_1778,N_1631);
and U1941 (N_1941,N_1604,N_1770);
nor U1942 (N_1942,N_1695,N_1749);
nor U1943 (N_1943,N_1605,N_1652);
xnor U1944 (N_1944,N_1728,N_1760);
xnor U1945 (N_1945,N_1646,N_1728);
and U1946 (N_1946,N_1698,N_1631);
nand U1947 (N_1947,N_1631,N_1780);
and U1948 (N_1948,N_1694,N_1645);
xor U1949 (N_1949,N_1612,N_1719);
nand U1950 (N_1950,N_1619,N_1649);
nand U1951 (N_1951,N_1773,N_1625);
nand U1952 (N_1952,N_1772,N_1783);
nand U1953 (N_1953,N_1713,N_1605);
nor U1954 (N_1954,N_1618,N_1738);
nor U1955 (N_1955,N_1768,N_1676);
nand U1956 (N_1956,N_1745,N_1636);
xor U1957 (N_1957,N_1770,N_1709);
and U1958 (N_1958,N_1767,N_1779);
nand U1959 (N_1959,N_1768,N_1701);
nand U1960 (N_1960,N_1622,N_1657);
and U1961 (N_1961,N_1790,N_1798);
nor U1962 (N_1962,N_1634,N_1606);
or U1963 (N_1963,N_1690,N_1614);
xnor U1964 (N_1964,N_1713,N_1751);
and U1965 (N_1965,N_1776,N_1741);
xnor U1966 (N_1966,N_1749,N_1785);
and U1967 (N_1967,N_1792,N_1791);
xor U1968 (N_1968,N_1799,N_1780);
nand U1969 (N_1969,N_1663,N_1677);
and U1970 (N_1970,N_1605,N_1791);
nand U1971 (N_1971,N_1721,N_1785);
nand U1972 (N_1972,N_1607,N_1783);
xor U1973 (N_1973,N_1752,N_1718);
and U1974 (N_1974,N_1746,N_1731);
or U1975 (N_1975,N_1702,N_1641);
xor U1976 (N_1976,N_1707,N_1751);
nor U1977 (N_1977,N_1625,N_1743);
nor U1978 (N_1978,N_1621,N_1681);
xor U1979 (N_1979,N_1763,N_1624);
xor U1980 (N_1980,N_1741,N_1612);
or U1981 (N_1981,N_1718,N_1769);
nand U1982 (N_1982,N_1763,N_1682);
and U1983 (N_1983,N_1772,N_1686);
or U1984 (N_1984,N_1767,N_1730);
xor U1985 (N_1985,N_1677,N_1794);
nand U1986 (N_1986,N_1622,N_1634);
xnor U1987 (N_1987,N_1680,N_1765);
xnor U1988 (N_1988,N_1652,N_1640);
xnor U1989 (N_1989,N_1685,N_1781);
xor U1990 (N_1990,N_1782,N_1733);
nor U1991 (N_1991,N_1694,N_1746);
nand U1992 (N_1992,N_1716,N_1630);
and U1993 (N_1993,N_1629,N_1607);
nand U1994 (N_1994,N_1603,N_1660);
xnor U1995 (N_1995,N_1756,N_1672);
nand U1996 (N_1996,N_1779,N_1694);
or U1997 (N_1997,N_1795,N_1793);
or U1998 (N_1998,N_1614,N_1768);
and U1999 (N_1999,N_1721,N_1678);
xnor U2000 (N_2000,N_1837,N_1976);
and U2001 (N_2001,N_1918,N_1978);
xor U2002 (N_2002,N_1925,N_1800);
or U2003 (N_2003,N_1871,N_1984);
xor U2004 (N_2004,N_1970,N_1852);
nand U2005 (N_2005,N_1945,N_1895);
xor U2006 (N_2006,N_1855,N_1841);
and U2007 (N_2007,N_1924,N_1839);
nand U2008 (N_2008,N_1894,N_1883);
nand U2009 (N_2009,N_1816,N_1957);
and U2010 (N_2010,N_1849,N_1864);
nor U2011 (N_2011,N_1949,N_1915);
or U2012 (N_2012,N_1926,N_1817);
or U2013 (N_2013,N_1827,N_1884);
xor U2014 (N_2014,N_1873,N_1810);
nor U2015 (N_2015,N_1980,N_1927);
nor U2016 (N_2016,N_1821,N_1846);
and U2017 (N_2017,N_1826,N_1994);
and U2018 (N_2018,N_1813,N_1922);
or U2019 (N_2019,N_1805,N_1896);
and U2020 (N_2020,N_1997,N_1844);
and U2021 (N_2021,N_1907,N_1989);
and U2022 (N_2022,N_1964,N_1876);
or U2023 (N_2023,N_1850,N_1904);
nand U2024 (N_2024,N_1912,N_1858);
nor U2025 (N_2025,N_1863,N_1906);
nand U2026 (N_2026,N_1804,N_1866);
xor U2027 (N_2027,N_1962,N_1942);
nand U2028 (N_2028,N_1809,N_1938);
or U2029 (N_2029,N_1992,N_1958);
nor U2030 (N_2030,N_1985,N_1899);
and U2031 (N_2031,N_1998,N_1819);
nor U2032 (N_2032,N_1947,N_1930);
and U2033 (N_2033,N_1851,N_1865);
and U2034 (N_2034,N_1908,N_1857);
nand U2035 (N_2035,N_1937,N_1854);
and U2036 (N_2036,N_1859,N_1950);
nor U2037 (N_2037,N_1961,N_1983);
nor U2038 (N_2038,N_1869,N_1903);
and U2039 (N_2039,N_1982,N_1888);
nor U2040 (N_2040,N_1952,N_1956);
and U2041 (N_2041,N_1823,N_1902);
nor U2042 (N_2042,N_1843,N_1975);
xnor U2043 (N_2043,N_1890,N_1909);
xnor U2044 (N_2044,N_1905,N_1911);
nor U2045 (N_2045,N_1808,N_1954);
or U2046 (N_2046,N_1987,N_1879);
nand U2047 (N_2047,N_1979,N_1824);
xnor U2048 (N_2048,N_1928,N_1867);
nor U2049 (N_2049,N_1814,N_1878);
xnor U2050 (N_2050,N_1932,N_1969);
xor U2051 (N_2051,N_1886,N_1960);
or U2052 (N_2052,N_1959,N_1936);
nor U2053 (N_2053,N_1948,N_1872);
and U2054 (N_2054,N_1853,N_1919);
nor U2055 (N_2055,N_1933,N_1973);
or U2056 (N_2056,N_1900,N_1941);
nand U2057 (N_2057,N_1955,N_1893);
nor U2058 (N_2058,N_1995,N_1934);
nor U2059 (N_2059,N_1860,N_1881);
nor U2060 (N_2060,N_1972,N_1921);
nor U2061 (N_2061,N_1870,N_1953);
or U2062 (N_2062,N_1977,N_1812);
and U2063 (N_2063,N_1929,N_1848);
xor U2064 (N_2064,N_1920,N_1874);
xor U2065 (N_2065,N_1991,N_1963);
nor U2066 (N_2066,N_1830,N_1861);
xor U2067 (N_2067,N_1939,N_1910);
xor U2068 (N_2068,N_1981,N_1845);
nand U2069 (N_2069,N_1880,N_1840);
or U2070 (N_2070,N_1965,N_1967);
xnor U2071 (N_2071,N_1811,N_1868);
and U2072 (N_2072,N_1885,N_1974);
nor U2073 (N_2073,N_1806,N_1877);
or U2074 (N_2074,N_1931,N_1951);
or U2075 (N_2075,N_1847,N_1986);
nor U2076 (N_2076,N_1897,N_1943);
and U2077 (N_2077,N_1901,N_1916);
nor U2078 (N_2078,N_1828,N_1835);
nand U2079 (N_2079,N_1968,N_1803);
or U2080 (N_2080,N_1836,N_1875);
nand U2081 (N_2081,N_1940,N_1807);
and U2082 (N_2082,N_1913,N_1882);
xnor U2083 (N_2083,N_1802,N_1822);
or U2084 (N_2084,N_1988,N_1834);
or U2085 (N_2085,N_1898,N_1971);
and U2086 (N_2086,N_1944,N_1917);
nor U2087 (N_2087,N_1946,N_1889);
nor U2088 (N_2088,N_1990,N_1829);
and U2089 (N_2089,N_1838,N_1825);
xor U2090 (N_2090,N_1801,N_1892);
or U2091 (N_2091,N_1923,N_1862);
xor U2092 (N_2092,N_1831,N_1999);
nor U2093 (N_2093,N_1856,N_1914);
or U2094 (N_2094,N_1820,N_1832);
and U2095 (N_2095,N_1935,N_1815);
nor U2096 (N_2096,N_1887,N_1993);
and U2097 (N_2097,N_1966,N_1842);
or U2098 (N_2098,N_1818,N_1833);
or U2099 (N_2099,N_1996,N_1891);
or U2100 (N_2100,N_1882,N_1983);
or U2101 (N_2101,N_1839,N_1838);
nand U2102 (N_2102,N_1807,N_1969);
and U2103 (N_2103,N_1891,N_1897);
and U2104 (N_2104,N_1980,N_1991);
nor U2105 (N_2105,N_1987,N_1954);
or U2106 (N_2106,N_1851,N_1811);
nor U2107 (N_2107,N_1916,N_1858);
nor U2108 (N_2108,N_1865,N_1838);
nor U2109 (N_2109,N_1970,N_1864);
nor U2110 (N_2110,N_1882,N_1855);
xnor U2111 (N_2111,N_1828,N_1886);
nor U2112 (N_2112,N_1900,N_1928);
and U2113 (N_2113,N_1861,N_1811);
nor U2114 (N_2114,N_1920,N_1902);
nor U2115 (N_2115,N_1807,N_1811);
xnor U2116 (N_2116,N_1911,N_1987);
or U2117 (N_2117,N_1896,N_1819);
nand U2118 (N_2118,N_1966,N_1910);
nand U2119 (N_2119,N_1838,N_1854);
xor U2120 (N_2120,N_1935,N_1838);
or U2121 (N_2121,N_1931,N_1881);
xnor U2122 (N_2122,N_1862,N_1964);
xnor U2123 (N_2123,N_1885,N_1994);
xor U2124 (N_2124,N_1820,N_1928);
xnor U2125 (N_2125,N_1886,N_1926);
nand U2126 (N_2126,N_1857,N_1834);
xnor U2127 (N_2127,N_1930,N_1920);
or U2128 (N_2128,N_1860,N_1890);
or U2129 (N_2129,N_1801,N_1887);
and U2130 (N_2130,N_1954,N_1891);
and U2131 (N_2131,N_1816,N_1953);
or U2132 (N_2132,N_1884,N_1970);
nor U2133 (N_2133,N_1920,N_1937);
nand U2134 (N_2134,N_1900,N_1818);
nor U2135 (N_2135,N_1846,N_1969);
and U2136 (N_2136,N_1828,N_1877);
nand U2137 (N_2137,N_1958,N_1881);
xnor U2138 (N_2138,N_1817,N_1819);
nor U2139 (N_2139,N_1974,N_1866);
nor U2140 (N_2140,N_1907,N_1946);
nand U2141 (N_2141,N_1909,N_1807);
nand U2142 (N_2142,N_1956,N_1800);
or U2143 (N_2143,N_1906,N_1867);
or U2144 (N_2144,N_1844,N_1903);
nand U2145 (N_2145,N_1955,N_1829);
or U2146 (N_2146,N_1866,N_1888);
nor U2147 (N_2147,N_1876,N_1941);
xor U2148 (N_2148,N_1893,N_1834);
nor U2149 (N_2149,N_1934,N_1955);
nor U2150 (N_2150,N_1818,N_1800);
or U2151 (N_2151,N_1978,N_1906);
nand U2152 (N_2152,N_1967,N_1947);
nand U2153 (N_2153,N_1889,N_1826);
nand U2154 (N_2154,N_1838,N_1937);
or U2155 (N_2155,N_1955,N_1967);
nand U2156 (N_2156,N_1892,N_1950);
or U2157 (N_2157,N_1826,N_1818);
nand U2158 (N_2158,N_1863,N_1989);
and U2159 (N_2159,N_1859,N_1970);
or U2160 (N_2160,N_1863,N_1883);
or U2161 (N_2161,N_1878,N_1964);
nand U2162 (N_2162,N_1936,N_1904);
nor U2163 (N_2163,N_1897,N_1858);
xor U2164 (N_2164,N_1912,N_1923);
nand U2165 (N_2165,N_1825,N_1981);
nand U2166 (N_2166,N_1801,N_1866);
nor U2167 (N_2167,N_1867,N_1912);
and U2168 (N_2168,N_1890,N_1821);
nor U2169 (N_2169,N_1845,N_1812);
nor U2170 (N_2170,N_1979,N_1949);
nand U2171 (N_2171,N_1914,N_1823);
or U2172 (N_2172,N_1881,N_1828);
or U2173 (N_2173,N_1933,N_1802);
or U2174 (N_2174,N_1802,N_1858);
nor U2175 (N_2175,N_1890,N_1871);
xor U2176 (N_2176,N_1809,N_1982);
xor U2177 (N_2177,N_1920,N_1876);
and U2178 (N_2178,N_1964,N_1971);
and U2179 (N_2179,N_1904,N_1803);
and U2180 (N_2180,N_1885,N_1978);
nor U2181 (N_2181,N_1886,N_1807);
or U2182 (N_2182,N_1880,N_1934);
xnor U2183 (N_2183,N_1879,N_1908);
and U2184 (N_2184,N_1893,N_1945);
or U2185 (N_2185,N_1804,N_1901);
or U2186 (N_2186,N_1984,N_1988);
or U2187 (N_2187,N_1981,N_1837);
nand U2188 (N_2188,N_1920,N_1879);
and U2189 (N_2189,N_1964,N_1987);
nand U2190 (N_2190,N_1978,N_1881);
or U2191 (N_2191,N_1964,N_1996);
nand U2192 (N_2192,N_1981,N_1876);
xnor U2193 (N_2193,N_1913,N_1962);
and U2194 (N_2194,N_1835,N_1994);
nor U2195 (N_2195,N_1950,N_1811);
and U2196 (N_2196,N_1878,N_1903);
and U2197 (N_2197,N_1806,N_1824);
nand U2198 (N_2198,N_1845,N_1808);
or U2199 (N_2199,N_1999,N_1880);
nand U2200 (N_2200,N_2128,N_2034);
xnor U2201 (N_2201,N_2022,N_2132);
nand U2202 (N_2202,N_2171,N_2043);
nand U2203 (N_2203,N_2179,N_2137);
xor U2204 (N_2204,N_2039,N_2008);
and U2205 (N_2205,N_2032,N_2119);
xnor U2206 (N_2206,N_2067,N_2002);
or U2207 (N_2207,N_2154,N_2096);
xnor U2208 (N_2208,N_2004,N_2031);
xnor U2209 (N_2209,N_2059,N_2101);
and U2210 (N_2210,N_2150,N_2057);
xor U2211 (N_2211,N_2056,N_2189);
and U2212 (N_2212,N_2165,N_2055);
or U2213 (N_2213,N_2087,N_2062);
and U2214 (N_2214,N_2076,N_2009);
nand U2215 (N_2215,N_2047,N_2162);
xnor U2216 (N_2216,N_2133,N_2116);
xnor U2217 (N_2217,N_2089,N_2103);
nand U2218 (N_2218,N_2065,N_2038);
xnor U2219 (N_2219,N_2113,N_2129);
and U2220 (N_2220,N_2003,N_2186);
and U2221 (N_2221,N_2066,N_2135);
and U2222 (N_2222,N_2078,N_2172);
or U2223 (N_2223,N_2035,N_2050);
or U2224 (N_2224,N_2177,N_2033);
and U2225 (N_2225,N_2090,N_2158);
or U2226 (N_2226,N_2104,N_2139);
xor U2227 (N_2227,N_2187,N_2130);
nand U2228 (N_2228,N_2016,N_2045);
nor U2229 (N_2229,N_2170,N_2125);
nand U2230 (N_2230,N_2083,N_2126);
xor U2231 (N_2231,N_2120,N_2143);
or U2232 (N_2232,N_2027,N_2086);
xor U2233 (N_2233,N_2106,N_2196);
or U2234 (N_2234,N_2159,N_2114);
xor U2235 (N_2235,N_2163,N_2088);
nor U2236 (N_2236,N_2107,N_2098);
xnor U2237 (N_2237,N_2193,N_2072);
or U2238 (N_2238,N_2079,N_2147);
nor U2239 (N_2239,N_2157,N_2138);
xor U2240 (N_2240,N_2148,N_2173);
nor U2241 (N_2241,N_2053,N_2077);
xnor U2242 (N_2242,N_2028,N_2102);
or U2243 (N_2243,N_2167,N_2197);
and U2244 (N_2244,N_2037,N_2085);
or U2245 (N_2245,N_2042,N_2095);
xnor U2246 (N_2246,N_2166,N_2176);
xor U2247 (N_2247,N_2142,N_2048);
and U2248 (N_2248,N_2069,N_2054);
nor U2249 (N_2249,N_2001,N_2024);
or U2250 (N_2250,N_2044,N_2180);
or U2251 (N_2251,N_2188,N_2017);
xnor U2252 (N_2252,N_2019,N_2000);
nand U2253 (N_2253,N_2012,N_2156);
and U2254 (N_2254,N_2131,N_2015);
or U2255 (N_2255,N_2068,N_2080);
nand U2256 (N_2256,N_2049,N_2190);
and U2257 (N_2257,N_2013,N_2127);
or U2258 (N_2258,N_2109,N_2155);
and U2259 (N_2259,N_2040,N_2018);
nor U2260 (N_2260,N_2005,N_2161);
or U2261 (N_2261,N_2075,N_2023);
nand U2262 (N_2262,N_2123,N_2182);
nor U2263 (N_2263,N_2121,N_2011);
nand U2264 (N_2264,N_2030,N_2152);
and U2265 (N_2265,N_2006,N_2071);
xnor U2266 (N_2266,N_2060,N_2140);
nand U2267 (N_2267,N_2007,N_2052);
nand U2268 (N_2268,N_2169,N_2149);
and U2269 (N_2269,N_2061,N_2191);
nor U2270 (N_2270,N_2036,N_2175);
and U2271 (N_2271,N_2051,N_2097);
xnor U2272 (N_2272,N_2074,N_2153);
and U2273 (N_2273,N_2014,N_2199);
or U2274 (N_2274,N_2070,N_2082);
and U2275 (N_2275,N_2168,N_2124);
or U2276 (N_2276,N_2112,N_2144);
nor U2277 (N_2277,N_2093,N_2164);
and U2278 (N_2278,N_2041,N_2118);
nor U2279 (N_2279,N_2084,N_2185);
or U2280 (N_2280,N_2025,N_2141);
and U2281 (N_2281,N_2099,N_2058);
nor U2282 (N_2282,N_2136,N_2020);
or U2283 (N_2283,N_2108,N_2174);
xnor U2284 (N_2284,N_2100,N_2192);
nor U2285 (N_2285,N_2183,N_2105);
and U2286 (N_2286,N_2184,N_2110);
nand U2287 (N_2287,N_2021,N_2029);
nor U2288 (N_2288,N_2091,N_2081);
or U2289 (N_2289,N_2010,N_2063);
or U2290 (N_2290,N_2198,N_2194);
nand U2291 (N_2291,N_2111,N_2160);
nor U2292 (N_2292,N_2026,N_2145);
nor U2293 (N_2293,N_2115,N_2117);
xor U2294 (N_2294,N_2181,N_2134);
nor U2295 (N_2295,N_2092,N_2064);
and U2296 (N_2296,N_2122,N_2195);
xnor U2297 (N_2297,N_2094,N_2073);
nand U2298 (N_2298,N_2178,N_2046);
and U2299 (N_2299,N_2151,N_2146);
nand U2300 (N_2300,N_2046,N_2160);
nor U2301 (N_2301,N_2198,N_2107);
or U2302 (N_2302,N_2102,N_2114);
or U2303 (N_2303,N_2103,N_2009);
nand U2304 (N_2304,N_2024,N_2199);
or U2305 (N_2305,N_2129,N_2128);
and U2306 (N_2306,N_2105,N_2171);
nand U2307 (N_2307,N_2028,N_2042);
xnor U2308 (N_2308,N_2097,N_2158);
xnor U2309 (N_2309,N_2124,N_2056);
nor U2310 (N_2310,N_2098,N_2010);
nor U2311 (N_2311,N_2000,N_2114);
xnor U2312 (N_2312,N_2108,N_2177);
xnor U2313 (N_2313,N_2135,N_2013);
or U2314 (N_2314,N_2001,N_2076);
nand U2315 (N_2315,N_2190,N_2088);
or U2316 (N_2316,N_2171,N_2050);
or U2317 (N_2317,N_2124,N_2096);
nand U2318 (N_2318,N_2119,N_2004);
nand U2319 (N_2319,N_2046,N_2039);
nor U2320 (N_2320,N_2056,N_2198);
xnor U2321 (N_2321,N_2098,N_2182);
nor U2322 (N_2322,N_2143,N_2150);
and U2323 (N_2323,N_2185,N_2009);
and U2324 (N_2324,N_2046,N_2005);
or U2325 (N_2325,N_2081,N_2153);
xor U2326 (N_2326,N_2121,N_2016);
or U2327 (N_2327,N_2158,N_2050);
nor U2328 (N_2328,N_2129,N_2093);
and U2329 (N_2329,N_2068,N_2188);
nand U2330 (N_2330,N_2094,N_2054);
nand U2331 (N_2331,N_2184,N_2064);
and U2332 (N_2332,N_2092,N_2003);
nand U2333 (N_2333,N_2157,N_2114);
nor U2334 (N_2334,N_2043,N_2100);
nand U2335 (N_2335,N_2104,N_2054);
and U2336 (N_2336,N_2042,N_2049);
or U2337 (N_2337,N_2047,N_2036);
nor U2338 (N_2338,N_2099,N_2029);
and U2339 (N_2339,N_2033,N_2024);
nand U2340 (N_2340,N_2141,N_2050);
nand U2341 (N_2341,N_2096,N_2002);
nand U2342 (N_2342,N_2115,N_2179);
nand U2343 (N_2343,N_2014,N_2194);
and U2344 (N_2344,N_2190,N_2110);
xor U2345 (N_2345,N_2057,N_2013);
nand U2346 (N_2346,N_2100,N_2135);
or U2347 (N_2347,N_2005,N_2179);
xor U2348 (N_2348,N_2005,N_2145);
nand U2349 (N_2349,N_2032,N_2106);
or U2350 (N_2350,N_2024,N_2079);
xor U2351 (N_2351,N_2016,N_2098);
xnor U2352 (N_2352,N_2125,N_2057);
nand U2353 (N_2353,N_2147,N_2178);
nor U2354 (N_2354,N_2191,N_2065);
or U2355 (N_2355,N_2156,N_2137);
and U2356 (N_2356,N_2127,N_2115);
nand U2357 (N_2357,N_2085,N_2137);
or U2358 (N_2358,N_2121,N_2155);
xor U2359 (N_2359,N_2162,N_2095);
xnor U2360 (N_2360,N_2158,N_2004);
or U2361 (N_2361,N_2100,N_2179);
or U2362 (N_2362,N_2140,N_2009);
and U2363 (N_2363,N_2167,N_2041);
nor U2364 (N_2364,N_2133,N_2120);
xnor U2365 (N_2365,N_2169,N_2144);
or U2366 (N_2366,N_2165,N_2109);
or U2367 (N_2367,N_2183,N_2004);
nor U2368 (N_2368,N_2038,N_2150);
nand U2369 (N_2369,N_2009,N_2125);
nor U2370 (N_2370,N_2190,N_2051);
xnor U2371 (N_2371,N_2046,N_2069);
or U2372 (N_2372,N_2193,N_2096);
nand U2373 (N_2373,N_2167,N_2194);
xnor U2374 (N_2374,N_2099,N_2163);
and U2375 (N_2375,N_2059,N_2098);
and U2376 (N_2376,N_2117,N_2062);
xor U2377 (N_2377,N_2052,N_2146);
or U2378 (N_2378,N_2021,N_2071);
nor U2379 (N_2379,N_2103,N_2110);
and U2380 (N_2380,N_2016,N_2001);
xnor U2381 (N_2381,N_2047,N_2015);
and U2382 (N_2382,N_2116,N_2128);
or U2383 (N_2383,N_2139,N_2012);
xor U2384 (N_2384,N_2118,N_2138);
nor U2385 (N_2385,N_2050,N_2162);
or U2386 (N_2386,N_2011,N_2108);
or U2387 (N_2387,N_2182,N_2008);
xor U2388 (N_2388,N_2189,N_2038);
or U2389 (N_2389,N_2041,N_2003);
xor U2390 (N_2390,N_2091,N_2153);
xnor U2391 (N_2391,N_2125,N_2027);
or U2392 (N_2392,N_2060,N_2152);
and U2393 (N_2393,N_2134,N_2033);
or U2394 (N_2394,N_2044,N_2050);
xor U2395 (N_2395,N_2094,N_2172);
nor U2396 (N_2396,N_2191,N_2062);
or U2397 (N_2397,N_2150,N_2181);
nand U2398 (N_2398,N_2089,N_2191);
or U2399 (N_2399,N_2081,N_2127);
nor U2400 (N_2400,N_2211,N_2264);
nand U2401 (N_2401,N_2352,N_2320);
nand U2402 (N_2402,N_2330,N_2285);
xnor U2403 (N_2403,N_2221,N_2299);
or U2404 (N_2404,N_2344,N_2387);
and U2405 (N_2405,N_2274,N_2391);
or U2406 (N_2406,N_2289,N_2226);
xnor U2407 (N_2407,N_2380,N_2362);
nand U2408 (N_2408,N_2331,N_2373);
nor U2409 (N_2409,N_2227,N_2287);
xor U2410 (N_2410,N_2388,N_2245);
or U2411 (N_2411,N_2209,N_2201);
nor U2412 (N_2412,N_2292,N_2350);
nor U2413 (N_2413,N_2389,N_2302);
nand U2414 (N_2414,N_2228,N_2343);
and U2415 (N_2415,N_2220,N_2323);
and U2416 (N_2416,N_2296,N_2318);
xor U2417 (N_2417,N_2239,N_2273);
or U2418 (N_2418,N_2231,N_2284);
nand U2419 (N_2419,N_2277,N_2392);
and U2420 (N_2420,N_2250,N_2263);
nor U2421 (N_2421,N_2313,N_2314);
and U2422 (N_2422,N_2203,N_2370);
nand U2423 (N_2423,N_2234,N_2257);
xnor U2424 (N_2424,N_2253,N_2233);
xor U2425 (N_2425,N_2351,N_2293);
nand U2426 (N_2426,N_2272,N_2241);
nor U2427 (N_2427,N_2256,N_2254);
nor U2428 (N_2428,N_2333,N_2283);
and U2429 (N_2429,N_2358,N_2282);
and U2430 (N_2430,N_2294,N_2360);
and U2431 (N_2431,N_2248,N_2204);
xnor U2432 (N_2432,N_2208,N_2332);
xor U2433 (N_2433,N_2255,N_2329);
and U2434 (N_2434,N_2281,N_2288);
and U2435 (N_2435,N_2308,N_2345);
xor U2436 (N_2436,N_2307,N_2390);
nor U2437 (N_2437,N_2202,N_2353);
nand U2438 (N_2438,N_2355,N_2368);
or U2439 (N_2439,N_2230,N_2361);
nand U2440 (N_2440,N_2270,N_2342);
nor U2441 (N_2441,N_2216,N_2275);
nand U2442 (N_2442,N_2229,N_2261);
xnor U2443 (N_2443,N_2300,N_2372);
nor U2444 (N_2444,N_2214,N_2371);
xor U2445 (N_2445,N_2269,N_2346);
nand U2446 (N_2446,N_2246,N_2398);
and U2447 (N_2447,N_2347,N_2240);
nand U2448 (N_2448,N_2365,N_2235);
and U2449 (N_2449,N_2315,N_2232);
nand U2450 (N_2450,N_2243,N_2238);
or U2451 (N_2451,N_2396,N_2359);
nand U2452 (N_2452,N_2339,N_2316);
or U2453 (N_2453,N_2236,N_2317);
and U2454 (N_2454,N_2306,N_2291);
nand U2455 (N_2455,N_2278,N_2384);
nand U2456 (N_2456,N_2335,N_2286);
and U2457 (N_2457,N_2354,N_2206);
nand U2458 (N_2458,N_2311,N_2376);
xnor U2459 (N_2459,N_2337,N_2295);
nand U2460 (N_2460,N_2377,N_2399);
and U2461 (N_2461,N_2212,N_2378);
nor U2462 (N_2462,N_2374,N_2309);
and U2463 (N_2463,N_2383,N_2259);
and U2464 (N_2464,N_2340,N_2215);
nand U2465 (N_2465,N_2262,N_2369);
nor U2466 (N_2466,N_2324,N_2382);
and U2467 (N_2467,N_2297,N_2322);
or U2468 (N_2468,N_2310,N_2224);
nand U2469 (N_2469,N_2207,N_2260);
and U2470 (N_2470,N_2321,N_2381);
xor U2471 (N_2471,N_2375,N_2213);
or U2472 (N_2472,N_2304,N_2356);
and U2473 (N_2473,N_2258,N_2319);
and U2474 (N_2474,N_2363,N_2348);
xor U2475 (N_2475,N_2366,N_2217);
or U2476 (N_2476,N_2237,N_2325);
nor U2477 (N_2477,N_2271,N_2397);
and U2478 (N_2478,N_2312,N_2268);
xor U2479 (N_2479,N_2303,N_2225);
or U2480 (N_2480,N_2298,N_2338);
xor U2481 (N_2481,N_2249,N_2219);
and U2482 (N_2482,N_2210,N_2267);
nor U2483 (N_2483,N_2247,N_2385);
xor U2484 (N_2484,N_2327,N_2251);
xnor U2485 (N_2485,N_2290,N_2364);
and U2486 (N_2486,N_2357,N_2280);
xor U2487 (N_2487,N_2266,N_2386);
and U2488 (N_2488,N_2223,N_2200);
xor U2489 (N_2489,N_2244,N_2305);
or U2490 (N_2490,N_2205,N_2222);
nand U2491 (N_2491,N_2279,N_2328);
and U2492 (N_2492,N_2395,N_2393);
and U2493 (N_2493,N_2301,N_2326);
or U2494 (N_2494,N_2218,N_2252);
or U2495 (N_2495,N_2336,N_2379);
and U2496 (N_2496,N_2242,N_2341);
nor U2497 (N_2497,N_2276,N_2394);
or U2498 (N_2498,N_2367,N_2349);
nor U2499 (N_2499,N_2334,N_2265);
or U2500 (N_2500,N_2307,N_2240);
nor U2501 (N_2501,N_2318,N_2205);
and U2502 (N_2502,N_2210,N_2242);
and U2503 (N_2503,N_2289,N_2251);
or U2504 (N_2504,N_2263,N_2349);
xor U2505 (N_2505,N_2339,N_2370);
or U2506 (N_2506,N_2270,N_2227);
nand U2507 (N_2507,N_2228,N_2267);
and U2508 (N_2508,N_2368,N_2261);
nor U2509 (N_2509,N_2252,N_2297);
nor U2510 (N_2510,N_2290,N_2385);
or U2511 (N_2511,N_2399,N_2272);
xnor U2512 (N_2512,N_2327,N_2370);
xnor U2513 (N_2513,N_2357,N_2396);
nor U2514 (N_2514,N_2345,N_2385);
and U2515 (N_2515,N_2225,N_2240);
and U2516 (N_2516,N_2390,N_2230);
or U2517 (N_2517,N_2308,N_2201);
nand U2518 (N_2518,N_2284,N_2384);
nand U2519 (N_2519,N_2231,N_2383);
xor U2520 (N_2520,N_2217,N_2358);
nand U2521 (N_2521,N_2319,N_2279);
xor U2522 (N_2522,N_2369,N_2388);
or U2523 (N_2523,N_2332,N_2256);
or U2524 (N_2524,N_2248,N_2334);
nand U2525 (N_2525,N_2234,N_2370);
xnor U2526 (N_2526,N_2352,N_2313);
nor U2527 (N_2527,N_2293,N_2256);
xor U2528 (N_2528,N_2392,N_2292);
nor U2529 (N_2529,N_2217,N_2377);
or U2530 (N_2530,N_2391,N_2279);
xor U2531 (N_2531,N_2229,N_2266);
and U2532 (N_2532,N_2220,N_2239);
and U2533 (N_2533,N_2380,N_2210);
and U2534 (N_2534,N_2362,N_2315);
xor U2535 (N_2535,N_2349,N_2260);
and U2536 (N_2536,N_2258,N_2379);
xnor U2537 (N_2537,N_2389,N_2255);
or U2538 (N_2538,N_2383,N_2299);
or U2539 (N_2539,N_2324,N_2384);
xnor U2540 (N_2540,N_2396,N_2316);
nand U2541 (N_2541,N_2349,N_2220);
or U2542 (N_2542,N_2207,N_2358);
or U2543 (N_2543,N_2368,N_2379);
nor U2544 (N_2544,N_2382,N_2360);
or U2545 (N_2545,N_2256,N_2201);
nor U2546 (N_2546,N_2220,N_2300);
nand U2547 (N_2547,N_2246,N_2395);
nand U2548 (N_2548,N_2317,N_2376);
and U2549 (N_2549,N_2342,N_2239);
nor U2550 (N_2550,N_2396,N_2321);
xnor U2551 (N_2551,N_2347,N_2251);
or U2552 (N_2552,N_2394,N_2293);
xor U2553 (N_2553,N_2376,N_2290);
nor U2554 (N_2554,N_2234,N_2224);
nand U2555 (N_2555,N_2214,N_2262);
nand U2556 (N_2556,N_2352,N_2384);
nor U2557 (N_2557,N_2313,N_2336);
nor U2558 (N_2558,N_2205,N_2244);
or U2559 (N_2559,N_2292,N_2326);
nor U2560 (N_2560,N_2325,N_2303);
nand U2561 (N_2561,N_2396,N_2257);
xnor U2562 (N_2562,N_2233,N_2346);
nor U2563 (N_2563,N_2381,N_2224);
xnor U2564 (N_2564,N_2373,N_2352);
xor U2565 (N_2565,N_2322,N_2357);
or U2566 (N_2566,N_2305,N_2269);
xor U2567 (N_2567,N_2262,N_2380);
or U2568 (N_2568,N_2268,N_2290);
nor U2569 (N_2569,N_2343,N_2398);
and U2570 (N_2570,N_2382,N_2288);
nor U2571 (N_2571,N_2254,N_2337);
and U2572 (N_2572,N_2300,N_2344);
nand U2573 (N_2573,N_2227,N_2291);
or U2574 (N_2574,N_2233,N_2283);
or U2575 (N_2575,N_2388,N_2249);
xnor U2576 (N_2576,N_2208,N_2377);
xnor U2577 (N_2577,N_2285,N_2331);
and U2578 (N_2578,N_2398,N_2272);
nand U2579 (N_2579,N_2319,N_2281);
nor U2580 (N_2580,N_2337,N_2285);
or U2581 (N_2581,N_2290,N_2277);
nor U2582 (N_2582,N_2353,N_2345);
and U2583 (N_2583,N_2325,N_2205);
xor U2584 (N_2584,N_2228,N_2239);
nor U2585 (N_2585,N_2390,N_2243);
nand U2586 (N_2586,N_2352,N_2284);
or U2587 (N_2587,N_2350,N_2358);
nor U2588 (N_2588,N_2309,N_2366);
or U2589 (N_2589,N_2386,N_2323);
xnor U2590 (N_2590,N_2279,N_2298);
or U2591 (N_2591,N_2318,N_2212);
xor U2592 (N_2592,N_2260,N_2325);
xnor U2593 (N_2593,N_2244,N_2372);
and U2594 (N_2594,N_2293,N_2289);
nor U2595 (N_2595,N_2388,N_2332);
and U2596 (N_2596,N_2329,N_2332);
nand U2597 (N_2597,N_2255,N_2335);
or U2598 (N_2598,N_2222,N_2204);
xor U2599 (N_2599,N_2390,N_2241);
xor U2600 (N_2600,N_2459,N_2594);
xor U2601 (N_2601,N_2525,N_2495);
xor U2602 (N_2602,N_2563,N_2585);
nor U2603 (N_2603,N_2415,N_2554);
or U2604 (N_2604,N_2434,N_2456);
xor U2605 (N_2605,N_2538,N_2552);
nand U2606 (N_2606,N_2413,N_2595);
and U2607 (N_2607,N_2590,N_2444);
nand U2608 (N_2608,N_2429,N_2584);
or U2609 (N_2609,N_2457,N_2482);
and U2610 (N_2610,N_2542,N_2446);
and U2611 (N_2611,N_2576,N_2416);
and U2612 (N_2612,N_2517,N_2515);
and U2613 (N_2613,N_2518,N_2427);
nand U2614 (N_2614,N_2534,N_2509);
nor U2615 (N_2615,N_2561,N_2469);
or U2616 (N_2616,N_2508,N_2420);
nor U2617 (N_2617,N_2581,N_2514);
or U2618 (N_2618,N_2436,N_2587);
and U2619 (N_2619,N_2502,N_2583);
nor U2620 (N_2620,N_2569,N_2491);
and U2621 (N_2621,N_2474,N_2507);
nand U2622 (N_2622,N_2567,N_2463);
or U2623 (N_2623,N_2564,N_2573);
and U2624 (N_2624,N_2405,N_2497);
xor U2625 (N_2625,N_2533,N_2532);
xor U2626 (N_2626,N_2557,N_2521);
nor U2627 (N_2627,N_2451,N_2575);
or U2628 (N_2628,N_2430,N_2522);
and U2629 (N_2629,N_2402,N_2473);
and U2630 (N_2630,N_2544,N_2545);
xor U2631 (N_2631,N_2513,N_2425);
nand U2632 (N_2632,N_2598,N_2528);
xor U2633 (N_2633,N_2455,N_2407);
nand U2634 (N_2634,N_2401,N_2445);
and U2635 (N_2635,N_2588,N_2454);
nor U2636 (N_2636,N_2537,N_2437);
nand U2637 (N_2637,N_2577,N_2486);
xnor U2638 (N_2638,N_2526,N_2597);
nand U2639 (N_2639,N_2535,N_2559);
or U2640 (N_2640,N_2406,N_2494);
nor U2641 (N_2641,N_2417,N_2505);
xor U2642 (N_2642,N_2452,N_2571);
or U2643 (N_2643,N_2589,N_2530);
nand U2644 (N_2644,N_2510,N_2547);
xor U2645 (N_2645,N_2476,N_2540);
nor U2646 (N_2646,N_2411,N_2499);
and U2647 (N_2647,N_2422,N_2516);
and U2648 (N_2648,N_2488,N_2492);
nand U2649 (N_2649,N_2479,N_2580);
xnor U2650 (N_2650,N_2501,N_2558);
or U2651 (N_2651,N_2438,N_2419);
or U2652 (N_2652,N_2440,N_2527);
and U2653 (N_2653,N_2593,N_2496);
and U2654 (N_2654,N_2565,N_2431);
nand U2655 (N_2655,N_2433,N_2471);
nor U2656 (N_2656,N_2465,N_2578);
or U2657 (N_2657,N_2566,N_2464);
nor U2658 (N_2658,N_2443,N_2477);
xor U2659 (N_2659,N_2448,N_2560);
or U2660 (N_2660,N_2493,N_2484);
nor U2661 (N_2661,N_2490,N_2550);
nor U2662 (N_2662,N_2582,N_2453);
nor U2663 (N_2663,N_2531,N_2400);
nor U2664 (N_2664,N_2414,N_2441);
or U2665 (N_2665,N_2487,N_2572);
nor U2666 (N_2666,N_2418,N_2475);
nand U2667 (N_2667,N_2504,N_2553);
or U2668 (N_2668,N_2480,N_2520);
xor U2669 (N_2669,N_2555,N_2403);
nor U2670 (N_2670,N_2548,N_2461);
xor U2671 (N_2671,N_2541,N_2543);
or U2672 (N_2672,N_2570,N_2460);
xnor U2673 (N_2673,N_2579,N_2549);
nand U2674 (N_2674,N_2519,N_2483);
or U2675 (N_2675,N_2592,N_2599);
xor U2676 (N_2676,N_2466,N_2503);
nand U2677 (N_2677,N_2439,N_2426);
nor U2678 (N_2678,N_2485,N_2404);
nand U2679 (N_2679,N_2539,N_2506);
xnor U2680 (N_2680,N_2586,N_2546);
or U2681 (N_2681,N_2432,N_2449);
nand U2682 (N_2682,N_2447,N_2489);
and U2683 (N_2683,N_2408,N_2450);
nor U2684 (N_2684,N_2511,N_2468);
xnor U2685 (N_2685,N_2512,N_2481);
and U2686 (N_2686,N_2467,N_2524);
nand U2687 (N_2687,N_2462,N_2428);
nor U2688 (N_2688,N_2568,N_2591);
xor U2689 (N_2689,N_2412,N_2556);
nor U2690 (N_2690,N_2596,N_2562);
and U2691 (N_2691,N_2423,N_2472);
nor U2692 (N_2692,N_2523,N_2409);
nand U2693 (N_2693,N_2421,N_2458);
xor U2694 (N_2694,N_2500,N_2574);
or U2695 (N_2695,N_2410,N_2498);
nand U2696 (N_2696,N_2536,N_2442);
or U2697 (N_2697,N_2529,N_2551);
or U2698 (N_2698,N_2435,N_2470);
or U2699 (N_2699,N_2424,N_2478);
nor U2700 (N_2700,N_2582,N_2534);
nor U2701 (N_2701,N_2483,N_2523);
nand U2702 (N_2702,N_2540,N_2539);
and U2703 (N_2703,N_2401,N_2558);
and U2704 (N_2704,N_2414,N_2537);
or U2705 (N_2705,N_2575,N_2505);
xor U2706 (N_2706,N_2591,N_2463);
xnor U2707 (N_2707,N_2492,N_2446);
xnor U2708 (N_2708,N_2575,N_2588);
nand U2709 (N_2709,N_2470,N_2444);
nor U2710 (N_2710,N_2557,N_2580);
xnor U2711 (N_2711,N_2509,N_2579);
nor U2712 (N_2712,N_2468,N_2447);
nand U2713 (N_2713,N_2527,N_2530);
nand U2714 (N_2714,N_2513,N_2437);
and U2715 (N_2715,N_2501,N_2408);
or U2716 (N_2716,N_2586,N_2486);
xnor U2717 (N_2717,N_2585,N_2430);
xnor U2718 (N_2718,N_2537,N_2448);
or U2719 (N_2719,N_2485,N_2480);
nand U2720 (N_2720,N_2502,N_2410);
nor U2721 (N_2721,N_2421,N_2450);
nor U2722 (N_2722,N_2530,N_2509);
and U2723 (N_2723,N_2535,N_2554);
and U2724 (N_2724,N_2425,N_2567);
nand U2725 (N_2725,N_2587,N_2544);
nand U2726 (N_2726,N_2491,N_2526);
or U2727 (N_2727,N_2482,N_2453);
or U2728 (N_2728,N_2548,N_2469);
or U2729 (N_2729,N_2522,N_2448);
nand U2730 (N_2730,N_2511,N_2529);
xnor U2731 (N_2731,N_2479,N_2548);
xnor U2732 (N_2732,N_2514,N_2526);
xor U2733 (N_2733,N_2576,N_2571);
nor U2734 (N_2734,N_2409,N_2558);
or U2735 (N_2735,N_2571,N_2437);
or U2736 (N_2736,N_2470,N_2446);
xnor U2737 (N_2737,N_2568,N_2430);
or U2738 (N_2738,N_2583,N_2489);
nor U2739 (N_2739,N_2592,N_2441);
xnor U2740 (N_2740,N_2432,N_2544);
xor U2741 (N_2741,N_2594,N_2545);
and U2742 (N_2742,N_2499,N_2568);
or U2743 (N_2743,N_2508,N_2576);
xnor U2744 (N_2744,N_2468,N_2491);
nor U2745 (N_2745,N_2507,N_2466);
or U2746 (N_2746,N_2550,N_2443);
nor U2747 (N_2747,N_2511,N_2483);
nor U2748 (N_2748,N_2565,N_2534);
or U2749 (N_2749,N_2574,N_2407);
or U2750 (N_2750,N_2580,N_2418);
or U2751 (N_2751,N_2520,N_2479);
nor U2752 (N_2752,N_2576,N_2456);
nor U2753 (N_2753,N_2523,N_2554);
nand U2754 (N_2754,N_2452,N_2474);
xnor U2755 (N_2755,N_2533,N_2541);
or U2756 (N_2756,N_2522,N_2586);
nand U2757 (N_2757,N_2559,N_2563);
or U2758 (N_2758,N_2476,N_2503);
xnor U2759 (N_2759,N_2581,N_2423);
xor U2760 (N_2760,N_2489,N_2411);
or U2761 (N_2761,N_2595,N_2562);
or U2762 (N_2762,N_2584,N_2453);
or U2763 (N_2763,N_2504,N_2581);
or U2764 (N_2764,N_2442,N_2551);
or U2765 (N_2765,N_2594,N_2489);
xnor U2766 (N_2766,N_2553,N_2471);
nor U2767 (N_2767,N_2483,N_2431);
or U2768 (N_2768,N_2449,N_2423);
or U2769 (N_2769,N_2596,N_2523);
and U2770 (N_2770,N_2448,N_2585);
xnor U2771 (N_2771,N_2497,N_2520);
and U2772 (N_2772,N_2586,N_2514);
or U2773 (N_2773,N_2583,N_2422);
nand U2774 (N_2774,N_2413,N_2577);
nor U2775 (N_2775,N_2565,N_2542);
and U2776 (N_2776,N_2419,N_2404);
and U2777 (N_2777,N_2557,N_2550);
or U2778 (N_2778,N_2543,N_2431);
nor U2779 (N_2779,N_2540,N_2458);
or U2780 (N_2780,N_2414,N_2543);
nor U2781 (N_2781,N_2591,N_2562);
or U2782 (N_2782,N_2527,N_2543);
and U2783 (N_2783,N_2560,N_2594);
nand U2784 (N_2784,N_2415,N_2476);
nand U2785 (N_2785,N_2538,N_2558);
or U2786 (N_2786,N_2411,N_2564);
xnor U2787 (N_2787,N_2428,N_2549);
nor U2788 (N_2788,N_2523,N_2577);
or U2789 (N_2789,N_2411,N_2555);
or U2790 (N_2790,N_2452,N_2483);
nor U2791 (N_2791,N_2461,N_2512);
or U2792 (N_2792,N_2455,N_2420);
nor U2793 (N_2793,N_2593,N_2590);
and U2794 (N_2794,N_2480,N_2400);
or U2795 (N_2795,N_2423,N_2468);
xnor U2796 (N_2796,N_2461,N_2550);
or U2797 (N_2797,N_2471,N_2509);
xnor U2798 (N_2798,N_2534,N_2414);
nor U2799 (N_2799,N_2492,N_2453);
xnor U2800 (N_2800,N_2690,N_2642);
or U2801 (N_2801,N_2683,N_2738);
nand U2802 (N_2802,N_2749,N_2723);
or U2803 (N_2803,N_2762,N_2793);
or U2804 (N_2804,N_2724,N_2663);
nor U2805 (N_2805,N_2713,N_2750);
and U2806 (N_2806,N_2633,N_2615);
or U2807 (N_2807,N_2791,N_2774);
or U2808 (N_2808,N_2781,N_2797);
and U2809 (N_2809,N_2602,N_2635);
nor U2810 (N_2810,N_2717,N_2659);
nor U2811 (N_2811,N_2621,N_2681);
xnor U2812 (N_2812,N_2655,N_2608);
or U2813 (N_2813,N_2623,N_2657);
xor U2814 (N_2814,N_2634,N_2771);
nor U2815 (N_2815,N_2695,N_2616);
nand U2816 (N_2816,N_2780,N_2798);
nand U2817 (N_2817,N_2753,N_2672);
and U2818 (N_2818,N_2628,N_2688);
and U2819 (N_2819,N_2669,N_2651);
nand U2820 (N_2820,N_2760,N_2700);
nand U2821 (N_2821,N_2676,N_2662);
or U2822 (N_2822,N_2728,N_2694);
nor U2823 (N_2823,N_2743,N_2629);
or U2824 (N_2824,N_2632,N_2747);
and U2825 (N_2825,N_2716,N_2752);
nor U2826 (N_2826,N_2773,N_2693);
and U2827 (N_2827,N_2714,N_2712);
xor U2828 (N_2828,N_2636,N_2610);
nand U2829 (N_2829,N_2618,N_2645);
xnor U2830 (N_2830,N_2718,N_2758);
or U2831 (N_2831,N_2653,N_2765);
nor U2832 (N_2832,N_2675,N_2764);
or U2833 (N_2833,N_2666,N_2748);
nand U2834 (N_2834,N_2609,N_2604);
and U2835 (N_2835,N_2667,N_2607);
and U2836 (N_2836,N_2674,N_2641);
nor U2837 (N_2837,N_2637,N_2689);
nand U2838 (N_2838,N_2703,N_2761);
nand U2839 (N_2839,N_2739,N_2770);
and U2840 (N_2840,N_2705,N_2744);
or U2841 (N_2841,N_2656,N_2601);
nor U2842 (N_2842,N_2660,N_2727);
xnor U2843 (N_2843,N_2782,N_2706);
or U2844 (N_2844,N_2730,N_2631);
and U2845 (N_2845,N_2790,N_2720);
xor U2846 (N_2846,N_2763,N_2686);
or U2847 (N_2847,N_2769,N_2684);
xnor U2848 (N_2848,N_2707,N_2670);
nor U2849 (N_2849,N_2643,N_2699);
nand U2850 (N_2850,N_2777,N_2679);
nand U2851 (N_2851,N_2691,N_2671);
nor U2852 (N_2852,N_2792,N_2711);
or U2853 (N_2853,N_2756,N_2673);
nand U2854 (N_2854,N_2665,N_2725);
nand U2855 (N_2855,N_2624,N_2605);
nor U2856 (N_2856,N_2622,N_2617);
xnor U2857 (N_2857,N_2726,N_2736);
nor U2858 (N_2858,N_2649,N_2625);
nand U2859 (N_2859,N_2692,N_2784);
nor U2860 (N_2860,N_2772,N_2620);
nor U2861 (N_2861,N_2611,N_2654);
and U2862 (N_2862,N_2627,N_2680);
or U2863 (N_2863,N_2799,N_2788);
nand U2864 (N_2864,N_2708,N_2619);
xor U2865 (N_2865,N_2600,N_2751);
nor U2866 (N_2866,N_2742,N_2704);
or U2867 (N_2867,N_2786,N_2735);
xnor U2868 (N_2868,N_2734,N_2687);
and U2869 (N_2869,N_2664,N_2644);
xor U2870 (N_2870,N_2768,N_2729);
xnor U2871 (N_2871,N_2698,N_2722);
or U2872 (N_2872,N_2766,N_2740);
and U2873 (N_2873,N_2759,N_2648);
nor U2874 (N_2874,N_2775,N_2741);
nor U2875 (N_2875,N_2685,N_2658);
xnor U2876 (N_2876,N_2613,N_2603);
and U2877 (N_2877,N_2626,N_2721);
nor U2878 (N_2878,N_2757,N_2640);
nor U2879 (N_2879,N_2606,N_2755);
xor U2880 (N_2880,N_2639,N_2682);
xnor U2881 (N_2881,N_2646,N_2787);
nand U2882 (N_2882,N_2612,N_2731);
nand U2883 (N_2883,N_2754,N_2677);
nand U2884 (N_2884,N_2737,N_2767);
nor U2885 (N_2885,N_2795,N_2785);
xor U2886 (N_2886,N_2745,N_2702);
nor U2887 (N_2887,N_2668,N_2696);
nor U2888 (N_2888,N_2647,N_2794);
nand U2889 (N_2889,N_2638,N_2701);
or U2890 (N_2890,N_2661,N_2710);
and U2891 (N_2891,N_2697,N_2709);
nand U2892 (N_2892,N_2678,N_2796);
nor U2893 (N_2893,N_2776,N_2746);
nand U2894 (N_2894,N_2778,N_2732);
nand U2895 (N_2895,N_2779,N_2719);
and U2896 (N_2896,N_2652,N_2614);
and U2897 (N_2897,N_2789,N_2733);
xor U2898 (N_2898,N_2630,N_2783);
xor U2899 (N_2899,N_2715,N_2650);
and U2900 (N_2900,N_2770,N_2611);
and U2901 (N_2901,N_2649,N_2772);
and U2902 (N_2902,N_2718,N_2771);
nor U2903 (N_2903,N_2635,N_2642);
or U2904 (N_2904,N_2645,N_2730);
nor U2905 (N_2905,N_2633,N_2767);
or U2906 (N_2906,N_2697,N_2636);
or U2907 (N_2907,N_2736,N_2670);
xor U2908 (N_2908,N_2668,N_2768);
or U2909 (N_2909,N_2766,N_2775);
xor U2910 (N_2910,N_2718,N_2723);
xnor U2911 (N_2911,N_2635,N_2627);
xor U2912 (N_2912,N_2761,N_2622);
and U2913 (N_2913,N_2700,N_2732);
or U2914 (N_2914,N_2699,N_2637);
nand U2915 (N_2915,N_2739,N_2654);
nand U2916 (N_2916,N_2690,N_2681);
nand U2917 (N_2917,N_2776,N_2759);
xnor U2918 (N_2918,N_2740,N_2783);
xor U2919 (N_2919,N_2628,N_2603);
xor U2920 (N_2920,N_2603,N_2605);
nand U2921 (N_2921,N_2624,N_2632);
and U2922 (N_2922,N_2633,N_2751);
nand U2923 (N_2923,N_2668,N_2665);
nand U2924 (N_2924,N_2709,N_2626);
nand U2925 (N_2925,N_2671,N_2776);
xor U2926 (N_2926,N_2755,N_2671);
nand U2927 (N_2927,N_2625,N_2615);
and U2928 (N_2928,N_2626,N_2719);
nor U2929 (N_2929,N_2711,N_2677);
and U2930 (N_2930,N_2796,N_2652);
and U2931 (N_2931,N_2602,N_2722);
xor U2932 (N_2932,N_2710,N_2708);
or U2933 (N_2933,N_2758,N_2748);
xnor U2934 (N_2934,N_2715,N_2603);
xor U2935 (N_2935,N_2796,N_2629);
or U2936 (N_2936,N_2604,N_2777);
nand U2937 (N_2937,N_2718,N_2712);
or U2938 (N_2938,N_2777,N_2618);
or U2939 (N_2939,N_2760,N_2612);
nand U2940 (N_2940,N_2701,N_2722);
nor U2941 (N_2941,N_2748,N_2709);
and U2942 (N_2942,N_2782,N_2759);
nand U2943 (N_2943,N_2626,N_2614);
xor U2944 (N_2944,N_2623,N_2632);
nor U2945 (N_2945,N_2775,N_2787);
and U2946 (N_2946,N_2685,N_2636);
xor U2947 (N_2947,N_2662,N_2683);
and U2948 (N_2948,N_2755,N_2787);
or U2949 (N_2949,N_2756,N_2615);
or U2950 (N_2950,N_2635,N_2658);
or U2951 (N_2951,N_2684,N_2612);
nor U2952 (N_2952,N_2705,N_2781);
nand U2953 (N_2953,N_2766,N_2687);
and U2954 (N_2954,N_2686,N_2621);
xnor U2955 (N_2955,N_2634,N_2707);
or U2956 (N_2956,N_2700,N_2715);
xor U2957 (N_2957,N_2661,N_2608);
xor U2958 (N_2958,N_2612,N_2699);
and U2959 (N_2959,N_2685,N_2611);
and U2960 (N_2960,N_2614,N_2682);
and U2961 (N_2961,N_2698,N_2709);
nand U2962 (N_2962,N_2722,N_2650);
or U2963 (N_2963,N_2671,N_2737);
or U2964 (N_2964,N_2620,N_2733);
and U2965 (N_2965,N_2611,N_2774);
nor U2966 (N_2966,N_2731,N_2771);
nand U2967 (N_2967,N_2671,N_2622);
and U2968 (N_2968,N_2634,N_2712);
nand U2969 (N_2969,N_2688,N_2670);
nor U2970 (N_2970,N_2675,N_2727);
and U2971 (N_2971,N_2711,N_2704);
nor U2972 (N_2972,N_2611,N_2637);
or U2973 (N_2973,N_2765,N_2741);
xnor U2974 (N_2974,N_2775,N_2677);
or U2975 (N_2975,N_2675,N_2661);
nor U2976 (N_2976,N_2740,N_2669);
or U2977 (N_2977,N_2605,N_2781);
nand U2978 (N_2978,N_2695,N_2684);
xnor U2979 (N_2979,N_2796,N_2634);
and U2980 (N_2980,N_2683,N_2753);
xor U2981 (N_2981,N_2610,N_2685);
nand U2982 (N_2982,N_2668,N_2681);
nor U2983 (N_2983,N_2724,N_2703);
nand U2984 (N_2984,N_2765,N_2701);
and U2985 (N_2985,N_2624,N_2692);
xor U2986 (N_2986,N_2760,N_2652);
xor U2987 (N_2987,N_2650,N_2718);
nor U2988 (N_2988,N_2709,N_2696);
xor U2989 (N_2989,N_2758,N_2720);
and U2990 (N_2990,N_2612,N_2630);
nor U2991 (N_2991,N_2710,N_2792);
nor U2992 (N_2992,N_2633,N_2653);
nor U2993 (N_2993,N_2667,N_2767);
or U2994 (N_2994,N_2670,N_2789);
nand U2995 (N_2995,N_2789,N_2672);
nor U2996 (N_2996,N_2672,N_2725);
xnor U2997 (N_2997,N_2673,N_2759);
nand U2998 (N_2998,N_2616,N_2691);
and U2999 (N_2999,N_2773,N_2670);
xnor U3000 (N_3000,N_2869,N_2901);
nor U3001 (N_3001,N_2964,N_2904);
and U3002 (N_3002,N_2882,N_2899);
and U3003 (N_3003,N_2974,N_2932);
nor U3004 (N_3004,N_2816,N_2886);
or U3005 (N_3005,N_2983,N_2988);
or U3006 (N_3006,N_2812,N_2960);
and U3007 (N_3007,N_2979,N_2860);
nand U3008 (N_3008,N_2863,N_2864);
nand U3009 (N_3009,N_2876,N_2908);
nor U3010 (N_3010,N_2889,N_2857);
xnor U3011 (N_3011,N_2871,N_2937);
xor U3012 (N_3012,N_2985,N_2829);
nor U3013 (N_3013,N_2827,N_2859);
xor U3014 (N_3014,N_2912,N_2892);
or U3015 (N_3015,N_2825,N_2893);
and U3016 (N_3016,N_2910,N_2994);
nand U3017 (N_3017,N_2890,N_2822);
and U3018 (N_3018,N_2956,N_2887);
nor U3019 (N_3019,N_2836,N_2920);
xnor U3020 (N_3020,N_2973,N_2903);
and U3021 (N_3021,N_2962,N_2971);
nand U3022 (N_3022,N_2996,N_2954);
nor U3023 (N_3023,N_2840,N_2843);
nand U3024 (N_3024,N_2959,N_2868);
or U3025 (N_3025,N_2870,N_2943);
xor U3026 (N_3026,N_2833,N_2936);
nor U3027 (N_3027,N_2966,N_2850);
and U3028 (N_3028,N_2938,N_2940);
nand U3029 (N_3029,N_2986,N_2969);
nor U3030 (N_3030,N_2953,N_2862);
nand U3031 (N_3031,N_2805,N_2809);
or U3032 (N_3032,N_2975,N_2838);
and U3033 (N_3033,N_2934,N_2849);
nand U3034 (N_3034,N_2928,N_2998);
xnor U3035 (N_3035,N_2902,N_2804);
or U3036 (N_3036,N_2949,N_2980);
and U3037 (N_3037,N_2841,N_2997);
nand U3038 (N_3038,N_2927,N_2929);
or U3039 (N_3039,N_2852,N_2967);
or U3040 (N_3040,N_2968,N_2948);
nand U3041 (N_3041,N_2925,N_2957);
xor U3042 (N_3042,N_2916,N_2880);
and U3043 (N_3043,N_2802,N_2832);
nand U3044 (N_3044,N_2917,N_2800);
nor U3045 (N_3045,N_2909,N_2877);
xnor U3046 (N_3046,N_2976,N_2879);
and U3047 (N_3047,N_2991,N_2978);
nand U3048 (N_3048,N_2820,N_2965);
or U3049 (N_3049,N_2963,N_2961);
nor U3050 (N_3050,N_2856,N_2945);
and U3051 (N_3051,N_2992,N_2989);
nand U3052 (N_3052,N_2922,N_2947);
xor U3053 (N_3053,N_2970,N_2995);
xor U3054 (N_3054,N_2801,N_2942);
nor U3055 (N_3055,N_2815,N_2896);
nor U3056 (N_3056,N_2999,N_2958);
or U3057 (N_3057,N_2918,N_2935);
nand U3058 (N_3058,N_2911,N_2872);
or U3059 (N_3059,N_2821,N_2834);
nor U3060 (N_3060,N_2982,N_2915);
and U3061 (N_3061,N_2895,N_2818);
xor U3062 (N_3062,N_2905,N_2885);
xor U3063 (N_3063,N_2831,N_2884);
nand U3064 (N_3064,N_2813,N_2823);
nor U3065 (N_3065,N_2853,N_2897);
xor U3066 (N_3066,N_2944,N_2977);
xor U3067 (N_3067,N_2814,N_2817);
nor U3068 (N_3068,N_2839,N_2867);
nand U3069 (N_3069,N_2913,N_2891);
nor U3070 (N_3070,N_2941,N_2808);
nor U3071 (N_3071,N_2984,N_2830);
or U3072 (N_3072,N_2924,N_2855);
nor U3073 (N_3073,N_2972,N_2828);
nor U3074 (N_3074,N_2990,N_2946);
nor U3075 (N_3075,N_2993,N_2865);
and U3076 (N_3076,N_2807,N_2881);
or U3077 (N_3077,N_2874,N_2848);
xor U3078 (N_3078,N_2861,N_2846);
nor U3079 (N_3079,N_2803,N_2894);
nand U3080 (N_3080,N_2931,N_2950);
and U3081 (N_3081,N_2835,N_2878);
or U3082 (N_3082,N_2914,N_2888);
xor U3083 (N_3083,N_2851,N_2854);
or U3084 (N_3084,N_2921,N_2873);
xnor U3085 (N_3085,N_2810,N_2930);
nor U3086 (N_3086,N_2952,N_2919);
or U3087 (N_3087,N_2981,N_2866);
or U3088 (N_3088,N_2824,N_2955);
nand U3089 (N_3089,N_2987,N_2806);
nor U3090 (N_3090,N_2858,N_2898);
or U3091 (N_3091,N_2923,N_2906);
and U3092 (N_3092,N_2811,N_2819);
or U3093 (N_3093,N_2842,N_2951);
or U3094 (N_3094,N_2907,N_2900);
nand U3095 (N_3095,N_2847,N_2826);
nor U3096 (N_3096,N_2933,N_2883);
or U3097 (N_3097,N_2875,N_2844);
or U3098 (N_3098,N_2926,N_2939);
nand U3099 (N_3099,N_2845,N_2837);
or U3100 (N_3100,N_2929,N_2808);
nor U3101 (N_3101,N_2888,N_2863);
or U3102 (N_3102,N_2870,N_2885);
nand U3103 (N_3103,N_2967,N_2935);
and U3104 (N_3104,N_2853,N_2990);
nand U3105 (N_3105,N_2992,N_2951);
nor U3106 (N_3106,N_2983,N_2813);
and U3107 (N_3107,N_2804,N_2890);
and U3108 (N_3108,N_2877,N_2905);
xnor U3109 (N_3109,N_2881,N_2895);
nand U3110 (N_3110,N_2820,N_2809);
or U3111 (N_3111,N_2901,N_2937);
and U3112 (N_3112,N_2915,N_2995);
nand U3113 (N_3113,N_2896,N_2897);
and U3114 (N_3114,N_2897,N_2975);
nor U3115 (N_3115,N_2864,N_2809);
nor U3116 (N_3116,N_2906,N_2862);
or U3117 (N_3117,N_2951,N_2958);
or U3118 (N_3118,N_2844,N_2924);
xnor U3119 (N_3119,N_2977,N_2952);
xnor U3120 (N_3120,N_2980,N_2846);
xor U3121 (N_3121,N_2930,N_2833);
and U3122 (N_3122,N_2875,N_2982);
or U3123 (N_3123,N_2968,N_2819);
nand U3124 (N_3124,N_2950,N_2862);
nor U3125 (N_3125,N_2913,N_2861);
nor U3126 (N_3126,N_2902,N_2899);
xor U3127 (N_3127,N_2871,N_2859);
nand U3128 (N_3128,N_2995,N_2823);
xor U3129 (N_3129,N_2946,N_2923);
xnor U3130 (N_3130,N_2883,N_2805);
and U3131 (N_3131,N_2988,N_2903);
nor U3132 (N_3132,N_2868,N_2940);
or U3133 (N_3133,N_2920,N_2857);
xnor U3134 (N_3134,N_2959,N_2891);
nand U3135 (N_3135,N_2921,N_2934);
and U3136 (N_3136,N_2816,N_2941);
nor U3137 (N_3137,N_2923,N_2893);
and U3138 (N_3138,N_2949,N_2996);
or U3139 (N_3139,N_2878,N_2842);
or U3140 (N_3140,N_2960,N_2869);
nand U3141 (N_3141,N_2964,N_2980);
nand U3142 (N_3142,N_2918,N_2824);
and U3143 (N_3143,N_2871,N_2990);
and U3144 (N_3144,N_2938,N_2832);
and U3145 (N_3145,N_2939,N_2911);
nand U3146 (N_3146,N_2926,N_2807);
xnor U3147 (N_3147,N_2815,N_2880);
and U3148 (N_3148,N_2879,N_2927);
and U3149 (N_3149,N_2889,N_2933);
nor U3150 (N_3150,N_2920,N_2989);
nor U3151 (N_3151,N_2977,N_2861);
xnor U3152 (N_3152,N_2809,N_2811);
and U3153 (N_3153,N_2934,N_2874);
or U3154 (N_3154,N_2898,N_2938);
nand U3155 (N_3155,N_2959,N_2885);
xor U3156 (N_3156,N_2917,N_2972);
xnor U3157 (N_3157,N_2969,N_2821);
and U3158 (N_3158,N_2891,N_2941);
nand U3159 (N_3159,N_2967,N_2891);
and U3160 (N_3160,N_2939,N_2856);
or U3161 (N_3161,N_2918,N_2838);
or U3162 (N_3162,N_2930,N_2946);
or U3163 (N_3163,N_2860,N_2959);
and U3164 (N_3164,N_2902,N_2861);
nand U3165 (N_3165,N_2967,N_2896);
nor U3166 (N_3166,N_2889,N_2856);
xnor U3167 (N_3167,N_2821,N_2980);
or U3168 (N_3168,N_2824,N_2938);
xor U3169 (N_3169,N_2814,N_2835);
nand U3170 (N_3170,N_2906,N_2982);
nand U3171 (N_3171,N_2822,N_2892);
nor U3172 (N_3172,N_2938,N_2950);
and U3173 (N_3173,N_2962,N_2825);
xnor U3174 (N_3174,N_2897,N_2806);
nor U3175 (N_3175,N_2875,N_2885);
xnor U3176 (N_3176,N_2820,N_2886);
xor U3177 (N_3177,N_2929,N_2825);
xnor U3178 (N_3178,N_2856,N_2910);
nand U3179 (N_3179,N_2944,N_2815);
or U3180 (N_3180,N_2870,N_2971);
xnor U3181 (N_3181,N_2863,N_2924);
xnor U3182 (N_3182,N_2930,N_2871);
or U3183 (N_3183,N_2832,N_2945);
and U3184 (N_3184,N_2907,N_2878);
or U3185 (N_3185,N_2997,N_2905);
nor U3186 (N_3186,N_2983,N_2928);
nand U3187 (N_3187,N_2912,N_2835);
or U3188 (N_3188,N_2977,N_2910);
xor U3189 (N_3189,N_2953,N_2917);
nand U3190 (N_3190,N_2832,N_2820);
nor U3191 (N_3191,N_2818,N_2840);
nand U3192 (N_3192,N_2808,N_2994);
or U3193 (N_3193,N_2903,N_2932);
and U3194 (N_3194,N_2991,N_2805);
and U3195 (N_3195,N_2831,N_2822);
xor U3196 (N_3196,N_2890,N_2905);
nor U3197 (N_3197,N_2923,N_2922);
or U3198 (N_3198,N_2936,N_2829);
nor U3199 (N_3199,N_2993,N_2859);
and U3200 (N_3200,N_3057,N_3171);
nor U3201 (N_3201,N_3160,N_3078);
nand U3202 (N_3202,N_3107,N_3106);
nor U3203 (N_3203,N_3101,N_3082);
nand U3204 (N_3204,N_3195,N_3175);
or U3205 (N_3205,N_3129,N_3115);
and U3206 (N_3206,N_3008,N_3026);
nor U3207 (N_3207,N_3164,N_3198);
or U3208 (N_3208,N_3173,N_3009);
nor U3209 (N_3209,N_3103,N_3169);
nor U3210 (N_3210,N_3095,N_3190);
xor U3211 (N_3211,N_3011,N_3109);
and U3212 (N_3212,N_3137,N_3077);
nor U3213 (N_3213,N_3093,N_3004);
xor U3214 (N_3214,N_3071,N_3127);
xnor U3215 (N_3215,N_3145,N_3174);
nor U3216 (N_3216,N_3079,N_3159);
nand U3217 (N_3217,N_3013,N_3100);
nand U3218 (N_3218,N_3142,N_3070);
or U3219 (N_3219,N_3177,N_3172);
or U3220 (N_3220,N_3181,N_3104);
and U3221 (N_3221,N_3135,N_3045);
nand U3222 (N_3222,N_3036,N_3182);
and U3223 (N_3223,N_3043,N_3199);
or U3224 (N_3224,N_3040,N_3147);
xnor U3225 (N_3225,N_3061,N_3167);
or U3226 (N_3226,N_3110,N_3179);
or U3227 (N_3227,N_3120,N_3131);
nor U3228 (N_3228,N_3000,N_3152);
xor U3229 (N_3229,N_3165,N_3053);
and U3230 (N_3230,N_3065,N_3023);
nor U3231 (N_3231,N_3184,N_3024);
or U3232 (N_3232,N_3039,N_3049);
and U3233 (N_3233,N_3192,N_3150);
or U3234 (N_3234,N_3168,N_3116);
or U3235 (N_3235,N_3016,N_3014);
or U3236 (N_3236,N_3094,N_3186);
and U3237 (N_3237,N_3075,N_3022);
xor U3238 (N_3238,N_3073,N_3037);
and U3239 (N_3239,N_3117,N_3090);
nor U3240 (N_3240,N_3108,N_3111);
and U3241 (N_3241,N_3193,N_3112);
xor U3242 (N_3242,N_3151,N_3149);
nand U3243 (N_3243,N_3085,N_3154);
or U3244 (N_3244,N_3146,N_3076);
nor U3245 (N_3245,N_3059,N_3069);
and U3246 (N_3246,N_3140,N_3124);
and U3247 (N_3247,N_3021,N_3087);
nor U3248 (N_3248,N_3178,N_3028);
xor U3249 (N_3249,N_3010,N_3047);
nor U3250 (N_3250,N_3044,N_3119);
and U3251 (N_3251,N_3084,N_3180);
nor U3252 (N_3252,N_3031,N_3089);
or U3253 (N_3253,N_3034,N_3176);
nor U3254 (N_3254,N_3126,N_3091);
nor U3255 (N_3255,N_3074,N_3088);
xor U3256 (N_3256,N_3144,N_3056);
xnor U3257 (N_3257,N_3033,N_3001);
and U3258 (N_3258,N_3003,N_3015);
xor U3259 (N_3259,N_3027,N_3141);
and U3260 (N_3260,N_3194,N_3157);
or U3261 (N_3261,N_3153,N_3136);
and U3262 (N_3262,N_3102,N_3122);
xnor U3263 (N_3263,N_3006,N_3138);
and U3264 (N_3264,N_3161,N_3187);
xor U3265 (N_3265,N_3098,N_3080);
and U3266 (N_3266,N_3051,N_3092);
and U3267 (N_3267,N_3018,N_3035);
nand U3268 (N_3268,N_3134,N_3196);
nand U3269 (N_3269,N_3066,N_3025);
nand U3270 (N_3270,N_3133,N_3096);
or U3271 (N_3271,N_3118,N_3029);
and U3272 (N_3272,N_3189,N_3019);
and U3273 (N_3273,N_3139,N_3097);
nand U3274 (N_3274,N_3060,N_3055);
xor U3275 (N_3275,N_3068,N_3067);
nand U3276 (N_3276,N_3185,N_3163);
or U3277 (N_3277,N_3063,N_3058);
or U3278 (N_3278,N_3128,N_3050);
nor U3279 (N_3279,N_3125,N_3064);
nor U3280 (N_3280,N_3046,N_3020);
and U3281 (N_3281,N_3072,N_3170);
nand U3282 (N_3282,N_3086,N_3123);
nand U3283 (N_3283,N_3042,N_3099);
nand U3284 (N_3284,N_3007,N_3143);
or U3285 (N_3285,N_3162,N_3155);
nor U3286 (N_3286,N_3197,N_3132);
or U3287 (N_3287,N_3062,N_3156);
nor U3288 (N_3288,N_3114,N_3002);
and U3289 (N_3289,N_3083,N_3191);
nand U3290 (N_3290,N_3121,N_3041);
nor U3291 (N_3291,N_3081,N_3048);
nand U3292 (N_3292,N_3030,N_3105);
or U3293 (N_3293,N_3183,N_3148);
xor U3294 (N_3294,N_3052,N_3054);
nor U3295 (N_3295,N_3032,N_3158);
nand U3296 (N_3296,N_3166,N_3005);
nand U3297 (N_3297,N_3012,N_3130);
xnor U3298 (N_3298,N_3038,N_3113);
and U3299 (N_3299,N_3188,N_3017);
and U3300 (N_3300,N_3163,N_3027);
xnor U3301 (N_3301,N_3079,N_3018);
and U3302 (N_3302,N_3182,N_3067);
nor U3303 (N_3303,N_3090,N_3093);
and U3304 (N_3304,N_3112,N_3002);
xnor U3305 (N_3305,N_3160,N_3092);
nor U3306 (N_3306,N_3121,N_3045);
nand U3307 (N_3307,N_3085,N_3046);
or U3308 (N_3308,N_3161,N_3083);
nand U3309 (N_3309,N_3092,N_3089);
or U3310 (N_3310,N_3011,N_3173);
or U3311 (N_3311,N_3033,N_3006);
xor U3312 (N_3312,N_3090,N_3122);
or U3313 (N_3313,N_3002,N_3190);
nor U3314 (N_3314,N_3089,N_3052);
nor U3315 (N_3315,N_3010,N_3082);
nor U3316 (N_3316,N_3103,N_3107);
and U3317 (N_3317,N_3068,N_3049);
and U3318 (N_3318,N_3006,N_3022);
or U3319 (N_3319,N_3058,N_3118);
nor U3320 (N_3320,N_3022,N_3154);
and U3321 (N_3321,N_3137,N_3075);
and U3322 (N_3322,N_3189,N_3015);
nor U3323 (N_3323,N_3026,N_3112);
nand U3324 (N_3324,N_3134,N_3168);
nor U3325 (N_3325,N_3193,N_3116);
or U3326 (N_3326,N_3054,N_3115);
and U3327 (N_3327,N_3167,N_3041);
or U3328 (N_3328,N_3132,N_3096);
and U3329 (N_3329,N_3042,N_3143);
nand U3330 (N_3330,N_3176,N_3166);
nand U3331 (N_3331,N_3173,N_3188);
or U3332 (N_3332,N_3041,N_3047);
nor U3333 (N_3333,N_3028,N_3144);
xnor U3334 (N_3334,N_3011,N_3107);
or U3335 (N_3335,N_3031,N_3155);
xor U3336 (N_3336,N_3002,N_3155);
nand U3337 (N_3337,N_3129,N_3152);
nand U3338 (N_3338,N_3043,N_3073);
and U3339 (N_3339,N_3185,N_3055);
xor U3340 (N_3340,N_3001,N_3101);
xor U3341 (N_3341,N_3001,N_3029);
and U3342 (N_3342,N_3110,N_3126);
xnor U3343 (N_3343,N_3069,N_3084);
xor U3344 (N_3344,N_3098,N_3084);
and U3345 (N_3345,N_3121,N_3197);
or U3346 (N_3346,N_3085,N_3111);
and U3347 (N_3347,N_3071,N_3178);
and U3348 (N_3348,N_3003,N_3027);
xnor U3349 (N_3349,N_3165,N_3036);
and U3350 (N_3350,N_3056,N_3018);
nor U3351 (N_3351,N_3031,N_3011);
xor U3352 (N_3352,N_3130,N_3187);
nand U3353 (N_3353,N_3120,N_3008);
and U3354 (N_3354,N_3029,N_3177);
xor U3355 (N_3355,N_3071,N_3106);
nor U3356 (N_3356,N_3062,N_3167);
nand U3357 (N_3357,N_3045,N_3138);
or U3358 (N_3358,N_3046,N_3194);
or U3359 (N_3359,N_3025,N_3173);
nor U3360 (N_3360,N_3152,N_3145);
xor U3361 (N_3361,N_3165,N_3070);
or U3362 (N_3362,N_3177,N_3021);
nand U3363 (N_3363,N_3160,N_3072);
xnor U3364 (N_3364,N_3177,N_3135);
and U3365 (N_3365,N_3182,N_3169);
nand U3366 (N_3366,N_3062,N_3189);
and U3367 (N_3367,N_3032,N_3120);
or U3368 (N_3368,N_3111,N_3183);
xor U3369 (N_3369,N_3143,N_3096);
xor U3370 (N_3370,N_3140,N_3040);
nand U3371 (N_3371,N_3125,N_3007);
nand U3372 (N_3372,N_3018,N_3048);
nor U3373 (N_3373,N_3053,N_3163);
and U3374 (N_3374,N_3044,N_3013);
nand U3375 (N_3375,N_3045,N_3009);
or U3376 (N_3376,N_3004,N_3032);
nor U3377 (N_3377,N_3140,N_3149);
or U3378 (N_3378,N_3078,N_3141);
and U3379 (N_3379,N_3064,N_3071);
nand U3380 (N_3380,N_3129,N_3195);
and U3381 (N_3381,N_3004,N_3185);
xnor U3382 (N_3382,N_3050,N_3129);
nor U3383 (N_3383,N_3017,N_3046);
nor U3384 (N_3384,N_3161,N_3060);
and U3385 (N_3385,N_3190,N_3147);
or U3386 (N_3386,N_3128,N_3082);
xnor U3387 (N_3387,N_3148,N_3068);
nor U3388 (N_3388,N_3185,N_3023);
nand U3389 (N_3389,N_3163,N_3064);
or U3390 (N_3390,N_3193,N_3170);
nand U3391 (N_3391,N_3123,N_3050);
nor U3392 (N_3392,N_3107,N_3169);
nand U3393 (N_3393,N_3172,N_3085);
nor U3394 (N_3394,N_3080,N_3177);
xor U3395 (N_3395,N_3134,N_3024);
and U3396 (N_3396,N_3174,N_3107);
nor U3397 (N_3397,N_3001,N_3066);
nand U3398 (N_3398,N_3067,N_3103);
nand U3399 (N_3399,N_3077,N_3058);
nand U3400 (N_3400,N_3285,N_3226);
nand U3401 (N_3401,N_3224,N_3336);
nand U3402 (N_3402,N_3225,N_3278);
and U3403 (N_3403,N_3311,N_3379);
xor U3404 (N_3404,N_3363,N_3389);
nand U3405 (N_3405,N_3206,N_3367);
xor U3406 (N_3406,N_3297,N_3323);
and U3407 (N_3407,N_3364,N_3240);
nand U3408 (N_3408,N_3228,N_3324);
nor U3409 (N_3409,N_3348,N_3231);
xor U3410 (N_3410,N_3306,N_3229);
and U3411 (N_3411,N_3244,N_3261);
xnor U3412 (N_3412,N_3316,N_3203);
nor U3413 (N_3413,N_3289,N_3235);
xor U3414 (N_3414,N_3345,N_3390);
or U3415 (N_3415,N_3309,N_3254);
nor U3416 (N_3416,N_3227,N_3330);
nand U3417 (N_3417,N_3239,N_3256);
nand U3418 (N_3418,N_3317,N_3201);
nor U3419 (N_3419,N_3214,N_3322);
or U3420 (N_3420,N_3283,N_3352);
xor U3421 (N_3421,N_3211,N_3304);
nor U3422 (N_3422,N_3359,N_3375);
and U3423 (N_3423,N_3313,N_3249);
or U3424 (N_3424,N_3277,N_3246);
nand U3425 (N_3425,N_3268,N_3370);
nor U3426 (N_3426,N_3286,N_3262);
xor U3427 (N_3427,N_3325,N_3288);
nand U3428 (N_3428,N_3310,N_3360);
nor U3429 (N_3429,N_3276,N_3343);
or U3430 (N_3430,N_3307,N_3340);
nand U3431 (N_3431,N_3368,N_3333);
nand U3432 (N_3432,N_3280,N_3314);
and U3433 (N_3433,N_3216,N_3346);
xnor U3434 (N_3434,N_3291,N_3386);
nor U3435 (N_3435,N_3397,N_3217);
nor U3436 (N_3436,N_3273,N_3385);
nor U3437 (N_3437,N_3362,N_3351);
and U3438 (N_3438,N_3237,N_3319);
and U3439 (N_3439,N_3296,N_3275);
nand U3440 (N_3440,N_3393,N_3308);
and U3441 (N_3441,N_3281,N_3234);
nor U3442 (N_3442,N_3326,N_3220);
and U3443 (N_3443,N_3335,N_3354);
nand U3444 (N_3444,N_3361,N_3248);
nand U3445 (N_3445,N_3315,N_3271);
xor U3446 (N_3446,N_3342,N_3259);
nor U3447 (N_3447,N_3384,N_3238);
nand U3448 (N_3448,N_3312,N_3236);
xnor U3449 (N_3449,N_3295,N_3202);
or U3450 (N_3450,N_3245,N_3210);
nand U3451 (N_3451,N_3394,N_3279);
and U3452 (N_3452,N_3301,N_3365);
xor U3453 (N_3453,N_3218,N_3318);
xor U3454 (N_3454,N_3358,N_3272);
nor U3455 (N_3455,N_3242,N_3221);
xnor U3456 (N_3456,N_3305,N_3392);
xnor U3457 (N_3457,N_3266,N_3327);
nor U3458 (N_3458,N_3264,N_3366);
nor U3459 (N_3459,N_3398,N_3356);
xnor U3460 (N_3460,N_3265,N_3292);
and U3461 (N_3461,N_3357,N_3294);
xor U3462 (N_3462,N_3208,N_3205);
and U3463 (N_3463,N_3267,N_3349);
or U3464 (N_3464,N_3391,N_3320);
xor U3465 (N_3465,N_3274,N_3223);
xor U3466 (N_3466,N_3269,N_3258);
or U3467 (N_3467,N_3230,N_3396);
xnor U3468 (N_3468,N_3353,N_3260);
nand U3469 (N_3469,N_3382,N_3350);
xor U3470 (N_3470,N_3251,N_3247);
nand U3471 (N_3471,N_3282,N_3290);
or U3472 (N_3472,N_3207,N_3383);
or U3473 (N_3473,N_3344,N_3388);
xnor U3474 (N_3474,N_3284,N_3222);
nand U3475 (N_3475,N_3334,N_3372);
or U3476 (N_3476,N_3253,N_3329);
xor U3477 (N_3477,N_3341,N_3232);
xnor U3478 (N_3478,N_3243,N_3300);
xor U3479 (N_3479,N_3212,N_3287);
and U3480 (N_3480,N_3255,N_3338);
nand U3481 (N_3481,N_3257,N_3250);
or U3482 (N_3482,N_3219,N_3378);
nand U3483 (N_3483,N_3399,N_3339);
nor U3484 (N_3484,N_3371,N_3215);
xor U3485 (N_3485,N_3328,N_3204);
xnor U3486 (N_3486,N_3270,N_3331);
or U3487 (N_3487,N_3387,N_3209);
nand U3488 (N_3488,N_3321,N_3263);
or U3489 (N_3489,N_3369,N_3302);
nor U3490 (N_3490,N_3380,N_3347);
nor U3491 (N_3491,N_3332,N_3355);
nand U3492 (N_3492,N_3303,N_3381);
or U3493 (N_3493,N_3241,N_3299);
and U3494 (N_3494,N_3252,N_3395);
nand U3495 (N_3495,N_3337,N_3293);
xor U3496 (N_3496,N_3200,N_3298);
and U3497 (N_3497,N_3376,N_3233);
nor U3498 (N_3498,N_3377,N_3213);
or U3499 (N_3499,N_3374,N_3373);
nand U3500 (N_3500,N_3318,N_3394);
nor U3501 (N_3501,N_3323,N_3368);
xnor U3502 (N_3502,N_3394,N_3334);
xor U3503 (N_3503,N_3216,N_3347);
nor U3504 (N_3504,N_3202,N_3382);
or U3505 (N_3505,N_3320,N_3363);
or U3506 (N_3506,N_3280,N_3381);
nand U3507 (N_3507,N_3298,N_3253);
nand U3508 (N_3508,N_3248,N_3360);
nor U3509 (N_3509,N_3251,N_3234);
and U3510 (N_3510,N_3262,N_3386);
nand U3511 (N_3511,N_3244,N_3307);
and U3512 (N_3512,N_3279,N_3241);
or U3513 (N_3513,N_3330,N_3344);
and U3514 (N_3514,N_3326,N_3292);
xor U3515 (N_3515,N_3303,N_3345);
nor U3516 (N_3516,N_3324,N_3346);
nor U3517 (N_3517,N_3285,N_3283);
and U3518 (N_3518,N_3382,N_3206);
xor U3519 (N_3519,N_3204,N_3386);
or U3520 (N_3520,N_3233,N_3294);
and U3521 (N_3521,N_3255,N_3292);
xnor U3522 (N_3522,N_3380,N_3393);
nand U3523 (N_3523,N_3292,N_3202);
nand U3524 (N_3524,N_3282,N_3210);
nand U3525 (N_3525,N_3345,N_3353);
nand U3526 (N_3526,N_3249,N_3225);
nor U3527 (N_3527,N_3216,N_3376);
nand U3528 (N_3528,N_3364,N_3369);
xnor U3529 (N_3529,N_3324,N_3311);
nand U3530 (N_3530,N_3239,N_3322);
xor U3531 (N_3531,N_3314,N_3340);
and U3532 (N_3532,N_3307,N_3320);
or U3533 (N_3533,N_3285,N_3372);
or U3534 (N_3534,N_3357,N_3380);
nand U3535 (N_3535,N_3207,N_3277);
and U3536 (N_3536,N_3216,N_3258);
xnor U3537 (N_3537,N_3322,N_3345);
or U3538 (N_3538,N_3219,N_3351);
nor U3539 (N_3539,N_3246,N_3398);
and U3540 (N_3540,N_3290,N_3387);
nand U3541 (N_3541,N_3316,N_3367);
nor U3542 (N_3542,N_3253,N_3275);
nand U3543 (N_3543,N_3245,N_3363);
or U3544 (N_3544,N_3320,N_3295);
nor U3545 (N_3545,N_3318,N_3385);
xnor U3546 (N_3546,N_3365,N_3312);
nor U3547 (N_3547,N_3346,N_3247);
or U3548 (N_3548,N_3332,N_3366);
nor U3549 (N_3549,N_3258,N_3252);
xnor U3550 (N_3550,N_3338,N_3208);
and U3551 (N_3551,N_3245,N_3300);
nand U3552 (N_3552,N_3235,N_3357);
nor U3553 (N_3553,N_3217,N_3325);
nand U3554 (N_3554,N_3327,N_3226);
nand U3555 (N_3555,N_3360,N_3279);
nand U3556 (N_3556,N_3297,N_3305);
nor U3557 (N_3557,N_3229,N_3257);
nand U3558 (N_3558,N_3245,N_3213);
or U3559 (N_3559,N_3384,N_3324);
and U3560 (N_3560,N_3222,N_3200);
or U3561 (N_3561,N_3241,N_3264);
nor U3562 (N_3562,N_3323,N_3202);
nand U3563 (N_3563,N_3249,N_3288);
nor U3564 (N_3564,N_3245,N_3351);
and U3565 (N_3565,N_3332,N_3309);
or U3566 (N_3566,N_3324,N_3304);
nand U3567 (N_3567,N_3209,N_3384);
nand U3568 (N_3568,N_3280,N_3210);
or U3569 (N_3569,N_3372,N_3295);
nor U3570 (N_3570,N_3204,N_3201);
and U3571 (N_3571,N_3284,N_3341);
and U3572 (N_3572,N_3346,N_3350);
nor U3573 (N_3573,N_3259,N_3399);
xor U3574 (N_3574,N_3204,N_3308);
nand U3575 (N_3575,N_3359,N_3336);
nand U3576 (N_3576,N_3322,N_3313);
xnor U3577 (N_3577,N_3279,N_3327);
or U3578 (N_3578,N_3368,N_3375);
xnor U3579 (N_3579,N_3302,N_3380);
nor U3580 (N_3580,N_3205,N_3250);
xor U3581 (N_3581,N_3366,N_3284);
or U3582 (N_3582,N_3390,N_3326);
xnor U3583 (N_3583,N_3358,N_3315);
and U3584 (N_3584,N_3260,N_3336);
nor U3585 (N_3585,N_3305,N_3364);
and U3586 (N_3586,N_3335,N_3273);
nand U3587 (N_3587,N_3327,N_3364);
and U3588 (N_3588,N_3231,N_3207);
nand U3589 (N_3589,N_3281,N_3212);
nor U3590 (N_3590,N_3202,N_3332);
or U3591 (N_3591,N_3340,N_3257);
nand U3592 (N_3592,N_3340,N_3342);
and U3593 (N_3593,N_3382,N_3277);
nand U3594 (N_3594,N_3317,N_3260);
nand U3595 (N_3595,N_3232,N_3226);
and U3596 (N_3596,N_3331,N_3328);
or U3597 (N_3597,N_3239,N_3295);
nand U3598 (N_3598,N_3214,N_3387);
and U3599 (N_3599,N_3279,N_3313);
and U3600 (N_3600,N_3490,N_3512);
nand U3601 (N_3601,N_3539,N_3535);
nand U3602 (N_3602,N_3408,N_3514);
nand U3603 (N_3603,N_3523,N_3592);
nor U3604 (N_3604,N_3566,N_3529);
nand U3605 (N_3605,N_3568,N_3434);
nand U3606 (N_3606,N_3530,N_3405);
or U3607 (N_3607,N_3465,N_3540);
nand U3608 (N_3608,N_3551,N_3517);
or U3609 (N_3609,N_3581,N_3435);
and U3610 (N_3610,N_3450,N_3491);
xnor U3611 (N_3611,N_3596,N_3467);
xnor U3612 (N_3612,N_3446,N_3502);
xnor U3613 (N_3613,N_3456,N_3474);
or U3614 (N_3614,N_3485,N_3559);
nand U3615 (N_3615,N_3426,N_3400);
xor U3616 (N_3616,N_3584,N_3580);
xor U3617 (N_3617,N_3532,N_3413);
nor U3618 (N_3618,N_3407,N_3455);
or U3619 (N_3619,N_3445,N_3571);
and U3620 (N_3620,N_3507,N_3578);
or U3621 (N_3621,N_3424,N_3531);
xor U3622 (N_3622,N_3401,N_3542);
nor U3623 (N_3623,N_3563,N_3573);
nor U3624 (N_3624,N_3481,N_3437);
and U3625 (N_3625,N_3569,N_3494);
nand U3626 (N_3626,N_3585,N_3545);
nor U3627 (N_3627,N_3546,N_3589);
or U3628 (N_3628,N_3564,N_3453);
nor U3629 (N_3629,N_3448,N_3582);
and U3630 (N_3630,N_3440,N_3489);
nor U3631 (N_3631,N_3417,N_3570);
nor U3632 (N_3632,N_3469,N_3537);
and U3633 (N_3633,N_3572,N_3479);
xnor U3634 (N_3634,N_3428,N_3493);
or U3635 (N_3635,N_3470,N_3510);
or U3636 (N_3636,N_3555,N_3526);
and U3637 (N_3637,N_3432,N_3567);
xor U3638 (N_3638,N_3454,N_3439);
nand U3639 (N_3639,N_3460,N_3499);
nor U3640 (N_3640,N_3548,N_3403);
nor U3641 (N_3641,N_3466,N_3505);
nand U3642 (N_3642,N_3597,N_3484);
nor U3643 (N_3643,N_3541,N_3519);
nor U3644 (N_3644,N_3420,N_3528);
and U3645 (N_3645,N_3444,N_3560);
xnor U3646 (N_3646,N_3482,N_3475);
and U3647 (N_3647,N_3588,N_3504);
nand U3648 (N_3648,N_3558,N_3521);
nor U3649 (N_3649,N_3509,N_3525);
or U3650 (N_3650,N_3503,N_3576);
nor U3651 (N_3651,N_3590,N_3462);
xor U3652 (N_3652,N_3463,N_3488);
nand U3653 (N_3653,N_3579,N_3561);
xor U3654 (N_3654,N_3430,N_3425);
xnor U3655 (N_3655,N_3511,N_3574);
nor U3656 (N_3656,N_3423,N_3552);
and U3657 (N_3657,N_3575,N_3508);
nor U3658 (N_3658,N_3506,N_3442);
nand U3659 (N_3659,N_3459,N_3583);
nand U3660 (N_3660,N_3543,N_3538);
nor U3661 (N_3661,N_3419,N_3477);
nand U3662 (N_3662,N_3422,N_3553);
or U3663 (N_3663,N_3410,N_3554);
nand U3664 (N_3664,N_3480,N_3468);
xor U3665 (N_3665,N_3565,N_3577);
nor U3666 (N_3666,N_3522,N_3486);
and U3667 (N_3667,N_3527,N_3429);
or U3668 (N_3668,N_3436,N_3472);
nor U3669 (N_3669,N_3595,N_3427);
nand U3670 (N_3670,N_3478,N_3449);
nor U3671 (N_3671,N_3498,N_3534);
and U3672 (N_3672,N_3515,N_3409);
or U3673 (N_3673,N_3536,N_3412);
and U3674 (N_3674,N_3587,N_3441);
or U3675 (N_3675,N_3451,N_3524);
or U3676 (N_3676,N_3549,N_3483);
or U3677 (N_3677,N_3495,N_3599);
nor U3678 (N_3678,N_3447,N_3402);
or U3679 (N_3679,N_3598,N_3418);
nand U3680 (N_3680,N_3421,N_3433);
and U3681 (N_3681,N_3438,N_3547);
xnor U3682 (N_3682,N_3458,N_3593);
nand U3683 (N_3683,N_3557,N_3594);
xor U3684 (N_3684,N_3520,N_3416);
nor U3685 (N_3685,N_3544,N_3591);
and U3686 (N_3686,N_3464,N_3586);
xor U3687 (N_3687,N_3501,N_3457);
nand U3688 (N_3688,N_3497,N_3518);
xnor U3689 (N_3689,N_3487,N_3533);
and U3690 (N_3690,N_3550,N_3473);
nor U3691 (N_3691,N_3496,N_3513);
nand U3692 (N_3692,N_3500,N_3406);
and U3693 (N_3693,N_3556,N_3404);
nand U3694 (N_3694,N_3411,N_3461);
xnor U3695 (N_3695,N_3443,N_3431);
nor U3696 (N_3696,N_3516,N_3476);
nand U3697 (N_3697,N_3492,N_3452);
and U3698 (N_3698,N_3415,N_3414);
or U3699 (N_3699,N_3562,N_3471);
or U3700 (N_3700,N_3419,N_3466);
nor U3701 (N_3701,N_3446,N_3568);
or U3702 (N_3702,N_3472,N_3457);
xor U3703 (N_3703,N_3416,N_3568);
and U3704 (N_3704,N_3509,N_3425);
nand U3705 (N_3705,N_3455,N_3599);
and U3706 (N_3706,N_3455,N_3558);
nand U3707 (N_3707,N_3488,N_3424);
xor U3708 (N_3708,N_3477,N_3476);
xor U3709 (N_3709,N_3489,N_3433);
nor U3710 (N_3710,N_3581,N_3575);
and U3711 (N_3711,N_3452,N_3453);
nor U3712 (N_3712,N_3467,N_3494);
and U3713 (N_3713,N_3587,N_3469);
or U3714 (N_3714,N_3521,N_3524);
xnor U3715 (N_3715,N_3442,N_3406);
or U3716 (N_3716,N_3469,N_3536);
nand U3717 (N_3717,N_3451,N_3458);
nor U3718 (N_3718,N_3402,N_3488);
xor U3719 (N_3719,N_3504,N_3584);
nand U3720 (N_3720,N_3550,N_3493);
or U3721 (N_3721,N_3452,N_3478);
or U3722 (N_3722,N_3547,N_3474);
xnor U3723 (N_3723,N_3552,N_3462);
nor U3724 (N_3724,N_3502,N_3499);
nand U3725 (N_3725,N_3491,N_3582);
xnor U3726 (N_3726,N_3494,N_3401);
nand U3727 (N_3727,N_3544,N_3419);
or U3728 (N_3728,N_3429,N_3508);
nor U3729 (N_3729,N_3464,N_3432);
and U3730 (N_3730,N_3530,N_3541);
xor U3731 (N_3731,N_3498,N_3592);
xnor U3732 (N_3732,N_3406,N_3529);
or U3733 (N_3733,N_3426,N_3526);
xor U3734 (N_3734,N_3538,N_3514);
or U3735 (N_3735,N_3480,N_3440);
or U3736 (N_3736,N_3537,N_3459);
or U3737 (N_3737,N_3480,N_3509);
nor U3738 (N_3738,N_3541,N_3460);
xor U3739 (N_3739,N_3470,N_3574);
nor U3740 (N_3740,N_3416,N_3536);
xor U3741 (N_3741,N_3528,N_3404);
nand U3742 (N_3742,N_3413,N_3558);
nor U3743 (N_3743,N_3499,N_3556);
nor U3744 (N_3744,N_3558,N_3587);
nand U3745 (N_3745,N_3473,N_3500);
and U3746 (N_3746,N_3534,N_3486);
nor U3747 (N_3747,N_3584,N_3402);
nand U3748 (N_3748,N_3467,N_3406);
and U3749 (N_3749,N_3534,N_3400);
and U3750 (N_3750,N_3553,N_3566);
xnor U3751 (N_3751,N_3529,N_3564);
or U3752 (N_3752,N_3526,N_3592);
or U3753 (N_3753,N_3543,N_3585);
or U3754 (N_3754,N_3516,N_3452);
nor U3755 (N_3755,N_3437,N_3514);
or U3756 (N_3756,N_3483,N_3545);
or U3757 (N_3757,N_3505,N_3584);
nor U3758 (N_3758,N_3441,N_3446);
or U3759 (N_3759,N_3451,N_3528);
or U3760 (N_3760,N_3543,N_3568);
and U3761 (N_3761,N_3464,N_3560);
xor U3762 (N_3762,N_3533,N_3445);
nand U3763 (N_3763,N_3404,N_3454);
nor U3764 (N_3764,N_3560,N_3406);
and U3765 (N_3765,N_3514,N_3400);
nand U3766 (N_3766,N_3468,N_3405);
nand U3767 (N_3767,N_3543,N_3508);
nor U3768 (N_3768,N_3534,N_3480);
or U3769 (N_3769,N_3518,N_3441);
nor U3770 (N_3770,N_3428,N_3474);
xnor U3771 (N_3771,N_3496,N_3431);
nand U3772 (N_3772,N_3516,N_3478);
nand U3773 (N_3773,N_3420,N_3407);
xor U3774 (N_3774,N_3509,N_3554);
or U3775 (N_3775,N_3445,N_3408);
and U3776 (N_3776,N_3554,N_3563);
nor U3777 (N_3777,N_3478,N_3412);
nor U3778 (N_3778,N_3529,N_3555);
or U3779 (N_3779,N_3487,N_3502);
or U3780 (N_3780,N_3535,N_3432);
or U3781 (N_3781,N_3494,N_3532);
nand U3782 (N_3782,N_3553,N_3530);
or U3783 (N_3783,N_3403,N_3549);
xor U3784 (N_3784,N_3446,N_3456);
nand U3785 (N_3785,N_3408,N_3569);
nand U3786 (N_3786,N_3572,N_3598);
nand U3787 (N_3787,N_3467,N_3443);
and U3788 (N_3788,N_3443,N_3474);
and U3789 (N_3789,N_3502,N_3556);
xnor U3790 (N_3790,N_3473,N_3414);
or U3791 (N_3791,N_3553,N_3406);
xnor U3792 (N_3792,N_3596,N_3468);
nor U3793 (N_3793,N_3546,N_3561);
nand U3794 (N_3794,N_3576,N_3573);
and U3795 (N_3795,N_3597,N_3459);
nor U3796 (N_3796,N_3572,N_3503);
nand U3797 (N_3797,N_3511,N_3556);
xor U3798 (N_3798,N_3412,N_3411);
nor U3799 (N_3799,N_3478,N_3528);
and U3800 (N_3800,N_3789,N_3631);
xor U3801 (N_3801,N_3669,N_3754);
and U3802 (N_3802,N_3647,N_3656);
xor U3803 (N_3803,N_3701,N_3751);
xnor U3804 (N_3804,N_3756,N_3663);
or U3805 (N_3805,N_3779,N_3630);
and U3806 (N_3806,N_3609,N_3627);
nand U3807 (N_3807,N_3739,N_3658);
nor U3808 (N_3808,N_3797,N_3712);
nand U3809 (N_3809,N_3752,N_3679);
nand U3810 (N_3810,N_3776,N_3649);
or U3811 (N_3811,N_3648,N_3675);
or U3812 (N_3812,N_3621,N_3721);
nor U3813 (N_3813,N_3623,N_3792);
or U3814 (N_3814,N_3693,N_3654);
nor U3815 (N_3815,N_3733,N_3676);
or U3816 (N_3816,N_3603,N_3750);
nand U3817 (N_3817,N_3662,N_3753);
and U3818 (N_3818,N_3683,N_3682);
xor U3819 (N_3819,N_3723,N_3601);
and U3820 (N_3820,N_3607,N_3747);
xor U3821 (N_3821,N_3722,N_3700);
or U3822 (N_3822,N_3742,N_3794);
xor U3823 (N_3823,N_3714,N_3695);
xor U3824 (N_3824,N_3681,N_3689);
xor U3825 (N_3825,N_3671,N_3674);
xnor U3826 (N_3826,N_3613,N_3771);
and U3827 (N_3827,N_3767,N_3760);
and U3828 (N_3828,N_3785,N_3705);
and U3829 (N_3829,N_3762,N_3680);
nor U3830 (N_3830,N_3636,N_3717);
nand U3831 (N_3831,N_3790,N_3773);
nor U3832 (N_3832,N_3659,N_3703);
nand U3833 (N_3833,N_3638,N_3637);
and U3834 (N_3834,N_3708,N_3726);
nand U3835 (N_3835,N_3799,N_3706);
nand U3836 (N_3836,N_3644,N_3634);
or U3837 (N_3837,N_3774,N_3786);
nor U3838 (N_3838,N_3670,N_3611);
or U3839 (N_3839,N_3687,N_3778);
or U3840 (N_3840,N_3657,N_3664);
nand U3841 (N_3841,N_3749,N_3718);
nor U3842 (N_3842,N_3617,N_3795);
and U3843 (N_3843,N_3653,N_3793);
nand U3844 (N_3844,N_3781,N_3748);
and U3845 (N_3845,N_3622,N_3612);
nor U3846 (N_3846,N_3764,N_3791);
xor U3847 (N_3847,N_3772,N_3672);
xnor U3848 (N_3848,N_3709,N_3650);
or U3849 (N_3849,N_3668,N_3602);
nand U3850 (N_3850,N_3730,N_3732);
xor U3851 (N_3851,N_3758,N_3645);
nand U3852 (N_3852,N_3796,N_3755);
or U3853 (N_3853,N_3608,N_3619);
xnor U3854 (N_3854,N_3702,N_3652);
nor U3855 (N_3855,N_3615,N_3735);
nand U3856 (N_3856,N_3620,N_3698);
or U3857 (N_3857,N_3690,N_3763);
or U3858 (N_3858,N_3677,N_3729);
and U3859 (N_3859,N_3624,N_3744);
and U3860 (N_3860,N_3770,N_3777);
nor U3861 (N_3861,N_3798,N_3741);
xor U3862 (N_3862,N_3768,N_3719);
nor U3863 (N_3863,N_3710,N_3605);
or U3864 (N_3864,N_3673,N_3745);
and U3865 (N_3865,N_3610,N_3699);
nand U3866 (N_3866,N_3655,N_3626);
and U3867 (N_3867,N_3736,N_3757);
xor U3868 (N_3868,N_3665,N_3784);
nand U3869 (N_3869,N_3775,N_3715);
nor U3870 (N_3870,N_3787,N_3720);
nor U3871 (N_3871,N_3604,N_3641);
xor U3872 (N_3872,N_3711,N_3704);
or U3873 (N_3873,N_3731,N_3783);
nand U3874 (N_3874,N_3625,N_3766);
xnor U3875 (N_3875,N_3628,N_3788);
nor U3876 (N_3876,N_3769,N_3614);
or U3877 (N_3877,N_3606,N_3684);
and U3878 (N_3878,N_3632,N_3643);
and U3879 (N_3879,N_3743,N_3651);
xnor U3880 (N_3880,N_3688,N_3780);
or U3881 (N_3881,N_3734,N_3765);
nor U3882 (N_3882,N_3759,N_3666);
and U3883 (N_3883,N_3691,N_3697);
or U3884 (N_3884,N_3782,N_3616);
or U3885 (N_3885,N_3633,N_3635);
or U3886 (N_3886,N_3678,N_3696);
and U3887 (N_3887,N_3737,N_3707);
or U3888 (N_3888,N_3728,N_3713);
and U3889 (N_3889,N_3642,N_3716);
and U3890 (N_3890,N_3740,N_3667);
nor U3891 (N_3891,N_3640,N_3738);
and U3892 (N_3892,N_3686,N_3725);
and U3893 (N_3893,N_3660,N_3761);
and U3894 (N_3894,N_3694,N_3724);
and U3895 (N_3895,N_3746,N_3646);
and U3896 (N_3896,N_3618,N_3661);
xnor U3897 (N_3897,N_3629,N_3692);
nor U3898 (N_3898,N_3600,N_3639);
and U3899 (N_3899,N_3727,N_3685);
or U3900 (N_3900,N_3747,N_3788);
nand U3901 (N_3901,N_3731,N_3793);
xnor U3902 (N_3902,N_3717,N_3777);
xor U3903 (N_3903,N_3703,N_3702);
nand U3904 (N_3904,N_3634,N_3696);
and U3905 (N_3905,N_3755,N_3624);
nor U3906 (N_3906,N_3670,N_3766);
or U3907 (N_3907,N_3656,N_3657);
and U3908 (N_3908,N_3649,N_3722);
and U3909 (N_3909,N_3692,N_3621);
nand U3910 (N_3910,N_3780,N_3673);
nor U3911 (N_3911,N_3788,N_3709);
nor U3912 (N_3912,N_3687,N_3710);
or U3913 (N_3913,N_3651,N_3641);
nor U3914 (N_3914,N_3790,N_3609);
and U3915 (N_3915,N_3725,N_3741);
and U3916 (N_3916,N_3719,N_3648);
nand U3917 (N_3917,N_3768,N_3684);
and U3918 (N_3918,N_3634,N_3648);
nor U3919 (N_3919,N_3674,N_3758);
nor U3920 (N_3920,N_3665,N_3652);
or U3921 (N_3921,N_3692,N_3757);
nand U3922 (N_3922,N_3771,N_3707);
nand U3923 (N_3923,N_3627,N_3774);
and U3924 (N_3924,N_3724,N_3761);
and U3925 (N_3925,N_3637,N_3713);
or U3926 (N_3926,N_3754,N_3724);
xor U3927 (N_3927,N_3641,N_3628);
nor U3928 (N_3928,N_3635,N_3701);
or U3929 (N_3929,N_3717,N_3715);
xor U3930 (N_3930,N_3762,N_3655);
or U3931 (N_3931,N_3645,N_3651);
and U3932 (N_3932,N_3779,N_3660);
nor U3933 (N_3933,N_3752,N_3730);
or U3934 (N_3934,N_3744,N_3746);
nand U3935 (N_3935,N_3668,N_3675);
and U3936 (N_3936,N_3751,N_3624);
and U3937 (N_3937,N_3743,N_3716);
xnor U3938 (N_3938,N_3634,N_3771);
nor U3939 (N_3939,N_3732,N_3745);
and U3940 (N_3940,N_3679,N_3716);
nor U3941 (N_3941,N_3793,N_3776);
nand U3942 (N_3942,N_3611,N_3704);
and U3943 (N_3943,N_3701,N_3663);
nor U3944 (N_3944,N_3696,N_3759);
nor U3945 (N_3945,N_3773,N_3642);
and U3946 (N_3946,N_3772,N_3708);
and U3947 (N_3947,N_3769,N_3764);
nand U3948 (N_3948,N_3756,N_3718);
or U3949 (N_3949,N_3794,N_3723);
nor U3950 (N_3950,N_3615,N_3696);
nor U3951 (N_3951,N_3668,N_3749);
and U3952 (N_3952,N_3740,N_3765);
nor U3953 (N_3953,N_3619,N_3749);
nand U3954 (N_3954,N_3654,N_3757);
xnor U3955 (N_3955,N_3703,N_3686);
xor U3956 (N_3956,N_3632,N_3647);
nand U3957 (N_3957,N_3785,N_3660);
xor U3958 (N_3958,N_3651,N_3610);
nor U3959 (N_3959,N_3676,N_3694);
and U3960 (N_3960,N_3763,N_3757);
or U3961 (N_3961,N_3690,N_3696);
or U3962 (N_3962,N_3644,N_3779);
nand U3963 (N_3963,N_3715,N_3609);
or U3964 (N_3964,N_3733,N_3794);
or U3965 (N_3965,N_3747,N_3660);
and U3966 (N_3966,N_3722,N_3784);
or U3967 (N_3967,N_3783,N_3796);
nor U3968 (N_3968,N_3796,N_3602);
nand U3969 (N_3969,N_3702,N_3642);
or U3970 (N_3970,N_3658,N_3758);
nor U3971 (N_3971,N_3705,N_3668);
or U3972 (N_3972,N_3758,N_3727);
nor U3973 (N_3973,N_3646,N_3612);
xor U3974 (N_3974,N_3706,N_3731);
or U3975 (N_3975,N_3621,N_3695);
or U3976 (N_3976,N_3772,N_3641);
nor U3977 (N_3977,N_3689,N_3795);
and U3978 (N_3978,N_3727,N_3601);
or U3979 (N_3979,N_3768,N_3623);
or U3980 (N_3980,N_3766,N_3770);
xnor U3981 (N_3981,N_3615,N_3796);
xnor U3982 (N_3982,N_3752,N_3795);
xnor U3983 (N_3983,N_3790,N_3612);
nor U3984 (N_3984,N_3717,N_3713);
nor U3985 (N_3985,N_3631,N_3655);
or U3986 (N_3986,N_3697,N_3630);
nand U3987 (N_3987,N_3789,N_3661);
or U3988 (N_3988,N_3605,N_3681);
xor U3989 (N_3989,N_3743,N_3722);
nand U3990 (N_3990,N_3682,N_3723);
xor U3991 (N_3991,N_3757,N_3708);
nor U3992 (N_3992,N_3647,N_3682);
and U3993 (N_3993,N_3613,N_3607);
or U3994 (N_3994,N_3644,N_3793);
nor U3995 (N_3995,N_3626,N_3693);
and U3996 (N_3996,N_3620,N_3641);
xnor U3997 (N_3997,N_3649,N_3760);
nand U3998 (N_3998,N_3696,N_3622);
and U3999 (N_3999,N_3793,N_3715);
nand U4000 (N_4000,N_3841,N_3960);
nand U4001 (N_4001,N_3923,N_3868);
and U4002 (N_4002,N_3954,N_3878);
nor U4003 (N_4003,N_3989,N_3850);
and U4004 (N_4004,N_3867,N_3958);
nand U4005 (N_4005,N_3908,N_3971);
and U4006 (N_4006,N_3838,N_3973);
nand U4007 (N_4007,N_3849,N_3826);
and U4008 (N_4008,N_3800,N_3986);
or U4009 (N_4009,N_3987,N_3982);
xor U4010 (N_4010,N_3992,N_3913);
and U4011 (N_4011,N_3802,N_3970);
xor U4012 (N_4012,N_3926,N_3824);
xnor U4013 (N_4013,N_3822,N_3904);
nor U4014 (N_4014,N_3962,N_3927);
nor U4015 (N_4015,N_3864,N_3993);
xnor U4016 (N_4016,N_3874,N_3832);
xnor U4017 (N_4017,N_3889,N_3944);
xnor U4018 (N_4018,N_3905,N_3968);
nor U4019 (N_4019,N_3862,N_3866);
xnor U4020 (N_4020,N_3803,N_3854);
xnor U4021 (N_4021,N_3843,N_3921);
xor U4022 (N_4022,N_3846,N_3865);
and U4023 (N_4023,N_3856,N_3895);
or U4024 (N_4024,N_3939,N_3976);
xnor U4025 (N_4025,N_3918,N_3897);
xor U4026 (N_4026,N_3806,N_3957);
or U4027 (N_4027,N_3901,N_3948);
and U4028 (N_4028,N_3951,N_3910);
or U4029 (N_4029,N_3855,N_3947);
xor U4030 (N_4030,N_3977,N_3880);
xnor U4031 (N_4031,N_3885,N_3835);
or U4032 (N_4032,N_3945,N_3881);
nor U4033 (N_4033,N_3999,N_3886);
or U4034 (N_4034,N_3828,N_3816);
xnor U4035 (N_4035,N_3848,N_3879);
nor U4036 (N_4036,N_3974,N_3810);
nor U4037 (N_4037,N_3840,N_3941);
xnor U4038 (N_4038,N_3814,N_3891);
nand U4039 (N_4039,N_3959,N_3946);
xnor U4040 (N_4040,N_3938,N_3887);
and U4041 (N_4041,N_3961,N_3831);
nand U4042 (N_4042,N_3847,N_3917);
nand U4043 (N_4043,N_3943,N_3861);
nand U4044 (N_4044,N_3820,N_3811);
and U4045 (N_4045,N_3922,N_3844);
nor U4046 (N_4046,N_3965,N_3937);
and U4047 (N_4047,N_3911,N_3884);
and U4048 (N_4048,N_3823,N_3869);
xor U4049 (N_4049,N_3892,N_3975);
and U4050 (N_4050,N_3893,N_3912);
nand U4051 (N_4051,N_3994,N_3899);
or U4052 (N_4052,N_3940,N_3863);
and U4053 (N_4053,N_3830,N_3845);
and U4054 (N_4054,N_3980,N_3859);
xnor U4055 (N_4055,N_3819,N_3876);
nand U4056 (N_4056,N_3930,N_3995);
nor U4057 (N_4057,N_3805,N_3981);
and U4058 (N_4058,N_3839,N_3966);
nor U4059 (N_4059,N_3984,N_3953);
xnor U4060 (N_4060,N_3920,N_3851);
or U4061 (N_4061,N_3964,N_3990);
nand U4062 (N_4062,N_3952,N_3907);
xor U4063 (N_4063,N_3928,N_3898);
nor U4064 (N_4064,N_3935,N_3860);
xor U4065 (N_4065,N_3870,N_3809);
xor U4066 (N_4066,N_3852,N_3933);
and U4067 (N_4067,N_3919,N_3890);
nor U4068 (N_4068,N_3996,N_3858);
and U4069 (N_4069,N_3978,N_3979);
or U4070 (N_4070,N_3888,N_3896);
nor U4071 (N_4071,N_3801,N_3827);
or U4072 (N_4072,N_3967,N_3817);
and U4073 (N_4073,N_3988,N_3829);
and U4074 (N_4074,N_3985,N_3997);
nand U4075 (N_4075,N_3836,N_3991);
xnor U4076 (N_4076,N_3818,N_3813);
or U4077 (N_4077,N_3821,N_3894);
and U4078 (N_4078,N_3983,N_3900);
nor U4079 (N_4079,N_3955,N_3909);
xor U4080 (N_4080,N_3842,N_3956);
xnor U4081 (N_4081,N_3837,N_3931);
or U4082 (N_4082,N_3925,N_3808);
and U4083 (N_4083,N_3902,N_3924);
nor U4084 (N_4084,N_3906,N_3972);
nor U4085 (N_4085,N_3825,N_3853);
xnor U4086 (N_4086,N_3934,N_3857);
xor U4087 (N_4087,N_3929,N_3804);
nor U4088 (N_4088,N_3916,N_3812);
nor U4089 (N_4089,N_3871,N_3882);
xor U4090 (N_4090,N_3963,N_3872);
and U4091 (N_4091,N_3942,N_3914);
nand U4092 (N_4092,N_3834,N_3950);
nor U4093 (N_4093,N_3903,N_3875);
nand U4094 (N_4094,N_3873,N_3883);
or U4095 (N_4095,N_3815,N_3998);
nand U4096 (N_4096,N_3833,N_3807);
xor U4097 (N_4097,N_3949,N_3877);
or U4098 (N_4098,N_3932,N_3936);
xor U4099 (N_4099,N_3915,N_3969);
xnor U4100 (N_4100,N_3838,N_3966);
or U4101 (N_4101,N_3992,N_3923);
nor U4102 (N_4102,N_3993,N_3847);
or U4103 (N_4103,N_3980,N_3985);
and U4104 (N_4104,N_3909,N_3835);
nand U4105 (N_4105,N_3944,N_3896);
nor U4106 (N_4106,N_3998,N_3848);
or U4107 (N_4107,N_3844,N_3905);
nor U4108 (N_4108,N_3859,N_3857);
nor U4109 (N_4109,N_3865,N_3830);
nand U4110 (N_4110,N_3918,N_3940);
nand U4111 (N_4111,N_3830,N_3925);
xor U4112 (N_4112,N_3894,N_3927);
nor U4113 (N_4113,N_3957,N_3907);
xor U4114 (N_4114,N_3960,N_3932);
or U4115 (N_4115,N_3928,N_3838);
and U4116 (N_4116,N_3833,N_3922);
or U4117 (N_4117,N_3987,N_3957);
nor U4118 (N_4118,N_3811,N_3822);
nor U4119 (N_4119,N_3860,N_3912);
and U4120 (N_4120,N_3997,N_3893);
or U4121 (N_4121,N_3904,N_3948);
or U4122 (N_4122,N_3944,N_3866);
or U4123 (N_4123,N_3995,N_3811);
xor U4124 (N_4124,N_3895,N_3992);
nand U4125 (N_4125,N_3907,N_3931);
and U4126 (N_4126,N_3993,N_3945);
nor U4127 (N_4127,N_3874,N_3934);
nor U4128 (N_4128,N_3873,N_3812);
nor U4129 (N_4129,N_3882,N_3984);
nand U4130 (N_4130,N_3897,N_3813);
nor U4131 (N_4131,N_3915,N_3940);
or U4132 (N_4132,N_3822,N_3912);
xor U4133 (N_4133,N_3918,N_3966);
nand U4134 (N_4134,N_3888,N_3905);
xnor U4135 (N_4135,N_3842,N_3821);
xor U4136 (N_4136,N_3855,N_3897);
or U4137 (N_4137,N_3904,N_3889);
and U4138 (N_4138,N_3804,N_3956);
xor U4139 (N_4139,N_3886,N_3923);
and U4140 (N_4140,N_3956,N_3948);
or U4141 (N_4141,N_3863,N_3907);
nand U4142 (N_4142,N_3966,N_3969);
nand U4143 (N_4143,N_3818,N_3872);
or U4144 (N_4144,N_3940,N_3824);
and U4145 (N_4145,N_3911,N_3928);
nor U4146 (N_4146,N_3851,N_3892);
xnor U4147 (N_4147,N_3870,N_3835);
xnor U4148 (N_4148,N_3999,N_3957);
xnor U4149 (N_4149,N_3804,N_3994);
nand U4150 (N_4150,N_3989,N_3991);
or U4151 (N_4151,N_3933,N_3968);
and U4152 (N_4152,N_3893,N_3892);
or U4153 (N_4153,N_3880,N_3854);
xor U4154 (N_4154,N_3860,N_3833);
xnor U4155 (N_4155,N_3909,N_3807);
or U4156 (N_4156,N_3900,N_3998);
nand U4157 (N_4157,N_3976,N_3943);
nor U4158 (N_4158,N_3888,N_3910);
and U4159 (N_4159,N_3978,N_3886);
xor U4160 (N_4160,N_3981,N_3962);
or U4161 (N_4161,N_3897,N_3965);
xnor U4162 (N_4162,N_3825,N_3855);
nand U4163 (N_4163,N_3996,N_3926);
or U4164 (N_4164,N_3867,N_3855);
xor U4165 (N_4165,N_3942,N_3848);
or U4166 (N_4166,N_3840,N_3935);
or U4167 (N_4167,N_3819,N_3868);
nor U4168 (N_4168,N_3850,N_3883);
nor U4169 (N_4169,N_3936,N_3858);
xor U4170 (N_4170,N_3918,N_3852);
xor U4171 (N_4171,N_3856,N_3989);
and U4172 (N_4172,N_3987,N_3999);
nand U4173 (N_4173,N_3907,N_3990);
or U4174 (N_4174,N_3879,N_3805);
nor U4175 (N_4175,N_3992,N_3914);
nor U4176 (N_4176,N_3801,N_3896);
or U4177 (N_4177,N_3861,N_3995);
xnor U4178 (N_4178,N_3908,N_3828);
nor U4179 (N_4179,N_3946,N_3930);
or U4180 (N_4180,N_3922,N_3868);
and U4181 (N_4181,N_3836,N_3825);
and U4182 (N_4182,N_3954,N_3854);
xor U4183 (N_4183,N_3935,N_3934);
nand U4184 (N_4184,N_3839,N_3897);
or U4185 (N_4185,N_3922,N_3952);
nor U4186 (N_4186,N_3810,N_3925);
or U4187 (N_4187,N_3997,N_3891);
and U4188 (N_4188,N_3869,N_3842);
xnor U4189 (N_4189,N_3989,N_3844);
nor U4190 (N_4190,N_3875,N_3801);
or U4191 (N_4191,N_3803,N_3936);
nand U4192 (N_4192,N_3885,N_3899);
nor U4193 (N_4193,N_3806,N_3889);
nor U4194 (N_4194,N_3960,N_3938);
nor U4195 (N_4195,N_3850,N_3897);
xnor U4196 (N_4196,N_3804,N_3937);
nand U4197 (N_4197,N_3950,N_3805);
or U4198 (N_4198,N_3824,N_3881);
xor U4199 (N_4199,N_3988,N_3910);
or U4200 (N_4200,N_4113,N_4009);
nand U4201 (N_4201,N_4086,N_4064);
and U4202 (N_4202,N_4198,N_4131);
nor U4203 (N_4203,N_4114,N_4096);
and U4204 (N_4204,N_4069,N_4022);
or U4205 (N_4205,N_4167,N_4088);
or U4206 (N_4206,N_4179,N_4141);
nor U4207 (N_4207,N_4162,N_4121);
or U4208 (N_4208,N_4102,N_4075);
xor U4209 (N_4209,N_4187,N_4100);
or U4210 (N_4210,N_4054,N_4067);
or U4211 (N_4211,N_4028,N_4109);
nor U4212 (N_4212,N_4148,N_4106);
nand U4213 (N_4213,N_4012,N_4010);
nand U4214 (N_4214,N_4043,N_4095);
xnor U4215 (N_4215,N_4154,N_4050);
nand U4216 (N_4216,N_4134,N_4058);
xor U4217 (N_4217,N_4180,N_4116);
nand U4218 (N_4218,N_4195,N_4140);
or U4219 (N_4219,N_4017,N_4165);
and U4220 (N_4220,N_4079,N_4078);
nor U4221 (N_4221,N_4184,N_4025);
and U4222 (N_4222,N_4164,N_4083);
nor U4223 (N_4223,N_4194,N_4048);
or U4224 (N_4224,N_4062,N_4019);
nor U4225 (N_4225,N_4097,N_4144);
and U4226 (N_4226,N_4125,N_4130);
nor U4227 (N_4227,N_4119,N_4132);
nand U4228 (N_4228,N_4163,N_4059);
nand U4229 (N_4229,N_4147,N_4128);
xor U4230 (N_4230,N_4020,N_4183);
nor U4231 (N_4231,N_4016,N_4173);
nand U4232 (N_4232,N_4138,N_4094);
nand U4233 (N_4233,N_4197,N_4133);
nand U4234 (N_4234,N_4135,N_4136);
or U4235 (N_4235,N_4011,N_4101);
or U4236 (N_4236,N_4000,N_4002);
and U4237 (N_4237,N_4199,N_4107);
nor U4238 (N_4238,N_4030,N_4171);
nor U4239 (N_4239,N_4077,N_4111);
and U4240 (N_4240,N_4076,N_4027);
nor U4241 (N_4241,N_4072,N_4026);
xor U4242 (N_4242,N_4152,N_4192);
nand U4243 (N_4243,N_4168,N_4150);
xor U4244 (N_4244,N_4196,N_4155);
nand U4245 (N_4245,N_4029,N_4018);
xnor U4246 (N_4246,N_4008,N_4166);
and U4247 (N_4247,N_4142,N_4047);
xnor U4248 (N_4248,N_4099,N_4188);
nor U4249 (N_4249,N_4161,N_4001);
and U4250 (N_4250,N_4031,N_4172);
or U4251 (N_4251,N_4104,N_4151);
xor U4252 (N_4252,N_4159,N_4080);
nand U4253 (N_4253,N_4024,N_4092);
and U4254 (N_4254,N_4063,N_4071);
xor U4255 (N_4255,N_4110,N_4093);
and U4256 (N_4256,N_4182,N_4089);
nor U4257 (N_4257,N_4117,N_4035);
and U4258 (N_4258,N_4174,N_4156);
nor U4259 (N_4259,N_4021,N_4177);
nand U4260 (N_4260,N_4045,N_4065);
nand U4261 (N_4261,N_4003,N_4189);
and U4262 (N_4262,N_4023,N_4040);
nand U4263 (N_4263,N_4175,N_4053);
or U4264 (N_4264,N_4032,N_4044);
nor U4265 (N_4265,N_4084,N_4123);
or U4266 (N_4266,N_4005,N_4073);
and U4267 (N_4267,N_4074,N_4015);
nand U4268 (N_4268,N_4052,N_4181);
xnor U4269 (N_4269,N_4042,N_4137);
nor U4270 (N_4270,N_4046,N_4120);
or U4271 (N_4271,N_4057,N_4124);
nor U4272 (N_4272,N_4039,N_4033);
nand U4273 (N_4273,N_4066,N_4146);
xnor U4274 (N_4274,N_4129,N_4157);
nor U4275 (N_4275,N_4176,N_4169);
or U4276 (N_4276,N_4036,N_4160);
nand U4277 (N_4277,N_4127,N_4186);
or U4278 (N_4278,N_4105,N_4178);
xor U4279 (N_4279,N_4049,N_4185);
nand U4280 (N_4280,N_4004,N_4122);
and U4281 (N_4281,N_4149,N_4014);
and U4282 (N_4282,N_4006,N_4068);
xnor U4283 (N_4283,N_4153,N_4038);
and U4284 (N_4284,N_4118,N_4158);
nor U4285 (N_4285,N_4037,N_4085);
or U4286 (N_4286,N_4108,N_4126);
and U4287 (N_4287,N_4081,N_4061);
and U4288 (N_4288,N_4193,N_4082);
and U4289 (N_4289,N_4055,N_4070);
nand U4290 (N_4290,N_4139,N_4115);
nand U4291 (N_4291,N_4034,N_4098);
or U4292 (N_4292,N_4103,N_4087);
nor U4293 (N_4293,N_4145,N_4112);
and U4294 (N_4294,N_4056,N_4191);
and U4295 (N_4295,N_4013,N_4091);
nand U4296 (N_4296,N_4170,N_4041);
nor U4297 (N_4297,N_4190,N_4051);
nand U4298 (N_4298,N_4143,N_4090);
xor U4299 (N_4299,N_4060,N_4007);
nor U4300 (N_4300,N_4079,N_4132);
nand U4301 (N_4301,N_4193,N_4138);
and U4302 (N_4302,N_4041,N_4089);
and U4303 (N_4303,N_4119,N_4156);
xnor U4304 (N_4304,N_4110,N_4148);
and U4305 (N_4305,N_4091,N_4064);
xnor U4306 (N_4306,N_4079,N_4140);
nor U4307 (N_4307,N_4181,N_4158);
and U4308 (N_4308,N_4047,N_4191);
xnor U4309 (N_4309,N_4088,N_4048);
xor U4310 (N_4310,N_4081,N_4186);
and U4311 (N_4311,N_4091,N_4156);
nand U4312 (N_4312,N_4154,N_4064);
xor U4313 (N_4313,N_4047,N_4192);
and U4314 (N_4314,N_4107,N_4034);
xor U4315 (N_4315,N_4020,N_4072);
and U4316 (N_4316,N_4025,N_4121);
nor U4317 (N_4317,N_4062,N_4126);
xnor U4318 (N_4318,N_4096,N_4134);
nor U4319 (N_4319,N_4144,N_4087);
nand U4320 (N_4320,N_4080,N_4082);
and U4321 (N_4321,N_4016,N_4103);
xnor U4322 (N_4322,N_4152,N_4036);
xor U4323 (N_4323,N_4112,N_4054);
and U4324 (N_4324,N_4085,N_4197);
xor U4325 (N_4325,N_4086,N_4134);
xor U4326 (N_4326,N_4145,N_4166);
and U4327 (N_4327,N_4022,N_4048);
and U4328 (N_4328,N_4019,N_4129);
xor U4329 (N_4329,N_4170,N_4198);
nand U4330 (N_4330,N_4124,N_4068);
or U4331 (N_4331,N_4003,N_4072);
xnor U4332 (N_4332,N_4080,N_4075);
or U4333 (N_4333,N_4178,N_4146);
and U4334 (N_4334,N_4120,N_4165);
or U4335 (N_4335,N_4172,N_4127);
xnor U4336 (N_4336,N_4006,N_4041);
or U4337 (N_4337,N_4096,N_4079);
nor U4338 (N_4338,N_4098,N_4045);
xnor U4339 (N_4339,N_4064,N_4161);
nand U4340 (N_4340,N_4031,N_4029);
xor U4341 (N_4341,N_4066,N_4009);
nor U4342 (N_4342,N_4004,N_4102);
or U4343 (N_4343,N_4195,N_4177);
xnor U4344 (N_4344,N_4089,N_4070);
and U4345 (N_4345,N_4075,N_4104);
nor U4346 (N_4346,N_4156,N_4092);
nor U4347 (N_4347,N_4179,N_4019);
or U4348 (N_4348,N_4088,N_4116);
or U4349 (N_4349,N_4008,N_4093);
nor U4350 (N_4350,N_4017,N_4015);
nor U4351 (N_4351,N_4006,N_4145);
or U4352 (N_4352,N_4060,N_4132);
xor U4353 (N_4353,N_4081,N_4184);
and U4354 (N_4354,N_4174,N_4029);
xor U4355 (N_4355,N_4073,N_4166);
or U4356 (N_4356,N_4080,N_4049);
nor U4357 (N_4357,N_4180,N_4163);
xnor U4358 (N_4358,N_4031,N_4019);
and U4359 (N_4359,N_4077,N_4105);
xor U4360 (N_4360,N_4155,N_4173);
nand U4361 (N_4361,N_4051,N_4072);
nand U4362 (N_4362,N_4177,N_4160);
and U4363 (N_4363,N_4016,N_4006);
xor U4364 (N_4364,N_4199,N_4026);
nand U4365 (N_4365,N_4087,N_4024);
xor U4366 (N_4366,N_4043,N_4157);
nor U4367 (N_4367,N_4117,N_4134);
xor U4368 (N_4368,N_4120,N_4071);
or U4369 (N_4369,N_4019,N_4053);
or U4370 (N_4370,N_4001,N_4170);
nand U4371 (N_4371,N_4048,N_4043);
nor U4372 (N_4372,N_4161,N_4027);
and U4373 (N_4373,N_4041,N_4175);
xnor U4374 (N_4374,N_4169,N_4029);
nor U4375 (N_4375,N_4080,N_4004);
nand U4376 (N_4376,N_4019,N_4121);
nand U4377 (N_4377,N_4036,N_4004);
xor U4378 (N_4378,N_4152,N_4143);
xor U4379 (N_4379,N_4058,N_4082);
and U4380 (N_4380,N_4012,N_4136);
xor U4381 (N_4381,N_4191,N_4156);
or U4382 (N_4382,N_4064,N_4173);
nand U4383 (N_4383,N_4141,N_4026);
xnor U4384 (N_4384,N_4160,N_4010);
and U4385 (N_4385,N_4140,N_4017);
xnor U4386 (N_4386,N_4183,N_4133);
and U4387 (N_4387,N_4024,N_4022);
or U4388 (N_4388,N_4006,N_4030);
nand U4389 (N_4389,N_4078,N_4075);
or U4390 (N_4390,N_4053,N_4024);
nand U4391 (N_4391,N_4085,N_4186);
or U4392 (N_4392,N_4057,N_4197);
nand U4393 (N_4393,N_4087,N_4005);
and U4394 (N_4394,N_4002,N_4059);
nor U4395 (N_4395,N_4010,N_4075);
and U4396 (N_4396,N_4057,N_4110);
nor U4397 (N_4397,N_4075,N_4107);
xnor U4398 (N_4398,N_4034,N_4009);
nor U4399 (N_4399,N_4174,N_4034);
xor U4400 (N_4400,N_4300,N_4271);
xnor U4401 (N_4401,N_4284,N_4324);
nand U4402 (N_4402,N_4399,N_4304);
nor U4403 (N_4403,N_4242,N_4306);
nor U4404 (N_4404,N_4236,N_4382);
nand U4405 (N_4405,N_4351,N_4257);
or U4406 (N_4406,N_4394,N_4252);
and U4407 (N_4407,N_4265,N_4230);
xor U4408 (N_4408,N_4392,N_4280);
nor U4409 (N_4409,N_4332,N_4371);
or U4410 (N_4410,N_4218,N_4295);
nand U4411 (N_4411,N_4212,N_4383);
nor U4412 (N_4412,N_4339,N_4363);
and U4413 (N_4413,N_4261,N_4210);
nand U4414 (N_4414,N_4299,N_4322);
nand U4415 (N_4415,N_4375,N_4369);
nand U4416 (N_4416,N_4333,N_4268);
or U4417 (N_4417,N_4227,N_4287);
or U4418 (N_4418,N_4229,N_4311);
nor U4419 (N_4419,N_4329,N_4398);
and U4420 (N_4420,N_4281,N_4319);
nand U4421 (N_4421,N_4272,N_4232);
nand U4422 (N_4422,N_4244,N_4397);
and U4423 (N_4423,N_4296,N_4207);
nand U4424 (N_4424,N_4327,N_4221);
nand U4425 (N_4425,N_4213,N_4205);
xor U4426 (N_4426,N_4288,N_4204);
xor U4427 (N_4427,N_4305,N_4285);
xor U4428 (N_4428,N_4346,N_4364);
xor U4429 (N_4429,N_4386,N_4235);
and U4430 (N_4430,N_4289,N_4331);
and U4431 (N_4431,N_4269,N_4313);
and U4432 (N_4432,N_4368,N_4350);
and U4433 (N_4433,N_4262,N_4309);
and U4434 (N_4434,N_4385,N_4275);
and U4435 (N_4435,N_4325,N_4373);
or U4436 (N_4436,N_4381,N_4348);
xnor U4437 (N_4437,N_4323,N_4302);
nor U4438 (N_4438,N_4372,N_4396);
nand U4439 (N_4439,N_4282,N_4370);
and U4440 (N_4440,N_4249,N_4314);
nand U4441 (N_4441,N_4395,N_4317);
and U4442 (N_4442,N_4316,N_4365);
nor U4443 (N_4443,N_4209,N_4225);
nand U4444 (N_4444,N_4224,N_4201);
or U4445 (N_4445,N_4307,N_4239);
nand U4446 (N_4446,N_4358,N_4376);
and U4447 (N_4447,N_4220,N_4200);
xor U4448 (N_4448,N_4214,N_4303);
nand U4449 (N_4449,N_4379,N_4208);
nor U4450 (N_4450,N_4255,N_4276);
nand U4451 (N_4451,N_4270,N_4367);
or U4452 (N_4452,N_4354,N_4222);
nor U4453 (N_4453,N_4263,N_4312);
or U4454 (N_4454,N_4228,N_4256);
and U4455 (N_4455,N_4231,N_4211);
nor U4456 (N_4456,N_4247,N_4347);
and U4457 (N_4457,N_4328,N_4384);
and U4458 (N_4458,N_4349,N_4273);
and U4459 (N_4459,N_4337,N_4240);
xnor U4460 (N_4460,N_4342,N_4253);
and U4461 (N_4461,N_4217,N_4290);
nand U4462 (N_4462,N_4389,N_4356);
or U4463 (N_4463,N_4391,N_4245);
and U4464 (N_4464,N_4219,N_4248);
xnor U4465 (N_4465,N_4310,N_4292);
and U4466 (N_4466,N_4359,N_4293);
or U4467 (N_4467,N_4226,N_4237);
nor U4468 (N_4468,N_4298,N_4340);
nand U4469 (N_4469,N_4266,N_4378);
or U4470 (N_4470,N_4320,N_4341);
xor U4471 (N_4471,N_4390,N_4335);
nor U4472 (N_4472,N_4377,N_4279);
and U4473 (N_4473,N_4286,N_4360);
xor U4474 (N_4474,N_4362,N_4274);
nor U4475 (N_4475,N_4361,N_4336);
xnor U4476 (N_4476,N_4393,N_4259);
nand U4477 (N_4477,N_4366,N_4260);
nor U4478 (N_4478,N_4294,N_4326);
nor U4479 (N_4479,N_4387,N_4315);
and U4480 (N_4480,N_4278,N_4250);
and U4481 (N_4481,N_4216,N_4374);
nor U4482 (N_4482,N_4352,N_4234);
and U4483 (N_4483,N_4241,N_4344);
nand U4484 (N_4484,N_4258,N_4283);
nor U4485 (N_4485,N_4353,N_4233);
xor U4486 (N_4486,N_4238,N_4264);
nand U4487 (N_4487,N_4206,N_4318);
or U4488 (N_4488,N_4357,N_4246);
nor U4489 (N_4489,N_4308,N_4345);
xnor U4490 (N_4490,N_4251,N_4223);
and U4491 (N_4491,N_4321,N_4334);
nand U4492 (N_4492,N_4203,N_4380);
or U4493 (N_4493,N_4343,N_4338);
nand U4494 (N_4494,N_4297,N_4254);
or U4495 (N_4495,N_4243,N_4330);
and U4496 (N_4496,N_4267,N_4301);
nor U4497 (N_4497,N_4388,N_4291);
nor U4498 (N_4498,N_4202,N_4215);
and U4499 (N_4499,N_4355,N_4277);
nand U4500 (N_4500,N_4319,N_4228);
or U4501 (N_4501,N_4201,N_4222);
nand U4502 (N_4502,N_4307,N_4305);
and U4503 (N_4503,N_4323,N_4367);
or U4504 (N_4504,N_4218,N_4325);
nand U4505 (N_4505,N_4270,N_4336);
and U4506 (N_4506,N_4231,N_4318);
nor U4507 (N_4507,N_4224,N_4223);
nor U4508 (N_4508,N_4367,N_4210);
nand U4509 (N_4509,N_4331,N_4275);
nand U4510 (N_4510,N_4213,N_4328);
xnor U4511 (N_4511,N_4332,N_4330);
nand U4512 (N_4512,N_4207,N_4276);
nand U4513 (N_4513,N_4287,N_4373);
nor U4514 (N_4514,N_4266,N_4308);
nor U4515 (N_4515,N_4379,N_4343);
and U4516 (N_4516,N_4346,N_4322);
and U4517 (N_4517,N_4399,N_4301);
or U4518 (N_4518,N_4310,N_4363);
nand U4519 (N_4519,N_4284,N_4396);
xor U4520 (N_4520,N_4379,N_4235);
or U4521 (N_4521,N_4374,N_4316);
xor U4522 (N_4522,N_4234,N_4280);
xnor U4523 (N_4523,N_4202,N_4351);
and U4524 (N_4524,N_4306,N_4261);
or U4525 (N_4525,N_4317,N_4332);
nand U4526 (N_4526,N_4342,N_4373);
xor U4527 (N_4527,N_4397,N_4219);
xnor U4528 (N_4528,N_4277,N_4309);
nand U4529 (N_4529,N_4367,N_4331);
and U4530 (N_4530,N_4373,N_4314);
nand U4531 (N_4531,N_4374,N_4390);
or U4532 (N_4532,N_4221,N_4369);
nor U4533 (N_4533,N_4394,N_4345);
nor U4534 (N_4534,N_4384,N_4294);
and U4535 (N_4535,N_4338,N_4312);
nand U4536 (N_4536,N_4366,N_4321);
nor U4537 (N_4537,N_4335,N_4273);
and U4538 (N_4538,N_4338,N_4365);
nand U4539 (N_4539,N_4286,N_4340);
xor U4540 (N_4540,N_4382,N_4352);
nor U4541 (N_4541,N_4385,N_4298);
and U4542 (N_4542,N_4226,N_4275);
xor U4543 (N_4543,N_4305,N_4312);
nand U4544 (N_4544,N_4397,N_4285);
or U4545 (N_4545,N_4241,N_4397);
nand U4546 (N_4546,N_4283,N_4250);
nand U4547 (N_4547,N_4367,N_4274);
nor U4548 (N_4548,N_4228,N_4234);
nand U4549 (N_4549,N_4335,N_4394);
xor U4550 (N_4550,N_4308,N_4314);
xnor U4551 (N_4551,N_4271,N_4350);
or U4552 (N_4552,N_4219,N_4238);
xor U4553 (N_4553,N_4308,N_4371);
nand U4554 (N_4554,N_4251,N_4220);
or U4555 (N_4555,N_4205,N_4341);
nand U4556 (N_4556,N_4205,N_4370);
or U4557 (N_4557,N_4269,N_4213);
nand U4558 (N_4558,N_4289,N_4376);
xnor U4559 (N_4559,N_4227,N_4250);
and U4560 (N_4560,N_4292,N_4296);
nand U4561 (N_4561,N_4364,N_4302);
and U4562 (N_4562,N_4277,N_4282);
and U4563 (N_4563,N_4387,N_4302);
nor U4564 (N_4564,N_4271,N_4260);
nand U4565 (N_4565,N_4238,N_4348);
and U4566 (N_4566,N_4379,N_4255);
nand U4567 (N_4567,N_4228,N_4238);
xnor U4568 (N_4568,N_4305,N_4371);
or U4569 (N_4569,N_4309,N_4256);
xor U4570 (N_4570,N_4218,N_4274);
and U4571 (N_4571,N_4372,N_4366);
or U4572 (N_4572,N_4297,N_4281);
nor U4573 (N_4573,N_4297,N_4290);
xor U4574 (N_4574,N_4334,N_4209);
and U4575 (N_4575,N_4201,N_4308);
nor U4576 (N_4576,N_4325,N_4277);
nor U4577 (N_4577,N_4398,N_4226);
or U4578 (N_4578,N_4235,N_4323);
xnor U4579 (N_4579,N_4370,N_4393);
xnor U4580 (N_4580,N_4366,N_4318);
and U4581 (N_4581,N_4337,N_4328);
nand U4582 (N_4582,N_4248,N_4265);
xnor U4583 (N_4583,N_4348,N_4227);
nand U4584 (N_4584,N_4365,N_4382);
xnor U4585 (N_4585,N_4203,N_4286);
or U4586 (N_4586,N_4314,N_4239);
nor U4587 (N_4587,N_4330,N_4338);
or U4588 (N_4588,N_4300,N_4285);
nand U4589 (N_4589,N_4227,N_4217);
xnor U4590 (N_4590,N_4351,N_4221);
nand U4591 (N_4591,N_4299,N_4395);
and U4592 (N_4592,N_4210,N_4357);
nand U4593 (N_4593,N_4302,N_4391);
nor U4594 (N_4594,N_4309,N_4328);
nand U4595 (N_4595,N_4204,N_4203);
nor U4596 (N_4596,N_4215,N_4325);
and U4597 (N_4597,N_4217,N_4226);
or U4598 (N_4598,N_4217,N_4334);
and U4599 (N_4599,N_4294,N_4305);
xnor U4600 (N_4600,N_4593,N_4594);
and U4601 (N_4601,N_4595,N_4529);
xnor U4602 (N_4602,N_4436,N_4586);
or U4603 (N_4603,N_4547,N_4518);
and U4604 (N_4604,N_4559,N_4445);
xor U4605 (N_4605,N_4455,N_4423);
and U4606 (N_4606,N_4499,N_4531);
nand U4607 (N_4607,N_4415,N_4427);
and U4608 (N_4608,N_4555,N_4466);
nand U4609 (N_4609,N_4503,N_4425);
xor U4610 (N_4610,N_4407,N_4442);
nand U4611 (N_4611,N_4494,N_4591);
nand U4612 (N_4612,N_4462,N_4465);
nand U4613 (N_4613,N_4471,N_4530);
or U4614 (N_4614,N_4554,N_4428);
xnor U4615 (N_4615,N_4482,N_4416);
or U4616 (N_4616,N_4438,N_4561);
xnor U4617 (N_4617,N_4583,N_4420);
xnor U4618 (N_4618,N_4504,N_4454);
nor U4619 (N_4619,N_4563,N_4562);
nor U4620 (N_4620,N_4448,N_4492);
nor U4621 (N_4621,N_4418,N_4549);
xnor U4622 (N_4622,N_4498,N_4433);
xnor U4623 (N_4623,N_4412,N_4553);
xor U4624 (N_4624,N_4525,N_4539);
and U4625 (N_4625,N_4488,N_4506);
nand U4626 (N_4626,N_4527,N_4575);
and U4627 (N_4627,N_4495,N_4443);
nor U4628 (N_4628,N_4572,N_4489);
and U4629 (N_4629,N_4523,N_4487);
xor U4630 (N_4630,N_4459,N_4484);
or U4631 (N_4631,N_4543,N_4551);
nor U4632 (N_4632,N_4474,N_4578);
nand U4633 (N_4633,N_4486,N_4431);
nand U4634 (N_4634,N_4509,N_4432);
nor U4635 (N_4635,N_4521,N_4515);
xnor U4636 (N_4636,N_4596,N_4537);
nand U4637 (N_4637,N_4571,N_4582);
xnor U4638 (N_4638,N_4452,N_4491);
nor U4639 (N_4639,N_4426,N_4403);
nor U4640 (N_4640,N_4532,N_4446);
nor U4641 (N_4641,N_4456,N_4508);
or U4642 (N_4642,N_4413,N_4450);
and U4643 (N_4643,N_4472,N_4469);
xnor U4644 (N_4644,N_4473,N_4587);
nor U4645 (N_4645,N_4577,N_4550);
nor U4646 (N_4646,N_4470,N_4584);
and U4647 (N_4647,N_4542,N_4599);
nand U4648 (N_4648,N_4510,N_4479);
and U4649 (N_4649,N_4406,N_4517);
nor U4650 (N_4650,N_4513,N_4500);
xnor U4651 (N_4651,N_4457,N_4405);
and U4652 (N_4652,N_4449,N_4585);
nand U4653 (N_4653,N_4434,N_4514);
nor U4654 (N_4654,N_4533,N_4460);
or U4655 (N_4655,N_4566,N_4520);
xnor U4656 (N_4656,N_4435,N_4580);
nor U4657 (N_4657,N_4524,N_4481);
xnor U4658 (N_4658,N_4589,N_4541);
or U4659 (N_4659,N_4536,N_4497);
or U4660 (N_4660,N_4534,N_4592);
or U4661 (N_4661,N_4598,N_4429);
xor U4662 (N_4662,N_4441,N_4409);
nand U4663 (N_4663,N_4496,N_4540);
or U4664 (N_4664,N_4400,N_4421);
xor U4665 (N_4665,N_4467,N_4461);
and U4666 (N_4666,N_4480,N_4573);
nand U4667 (N_4667,N_4401,N_4437);
nor U4668 (N_4668,N_4478,N_4502);
nor U4669 (N_4669,N_4451,N_4546);
or U4670 (N_4670,N_4576,N_4483);
xnor U4671 (N_4671,N_4557,N_4463);
and U4672 (N_4672,N_4526,N_4570);
xor U4673 (N_4673,N_4430,N_4522);
and U4674 (N_4674,N_4574,N_4404);
and U4675 (N_4675,N_4516,N_4468);
nor U4676 (N_4676,N_4569,N_4597);
or U4677 (N_4677,N_4464,N_4447);
and U4678 (N_4678,N_4519,N_4558);
nor U4679 (N_4679,N_4444,N_4439);
and U4680 (N_4680,N_4567,N_4579);
or U4681 (N_4681,N_4424,N_4458);
nor U4682 (N_4682,N_4417,N_4511);
nor U4683 (N_4683,N_4501,N_4485);
xnor U4684 (N_4684,N_4419,N_4453);
nor U4685 (N_4685,N_4535,N_4490);
xor U4686 (N_4686,N_4560,N_4414);
or U4687 (N_4687,N_4410,N_4568);
or U4688 (N_4688,N_4505,N_4588);
nand U4689 (N_4689,N_4545,N_4564);
xnor U4690 (N_4690,N_4411,N_4422);
nand U4691 (N_4691,N_4512,N_4408);
nand U4692 (N_4692,N_4477,N_4440);
or U4693 (N_4693,N_4493,N_4402);
nand U4694 (N_4694,N_4590,N_4475);
nand U4695 (N_4695,N_4581,N_4476);
nor U4696 (N_4696,N_4565,N_4556);
nor U4697 (N_4697,N_4507,N_4528);
and U4698 (N_4698,N_4552,N_4548);
and U4699 (N_4699,N_4544,N_4538);
and U4700 (N_4700,N_4556,N_4580);
nor U4701 (N_4701,N_4473,N_4531);
nor U4702 (N_4702,N_4464,N_4565);
nor U4703 (N_4703,N_4498,N_4503);
xor U4704 (N_4704,N_4540,N_4471);
xnor U4705 (N_4705,N_4527,N_4481);
xor U4706 (N_4706,N_4506,N_4476);
xnor U4707 (N_4707,N_4405,N_4428);
and U4708 (N_4708,N_4516,N_4449);
nand U4709 (N_4709,N_4556,N_4515);
nor U4710 (N_4710,N_4449,N_4533);
nor U4711 (N_4711,N_4419,N_4443);
nand U4712 (N_4712,N_4539,N_4582);
nor U4713 (N_4713,N_4546,N_4419);
xor U4714 (N_4714,N_4468,N_4414);
nand U4715 (N_4715,N_4545,N_4425);
and U4716 (N_4716,N_4478,N_4457);
and U4717 (N_4717,N_4407,N_4481);
nand U4718 (N_4718,N_4496,N_4441);
and U4719 (N_4719,N_4498,N_4427);
or U4720 (N_4720,N_4540,N_4421);
xnor U4721 (N_4721,N_4451,N_4403);
nor U4722 (N_4722,N_4445,N_4578);
or U4723 (N_4723,N_4407,N_4428);
or U4724 (N_4724,N_4431,N_4528);
or U4725 (N_4725,N_4472,N_4487);
nor U4726 (N_4726,N_4582,N_4497);
nor U4727 (N_4727,N_4484,N_4450);
nand U4728 (N_4728,N_4559,N_4400);
xor U4729 (N_4729,N_4463,N_4411);
xnor U4730 (N_4730,N_4565,N_4450);
or U4731 (N_4731,N_4592,N_4415);
nor U4732 (N_4732,N_4473,N_4541);
nand U4733 (N_4733,N_4526,N_4482);
nand U4734 (N_4734,N_4567,N_4499);
or U4735 (N_4735,N_4573,N_4533);
xor U4736 (N_4736,N_4507,N_4446);
or U4737 (N_4737,N_4449,N_4577);
xor U4738 (N_4738,N_4504,N_4470);
nor U4739 (N_4739,N_4582,N_4489);
nor U4740 (N_4740,N_4534,N_4510);
or U4741 (N_4741,N_4562,N_4467);
or U4742 (N_4742,N_4587,N_4402);
xnor U4743 (N_4743,N_4493,N_4443);
or U4744 (N_4744,N_4464,N_4510);
or U4745 (N_4745,N_4455,N_4595);
or U4746 (N_4746,N_4467,N_4482);
and U4747 (N_4747,N_4422,N_4445);
xor U4748 (N_4748,N_4449,N_4590);
or U4749 (N_4749,N_4438,N_4579);
or U4750 (N_4750,N_4479,N_4468);
or U4751 (N_4751,N_4528,N_4436);
nor U4752 (N_4752,N_4533,N_4446);
or U4753 (N_4753,N_4426,N_4536);
and U4754 (N_4754,N_4429,N_4483);
nor U4755 (N_4755,N_4451,N_4594);
xnor U4756 (N_4756,N_4489,N_4451);
xor U4757 (N_4757,N_4424,N_4460);
nor U4758 (N_4758,N_4586,N_4536);
nor U4759 (N_4759,N_4557,N_4403);
nor U4760 (N_4760,N_4433,N_4461);
nor U4761 (N_4761,N_4469,N_4585);
nand U4762 (N_4762,N_4501,N_4527);
or U4763 (N_4763,N_4543,N_4594);
xnor U4764 (N_4764,N_4543,N_4563);
nor U4765 (N_4765,N_4424,N_4475);
xnor U4766 (N_4766,N_4500,N_4557);
nor U4767 (N_4767,N_4425,N_4434);
or U4768 (N_4768,N_4406,N_4528);
xor U4769 (N_4769,N_4587,N_4429);
xnor U4770 (N_4770,N_4419,N_4470);
nand U4771 (N_4771,N_4512,N_4543);
nand U4772 (N_4772,N_4550,N_4423);
nor U4773 (N_4773,N_4540,N_4508);
xnor U4774 (N_4774,N_4508,N_4564);
or U4775 (N_4775,N_4529,N_4406);
or U4776 (N_4776,N_4464,N_4419);
or U4777 (N_4777,N_4414,N_4476);
xnor U4778 (N_4778,N_4425,N_4486);
xnor U4779 (N_4779,N_4461,N_4522);
nor U4780 (N_4780,N_4458,N_4403);
nor U4781 (N_4781,N_4508,N_4469);
and U4782 (N_4782,N_4498,N_4559);
nand U4783 (N_4783,N_4510,N_4474);
and U4784 (N_4784,N_4440,N_4501);
and U4785 (N_4785,N_4492,N_4465);
and U4786 (N_4786,N_4412,N_4470);
and U4787 (N_4787,N_4487,N_4437);
xor U4788 (N_4788,N_4419,N_4472);
nor U4789 (N_4789,N_4551,N_4415);
and U4790 (N_4790,N_4458,N_4527);
nand U4791 (N_4791,N_4401,N_4414);
nand U4792 (N_4792,N_4412,N_4527);
xor U4793 (N_4793,N_4532,N_4506);
xor U4794 (N_4794,N_4460,N_4481);
or U4795 (N_4795,N_4567,N_4478);
nand U4796 (N_4796,N_4581,N_4481);
and U4797 (N_4797,N_4574,N_4570);
or U4798 (N_4798,N_4585,N_4447);
nand U4799 (N_4799,N_4549,N_4461);
nand U4800 (N_4800,N_4720,N_4710);
nand U4801 (N_4801,N_4769,N_4636);
xnor U4802 (N_4802,N_4723,N_4740);
xnor U4803 (N_4803,N_4702,N_4748);
nand U4804 (N_4804,N_4680,N_4618);
or U4805 (N_4805,N_4716,N_4685);
or U4806 (N_4806,N_4608,N_4721);
nor U4807 (N_4807,N_4719,N_4777);
nor U4808 (N_4808,N_4639,N_4621);
xor U4809 (N_4809,N_4738,N_4665);
nor U4810 (N_4810,N_4656,N_4712);
and U4811 (N_4811,N_4610,N_4774);
nor U4812 (N_4812,N_4762,N_4708);
xnor U4813 (N_4813,N_4641,N_4638);
xnor U4814 (N_4814,N_4786,N_4755);
and U4815 (N_4815,N_4775,N_4739);
or U4816 (N_4816,N_4686,N_4632);
and U4817 (N_4817,N_4732,N_4707);
nand U4818 (N_4818,N_4790,N_4699);
or U4819 (N_4819,N_4772,N_4626);
nor U4820 (N_4820,N_4698,N_4795);
xnor U4821 (N_4821,N_4684,N_4747);
nor U4822 (N_4822,N_4696,N_4797);
xnor U4823 (N_4823,N_4767,N_4779);
nor U4824 (N_4824,N_4659,N_4788);
nand U4825 (N_4825,N_4727,N_4616);
nor U4826 (N_4826,N_4613,N_4657);
xor U4827 (N_4827,N_4751,N_4683);
or U4828 (N_4828,N_4736,N_4635);
xnor U4829 (N_4829,N_4681,N_4765);
xor U4830 (N_4830,N_4653,N_4624);
and U4831 (N_4831,N_4660,N_4749);
and U4832 (N_4832,N_4654,N_4674);
xnor U4833 (N_4833,N_4631,N_4630);
xnor U4834 (N_4834,N_4700,N_4644);
and U4835 (N_4835,N_4649,N_4766);
nor U4836 (N_4836,N_4643,N_4697);
and U4837 (N_4837,N_4612,N_4668);
and U4838 (N_4838,N_4776,N_4717);
or U4839 (N_4839,N_4715,N_4750);
or U4840 (N_4840,N_4648,N_4734);
nand U4841 (N_4841,N_4725,N_4675);
nand U4842 (N_4842,N_4693,N_4620);
nor U4843 (N_4843,N_4600,N_4672);
nor U4844 (N_4844,N_4763,N_4694);
nor U4845 (N_4845,N_4745,N_4780);
or U4846 (N_4846,N_4728,N_4652);
nor U4847 (N_4847,N_4718,N_4679);
xor U4848 (N_4848,N_4709,N_4733);
and U4849 (N_4849,N_4722,N_4617);
nor U4850 (N_4850,N_4677,N_4758);
and U4851 (N_4851,N_4705,N_4687);
nand U4852 (N_4852,N_4666,N_4604);
and U4853 (N_4853,N_4793,N_4601);
nand U4854 (N_4854,N_4798,N_4628);
and U4855 (N_4855,N_4744,N_4796);
or U4856 (N_4856,N_4682,N_4752);
nand U4857 (N_4857,N_4603,N_4671);
and U4858 (N_4858,N_4784,N_4609);
nand U4859 (N_4859,N_4678,N_4791);
nand U4860 (N_4860,N_4737,N_4670);
nor U4861 (N_4861,N_4690,N_4783);
or U4862 (N_4862,N_4622,N_4764);
nor U4863 (N_4863,N_4753,N_4730);
nor U4864 (N_4864,N_4781,N_4789);
and U4865 (N_4865,N_4640,N_4704);
nor U4866 (N_4866,N_4778,N_4787);
or U4867 (N_4867,N_4703,N_4714);
xor U4868 (N_4868,N_4757,N_4650);
and U4869 (N_4869,N_4602,N_4605);
or U4870 (N_4870,N_4689,N_4724);
or U4871 (N_4871,N_4646,N_4664);
and U4872 (N_4872,N_4760,N_4629);
nor U4873 (N_4873,N_4669,N_4691);
nand U4874 (N_4874,N_4773,N_4761);
xnor U4875 (N_4875,N_4688,N_4706);
or U4876 (N_4876,N_4729,N_4655);
xnor U4877 (N_4877,N_4771,N_4625);
xnor U4878 (N_4878,N_4637,N_4663);
nand U4879 (N_4879,N_4792,N_4759);
or U4880 (N_4880,N_4726,N_4627);
or U4881 (N_4881,N_4713,N_4799);
or U4882 (N_4882,N_4615,N_4754);
xnor U4883 (N_4883,N_4606,N_4619);
and U4884 (N_4884,N_4667,N_4651);
and U4885 (N_4885,N_4692,N_4614);
nor U4886 (N_4886,N_4611,N_4633);
nor U4887 (N_4887,N_4770,N_4642);
or U4888 (N_4888,N_4645,N_4746);
or U4889 (N_4889,N_4658,N_4768);
and U4890 (N_4890,N_4701,N_4662);
xnor U4891 (N_4891,N_4634,N_4756);
or U4892 (N_4892,N_4673,N_4741);
xnor U4893 (N_4893,N_4695,N_4647);
xor U4894 (N_4894,N_4623,N_4742);
nor U4895 (N_4895,N_4711,N_4731);
xor U4896 (N_4896,N_4676,N_4661);
or U4897 (N_4897,N_4607,N_4743);
or U4898 (N_4898,N_4735,N_4785);
nor U4899 (N_4899,N_4794,N_4782);
nand U4900 (N_4900,N_4653,N_4772);
nor U4901 (N_4901,N_4702,N_4695);
nor U4902 (N_4902,N_4632,N_4793);
nand U4903 (N_4903,N_4664,N_4713);
nand U4904 (N_4904,N_4678,N_4652);
xnor U4905 (N_4905,N_4637,N_4715);
nor U4906 (N_4906,N_4774,N_4777);
nor U4907 (N_4907,N_4623,N_4694);
or U4908 (N_4908,N_4771,N_4708);
nor U4909 (N_4909,N_4709,N_4669);
nor U4910 (N_4910,N_4770,N_4705);
xnor U4911 (N_4911,N_4697,N_4607);
nand U4912 (N_4912,N_4753,N_4703);
and U4913 (N_4913,N_4689,N_4615);
nor U4914 (N_4914,N_4674,N_4777);
xor U4915 (N_4915,N_4705,N_4742);
xnor U4916 (N_4916,N_4714,N_4691);
nand U4917 (N_4917,N_4763,N_4696);
nor U4918 (N_4918,N_4769,N_4605);
nand U4919 (N_4919,N_4693,N_4644);
or U4920 (N_4920,N_4775,N_4712);
xnor U4921 (N_4921,N_4637,N_4682);
nand U4922 (N_4922,N_4701,N_4669);
xnor U4923 (N_4923,N_4698,N_4738);
and U4924 (N_4924,N_4668,N_4642);
nor U4925 (N_4925,N_4614,N_4793);
xor U4926 (N_4926,N_4640,N_4619);
nand U4927 (N_4927,N_4773,N_4673);
or U4928 (N_4928,N_4659,N_4782);
or U4929 (N_4929,N_4711,N_4743);
nor U4930 (N_4930,N_4665,N_4716);
nand U4931 (N_4931,N_4766,N_4722);
or U4932 (N_4932,N_4733,N_4642);
or U4933 (N_4933,N_4655,N_4606);
nand U4934 (N_4934,N_4714,N_4740);
or U4935 (N_4935,N_4695,N_4699);
or U4936 (N_4936,N_4613,N_4781);
nand U4937 (N_4937,N_4645,N_4650);
nand U4938 (N_4938,N_4627,N_4623);
or U4939 (N_4939,N_4740,N_4777);
or U4940 (N_4940,N_4605,N_4693);
xnor U4941 (N_4941,N_4780,N_4778);
nand U4942 (N_4942,N_4675,N_4602);
or U4943 (N_4943,N_4670,N_4652);
and U4944 (N_4944,N_4633,N_4725);
nand U4945 (N_4945,N_4724,N_4720);
nand U4946 (N_4946,N_4731,N_4610);
or U4947 (N_4947,N_4770,N_4771);
xor U4948 (N_4948,N_4781,N_4675);
and U4949 (N_4949,N_4713,N_4706);
and U4950 (N_4950,N_4649,N_4693);
nor U4951 (N_4951,N_4679,N_4697);
or U4952 (N_4952,N_4712,N_4626);
and U4953 (N_4953,N_4753,N_4745);
or U4954 (N_4954,N_4606,N_4709);
nor U4955 (N_4955,N_4630,N_4710);
nand U4956 (N_4956,N_4602,N_4769);
xnor U4957 (N_4957,N_4611,N_4681);
or U4958 (N_4958,N_4711,N_4704);
or U4959 (N_4959,N_4764,N_4758);
nor U4960 (N_4960,N_4772,N_4727);
and U4961 (N_4961,N_4634,N_4708);
and U4962 (N_4962,N_4736,N_4651);
or U4963 (N_4963,N_4720,N_4749);
xor U4964 (N_4964,N_4693,N_4732);
nand U4965 (N_4965,N_4652,N_4751);
xor U4966 (N_4966,N_4760,N_4730);
nor U4967 (N_4967,N_4678,N_4611);
nor U4968 (N_4968,N_4719,N_4654);
nor U4969 (N_4969,N_4737,N_4607);
nand U4970 (N_4970,N_4633,N_4745);
and U4971 (N_4971,N_4601,N_4783);
nor U4972 (N_4972,N_4708,N_4743);
and U4973 (N_4973,N_4792,N_4634);
nor U4974 (N_4974,N_4636,N_4683);
xnor U4975 (N_4975,N_4733,N_4674);
and U4976 (N_4976,N_4703,N_4726);
and U4977 (N_4977,N_4602,N_4694);
and U4978 (N_4978,N_4604,N_4780);
xor U4979 (N_4979,N_4770,N_4692);
nand U4980 (N_4980,N_4749,N_4715);
nand U4981 (N_4981,N_4640,N_4691);
and U4982 (N_4982,N_4787,N_4713);
and U4983 (N_4983,N_4619,N_4699);
or U4984 (N_4984,N_4671,N_4750);
and U4985 (N_4985,N_4792,N_4693);
nand U4986 (N_4986,N_4753,N_4650);
nand U4987 (N_4987,N_4716,N_4654);
and U4988 (N_4988,N_4788,N_4784);
nand U4989 (N_4989,N_4706,N_4658);
or U4990 (N_4990,N_4681,N_4794);
and U4991 (N_4991,N_4677,N_4749);
and U4992 (N_4992,N_4606,N_4652);
and U4993 (N_4993,N_4684,N_4609);
and U4994 (N_4994,N_4798,N_4624);
or U4995 (N_4995,N_4759,N_4696);
and U4996 (N_4996,N_4658,N_4764);
nor U4997 (N_4997,N_4782,N_4709);
nand U4998 (N_4998,N_4731,N_4756);
and U4999 (N_4999,N_4697,N_4677);
and U5000 (N_5000,N_4990,N_4953);
and U5001 (N_5001,N_4995,N_4988);
xor U5002 (N_5002,N_4964,N_4820);
and U5003 (N_5003,N_4884,N_4965);
xor U5004 (N_5004,N_4868,N_4892);
xor U5005 (N_5005,N_4937,N_4998);
xnor U5006 (N_5006,N_4913,N_4922);
xnor U5007 (N_5007,N_4908,N_4911);
nor U5008 (N_5008,N_4959,N_4983);
and U5009 (N_5009,N_4840,N_4854);
nor U5010 (N_5010,N_4993,N_4873);
nor U5011 (N_5011,N_4980,N_4976);
nor U5012 (N_5012,N_4896,N_4888);
and U5013 (N_5013,N_4999,N_4800);
nor U5014 (N_5014,N_4935,N_4902);
xor U5015 (N_5015,N_4994,N_4914);
or U5016 (N_5016,N_4844,N_4871);
nor U5017 (N_5017,N_4987,N_4938);
xnor U5018 (N_5018,N_4872,N_4897);
and U5019 (N_5019,N_4809,N_4822);
or U5020 (N_5020,N_4931,N_4961);
nand U5021 (N_5021,N_4952,N_4958);
xor U5022 (N_5022,N_4962,N_4904);
xnor U5023 (N_5023,N_4936,N_4954);
and U5024 (N_5024,N_4816,N_4882);
xor U5025 (N_5025,N_4894,N_4975);
nor U5026 (N_5026,N_4857,N_4905);
and U5027 (N_5027,N_4806,N_4972);
nor U5028 (N_5028,N_4803,N_4869);
nand U5029 (N_5029,N_4891,N_4997);
nand U5030 (N_5030,N_4812,N_4824);
nand U5031 (N_5031,N_4819,N_4927);
and U5032 (N_5032,N_4890,N_4880);
and U5033 (N_5033,N_4862,N_4957);
and U5034 (N_5034,N_4917,N_4989);
or U5035 (N_5035,N_4855,N_4901);
or U5036 (N_5036,N_4867,N_4808);
nand U5037 (N_5037,N_4861,N_4838);
nand U5038 (N_5038,N_4996,N_4810);
or U5039 (N_5039,N_4841,N_4918);
nand U5040 (N_5040,N_4848,N_4837);
and U5041 (N_5041,N_4856,N_4977);
or U5042 (N_5042,N_4864,N_4924);
xnor U5043 (N_5043,N_4916,N_4992);
and U5044 (N_5044,N_4991,N_4955);
nor U5045 (N_5045,N_4852,N_4984);
nand U5046 (N_5046,N_4912,N_4876);
nand U5047 (N_5047,N_4960,N_4889);
xor U5048 (N_5048,N_4831,N_4865);
nor U5049 (N_5049,N_4971,N_4932);
nor U5050 (N_5050,N_4826,N_4944);
xor U5051 (N_5051,N_4879,N_4947);
and U5052 (N_5052,N_4970,N_4827);
nand U5053 (N_5053,N_4832,N_4893);
nor U5054 (N_5054,N_4823,N_4877);
xnor U5055 (N_5055,N_4828,N_4860);
and U5056 (N_5056,N_4870,N_4900);
xnor U5057 (N_5057,N_4982,N_4829);
nand U5058 (N_5058,N_4839,N_4811);
nor U5059 (N_5059,N_4863,N_4951);
xor U5060 (N_5060,N_4875,N_4858);
nand U5061 (N_5061,N_4898,N_4886);
and U5062 (N_5062,N_4981,N_4928);
xor U5063 (N_5063,N_4986,N_4802);
xnor U5064 (N_5064,N_4859,N_4929);
nand U5065 (N_5065,N_4942,N_4887);
or U5066 (N_5066,N_4847,N_4836);
xnor U5067 (N_5067,N_4807,N_4830);
or U5068 (N_5068,N_4801,N_4866);
or U5069 (N_5069,N_4910,N_4883);
nand U5070 (N_5070,N_4814,N_4946);
nor U5071 (N_5071,N_4907,N_4849);
xor U5072 (N_5072,N_4950,N_4973);
and U5073 (N_5073,N_4850,N_4956);
nor U5074 (N_5074,N_4940,N_4949);
nand U5075 (N_5075,N_4969,N_4851);
xor U5076 (N_5076,N_4853,N_4926);
or U5077 (N_5077,N_4821,N_4881);
and U5078 (N_5078,N_4845,N_4817);
nor U5079 (N_5079,N_4925,N_4943);
nor U5080 (N_5080,N_4920,N_4923);
nand U5081 (N_5081,N_4874,N_4948);
or U5082 (N_5082,N_4919,N_4915);
xor U5083 (N_5083,N_4818,N_4966);
and U5084 (N_5084,N_4835,N_4805);
or U5085 (N_5085,N_4842,N_4941);
nor U5086 (N_5086,N_4843,N_4878);
nor U5087 (N_5087,N_4967,N_4903);
or U5088 (N_5088,N_4815,N_4909);
and U5089 (N_5089,N_4899,N_4921);
nand U5090 (N_5090,N_4974,N_4895);
nor U5091 (N_5091,N_4930,N_4834);
nand U5092 (N_5092,N_4945,N_4885);
or U5093 (N_5093,N_4813,N_4846);
nor U5094 (N_5094,N_4825,N_4934);
xor U5095 (N_5095,N_4978,N_4833);
xor U5096 (N_5096,N_4979,N_4963);
nand U5097 (N_5097,N_4804,N_4933);
nand U5098 (N_5098,N_4906,N_4968);
nor U5099 (N_5099,N_4985,N_4939);
nand U5100 (N_5100,N_4856,N_4876);
nand U5101 (N_5101,N_4818,N_4801);
nand U5102 (N_5102,N_4853,N_4852);
or U5103 (N_5103,N_4997,N_4930);
nand U5104 (N_5104,N_4904,N_4873);
or U5105 (N_5105,N_4843,N_4897);
xnor U5106 (N_5106,N_4860,N_4864);
or U5107 (N_5107,N_4990,N_4951);
or U5108 (N_5108,N_4805,N_4856);
or U5109 (N_5109,N_4801,N_4809);
xor U5110 (N_5110,N_4811,N_4924);
xor U5111 (N_5111,N_4974,N_4828);
nor U5112 (N_5112,N_4950,N_4991);
nor U5113 (N_5113,N_4891,N_4807);
and U5114 (N_5114,N_4841,N_4933);
nand U5115 (N_5115,N_4895,N_4897);
nor U5116 (N_5116,N_4953,N_4995);
or U5117 (N_5117,N_4824,N_4922);
and U5118 (N_5118,N_4897,N_4818);
and U5119 (N_5119,N_4830,N_4957);
xor U5120 (N_5120,N_4869,N_4879);
and U5121 (N_5121,N_4926,N_4869);
nand U5122 (N_5122,N_4826,N_4832);
xnor U5123 (N_5123,N_4862,N_4910);
nor U5124 (N_5124,N_4873,N_4945);
xnor U5125 (N_5125,N_4982,N_4873);
xnor U5126 (N_5126,N_4958,N_4902);
nand U5127 (N_5127,N_4805,N_4941);
xnor U5128 (N_5128,N_4884,N_4803);
and U5129 (N_5129,N_4901,N_4998);
xor U5130 (N_5130,N_4893,N_4977);
nor U5131 (N_5131,N_4846,N_4960);
xor U5132 (N_5132,N_4975,N_4868);
or U5133 (N_5133,N_4973,N_4893);
xnor U5134 (N_5134,N_4827,N_4832);
and U5135 (N_5135,N_4979,N_4998);
or U5136 (N_5136,N_4964,N_4838);
nand U5137 (N_5137,N_4967,N_4816);
nand U5138 (N_5138,N_4805,N_4935);
or U5139 (N_5139,N_4875,N_4922);
and U5140 (N_5140,N_4882,N_4851);
nor U5141 (N_5141,N_4828,N_4977);
or U5142 (N_5142,N_4976,N_4863);
xnor U5143 (N_5143,N_4954,N_4934);
nand U5144 (N_5144,N_4945,N_4962);
or U5145 (N_5145,N_4936,N_4818);
nor U5146 (N_5146,N_4863,N_4884);
or U5147 (N_5147,N_4893,N_4860);
nand U5148 (N_5148,N_4953,N_4867);
nor U5149 (N_5149,N_4929,N_4919);
xnor U5150 (N_5150,N_4941,N_4848);
xor U5151 (N_5151,N_4945,N_4989);
nor U5152 (N_5152,N_4961,N_4906);
and U5153 (N_5153,N_4977,N_4841);
nand U5154 (N_5154,N_4853,N_4955);
and U5155 (N_5155,N_4836,N_4962);
and U5156 (N_5156,N_4817,N_4847);
nand U5157 (N_5157,N_4860,N_4824);
nor U5158 (N_5158,N_4894,N_4981);
nand U5159 (N_5159,N_4964,N_4897);
xnor U5160 (N_5160,N_4901,N_4906);
xnor U5161 (N_5161,N_4848,N_4853);
and U5162 (N_5162,N_4997,N_4864);
and U5163 (N_5163,N_4800,N_4878);
xor U5164 (N_5164,N_4932,N_4878);
and U5165 (N_5165,N_4980,N_4810);
nor U5166 (N_5166,N_4801,N_4867);
and U5167 (N_5167,N_4972,N_4938);
xor U5168 (N_5168,N_4832,N_4972);
nand U5169 (N_5169,N_4810,N_4809);
or U5170 (N_5170,N_4825,N_4909);
xor U5171 (N_5171,N_4880,N_4879);
xnor U5172 (N_5172,N_4859,N_4846);
and U5173 (N_5173,N_4999,N_4951);
xnor U5174 (N_5174,N_4938,N_4934);
or U5175 (N_5175,N_4803,N_4969);
and U5176 (N_5176,N_4853,N_4972);
nand U5177 (N_5177,N_4829,N_4925);
or U5178 (N_5178,N_4956,N_4960);
and U5179 (N_5179,N_4848,N_4849);
nand U5180 (N_5180,N_4824,N_4972);
nand U5181 (N_5181,N_4917,N_4942);
and U5182 (N_5182,N_4965,N_4858);
xnor U5183 (N_5183,N_4993,N_4998);
and U5184 (N_5184,N_4953,N_4860);
or U5185 (N_5185,N_4957,N_4840);
nor U5186 (N_5186,N_4896,N_4980);
nand U5187 (N_5187,N_4950,N_4882);
or U5188 (N_5188,N_4921,N_4834);
and U5189 (N_5189,N_4868,N_4851);
or U5190 (N_5190,N_4984,N_4803);
and U5191 (N_5191,N_4824,N_4890);
or U5192 (N_5192,N_4885,N_4835);
or U5193 (N_5193,N_4853,N_4881);
or U5194 (N_5194,N_4871,N_4846);
xnor U5195 (N_5195,N_4987,N_4947);
xnor U5196 (N_5196,N_4800,N_4908);
and U5197 (N_5197,N_4992,N_4927);
and U5198 (N_5198,N_4857,N_4829);
xor U5199 (N_5199,N_4914,N_4920);
nand U5200 (N_5200,N_5128,N_5053);
or U5201 (N_5201,N_5129,N_5119);
xnor U5202 (N_5202,N_5165,N_5180);
or U5203 (N_5203,N_5127,N_5070);
or U5204 (N_5204,N_5090,N_5025);
nor U5205 (N_5205,N_5175,N_5142);
xor U5206 (N_5206,N_5084,N_5140);
nor U5207 (N_5207,N_5195,N_5063);
and U5208 (N_5208,N_5011,N_5033);
or U5209 (N_5209,N_5081,N_5174);
nand U5210 (N_5210,N_5169,N_5096);
nor U5211 (N_5211,N_5125,N_5132);
xnor U5212 (N_5212,N_5173,N_5170);
or U5213 (N_5213,N_5130,N_5167);
xnor U5214 (N_5214,N_5027,N_5186);
or U5215 (N_5215,N_5143,N_5137);
xor U5216 (N_5216,N_5041,N_5120);
and U5217 (N_5217,N_5021,N_5079);
nor U5218 (N_5218,N_5184,N_5089);
or U5219 (N_5219,N_5156,N_5022);
nand U5220 (N_5220,N_5133,N_5150);
or U5221 (N_5221,N_5151,N_5073);
xor U5222 (N_5222,N_5005,N_5039);
or U5223 (N_5223,N_5057,N_5026);
or U5224 (N_5224,N_5135,N_5024);
nand U5225 (N_5225,N_5122,N_5048);
xor U5226 (N_5226,N_5091,N_5123);
xnor U5227 (N_5227,N_5064,N_5077);
xor U5228 (N_5228,N_5065,N_5109);
nor U5229 (N_5229,N_5160,N_5062);
or U5230 (N_5230,N_5056,N_5043);
nand U5231 (N_5231,N_5085,N_5115);
nand U5232 (N_5232,N_5030,N_5074);
xnor U5233 (N_5233,N_5076,N_5016);
nor U5234 (N_5234,N_5078,N_5072);
nor U5235 (N_5235,N_5094,N_5032);
nor U5236 (N_5236,N_5162,N_5001);
or U5237 (N_5237,N_5055,N_5058);
nand U5238 (N_5238,N_5023,N_5116);
xnor U5239 (N_5239,N_5161,N_5112);
xnor U5240 (N_5240,N_5187,N_5188);
nand U5241 (N_5241,N_5059,N_5158);
and U5242 (N_5242,N_5000,N_5086);
xnor U5243 (N_5243,N_5110,N_5189);
or U5244 (N_5244,N_5052,N_5003);
nand U5245 (N_5245,N_5098,N_5149);
or U5246 (N_5246,N_5136,N_5080);
and U5247 (N_5247,N_5154,N_5019);
or U5248 (N_5248,N_5159,N_5017);
or U5249 (N_5249,N_5177,N_5002);
xor U5250 (N_5250,N_5199,N_5102);
nand U5251 (N_5251,N_5126,N_5181);
nand U5252 (N_5252,N_5100,N_5166);
xnor U5253 (N_5253,N_5157,N_5147);
nor U5254 (N_5254,N_5131,N_5028);
nand U5255 (N_5255,N_5018,N_5145);
nand U5256 (N_5256,N_5164,N_5050);
nor U5257 (N_5257,N_5108,N_5038);
and U5258 (N_5258,N_5067,N_5106);
xnor U5259 (N_5259,N_5117,N_5095);
and U5260 (N_5260,N_5071,N_5104);
nand U5261 (N_5261,N_5172,N_5114);
xnor U5262 (N_5262,N_5118,N_5113);
xnor U5263 (N_5263,N_5191,N_5182);
xnor U5264 (N_5264,N_5007,N_5168);
xor U5265 (N_5265,N_5049,N_5082);
nand U5266 (N_5266,N_5178,N_5008);
and U5267 (N_5267,N_5068,N_5171);
nand U5268 (N_5268,N_5193,N_5034);
nand U5269 (N_5269,N_5141,N_5031);
nand U5270 (N_5270,N_5146,N_5006);
nor U5271 (N_5271,N_5045,N_5066);
or U5272 (N_5272,N_5036,N_5107);
nor U5273 (N_5273,N_5144,N_5183);
xor U5274 (N_5274,N_5194,N_5051);
or U5275 (N_5275,N_5035,N_5179);
xnor U5276 (N_5276,N_5185,N_5138);
or U5277 (N_5277,N_5020,N_5139);
and U5278 (N_5278,N_5097,N_5015);
nor U5279 (N_5279,N_5013,N_5037);
or U5280 (N_5280,N_5010,N_5155);
nor U5281 (N_5281,N_5190,N_5121);
xor U5282 (N_5282,N_5069,N_5029);
or U5283 (N_5283,N_5103,N_5040);
and U5284 (N_5284,N_5152,N_5101);
nor U5285 (N_5285,N_5192,N_5044);
nand U5286 (N_5286,N_5099,N_5093);
nand U5287 (N_5287,N_5153,N_5105);
or U5288 (N_5288,N_5054,N_5092);
xnor U5289 (N_5289,N_5060,N_5088);
and U5290 (N_5290,N_5124,N_5012);
nand U5291 (N_5291,N_5134,N_5196);
or U5292 (N_5292,N_5176,N_5042);
nor U5293 (N_5293,N_5148,N_5061);
or U5294 (N_5294,N_5046,N_5087);
and U5295 (N_5295,N_5163,N_5198);
or U5296 (N_5296,N_5075,N_5014);
nor U5297 (N_5297,N_5047,N_5083);
or U5298 (N_5298,N_5111,N_5009);
or U5299 (N_5299,N_5004,N_5197);
nor U5300 (N_5300,N_5016,N_5107);
xnor U5301 (N_5301,N_5132,N_5180);
and U5302 (N_5302,N_5050,N_5091);
nand U5303 (N_5303,N_5154,N_5190);
and U5304 (N_5304,N_5110,N_5028);
or U5305 (N_5305,N_5154,N_5101);
nor U5306 (N_5306,N_5087,N_5153);
nor U5307 (N_5307,N_5079,N_5085);
nand U5308 (N_5308,N_5161,N_5169);
xnor U5309 (N_5309,N_5003,N_5014);
and U5310 (N_5310,N_5103,N_5034);
nor U5311 (N_5311,N_5074,N_5152);
nand U5312 (N_5312,N_5090,N_5154);
xnor U5313 (N_5313,N_5115,N_5062);
or U5314 (N_5314,N_5102,N_5183);
or U5315 (N_5315,N_5190,N_5103);
nor U5316 (N_5316,N_5095,N_5154);
and U5317 (N_5317,N_5091,N_5004);
and U5318 (N_5318,N_5126,N_5111);
nor U5319 (N_5319,N_5148,N_5179);
nor U5320 (N_5320,N_5084,N_5077);
xnor U5321 (N_5321,N_5181,N_5197);
nor U5322 (N_5322,N_5162,N_5033);
or U5323 (N_5323,N_5000,N_5155);
nand U5324 (N_5324,N_5149,N_5000);
xnor U5325 (N_5325,N_5034,N_5165);
and U5326 (N_5326,N_5155,N_5077);
xor U5327 (N_5327,N_5157,N_5003);
or U5328 (N_5328,N_5182,N_5019);
or U5329 (N_5329,N_5131,N_5082);
xor U5330 (N_5330,N_5113,N_5168);
and U5331 (N_5331,N_5173,N_5162);
nor U5332 (N_5332,N_5018,N_5136);
or U5333 (N_5333,N_5168,N_5000);
nor U5334 (N_5334,N_5098,N_5173);
nor U5335 (N_5335,N_5118,N_5042);
xnor U5336 (N_5336,N_5058,N_5060);
nor U5337 (N_5337,N_5018,N_5097);
xor U5338 (N_5338,N_5051,N_5039);
or U5339 (N_5339,N_5160,N_5002);
and U5340 (N_5340,N_5033,N_5024);
or U5341 (N_5341,N_5100,N_5147);
nor U5342 (N_5342,N_5057,N_5136);
nor U5343 (N_5343,N_5099,N_5143);
and U5344 (N_5344,N_5116,N_5043);
xor U5345 (N_5345,N_5050,N_5166);
nor U5346 (N_5346,N_5171,N_5046);
xor U5347 (N_5347,N_5028,N_5164);
and U5348 (N_5348,N_5161,N_5029);
xor U5349 (N_5349,N_5097,N_5118);
nor U5350 (N_5350,N_5137,N_5154);
and U5351 (N_5351,N_5124,N_5075);
or U5352 (N_5352,N_5177,N_5011);
or U5353 (N_5353,N_5074,N_5131);
and U5354 (N_5354,N_5128,N_5085);
nor U5355 (N_5355,N_5005,N_5152);
xnor U5356 (N_5356,N_5074,N_5108);
nor U5357 (N_5357,N_5045,N_5010);
and U5358 (N_5358,N_5196,N_5089);
nand U5359 (N_5359,N_5070,N_5185);
and U5360 (N_5360,N_5045,N_5131);
and U5361 (N_5361,N_5183,N_5150);
nand U5362 (N_5362,N_5001,N_5149);
and U5363 (N_5363,N_5071,N_5018);
and U5364 (N_5364,N_5157,N_5124);
or U5365 (N_5365,N_5179,N_5178);
xor U5366 (N_5366,N_5071,N_5024);
nand U5367 (N_5367,N_5118,N_5018);
and U5368 (N_5368,N_5126,N_5034);
or U5369 (N_5369,N_5191,N_5108);
nor U5370 (N_5370,N_5040,N_5008);
xnor U5371 (N_5371,N_5109,N_5087);
and U5372 (N_5372,N_5103,N_5141);
or U5373 (N_5373,N_5077,N_5161);
nand U5374 (N_5374,N_5080,N_5115);
nor U5375 (N_5375,N_5071,N_5154);
nor U5376 (N_5376,N_5129,N_5160);
xor U5377 (N_5377,N_5082,N_5164);
nand U5378 (N_5378,N_5151,N_5108);
or U5379 (N_5379,N_5193,N_5081);
and U5380 (N_5380,N_5127,N_5061);
and U5381 (N_5381,N_5065,N_5119);
nor U5382 (N_5382,N_5055,N_5077);
xnor U5383 (N_5383,N_5053,N_5161);
or U5384 (N_5384,N_5167,N_5150);
nand U5385 (N_5385,N_5152,N_5048);
or U5386 (N_5386,N_5110,N_5175);
or U5387 (N_5387,N_5149,N_5164);
nor U5388 (N_5388,N_5135,N_5056);
xor U5389 (N_5389,N_5006,N_5068);
or U5390 (N_5390,N_5058,N_5092);
nor U5391 (N_5391,N_5180,N_5187);
or U5392 (N_5392,N_5171,N_5120);
xnor U5393 (N_5393,N_5071,N_5050);
or U5394 (N_5394,N_5186,N_5126);
nor U5395 (N_5395,N_5165,N_5166);
xor U5396 (N_5396,N_5004,N_5130);
xnor U5397 (N_5397,N_5170,N_5176);
nor U5398 (N_5398,N_5075,N_5083);
xnor U5399 (N_5399,N_5164,N_5084);
xnor U5400 (N_5400,N_5326,N_5368);
or U5401 (N_5401,N_5374,N_5243);
nor U5402 (N_5402,N_5277,N_5349);
nor U5403 (N_5403,N_5288,N_5360);
nand U5404 (N_5404,N_5299,N_5268);
and U5405 (N_5405,N_5208,N_5332);
nor U5406 (N_5406,N_5227,N_5209);
nand U5407 (N_5407,N_5260,N_5356);
and U5408 (N_5408,N_5369,N_5265);
and U5409 (N_5409,N_5397,N_5234);
xnor U5410 (N_5410,N_5310,N_5351);
xnor U5411 (N_5411,N_5314,N_5372);
nand U5412 (N_5412,N_5235,N_5335);
nor U5413 (N_5413,N_5334,N_5321);
nand U5414 (N_5414,N_5377,N_5366);
nor U5415 (N_5415,N_5245,N_5279);
xnor U5416 (N_5416,N_5328,N_5283);
nor U5417 (N_5417,N_5363,N_5286);
or U5418 (N_5418,N_5304,N_5207);
and U5419 (N_5419,N_5362,N_5340);
nor U5420 (N_5420,N_5239,N_5284);
nand U5421 (N_5421,N_5350,N_5364);
or U5422 (N_5422,N_5224,N_5318);
nor U5423 (N_5423,N_5223,N_5258);
nor U5424 (N_5424,N_5355,N_5342);
nor U5425 (N_5425,N_5202,N_5359);
or U5426 (N_5426,N_5385,N_5241);
xnor U5427 (N_5427,N_5222,N_5232);
nand U5428 (N_5428,N_5389,N_5343);
or U5429 (N_5429,N_5201,N_5392);
xnor U5430 (N_5430,N_5386,N_5327);
xnor U5431 (N_5431,N_5300,N_5252);
nand U5432 (N_5432,N_5253,N_5383);
xnor U5433 (N_5433,N_5290,N_5256);
nand U5434 (N_5434,N_5379,N_5278);
and U5435 (N_5435,N_5200,N_5229);
and U5436 (N_5436,N_5352,N_5302);
or U5437 (N_5437,N_5308,N_5271);
nor U5438 (N_5438,N_5275,N_5262);
or U5439 (N_5439,N_5396,N_5249);
nand U5440 (N_5440,N_5269,N_5338);
nand U5441 (N_5441,N_5381,N_5387);
or U5442 (N_5442,N_5344,N_5367);
nor U5443 (N_5443,N_5211,N_5373);
nand U5444 (N_5444,N_5212,N_5358);
and U5445 (N_5445,N_5305,N_5226);
nand U5446 (N_5446,N_5390,N_5274);
nor U5447 (N_5447,N_5217,N_5330);
xor U5448 (N_5448,N_5345,N_5388);
xnor U5449 (N_5449,N_5320,N_5393);
nand U5450 (N_5450,N_5233,N_5336);
xor U5451 (N_5451,N_5246,N_5218);
nand U5452 (N_5452,N_5398,N_5382);
and U5453 (N_5453,N_5376,N_5228);
xor U5454 (N_5454,N_5337,N_5339);
nand U5455 (N_5455,N_5316,N_5216);
or U5456 (N_5456,N_5296,N_5206);
nor U5457 (N_5457,N_5251,N_5348);
and U5458 (N_5458,N_5357,N_5214);
nor U5459 (N_5459,N_5293,N_5213);
xor U5460 (N_5460,N_5298,N_5231);
nand U5461 (N_5461,N_5255,N_5248);
or U5462 (N_5462,N_5378,N_5365);
and U5463 (N_5463,N_5261,N_5282);
nor U5464 (N_5464,N_5322,N_5267);
xor U5465 (N_5465,N_5325,N_5259);
nand U5466 (N_5466,N_5230,N_5303);
and U5467 (N_5467,N_5242,N_5311);
xnor U5468 (N_5468,N_5399,N_5263);
nor U5469 (N_5469,N_5394,N_5204);
nand U5470 (N_5470,N_5354,N_5346);
nor U5471 (N_5471,N_5341,N_5347);
nand U5472 (N_5472,N_5323,N_5301);
nand U5473 (N_5473,N_5375,N_5391);
xnor U5474 (N_5474,N_5315,N_5287);
nor U5475 (N_5475,N_5395,N_5295);
nand U5476 (N_5476,N_5281,N_5240);
nor U5477 (N_5477,N_5220,N_5370);
xnor U5478 (N_5478,N_5225,N_5333);
xnor U5479 (N_5479,N_5210,N_5292);
nand U5480 (N_5480,N_5331,N_5294);
and U5481 (N_5481,N_5264,N_5247);
nor U5482 (N_5482,N_5306,N_5270);
nand U5483 (N_5483,N_5238,N_5254);
nor U5484 (N_5484,N_5312,N_5319);
or U5485 (N_5485,N_5280,N_5205);
nand U5486 (N_5486,N_5324,N_5380);
or U5487 (N_5487,N_5250,N_5329);
xor U5488 (N_5488,N_5297,N_5203);
or U5489 (N_5489,N_5236,N_5371);
nor U5490 (N_5490,N_5285,N_5289);
nor U5491 (N_5491,N_5257,N_5353);
nand U5492 (N_5492,N_5309,N_5273);
nand U5493 (N_5493,N_5266,N_5272);
and U5494 (N_5494,N_5317,N_5361);
nand U5495 (N_5495,N_5291,N_5307);
xnor U5496 (N_5496,N_5215,N_5313);
nand U5497 (N_5497,N_5237,N_5244);
xor U5498 (N_5498,N_5384,N_5219);
or U5499 (N_5499,N_5221,N_5276);
nand U5500 (N_5500,N_5308,N_5217);
nand U5501 (N_5501,N_5281,N_5233);
or U5502 (N_5502,N_5303,N_5203);
xnor U5503 (N_5503,N_5369,N_5289);
and U5504 (N_5504,N_5363,N_5306);
or U5505 (N_5505,N_5271,N_5374);
nor U5506 (N_5506,N_5213,N_5389);
or U5507 (N_5507,N_5323,N_5353);
and U5508 (N_5508,N_5245,N_5241);
and U5509 (N_5509,N_5370,N_5291);
nand U5510 (N_5510,N_5379,N_5367);
nand U5511 (N_5511,N_5313,N_5211);
and U5512 (N_5512,N_5281,N_5378);
or U5513 (N_5513,N_5306,N_5284);
and U5514 (N_5514,N_5304,N_5213);
nand U5515 (N_5515,N_5220,N_5365);
xnor U5516 (N_5516,N_5330,N_5295);
and U5517 (N_5517,N_5236,N_5272);
xor U5518 (N_5518,N_5287,N_5378);
xor U5519 (N_5519,N_5247,N_5256);
and U5520 (N_5520,N_5365,N_5342);
and U5521 (N_5521,N_5264,N_5356);
nor U5522 (N_5522,N_5203,N_5252);
nor U5523 (N_5523,N_5224,N_5354);
and U5524 (N_5524,N_5270,N_5245);
and U5525 (N_5525,N_5204,N_5365);
xor U5526 (N_5526,N_5394,N_5352);
nor U5527 (N_5527,N_5357,N_5332);
or U5528 (N_5528,N_5236,N_5283);
xor U5529 (N_5529,N_5391,N_5268);
and U5530 (N_5530,N_5354,N_5272);
xnor U5531 (N_5531,N_5202,N_5255);
and U5532 (N_5532,N_5279,N_5274);
xor U5533 (N_5533,N_5273,N_5318);
nand U5534 (N_5534,N_5353,N_5284);
xor U5535 (N_5535,N_5398,N_5315);
nor U5536 (N_5536,N_5246,N_5217);
xor U5537 (N_5537,N_5357,N_5378);
and U5538 (N_5538,N_5241,N_5359);
nor U5539 (N_5539,N_5349,N_5226);
nor U5540 (N_5540,N_5348,N_5253);
xnor U5541 (N_5541,N_5346,N_5231);
or U5542 (N_5542,N_5252,N_5278);
or U5543 (N_5543,N_5264,N_5366);
and U5544 (N_5544,N_5319,N_5285);
or U5545 (N_5545,N_5301,N_5328);
nand U5546 (N_5546,N_5397,N_5317);
and U5547 (N_5547,N_5376,N_5282);
and U5548 (N_5548,N_5332,N_5281);
or U5549 (N_5549,N_5267,N_5332);
xnor U5550 (N_5550,N_5274,N_5230);
nand U5551 (N_5551,N_5306,N_5328);
or U5552 (N_5552,N_5216,N_5348);
nand U5553 (N_5553,N_5213,N_5210);
and U5554 (N_5554,N_5389,N_5226);
nor U5555 (N_5555,N_5259,N_5204);
and U5556 (N_5556,N_5284,N_5214);
and U5557 (N_5557,N_5218,N_5317);
nor U5558 (N_5558,N_5386,N_5286);
or U5559 (N_5559,N_5223,N_5347);
nand U5560 (N_5560,N_5322,N_5352);
nand U5561 (N_5561,N_5362,N_5236);
xor U5562 (N_5562,N_5242,N_5398);
xnor U5563 (N_5563,N_5270,N_5264);
nor U5564 (N_5564,N_5269,N_5339);
nor U5565 (N_5565,N_5337,N_5282);
and U5566 (N_5566,N_5364,N_5323);
or U5567 (N_5567,N_5318,N_5235);
or U5568 (N_5568,N_5222,N_5209);
nand U5569 (N_5569,N_5375,N_5237);
and U5570 (N_5570,N_5286,N_5367);
xor U5571 (N_5571,N_5263,N_5350);
xor U5572 (N_5572,N_5244,N_5388);
or U5573 (N_5573,N_5392,N_5358);
or U5574 (N_5574,N_5376,N_5223);
or U5575 (N_5575,N_5248,N_5291);
xnor U5576 (N_5576,N_5275,N_5316);
and U5577 (N_5577,N_5297,N_5277);
nor U5578 (N_5578,N_5357,N_5369);
and U5579 (N_5579,N_5349,N_5396);
and U5580 (N_5580,N_5328,N_5206);
xor U5581 (N_5581,N_5222,N_5394);
nor U5582 (N_5582,N_5271,N_5389);
or U5583 (N_5583,N_5290,N_5302);
nor U5584 (N_5584,N_5209,N_5352);
nor U5585 (N_5585,N_5308,N_5391);
xor U5586 (N_5586,N_5280,N_5335);
xor U5587 (N_5587,N_5204,N_5205);
or U5588 (N_5588,N_5244,N_5269);
and U5589 (N_5589,N_5320,N_5388);
nor U5590 (N_5590,N_5227,N_5384);
and U5591 (N_5591,N_5298,N_5271);
or U5592 (N_5592,N_5369,N_5294);
or U5593 (N_5593,N_5260,N_5279);
and U5594 (N_5594,N_5223,N_5231);
nand U5595 (N_5595,N_5355,N_5285);
and U5596 (N_5596,N_5229,N_5396);
and U5597 (N_5597,N_5301,N_5399);
nor U5598 (N_5598,N_5328,N_5251);
nor U5599 (N_5599,N_5307,N_5233);
nand U5600 (N_5600,N_5555,N_5547);
nor U5601 (N_5601,N_5494,N_5435);
nor U5602 (N_5602,N_5585,N_5451);
xor U5603 (N_5603,N_5568,N_5471);
nor U5604 (N_5604,N_5535,N_5488);
or U5605 (N_5605,N_5592,N_5566);
nand U5606 (N_5606,N_5482,N_5407);
xnor U5607 (N_5607,N_5405,N_5519);
and U5608 (N_5608,N_5586,N_5560);
and U5609 (N_5609,N_5443,N_5591);
and U5610 (N_5610,N_5543,N_5480);
or U5611 (N_5611,N_5453,N_5576);
or U5612 (N_5612,N_5424,N_5550);
nor U5613 (N_5613,N_5595,N_5511);
nor U5614 (N_5614,N_5402,N_5489);
and U5615 (N_5615,N_5524,N_5452);
xor U5616 (N_5616,N_5504,N_5593);
nor U5617 (N_5617,N_5573,N_5429);
xor U5618 (N_5618,N_5571,N_5532);
xor U5619 (N_5619,N_5458,N_5470);
nor U5620 (N_5620,N_5438,N_5503);
or U5621 (N_5621,N_5523,N_5401);
or U5622 (N_5622,N_5469,N_5414);
and U5623 (N_5623,N_5428,N_5427);
or U5624 (N_5624,N_5439,N_5588);
nor U5625 (N_5625,N_5485,N_5520);
or U5626 (N_5626,N_5589,N_5587);
nor U5627 (N_5627,N_5477,N_5457);
or U5628 (N_5628,N_5476,N_5446);
or U5629 (N_5629,N_5464,N_5490);
nand U5630 (N_5630,N_5516,N_5472);
and U5631 (N_5631,N_5584,N_5580);
and U5632 (N_5632,N_5509,N_5463);
nor U5633 (N_5633,N_5468,N_5487);
xnor U5634 (N_5634,N_5556,N_5459);
and U5635 (N_5635,N_5409,N_5534);
nor U5636 (N_5636,N_5531,N_5411);
nor U5637 (N_5637,N_5492,N_5542);
nor U5638 (N_5638,N_5575,N_5467);
or U5639 (N_5639,N_5403,N_5473);
or U5640 (N_5640,N_5420,N_5456);
and U5641 (N_5641,N_5474,N_5538);
and U5642 (N_5642,N_5551,N_5594);
and U5643 (N_5643,N_5508,N_5436);
or U5644 (N_5644,N_5440,N_5572);
or U5645 (N_5645,N_5537,N_5599);
nor U5646 (N_5646,N_5400,N_5583);
or U5647 (N_5647,N_5433,N_5430);
or U5648 (N_5648,N_5559,N_5522);
xor U5649 (N_5649,N_5525,N_5431);
and U5650 (N_5650,N_5496,N_5432);
xor U5651 (N_5651,N_5505,N_5499);
and U5652 (N_5652,N_5455,N_5461);
nand U5653 (N_5653,N_5478,N_5521);
nor U5654 (N_5654,N_5421,N_5422);
nor U5655 (N_5655,N_5491,N_5527);
nand U5656 (N_5656,N_5404,N_5413);
xnor U5657 (N_5657,N_5498,N_5481);
nor U5658 (N_5658,N_5416,N_5529);
nor U5659 (N_5659,N_5483,N_5449);
nand U5660 (N_5660,N_5500,N_5465);
or U5661 (N_5661,N_5544,N_5493);
nand U5662 (N_5662,N_5526,N_5581);
nor U5663 (N_5663,N_5513,N_5501);
or U5664 (N_5664,N_5548,N_5558);
nor U5665 (N_5665,N_5450,N_5442);
xnor U5666 (N_5666,N_5484,N_5475);
nand U5667 (N_5667,N_5530,N_5466);
nor U5668 (N_5668,N_5553,N_5408);
or U5669 (N_5669,N_5512,N_5495);
xor U5670 (N_5670,N_5417,N_5445);
and U5671 (N_5671,N_5574,N_5486);
xnor U5672 (N_5672,N_5539,N_5561);
and U5673 (N_5673,N_5460,N_5517);
and U5674 (N_5674,N_5418,N_5447);
or U5675 (N_5675,N_5506,N_5406);
or U5676 (N_5676,N_5444,N_5565);
xor U5677 (N_5677,N_5582,N_5514);
xor U5678 (N_5678,N_5552,N_5557);
or U5679 (N_5679,N_5410,N_5567);
nor U5680 (N_5680,N_5549,N_5545);
xor U5681 (N_5681,N_5518,N_5579);
nor U5682 (N_5682,N_5578,N_5415);
xor U5683 (N_5683,N_5454,N_5448);
or U5684 (N_5684,N_5597,N_5541);
and U5685 (N_5685,N_5564,N_5510);
or U5686 (N_5686,N_5554,N_5441);
or U5687 (N_5687,N_5412,N_5590);
and U5688 (N_5688,N_5507,N_5528);
nor U5689 (N_5689,N_5540,N_5479);
nor U5690 (N_5690,N_5434,N_5536);
or U5691 (N_5691,N_5569,N_5462);
and U5692 (N_5692,N_5563,N_5562);
nor U5693 (N_5693,N_5577,N_5570);
and U5694 (N_5694,N_5596,N_5426);
nand U5695 (N_5695,N_5437,N_5497);
and U5696 (N_5696,N_5423,N_5598);
and U5697 (N_5697,N_5546,N_5425);
nand U5698 (N_5698,N_5533,N_5419);
and U5699 (N_5699,N_5502,N_5515);
nor U5700 (N_5700,N_5543,N_5484);
and U5701 (N_5701,N_5530,N_5522);
xnor U5702 (N_5702,N_5583,N_5512);
nor U5703 (N_5703,N_5574,N_5591);
or U5704 (N_5704,N_5433,N_5584);
or U5705 (N_5705,N_5440,N_5599);
or U5706 (N_5706,N_5499,N_5431);
or U5707 (N_5707,N_5538,N_5436);
or U5708 (N_5708,N_5412,N_5450);
xnor U5709 (N_5709,N_5567,N_5542);
nand U5710 (N_5710,N_5480,N_5420);
xnor U5711 (N_5711,N_5524,N_5422);
xnor U5712 (N_5712,N_5439,N_5558);
xor U5713 (N_5713,N_5501,N_5511);
nand U5714 (N_5714,N_5539,N_5453);
nor U5715 (N_5715,N_5596,N_5587);
and U5716 (N_5716,N_5483,N_5562);
and U5717 (N_5717,N_5548,N_5567);
or U5718 (N_5718,N_5476,N_5554);
nand U5719 (N_5719,N_5470,N_5531);
nor U5720 (N_5720,N_5429,N_5435);
and U5721 (N_5721,N_5489,N_5515);
and U5722 (N_5722,N_5557,N_5567);
nor U5723 (N_5723,N_5565,N_5496);
nor U5724 (N_5724,N_5416,N_5504);
xor U5725 (N_5725,N_5556,N_5409);
xnor U5726 (N_5726,N_5596,N_5568);
nor U5727 (N_5727,N_5400,N_5512);
or U5728 (N_5728,N_5411,N_5463);
or U5729 (N_5729,N_5529,N_5460);
nand U5730 (N_5730,N_5556,N_5581);
and U5731 (N_5731,N_5406,N_5494);
nor U5732 (N_5732,N_5445,N_5433);
nand U5733 (N_5733,N_5488,N_5565);
nand U5734 (N_5734,N_5482,N_5577);
or U5735 (N_5735,N_5452,N_5482);
xnor U5736 (N_5736,N_5416,N_5574);
xor U5737 (N_5737,N_5442,N_5408);
and U5738 (N_5738,N_5566,N_5491);
nor U5739 (N_5739,N_5563,N_5427);
nand U5740 (N_5740,N_5580,N_5536);
nor U5741 (N_5741,N_5417,N_5551);
or U5742 (N_5742,N_5507,N_5416);
nand U5743 (N_5743,N_5497,N_5501);
nand U5744 (N_5744,N_5586,N_5419);
xnor U5745 (N_5745,N_5471,N_5456);
xnor U5746 (N_5746,N_5509,N_5538);
xnor U5747 (N_5747,N_5524,N_5562);
and U5748 (N_5748,N_5485,N_5549);
xor U5749 (N_5749,N_5420,N_5557);
nand U5750 (N_5750,N_5433,N_5406);
nand U5751 (N_5751,N_5418,N_5431);
nor U5752 (N_5752,N_5589,N_5404);
nor U5753 (N_5753,N_5490,N_5494);
or U5754 (N_5754,N_5436,N_5462);
nand U5755 (N_5755,N_5503,N_5555);
and U5756 (N_5756,N_5522,N_5510);
nand U5757 (N_5757,N_5469,N_5464);
nor U5758 (N_5758,N_5406,N_5530);
xnor U5759 (N_5759,N_5567,N_5464);
or U5760 (N_5760,N_5575,N_5555);
and U5761 (N_5761,N_5548,N_5501);
and U5762 (N_5762,N_5405,N_5521);
or U5763 (N_5763,N_5567,N_5466);
or U5764 (N_5764,N_5564,N_5546);
nand U5765 (N_5765,N_5404,N_5487);
and U5766 (N_5766,N_5475,N_5476);
and U5767 (N_5767,N_5402,N_5438);
and U5768 (N_5768,N_5425,N_5548);
nand U5769 (N_5769,N_5437,N_5400);
and U5770 (N_5770,N_5478,N_5524);
nor U5771 (N_5771,N_5478,N_5471);
xor U5772 (N_5772,N_5587,N_5549);
nand U5773 (N_5773,N_5471,N_5476);
nand U5774 (N_5774,N_5431,N_5407);
nand U5775 (N_5775,N_5438,N_5578);
or U5776 (N_5776,N_5408,N_5504);
nand U5777 (N_5777,N_5561,N_5579);
xor U5778 (N_5778,N_5522,N_5450);
xnor U5779 (N_5779,N_5567,N_5458);
and U5780 (N_5780,N_5599,N_5487);
and U5781 (N_5781,N_5456,N_5445);
nand U5782 (N_5782,N_5579,N_5467);
nor U5783 (N_5783,N_5437,N_5549);
and U5784 (N_5784,N_5425,N_5480);
or U5785 (N_5785,N_5478,N_5568);
nand U5786 (N_5786,N_5576,N_5528);
or U5787 (N_5787,N_5494,N_5461);
or U5788 (N_5788,N_5501,N_5471);
and U5789 (N_5789,N_5502,N_5571);
or U5790 (N_5790,N_5541,N_5575);
nor U5791 (N_5791,N_5519,N_5415);
nand U5792 (N_5792,N_5572,N_5494);
and U5793 (N_5793,N_5552,N_5486);
nand U5794 (N_5794,N_5497,N_5408);
nand U5795 (N_5795,N_5499,N_5488);
nand U5796 (N_5796,N_5434,N_5537);
nand U5797 (N_5797,N_5431,N_5503);
nor U5798 (N_5798,N_5527,N_5509);
nor U5799 (N_5799,N_5570,N_5402);
and U5800 (N_5800,N_5661,N_5718);
xnor U5801 (N_5801,N_5728,N_5615);
or U5802 (N_5802,N_5771,N_5726);
xnor U5803 (N_5803,N_5622,N_5732);
and U5804 (N_5804,N_5616,N_5768);
and U5805 (N_5805,N_5750,N_5690);
nand U5806 (N_5806,N_5647,N_5796);
or U5807 (N_5807,N_5601,N_5749);
or U5808 (N_5808,N_5740,N_5652);
or U5809 (N_5809,N_5669,N_5610);
and U5810 (N_5810,N_5767,N_5735);
xor U5811 (N_5811,N_5675,N_5739);
xnor U5812 (N_5812,N_5751,N_5752);
nand U5813 (N_5813,N_5632,N_5762);
or U5814 (N_5814,N_5613,N_5797);
nor U5815 (N_5815,N_5788,N_5758);
and U5816 (N_5816,N_5780,N_5608);
nand U5817 (N_5817,N_5686,N_5784);
nand U5818 (N_5818,N_5623,N_5600);
and U5819 (N_5819,N_5770,N_5748);
nor U5820 (N_5820,N_5603,N_5703);
xor U5821 (N_5821,N_5745,N_5799);
nor U5822 (N_5822,N_5709,N_5654);
nand U5823 (N_5823,N_5755,N_5756);
nor U5824 (N_5824,N_5629,N_5602);
or U5825 (N_5825,N_5787,N_5704);
or U5826 (N_5826,N_5697,N_5783);
nor U5827 (N_5827,N_5611,N_5667);
nor U5828 (N_5828,N_5636,N_5722);
nor U5829 (N_5829,N_5638,N_5618);
xor U5830 (N_5830,N_5798,N_5607);
nor U5831 (N_5831,N_5720,N_5736);
or U5832 (N_5832,N_5717,N_5640);
xnor U5833 (N_5833,N_5766,N_5625);
xor U5834 (N_5834,N_5769,N_5648);
nand U5835 (N_5835,N_5782,N_5664);
xnor U5836 (N_5836,N_5670,N_5668);
xor U5837 (N_5837,N_5702,N_5719);
xnor U5838 (N_5838,N_5694,N_5683);
or U5839 (N_5839,N_5662,N_5738);
xor U5840 (N_5840,N_5671,N_5680);
xnor U5841 (N_5841,N_5689,N_5646);
xnor U5842 (N_5842,N_5612,N_5653);
nand U5843 (N_5843,N_5674,N_5743);
or U5844 (N_5844,N_5777,N_5725);
and U5845 (N_5845,N_5779,N_5630);
nand U5846 (N_5846,N_5637,N_5757);
nand U5847 (N_5847,N_5711,N_5744);
nand U5848 (N_5848,N_5715,N_5781);
and U5849 (N_5849,N_5700,N_5631);
xor U5850 (N_5850,N_5692,N_5656);
xnor U5851 (N_5851,N_5775,N_5724);
and U5852 (N_5852,N_5706,N_5685);
nand U5853 (N_5853,N_5641,N_5604);
and U5854 (N_5854,N_5649,N_5624);
nor U5855 (N_5855,N_5655,N_5753);
and U5856 (N_5856,N_5764,N_5672);
nor U5857 (N_5857,N_5731,N_5776);
xor U5858 (N_5858,N_5606,N_5660);
or U5859 (N_5859,N_5733,N_5627);
nand U5860 (N_5860,N_5786,N_5687);
and U5861 (N_5861,N_5614,N_5696);
nor U5862 (N_5862,N_5712,N_5651);
and U5863 (N_5863,N_5737,N_5723);
or U5864 (N_5864,N_5681,N_5794);
nor U5865 (N_5865,N_5679,N_5795);
and U5866 (N_5866,N_5773,N_5609);
and U5867 (N_5867,N_5663,N_5699);
xnor U5868 (N_5868,N_5617,N_5634);
xnor U5869 (N_5869,N_5639,N_5754);
nand U5870 (N_5870,N_5772,N_5730);
nand U5871 (N_5871,N_5716,N_5790);
xnor U5872 (N_5872,N_5642,N_5774);
nor U5873 (N_5873,N_5665,N_5693);
xnor U5874 (N_5874,N_5666,N_5721);
xnor U5875 (N_5875,N_5605,N_5620);
nand U5876 (N_5876,N_5729,N_5676);
or U5877 (N_5877,N_5650,N_5658);
xnor U5878 (N_5878,N_5691,N_5778);
or U5879 (N_5879,N_5727,N_5742);
or U5880 (N_5880,N_5682,N_5761);
nor U5881 (N_5881,N_5759,N_5619);
or U5882 (N_5882,N_5785,N_5714);
nor U5883 (N_5883,N_5747,N_5695);
or U5884 (N_5884,N_5741,N_5791);
and U5885 (N_5885,N_5698,N_5621);
or U5886 (N_5886,N_5684,N_5792);
nor U5887 (N_5887,N_5688,N_5705);
or U5888 (N_5888,N_5710,N_5765);
nand U5889 (N_5889,N_5707,N_5713);
nor U5890 (N_5890,N_5789,N_5628);
nor U5891 (N_5891,N_5708,N_5673);
or U5892 (N_5892,N_5626,N_5746);
or U5893 (N_5893,N_5659,N_5763);
nor U5894 (N_5894,N_5643,N_5677);
nand U5895 (N_5895,N_5760,N_5734);
nor U5896 (N_5896,N_5678,N_5793);
nand U5897 (N_5897,N_5633,N_5644);
xnor U5898 (N_5898,N_5657,N_5635);
or U5899 (N_5899,N_5645,N_5701);
or U5900 (N_5900,N_5726,N_5784);
nand U5901 (N_5901,N_5645,N_5732);
and U5902 (N_5902,N_5717,N_5714);
or U5903 (N_5903,N_5724,N_5790);
and U5904 (N_5904,N_5602,N_5616);
nor U5905 (N_5905,N_5791,N_5682);
or U5906 (N_5906,N_5695,N_5722);
xnor U5907 (N_5907,N_5685,N_5679);
or U5908 (N_5908,N_5645,N_5670);
and U5909 (N_5909,N_5651,N_5786);
or U5910 (N_5910,N_5670,N_5769);
nand U5911 (N_5911,N_5753,N_5748);
nor U5912 (N_5912,N_5733,N_5629);
or U5913 (N_5913,N_5761,N_5695);
and U5914 (N_5914,N_5737,N_5710);
nand U5915 (N_5915,N_5600,N_5622);
and U5916 (N_5916,N_5721,N_5635);
nor U5917 (N_5917,N_5796,N_5765);
and U5918 (N_5918,N_5680,N_5664);
xnor U5919 (N_5919,N_5690,N_5760);
nor U5920 (N_5920,N_5702,N_5645);
nand U5921 (N_5921,N_5603,N_5712);
or U5922 (N_5922,N_5700,N_5703);
nor U5923 (N_5923,N_5794,N_5617);
and U5924 (N_5924,N_5722,N_5664);
and U5925 (N_5925,N_5658,N_5649);
or U5926 (N_5926,N_5626,N_5630);
xor U5927 (N_5927,N_5652,N_5606);
xor U5928 (N_5928,N_5670,N_5734);
nor U5929 (N_5929,N_5669,N_5764);
xor U5930 (N_5930,N_5752,N_5656);
nor U5931 (N_5931,N_5661,N_5779);
or U5932 (N_5932,N_5777,N_5696);
or U5933 (N_5933,N_5736,N_5787);
nand U5934 (N_5934,N_5683,N_5790);
and U5935 (N_5935,N_5638,N_5681);
nand U5936 (N_5936,N_5782,N_5777);
or U5937 (N_5937,N_5708,N_5795);
or U5938 (N_5938,N_5779,N_5689);
and U5939 (N_5939,N_5735,N_5796);
and U5940 (N_5940,N_5738,N_5741);
and U5941 (N_5941,N_5601,N_5754);
or U5942 (N_5942,N_5731,N_5796);
nand U5943 (N_5943,N_5696,N_5734);
nand U5944 (N_5944,N_5650,N_5789);
nand U5945 (N_5945,N_5655,N_5787);
xnor U5946 (N_5946,N_5637,N_5724);
or U5947 (N_5947,N_5747,N_5626);
and U5948 (N_5948,N_5642,N_5735);
and U5949 (N_5949,N_5795,N_5780);
or U5950 (N_5950,N_5735,N_5641);
xnor U5951 (N_5951,N_5640,N_5697);
and U5952 (N_5952,N_5717,N_5651);
nand U5953 (N_5953,N_5612,N_5623);
and U5954 (N_5954,N_5639,N_5702);
or U5955 (N_5955,N_5723,N_5784);
xnor U5956 (N_5956,N_5744,N_5796);
nand U5957 (N_5957,N_5689,N_5622);
nand U5958 (N_5958,N_5771,N_5638);
and U5959 (N_5959,N_5693,N_5601);
or U5960 (N_5960,N_5748,N_5745);
and U5961 (N_5961,N_5792,N_5682);
or U5962 (N_5962,N_5729,N_5626);
and U5963 (N_5963,N_5641,N_5696);
nand U5964 (N_5964,N_5710,N_5771);
and U5965 (N_5965,N_5777,N_5741);
or U5966 (N_5966,N_5613,N_5799);
nor U5967 (N_5967,N_5798,N_5634);
nand U5968 (N_5968,N_5668,N_5651);
and U5969 (N_5969,N_5668,N_5667);
nand U5970 (N_5970,N_5721,N_5692);
xnor U5971 (N_5971,N_5727,N_5779);
nand U5972 (N_5972,N_5747,N_5704);
and U5973 (N_5973,N_5671,N_5704);
xor U5974 (N_5974,N_5745,N_5782);
xor U5975 (N_5975,N_5672,N_5684);
or U5976 (N_5976,N_5638,N_5637);
or U5977 (N_5977,N_5746,N_5719);
nand U5978 (N_5978,N_5702,N_5759);
xnor U5979 (N_5979,N_5601,N_5727);
nand U5980 (N_5980,N_5781,N_5787);
xnor U5981 (N_5981,N_5789,N_5607);
xnor U5982 (N_5982,N_5747,N_5738);
and U5983 (N_5983,N_5616,N_5737);
nor U5984 (N_5984,N_5603,N_5655);
nor U5985 (N_5985,N_5602,N_5768);
nand U5986 (N_5986,N_5692,N_5682);
nor U5987 (N_5987,N_5744,N_5720);
xor U5988 (N_5988,N_5625,N_5637);
nor U5989 (N_5989,N_5681,N_5734);
or U5990 (N_5990,N_5717,N_5617);
and U5991 (N_5991,N_5758,N_5653);
and U5992 (N_5992,N_5751,N_5744);
xor U5993 (N_5993,N_5742,N_5733);
xnor U5994 (N_5994,N_5711,N_5608);
nor U5995 (N_5995,N_5755,N_5760);
and U5996 (N_5996,N_5703,N_5638);
and U5997 (N_5997,N_5775,N_5706);
nand U5998 (N_5998,N_5654,N_5794);
xnor U5999 (N_5999,N_5744,N_5640);
nand U6000 (N_6000,N_5856,N_5994);
xor U6001 (N_6001,N_5952,N_5962);
nor U6002 (N_6002,N_5995,N_5888);
and U6003 (N_6003,N_5875,N_5967);
and U6004 (N_6004,N_5887,N_5928);
and U6005 (N_6005,N_5873,N_5997);
xor U6006 (N_6006,N_5863,N_5963);
xnor U6007 (N_6007,N_5965,N_5883);
and U6008 (N_6008,N_5882,N_5912);
nor U6009 (N_6009,N_5946,N_5972);
nor U6010 (N_6010,N_5868,N_5893);
nor U6011 (N_6011,N_5884,N_5948);
nor U6012 (N_6012,N_5927,N_5907);
xor U6013 (N_6013,N_5957,N_5989);
nor U6014 (N_6014,N_5889,N_5959);
xor U6015 (N_6015,N_5804,N_5854);
nand U6016 (N_6016,N_5853,N_5980);
nand U6017 (N_6017,N_5913,N_5852);
or U6018 (N_6018,N_5945,N_5820);
and U6019 (N_6019,N_5930,N_5845);
and U6020 (N_6020,N_5911,N_5847);
xor U6021 (N_6021,N_5988,N_5809);
and U6022 (N_6022,N_5982,N_5987);
or U6023 (N_6023,N_5929,N_5996);
nor U6024 (N_6024,N_5859,N_5978);
and U6025 (N_6025,N_5814,N_5841);
or U6026 (N_6026,N_5943,N_5885);
or U6027 (N_6027,N_5942,N_5956);
and U6028 (N_6028,N_5899,N_5905);
xor U6029 (N_6029,N_5971,N_5909);
nand U6030 (N_6030,N_5827,N_5810);
or U6031 (N_6031,N_5811,N_5832);
nor U6032 (N_6032,N_5805,N_5984);
nor U6033 (N_6033,N_5917,N_5991);
xnor U6034 (N_6034,N_5834,N_5844);
and U6035 (N_6035,N_5896,N_5937);
nor U6036 (N_6036,N_5877,N_5803);
or U6037 (N_6037,N_5802,N_5822);
and U6038 (N_6038,N_5900,N_5829);
nor U6039 (N_6039,N_5949,N_5955);
or U6040 (N_6040,N_5979,N_5800);
nand U6041 (N_6041,N_5933,N_5990);
or U6042 (N_6042,N_5966,N_5871);
or U6043 (N_6043,N_5861,N_5892);
nor U6044 (N_6044,N_5923,N_5904);
nand U6045 (N_6045,N_5801,N_5813);
or U6046 (N_6046,N_5920,N_5886);
or U6047 (N_6047,N_5842,N_5816);
or U6048 (N_6048,N_5926,N_5993);
or U6049 (N_6049,N_5998,N_5934);
and U6050 (N_6050,N_5817,N_5922);
or U6051 (N_6051,N_5964,N_5910);
nor U6052 (N_6052,N_5869,N_5879);
and U6053 (N_6053,N_5826,N_5823);
nand U6054 (N_6054,N_5846,N_5931);
nand U6055 (N_6055,N_5838,N_5894);
nor U6056 (N_6056,N_5973,N_5936);
nor U6057 (N_6057,N_5836,N_5944);
xnor U6058 (N_6058,N_5858,N_5951);
nand U6059 (N_6059,N_5872,N_5954);
xnor U6060 (N_6060,N_5916,N_5812);
or U6061 (N_6061,N_5968,N_5866);
and U6062 (N_6062,N_5941,N_5881);
and U6063 (N_6063,N_5850,N_5906);
xnor U6064 (N_6064,N_5921,N_5865);
nor U6065 (N_6065,N_5891,N_5862);
or U6066 (N_6066,N_5831,N_5958);
xor U6067 (N_6067,N_5815,N_5870);
nor U6068 (N_6068,N_5953,N_5855);
nand U6069 (N_6069,N_5828,N_5878);
or U6070 (N_6070,N_5821,N_5835);
or U6071 (N_6071,N_5833,N_5938);
nand U6072 (N_6072,N_5864,N_5807);
nand U6073 (N_6073,N_5849,N_5806);
nand U6074 (N_6074,N_5903,N_5975);
xor U6075 (N_6075,N_5901,N_5940);
and U6076 (N_6076,N_5898,N_5919);
or U6077 (N_6077,N_5961,N_5808);
or U6078 (N_6078,N_5969,N_5848);
and U6079 (N_6079,N_5839,N_5867);
and U6080 (N_6080,N_5818,N_5895);
nor U6081 (N_6081,N_5914,N_5939);
xnor U6082 (N_6082,N_5857,N_5897);
xnor U6083 (N_6083,N_5999,N_5851);
nand U6084 (N_6084,N_5976,N_5970);
or U6085 (N_6085,N_5819,N_5837);
or U6086 (N_6086,N_5880,N_5925);
or U6087 (N_6087,N_5840,N_5908);
xor U6088 (N_6088,N_5915,N_5950);
nor U6089 (N_6089,N_5974,N_5830);
xnor U6090 (N_6090,N_5902,N_5947);
and U6091 (N_6091,N_5918,N_5932);
xor U6092 (N_6092,N_5960,N_5924);
and U6093 (N_6093,N_5986,N_5890);
nand U6094 (N_6094,N_5981,N_5824);
or U6095 (N_6095,N_5983,N_5843);
nand U6096 (N_6096,N_5874,N_5825);
nand U6097 (N_6097,N_5977,N_5860);
or U6098 (N_6098,N_5992,N_5935);
nand U6099 (N_6099,N_5876,N_5985);
or U6100 (N_6100,N_5960,N_5866);
and U6101 (N_6101,N_5947,N_5940);
nand U6102 (N_6102,N_5912,N_5868);
nor U6103 (N_6103,N_5939,N_5876);
nand U6104 (N_6104,N_5812,N_5893);
nor U6105 (N_6105,N_5851,N_5811);
nand U6106 (N_6106,N_5973,N_5985);
xor U6107 (N_6107,N_5917,N_5871);
and U6108 (N_6108,N_5818,N_5944);
or U6109 (N_6109,N_5821,N_5985);
xnor U6110 (N_6110,N_5829,N_5813);
xnor U6111 (N_6111,N_5994,N_5872);
and U6112 (N_6112,N_5841,N_5940);
nor U6113 (N_6113,N_5879,N_5801);
nand U6114 (N_6114,N_5874,N_5960);
or U6115 (N_6115,N_5938,N_5928);
xnor U6116 (N_6116,N_5865,N_5876);
nor U6117 (N_6117,N_5850,N_5823);
and U6118 (N_6118,N_5822,N_5943);
nor U6119 (N_6119,N_5808,N_5856);
xnor U6120 (N_6120,N_5922,N_5944);
and U6121 (N_6121,N_5818,N_5830);
nor U6122 (N_6122,N_5829,N_5993);
or U6123 (N_6123,N_5807,N_5991);
nand U6124 (N_6124,N_5817,N_5920);
nand U6125 (N_6125,N_5976,N_5896);
xnor U6126 (N_6126,N_5988,N_5807);
and U6127 (N_6127,N_5994,N_5917);
nand U6128 (N_6128,N_5975,N_5930);
nor U6129 (N_6129,N_5820,N_5866);
or U6130 (N_6130,N_5850,N_5946);
nor U6131 (N_6131,N_5961,N_5990);
nor U6132 (N_6132,N_5980,N_5906);
and U6133 (N_6133,N_5970,N_5948);
or U6134 (N_6134,N_5997,N_5838);
and U6135 (N_6135,N_5811,N_5991);
nor U6136 (N_6136,N_5867,N_5922);
and U6137 (N_6137,N_5864,N_5868);
or U6138 (N_6138,N_5941,N_5855);
or U6139 (N_6139,N_5874,N_5831);
nand U6140 (N_6140,N_5836,N_5983);
nor U6141 (N_6141,N_5866,N_5842);
nand U6142 (N_6142,N_5963,N_5962);
and U6143 (N_6143,N_5908,N_5950);
or U6144 (N_6144,N_5870,N_5826);
xor U6145 (N_6145,N_5892,N_5828);
xnor U6146 (N_6146,N_5829,N_5942);
nand U6147 (N_6147,N_5982,N_5914);
or U6148 (N_6148,N_5972,N_5884);
nand U6149 (N_6149,N_5843,N_5940);
and U6150 (N_6150,N_5917,N_5941);
nand U6151 (N_6151,N_5843,N_5978);
nand U6152 (N_6152,N_5967,N_5974);
and U6153 (N_6153,N_5943,N_5836);
nor U6154 (N_6154,N_5849,N_5917);
nor U6155 (N_6155,N_5811,N_5979);
or U6156 (N_6156,N_5895,N_5810);
and U6157 (N_6157,N_5876,N_5955);
nor U6158 (N_6158,N_5840,N_5946);
xor U6159 (N_6159,N_5845,N_5806);
nor U6160 (N_6160,N_5883,N_5940);
or U6161 (N_6161,N_5956,N_5904);
nand U6162 (N_6162,N_5848,N_5905);
and U6163 (N_6163,N_5966,N_5998);
or U6164 (N_6164,N_5846,N_5894);
nand U6165 (N_6165,N_5849,N_5978);
nor U6166 (N_6166,N_5875,N_5857);
nand U6167 (N_6167,N_5943,N_5830);
xnor U6168 (N_6168,N_5984,N_5980);
and U6169 (N_6169,N_5916,N_5887);
nor U6170 (N_6170,N_5934,N_5854);
xor U6171 (N_6171,N_5848,N_5984);
nand U6172 (N_6172,N_5959,N_5997);
nor U6173 (N_6173,N_5867,N_5977);
or U6174 (N_6174,N_5852,N_5946);
xor U6175 (N_6175,N_5943,N_5947);
xnor U6176 (N_6176,N_5836,N_5892);
nor U6177 (N_6177,N_5914,N_5920);
xnor U6178 (N_6178,N_5827,N_5975);
or U6179 (N_6179,N_5959,N_5993);
xnor U6180 (N_6180,N_5875,N_5999);
nand U6181 (N_6181,N_5815,N_5878);
nor U6182 (N_6182,N_5925,N_5864);
and U6183 (N_6183,N_5879,N_5901);
nand U6184 (N_6184,N_5822,N_5999);
xor U6185 (N_6185,N_5834,N_5849);
and U6186 (N_6186,N_5989,N_5925);
nor U6187 (N_6187,N_5949,N_5951);
and U6188 (N_6188,N_5874,N_5950);
and U6189 (N_6189,N_5967,N_5866);
nand U6190 (N_6190,N_5837,N_5957);
nor U6191 (N_6191,N_5949,N_5891);
nand U6192 (N_6192,N_5887,N_5871);
xor U6193 (N_6193,N_5949,N_5965);
nor U6194 (N_6194,N_5946,N_5958);
nand U6195 (N_6195,N_5808,N_5841);
nor U6196 (N_6196,N_5903,N_5921);
nand U6197 (N_6197,N_5885,N_5824);
xor U6198 (N_6198,N_5985,N_5989);
and U6199 (N_6199,N_5947,N_5916);
nand U6200 (N_6200,N_6183,N_6169);
nor U6201 (N_6201,N_6103,N_6058);
and U6202 (N_6202,N_6082,N_6001);
nand U6203 (N_6203,N_6122,N_6100);
nor U6204 (N_6204,N_6187,N_6197);
nor U6205 (N_6205,N_6036,N_6070);
xnor U6206 (N_6206,N_6092,N_6008);
nand U6207 (N_6207,N_6029,N_6031);
nand U6208 (N_6208,N_6019,N_6140);
and U6209 (N_6209,N_6119,N_6000);
or U6210 (N_6210,N_6083,N_6181);
xnor U6211 (N_6211,N_6113,N_6193);
or U6212 (N_6212,N_6020,N_6054);
or U6213 (N_6213,N_6114,N_6014);
and U6214 (N_6214,N_6060,N_6132);
and U6215 (N_6215,N_6035,N_6079);
xor U6216 (N_6216,N_6097,N_6033);
nor U6217 (N_6217,N_6134,N_6024);
xor U6218 (N_6218,N_6048,N_6121);
xnor U6219 (N_6219,N_6042,N_6088);
xor U6220 (N_6220,N_6126,N_6022);
or U6221 (N_6221,N_6040,N_6018);
and U6222 (N_6222,N_6117,N_6073);
nor U6223 (N_6223,N_6105,N_6072);
or U6224 (N_6224,N_6120,N_6163);
xor U6225 (N_6225,N_6130,N_6170);
or U6226 (N_6226,N_6049,N_6098);
or U6227 (N_6227,N_6050,N_6017);
or U6228 (N_6228,N_6115,N_6127);
xor U6229 (N_6229,N_6086,N_6063);
xor U6230 (N_6230,N_6177,N_6186);
or U6231 (N_6231,N_6030,N_6133);
xor U6232 (N_6232,N_6131,N_6179);
or U6233 (N_6233,N_6046,N_6157);
or U6234 (N_6234,N_6006,N_6009);
xnor U6235 (N_6235,N_6087,N_6081);
nor U6236 (N_6236,N_6165,N_6067);
or U6237 (N_6237,N_6154,N_6023);
nor U6238 (N_6238,N_6153,N_6106);
xor U6239 (N_6239,N_6043,N_6176);
nand U6240 (N_6240,N_6175,N_6016);
xor U6241 (N_6241,N_6109,N_6028);
xor U6242 (N_6242,N_6141,N_6002);
xor U6243 (N_6243,N_6111,N_6041);
nor U6244 (N_6244,N_6150,N_6116);
and U6245 (N_6245,N_6013,N_6032);
nor U6246 (N_6246,N_6160,N_6144);
and U6247 (N_6247,N_6155,N_6012);
and U6248 (N_6248,N_6044,N_6172);
or U6249 (N_6249,N_6069,N_6191);
nand U6250 (N_6250,N_6196,N_6108);
and U6251 (N_6251,N_6164,N_6015);
xor U6252 (N_6252,N_6138,N_6093);
and U6253 (N_6253,N_6107,N_6182);
xor U6254 (N_6254,N_6027,N_6142);
nand U6255 (N_6255,N_6135,N_6156);
or U6256 (N_6256,N_6136,N_6052);
nor U6257 (N_6257,N_6199,N_6077);
nor U6258 (N_6258,N_6146,N_6198);
xor U6259 (N_6259,N_6021,N_6096);
xor U6260 (N_6260,N_6062,N_6034);
or U6261 (N_6261,N_6180,N_6068);
and U6262 (N_6262,N_6104,N_6061);
and U6263 (N_6263,N_6128,N_6192);
xnor U6264 (N_6264,N_6101,N_6149);
nand U6265 (N_6265,N_6089,N_6084);
xnor U6266 (N_6266,N_6037,N_6004);
and U6267 (N_6267,N_6162,N_6059);
xnor U6268 (N_6268,N_6025,N_6074);
or U6269 (N_6269,N_6075,N_6056);
nor U6270 (N_6270,N_6151,N_6064);
nand U6271 (N_6271,N_6152,N_6102);
nand U6272 (N_6272,N_6038,N_6188);
nand U6273 (N_6273,N_6167,N_6085);
and U6274 (N_6274,N_6051,N_6159);
nand U6275 (N_6275,N_6055,N_6005);
or U6276 (N_6276,N_6125,N_6145);
nand U6277 (N_6277,N_6045,N_6112);
or U6278 (N_6278,N_6195,N_6174);
nand U6279 (N_6279,N_6168,N_6010);
xor U6280 (N_6280,N_6053,N_6065);
nand U6281 (N_6281,N_6076,N_6137);
and U6282 (N_6282,N_6094,N_6139);
nor U6283 (N_6283,N_6091,N_6007);
or U6284 (N_6284,N_6147,N_6095);
or U6285 (N_6285,N_6047,N_6099);
nor U6286 (N_6286,N_6118,N_6124);
or U6287 (N_6287,N_6090,N_6066);
nand U6288 (N_6288,N_6148,N_6189);
xnor U6289 (N_6289,N_6184,N_6129);
or U6290 (N_6290,N_6166,N_6185);
nor U6291 (N_6291,N_6110,N_6171);
xnor U6292 (N_6292,N_6190,N_6173);
and U6293 (N_6293,N_6011,N_6003);
and U6294 (N_6294,N_6143,N_6057);
and U6295 (N_6295,N_6194,N_6080);
nor U6296 (N_6296,N_6026,N_6078);
nor U6297 (N_6297,N_6039,N_6158);
or U6298 (N_6298,N_6178,N_6161);
and U6299 (N_6299,N_6123,N_6071);
nand U6300 (N_6300,N_6143,N_6054);
nor U6301 (N_6301,N_6107,N_6193);
nand U6302 (N_6302,N_6165,N_6008);
or U6303 (N_6303,N_6167,N_6027);
nand U6304 (N_6304,N_6074,N_6164);
nor U6305 (N_6305,N_6020,N_6187);
nor U6306 (N_6306,N_6024,N_6053);
xor U6307 (N_6307,N_6036,N_6042);
xor U6308 (N_6308,N_6071,N_6173);
xor U6309 (N_6309,N_6109,N_6003);
or U6310 (N_6310,N_6054,N_6144);
nor U6311 (N_6311,N_6048,N_6167);
nor U6312 (N_6312,N_6089,N_6015);
nor U6313 (N_6313,N_6028,N_6144);
and U6314 (N_6314,N_6115,N_6041);
or U6315 (N_6315,N_6177,N_6076);
and U6316 (N_6316,N_6127,N_6038);
nor U6317 (N_6317,N_6151,N_6173);
and U6318 (N_6318,N_6138,N_6115);
nand U6319 (N_6319,N_6110,N_6175);
nor U6320 (N_6320,N_6116,N_6115);
nand U6321 (N_6321,N_6142,N_6042);
nand U6322 (N_6322,N_6003,N_6054);
and U6323 (N_6323,N_6029,N_6049);
nor U6324 (N_6324,N_6145,N_6132);
or U6325 (N_6325,N_6034,N_6096);
nor U6326 (N_6326,N_6135,N_6103);
xnor U6327 (N_6327,N_6003,N_6055);
and U6328 (N_6328,N_6082,N_6019);
nand U6329 (N_6329,N_6190,N_6080);
or U6330 (N_6330,N_6013,N_6162);
xnor U6331 (N_6331,N_6154,N_6075);
xor U6332 (N_6332,N_6113,N_6029);
xnor U6333 (N_6333,N_6113,N_6006);
nor U6334 (N_6334,N_6022,N_6181);
xnor U6335 (N_6335,N_6025,N_6022);
xnor U6336 (N_6336,N_6028,N_6081);
nand U6337 (N_6337,N_6082,N_6137);
nor U6338 (N_6338,N_6087,N_6120);
xnor U6339 (N_6339,N_6054,N_6059);
and U6340 (N_6340,N_6045,N_6188);
xnor U6341 (N_6341,N_6002,N_6132);
and U6342 (N_6342,N_6158,N_6101);
nor U6343 (N_6343,N_6045,N_6070);
nor U6344 (N_6344,N_6046,N_6020);
or U6345 (N_6345,N_6155,N_6001);
and U6346 (N_6346,N_6095,N_6121);
and U6347 (N_6347,N_6116,N_6155);
and U6348 (N_6348,N_6026,N_6180);
xor U6349 (N_6349,N_6071,N_6080);
and U6350 (N_6350,N_6189,N_6158);
xnor U6351 (N_6351,N_6068,N_6192);
and U6352 (N_6352,N_6043,N_6114);
nor U6353 (N_6353,N_6122,N_6095);
xor U6354 (N_6354,N_6019,N_6130);
xnor U6355 (N_6355,N_6056,N_6173);
xnor U6356 (N_6356,N_6052,N_6001);
xor U6357 (N_6357,N_6108,N_6139);
nand U6358 (N_6358,N_6055,N_6133);
and U6359 (N_6359,N_6066,N_6086);
or U6360 (N_6360,N_6005,N_6160);
and U6361 (N_6361,N_6166,N_6014);
nand U6362 (N_6362,N_6192,N_6190);
nand U6363 (N_6363,N_6068,N_6022);
and U6364 (N_6364,N_6135,N_6083);
and U6365 (N_6365,N_6194,N_6047);
or U6366 (N_6366,N_6061,N_6195);
xnor U6367 (N_6367,N_6198,N_6110);
or U6368 (N_6368,N_6154,N_6158);
xor U6369 (N_6369,N_6047,N_6006);
nand U6370 (N_6370,N_6065,N_6193);
or U6371 (N_6371,N_6176,N_6186);
or U6372 (N_6372,N_6141,N_6085);
xor U6373 (N_6373,N_6040,N_6011);
nand U6374 (N_6374,N_6063,N_6087);
and U6375 (N_6375,N_6190,N_6161);
nor U6376 (N_6376,N_6010,N_6120);
nand U6377 (N_6377,N_6162,N_6192);
xnor U6378 (N_6378,N_6082,N_6105);
or U6379 (N_6379,N_6134,N_6180);
nor U6380 (N_6380,N_6128,N_6029);
and U6381 (N_6381,N_6008,N_6183);
or U6382 (N_6382,N_6014,N_6069);
and U6383 (N_6383,N_6118,N_6066);
and U6384 (N_6384,N_6169,N_6174);
nor U6385 (N_6385,N_6048,N_6194);
or U6386 (N_6386,N_6036,N_6037);
or U6387 (N_6387,N_6014,N_6096);
nand U6388 (N_6388,N_6011,N_6076);
or U6389 (N_6389,N_6161,N_6196);
and U6390 (N_6390,N_6022,N_6137);
or U6391 (N_6391,N_6143,N_6196);
xor U6392 (N_6392,N_6177,N_6063);
nand U6393 (N_6393,N_6108,N_6031);
and U6394 (N_6394,N_6166,N_6114);
and U6395 (N_6395,N_6121,N_6120);
nand U6396 (N_6396,N_6172,N_6179);
or U6397 (N_6397,N_6110,N_6037);
xor U6398 (N_6398,N_6052,N_6166);
or U6399 (N_6399,N_6133,N_6177);
nor U6400 (N_6400,N_6339,N_6205);
and U6401 (N_6401,N_6367,N_6295);
nor U6402 (N_6402,N_6224,N_6371);
and U6403 (N_6403,N_6238,N_6252);
xor U6404 (N_6404,N_6234,N_6341);
and U6405 (N_6405,N_6322,N_6337);
xor U6406 (N_6406,N_6369,N_6290);
nand U6407 (N_6407,N_6316,N_6247);
nor U6408 (N_6408,N_6333,N_6354);
or U6409 (N_6409,N_6397,N_6288);
or U6410 (N_6410,N_6267,N_6216);
and U6411 (N_6411,N_6261,N_6273);
xnor U6412 (N_6412,N_6345,N_6230);
or U6413 (N_6413,N_6235,N_6246);
nand U6414 (N_6414,N_6237,N_6298);
and U6415 (N_6415,N_6262,N_6285);
xor U6416 (N_6416,N_6223,N_6289);
and U6417 (N_6417,N_6349,N_6395);
nand U6418 (N_6418,N_6385,N_6313);
or U6419 (N_6419,N_6356,N_6326);
nand U6420 (N_6420,N_6274,N_6379);
and U6421 (N_6421,N_6372,N_6200);
and U6422 (N_6422,N_6244,N_6324);
and U6423 (N_6423,N_6240,N_6293);
nor U6424 (N_6424,N_6222,N_6334);
and U6425 (N_6425,N_6399,N_6310);
and U6426 (N_6426,N_6355,N_6377);
nor U6427 (N_6427,N_6256,N_6229);
xor U6428 (N_6428,N_6347,N_6281);
nor U6429 (N_6429,N_6340,N_6357);
and U6430 (N_6430,N_6375,N_6306);
and U6431 (N_6431,N_6210,N_6228);
or U6432 (N_6432,N_6232,N_6382);
xnor U6433 (N_6433,N_6364,N_6388);
xor U6434 (N_6434,N_6396,N_6330);
nor U6435 (N_6435,N_6358,N_6265);
nand U6436 (N_6436,N_6319,N_6378);
and U6437 (N_6437,N_6268,N_6303);
xnor U6438 (N_6438,N_6314,N_6329);
xnor U6439 (N_6439,N_6374,N_6225);
or U6440 (N_6440,N_6207,N_6226);
nand U6441 (N_6441,N_6266,N_6325);
and U6442 (N_6442,N_6271,N_6346);
nor U6443 (N_6443,N_6211,N_6227);
nand U6444 (N_6444,N_6208,N_6243);
or U6445 (N_6445,N_6221,N_6304);
nor U6446 (N_6446,N_6391,N_6383);
nand U6447 (N_6447,N_6318,N_6296);
nor U6448 (N_6448,N_6327,N_6352);
nor U6449 (N_6449,N_6250,N_6309);
xor U6450 (N_6450,N_6320,N_6217);
xor U6451 (N_6451,N_6368,N_6203);
xnor U6452 (N_6452,N_6263,N_6373);
and U6453 (N_6453,N_6389,N_6370);
xnor U6454 (N_6454,N_6231,N_6215);
nor U6455 (N_6455,N_6287,N_6251);
xnor U6456 (N_6456,N_6253,N_6301);
or U6457 (N_6457,N_6264,N_6308);
nor U6458 (N_6458,N_6258,N_6311);
nand U6459 (N_6459,N_6393,N_6343);
nor U6460 (N_6460,N_6241,N_6365);
or U6461 (N_6461,N_6328,N_6276);
and U6462 (N_6462,N_6392,N_6272);
or U6463 (N_6463,N_6255,N_6282);
nand U6464 (N_6464,N_6342,N_6362);
xnor U6465 (N_6465,N_6338,N_6348);
xnor U6466 (N_6466,N_6332,N_6218);
nand U6467 (N_6467,N_6291,N_6351);
or U6468 (N_6468,N_6202,N_6321);
and U6469 (N_6469,N_6213,N_6307);
or U6470 (N_6470,N_6353,N_6300);
nor U6471 (N_6471,N_6335,N_6269);
and U6472 (N_6472,N_6380,N_6277);
xnor U6473 (N_6473,N_6279,N_6361);
nor U6474 (N_6474,N_6363,N_6336);
nor U6475 (N_6475,N_6212,N_6220);
xnor U6476 (N_6476,N_6249,N_6359);
xnor U6477 (N_6477,N_6233,N_6236);
nor U6478 (N_6478,N_6315,N_6360);
or U6479 (N_6479,N_6201,N_6317);
and U6480 (N_6480,N_6305,N_6312);
nor U6481 (N_6481,N_6294,N_6254);
and U6482 (N_6482,N_6387,N_6278);
or U6483 (N_6483,N_6283,N_6248);
and U6484 (N_6484,N_6280,N_6214);
or U6485 (N_6485,N_6344,N_6257);
xor U6486 (N_6486,N_6206,N_6390);
or U6487 (N_6487,N_6302,N_6292);
or U6488 (N_6488,N_6398,N_6209);
nand U6489 (N_6489,N_6366,N_6381);
nor U6490 (N_6490,N_6245,N_6331);
nor U6491 (N_6491,N_6394,N_6219);
nor U6492 (N_6492,N_6384,N_6376);
nor U6493 (N_6493,N_6275,N_6239);
nand U6494 (N_6494,N_6242,N_6286);
or U6495 (N_6495,N_6204,N_6386);
or U6496 (N_6496,N_6297,N_6284);
nand U6497 (N_6497,N_6270,N_6259);
nand U6498 (N_6498,N_6260,N_6323);
and U6499 (N_6499,N_6350,N_6299);
or U6500 (N_6500,N_6257,N_6393);
and U6501 (N_6501,N_6314,N_6260);
and U6502 (N_6502,N_6249,N_6221);
nand U6503 (N_6503,N_6282,N_6284);
xnor U6504 (N_6504,N_6377,N_6364);
xnor U6505 (N_6505,N_6236,N_6382);
xor U6506 (N_6506,N_6343,N_6260);
nand U6507 (N_6507,N_6366,N_6221);
or U6508 (N_6508,N_6288,N_6361);
or U6509 (N_6509,N_6320,N_6389);
and U6510 (N_6510,N_6263,N_6236);
nand U6511 (N_6511,N_6239,N_6295);
and U6512 (N_6512,N_6212,N_6338);
xnor U6513 (N_6513,N_6204,N_6281);
nand U6514 (N_6514,N_6369,N_6368);
or U6515 (N_6515,N_6363,N_6347);
nand U6516 (N_6516,N_6370,N_6297);
nor U6517 (N_6517,N_6291,N_6206);
nor U6518 (N_6518,N_6306,N_6213);
and U6519 (N_6519,N_6234,N_6364);
and U6520 (N_6520,N_6233,N_6351);
and U6521 (N_6521,N_6359,N_6397);
and U6522 (N_6522,N_6206,N_6372);
nand U6523 (N_6523,N_6308,N_6381);
nor U6524 (N_6524,N_6282,N_6209);
and U6525 (N_6525,N_6366,N_6370);
xor U6526 (N_6526,N_6288,N_6276);
nand U6527 (N_6527,N_6207,N_6225);
and U6528 (N_6528,N_6281,N_6223);
or U6529 (N_6529,N_6237,N_6384);
xnor U6530 (N_6530,N_6318,N_6246);
nand U6531 (N_6531,N_6292,N_6288);
nor U6532 (N_6532,N_6272,N_6399);
or U6533 (N_6533,N_6313,N_6256);
nor U6534 (N_6534,N_6379,N_6200);
nor U6535 (N_6535,N_6330,N_6240);
xor U6536 (N_6536,N_6291,N_6271);
nor U6537 (N_6537,N_6390,N_6325);
or U6538 (N_6538,N_6316,N_6311);
and U6539 (N_6539,N_6359,N_6312);
nor U6540 (N_6540,N_6223,N_6207);
xnor U6541 (N_6541,N_6308,N_6280);
xnor U6542 (N_6542,N_6296,N_6323);
and U6543 (N_6543,N_6254,N_6336);
nor U6544 (N_6544,N_6371,N_6314);
or U6545 (N_6545,N_6247,N_6386);
and U6546 (N_6546,N_6277,N_6387);
xor U6547 (N_6547,N_6247,N_6245);
nor U6548 (N_6548,N_6358,N_6322);
or U6549 (N_6549,N_6217,N_6336);
or U6550 (N_6550,N_6394,N_6397);
and U6551 (N_6551,N_6299,N_6282);
or U6552 (N_6552,N_6379,N_6321);
and U6553 (N_6553,N_6285,N_6389);
nor U6554 (N_6554,N_6217,N_6382);
and U6555 (N_6555,N_6374,N_6207);
xnor U6556 (N_6556,N_6373,N_6375);
xnor U6557 (N_6557,N_6264,N_6213);
nand U6558 (N_6558,N_6384,N_6261);
or U6559 (N_6559,N_6206,N_6356);
xor U6560 (N_6560,N_6270,N_6279);
xnor U6561 (N_6561,N_6235,N_6264);
nand U6562 (N_6562,N_6379,N_6309);
nor U6563 (N_6563,N_6357,N_6358);
xor U6564 (N_6564,N_6336,N_6238);
or U6565 (N_6565,N_6323,N_6338);
and U6566 (N_6566,N_6283,N_6394);
nand U6567 (N_6567,N_6365,N_6267);
and U6568 (N_6568,N_6307,N_6372);
and U6569 (N_6569,N_6340,N_6215);
nor U6570 (N_6570,N_6325,N_6331);
xnor U6571 (N_6571,N_6312,N_6309);
or U6572 (N_6572,N_6305,N_6295);
xnor U6573 (N_6573,N_6307,N_6239);
nor U6574 (N_6574,N_6362,N_6274);
nor U6575 (N_6575,N_6277,N_6327);
nand U6576 (N_6576,N_6206,N_6326);
xor U6577 (N_6577,N_6370,N_6352);
nor U6578 (N_6578,N_6302,N_6386);
and U6579 (N_6579,N_6286,N_6290);
xor U6580 (N_6580,N_6277,N_6231);
and U6581 (N_6581,N_6215,N_6351);
and U6582 (N_6582,N_6224,N_6368);
and U6583 (N_6583,N_6336,N_6397);
and U6584 (N_6584,N_6383,N_6238);
nor U6585 (N_6585,N_6391,N_6395);
and U6586 (N_6586,N_6356,N_6203);
nor U6587 (N_6587,N_6365,N_6252);
or U6588 (N_6588,N_6268,N_6358);
nand U6589 (N_6589,N_6318,N_6374);
nand U6590 (N_6590,N_6298,N_6270);
and U6591 (N_6591,N_6207,N_6338);
nor U6592 (N_6592,N_6269,N_6381);
or U6593 (N_6593,N_6253,N_6370);
or U6594 (N_6594,N_6355,N_6339);
and U6595 (N_6595,N_6272,N_6215);
or U6596 (N_6596,N_6255,N_6234);
nor U6597 (N_6597,N_6286,N_6389);
and U6598 (N_6598,N_6239,N_6223);
or U6599 (N_6599,N_6352,N_6218);
or U6600 (N_6600,N_6490,N_6473);
or U6601 (N_6601,N_6402,N_6599);
xor U6602 (N_6602,N_6489,N_6522);
xor U6603 (N_6603,N_6432,N_6420);
nor U6604 (N_6604,N_6434,N_6429);
nand U6605 (N_6605,N_6443,N_6463);
or U6606 (N_6606,N_6447,N_6554);
xnor U6607 (N_6607,N_6435,N_6511);
nor U6608 (N_6608,N_6454,N_6530);
xor U6609 (N_6609,N_6566,N_6568);
nor U6610 (N_6610,N_6410,N_6456);
or U6611 (N_6611,N_6567,N_6519);
and U6612 (N_6612,N_6497,N_6563);
nand U6613 (N_6613,N_6585,N_6541);
nand U6614 (N_6614,N_6483,N_6482);
nor U6615 (N_6615,N_6424,N_6527);
nor U6616 (N_6616,N_6575,N_6478);
or U6617 (N_6617,N_6540,N_6413);
and U6618 (N_6618,N_6405,N_6477);
nor U6619 (N_6619,N_6464,N_6593);
xnor U6620 (N_6620,N_6484,N_6556);
xnor U6621 (N_6621,N_6523,N_6553);
and U6622 (N_6622,N_6470,N_6532);
and U6623 (N_6623,N_6516,N_6544);
nor U6624 (N_6624,N_6588,N_6572);
xnor U6625 (N_6625,N_6557,N_6584);
nor U6626 (N_6626,N_6417,N_6573);
and U6627 (N_6627,N_6494,N_6471);
nand U6628 (N_6628,N_6465,N_6431);
nand U6629 (N_6629,N_6472,N_6580);
nand U6630 (N_6630,N_6441,N_6551);
xnor U6631 (N_6631,N_6408,N_6481);
and U6632 (N_6632,N_6550,N_6546);
and U6633 (N_6633,N_6493,N_6533);
or U6634 (N_6634,N_6491,N_6538);
nor U6635 (N_6635,N_6510,N_6590);
and U6636 (N_6636,N_6462,N_6409);
xnor U6637 (N_6637,N_6461,N_6521);
nor U6638 (N_6638,N_6587,N_6440);
and U6639 (N_6639,N_6437,N_6488);
or U6640 (N_6640,N_6452,N_6503);
nand U6641 (N_6641,N_6578,N_6415);
xnor U6642 (N_6642,N_6504,N_6467);
xnor U6643 (N_6643,N_6592,N_6425);
or U6644 (N_6644,N_6555,N_6449);
or U6645 (N_6645,N_6508,N_6496);
nor U6646 (N_6646,N_6535,N_6598);
nand U6647 (N_6647,N_6525,N_6586);
or U6648 (N_6648,N_6559,N_6583);
xor U6649 (N_6649,N_6495,N_6517);
and U6650 (N_6650,N_6547,N_6445);
and U6651 (N_6651,N_6427,N_6597);
xnor U6652 (N_6652,N_6487,N_6562);
nand U6653 (N_6653,N_6529,N_6536);
nand U6654 (N_6654,N_6524,N_6502);
or U6655 (N_6655,N_6401,N_6439);
nand U6656 (N_6656,N_6423,N_6406);
xor U6657 (N_6657,N_6468,N_6560);
nand U6658 (N_6658,N_6499,N_6564);
nor U6659 (N_6659,N_6416,N_6591);
nor U6660 (N_6660,N_6466,N_6596);
nand U6661 (N_6661,N_6561,N_6421);
nand U6662 (N_6662,N_6542,N_6438);
xor U6663 (N_6663,N_6539,N_6528);
nand U6664 (N_6664,N_6512,N_6426);
or U6665 (N_6665,N_6430,N_6507);
nand U6666 (N_6666,N_6419,N_6422);
nand U6667 (N_6667,N_6569,N_6433);
or U6668 (N_6668,N_6428,N_6549);
and U6669 (N_6669,N_6485,N_6534);
and U6670 (N_6670,N_6450,N_6548);
nor U6671 (N_6671,N_6558,N_6595);
and U6672 (N_6672,N_6475,N_6457);
and U6673 (N_6673,N_6436,N_6498);
xor U6674 (N_6674,N_6565,N_6531);
nand U6675 (N_6675,N_6581,N_6412);
xor U6676 (N_6676,N_6492,N_6403);
or U6677 (N_6677,N_6442,N_6509);
or U6678 (N_6678,N_6526,N_6577);
and U6679 (N_6679,N_6543,N_6444);
xor U6680 (N_6680,N_6514,N_6459);
nand U6681 (N_6681,N_6448,N_6513);
or U6682 (N_6682,N_6574,N_6480);
or U6683 (N_6683,N_6506,N_6505);
nand U6684 (N_6684,N_6414,N_6576);
xor U6685 (N_6685,N_6446,N_6469);
nand U6686 (N_6686,N_6537,N_6474);
and U6687 (N_6687,N_6571,N_6453);
and U6688 (N_6688,N_6411,N_6500);
nand U6689 (N_6689,N_6458,N_6552);
nand U6690 (N_6690,N_6589,N_6545);
nor U6691 (N_6691,N_6451,N_6582);
and U6692 (N_6692,N_6520,N_6479);
nor U6693 (N_6693,N_6400,N_6570);
xnor U6694 (N_6694,N_6407,N_6594);
nand U6695 (N_6695,N_6579,N_6404);
or U6696 (N_6696,N_6455,N_6501);
nor U6697 (N_6697,N_6418,N_6515);
and U6698 (N_6698,N_6486,N_6460);
nor U6699 (N_6699,N_6476,N_6518);
and U6700 (N_6700,N_6576,N_6526);
xor U6701 (N_6701,N_6528,N_6585);
xor U6702 (N_6702,N_6462,N_6517);
nand U6703 (N_6703,N_6441,N_6522);
and U6704 (N_6704,N_6444,N_6590);
or U6705 (N_6705,N_6401,N_6455);
xnor U6706 (N_6706,N_6429,N_6416);
or U6707 (N_6707,N_6471,N_6401);
xor U6708 (N_6708,N_6446,N_6574);
or U6709 (N_6709,N_6529,N_6565);
nand U6710 (N_6710,N_6501,N_6513);
nand U6711 (N_6711,N_6497,N_6487);
or U6712 (N_6712,N_6559,N_6580);
nor U6713 (N_6713,N_6417,N_6404);
nand U6714 (N_6714,N_6538,N_6455);
or U6715 (N_6715,N_6575,N_6479);
or U6716 (N_6716,N_6452,N_6457);
or U6717 (N_6717,N_6435,N_6472);
nand U6718 (N_6718,N_6448,N_6523);
and U6719 (N_6719,N_6441,N_6536);
or U6720 (N_6720,N_6423,N_6598);
or U6721 (N_6721,N_6573,N_6463);
nor U6722 (N_6722,N_6583,N_6576);
or U6723 (N_6723,N_6426,N_6535);
or U6724 (N_6724,N_6493,N_6594);
nor U6725 (N_6725,N_6522,N_6544);
xor U6726 (N_6726,N_6470,N_6537);
nor U6727 (N_6727,N_6535,N_6586);
xnor U6728 (N_6728,N_6595,N_6414);
xnor U6729 (N_6729,N_6436,N_6427);
nand U6730 (N_6730,N_6571,N_6547);
or U6731 (N_6731,N_6453,N_6413);
and U6732 (N_6732,N_6451,N_6439);
nor U6733 (N_6733,N_6427,N_6441);
xor U6734 (N_6734,N_6590,N_6407);
xor U6735 (N_6735,N_6524,N_6538);
nand U6736 (N_6736,N_6498,N_6450);
xor U6737 (N_6737,N_6509,N_6592);
nand U6738 (N_6738,N_6505,N_6521);
nor U6739 (N_6739,N_6592,N_6586);
nand U6740 (N_6740,N_6415,N_6404);
and U6741 (N_6741,N_6480,N_6599);
nor U6742 (N_6742,N_6492,N_6464);
and U6743 (N_6743,N_6472,N_6469);
nor U6744 (N_6744,N_6598,N_6418);
xor U6745 (N_6745,N_6464,N_6459);
nand U6746 (N_6746,N_6498,N_6405);
xor U6747 (N_6747,N_6436,N_6424);
nand U6748 (N_6748,N_6520,N_6590);
or U6749 (N_6749,N_6422,N_6570);
xor U6750 (N_6750,N_6536,N_6463);
or U6751 (N_6751,N_6432,N_6503);
nand U6752 (N_6752,N_6429,N_6443);
xor U6753 (N_6753,N_6561,N_6415);
nor U6754 (N_6754,N_6483,N_6408);
xor U6755 (N_6755,N_6502,N_6408);
nand U6756 (N_6756,N_6405,N_6489);
nand U6757 (N_6757,N_6490,N_6596);
and U6758 (N_6758,N_6549,N_6456);
and U6759 (N_6759,N_6540,N_6490);
and U6760 (N_6760,N_6546,N_6594);
xnor U6761 (N_6761,N_6477,N_6457);
or U6762 (N_6762,N_6495,N_6463);
xor U6763 (N_6763,N_6479,N_6468);
and U6764 (N_6764,N_6571,N_6412);
or U6765 (N_6765,N_6402,N_6458);
or U6766 (N_6766,N_6451,N_6405);
nand U6767 (N_6767,N_6489,N_6411);
and U6768 (N_6768,N_6536,N_6476);
nor U6769 (N_6769,N_6493,N_6555);
and U6770 (N_6770,N_6425,N_6489);
and U6771 (N_6771,N_6516,N_6491);
xor U6772 (N_6772,N_6570,N_6404);
or U6773 (N_6773,N_6548,N_6415);
xor U6774 (N_6774,N_6587,N_6432);
or U6775 (N_6775,N_6510,N_6592);
nand U6776 (N_6776,N_6556,N_6532);
or U6777 (N_6777,N_6528,N_6572);
nor U6778 (N_6778,N_6537,N_6586);
and U6779 (N_6779,N_6406,N_6414);
and U6780 (N_6780,N_6416,N_6411);
or U6781 (N_6781,N_6488,N_6560);
and U6782 (N_6782,N_6517,N_6493);
or U6783 (N_6783,N_6535,N_6548);
and U6784 (N_6784,N_6562,N_6447);
nor U6785 (N_6785,N_6497,N_6587);
xnor U6786 (N_6786,N_6564,N_6576);
xnor U6787 (N_6787,N_6460,N_6488);
and U6788 (N_6788,N_6570,N_6545);
xor U6789 (N_6789,N_6451,N_6526);
or U6790 (N_6790,N_6510,N_6591);
nor U6791 (N_6791,N_6474,N_6407);
nor U6792 (N_6792,N_6577,N_6435);
and U6793 (N_6793,N_6541,N_6575);
and U6794 (N_6794,N_6434,N_6526);
nor U6795 (N_6795,N_6430,N_6541);
or U6796 (N_6796,N_6498,N_6428);
nor U6797 (N_6797,N_6499,N_6459);
nand U6798 (N_6798,N_6442,N_6567);
or U6799 (N_6799,N_6426,N_6405);
xnor U6800 (N_6800,N_6742,N_6662);
or U6801 (N_6801,N_6747,N_6652);
nor U6802 (N_6802,N_6791,N_6778);
nor U6803 (N_6803,N_6776,N_6632);
or U6804 (N_6804,N_6725,N_6702);
nand U6805 (N_6805,N_6784,N_6671);
or U6806 (N_6806,N_6658,N_6706);
xor U6807 (N_6807,N_6688,N_6686);
nor U6808 (N_6808,N_6676,N_6746);
xnor U6809 (N_6809,N_6728,N_6783);
nor U6810 (N_6810,N_6796,N_6756);
or U6811 (N_6811,N_6645,N_6714);
or U6812 (N_6812,N_6642,N_6698);
and U6813 (N_6813,N_6692,N_6724);
nand U6814 (N_6814,N_6669,N_6607);
or U6815 (N_6815,N_6666,N_6610);
xor U6816 (N_6816,N_6797,N_6754);
and U6817 (N_6817,N_6628,N_6782);
nand U6818 (N_6818,N_6637,N_6694);
and U6819 (N_6819,N_6729,N_6700);
and U6820 (N_6820,N_6765,N_6624);
xnor U6821 (N_6821,N_6745,N_6731);
or U6822 (N_6822,N_6741,N_6708);
nand U6823 (N_6823,N_6613,N_6744);
or U6824 (N_6824,N_6685,N_6774);
or U6825 (N_6825,N_6654,N_6608);
xnor U6826 (N_6826,N_6718,N_6717);
nor U6827 (N_6827,N_6604,N_6673);
and U6828 (N_6828,N_6674,N_6766);
nor U6829 (N_6829,N_6684,N_6660);
and U6830 (N_6830,N_6722,N_6735);
nand U6831 (N_6831,N_6710,N_6738);
and U6832 (N_6832,N_6627,N_6665);
nor U6833 (N_6833,N_6629,N_6723);
xor U6834 (N_6834,N_6683,N_6643);
and U6835 (N_6835,N_6730,N_6649);
or U6836 (N_6836,N_6733,N_6602);
nand U6837 (N_6837,N_6657,N_6603);
nor U6838 (N_6838,N_6672,N_6650);
and U6839 (N_6839,N_6720,N_6734);
nor U6840 (N_6840,N_6612,N_6701);
and U6841 (N_6841,N_6606,N_6601);
or U6842 (N_6842,N_6775,N_6768);
and U6843 (N_6843,N_6737,N_6758);
nor U6844 (N_6844,N_6677,N_6771);
nor U6845 (N_6845,N_6787,N_6630);
nor U6846 (N_6846,N_6634,N_6795);
nor U6847 (N_6847,N_6689,N_6696);
xor U6848 (N_6848,N_6668,N_6640);
xnor U6849 (N_6849,N_6697,N_6679);
and U6850 (N_6850,N_6616,N_6740);
or U6851 (N_6851,N_6693,N_6777);
or U6852 (N_6852,N_6626,N_6793);
or U6853 (N_6853,N_6681,N_6709);
nor U6854 (N_6854,N_6661,N_6614);
or U6855 (N_6855,N_6769,N_6605);
and U6856 (N_6856,N_6785,N_6799);
and U6857 (N_6857,N_6750,N_6726);
xnor U6858 (N_6858,N_6611,N_6703);
nand U6859 (N_6859,N_6699,N_6759);
and U6860 (N_6860,N_6633,N_6653);
nand U6861 (N_6861,N_6786,N_6760);
nor U6862 (N_6862,N_6682,N_6620);
and U6863 (N_6863,N_6675,N_6625);
or U6864 (N_6864,N_6617,N_6623);
nor U6865 (N_6865,N_6656,N_6764);
nor U6866 (N_6866,N_6631,N_6752);
xnor U6867 (N_6867,N_6773,N_6711);
nor U6868 (N_6868,N_6794,N_6749);
nor U6869 (N_6869,N_6655,N_6646);
and U6870 (N_6870,N_6651,N_6790);
nand U6871 (N_6871,N_6712,N_6687);
and U6872 (N_6872,N_6600,N_6609);
xnor U6873 (N_6873,N_6762,N_6788);
nor U6874 (N_6874,N_6664,N_6727);
nor U6875 (N_6875,N_6678,N_6648);
xor U6876 (N_6876,N_6704,N_6767);
and U6877 (N_6877,N_6621,N_6753);
xor U6878 (N_6878,N_6721,N_6715);
and U6879 (N_6879,N_6732,N_6792);
nor U6880 (N_6880,N_6780,N_6736);
nand U6881 (N_6881,N_6667,N_6695);
xor U6882 (N_6882,N_6639,N_6635);
or U6883 (N_6883,N_6798,N_6618);
nand U6884 (N_6884,N_6716,N_6719);
and U6885 (N_6885,N_6779,N_6636);
and U6886 (N_6886,N_6691,N_6644);
nand U6887 (N_6887,N_6713,N_6680);
nor U6888 (N_6888,N_6789,N_6622);
and U6889 (N_6889,N_6663,N_6743);
nor U6890 (N_6890,N_6772,N_6748);
and U6891 (N_6891,N_6770,N_6739);
nor U6892 (N_6892,N_6751,N_6659);
nor U6893 (N_6893,N_6755,N_6763);
xor U6894 (N_6894,N_6690,N_6781);
xnor U6895 (N_6895,N_6615,N_6641);
nand U6896 (N_6896,N_6757,N_6619);
or U6897 (N_6897,N_6638,N_6705);
or U6898 (N_6898,N_6707,N_6647);
and U6899 (N_6899,N_6670,N_6761);
xnor U6900 (N_6900,N_6761,N_6626);
nor U6901 (N_6901,N_6608,N_6732);
and U6902 (N_6902,N_6632,N_6651);
or U6903 (N_6903,N_6772,N_6692);
xor U6904 (N_6904,N_6740,N_6663);
or U6905 (N_6905,N_6741,N_6656);
or U6906 (N_6906,N_6616,N_6701);
and U6907 (N_6907,N_6743,N_6769);
nand U6908 (N_6908,N_6650,N_6638);
nand U6909 (N_6909,N_6607,N_6689);
nor U6910 (N_6910,N_6703,N_6762);
nor U6911 (N_6911,N_6682,N_6765);
or U6912 (N_6912,N_6734,N_6695);
or U6913 (N_6913,N_6643,N_6661);
and U6914 (N_6914,N_6643,N_6704);
and U6915 (N_6915,N_6796,N_6779);
nor U6916 (N_6916,N_6694,N_6785);
nand U6917 (N_6917,N_6613,N_6741);
xnor U6918 (N_6918,N_6714,N_6769);
or U6919 (N_6919,N_6794,N_6787);
nor U6920 (N_6920,N_6697,N_6635);
xnor U6921 (N_6921,N_6752,N_6758);
and U6922 (N_6922,N_6798,N_6757);
xor U6923 (N_6923,N_6603,N_6650);
xor U6924 (N_6924,N_6642,N_6759);
or U6925 (N_6925,N_6670,N_6626);
nand U6926 (N_6926,N_6673,N_6623);
nand U6927 (N_6927,N_6765,N_6794);
xnor U6928 (N_6928,N_6608,N_6701);
and U6929 (N_6929,N_6680,N_6736);
nor U6930 (N_6930,N_6778,N_6712);
nand U6931 (N_6931,N_6604,N_6741);
nor U6932 (N_6932,N_6789,N_6686);
nand U6933 (N_6933,N_6676,N_6636);
and U6934 (N_6934,N_6682,N_6638);
nand U6935 (N_6935,N_6658,N_6736);
nand U6936 (N_6936,N_6793,N_6783);
or U6937 (N_6937,N_6615,N_6636);
or U6938 (N_6938,N_6754,N_6665);
nand U6939 (N_6939,N_6753,N_6760);
or U6940 (N_6940,N_6738,N_6712);
and U6941 (N_6941,N_6779,N_6717);
or U6942 (N_6942,N_6736,N_6727);
xor U6943 (N_6943,N_6763,N_6726);
nand U6944 (N_6944,N_6706,N_6681);
or U6945 (N_6945,N_6745,N_6612);
or U6946 (N_6946,N_6709,N_6623);
or U6947 (N_6947,N_6676,N_6613);
nor U6948 (N_6948,N_6761,N_6601);
nor U6949 (N_6949,N_6728,N_6704);
and U6950 (N_6950,N_6651,N_6682);
nor U6951 (N_6951,N_6652,N_6769);
nand U6952 (N_6952,N_6610,N_6716);
or U6953 (N_6953,N_6781,N_6712);
or U6954 (N_6954,N_6737,N_6709);
nand U6955 (N_6955,N_6611,N_6690);
and U6956 (N_6956,N_6756,N_6757);
nand U6957 (N_6957,N_6736,N_6701);
nor U6958 (N_6958,N_6771,N_6749);
nor U6959 (N_6959,N_6748,N_6650);
xnor U6960 (N_6960,N_6647,N_6739);
or U6961 (N_6961,N_6624,N_6691);
and U6962 (N_6962,N_6603,N_6666);
and U6963 (N_6963,N_6758,N_6641);
nor U6964 (N_6964,N_6715,N_6716);
and U6965 (N_6965,N_6787,N_6687);
or U6966 (N_6966,N_6625,N_6633);
nand U6967 (N_6967,N_6790,N_6714);
nand U6968 (N_6968,N_6666,N_6629);
xor U6969 (N_6969,N_6703,N_6788);
or U6970 (N_6970,N_6701,N_6786);
nor U6971 (N_6971,N_6701,N_6690);
nand U6972 (N_6972,N_6779,N_6639);
nor U6973 (N_6973,N_6696,N_6652);
nand U6974 (N_6974,N_6716,N_6644);
xnor U6975 (N_6975,N_6712,N_6779);
and U6976 (N_6976,N_6629,N_6684);
or U6977 (N_6977,N_6720,N_6775);
nand U6978 (N_6978,N_6786,N_6656);
or U6979 (N_6979,N_6755,N_6655);
nand U6980 (N_6980,N_6641,N_6619);
nor U6981 (N_6981,N_6675,N_6731);
nand U6982 (N_6982,N_6734,N_6783);
or U6983 (N_6983,N_6709,N_6640);
nor U6984 (N_6984,N_6765,N_6627);
nor U6985 (N_6985,N_6628,N_6794);
or U6986 (N_6986,N_6782,N_6759);
nor U6987 (N_6987,N_6781,N_6740);
or U6988 (N_6988,N_6795,N_6747);
nor U6989 (N_6989,N_6659,N_6739);
nand U6990 (N_6990,N_6706,N_6769);
and U6991 (N_6991,N_6768,N_6602);
or U6992 (N_6992,N_6639,N_6717);
or U6993 (N_6993,N_6761,N_6609);
or U6994 (N_6994,N_6626,N_6603);
nand U6995 (N_6995,N_6606,N_6711);
nor U6996 (N_6996,N_6788,N_6625);
nor U6997 (N_6997,N_6677,N_6670);
nand U6998 (N_6998,N_6702,N_6710);
and U6999 (N_6999,N_6762,N_6719);
nand U7000 (N_7000,N_6999,N_6920);
nor U7001 (N_7001,N_6938,N_6951);
nand U7002 (N_7002,N_6950,N_6902);
nor U7003 (N_7003,N_6857,N_6995);
or U7004 (N_7004,N_6841,N_6947);
or U7005 (N_7005,N_6824,N_6815);
nand U7006 (N_7006,N_6875,N_6946);
nand U7007 (N_7007,N_6819,N_6915);
and U7008 (N_7008,N_6897,N_6944);
xor U7009 (N_7009,N_6949,N_6973);
nand U7010 (N_7010,N_6901,N_6834);
or U7011 (N_7011,N_6921,N_6983);
nand U7012 (N_7012,N_6977,N_6993);
or U7013 (N_7013,N_6856,N_6948);
or U7014 (N_7014,N_6971,N_6894);
nand U7015 (N_7015,N_6839,N_6854);
xor U7016 (N_7016,N_6932,N_6827);
or U7017 (N_7017,N_6840,N_6900);
xnor U7018 (N_7018,N_6838,N_6868);
and U7019 (N_7019,N_6970,N_6805);
and U7020 (N_7020,N_6860,N_6830);
and U7021 (N_7021,N_6982,N_6928);
and U7022 (N_7022,N_6821,N_6810);
xor U7023 (N_7023,N_6986,N_6957);
nand U7024 (N_7024,N_6903,N_6812);
or U7025 (N_7025,N_6861,N_6800);
nor U7026 (N_7026,N_6822,N_6814);
nor U7027 (N_7027,N_6855,N_6943);
xnor U7028 (N_7028,N_6811,N_6828);
nand U7029 (N_7029,N_6876,N_6809);
or U7030 (N_7030,N_6836,N_6833);
nand U7031 (N_7031,N_6985,N_6823);
nand U7032 (N_7032,N_6904,N_6933);
nand U7033 (N_7033,N_6942,N_6955);
and U7034 (N_7034,N_6885,N_6899);
and U7035 (N_7035,N_6882,N_6835);
nor U7036 (N_7036,N_6818,N_6910);
or U7037 (N_7037,N_6887,N_6998);
nor U7038 (N_7038,N_6871,N_6994);
or U7039 (N_7039,N_6848,N_6870);
and U7040 (N_7040,N_6813,N_6969);
nand U7041 (N_7041,N_6892,N_6945);
xor U7042 (N_7042,N_6908,N_6953);
xor U7043 (N_7043,N_6888,N_6865);
nand U7044 (N_7044,N_6852,N_6979);
xor U7045 (N_7045,N_6873,N_6914);
nor U7046 (N_7046,N_6864,N_6867);
xor U7047 (N_7047,N_6962,N_6936);
or U7048 (N_7048,N_6990,N_6826);
or U7049 (N_7049,N_6804,N_6940);
xor U7050 (N_7050,N_6842,N_6924);
and U7051 (N_7051,N_6922,N_6845);
nand U7052 (N_7052,N_6858,N_6803);
xnor U7053 (N_7053,N_6843,N_6992);
and U7054 (N_7054,N_6996,N_6958);
or U7055 (N_7055,N_6967,N_6961);
xor U7056 (N_7056,N_6891,N_6898);
or U7057 (N_7057,N_6987,N_6816);
nand U7058 (N_7058,N_6817,N_6877);
nand U7059 (N_7059,N_6937,N_6984);
or U7060 (N_7060,N_6917,N_6907);
nand U7061 (N_7061,N_6807,N_6906);
nand U7062 (N_7062,N_6976,N_6959);
nor U7063 (N_7063,N_6916,N_6931);
nand U7064 (N_7064,N_6905,N_6978);
or U7065 (N_7065,N_6918,N_6808);
and U7066 (N_7066,N_6954,N_6934);
and U7067 (N_7067,N_6988,N_6863);
nand U7068 (N_7068,N_6896,N_6880);
nor U7069 (N_7069,N_6844,N_6923);
and U7070 (N_7070,N_6884,N_6879);
nand U7071 (N_7071,N_6926,N_6859);
nor U7072 (N_7072,N_6831,N_6929);
or U7073 (N_7073,N_6849,N_6866);
nand U7074 (N_7074,N_6989,N_6832);
xor U7075 (N_7075,N_6980,N_6963);
xor U7076 (N_7076,N_6966,N_6846);
and U7077 (N_7077,N_6935,N_6802);
xnor U7078 (N_7078,N_6853,N_6965);
or U7079 (N_7079,N_6862,N_6952);
nor U7080 (N_7080,N_6939,N_6930);
and U7081 (N_7081,N_6890,N_6893);
xor U7082 (N_7082,N_6869,N_6964);
and U7083 (N_7083,N_6960,N_6968);
nand U7084 (N_7084,N_6927,N_6991);
and U7085 (N_7085,N_6806,N_6847);
nor U7086 (N_7086,N_6919,N_6925);
nand U7087 (N_7087,N_6874,N_6974);
and U7088 (N_7088,N_6911,N_6886);
nand U7089 (N_7089,N_6909,N_6801);
and U7090 (N_7090,N_6850,N_6895);
xnor U7091 (N_7091,N_6889,N_6825);
and U7092 (N_7092,N_6881,N_6972);
xor U7093 (N_7093,N_6883,N_6981);
nand U7094 (N_7094,N_6851,N_6829);
xnor U7095 (N_7095,N_6872,N_6941);
nand U7096 (N_7096,N_6913,N_6878);
nand U7097 (N_7097,N_6912,N_6956);
and U7098 (N_7098,N_6975,N_6837);
and U7099 (N_7099,N_6820,N_6997);
or U7100 (N_7100,N_6979,N_6986);
nand U7101 (N_7101,N_6995,N_6911);
or U7102 (N_7102,N_6923,N_6932);
or U7103 (N_7103,N_6860,N_6992);
or U7104 (N_7104,N_6984,N_6844);
and U7105 (N_7105,N_6867,N_6968);
and U7106 (N_7106,N_6870,N_6882);
and U7107 (N_7107,N_6911,N_6824);
nand U7108 (N_7108,N_6962,N_6933);
nor U7109 (N_7109,N_6977,N_6885);
xnor U7110 (N_7110,N_6813,N_6886);
nand U7111 (N_7111,N_6876,N_6953);
nor U7112 (N_7112,N_6912,N_6847);
xor U7113 (N_7113,N_6884,N_6944);
nand U7114 (N_7114,N_6910,N_6966);
nand U7115 (N_7115,N_6948,N_6973);
xor U7116 (N_7116,N_6880,N_6872);
and U7117 (N_7117,N_6927,N_6957);
xnor U7118 (N_7118,N_6844,N_6895);
nor U7119 (N_7119,N_6893,N_6807);
and U7120 (N_7120,N_6817,N_6805);
nor U7121 (N_7121,N_6993,N_6948);
nor U7122 (N_7122,N_6954,N_6834);
xor U7123 (N_7123,N_6810,N_6952);
and U7124 (N_7124,N_6814,N_6971);
or U7125 (N_7125,N_6930,N_6943);
or U7126 (N_7126,N_6887,N_6805);
and U7127 (N_7127,N_6893,N_6860);
nor U7128 (N_7128,N_6966,N_6862);
or U7129 (N_7129,N_6836,N_6919);
nand U7130 (N_7130,N_6902,N_6964);
nor U7131 (N_7131,N_6890,N_6836);
and U7132 (N_7132,N_6832,N_6810);
xor U7133 (N_7133,N_6984,N_6836);
nand U7134 (N_7134,N_6909,N_6905);
nand U7135 (N_7135,N_6946,N_6903);
and U7136 (N_7136,N_6923,N_6882);
or U7137 (N_7137,N_6960,N_6830);
nand U7138 (N_7138,N_6906,N_6959);
xor U7139 (N_7139,N_6889,N_6826);
nor U7140 (N_7140,N_6819,N_6960);
nand U7141 (N_7141,N_6915,N_6842);
and U7142 (N_7142,N_6948,N_6934);
or U7143 (N_7143,N_6801,N_6882);
xnor U7144 (N_7144,N_6837,N_6962);
and U7145 (N_7145,N_6979,N_6815);
or U7146 (N_7146,N_6924,N_6926);
and U7147 (N_7147,N_6931,N_6861);
nand U7148 (N_7148,N_6826,N_6848);
nand U7149 (N_7149,N_6858,N_6888);
and U7150 (N_7150,N_6915,N_6810);
nor U7151 (N_7151,N_6967,N_6872);
nand U7152 (N_7152,N_6835,N_6877);
or U7153 (N_7153,N_6851,N_6895);
and U7154 (N_7154,N_6840,N_6990);
or U7155 (N_7155,N_6925,N_6975);
or U7156 (N_7156,N_6869,N_6960);
nand U7157 (N_7157,N_6927,N_6955);
xor U7158 (N_7158,N_6988,N_6954);
nor U7159 (N_7159,N_6977,N_6936);
xnor U7160 (N_7160,N_6831,N_6822);
nor U7161 (N_7161,N_6928,N_6910);
xor U7162 (N_7162,N_6821,N_6846);
xor U7163 (N_7163,N_6810,N_6984);
xor U7164 (N_7164,N_6941,N_6983);
or U7165 (N_7165,N_6978,N_6923);
xnor U7166 (N_7166,N_6971,N_6861);
nor U7167 (N_7167,N_6859,N_6881);
xnor U7168 (N_7168,N_6855,N_6958);
and U7169 (N_7169,N_6850,N_6829);
nor U7170 (N_7170,N_6901,N_6819);
or U7171 (N_7171,N_6976,N_6991);
and U7172 (N_7172,N_6839,N_6992);
nand U7173 (N_7173,N_6920,N_6911);
nand U7174 (N_7174,N_6938,N_6823);
and U7175 (N_7175,N_6875,N_6828);
nor U7176 (N_7176,N_6881,N_6994);
xor U7177 (N_7177,N_6832,N_6835);
xnor U7178 (N_7178,N_6904,N_6974);
nor U7179 (N_7179,N_6863,N_6898);
nor U7180 (N_7180,N_6929,N_6973);
nand U7181 (N_7181,N_6924,N_6901);
or U7182 (N_7182,N_6960,N_6964);
nor U7183 (N_7183,N_6881,N_6860);
xor U7184 (N_7184,N_6939,N_6863);
nor U7185 (N_7185,N_6863,N_6855);
xnor U7186 (N_7186,N_6836,N_6929);
nor U7187 (N_7187,N_6903,N_6937);
and U7188 (N_7188,N_6825,N_6944);
nand U7189 (N_7189,N_6824,N_6809);
or U7190 (N_7190,N_6970,N_6830);
xnor U7191 (N_7191,N_6910,N_6957);
xor U7192 (N_7192,N_6924,N_6870);
and U7193 (N_7193,N_6936,N_6967);
or U7194 (N_7194,N_6980,N_6830);
nand U7195 (N_7195,N_6997,N_6907);
or U7196 (N_7196,N_6948,N_6952);
nand U7197 (N_7197,N_6910,N_6983);
nor U7198 (N_7198,N_6880,N_6918);
xor U7199 (N_7199,N_6861,N_6966);
xnor U7200 (N_7200,N_7147,N_7179);
nand U7201 (N_7201,N_7092,N_7186);
nand U7202 (N_7202,N_7136,N_7075);
or U7203 (N_7203,N_7199,N_7053);
and U7204 (N_7204,N_7002,N_7120);
xnor U7205 (N_7205,N_7030,N_7168);
or U7206 (N_7206,N_7054,N_7141);
or U7207 (N_7207,N_7088,N_7081);
and U7208 (N_7208,N_7072,N_7145);
and U7209 (N_7209,N_7099,N_7027);
xor U7210 (N_7210,N_7070,N_7177);
nor U7211 (N_7211,N_7171,N_7071);
and U7212 (N_7212,N_7082,N_7011);
or U7213 (N_7213,N_7029,N_7163);
xnor U7214 (N_7214,N_7160,N_7013);
xor U7215 (N_7215,N_7045,N_7197);
or U7216 (N_7216,N_7127,N_7178);
or U7217 (N_7217,N_7109,N_7134);
and U7218 (N_7218,N_7187,N_7084);
nand U7219 (N_7219,N_7114,N_7161);
nand U7220 (N_7220,N_7009,N_7050);
nor U7221 (N_7221,N_7035,N_7198);
nor U7222 (N_7222,N_7062,N_7043);
or U7223 (N_7223,N_7193,N_7005);
nand U7224 (N_7224,N_7181,N_7041);
nand U7225 (N_7225,N_7155,N_7176);
or U7226 (N_7226,N_7023,N_7060);
nor U7227 (N_7227,N_7128,N_7095);
or U7228 (N_7228,N_7015,N_7090);
nand U7229 (N_7229,N_7059,N_7056);
and U7230 (N_7230,N_7113,N_7103);
nor U7231 (N_7231,N_7138,N_7052);
and U7232 (N_7232,N_7094,N_7026);
xnor U7233 (N_7233,N_7042,N_7164);
and U7234 (N_7234,N_7038,N_7018);
nor U7235 (N_7235,N_7058,N_7121);
xnor U7236 (N_7236,N_7125,N_7012);
nor U7237 (N_7237,N_7174,N_7152);
nor U7238 (N_7238,N_7000,N_7061);
nor U7239 (N_7239,N_7157,N_7089);
and U7240 (N_7240,N_7185,N_7016);
nand U7241 (N_7241,N_7022,N_7007);
or U7242 (N_7242,N_7166,N_7020);
and U7243 (N_7243,N_7087,N_7083);
xnor U7244 (N_7244,N_7182,N_7001);
and U7245 (N_7245,N_7107,N_7024);
and U7246 (N_7246,N_7133,N_7137);
xor U7247 (N_7247,N_7017,N_7108);
or U7248 (N_7248,N_7057,N_7142);
nand U7249 (N_7249,N_7014,N_7190);
or U7250 (N_7250,N_7055,N_7115);
nor U7251 (N_7251,N_7135,N_7093);
nand U7252 (N_7252,N_7032,N_7124);
and U7253 (N_7253,N_7149,N_7008);
and U7254 (N_7254,N_7167,N_7144);
xnor U7255 (N_7255,N_7086,N_7188);
nor U7256 (N_7256,N_7119,N_7006);
or U7257 (N_7257,N_7080,N_7037);
and U7258 (N_7258,N_7154,N_7079);
xnor U7259 (N_7259,N_7194,N_7195);
or U7260 (N_7260,N_7047,N_7048);
or U7261 (N_7261,N_7078,N_7076);
or U7262 (N_7262,N_7189,N_7126);
nor U7263 (N_7263,N_7021,N_7158);
nor U7264 (N_7264,N_7116,N_7146);
and U7265 (N_7265,N_7097,N_7196);
xor U7266 (N_7266,N_7104,N_7064);
and U7267 (N_7267,N_7173,N_7051);
nor U7268 (N_7268,N_7156,N_7153);
xnor U7269 (N_7269,N_7067,N_7003);
nand U7270 (N_7270,N_7112,N_7025);
and U7271 (N_7271,N_7192,N_7098);
nand U7272 (N_7272,N_7165,N_7085);
xnor U7273 (N_7273,N_7034,N_7184);
xnor U7274 (N_7274,N_7073,N_7139);
xnor U7275 (N_7275,N_7004,N_7159);
nor U7276 (N_7276,N_7091,N_7183);
and U7277 (N_7277,N_7031,N_7132);
nor U7278 (N_7278,N_7111,N_7151);
nand U7279 (N_7279,N_7191,N_7150);
or U7280 (N_7280,N_7180,N_7096);
xnor U7281 (N_7281,N_7033,N_7129);
nand U7282 (N_7282,N_7019,N_7068);
or U7283 (N_7283,N_7123,N_7131);
or U7284 (N_7284,N_7100,N_7117);
nor U7285 (N_7285,N_7118,N_7143);
and U7286 (N_7286,N_7077,N_7172);
nand U7287 (N_7287,N_7074,N_7148);
xnor U7288 (N_7288,N_7162,N_7122);
or U7289 (N_7289,N_7049,N_7102);
nor U7290 (N_7290,N_7175,N_7040);
nor U7291 (N_7291,N_7066,N_7065);
nand U7292 (N_7292,N_7028,N_7110);
or U7293 (N_7293,N_7169,N_7106);
or U7294 (N_7294,N_7130,N_7140);
and U7295 (N_7295,N_7046,N_7069);
or U7296 (N_7296,N_7105,N_7170);
nor U7297 (N_7297,N_7036,N_7039);
nand U7298 (N_7298,N_7063,N_7101);
xor U7299 (N_7299,N_7044,N_7010);
nand U7300 (N_7300,N_7007,N_7103);
and U7301 (N_7301,N_7051,N_7084);
nor U7302 (N_7302,N_7140,N_7122);
nor U7303 (N_7303,N_7118,N_7055);
xor U7304 (N_7304,N_7190,N_7196);
xor U7305 (N_7305,N_7016,N_7192);
and U7306 (N_7306,N_7086,N_7101);
xnor U7307 (N_7307,N_7018,N_7172);
and U7308 (N_7308,N_7106,N_7109);
nor U7309 (N_7309,N_7034,N_7166);
xnor U7310 (N_7310,N_7125,N_7105);
or U7311 (N_7311,N_7184,N_7176);
nand U7312 (N_7312,N_7163,N_7077);
xnor U7313 (N_7313,N_7133,N_7040);
nor U7314 (N_7314,N_7082,N_7193);
nand U7315 (N_7315,N_7134,N_7117);
and U7316 (N_7316,N_7051,N_7148);
or U7317 (N_7317,N_7030,N_7109);
nand U7318 (N_7318,N_7112,N_7198);
and U7319 (N_7319,N_7092,N_7173);
nor U7320 (N_7320,N_7120,N_7027);
and U7321 (N_7321,N_7133,N_7199);
or U7322 (N_7322,N_7148,N_7139);
and U7323 (N_7323,N_7117,N_7102);
xnor U7324 (N_7324,N_7065,N_7129);
and U7325 (N_7325,N_7059,N_7062);
or U7326 (N_7326,N_7029,N_7169);
nand U7327 (N_7327,N_7117,N_7120);
and U7328 (N_7328,N_7058,N_7074);
and U7329 (N_7329,N_7102,N_7183);
nand U7330 (N_7330,N_7011,N_7125);
or U7331 (N_7331,N_7119,N_7136);
nand U7332 (N_7332,N_7146,N_7057);
xor U7333 (N_7333,N_7108,N_7080);
xnor U7334 (N_7334,N_7044,N_7047);
xnor U7335 (N_7335,N_7036,N_7195);
or U7336 (N_7336,N_7002,N_7173);
and U7337 (N_7337,N_7020,N_7133);
nand U7338 (N_7338,N_7198,N_7158);
or U7339 (N_7339,N_7013,N_7158);
nand U7340 (N_7340,N_7020,N_7034);
or U7341 (N_7341,N_7181,N_7045);
and U7342 (N_7342,N_7049,N_7157);
xnor U7343 (N_7343,N_7186,N_7086);
and U7344 (N_7344,N_7093,N_7009);
or U7345 (N_7345,N_7181,N_7080);
nand U7346 (N_7346,N_7048,N_7193);
nand U7347 (N_7347,N_7051,N_7032);
xnor U7348 (N_7348,N_7122,N_7152);
nor U7349 (N_7349,N_7029,N_7076);
or U7350 (N_7350,N_7189,N_7171);
or U7351 (N_7351,N_7171,N_7023);
xnor U7352 (N_7352,N_7160,N_7006);
nand U7353 (N_7353,N_7125,N_7020);
nor U7354 (N_7354,N_7198,N_7191);
nor U7355 (N_7355,N_7141,N_7178);
nand U7356 (N_7356,N_7015,N_7128);
or U7357 (N_7357,N_7113,N_7159);
nor U7358 (N_7358,N_7189,N_7012);
and U7359 (N_7359,N_7027,N_7028);
and U7360 (N_7360,N_7071,N_7045);
or U7361 (N_7361,N_7055,N_7129);
xor U7362 (N_7362,N_7071,N_7081);
or U7363 (N_7363,N_7088,N_7135);
xnor U7364 (N_7364,N_7036,N_7042);
or U7365 (N_7365,N_7034,N_7159);
nor U7366 (N_7366,N_7144,N_7050);
nor U7367 (N_7367,N_7173,N_7072);
or U7368 (N_7368,N_7155,N_7067);
xor U7369 (N_7369,N_7049,N_7084);
nand U7370 (N_7370,N_7000,N_7112);
and U7371 (N_7371,N_7135,N_7074);
nor U7372 (N_7372,N_7157,N_7181);
and U7373 (N_7373,N_7154,N_7042);
xnor U7374 (N_7374,N_7156,N_7023);
nand U7375 (N_7375,N_7139,N_7143);
xor U7376 (N_7376,N_7103,N_7017);
or U7377 (N_7377,N_7181,N_7091);
or U7378 (N_7378,N_7181,N_7088);
xor U7379 (N_7379,N_7115,N_7059);
or U7380 (N_7380,N_7131,N_7052);
and U7381 (N_7381,N_7065,N_7047);
and U7382 (N_7382,N_7040,N_7132);
xnor U7383 (N_7383,N_7131,N_7137);
or U7384 (N_7384,N_7020,N_7139);
xor U7385 (N_7385,N_7170,N_7181);
nand U7386 (N_7386,N_7151,N_7080);
xnor U7387 (N_7387,N_7021,N_7028);
nor U7388 (N_7388,N_7087,N_7179);
or U7389 (N_7389,N_7108,N_7096);
xor U7390 (N_7390,N_7108,N_7180);
and U7391 (N_7391,N_7127,N_7009);
and U7392 (N_7392,N_7138,N_7104);
nor U7393 (N_7393,N_7137,N_7192);
and U7394 (N_7394,N_7101,N_7137);
nor U7395 (N_7395,N_7106,N_7137);
xor U7396 (N_7396,N_7028,N_7046);
xor U7397 (N_7397,N_7087,N_7050);
xor U7398 (N_7398,N_7008,N_7066);
nand U7399 (N_7399,N_7033,N_7125);
nand U7400 (N_7400,N_7332,N_7303);
and U7401 (N_7401,N_7293,N_7216);
nor U7402 (N_7402,N_7242,N_7399);
and U7403 (N_7403,N_7215,N_7246);
xor U7404 (N_7404,N_7255,N_7367);
xnor U7405 (N_7405,N_7382,N_7254);
and U7406 (N_7406,N_7210,N_7366);
nand U7407 (N_7407,N_7395,N_7238);
nand U7408 (N_7408,N_7334,N_7387);
xnor U7409 (N_7409,N_7314,N_7225);
and U7410 (N_7410,N_7240,N_7282);
nor U7411 (N_7411,N_7275,N_7221);
xor U7412 (N_7412,N_7259,N_7381);
xor U7413 (N_7413,N_7209,N_7241);
nor U7414 (N_7414,N_7397,N_7388);
nand U7415 (N_7415,N_7355,N_7280);
and U7416 (N_7416,N_7260,N_7386);
nor U7417 (N_7417,N_7217,N_7219);
nor U7418 (N_7418,N_7318,N_7304);
nor U7419 (N_7419,N_7393,N_7291);
nor U7420 (N_7420,N_7272,N_7383);
xnor U7421 (N_7421,N_7268,N_7370);
or U7422 (N_7422,N_7317,N_7392);
or U7423 (N_7423,N_7305,N_7287);
and U7424 (N_7424,N_7294,N_7292);
or U7425 (N_7425,N_7265,N_7297);
nor U7426 (N_7426,N_7371,N_7389);
and U7427 (N_7427,N_7345,N_7251);
nor U7428 (N_7428,N_7234,N_7358);
xnor U7429 (N_7429,N_7247,N_7340);
xnor U7430 (N_7430,N_7273,N_7306);
nor U7431 (N_7431,N_7329,N_7351);
xor U7432 (N_7432,N_7203,N_7374);
xor U7433 (N_7433,N_7330,N_7361);
xor U7434 (N_7434,N_7249,N_7200);
nand U7435 (N_7435,N_7266,N_7201);
xor U7436 (N_7436,N_7245,N_7222);
and U7437 (N_7437,N_7220,N_7365);
or U7438 (N_7438,N_7325,N_7269);
or U7439 (N_7439,N_7341,N_7312);
nor U7440 (N_7440,N_7310,N_7313);
nand U7441 (N_7441,N_7253,N_7307);
nand U7442 (N_7442,N_7384,N_7333);
and U7443 (N_7443,N_7300,N_7232);
nor U7444 (N_7444,N_7349,N_7331);
xor U7445 (N_7445,N_7264,N_7327);
nor U7446 (N_7446,N_7237,N_7396);
and U7447 (N_7447,N_7343,N_7233);
or U7448 (N_7448,N_7230,N_7295);
xor U7449 (N_7449,N_7385,N_7398);
and U7450 (N_7450,N_7390,N_7218);
xnor U7451 (N_7451,N_7202,N_7243);
and U7452 (N_7452,N_7208,N_7350);
nand U7453 (N_7453,N_7336,N_7258);
and U7454 (N_7454,N_7286,N_7270);
or U7455 (N_7455,N_7356,N_7347);
nor U7456 (N_7456,N_7378,N_7223);
or U7457 (N_7457,N_7311,N_7373);
and U7458 (N_7458,N_7277,N_7267);
or U7459 (N_7459,N_7302,N_7360);
xnor U7460 (N_7460,N_7283,N_7346);
nor U7461 (N_7461,N_7364,N_7352);
and U7462 (N_7462,N_7298,N_7226);
or U7463 (N_7463,N_7379,N_7288);
nor U7464 (N_7464,N_7281,N_7284);
nand U7465 (N_7465,N_7368,N_7279);
nand U7466 (N_7466,N_7344,N_7362);
nand U7467 (N_7467,N_7227,N_7213);
nand U7468 (N_7468,N_7252,N_7316);
and U7469 (N_7469,N_7212,N_7359);
nor U7470 (N_7470,N_7262,N_7319);
and U7471 (N_7471,N_7231,N_7301);
xor U7472 (N_7472,N_7376,N_7348);
xor U7473 (N_7473,N_7235,N_7274);
and U7474 (N_7474,N_7375,N_7372);
xor U7475 (N_7475,N_7211,N_7257);
xnor U7476 (N_7476,N_7323,N_7309);
xnor U7477 (N_7477,N_7214,N_7320);
xnor U7478 (N_7478,N_7363,N_7357);
xor U7479 (N_7479,N_7289,N_7342);
xor U7480 (N_7480,N_7206,N_7321);
and U7481 (N_7481,N_7322,N_7244);
nor U7482 (N_7482,N_7377,N_7369);
xor U7483 (N_7483,N_7205,N_7339);
nor U7484 (N_7484,N_7394,N_7391);
xor U7485 (N_7485,N_7315,N_7224);
nand U7486 (N_7486,N_7263,N_7328);
nand U7487 (N_7487,N_7324,N_7271);
or U7488 (N_7488,N_7228,N_7290);
and U7489 (N_7489,N_7337,N_7250);
or U7490 (N_7490,N_7278,N_7285);
nor U7491 (N_7491,N_7326,N_7308);
or U7492 (N_7492,N_7204,N_7239);
nor U7493 (N_7493,N_7354,N_7248);
xnor U7494 (N_7494,N_7335,N_7296);
and U7495 (N_7495,N_7380,N_7207);
or U7496 (N_7496,N_7256,N_7276);
nor U7497 (N_7497,N_7338,N_7229);
nor U7498 (N_7498,N_7353,N_7261);
and U7499 (N_7499,N_7236,N_7299);
nand U7500 (N_7500,N_7258,N_7379);
xor U7501 (N_7501,N_7216,N_7362);
and U7502 (N_7502,N_7210,N_7263);
nor U7503 (N_7503,N_7235,N_7228);
and U7504 (N_7504,N_7392,N_7204);
nand U7505 (N_7505,N_7275,N_7386);
xor U7506 (N_7506,N_7238,N_7316);
or U7507 (N_7507,N_7301,N_7258);
xor U7508 (N_7508,N_7329,N_7299);
xnor U7509 (N_7509,N_7353,N_7229);
xnor U7510 (N_7510,N_7389,N_7358);
and U7511 (N_7511,N_7265,N_7302);
and U7512 (N_7512,N_7366,N_7333);
nor U7513 (N_7513,N_7302,N_7309);
or U7514 (N_7514,N_7377,N_7354);
xor U7515 (N_7515,N_7257,N_7320);
nor U7516 (N_7516,N_7283,N_7390);
nand U7517 (N_7517,N_7269,N_7263);
and U7518 (N_7518,N_7251,N_7260);
nor U7519 (N_7519,N_7343,N_7381);
nor U7520 (N_7520,N_7373,N_7278);
xnor U7521 (N_7521,N_7304,N_7227);
and U7522 (N_7522,N_7277,N_7295);
or U7523 (N_7523,N_7238,N_7257);
nand U7524 (N_7524,N_7384,N_7269);
or U7525 (N_7525,N_7385,N_7387);
and U7526 (N_7526,N_7397,N_7203);
nand U7527 (N_7527,N_7304,N_7389);
nand U7528 (N_7528,N_7380,N_7212);
nor U7529 (N_7529,N_7308,N_7335);
nand U7530 (N_7530,N_7241,N_7319);
nor U7531 (N_7531,N_7352,N_7237);
or U7532 (N_7532,N_7203,N_7276);
nand U7533 (N_7533,N_7315,N_7204);
and U7534 (N_7534,N_7265,N_7358);
nand U7535 (N_7535,N_7380,N_7344);
and U7536 (N_7536,N_7365,N_7212);
and U7537 (N_7537,N_7245,N_7269);
nor U7538 (N_7538,N_7237,N_7285);
and U7539 (N_7539,N_7358,N_7295);
xnor U7540 (N_7540,N_7395,N_7361);
or U7541 (N_7541,N_7214,N_7366);
nor U7542 (N_7542,N_7351,N_7280);
nand U7543 (N_7543,N_7276,N_7297);
nor U7544 (N_7544,N_7286,N_7243);
or U7545 (N_7545,N_7287,N_7215);
nand U7546 (N_7546,N_7350,N_7318);
nor U7547 (N_7547,N_7255,N_7209);
xor U7548 (N_7548,N_7245,N_7205);
or U7549 (N_7549,N_7325,N_7355);
nor U7550 (N_7550,N_7399,N_7369);
nand U7551 (N_7551,N_7348,N_7375);
nand U7552 (N_7552,N_7340,N_7389);
or U7553 (N_7553,N_7378,N_7336);
nor U7554 (N_7554,N_7325,N_7224);
nand U7555 (N_7555,N_7238,N_7335);
nand U7556 (N_7556,N_7245,N_7313);
nand U7557 (N_7557,N_7221,N_7281);
and U7558 (N_7558,N_7303,N_7372);
or U7559 (N_7559,N_7279,N_7223);
or U7560 (N_7560,N_7278,N_7346);
nand U7561 (N_7561,N_7347,N_7375);
nor U7562 (N_7562,N_7354,N_7297);
nand U7563 (N_7563,N_7252,N_7207);
nor U7564 (N_7564,N_7348,N_7306);
xnor U7565 (N_7565,N_7372,N_7210);
nand U7566 (N_7566,N_7384,N_7301);
nor U7567 (N_7567,N_7265,N_7295);
nand U7568 (N_7568,N_7399,N_7248);
nor U7569 (N_7569,N_7278,N_7317);
and U7570 (N_7570,N_7289,N_7236);
or U7571 (N_7571,N_7296,N_7275);
xor U7572 (N_7572,N_7323,N_7270);
nand U7573 (N_7573,N_7218,N_7352);
nor U7574 (N_7574,N_7292,N_7354);
and U7575 (N_7575,N_7357,N_7325);
nor U7576 (N_7576,N_7330,N_7347);
and U7577 (N_7577,N_7379,N_7250);
xnor U7578 (N_7578,N_7241,N_7207);
nand U7579 (N_7579,N_7318,N_7364);
or U7580 (N_7580,N_7225,N_7303);
or U7581 (N_7581,N_7214,N_7253);
or U7582 (N_7582,N_7250,N_7207);
nor U7583 (N_7583,N_7347,N_7313);
or U7584 (N_7584,N_7226,N_7268);
or U7585 (N_7585,N_7219,N_7234);
nand U7586 (N_7586,N_7275,N_7249);
xnor U7587 (N_7587,N_7398,N_7280);
nand U7588 (N_7588,N_7273,N_7222);
nor U7589 (N_7589,N_7384,N_7265);
nor U7590 (N_7590,N_7371,N_7395);
or U7591 (N_7591,N_7378,N_7213);
nor U7592 (N_7592,N_7290,N_7226);
nand U7593 (N_7593,N_7342,N_7354);
xnor U7594 (N_7594,N_7242,N_7362);
nor U7595 (N_7595,N_7204,N_7377);
nand U7596 (N_7596,N_7292,N_7301);
nand U7597 (N_7597,N_7311,N_7266);
xor U7598 (N_7598,N_7334,N_7225);
nor U7599 (N_7599,N_7213,N_7285);
xor U7600 (N_7600,N_7450,N_7531);
or U7601 (N_7601,N_7448,N_7523);
nor U7602 (N_7602,N_7473,N_7457);
and U7603 (N_7603,N_7479,N_7561);
nand U7604 (N_7604,N_7494,N_7516);
or U7605 (N_7605,N_7495,N_7486);
nor U7606 (N_7606,N_7560,N_7546);
xor U7607 (N_7607,N_7583,N_7466);
xnor U7608 (N_7608,N_7573,N_7585);
xor U7609 (N_7609,N_7528,N_7465);
or U7610 (N_7610,N_7496,N_7570);
and U7611 (N_7611,N_7504,N_7551);
xnor U7612 (N_7612,N_7521,N_7430);
xnor U7613 (N_7613,N_7499,N_7547);
nor U7614 (N_7614,N_7597,N_7468);
or U7615 (N_7615,N_7446,N_7431);
nand U7616 (N_7616,N_7580,N_7598);
nor U7617 (N_7617,N_7549,N_7405);
or U7618 (N_7618,N_7423,N_7595);
nand U7619 (N_7619,N_7437,N_7497);
xor U7620 (N_7620,N_7581,N_7480);
nand U7621 (N_7621,N_7487,N_7427);
nor U7622 (N_7622,N_7519,N_7433);
nor U7623 (N_7623,N_7471,N_7505);
or U7624 (N_7624,N_7532,N_7567);
nand U7625 (N_7625,N_7447,N_7591);
xor U7626 (N_7626,N_7540,N_7436);
or U7627 (N_7627,N_7449,N_7593);
nand U7628 (N_7628,N_7445,N_7484);
xnor U7629 (N_7629,N_7439,N_7441);
xor U7630 (N_7630,N_7525,N_7482);
nand U7631 (N_7631,N_7403,N_7550);
or U7632 (N_7632,N_7488,N_7510);
or U7633 (N_7633,N_7442,N_7438);
xnor U7634 (N_7634,N_7464,N_7563);
or U7635 (N_7635,N_7422,N_7556);
or U7636 (N_7636,N_7420,N_7416);
or U7637 (N_7637,N_7534,N_7490);
xor U7638 (N_7638,N_7564,N_7460);
nor U7639 (N_7639,N_7548,N_7467);
xnor U7640 (N_7640,N_7415,N_7409);
or U7641 (N_7641,N_7493,N_7404);
nor U7642 (N_7642,N_7435,N_7535);
xor U7643 (N_7643,N_7545,N_7407);
nand U7644 (N_7644,N_7424,N_7577);
nand U7645 (N_7645,N_7524,N_7578);
nand U7646 (N_7646,N_7558,N_7518);
nand U7647 (N_7647,N_7414,N_7584);
xnor U7648 (N_7648,N_7477,N_7429);
nor U7649 (N_7649,N_7472,N_7470);
or U7650 (N_7650,N_7411,N_7553);
and U7651 (N_7651,N_7542,N_7544);
and U7652 (N_7652,N_7508,N_7569);
or U7653 (N_7653,N_7541,N_7555);
and U7654 (N_7654,N_7453,N_7461);
xnor U7655 (N_7655,N_7506,N_7458);
and U7656 (N_7656,N_7452,N_7582);
and U7657 (N_7657,N_7513,N_7594);
nor U7658 (N_7658,N_7419,N_7515);
nor U7659 (N_7659,N_7512,N_7522);
xnor U7660 (N_7660,N_7574,N_7443);
and U7661 (N_7661,N_7434,N_7589);
nand U7662 (N_7662,N_7451,N_7440);
and U7663 (N_7663,N_7408,N_7417);
nand U7664 (N_7664,N_7539,N_7554);
xor U7665 (N_7665,N_7410,N_7456);
nand U7666 (N_7666,N_7402,N_7463);
or U7667 (N_7667,N_7432,N_7588);
nor U7668 (N_7668,N_7418,N_7559);
and U7669 (N_7669,N_7529,N_7489);
nand U7670 (N_7670,N_7517,N_7509);
and U7671 (N_7671,N_7485,N_7511);
nand U7672 (N_7672,N_7575,N_7562);
nand U7673 (N_7673,N_7413,N_7428);
nand U7674 (N_7674,N_7478,N_7503);
nor U7675 (N_7675,N_7572,N_7502);
xnor U7676 (N_7676,N_7527,N_7536);
nand U7677 (N_7677,N_7520,N_7552);
xnor U7678 (N_7678,N_7590,N_7426);
or U7679 (N_7679,N_7474,N_7530);
nand U7680 (N_7680,N_7459,N_7421);
or U7681 (N_7681,N_7491,N_7401);
xnor U7682 (N_7682,N_7514,N_7576);
xnor U7683 (N_7683,N_7492,N_7425);
xnor U7684 (N_7684,N_7586,N_7475);
xnor U7685 (N_7685,N_7526,N_7483);
nand U7686 (N_7686,N_7455,N_7444);
xnor U7687 (N_7687,N_7462,N_7476);
or U7688 (N_7688,N_7533,N_7557);
and U7689 (N_7689,N_7596,N_7406);
or U7690 (N_7690,N_7537,N_7454);
xnor U7691 (N_7691,N_7566,N_7571);
or U7692 (N_7692,N_7469,N_7543);
xnor U7693 (N_7693,N_7498,N_7507);
or U7694 (N_7694,N_7579,N_7481);
nor U7695 (N_7695,N_7592,N_7587);
nand U7696 (N_7696,N_7412,N_7599);
and U7697 (N_7697,N_7568,N_7400);
nor U7698 (N_7698,N_7501,N_7565);
or U7699 (N_7699,N_7538,N_7500);
or U7700 (N_7700,N_7461,N_7507);
xor U7701 (N_7701,N_7599,N_7478);
and U7702 (N_7702,N_7457,N_7539);
nor U7703 (N_7703,N_7560,N_7487);
nor U7704 (N_7704,N_7555,N_7463);
and U7705 (N_7705,N_7516,N_7416);
nor U7706 (N_7706,N_7520,N_7579);
and U7707 (N_7707,N_7414,N_7494);
or U7708 (N_7708,N_7574,N_7523);
nand U7709 (N_7709,N_7557,N_7445);
and U7710 (N_7710,N_7415,N_7493);
xnor U7711 (N_7711,N_7571,N_7510);
nand U7712 (N_7712,N_7408,N_7557);
or U7713 (N_7713,N_7425,N_7421);
xnor U7714 (N_7714,N_7474,N_7439);
and U7715 (N_7715,N_7467,N_7569);
nand U7716 (N_7716,N_7509,N_7488);
or U7717 (N_7717,N_7462,N_7417);
and U7718 (N_7718,N_7536,N_7520);
xnor U7719 (N_7719,N_7455,N_7422);
nand U7720 (N_7720,N_7594,N_7572);
or U7721 (N_7721,N_7562,N_7459);
or U7722 (N_7722,N_7508,N_7408);
nand U7723 (N_7723,N_7444,N_7435);
or U7724 (N_7724,N_7460,N_7471);
nor U7725 (N_7725,N_7422,N_7503);
nand U7726 (N_7726,N_7549,N_7495);
xor U7727 (N_7727,N_7409,N_7502);
nor U7728 (N_7728,N_7462,N_7583);
nor U7729 (N_7729,N_7537,N_7434);
or U7730 (N_7730,N_7442,N_7529);
nor U7731 (N_7731,N_7410,N_7573);
xor U7732 (N_7732,N_7450,N_7448);
xor U7733 (N_7733,N_7581,N_7431);
xnor U7734 (N_7734,N_7449,N_7573);
nand U7735 (N_7735,N_7492,N_7431);
nand U7736 (N_7736,N_7459,N_7412);
or U7737 (N_7737,N_7409,N_7462);
and U7738 (N_7738,N_7472,N_7495);
nor U7739 (N_7739,N_7413,N_7432);
nor U7740 (N_7740,N_7596,N_7462);
nand U7741 (N_7741,N_7570,N_7557);
nand U7742 (N_7742,N_7570,N_7447);
and U7743 (N_7743,N_7460,N_7544);
and U7744 (N_7744,N_7586,N_7502);
or U7745 (N_7745,N_7536,N_7451);
nor U7746 (N_7746,N_7405,N_7547);
nand U7747 (N_7747,N_7435,N_7427);
nor U7748 (N_7748,N_7440,N_7495);
nand U7749 (N_7749,N_7527,N_7579);
xnor U7750 (N_7750,N_7509,N_7598);
or U7751 (N_7751,N_7557,N_7510);
xor U7752 (N_7752,N_7564,N_7500);
xnor U7753 (N_7753,N_7424,N_7545);
nor U7754 (N_7754,N_7532,N_7594);
xor U7755 (N_7755,N_7405,N_7491);
xnor U7756 (N_7756,N_7475,N_7415);
xor U7757 (N_7757,N_7463,N_7497);
xor U7758 (N_7758,N_7578,N_7521);
and U7759 (N_7759,N_7418,N_7504);
nor U7760 (N_7760,N_7553,N_7583);
and U7761 (N_7761,N_7475,N_7486);
nand U7762 (N_7762,N_7522,N_7410);
or U7763 (N_7763,N_7559,N_7531);
nand U7764 (N_7764,N_7514,N_7555);
or U7765 (N_7765,N_7496,N_7566);
or U7766 (N_7766,N_7495,N_7503);
xor U7767 (N_7767,N_7491,N_7559);
or U7768 (N_7768,N_7422,N_7498);
and U7769 (N_7769,N_7599,N_7584);
nand U7770 (N_7770,N_7513,N_7503);
xor U7771 (N_7771,N_7584,N_7492);
nand U7772 (N_7772,N_7407,N_7506);
nand U7773 (N_7773,N_7526,N_7465);
or U7774 (N_7774,N_7414,N_7530);
or U7775 (N_7775,N_7580,N_7455);
xnor U7776 (N_7776,N_7520,N_7587);
nor U7777 (N_7777,N_7554,N_7462);
or U7778 (N_7778,N_7511,N_7510);
xor U7779 (N_7779,N_7448,N_7438);
and U7780 (N_7780,N_7596,N_7407);
and U7781 (N_7781,N_7412,N_7563);
or U7782 (N_7782,N_7508,N_7513);
and U7783 (N_7783,N_7447,N_7470);
and U7784 (N_7784,N_7413,N_7594);
xnor U7785 (N_7785,N_7421,N_7535);
xnor U7786 (N_7786,N_7460,N_7419);
nand U7787 (N_7787,N_7467,N_7553);
nor U7788 (N_7788,N_7519,N_7524);
nor U7789 (N_7789,N_7511,N_7568);
nand U7790 (N_7790,N_7584,N_7526);
nor U7791 (N_7791,N_7582,N_7527);
or U7792 (N_7792,N_7597,N_7426);
nand U7793 (N_7793,N_7492,N_7467);
xnor U7794 (N_7794,N_7556,N_7416);
nor U7795 (N_7795,N_7482,N_7533);
and U7796 (N_7796,N_7435,N_7570);
or U7797 (N_7797,N_7577,N_7430);
nor U7798 (N_7798,N_7431,N_7437);
or U7799 (N_7799,N_7407,N_7406);
nor U7800 (N_7800,N_7792,N_7603);
xor U7801 (N_7801,N_7759,N_7726);
or U7802 (N_7802,N_7740,N_7743);
nor U7803 (N_7803,N_7728,N_7748);
or U7804 (N_7804,N_7765,N_7669);
nand U7805 (N_7805,N_7732,N_7701);
and U7806 (N_7806,N_7786,N_7653);
and U7807 (N_7807,N_7737,N_7711);
nor U7808 (N_7808,N_7727,N_7641);
xnor U7809 (N_7809,N_7686,N_7793);
xor U7810 (N_7810,N_7702,N_7689);
or U7811 (N_7811,N_7601,N_7657);
xor U7812 (N_7812,N_7720,N_7630);
nor U7813 (N_7813,N_7623,N_7618);
nand U7814 (N_7814,N_7662,N_7738);
or U7815 (N_7815,N_7664,N_7712);
nand U7816 (N_7816,N_7672,N_7692);
or U7817 (N_7817,N_7767,N_7665);
nor U7818 (N_7818,N_7721,N_7744);
xnor U7819 (N_7819,N_7784,N_7687);
nand U7820 (N_7820,N_7602,N_7753);
and U7821 (N_7821,N_7619,N_7627);
nand U7822 (N_7822,N_7681,N_7787);
xor U7823 (N_7823,N_7696,N_7610);
nor U7824 (N_7824,N_7659,N_7782);
xor U7825 (N_7825,N_7683,N_7690);
nor U7826 (N_7826,N_7779,N_7663);
xnor U7827 (N_7827,N_7635,N_7795);
nand U7828 (N_7828,N_7629,N_7661);
or U7829 (N_7829,N_7673,N_7745);
and U7830 (N_7830,N_7706,N_7785);
nand U7831 (N_7831,N_7707,N_7719);
xnor U7832 (N_7832,N_7718,N_7791);
and U7833 (N_7833,N_7652,N_7632);
nor U7834 (N_7834,N_7723,N_7647);
and U7835 (N_7835,N_7611,N_7671);
nand U7836 (N_7836,N_7695,N_7656);
nor U7837 (N_7837,N_7644,N_7796);
and U7838 (N_7838,N_7774,N_7691);
nor U7839 (N_7839,N_7639,N_7797);
or U7840 (N_7840,N_7607,N_7633);
nor U7841 (N_7841,N_7654,N_7788);
or U7842 (N_7842,N_7735,N_7693);
xnor U7843 (N_7843,N_7668,N_7608);
or U7844 (N_7844,N_7651,N_7645);
xor U7845 (N_7845,N_7667,N_7747);
or U7846 (N_7846,N_7688,N_7617);
xor U7847 (N_7847,N_7698,N_7799);
or U7848 (N_7848,N_7642,N_7600);
nand U7849 (N_7849,N_7604,N_7798);
and U7850 (N_7850,N_7631,N_7697);
xnor U7851 (N_7851,N_7708,N_7622);
nor U7852 (N_7852,N_7620,N_7679);
xor U7853 (N_7853,N_7762,N_7624);
nand U7854 (N_7854,N_7704,N_7746);
nand U7855 (N_7855,N_7715,N_7714);
xor U7856 (N_7856,N_7703,N_7724);
nand U7857 (N_7857,N_7677,N_7612);
nor U7858 (N_7858,N_7769,N_7768);
xnor U7859 (N_7859,N_7621,N_7650);
xor U7860 (N_7860,N_7694,N_7754);
or U7861 (N_7861,N_7626,N_7648);
nor U7862 (N_7862,N_7783,N_7773);
and U7863 (N_7863,N_7615,N_7638);
xor U7864 (N_7864,N_7705,N_7709);
xnor U7865 (N_7865,N_7757,N_7684);
or U7866 (N_7866,N_7640,N_7780);
xor U7867 (N_7867,N_7678,N_7625);
nor U7868 (N_7868,N_7674,N_7771);
and U7869 (N_7869,N_7751,N_7794);
and U7870 (N_7870,N_7734,N_7658);
nor U7871 (N_7871,N_7676,N_7750);
and U7872 (N_7872,N_7606,N_7646);
xnor U7873 (N_7873,N_7613,N_7731);
nand U7874 (N_7874,N_7713,N_7700);
or U7875 (N_7875,N_7733,N_7699);
nand U7876 (N_7876,N_7634,N_7605);
or U7877 (N_7877,N_7790,N_7761);
or U7878 (N_7878,N_7758,N_7756);
or U7879 (N_7879,N_7643,N_7682);
nor U7880 (N_7880,N_7725,N_7755);
nor U7881 (N_7881,N_7775,N_7770);
nand U7882 (N_7882,N_7636,N_7742);
nor U7883 (N_7883,N_7628,N_7739);
nor U7884 (N_7884,N_7717,N_7729);
xnor U7885 (N_7885,N_7789,N_7763);
and U7886 (N_7886,N_7649,N_7776);
nand U7887 (N_7887,N_7616,N_7675);
nor U7888 (N_7888,N_7614,N_7670);
xor U7889 (N_7889,N_7710,N_7736);
or U7890 (N_7890,N_7764,N_7760);
or U7891 (N_7891,N_7766,N_7655);
xor U7892 (N_7892,N_7752,N_7722);
and U7893 (N_7893,N_7772,N_7680);
xnor U7894 (N_7894,N_7730,N_7749);
nor U7895 (N_7895,N_7716,N_7660);
nor U7896 (N_7896,N_7778,N_7685);
and U7897 (N_7897,N_7741,N_7777);
or U7898 (N_7898,N_7666,N_7637);
xnor U7899 (N_7899,N_7781,N_7609);
nor U7900 (N_7900,N_7641,N_7604);
or U7901 (N_7901,N_7650,N_7788);
xnor U7902 (N_7902,N_7643,N_7764);
nand U7903 (N_7903,N_7660,N_7680);
nor U7904 (N_7904,N_7683,N_7620);
xor U7905 (N_7905,N_7662,N_7759);
nor U7906 (N_7906,N_7625,N_7734);
or U7907 (N_7907,N_7779,N_7640);
and U7908 (N_7908,N_7642,N_7748);
or U7909 (N_7909,N_7652,N_7659);
xnor U7910 (N_7910,N_7661,N_7777);
xnor U7911 (N_7911,N_7649,N_7702);
xor U7912 (N_7912,N_7669,N_7664);
or U7913 (N_7913,N_7683,N_7710);
or U7914 (N_7914,N_7644,N_7763);
and U7915 (N_7915,N_7657,N_7632);
and U7916 (N_7916,N_7714,N_7639);
nor U7917 (N_7917,N_7794,N_7795);
nor U7918 (N_7918,N_7654,N_7712);
or U7919 (N_7919,N_7779,N_7659);
nor U7920 (N_7920,N_7606,N_7632);
or U7921 (N_7921,N_7708,N_7712);
nand U7922 (N_7922,N_7624,N_7675);
xnor U7923 (N_7923,N_7645,N_7638);
and U7924 (N_7924,N_7621,N_7715);
xnor U7925 (N_7925,N_7793,N_7722);
or U7926 (N_7926,N_7781,N_7724);
and U7927 (N_7927,N_7754,N_7675);
nand U7928 (N_7928,N_7663,N_7696);
xnor U7929 (N_7929,N_7795,N_7608);
xor U7930 (N_7930,N_7752,N_7711);
nor U7931 (N_7931,N_7657,N_7651);
or U7932 (N_7932,N_7726,N_7637);
nor U7933 (N_7933,N_7633,N_7761);
xor U7934 (N_7934,N_7689,N_7735);
nor U7935 (N_7935,N_7774,N_7696);
xor U7936 (N_7936,N_7608,N_7632);
xor U7937 (N_7937,N_7702,N_7782);
or U7938 (N_7938,N_7724,N_7708);
and U7939 (N_7939,N_7636,N_7669);
nor U7940 (N_7940,N_7653,N_7658);
nor U7941 (N_7941,N_7644,N_7606);
nand U7942 (N_7942,N_7674,N_7783);
or U7943 (N_7943,N_7683,N_7779);
nand U7944 (N_7944,N_7791,N_7617);
or U7945 (N_7945,N_7765,N_7610);
or U7946 (N_7946,N_7631,N_7621);
and U7947 (N_7947,N_7668,N_7601);
nor U7948 (N_7948,N_7650,N_7734);
nor U7949 (N_7949,N_7792,N_7747);
nor U7950 (N_7950,N_7607,N_7725);
xor U7951 (N_7951,N_7764,N_7644);
and U7952 (N_7952,N_7674,N_7796);
nand U7953 (N_7953,N_7707,N_7772);
or U7954 (N_7954,N_7778,N_7604);
or U7955 (N_7955,N_7604,N_7756);
nor U7956 (N_7956,N_7770,N_7616);
and U7957 (N_7957,N_7719,N_7731);
and U7958 (N_7958,N_7630,N_7698);
and U7959 (N_7959,N_7797,N_7763);
and U7960 (N_7960,N_7729,N_7793);
and U7961 (N_7961,N_7779,N_7607);
nor U7962 (N_7962,N_7779,N_7766);
or U7963 (N_7963,N_7754,N_7676);
nand U7964 (N_7964,N_7637,N_7633);
and U7965 (N_7965,N_7614,N_7769);
xnor U7966 (N_7966,N_7721,N_7692);
or U7967 (N_7967,N_7723,N_7629);
nor U7968 (N_7968,N_7657,N_7733);
nor U7969 (N_7969,N_7617,N_7694);
and U7970 (N_7970,N_7793,N_7718);
nand U7971 (N_7971,N_7622,N_7722);
or U7972 (N_7972,N_7676,N_7685);
xnor U7973 (N_7973,N_7606,N_7663);
xor U7974 (N_7974,N_7650,N_7696);
xor U7975 (N_7975,N_7657,N_7719);
nand U7976 (N_7976,N_7691,N_7653);
or U7977 (N_7977,N_7743,N_7651);
nand U7978 (N_7978,N_7627,N_7673);
and U7979 (N_7979,N_7664,N_7746);
and U7980 (N_7980,N_7757,N_7719);
or U7981 (N_7981,N_7793,N_7697);
or U7982 (N_7982,N_7771,N_7797);
xor U7983 (N_7983,N_7663,N_7677);
xor U7984 (N_7984,N_7658,N_7750);
or U7985 (N_7985,N_7648,N_7671);
and U7986 (N_7986,N_7628,N_7649);
nand U7987 (N_7987,N_7791,N_7623);
nand U7988 (N_7988,N_7722,N_7666);
and U7989 (N_7989,N_7648,N_7654);
xor U7990 (N_7990,N_7627,N_7775);
nand U7991 (N_7991,N_7797,N_7675);
nor U7992 (N_7992,N_7678,N_7607);
nor U7993 (N_7993,N_7617,N_7716);
nor U7994 (N_7994,N_7626,N_7603);
nor U7995 (N_7995,N_7781,N_7744);
or U7996 (N_7996,N_7737,N_7709);
nand U7997 (N_7997,N_7727,N_7674);
nand U7998 (N_7998,N_7771,N_7799);
and U7999 (N_7999,N_7614,N_7780);
nand U8000 (N_8000,N_7992,N_7850);
nand U8001 (N_8001,N_7990,N_7802);
or U8002 (N_8002,N_7954,N_7997);
or U8003 (N_8003,N_7816,N_7915);
nand U8004 (N_8004,N_7809,N_7844);
nor U8005 (N_8005,N_7876,N_7932);
xnor U8006 (N_8006,N_7808,N_7983);
nor U8007 (N_8007,N_7975,N_7886);
nand U8008 (N_8008,N_7971,N_7981);
or U8009 (N_8009,N_7928,N_7925);
nor U8010 (N_8010,N_7953,N_7859);
xor U8011 (N_8011,N_7814,N_7870);
xor U8012 (N_8012,N_7828,N_7896);
nand U8013 (N_8013,N_7994,N_7831);
and U8014 (N_8014,N_7962,N_7940);
or U8015 (N_8015,N_7840,N_7817);
xnor U8016 (N_8016,N_7911,N_7908);
nand U8017 (N_8017,N_7813,N_7945);
and U8018 (N_8018,N_7972,N_7974);
nor U8019 (N_8019,N_7993,N_7939);
and U8020 (N_8020,N_7871,N_7913);
nor U8021 (N_8021,N_7811,N_7881);
or U8022 (N_8022,N_7875,N_7955);
and U8023 (N_8023,N_7861,N_7883);
xor U8024 (N_8024,N_7984,N_7819);
xnor U8025 (N_8025,N_7853,N_7845);
nand U8026 (N_8026,N_7988,N_7989);
or U8027 (N_8027,N_7986,N_7815);
xnor U8028 (N_8028,N_7897,N_7929);
or U8029 (N_8029,N_7907,N_7880);
xnor U8030 (N_8030,N_7833,N_7982);
or U8031 (N_8031,N_7827,N_7849);
nand U8032 (N_8032,N_7892,N_7977);
xnor U8033 (N_8033,N_7856,N_7807);
or U8034 (N_8034,N_7961,N_7874);
and U8035 (N_8035,N_7930,N_7848);
nand U8036 (N_8036,N_7841,N_7951);
and U8037 (N_8037,N_7866,N_7905);
and U8038 (N_8038,N_7812,N_7898);
nand U8039 (N_8039,N_7947,N_7862);
xnor U8040 (N_8040,N_7917,N_7923);
nor U8041 (N_8041,N_7843,N_7824);
or U8042 (N_8042,N_7837,N_7826);
xor U8043 (N_8043,N_7999,N_7933);
xnor U8044 (N_8044,N_7901,N_7851);
nor U8045 (N_8045,N_7966,N_7852);
or U8046 (N_8046,N_7952,N_7893);
nor U8047 (N_8047,N_7867,N_7835);
nor U8048 (N_8048,N_7864,N_7872);
and U8049 (N_8049,N_7804,N_7887);
or U8050 (N_8050,N_7879,N_7818);
or U8051 (N_8051,N_7855,N_7904);
nand U8052 (N_8052,N_7922,N_7842);
or U8053 (N_8053,N_7964,N_7884);
or U8054 (N_8054,N_7832,N_7878);
nand U8055 (N_8055,N_7937,N_7903);
nand U8056 (N_8056,N_7941,N_7823);
nand U8057 (N_8057,N_7973,N_7863);
nand U8058 (N_8058,N_7810,N_7909);
nand U8059 (N_8059,N_7829,N_7877);
nand U8060 (N_8060,N_7985,N_7885);
or U8061 (N_8061,N_7931,N_7919);
and U8062 (N_8062,N_7894,N_7869);
and U8063 (N_8063,N_7890,N_7918);
and U8064 (N_8064,N_7803,N_7959);
nor U8065 (N_8065,N_7805,N_7960);
xor U8066 (N_8066,N_7938,N_7806);
or U8067 (N_8067,N_7934,N_7873);
or U8068 (N_8068,N_7854,N_7868);
xnor U8069 (N_8069,N_7834,N_7944);
nand U8070 (N_8070,N_7995,N_7821);
nand U8071 (N_8071,N_7860,N_7882);
xnor U8072 (N_8072,N_7891,N_7921);
and U8073 (N_8073,N_7998,N_7979);
xor U8074 (N_8074,N_7943,N_7889);
nand U8075 (N_8075,N_7910,N_7846);
nor U8076 (N_8076,N_7927,N_7895);
and U8077 (N_8077,N_7935,N_7936);
or U8078 (N_8078,N_7958,N_7838);
xor U8079 (N_8079,N_7946,N_7968);
nand U8080 (N_8080,N_7822,N_7847);
nand U8081 (N_8081,N_7899,N_7888);
xor U8082 (N_8082,N_7987,N_7836);
nand U8083 (N_8083,N_7865,N_7965);
nor U8084 (N_8084,N_7956,N_7957);
xor U8085 (N_8085,N_7970,N_7820);
xor U8086 (N_8086,N_7858,N_7906);
nor U8087 (N_8087,N_7942,N_7980);
xor U8088 (N_8088,N_7801,N_7978);
nor U8089 (N_8089,N_7839,N_7914);
nand U8090 (N_8090,N_7949,N_7924);
xnor U8091 (N_8091,N_7916,N_7969);
xor U8092 (N_8092,N_7902,N_7967);
nor U8093 (N_8093,N_7900,N_7920);
and U8094 (N_8094,N_7996,N_7825);
xnor U8095 (N_8095,N_7800,N_7948);
or U8096 (N_8096,N_7926,N_7912);
nand U8097 (N_8097,N_7830,N_7976);
and U8098 (N_8098,N_7950,N_7991);
nand U8099 (N_8099,N_7857,N_7963);
nand U8100 (N_8100,N_7988,N_7991);
or U8101 (N_8101,N_7896,N_7923);
and U8102 (N_8102,N_7925,N_7841);
and U8103 (N_8103,N_7852,N_7973);
and U8104 (N_8104,N_7837,N_7829);
and U8105 (N_8105,N_7978,N_7959);
and U8106 (N_8106,N_7886,N_7890);
or U8107 (N_8107,N_7930,N_7827);
nand U8108 (N_8108,N_7909,N_7825);
nor U8109 (N_8109,N_7896,N_7934);
or U8110 (N_8110,N_7910,N_7941);
xor U8111 (N_8111,N_7904,N_7984);
or U8112 (N_8112,N_7965,N_7916);
and U8113 (N_8113,N_7907,N_7999);
and U8114 (N_8114,N_7843,N_7807);
or U8115 (N_8115,N_7843,N_7808);
nand U8116 (N_8116,N_7954,N_7932);
or U8117 (N_8117,N_7902,N_7913);
xnor U8118 (N_8118,N_7960,N_7954);
nand U8119 (N_8119,N_7971,N_7839);
xor U8120 (N_8120,N_7818,N_7803);
xnor U8121 (N_8121,N_7930,N_7889);
and U8122 (N_8122,N_7819,N_7970);
xor U8123 (N_8123,N_7926,N_7933);
nor U8124 (N_8124,N_7841,N_7966);
nor U8125 (N_8125,N_7908,N_7810);
xor U8126 (N_8126,N_7941,N_7989);
nand U8127 (N_8127,N_7891,N_7893);
nand U8128 (N_8128,N_7880,N_7925);
or U8129 (N_8129,N_7924,N_7811);
nand U8130 (N_8130,N_7922,N_7938);
xor U8131 (N_8131,N_7953,N_7871);
nand U8132 (N_8132,N_7987,N_7835);
nor U8133 (N_8133,N_7883,N_7840);
nor U8134 (N_8134,N_7946,N_7880);
or U8135 (N_8135,N_7967,N_7850);
nand U8136 (N_8136,N_7960,N_7909);
nor U8137 (N_8137,N_7933,N_7961);
nand U8138 (N_8138,N_7923,N_7958);
and U8139 (N_8139,N_7836,N_7827);
or U8140 (N_8140,N_7902,N_7877);
nor U8141 (N_8141,N_7882,N_7843);
or U8142 (N_8142,N_7925,N_7942);
nand U8143 (N_8143,N_7938,N_7828);
or U8144 (N_8144,N_7932,N_7914);
and U8145 (N_8145,N_7825,N_7990);
nand U8146 (N_8146,N_7899,N_7991);
xnor U8147 (N_8147,N_7868,N_7872);
or U8148 (N_8148,N_7818,N_7808);
or U8149 (N_8149,N_7917,N_7815);
and U8150 (N_8150,N_7936,N_7801);
xnor U8151 (N_8151,N_7959,N_7836);
xnor U8152 (N_8152,N_7841,N_7888);
xnor U8153 (N_8153,N_7841,N_7858);
nor U8154 (N_8154,N_7874,N_7800);
and U8155 (N_8155,N_7818,N_7885);
nor U8156 (N_8156,N_7802,N_7998);
nor U8157 (N_8157,N_7997,N_7807);
and U8158 (N_8158,N_7909,N_7986);
nor U8159 (N_8159,N_7858,N_7860);
nor U8160 (N_8160,N_7961,N_7965);
and U8161 (N_8161,N_7968,N_7917);
nor U8162 (N_8162,N_7877,N_7957);
nand U8163 (N_8163,N_7905,N_7970);
nand U8164 (N_8164,N_7967,N_7910);
nor U8165 (N_8165,N_7897,N_7923);
nand U8166 (N_8166,N_7904,N_7926);
xor U8167 (N_8167,N_7945,N_7849);
nand U8168 (N_8168,N_7896,N_7912);
nand U8169 (N_8169,N_7869,N_7855);
xnor U8170 (N_8170,N_7815,N_7920);
and U8171 (N_8171,N_7931,N_7985);
nor U8172 (N_8172,N_7883,N_7897);
xnor U8173 (N_8173,N_7862,N_7828);
xnor U8174 (N_8174,N_7968,N_7990);
and U8175 (N_8175,N_7929,N_7973);
nand U8176 (N_8176,N_7843,N_7850);
and U8177 (N_8177,N_7831,N_7927);
and U8178 (N_8178,N_7942,N_7970);
xnor U8179 (N_8179,N_7815,N_7816);
and U8180 (N_8180,N_7979,N_7852);
xnor U8181 (N_8181,N_7878,N_7933);
xor U8182 (N_8182,N_7868,N_7865);
or U8183 (N_8183,N_7942,N_7866);
nand U8184 (N_8184,N_7920,N_7862);
nand U8185 (N_8185,N_7996,N_7905);
and U8186 (N_8186,N_7986,N_7958);
nand U8187 (N_8187,N_7809,N_7881);
or U8188 (N_8188,N_7913,N_7882);
nor U8189 (N_8189,N_7825,N_7821);
and U8190 (N_8190,N_7949,N_7852);
and U8191 (N_8191,N_7927,N_7840);
xnor U8192 (N_8192,N_7885,N_7869);
or U8193 (N_8193,N_7858,N_7859);
nand U8194 (N_8194,N_7937,N_7827);
xor U8195 (N_8195,N_7933,N_7927);
and U8196 (N_8196,N_7982,N_7911);
and U8197 (N_8197,N_7854,N_7952);
xnor U8198 (N_8198,N_7848,N_7900);
nor U8199 (N_8199,N_7889,N_7894);
nor U8200 (N_8200,N_8016,N_8192);
or U8201 (N_8201,N_8101,N_8126);
or U8202 (N_8202,N_8061,N_8131);
xor U8203 (N_8203,N_8007,N_8173);
nand U8204 (N_8204,N_8193,N_8092);
and U8205 (N_8205,N_8179,N_8098);
and U8206 (N_8206,N_8075,N_8198);
or U8207 (N_8207,N_8142,N_8033);
xnor U8208 (N_8208,N_8153,N_8029);
xor U8209 (N_8209,N_8130,N_8162);
nand U8210 (N_8210,N_8189,N_8084);
and U8211 (N_8211,N_8129,N_8058);
nor U8212 (N_8212,N_8125,N_8168);
and U8213 (N_8213,N_8062,N_8004);
nand U8214 (N_8214,N_8134,N_8091);
nor U8215 (N_8215,N_8115,N_8077);
and U8216 (N_8216,N_8104,N_8139);
nor U8217 (N_8217,N_8022,N_8049);
or U8218 (N_8218,N_8155,N_8013);
and U8219 (N_8219,N_8119,N_8071);
nand U8220 (N_8220,N_8078,N_8197);
nor U8221 (N_8221,N_8086,N_8100);
and U8222 (N_8222,N_8145,N_8018);
and U8223 (N_8223,N_8147,N_8178);
or U8224 (N_8224,N_8060,N_8037);
nand U8225 (N_8225,N_8132,N_8122);
or U8226 (N_8226,N_8118,N_8081);
or U8227 (N_8227,N_8056,N_8158);
or U8228 (N_8228,N_8065,N_8008);
nand U8229 (N_8229,N_8025,N_8074);
or U8230 (N_8230,N_8123,N_8076);
or U8231 (N_8231,N_8034,N_8050);
nor U8232 (N_8232,N_8047,N_8048);
nor U8233 (N_8233,N_8040,N_8113);
nand U8234 (N_8234,N_8127,N_8088);
xor U8235 (N_8235,N_8166,N_8044);
or U8236 (N_8236,N_8090,N_8176);
nand U8237 (N_8237,N_8096,N_8128);
or U8238 (N_8238,N_8045,N_8114);
nor U8239 (N_8239,N_8159,N_8021);
xor U8240 (N_8240,N_8046,N_8140);
xnor U8241 (N_8241,N_8195,N_8059);
nor U8242 (N_8242,N_8121,N_8180);
or U8243 (N_8243,N_8106,N_8185);
and U8244 (N_8244,N_8188,N_8035);
or U8245 (N_8245,N_8111,N_8093);
xnor U8246 (N_8246,N_8082,N_8141);
nand U8247 (N_8247,N_8102,N_8136);
or U8248 (N_8248,N_8068,N_8097);
xor U8249 (N_8249,N_8023,N_8135);
or U8250 (N_8250,N_8160,N_8175);
xnor U8251 (N_8251,N_8154,N_8053);
and U8252 (N_8252,N_8066,N_8199);
and U8253 (N_8253,N_8027,N_8003);
or U8254 (N_8254,N_8112,N_8042);
nor U8255 (N_8255,N_8187,N_8030);
nand U8256 (N_8256,N_8087,N_8038);
or U8257 (N_8257,N_8182,N_8172);
nor U8258 (N_8258,N_8064,N_8005);
or U8259 (N_8259,N_8149,N_8107);
nor U8260 (N_8260,N_8117,N_8000);
and U8261 (N_8261,N_8020,N_8026);
nand U8262 (N_8262,N_8039,N_8085);
xnor U8263 (N_8263,N_8052,N_8024);
nand U8264 (N_8264,N_8014,N_8001);
xor U8265 (N_8265,N_8073,N_8051);
xnor U8266 (N_8266,N_8006,N_8012);
or U8267 (N_8267,N_8138,N_8186);
and U8268 (N_8268,N_8184,N_8057);
nand U8269 (N_8269,N_8144,N_8011);
or U8270 (N_8270,N_8009,N_8110);
or U8271 (N_8271,N_8070,N_8157);
xor U8272 (N_8272,N_8191,N_8167);
nand U8273 (N_8273,N_8165,N_8063);
and U8274 (N_8274,N_8094,N_8010);
xnor U8275 (N_8275,N_8067,N_8171);
and U8276 (N_8276,N_8072,N_8054);
and U8277 (N_8277,N_8124,N_8163);
or U8278 (N_8278,N_8089,N_8151);
nand U8279 (N_8279,N_8109,N_8143);
nand U8280 (N_8280,N_8181,N_8108);
xor U8281 (N_8281,N_8148,N_8169);
xnor U8282 (N_8282,N_8161,N_8017);
xnor U8283 (N_8283,N_8105,N_8170);
and U8284 (N_8284,N_8164,N_8043);
nand U8285 (N_8285,N_8196,N_8041);
or U8286 (N_8286,N_8146,N_8036);
nand U8287 (N_8287,N_8116,N_8183);
nand U8288 (N_8288,N_8069,N_8137);
or U8289 (N_8289,N_8032,N_8152);
nand U8290 (N_8290,N_8095,N_8031);
xor U8291 (N_8291,N_8177,N_8002);
xor U8292 (N_8292,N_8015,N_8133);
xor U8293 (N_8293,N_8083,N_8055);
and U8294 (N_8294,N_8194,N_8120);
nand U8295 (N_8295,N_8174,N_8080);
nor U8296 (N_8296,N_8019,N_8156);
and U8297 (N_8297,N_8190,N_8103);
nor U8298 (N_8298,N_8079,N_8099);
and U8299 (N_8299,N_8028,N_8150);
or U8300 (N_8300,N_8044,N_8199);
xor U8301 (N_8301,N_8006,N_8192);
nand U8302 (N_8302,N_8005,N_8159);
or U8303 (N_8303,N_8048,N_8101);
or U8304 (N_8304,N_8016,N_8195);
or U8305 (N_8305,N_8184,N_8079);
nand U8306 (N_8306,N_8091,N_8063);
nor U8307 (N_8307,N_8175,N_8052);
nor U8308 (N_8308,N_8168,N_8185);
nor U8309 (N_8309,N_8121,N_8094);
xnor U8310 (N_8310,N_8157,N_8133);
or U8311 (N_8311,N_8038,N_8099);
nand U8312 (N_8312,N_8017,N_8086);
nor U8313 (N_8313,N_8072,N_8082);
nand U8314 (N_8314,N_8137,N_8116);
and U8315 (N_8315,N_8045,N_8137);
nor U8316 (N_8316,N_8123,N_8165);
and U8317 (N_8317,N_8174,N_8079);
nand U8318 (N_8318,N_8169,N_8189);
nand U8319 (N_8319,N_8080,N_8043);
or U8320 (N_8320,N_8166,N_8189);
nand U8321 (N_8321,N_8084,N_8155);
nand U8322 (N_8322,N_8122,N_8003);
nand U8323 (N_8323,N_8043,N_8069);
nand U8324 (N_8324,N_8160,N_8021);
nor U8325 (N_8325,N_8074,N_8020);
nand U8326 (N_8326,N_8163,N_8031);
nor U8327 (N_8327,N_8197,N_8035);
xnor U8328 (N_8328,N_8042,N_8001);
and U8329 (N_8329,N_8164,N_8143);
and U8330 (N_8330,N_8164,N_8167);
xor U8331 (N_8331,N_8042,N_8123);
and U8332 (N_8332,N_8179,N_8053);
xor U8333 (N_8333,N_8115,N_8192);
or U8334 (N_8334,N_8099,N_8117);
nor U8335 (N_8335,N_8043,N_8046);
xnor U8336 (N_8336,N_8082,N_8035);
xor U8337 (N_8337,N_8116,N_8141);
and U8338 (N_8338,N_8073,N_8180);
nand U8339 (N_8339,N_8171,N_8139);
nor U8340 (N_8340,N_8154,N_8173);
nand U8341 (N_8341,N_8142,N_8040);
or U8342 (N_8342,N_8015,N_8141);
or U8343 (N_8343,N_8036,N_8103);
or U8344 (N_8344,N_8133,N_8079);
xnor U8345 (N_8345,N_8049,N_8074);
nand U8346 (N_8346,N_8103,N_8030);
or U8347 (N_8347,N_8087,N_8024);
xnor U8348 (N_8348,N_8048,N_8152);
and U8349 (N_8349,N_8046,N_8117);
or U8350 (N_8350,N_8079,N_8136);
nand U8351 (N_8351,N_8048,N_8023);
or U8352 (N_8352,N_8189,N_8018);
and U8353 (N_8353,N_8031,N_8171);
xnor U8354 (N_8354,N_8128,N_8067);
xnor U8355 (N_8355,N_8105,N_8180);
and U8356 (N_8356,N_8045,N_8169);
or U8357 (N_8357,N_8087,N_8054);
nor U8358 (N_8358,N_8014,N_8144);
or U8359 (N_8359,N_8026,N_8050);
xor U8360 (N_8360,N_8027,N_8080);
xnor U8361 (N_8361,N_8063,N_8052);
nor U8362 (N_8362,N_8085,N_8126);
and U8363 (N_8363,N_8063,N_8193);
nor U8364 (N_8364,N_8124,N_8044);
and U8365 (N_8365,N_8083,N_8063);
and U8366 (N_8366,N_8151,N_8157);
or U8367 (N_8367,N_8173,N_8143);
xor U8368 (N_8368,N_8146,N_8119);
nor U8369 (N_8369,N_8047,N_8146);
xor U8370 (N_8370,N_8021,N_8146);
xor U8371 (N_8371,N_8178,N_8006);
nand U8372 (N_8372,N_8195,N_8116);
nor U8373 (N_8373,N_8016,N_8069);
or U8374 (N_8374,N_8035,N_8101);
or U8375 (N_8375,N_8047,N_8088);
or U8376 (N_8376,N_8026,N_8027);
nand U8377 (N_8377,N_8022,N_8149);
nor U8378 (N_8378,N_8088,N_8176);
or U8379 (N_8379,N_8025,N_8079);
xor U8380 (N_8380,N_8158,N_8051);
nor U8381 (N_8381,N_8058,N_8154);
and U8382 (N_8382,N_8026,N_8192);
nand U8383 (N_8383,N_8028,N_8152);
xor U8384 (N_8384,N_8094,N_8056);
nor U8385 (N_8385,N_8004,N_8126);
nand U8386 (N_8386,N_8075,N_8004);
nand U8387 (N_8387,N_8139,N_8184);
and U8388 (N_8388,N_8171,N_8020);
nand U8389 (N_8389,N_8140,N_8157);
and U8390 (N_8390,N_8025,N_8174);
or U8391 (N_8391,N_8169,N_8178);
nand U8392 (N_8392,N_8193,N_8081);
xor U8393 (N_8393,N_8167,N_8128);
xor U8394 (N_8394,N_8146,N_8059);
xnor U8395 (N_8395,N_8017,N_8140);
or U8396 (N_8396,N_8085,N_8199);
xnor U8397 (N_8397,N_8009,N_8139);
nand U8398 (N_8398,N_8161,N_8103);
xnor U8399 (N_8399,N_8084,N_8156);
nand U8400 (N_8400,N_8216,N_8290);
or U8401 (N_8401,N_8388,N_8285);
and U8402 (N_8402,N_8293,N_8226);
or U8403 (N_8403,N_8259,N_8297);
or U8404 (N_8404,N_8304,N_8294);
or U8405 (N_8405,N_8397,N_8282);
or U8406 (N_8406,N_8344,N_8278);
xnor U8407 (N_8407,N_8224,N_8366);
and U8408 (N_8408,N_8398,N_8387);
xnor U8409 (N_8409,N_8205,N_8233);
or U8410 (N_8410,N_8238,N_8279);
nor U8411 (N_8411,N_8303,N_8325);
xor U8412 (N_8412,N_8383,N_8322);
xnor U8413 (N_8413,N_8234,N_8220);
and U8414 (N_8414,N_8335,N_8330);
or U8415 (N_8415,N_8360,N_8345);
or U8416 (N_8416,N_8207,N_8248);
nand U8417 (N_8417,N_8200,N_8256);
xor U8418 (N_8418,N_8312,N_8318);
xor U8419 (N_8419,N_8370,N_8362);
xnor U8420 (N_8420,N_8310,N_8311);
nor U8421 (N_8421,N_8242,N_8378);
xor U8422 (N_8422,N_8382,N_8340);
nand U8423 (N_8423,N_8308,N_8301);
nand U8424 (N_8424,N_8280,N_8392);
or U8425 (N_8425,N_8288,N_8327);
nand U8426 (N_8426,N_8355,N_8385);
xor U8427 (N_8427,N_8295,N_8246);
xor U8428 (N_8428,N_8269,N_8346);
nor U8429 (N_8429,N_8323,N_8331);
nor U8430 (N_8430,N_8391,N_8271);
or U8431 (N_8431,N_8237,N_8364);
nand U8432 (N_8432,N_8263,N_8296);
or U8433 (N_8433,N_8365,N_8374);
xor U8434 (N_8434,N_8321,N_8396);
and U8435 (N_8435,N_8343,N_8229);
or U8436 (N_8436,N_8265,N_8257);
or U8437 (N_8437,N_8316,N_8268);
or U8438 (N_8438,N_8291,N_8299);
or U8439 (N_8439,N_8266,N_8314);
or U8440 (N_8440,N_8337,N_8375);
or U8441 (N_8441,N_8206,N_8390);
nand U8442 (N_8442,N_8223,N_8239);
nand U8443 (N_8443,N_8394,N_8326);
xnor U8444 (N_8444,N_8332,N_8358);
xnor U8445 (N_8445,N_8247,N_8250);
nor U8446 (N_8446,N_8222,N_8252);
and U8447 (N_8447,N_8272,N_8381);
xor U8448 (N_8448,N_8244,N_8212);
nor U8449 (N_8449,N_8399,N_8315);
nand U8450 (N_8450,N_8211,N_8363);
nand U8451 (N_8451,N_8320,N_8249);
nand U8452 (N_8452,N_8210,N_8262);
or U8453 (N_8453,N_8348,N_8228);
xnor U8454 (N_8454,N_8350,N_8329);
and U8455 (N_8455,N_8328,N_8349);
or U8456 (N_8456,N_8384,N_8264);
and U8457 (N_8457,N_8219,N_8339);
and U8458 (N_8458,N_8359,N_8251);
nand U8459 (N_8459,N_8277,N_8276);
nand U8460 (N_8460,N_8319,N_8231);
or U8461 (N_8461,N_8351,N_8204);
nand U8462 (N_8462,N_8334,N_8214);
xnor U8463 (N_8463,N_8217,N_8209);
or U8464 (N_8464,N_8313,N_8267);
xnor U8465 (N_8465,N_8286,N_8243);
nor U8466 (N_8466,N_8241,N_8386);
nand U8467 (N_8467,N_8347,N_8361);
nor U8468 (N_8468,N_8369,N_8305);
and U8469 (N_8469,N_8302,N_8274);
xnor U8470 (N_8470,N_8281,N_8232);
nor U8471 (N_8471,N_8289,N_8373);
or U8472 (N_8472,N_8356,N_8379);
nand U8473 (N_8473,N_8357,N_8253);
nand U8474 (N_8474,N_8225,N_8218);
and U8475 (N_8475,N_8300,N_8372);
or U8476 (N_8476,N_8201,N_8393);
nor U8477 (N_8477,N_8306,N_8338);
xor U8478 (N_8478,N_8284,N_8307);
and U8479 (N_8479,N_8227,N_8236);
and U8480 (N_8480,N_8367,N_8317);
and U8481 (N_8481,N_8202,N_8377);
nand U8482 (N_8482,N_8258,N_8287);
nand U8483 (N_8483,N_8342,N_8324);
nor U8484 (N_8484,N_8235,N_8352);
or U8485 (N_8485,N_8341,N_8245);
or U8486 (N_8486,N_8333,N_8292);
xnor U8487 (N_8487,N_8203,N_8255);
nor U8488 (N_8488,N_8213,N_8215);
xnor U8489 (N_8489,N_8371,N_8260);
nor U8490 (N_8490,N_8254,N_8273);
nor U8491 (N_8491,N_8380,N_8368);
nor U8492 (N_8492,N_8240,N_8336);
xor U8493 (N_8493,N_8353,N_8389);
nor U8494 (N_8494,N_8298,N_8395);
xor U8495 (N_8495,N_8376,N_8309);
and U8496 (N_8496,N_8270,N_8208);
nor U8497 (N_8497,N_8261,N_8275);
xor U8498 (N_8498,N_8283,N_8221);
nand U8499 (N_8499,N_8230,N_8354);
or U8500 (N_8500,N_8303,N_8201);
xnor U8501 (N_8501,N_8232,N_8325);
and U8502 (N_8502,N_8345,N_8234);
nand U8503 (N_8503,N_8381,N_8383);
nand U8504 (N_8504,N_8356,N_8277);
xnor U8505 (N_8505,N_8214,N_8333);
nand U8506 (N_8506,N_8289,N_8272);
nor U8507 (N_8507,N_8297,N_8350);
and U8508 (N_8508,N_8251,N_8205);
nor U8509 (N_8509,N_8340,N_8397);
and U8510 (N_8510,N_8217,N_8240);
or U8511 (N_8511,N_8213,N_8276);
and U8512 (N_8512,N_8322,N_8386);
xnor U8513 (N_8513,N_8213,N_8310);
xnor U8514 (N_8514,N_8263,N_8246);
and U8515 (N_8515,N_8205,N_8297);
xor U8516 (N_8516,N_8356,N_8208);
or U8517 (N_8517,N_8346,N_8287);
nand U8518 (N_8518,N_8275,N_8296);
nand U8519 (N_8519,N_8366,N_8277);
nand U8520 (N_8520,N_8339,N_8384);
xor U8521 (N_8521,N_8363,N_8220);
xor U8522 (N_8522,N_8399,N_8387);
xnor U8523 (N_8523,N_8251,N_8357);
and U8524 (N_8524,N_8270,N_8350);
nand U8525 (N_8525,N_8311,N_8355);
xor U8526 (N_8526,N_8222,N_8257);
nand U8527 (N_8527,N_8200,N_8305);
or U8528 (N_8528,N_8252,N_8201);
nand U8529 (N_8529,N_8261,N_8312);
and U8530 (N_8530,N_8222,N_8391);
nand U8531 (N_8531,N_8383,N_8331);
nor U8532 (N_8532,N_8275,N_8203);
nand U8533 (N_8533,N_8290,N_8328);
nand U8534 (N_8534,N_8337,N_8345);
or U8535 (N_8535,N_8277,N_8319);
nand U8536 (N_8536,N_8382,N_8374);
or U8537 (N_8537,N_8241,N_8295);
xnor U8538 (N_8538,N_8233,N_8249);
xor U8539 (N_8539,N_8339,N_8247);
xnor U8540 (N_8540,N_8322,N_8262);
nand U8541 (N_8541,N_8365,N_8202);
nand U8542 (N_8542,N_8252,N_8366);
nand U8543 (N_8543,N_8261,N_8304);
xnor U8544 (N_8544,N_8361,N_8206);
and U8545 (N_8545,N_8341,N_8282);
and U8546 (N_8546,N_8399,N_8366);
xor U8547 (N_8547,N_8338,N_8260);
nand U8548 (N_8548,N_8347,N_8218);
and U8549 (N_8549,N_8202,N_8229);
and U8550 (N_8550,N_8235,N_8201);
and U8551 (N_8551,N_8330,N_8354);
and U8552 (N_8552,N_8318,N_8275);
nor U8553 (N_8553,N_8356,N_8219);
xnor U8554 (N_8554,N_8367,N_8370);
xor U8555 (N_8555,N_8346,N_8211);
nor U8556 (N_8556,N_8261,N_8253);
xor U8557 (N_8557,N_8313,N_8316);
and U8558 (N_8558,N_8361,N_8358);
and U8559 (N_8559,N_8330,N_8303);
and U8560 (N_8560,N_8297,N_8286);
nor U8561 (N_8561,N_8256,N_8355);
and U8562 (N_8562,N_8310,N_8238);
nor U8563 (N_8563,N_8233,N_8262);
nor U8564 (N_8564,N_8237,N_8213);
nand U8565 (N_8565,N_8276,N_8383);
and U8566 (N_8566,N_8363,N_8237);
nand U8567 (N_8567,N_8284,N_8238);
and U8568 (N_8568,N_8249,N_8212);
xnor U8569 (N_8569,N_8210,N_8304);
xor U8570 (N_8570,N_8329,N_8359);
nand U8571 (N_8571,N_8375,N_8355);
nand U8572 (N_8572,N_8271,N_8202);
xor U8573 (N_8573,N_8304,N_8333);
or U8574 (N_8574,N_8256,N_8244);
nand U8575 (N_8575,N_8286,N_8288);
xnor U8576 (N_8576,N_8369,N_8217);
xor U8577 (N_8577,N_8295,N_8305);
and U8578 (N_8578,N_8309,N_8279);
xor U8579 (N_8579,N_8367,N_8298);
xnor U8580 (N_8580,N_8285,N_8312);
or U8581 (N_8581,N_8317,N_8339);
nor U8582 (N_8582,N_8316,N_8310);
nor U8583 (N_8583,N_8270,N_8305);
and U8584 (N_8584,N_8342,N_8360);
and U8585 (N_8585,N_8212,N_8319);
and U8586 (N_8586,N_8263,N_8216);
and U8587 (N_8587,N_8380,N_8396);
xnor U8588 (N_8588,N_8355,N_8318);
nand U8589 (N_8589,N_8273,N_8256);
nor U8590 (N_8590,N_8285,N_8303);
nand U8591 (N_8591,N_8242,N_8308);
or U8592 (N_8592,N_8232,N_8299);
or U8593 (N_8593,N_8342,N_8200);
xor U8594 (N_8594,N_8245,N_8322);
xor U8595 (N_8595,N_8284,N_8363);
nor U8596 (N_8596,N_8234,N_8368);
or U8597 (N_8597,N_8336,N_8332);
nor U8598 (N_8598,N_8244,N_8201);
nand U8599 (N_8599,N_8334,N_8206);
and U8600 (N_8600,N_8414,N_8454);
nor U8601 (N_8601,N_8550,N_8530);
nor U8602 (N_8602,N_8419,N_8497);
xor U8603 (N_8603,N_8468,N_8491);
or U8604 (N_8604,N_8511,N_8416);
nand U8605 (N_8605,N_8555,N_8580);
or U8606 (N_8606,N_8574,N_8589);
xnor U8607 (N_8607,N_8409,N_8552);
and U8608 (N_8608,N_8439,N_8400);
nor U8609 (N_8609,N_8449,N_8532);
nand U8610 (N_8610,N_8518,N_8429);
nor U8611 (N_8611,N_8551,N_8411);
nor U8612 (N_8612,N_8458,N_8421);
nor U8613 (N_8613,N_8540,N_8443);
nor U8614 (N_8614,N_8598,N_8542);
nor U8615 (N_8615,N_8565,N_8592);
or U8616 (N_8616,N_8405,N_8436);
or U8617 (N_8617,N_8466,N_8403);
xor U8618 (N_8618,N_8402,N_8517);
nand U8619 (N_8619,N_8410,N_8432);
or U8620 (N_8620,N_8445,N_8545);
and U8621 (N_8621,N_8450,N_8437);
nand U8622 (N_8622,N_8461,N_8418);
nor U8623 (N_8623,N_8577,N_8506);
xnor U8624 (N_8624,N_8544,N_8539);
xor U8625 (N_8625,N_8498,N_8459);
nand U8626 (N_8626,N_8549,N_8590);
nand U8627 (N_8627,N_8487,N_8425);
and U8628 (N_8628,N_8509,N_8528);
nand U8629 (N_8629,N_8512,N_8452);
and U8630 (N_8630,N_8541,N_8486);
nor U8631 (N_8631,N_8470,N_8538);
nor U8632 (N_8632,N_8407,N_8440);
and U8633 (N_8633,N_8571,N_8529);
or U8634 (N_8634,N_8561,N_8430);
nor U8635 (N_8635,N_8569,N_8547);
and U8636 (N_8636,N_8485,N_8501);
or U8637 (N_8637,N_8490,N_8438);
or U8638 (N_8638,N_8558,N_8424);
nor U8639 (N_8639,N_8570,N_8441);
nor U8640 (N_8640,N_8502,N_8460);
and U8641 (N_8641,N_8464,N_8453);
or U8642 (N_8642,N_8427,N_8448);
or U8643 (N_8643,N_8428,N_8478);
nand U8644 (N_8644,N_8423,N_8499);
nand U8645 (N_8645,N_8557,N_8493);
nand U8646 (N_8646,N_8472,N_8479);
and U8647 (N_8647,N_8465,N_8447);
nor U8648 (N_8648,N_8568,N_8508);
nand U8649 (N_8649,N_8554,N_8520);
xor U8650 (N_8650,N_8431,N_8401);
nand U8651 (N_8651,N_8417,N_8583);
or U8652 (N_8652,N_8484,N_8467);
nand U8653 (N_8653,N_8455,N_8489);
nand U8654 (N_8654,N_8599,N_8471);
xor U8655 (N_8655,N_8474,N_8516);
nor U8656 (N_8656,N_8514,N_8560);
or U8657 (N_8657,N_8567,N_8513);
nand U8658 (N_8658,N_8531,N_8579);
nand U8659 (N_8659,N_8559,N_8475);
and U8660 (N_8660,N_8537,N_8462);
nand U8661 (N_8661,N_8413,N_8488);
nand U8662 (N_8662,N_8563,N_8593);
nor U8663 (N_8663,N_8519,N_8482);
xor U8664 (N_8664,N_8523,N_8535);
nand U8665 (N_8665,N_8585,N_8426);
or U8666 (N_8666,N_8435,N_8446);
or U8667 (N_8667,N_8481,N_8507);
and U8668 (N_8668,N_8534,N_8548);
xnor U8669 (N_8669,N_8463,N_8573);
and U8670 (N_8670,N_8503,N_8433);
or U8671 (N_8671,N_8553,N_8596);
nor U8672 (N_8672,N_8584,N_8406);
and U8673 (N_8673,N_8556,N_8522);
xor U8674 (N_8674,N_8576,N_8526);
or U8675 (N_8675,N_8527,N_8456);
nor U8676 (N_8676,N_8543,N_8510);
and U8677 (N_8677,N_8496,N_8494);
xor U8678 (N_8678,N_8578,N_8586);
nand U8679 (N_8679,N_8524,N_8536);
nor U8680 (N_8680,N_8587,N_8595);
nand U8681 (N_8681,N_8404,N_8451);
or U8682 (N_8682,N_8469,N_8515);
and U8683 (N_8683,N_8500,N_8476);
and U8684 (N_8684,N_8477,N_8566);
nand U8685 (N_8685,N_8572,N_8582);
and U8686 (N_8686,N_8575,N_8505);
or U8687 (N_8687,N_8495,N_8564);
or U8688 (N_8688,N_8422,N_8412);
and U8689 (N_8689,N_8480,N_8562);
nor U8690 (N_8690,N_8591,N_8444);
nand U8691 (N_8691,N_8415,N_8442);
xor U8692 (N_8692,N_8594,N_8588);
nand U8693 (N_8693,N_8408,N_8492);
or U8694 (N_8694,N_8483,N_8546);
xnor U8695 (N_8695,N_8434,N_8457);
and U8696 (N_8696,N_8521,N_8473);
nor U8697 (N_8697,N_8420,N_8525);
nor U8698 (N_8698,N_8581,N_8597);
nand U8699 (N_8699,N_8504,N_8533);
or U8700 (N_8700,N_8559,N_8505);
nand U8701 (N_8701,N_8588,N_8461);
or U8702 (N_8702,N_8583,N_8530);
or U8703 (N_8703,N_8494,N_8513);
nand U8704 (N_8704,N_8411,N_8500);
or U8705 (N_8705,N_8578,N_8420);
nand U8706 (N_8706,N_8402,N_8443);
nand U8707 (N_8707,N_8517,N_8418);
xnor U8708 (N_8708,N_8546,N_8435);
nand U8709 (N_8709,N_8510,N_8495);
and U8710 (N_8710,N_8443,N_8442);
nand U8711 (N_8711,N_8543,N_8409);
xnor U8712 (N_8712,N_8420,N_8505);
nor U8713 (N_8713,N_8561,N_8596);
or U8714 (N_8714,N_8482,N_8412);
nand U8715 (N_8715,N_8512,N_8455);
and U8716 (N_8716,N_8519,N_8489);
and U8717 (N_8717,N_8521,N_8447);
nand U8718 (N_8718,N_8508,N_8548);
xnor U8719 (N_8719,N_8591,N_8456);
nor U8720 (N_8720,N_8581,N_8491);
xor U8721 (N_8721,N_8575,N_8538);
and U8722 (N_8722,N_8441,N_8461);
nor U8723 (N_8723,N_8506,N_8515);
and U8724 (N_8724,N_8570,N_8596);
nand U8725 (N_8725,N_8537,N_8453);
xnor U8726 (N_8726,N_8599,N_8464);
nand U8727 (N_8727,N_8547,N_8499);
nor U8728 (N_8728,N_8581,N_8579);
xor U8729 (N_8729,N_8569,N_8507);
and U8730 (N_8730,N_8462,N_8531);
nor U8731 (N_8731,N_8429,N_8507);
xnor U8732 (N_8732,N_8423,N_8592);
and U8733 (N_8733,N_8559,N_8560);
nand U8734 (N_8734,N_8525,N_8563);
and U8735 (N_8735,N_8444,N_8563);
nand U8736 (N_8736,N_8506,N_8592);
or U8737 (N_8737,N_8585,N_8458);
nor U8738 (N_8738,N_8456,N_8453);
and U8739 (N_8739,N_8559,N_8541);
nor U8740 (N_8740,N_8565,N_8532);
xnor U8741 (N_8741,N_8540,N_8449);
xor U8742 (N_8742,N_8418,N_8552);
and U8743 (N_8743,N_8457,N_8579);
and U8744 (N_8744,N_8424,N_8413);
or U8745 (N_8745,N_8590,N_8427);
nand U8746 (N_8746,N_8476,N_8417);
nor U8747 (N_8747,N_8448,N_8413);
nor U8748 (N_8748,N_8502,N_8564);
nor U8749 (N_8749,N_8436,N_8438);
or U8750 (N_8750,N_8438,N_8584);
xnor U8751 (N_8751,N_8540,N_8455);
and U8752 (N_8752,N_8413,N_8548);
nand U8753 (N_8753,N_8563,N_8518);
nor U8754 (N_8754,N_8536,N_8452);
or U8755 (N_8755,N_8556,N_8407);
xor U8756 (N_8756,N_8566,N_8491);
or U8757 (N_8757,N_8535,N_8462);
xor U8758 (N_8758,N_8531,N_8537);
and U8759 (N_8759,N_8532,N_8552);
and U8760 (N_8760,N_8585,N_8439);
and U8761 (N_8761,N_8409,N_8519);
or U8762 (N_8762,N_8408,N_8579);
nand U8763 (N_8763,N_8449,N_8466);
nand U8764 (N_8764,N_8537,N_8493);
nand U8765 (N_8765,N_8443,N_8573);
or U8766 (N_8766,N_8401,N_8560);
or U8767 (N_8767,N_8534,N_8494);
nand U8768 (N_8768,N_8557,N_8492);
nor U8769 (N_8769,N_8494,N_8464);
xnor U8770 (N_8770,N_8563,N_8496);
and U8771 (N_8771,N_8515,N_8594);
and U8772 (N_8772,N_8442,N_8451);
nor U8773 (N_8773,N_8440,N_8586);
and U8774 (N_8774,N_8409,N_8491);
xnor U8775 (N_8775,N_8550,N_8457);
xor U8776 (N_8776,N_8589,N_8593);
nand U8777 (N_8777,N_8580,N_8564);
xnor U8778 (N_8778,N_8584,N_8595);
or U8779 (N_8779,N_8409,N_8584);
and U8780 (N_8780,N_8478,N_8546);
and U8781 (N_8781,N_8431,N_8543);
nand U8782 (N_8782,N_8513,N_8440);
or U8783 (N_8783,N_8497,N_8491);
or U8784 (N_8784,N_8584,N_8515);
or U8785 (N_8785,N_8489,N_8569);
or U8786 (N_8786,N_8575,N_8416);
xor U8787 (N_8787,N_8564,N_8560);
xor U8788 (N_8788,N_8494,N_8549);
or U8789 (N_8789,N_8495,N_8400);
nor U8790 (N_8790,N_8551,N_8520);
nor U8791 (N_8791,N_8413,N_8592);
and U8792 (N_8792,N_8493,N_8447);
nor U8793 (N_8793,N_8509,N_8497);
and U8794 (N_8794,N_8596,N_8575);
or U8795 (N_8795,N_8546,N_8547);
nand U8796 (N_8796,N_8452,N_8427);
and U8797 (N_8797,N_8522,N_8582);
and U8798 (N_8798,N_8402,N_8448);
nor U8799 (N_8799,N_8494,N_8480);
nand U8800 (N_8800,N_8668,N_8712);
xnor U8801 (N_8801,N_8707,N_8735);
nand U8802 (N_8802,N_8738,N_8676);
and U8803 (N_8803,N_8752,N_8736);
or U8804 (N_8804,N_8695,N_8797);
or U8805 (N_8805,N_8799,N_8772);
and U8806 (N_8806,N_8673,N_8764);
and U8807 (N_8807,N_8766,N_8775);
xor U8808 (N_8808,N_8776,N_8606);
or U8809 (N_8809,N_8777,N_8779);
and U8810 (N_8810,N_8617,N_8696);
and U8811 (N_8811,N_8742,N_8615);
nand U8812 (N_8812,N_8630,N_8732);
and U8813 (N_8813,N_8678,N_8651);
and U8814 (N_8814,N_8748,N_8619);
or U8815 (N_8815,N_8734,N_8773);
nor U8816 (N_8816,N_8758,N_8768);
or U8817 (N_8817,N_8697,N_8703);
and U8818 (N_8818,N_8716,N_8719);
xnor U8819 (N_8819,N_8746,N_8622);
and U8820 (N_8820,N_8770,N_8715);
nor U8821 (N_8821,N_8756,N_8739);
nor U8822 (N_8822,N_8755,N_8687);
nand U8823 (N_8823,N_8740,N_8643);
xor U8824 (N_8824,N_8623,N_8637);
or U8825 (N_8825,N_8650,N_8692);
nand U8826 (N_8826,N_8642,N_8761);
nor U8827 (N_8827,N_8753,N_8733);
and U8828 (N_8828,N_8689,N_8724);
xnor U8829 (N_8829,N_8728,N_8665);
xor U8830 (N_8830,N_8620,N_8627);
nand U8831 (N_8831,N_8634,N_8647);
or U8832 (N_8832,N_8691,N_8674);
and U8833 (N_8833,N_8677,N_8771);
nand U8834 (N_8834,N_8760,N_8635);
nor U8835 (N_8835,N_8693,N_8618);
nor U8836 (N_8836,N_8745,N_8708);
nand U8837 (N_8837,N_8671,N_8640);
or U8838 (N_8838,N_8655,N_8602);
and U8839 (N_8839,N_8607,N_8645);
nand U8840 (N_8840,N_8667,N_8683);
nor U8841 (N_8841,N_8699,N_8616);
nand U8842 (N_8842,N_8791,N_8639);
xor U8843 (N_8843,N_8744,N_8611);
xor U8844 (N_8844,N_8631,N_8790);
xnor U8845 (N_8845,N_8721,N_8788);
and U8846 (N_8846,N_8723,N_8730);
nand U8847 (N_8847,N_8741,N_8722);
or U8848 (N_8848,N_8609,N_8751);
or U8849 (N_8849,N_8762,N_8613);
xor U8850 (N_8850,N_8653,N_8660);
nand U8851 (N_8851,N_8688,N_8626);
xnor U8852 (N_8852,N_8600,N_8601);
xnor U8853 (N_8853,N_8654,N_8737);
nor U8854 (N_8854,N_8686,N_8664);
xor U8855 (N_8855,N_8782,N_8648);
or U8856 (N_8856,N_8749,N_8612);
xor U8857 (N_8857,N_8670,N_8632);
xnor U8858 (N_8858,N_8731,N_8785);
xor U8859 (N_8859,N_8750,N_8657);
or U8860 (N_8860,N_8661,N_8763);
or U8861 (N_8861,N_8701,N_8796);
xnor U8862 (N_8862,N_8694,N_8684);
or U8863 (N_8863,N_8793,N_8680);
nand U8864 (N_8864,N_8787,N_8685);
and U8865 (N_8865,N_8649,N_8786);
xor U8866 (N_8866,N_8672,N_8646);
xnor U8867 (N_8867,N_8765,N_8629);
xor U8868 (N_8868,N_8713,N_8628);
or U8869 (N_8869,N_8767,N_8604);
or U8870 (N_8870,N_8666,N_8690);
and U8871 (N_8871,N_8705,N_8780);
nand U8872 (N_8872,N_8704,N_8636);
and U8873 (N_8873,N_8718,N_8698);
nor U8874 (N_8874,N_8727,N_8709);
and U8875 (N_8875,N_8603,N_8729);
xor U8876 (N_8876,N_8711,N_8795);
nand U8877 (N_8877,N_8717,N_8781);
and U8878 (N_8878,N_8659,N_8669);
xnor U8879 (N_8879,N_8794,N_8792);
or U8880 (N_8880,N_8641,N_8778);
or U8881 (N_8881,N_8784,N_8605);
nand U8882 (N_8882,N_8614,N_8644);
nor U8883 (N_8883,N_8662,N_8726);
xnor U8884 (N_8884,N_8675,N_8710);
nor U8885 (N_8885,N_8663,N_8769);
nand U8886 (N_8886,N_8624,N_8682);
xnor U8887 (N_8887,N_8656,N_8706);
nor U8888 (N_8888,N_8798,N_8714);
xor U8889 (N_8889,N_8725,N_8754);
and U8890 (N_8890,N_8783,N_8638);
or U8891 (N_8891,N_8625,N_8633);
and U8892 (N_8892,N_8681,N_8608);
nor U8893 (N_8893,N_8610,N_8757);
nor U8894 (N_8894,N_8747,N_8759);
nor U8895 (N_8895,N_8621,N_8679);
nand U8896 (N_8896,N_8743,N_8702);
and U8897 (N_8897,N_8658,N_8700);
nand U8898 (N_8898,N_8774,N_8720);
xor U8899 (N_8899,N_8652,N_8789);
nand U8900 (N_8900,N_8621,N_8657);
nand U8901 (N_8901,N_8725,N_8638);
and U8902 (N_8902,N_8641,N_8708);
and U8903 (N_8903,N_8698,N_8652);
and U8904 (N_8904,N_8797,N_8697);
nor U8905 (N_8905,N_8757,N_8632);
and U8906 (N_8906,N_8652,N_8691);
nor U8907 (N_8907,N_8763,N_8774);
nand U8908 (N_8908,N_8690,N_8775);
nor U8909 (N_8909,N_8701,N_8646);
nand U8910 (N_8910,N_8614,N_8774);
nand U8911 (N_8911,N_8712,N_8654);
xor U8912 (N_8912,N_8706,N_8676);
nand U8913 (N_8913,N_8648,N_8705);
nor U8914 (N_8914,N_8765,N_8618);
nor U8915 (N_8915,N_8675,N_8789);
xnor U8916 (N_8916,N_8744,N_8604);
or U8917 (N_8917,N_8706,N_8793);
nand U8918 (N_8918,N_8613,N_8781);
nand U8919 (N_8919,N_8663,N_8754);
and U8920 (N_8920,N_8762,N_8643);
nor U8921 (N_8921,N_8641,N_8638);
nand U8922 (N_8922,N_8635,N_8643);
and U8923 (N_8923,N_8718,N_8602);
nor U8924 (N_8924,N_8681,N_8658);
nand U8925 (N_8925,N_8621,N_8649);
nor U8926 (N_8926,N_8752,N_8791);
nand U8927 (N_8927,N_8697,N_8787);
and U8928 (N_8928,N_8628,N_8722);
and U8929 (N_8929,N_8755,N_8655);
or U8930 (N_8930,N_8711,N_8609);
nand U8931 (N_8931,N_8654,N_8612);
or U8932 (N_8932,N_8730,N_8758);
xnor U8933 (N_8933,N_8787,N_8744);
and U8934 (N_8934,N_8787,N_8683);
or U8935 (N_8935,N_8722,N_8650);
nand U8936 (N_8936,N_8763,N_8708);
nand U8937 (N_8937,N_8789,N_8705);
or U8938 (N_8938,N_8799,N_8684);
and U8939 (N_8939,N_8750,N_8789);
or U8940 (N_8940,N_8655,N_8761);
or U8941 (N_8941,N_8621,N_8700);
xnor U8942 (N_8942,N_8716,N_8641);
nand U8943 (N_8943,N_8618,N_8668);
nand U8944 (N_8944,N_8726,N_8617);
nor U8945 (N_8945,N_8715,N_8619);
nor U8946 (N_8946,N_8798,N_8726);
or U8947 (N_8947,N_8743,N_8793);
nor U8948 (N_8948,N_8601,N_8642);
nor U8949 (N_8949,N_8710,N_8785);
or U8950 (N_8950,N_8663,N_8759);
nor U8951 (N_8951,N_8793,N_8739);
nor U8952 (N_8952,N_8634,N_8752);
or U8953 (N_8953,N_8706,N_8644);
xor U8954 (N_8954,N_8750,N_8634);
and U8955 (N_8955,N_8605,N_8721);
or U8956 (N_8956,N_8740,N_8711);
nor U8957 (N_8957,N_8722,N_8632);
and U8958 (N_8958,N_8737,N_8795);
or U8959 (N_8959,N_8781,N_8779);
xor U8960 (N_8960,N_8715,N_8719);
xor U8961 (N_8961,N_8618,N_8798);
nand U8962 (N_8962,N_8757,N_8709);
and U8963 (N_8963,N_8666,N_8709);
or U8964 (N_8964,N_8651,N_8739);
or U8965 (N_8965,N_8668,N_8608);
xnor U8966 (N_8966,N_8697,N_8664);
nand U8967 (N_8967,N_8660,N_8673);
xor U8968 (N_8968,N_8702,N_8657);
nand U8969 (N_8969,N_8680,N_8682);
nand U8970 (N_8970,N_8632,N_8707);
and U8971 (N_8971,N_8769,N_8789);
nor U8972 (N_8972,N_8796,N_8751);
nand U8973 (N_8973,N_8658,N_8754);
nand U8974 (N_8974,N_8681,N_8609);
nand U8975 (N_8975,N_8653,N_8766);
xor U8976 (N_8976,N_8737,N_8787);
xnor U8977 (N_8977,N_8600,N_8711);
nand U8978 (N_8978,N_8633,N_8709);
nor U8979 (N_8979,N_8735,N_8656);
and U8980 (N_8980,N_8631,N_8658);
nor U8981 (N_8981,N_8655,N_8735);
nor U8982 (N_8982,N_8725,N_8684);
xor U8983 (N_8983,N_8770,N_8664);
or U8984 (N_8984,N_8794,N_8661);
and U8985 (N_8985,N_8629,N_8658);
nand U8986 (N_8986,N_8730,N_8638);
xor U8987 (N_8987,N_8713,N_8708);
and U8988 (N_8988,N_8774,N_8669);
nor U8989 (N_8989,N_8748,N_8753);
and U8990 (N_8990,N_8600,N_8714);
nor U8991 (N_8991,N_8784,N_8708);
nor U8992 (N_8992,N_8751,N_8667);
and U8993 (N_8993,N_8741,N_8670);
xnor U8994 (N_8994,N_8689,N_8643);
xnor U8995 (N_8995,N_8665,N_8732);
and U8996 (N_8996,N_8769,N_8664);
nand U8997 (N_8997,N_8637,N_8612);
nor U8998 (N_8998,N_8795,N_8630);
and U8999 (N_8999,N_8756,N_8700);
and U9000 (N_9000,N_8902,N_8989);
xnor U9001 (N_9001,N_8827,N_8905);
nand U9002 (N_9002,N_8993,N_8966);
nand U9003 (N_9003,N_8937,N_8988);
nand U9004 (N_9004,N_8978,N_8889);
xnor U9005 (N_9005,N_8810,N_8880);
nor U9006 (N_9006,N_8939,N_8948);
and U9007 (N_9007,N_8938,N_8881);
nor U9008 (N_9008,N_8912,N_8949);
and U9009 (N_9009,N_8932,N_8825);
or U9010 (N_9010,N_8942,N_8903);
and U9011 (N_9011,N_8924,N_8872);
or U9012 (N_9012,N_8958,N_8951);
nor U9013 (N_9013,N_8990,N_8998);
nand U9014 (N_9014,N_8934,N_8830);
nor U9015 (N_9015,N_8960,N_8916);
nor U9016 (N_9016,N_8831,N_8955);
nand U9017 (N_9017,N_8922,N_8931);
or U9018 (N_9018,N_8814,N_8813);
xor U9019 (N_9019,N_8835,N_8879);
nor U9020 (N_9020,N_8962,N_8997);
or U9021 (N_9021,N_8877,N_8908);
and U9022 (N_9022,N_8848,N_8944);
nor U9023 (N_9023,N_8979,N_8929);
nor U9024 (N_9024,N_8809,N_8975);
or U9025 (N_9025,N_8909,N_8984);
nor U9026 (N_9026,N_8833,N_8926);
or U9027 (N_9027,N_8935,N_8928);
nand U9028 (N_9028,N_8952,N_8985);
nor U9029 (N_9029,N_8856,N_8802);
xnor U9030 (N_9030,N_8987,N_8846);
nand U9031 (N_9031,N_8967,N_8900);
or U9032 (N_9032,N_8961,N_8884);
xor U9033 (N_9033,N_8834,N_8826);
and U9034 (N_9034,N_8971,N_8841);
xor U9035 (N_9035,N_8973,N_8849);
or U9036 (N_9036,N_8991,N_8977);
or U9037 (N_9037,N_8890,N_8911);
nand U9038 (N_9038,N_8875,N_8886);
and U9039 (N_9039,N_8950,N_8815);
and U9040 (N_9040,N_8805,N_8898);
or U9041 (N_9041,N_8828,N_8844);
nor U9042 (N_9042,N_8850,N_8906);
xor U9043 (N_9043,N_8843,N_8963);
xnor U9044 (N_9044,N_8918,N_8878);
nor U9045 (N_9045,N_8974,N_8859);
and U9046 (N_9046,N_8839,N_8824);
or U9047 (N_9047,N_8838,N_8804);
and U9048 (N_9048,N_8921,N_8874);
xor U9049 (N_9049,N_8965,N_8959);
xor U9050 (N_9050,N_8980,N_8956);
xnor U9051 (N_9051,N_8837,N_8970);
nor U9052 (N_9052,N_8894,N_8851);
nor U9053 (N_9053,N_8941,N_8917);
xor U9054 (N_9054,N_8891,N_8983);
nor U9055 (N_9055,N_8899,N_8852);
xnor U9056 (N_9056,N_8999,N_8888);
xnor U9057 (N_9057,N_8995,N_8869);
nand U9058 (N_9058,N_8818,N_8883);
and U9059 (N_9059,N_8873,N_8800);
nor U9060 (N_9060,N_8896,N_8822);
nor U9061 (N_9061,N_8871,N_8882);
and U9062 (N_9062,N_8808,N_8914);
nand U9063 (N_9063,N_8933,N_8968);
nand U9064 (N_9064,N_8892,N_8845);
and U9065 (N_9065,N_8847,N_8867);
or U9066 (N_9066,N_8865,N_8863);
and U9067 (N_9067,N_8996,N_8943);
nand U9068 (N_9068,N_8817,N_8901);
and U9069 (N_9069,N_8887,N_8982);
xor U9070 (N_9070,N_8897,N_8806);
nor U9071 (N_9071,N_8930,N_8910);
nor U9072 (N_9072,N_8857,N_8992);
nand U9073 (N_9073,N_8986,N_8940);
or U9074 (N_9074,N_8832,N_8866);
nand U9075 (N_9075,N_8870,N_8860);
nor U9076 (N_9076,N_8981,N_8895);
nor U9077 (N_9077,N_8893,N_8957);
and U9078 (N_9078,N_8821,N_8855);
or U9079 (N_9079,N_8904,N_8936);
or U9080 (N_9080,N_8919,N_8861);
or U9081 (N_9081,N_8858,N_8836);
and U9082 (N_9082,N_8829,N_8820);
nor U9083 (N_9083,N_8864,N_8868);
nand U9084 (N_9084,N_8819,N_8920);
nand U9085 (N_9085,N_8923,N_8842);
nor U9086 (N_9086,N_8946,N_8972);
nor U9087 (N_9087,N_8840,N_8854);
or U9088 (N_9088,N_8811,N_8876);
nor U9089 (N_9089,N_8816,N_8807);
nor U9090 (N_9090,N_8885,N_8925);
xor U9091 (N_9091,N_8823,N_8954);
and U9092 (N_9092,N_8994,N_8803);
xor U9093 (N_9093,N_8964,N_8947);
and U9094 (N_9094,N_8853,N_8945);
and U9095 (N_9095,N_8927,N_8801);
nor U9096 (N_9096,N_8915,N_8976);
and U9097 (N_9097,N_8907,N_8953);
or U9098 (N_9098,N_8913,N_8862);
and U9099 (N_9099,N_8812,N_8969);
or U9100 (N_9100,N_8822,N_8826);
or U9101 (N_9101,N_8942,N_8992);
or U9102 (N_9102,N_8807,N_8898);
and U9103 (N_9103,N_8907,N_8994);
nand U9104 (N_9104,N_8840,N_8832);
nor U9105 (N_9105,N_8843,N_8865);
nor U9106 (N_9106,N_8983,N_8836);
nand U9107 (N_9107,N_8812,N_8878);
nand U9108 (N_9108,N_8801,N_8807);
nor U9109 (N_9109,N_8943,N_8906);
nor U9110 (N_9110,N_8844,N_8889);
nor U9111 (N_9111,N_8817,N_8899);
or U9112 (N_9112,N_8970,N_8825);
or U9113 (N_9113,N_8891,N_8920);
or U9114 (N_9114,N_8866,N_8958);
or U9115 (N_9115,N_8823,N_8894);
or U9116 (N_9116,N_8876,N_8800);
nor U9117 (N_9117,N_8890,N_8807);
nand U9118 (N_9118,N_8901,N_8987);
xnor U9119 (N_9119,N_8852,N_8946);
xnor U9120 (N_9120,N_8896,N_8871);
xor U9121 (N_9121,N_8882,N_8881);
nand U9122 (N_9122,N_8857,N_8985);
xor U9123 (N_9123,N_8959,N_8819);
nor U9124 (N_9124,N_8968,N_8980);
and U9125 (N_9125,N_8901,N_8936);
nand U9126 (N_9126,N_8969,N_8827);
nor U9127 (N_9127,N_8833,N_8908);
and U9128 (N_9128,N_8888,N_8868);
xnor U9129 (N_9129,N_8922,N_8936);
or U9130 (N_9130,N_8971,N_8929);
xor U9131 (N_9131,N_8909,N_8904);
and U9132 (N_9132,N_8862,N_8977);
and U9133 (N_9133,N_8890,N_8953);
nor U9134 (N_9134,N_8931,N_8980);
or U9135 (N_9135,N_8892,N_8953);
xor U9136 (N_9136,N_8988,N_8923);
and U9137 (N_9137,N_8849,N_8897);
or U9138 (N_9138,N_8901,N_8917);
or U9139 (N_9139,N_8998,N_8901);
and U9140 (N_9140,N_8856,N_8922);
and U9141 (N_9141,N_8843,N_8812);
nor U9142 (N_9142,N_8981,N_8915);
xnor U9143 (N_9143,N_8808,N_8935);
nand U9144 (N_9144,N_8910,N_8974);
xnor U9145 (N_9145,N_8898,N_8913);
or U9146 (N_9146,N_8952,N_8955);
xnor U9147 (N_9147,N_8807,N_8981);
nor U9148 (N_9148,N_8960,N_8926);
nor U9149 (N_9149,N_8935,N_8822);
and U9150 (N_9150,N_8837,N_8806);
xor U9151 (N_9151,N_8828,N_8927);
nor U9152 (N_9152,N_8948,N_8995);
or U9153 (N_9153,N_8801,N_8916);
or U9154 (N_9154,N_8964,N_8988);
nand U9155 (N_9155,N_8873,N_8819);
nor U9156 (N_9156,N_8917,N_8813);
nor U9157 (N_9157,N_8932,N_8984);
xor U9158 (N_9158,N_8848,N_8835);
or U9159 (N_9159,N_8994,N_8841);
or U9160 (N_9160,N_8870,N_8904);
or U9161 (N_9161,N_8941,N_8958);
or U9162 (N_9162,N_8970,N_8975);
nor U9163 (N_9163,N_8860,N_8832);
nand U9164 (N_9164,N_8975,N_8950);
nand U9165 (N_9165,N_8977,N_8925);
nand U9166 (N_9166,N_8901,N_8808);
nand U9167 (N_9167,N_8958,N_8807);
or U9168 (N_9168,N_8944,N_8982);
nand U9169 (N_9169,N_8925,N_8808);
and U9170 (N_9170,N_8951,N_8900);
or U9171 (N_9171,N_8820,N_8860);
xnor U9172 (N_9172,N_8927,N_8915);
or U9173 (N_9173,N_8859,N_8861);
xnor U9174 (N_9174,N_8917,N_8929);
nand U9175 (N_9175,N_8875,N_8938);
and U9176 (N_9176,N_8903,N_8848);
nor U9177 (N_9177,N_8982,N_8833);
and U9178 (N_9178,N_8949,N_8915);
xnor U9179 (N_9179,N_8986,N_8887);
xor U9180 (N_9180,N_8823,N_8830);
nand U9181 (N_9181,N_8944,N_8873);
nor U9182 (N_9182,N_8969,N_8816);
and U9183 (N_9183,N_8879,N_8984);
or U9184 (N_9184,N_8871,N_8838);
xor U9185 (N_9185,N_8868,N_8837);
and U9186 (N_9186,N_8929,N_8911);
nor U9187 (N_9187,N_8827,N_8951);
nand U9188 (N_9188,N_8974,N_8971);
nor U9189 (N_9189,N_8966,N_8892);
xnor U9190 (N_9190,N_8887,N_8837);
or U9191 (N_9191,N_8905,N_8928);
nand U9192 (N_9192,N_8996,N_8848);
xnor U9193 (N_9193,N_8962,N_8833);
and U9194 (N_9194,N_8962,N_8941);
or U9195 (N_9195,N_8962,N_8873);
or U9196 (N_9196,N_8845,N_8978);
or U9197 (N_9197,N_8986,N_8902);
or U9198 (N_9198,N_8934,N_8956);
or U9199 (N_9199,N_8828,N_8937);
xor U9200 (N_9200,N_9023,N_9114);
or U9201 (N_9201,N_9060,N_9126);
and U9202 (N_9202,N_9101,N_9070);
nand U9203 (N_9203,N_9152,N_9011);
and U9204 (N_9204,N_9135,N_9032);
or U9205 (N_9205,N_9171,N_9065);
xor U9206 (N_9206,N_9054,N_9165);
or U9207 (N_9207,N_9094,N_9069);
xor U9208 (N_9208,N_9064,N_9052);
nor U9209 (N_9209,N_9156,N_9113);
nor U9210 (N_9210,N_9087,N_9047);
nor U9211 (N_9211,N_9058,N_9166);
nor U9212 (N_9212,N_9116,N_9007);
and U9213 (N_9213,N_9189,N_9012);
or U9214 (N_9214,N_9105,N_9157);
or U9215 (N_9215,N_9084,N_9088);
nor U9216 (N_9216,N_9035,N_9091);
xor U9217 (N_9217,N_9009,N_9083);
or U9218 (N_9218,N_9123,N_9045);
xor U9219 (N_9219,N_9059,N_9042);
xor U9220 (N_9220,N_9085,N_9178);
nor U9221 (N_9221,N_9097,N_9017);
nor U9222 (N_9222,N_9143,N_9075);
nand U9223 (N_9223,N_9079,N_9130);
nor U9224 (N_9224,N_9191,N_9026);
or U9225 (N_9225,N_9112,N_9163);
nor U9226 (N_9226,N_9038,N_9120);
xnor U9227 (N_9227,N_9153,N_9115);
and U9228 (N_9228,N_9076,N_9066);
and U9229 (N_9229,N_9182,N_9024);
or U9230 (N_9230,N_9080,N_9073);
or U9231 (N_9231,N_9129,N_9198);
nor U9232 (N_9232,N_9095,N_9110);
nor U9233 (N_9233,N_9093,N_9179);
and U9234 (N_9234,N_9049,N_9001);
nand U9235 (N_9235,N_9140,N_9159);
or U9236 (N_9236,N_9164,N_9186);
nor U9237 (N_9237,N_9034,N_9193);
xnor U9238 (N_9238,N_9004,N_9127);
or U9239 (N_9239,N_9051,N_9008);
and U9240 (N_9240,N_9148,N_9013);
xnor U9241 (N_9241,N_9025,N_9176);
and U9242 (N_9242,N_9136,N_9072);
nand U9243 (N_9243,N_9133,N_9134);
or U9244 (N_9244,N_9117,N_9003);
nor U9245 (N_9245,N_9173,N_9063);
and U9246 (N_9246,N_9139,N_9188);
nor U9247 (N_9247,N_9138,N_9167);
or U9248 (N_9248,N_9030,N_9041);
and U9249 (N_9249,N_9168,N_9172);
nand U9250 (N_9250,N_9040,N_9096);
and U9251 (N_9251,N_9197,N_9192);
xor U9252 (N_9252,N_9102,N_9108);
nor U9253 (N_9253,N_9183,N_9147);
nand U9254 (N_9254,N_9019,N_9106);
nor U9255 (N_9255,N_9149,N_9196);
nor U9256 (N_9256,N_9014,N_9177);
nor U9257 (N_9257,N_9119,N_9124);
or U9258 (N_9258,N_9081,N_9181);
nor U9259 (N_9259,N_9131,N_9067);
nand U9260 (N_9260,N_9010,N_9078);
xnor U9261 (N_9261,N_9100,N_9174);
xor U9262 (N_9262,N_9111,N_9154);
or U9263 (N_9263,N_9027,N_9053);
and U9264 (N_9264,N_9175,N_9128);
or U9265 (N_9265,N_9155,N_9020);
or U9266 (N_9266,N_9068,N_9016);
or U9267 (N_9267,N_9018,N_9089);
and U9268 (N_9268,N_9169,N_9000);
xor U9269 (N_9269,N_9122,N_9033);
or U9270 (N_9270,N_9057,N_9146);
xnor U9271 (N_9271,N_9046,N_9006);
xor U9272 (N_9272,N_9184,N_9044);
or U9273 (N_9273,N_9002,N_9195);
nand U9274 (N_9274,N_9056,N_9043);
nand U9275 (N_9275,N_9061,N_9185);
xnor U9276 (N_9276,N_9118,N_9107);
and U9277 (N_9277,N_9005,N_9086);
and U9278 (N_9278,N_9048,N_9074);
nand U9279 (N_9279,N_9145,N_9121);
nand U9280 (N_9280,N_9090,N_9103);
and U9281 (N_9281,N_9055,N_9039);
nor U9282 (N_9282,N_9190,N_9142);
nor U9283 (N_9283,N_9132,N_9161);
nand U9284 (N_9284,N_9160,N_9028);
nand U9285 (N_9285,N_9021,N_9092);
nand U9286 (N_9286,N_9125,N_9158);
nand U9287 (N_9287,N_9137,N_9162);
nand U9288 (N_9288,N_9187,N_9109);
and U9289 (N_9289,N_9037,N_9151);
nor U9290 (N_9290,N_9022,N_9170);
nand U9291 (N_9291,N_9098,N_9082);
xnor U9292 (N_9292,N_9150,N_9031);
xor U9293 (N_9293,N_9071,N_9194);
xnor U9294 (N_9294,N_9036,N_9104);
and U9295 (N_9295,N_9099,N_9144);
xnor U9296 (N_9296,N_9050,N_9029);
and U9297 (N_9297,N_9141,N_9199);
nand U9298 (N_9298,N_9180,N_9062);
and U9299 (N_9299,N_9015,N_9077);
xor U9300 (N_9300,N_9132,N_9196);
nor U9301 (N_9301,N_9071,N_9005);
nand U9302 (N_9302,N_9006,N_9014);
nor U9303 (N_9303,N_9048,N_9002);
nor U9304 (N_9304,N_9197,N_9114);
nor U9305 (N_9305,N_9014,N_9096);
nor U9306 (N_9306,N_9099,N_9121);
xnor U9307 (N_9307,N_9057,N_9118);
or U9308 (N_9308,N_9080,N_9001);
xnor U9309 (N_9309,N_9000,N_9109);
nand U9310 (N_9310,N_9109,N_9125);
and U9311 (N_9311,N_9128,N_9013);
nand U9312 (N_9312,N_9137,N_9164);
nand U9313 (N_9313,N_9177,N_9163);
or U9314 (N_9314,N_9004,N_9095);
nand U9315 (N_9315,N_9089,N_9163);
or U9316 (N_9316,N_9036,N_9129);
nor U9317 (N_9317,N_9075,N_9109);
nand U9318 (N_9318,N_9109,N_9004);
nand U9319 (N_9319,N_9102,N_9027);
nand U9320 (N_9320,N_9074,N_9001);
xor U9321 (N_9321,N_9050,N_9096);
xor U9322 (N_9322,N_9050,N_9022);
xnor U9323 (N_9323,N_9046,N_9152);
and U9324 (N_9324,N_9188,N_9168);
and U9325 (N_9325,N_9131,N_9027);
xnor U9326 (N_9326,N_9193,N_9043);
nand U9327 (N_9327,N_9123,N_9062);
xor U9328 (N_9328,N_9131,N_9070);
or U9329 (N_9329,N_9124,N_9002);
nand U9330 (N_9330,N_9147,N_9174);
or U9331 (N_9331,N_9042,N_9147);
nor U9332 (N_9332,N_9190,N_9188);
and U9333 (N_9333,N_9070,N_9001);
or U9334 (N_9334,N_9123,N_9010);
or U9335 (N_9335,N_9170,N_9048);
or U9336 (N_9336,N_9161,N_9159);
or U9337 (N_9337,N_9120,N_9075);
nand U9338 (N_9338,N_9184,N_9118);
nor U9339 (N_9339,N_9144,N_9168);
nand U9340 (N_9340,N_9094,N_9180);
nand U9341 (N_9341,N_9146,N_9145);
nor U9342 (N_9342,N_9125,N_9184);
or U9343 (N_9343,N_9113,N_9106);
nor U9344 (N_9344,N_9051,N_9009);
and U9345 (N_9345,N_9141,N_9041);
and U9346 (N_9346,N_9089,N_9020);
or U9347 (N_9347,N_9139,N_9190);
nand U9348 (N_9348,N_9174,N_9136);
nand U9349 (N_9349,N_9005,N_9108);
nor U9350 (N_9350,N_9143,N_9069);
nand U9351 (N_9351,N_9073,N_9163);
nor U9352 (N_9352,N_9068,N_9059);
nor U9353 (N_9353,N_9096,N_9066);
xor U9354 (N_9354,N_9124,N_9128);
nor U9355 (N_9355,N_9101,N_9025);
nand U9356 (N_9356,N_9048,N_9059);
nand U9357 (N_9357,N_9193,N_9033);
xor U9358 (N_9358,N_9073,N_9077);
and U9359 (N_9359,N_9072,N_9093);
nand U9360 (N_9360,N_9027,N_9045);
or U9361 (N_9361,N_9037,N_9073);
nor U9362 (N_9362,N_9119,N_9062);
nor U9363 (N_9363,N_9121,N_9005);
nand U9364 (N_9364,N_9025,N_9058);
and U9365 (N_9365,N_9119,N_9036);
or U9366 (N_9366,N_9017,N_9108);
nor U9367 (N_9367,N_9194,N_9057);
and U9368 (N_9368,N_9155,N_9062);
nand U9369 (N_9369,N_9171,N_9036);
xor U9370 (N_9370,N_9193,N_9119);
or U9371 (N_9371,N_9003,N_9104);
nor U9372 (N_9372,N_9194,N_9078);
or U9373 (N_9373,N_9163,N_9051);
nor U9374 (N_9374,N_9024,N_9133);
nand U9375 (N_9375,N_9006,N_9044);
or U9376 (N_9376,N_9079,N_9170);
nand U9377 (N_9377,N_9176,N_9194);
xnor U9378 (N_9378,N_9187,N_9028);
and U9379 (N_9379,N_9064,N_9081);
nand U9380 (N_9380,N_9025,N_9131);
nand U9381 (N_9381,N_9030,N_9092);
nor U9382 (N_9382,N_9133,N_9163);
nor U9383 (N_9383,N_9080,N_9175);
or U9384 (N_9384,N_9140,N_9169);
or U9385 (N_9385,N_9199,N_9196);
xnor U9386 (N_9386,N_9102,N_9133);
nand U9387 (N_9387,N_9091,N_9021);
nor U9388 (N_9388,N_9054,N_9052);
or U9389 (N_9389,N_9042,N_9140);
nor U9390 (N_9390,N_9174,N_9068);
xor U9391 (N_9391,N_9164,N_9047);
and U9392 (N_9392,N_9005,N_9097);
and U9393 (N_9393,N_9024,N_9193);
nor U9394 (N_9394,N_9181,N_9104);
and U9395 (N_9395,N_9065,N_9027);
nor U9396 (N_9396,N_9193,N_9112);
and U9397 (N_9397,N_9141,N_9126);
and U9398 (N_9398,N_9186,N_9075);
or U9399 (N_9399,N_9139,N_9048);
nand U9400 (N_9400,N_9225,N_9266);
or U9401 (N_9401,N_9354,N_9209);
and U9402 (N_9402,N_9386,N_9319);
nor U9403 (N_9403,N_9292,N_9206);
xor U9404 (N_9404,N_9372,N_9373);
nand U9405 (N_9405,N_9214,N_9342);
nor U9406 (N_9406,N_9391,N_9326);
xor U9407 (N_9407,N_9339,N_9378);
nand U9408 (N_9408,N_9324,N_9230);
nor U9409 (N_9409,N_9238,N_9335);
or U9410 (N_9410,N_9264,N_9389);
and U9411 (N_9411,N_9345,N_9205);
nor U9412 (N_9412,N_9215,N_9255);
and U9413 (N_9413,N_9229,N_9274);
nor U9414 (N_9414,N_9227,N_9239);
nor U9415 (N_9415,N_9394,N_9341);
and U9416 (N_9416,N_9259,N_9248);
nand U9417 (N_9417,N_9291,N_9396);
or U9418 (N_9418,N_9343,N_9216);
nor U9419 (N_9419,N_9219,N_9382);
xnor U9420 (N_9420,N_9243,N_9320);
or U9421 (N_9421,N_9231,N_9361);
and U9422 (N_9422,N_9217,N_9332);
nand U9423 (N_9423,N_9256,N_9221);
xnor U9424 (N_9424,N_9374,N_9363);
or U9425 (N_9425,N_9375,N_9353);
nor U9426 (N_9426,N_9237,N_9287);
nand U9427 (N_9427,N_9338,N_9397);
xor U9428 (N_9428,N_9285,N_9370);
and U9429 (N_9429,N_9288,N_9220);
nand U9430 (N_9430,N_9351,N_9340);
or U9431 (N_9431,N_9307,N_9312);
nor U9432 (N_9432,N_9384,N_9388);
xor U9433 (N_9433,N_9306,N_9376);
and U9434 (N_9434,N_9327,N_9210);
nor U9435 (N_9435,N_9267,N_9395);
and U9436 (N_9436,N_9222,N_9289);
nand U9437 (N_9437,N_9301,N_9311);
or U9438 (N_9438,N_9250,N_9202);
xnor U9439 (N_9439,N_9295,N_9357);
or U9440 (N_9440,N_9317,N_9276);
nand U9441 (N_9441,N_9201,N_9365);
nand U9442 (N_9442,N_9269,N_9280);
nor U9443 (N_9443,N_9393,N_9241);
nand U9444 (N_9444,N_9294,N_9275);
xnor U9445 (N_9445,N_9242,N_9359);
xor U9446 (N_9446,N_9337,N_9253);
and U9447 (N_9447,N_9352,N_9358);
nor U9448 (N_9448,N_9286,N_9371);
nand U9449 (N_9449,N_9297,N_9387);
nand U9450 (N_9450,N_9362,N_9380);
xnor U9451 (N_9451,N_9279,N_9218);
and U9452 (N_9452,N_9245,N_9398);
or U9453 (N_9453,N_9329,N_9315);
nor U9454 (N_9454,N_9235,N_9223);
and U9455 (N_9455,N_9270,N_9244);
nor U9456 (N_9456,N_9257,N_9344);
nand U9457 (N_9457,N_9200,N_9268);
nor U9458 (N_9458,N_9261,N_9355);
nand U9459 (N_9459,N_9313,N_9302);
nand U9460 (N_9460,N_9258,N_9272);
xnor U9461 (N_9461,N_9381,N_9316);
nand U9462 (N_9462,N_9325,N_9390);
nand U9463 (N_9463,N_9299,N_9273);
nand U9464 (N_9464,N_9318,N_9203);
or U9465 (N_9465,N_9207,N_9265);
and U9466 (N_9466,N_9271,N_9364);
nor U9467 (N_9467,N_9314,N_9369);
or U9468 (N_9468,N_9212,N_9377);
xnor U9469 (N_9469,N_9254,N_9226);
or U9470 (N_9470,N_9366,N_9356);
nor U9471 (N_9471,N_9346,N_9336);
nor U9472 (N_9472,N_9304,N_9350);
nand U9473 (N_9473,N_9211,N_9208);
and U9474 (N_9474,N_9300,N_9309);
nor U9475 (N_9475,N_9305,N_9290);
nand U9476 (N_9476,N_9281,N_9263);
and U9477 (N_9477,N_9233,N_9349);
and U9478 (N_9478,N_9334,N_9368);
or U9479 (N_9479,N_9252,N_9240);
nor U9480 (N_9480,N_9367,N_9234);
or U9481 (N_9481,N_9379,N_9330);
or U9482 (N_9482,N_9282,N_9322);
and U9483 (N_9483,N_9303,N_9298);
nand U9484 (N_9484,N_9347,N_9385);
or U9485 (N_9485,N_9399,N_9308);
or U9486 (N_9486,N_9224,N_9284);
xnor U9487 (N_9487,N_9260,N_9246);
or U9488 (N_9488,N_9262,N_9247);
and U9489 (N_9489,N_9328,N_9360);
and U9490 (N_9490,N_9228,N_9232);
nand U9491 (N_9491,N_9331,N_9293);
nand U9492 (N_9492,N_9323,N_9383);
nand U9493 (N_9493,N_9249,N_9283);
or U9494 (N_9494,N_9251,N_9236);
xor U9495 (N_9495,N_9277,N_9213);
or U9496 (N_9496,N_9296,N_9333);
or U9497 (N_9497,N_9321,N_9348);
nand U9498 (N_9498,N_9278,N_9204);
nand U9499 (N_9499,N_9392,N_9310);
and U9500 (N_9500,N_9238,N_9280);
nor U9501 (N_9501,N_9299,N_9292);
nor U9502 (N_9502,N_9241,N_9331);
or U9503 (N_9503,N_9244,N_9347);
nand U9504 (N_9504,N_9330,N_9361);
and U9505 (N_9505,N_9230,N_9333);
and U9506 (N_9506,N_9342,N_9375);
xnor U9507 (N_9507,N_9282,N_9352);
nor U9508 (N_9508,N_9389,N_9283);
or U9509 (N_9509,N_9332,N_9287);
and U9510 (N_9510,N_9258,N_9347);
or U9511 (N_9511,N_9323,N_9346);
and U9512 (N_9512,N_9342,N_9353);
and U9513 (N_9513,N_9355,N_9329);
or U9514 (N_9514,N_9244,N_9233);
and U9515 (N_9515,N_9280,N_9360);
xor U9516 (N_9516,N_9215,N_9392);
or U9517 (N_9517,N_9224,N_9263);
and U9518 (N_9518,N_9234,N_9209);
or U9519 (N_9519,N_9296,N_9347);
xor U9520 (N_9520,N_9300,N_9320);
nor U9521 (N_9521,N_9361,N_9305);
or U9522 (N_9522,N_9208,N_9331);
nand U9523 (N_9523,N_9355,N_9273);
or U9524 (N_9524,N_9248,N_9213);
nand U9525 (N_9525,N_9398,N_9256);
or U9526 (N_9526,N_9274,N_9317);
xnor U9527 (N_9527,N_9361,N_9325);
and U9528 (N_9528,N_9294,N_9224);
xnor U9529 (N_9529,N_9359,N_9304);
nand U9530 (N_9530,N_9374,N_9294);
xor U9531 (N_9531,N_9334,N_9242);
xnor U9532 (N_9532,N_9353,N_9372);
nand U9533 (N_9533,N_9377,N_9342);
xor U9534 (N_9534,N_9318,N_9276);
or U9535 (N_9535,N_9205,N_9317);
or U9536 (N_9536,N_9238,N_9217);
or U9537 (N_9537,N_9211,N_9210);
nor U9538 (N_9538,N_9296,N_9357);
xnor U9539 (N_9539,N_9303,N_9253);
nand U9540 (N_9540,N_9258,N_9232);
nand U9541 (N_9541,N_9246,N_9377);
and U9542 (N_9542,N_9328,N_9312);
or U9543 (N_9543,N_9283,N_9373);
and U9544 (N_9544,N_9291,N_9266);
nor U9545 (N_9545,N_9370,N_9332);
nor U9546 (N_9546,N_9228,N_9289);
and U9547 (N_9547,N_9374,N_9225);
nor U9548 (N_9548,N_9221,N_9314);
nand U9549 (N_9549,N_9233,N_9203);
nor U9550 (N_9550,N_9265,N_9312);
or U9551 (N_9551,N_9221,N_9263);
nor U9552 (N_9552,N_9271,N_9260);
and U9553 (N_9553,N_9337,N_9254);
or U9554 (N_9554,N_9313,N_9319);
or U9555 (N_9555,N_9366,N_9343);
and U9556 (N_9556,N_9205,N_9390);
and U9557 (N_9557,N_9369,N_9382);
nand U9558 (N_9558,N_9340,N_9311);
and U9559 (N_9559,N_9369,N_9308);
and U9560 (N_9560,N_9229,N_9240);
xor U9561 (N_9561,N_9210,N_9295);
or U9562 (N_9562,N_9299,N_9310);
and U9563 (N_9563,N_9249,N_9354);
nor U9564 (N_9564,N_9268,N_9348);
and U9565 (N_9565,N_9375,N_9303);
or U9566 (N_9566,N_9216,N_9370);
and U9567 (N_9567,N_9338,N_9204);
xor U9568 (N_9568,N_9308,N_9268);
nand U9569 (N_9569,N_9392,N_9384);
xnor U9570 (N_9570,N_9297,N_9227);
and U9571 (N_9571,N_9371,N_9212);
nor U9572 (N_9572,N_9396,N_9337);
nand U9573 (N_9573,N_9258,N_9242);
and U9574 (N_9574,N_9331,N_9276);
nand U9575 (N_9575,N_9368,N_9388);
nor U9576 (N_9576,N_9382,N_9335);
xnor U9577 (N_9577,N_9269,N_9312);
nand U9578 (N_9578,N_9371,N_9283);
xnor U9579 (N_9579,N_9269,N_9359);
and U9580 (N_9580,N_9215,N_9328);
and U9581 (N_9581,N_9214,N_9266);
nor U9582 (N_9582,N_9208,N_9312);
xnor U9583 (N_9583,N_9350,N_9285);
xor U9584 (N_9584,N_9235,N_9293);
nor U9585 (N_9585,N_9202,N_9364);
nor U9586 (N_9586,N_9216,N_9387);
and U9587 (N_9587,N_9392,N_9334);
nand U9588 (N_9588,N_9366,N_9331);
xor U9589 (N_9589,N_9272,N_9389);
nor U9590 (N_9590,N_9286,N_9372);
or U9591 (N_9591,N_9203,N_9259);
or U9592 (N_9592,N_9342,N_9324);
and U9593 (N_9593,N_9324,N_9304);
or U9594 (N_9594,N_9231,N_9364);
and U9595 (N_9595,N_9256,N_9389);
xor U9596 (N_9596,N_9206,N_9300);
or U9597 (N_9597,N_9267,N_9325);
and U9598 (N_9598,N_9261,N_9377);
xor U9599 (N_9599,N_9362,N_9236);
and U9600 (N_9600,N_9518,N_9409);
nor U9601 (N_9601,N_9529,N_9422);
nor U9602 (N_9602,N_9507,N_9432);
nand U9603 (N_9603,N_9462,N_9512);
xor U9604 (N_9604,N_9550,N_9571);
xnor U9605 (N_9605,N_9481,N_9514);
nor U9606 (N_9606,N_9584,N_9457);
and U9607 (N_9607,N_9505,N_9577);
nand U9608 (N_9608,N_9598,N_9458);
or U9609 (N_9609,N_9542,N_9556);
nand U9610 (N_9610,N_9434,N_9403);
xor U9611 (N_9611,N_9410,N_9506);
xnor U9612 (N_9612,N_9450,N_9472);
and U9613 (N_9613,N_9561,N_9499);
nand U9614 (N_9614,N_9420,N_9504);
xnor U9615 (N_9615,N_9595,N_9401);
nand U9616 (N_9616,N_9549,N_9438);
nor U9617 (N_9617,N_9439,N_9490);
or U9618 (N_9618,N_9528,N_9485);
xor U9619 (N_9619,N_9452,N_9510);
or U9620 (N_9620,N_9560,N_9597);
or U9621 (N_9621,N_9535,N_9574);
xnor U9622 (N_9622,N_9592,N_9565);
and U9623 (N_9623,N_9520,N_9516);
nand U9624 (N_9624,N_9469,N_9407);
nor U9625 (N_9625,N_9412,N_9473);
or U9626 (N_9626,N_9415,N_9443);
and U9627 (N_9627,N_9447,N_9502);
nor U9628 (N_9628,N_9468,N_9495);
and U9629 (N_9629,N_9475,N_9425);
nor U9630 (N_9630,N_9427,N_9444);
nand U9631 (N_9631,N_9416,N_9527);
and U9632 (N_9632,N_9503,N_9579);
nand U9633 (N_9633,N_9460,N_9523);
or U9634 (N_9634,N_9451,N_9467);
and U9635 (N_9635,N_9446,N_9546);
nor U9636 (N_9636,N_9539,N_9586);
and U9637 (N_9637,N_9570,N_9572);
nor U9638 (N_9638,N_9406,N_9448);
nor U9639 (N_9639,N_9531,N_9538);
xor U9640 (N_9640,N_9559,N_9479);
nor U9641 (N_9641,N_9449,N_9508);
nor U9642 (N_9642,N_9594,N_9522);
xnor U9643 (N_9643,N_9567,N_9429);
and U9644 (N_9644,N_9513,N_9402);
nand U9645 (N_9645,N_9515,N_9590);
nand U9646 (N_9646,N_9445,N_9562);
or U9647 (N_9647,N_9541,N_9424);
or U9648 (N_9648,N_9436,N_9545);
or U9649 (N_9649,N_9430,N_9509);
and U9650 (N_9650,N_9471,N_9587);
nand U9651 (N_9651,N_9431,N_9593);
nand U9652 (N_9652,N_9551,N_9552);
nand U9653 (N_9653,N_9440,N_9575);
and U9654 (N_9654,N_9532,N_9500);
xor U9655 (N_9655,N_9476,N_9578);
xnor U9656 (N_9656,N_9465,N_9573);
nand U9657 (N_9657,N_9489,N_9453);
nor U9658 (N_9658,N_9461,N_9404);
nor U9659 (N_9659,N_9470,N_9580);
xnor U9660 (N_9660,N_9482,N_9493);
and U9661 (N_9661,N_9558,N_9498);
and U9662 (N_9662,N_9501,N_9414);
and U9663 (N_9663,N_9525,N_9413);
nor U9664 (N_9664,N_9477,N_9588);
xnor U9665 (N_9665,N_9437,N_9543);
and U9666 (N_9666,N_9524,N_9599);
and U9667 (N_9667,N_9442,N_9418);
and U9668 (N_9668,N_9585,N_9486);
nand U9669 (N_9669,N_9517,N_9530);
or U9670 (N_9670,N_9555,N_9478);
nor U9671 (N_9671,N_9576,N_9540);
or U9672 (N_9672,N_9488,N_9497);
xor U9673 (N_9673,N_9534,N_9426);
and U9674 (N_9674,N_9408,N_9480);
xnor U9675 (N_9675,N_9405,N_9564);
xnor U9676 (N_9676,N_9554,N_9466);
nand U9677 (N_9677,N_9544,N_9496);
xor U9678 (N_9678,N_9582,N_9563);
nand U9679 (N_9679,N_9581,N_9474);
xnor U9680 (N_9680,N_9456,N_9533);
nor U9681 (N_9681,N_9537,N_9400);
nand U9682 (N_9682,N_9583,N_9568);
nand U9683 (N_9683,N_9553,N_9435);
nand U9684 (N_9684,N_9483,N_9494);
nor U9685 (N_9685,N_9411,N_9596);
nor U9686 (N_9686,N_9566,N_9454);
xor U9687 (N_9687,N_9547,N_9464);
nor U9688 (N_9688,N_9548,N_9521);
xnor U9689 (N_9689,N_9419,N_9492);
xnor U9690 (N_9690,N_9433,N_9441);
nor U9691 (N_9691,N_9455,N_9591);
or U9692 (N_9692,N_9417,N_9589);
xnor U9693 (N_9693,N_9463,N_9526);
nand U9694 (N_9694,N_9491,N_9519);
nand U9695 (N_9695,N_9557,N_9421);
and U9696 (N_9696,N_9511,N_9536);
nand U9697 (N_9697,N_9459,N_9569);
nand U9698 (N_9698,N_9487,N_9428);
nand U9699 (N_9699,N_9423,N_9484);
or U9700 (N_9700,N_9522,N_9523);
or U9701 (N_9701,N_9425,N_9579);
nand U9702 (N_9702,N_9422,N_9453);
nand U9703 (N_9703,N_9507,N_9400);
xor U9704 (N_9704,N_9421,N_9450);
xnor U9705 (N_9705,N_9496,N_9435);
nand U9706 (N_9706,N_9446,N_9498);
or U9707 (N_9707,N_9450,N_9569);
nor U9708 (N_9708,N_9582,N_9454);
nor U9709 (N_9709,N_9476,N_9454);
nor U9710 (N_9710,N_9549,N_9519);
nor U9711 (N_9711,N_9428,N_9512);
nand U9712 (N_9712,N_9597,N_9582);
xnor U9713 (N_9713,N_9503,N_9580);
nand U9714 (N_9714,N_9450,N_9418);
nand U9715 (N_9715,N_9514,N_9448);
nor U9716 (N_9716,N_9564,N_9455);
and U9717 (N_9717,N_9400,N_9500);
and U9718 (N_9718,N_9480,N_9535);
nand U9719 (N_9719,N_9458,N_9432);
nand U9720 (N_9720,N_9550,N_9596);
nand U9721 (N_9721,N_9546,N_9531);
and U9722 (N_9722,N_9407,N_9529);
nand U9723 (N_9723,N_9590,N_9580);
nor U9724 (N_9724,N_9466,N_9595);
xnor U9725 (N_9725,N_9586,N_9571);
nand U9726 (N_9726,N_9421,N_9497);
nor U9727 (N_9727,N_9421,N_9490);
and U9728 (N_9728,N_9454,N_9530);
xor U9729 (N_9729,N_9505,N_9482);
or U9730 (N_9730,N_9438,N_9500);
nor U9731 (N_9731,N_9563,N_9440);
xor U9732 (N_9732,N_9585,N_9471);
and U9733 (N_9733,N_9538,N_9567);
nand U9734 (N_9734,N_9465,N_9414);
or U9735 (N_9735,N_9567,N_9532);
nor U9736 (N_9736,N_9525,N_9414);
and U9737 (N_9737,N_9450,N_9411);
xnor U9738 (N_9738,N_9583,N_9466);
or U9739 (N_9739,N_9515,N_9523);
xnor U9740 (N_9740,N_9452,N_9492);
nand U9741 (N_9741,N_9477,N_9553);
and U9742 (N_9742,N_9529,N_9497);
nand U9743 (N_9743,N_9546,N_9401);
nor U9744 (N_9744,N_9513,N_9413);
or U9745 (N_9745,N_9544,N_9450);
and U9746 (N_9746,N_9525,N_9568);
xor U9747 (N_9747,N_9555,N_9464);
nand U9748 (N_9748,N_9472,N_9499);
or U9749 (N_9749,N_9551,N_9540);
xnor U9750 (N_9750,N_9409,N_9592);
nor U9751 (N_9751,N_9433,N_9527);
nand U9752 (N_9752,N_9411,N_9530);
or U9753 (N_9753,N_9589,N_9521);
nor U9754 (N_9754,N_9488,N_9566);
nand U9755 (N_9755,N_9507,N_9525);
xor U9756 (N_9756,N_9585,N_9590);
and U9757 (N_9757,N_9515,N_9532);
nor U9758 (N_9758,N_9436,N_9403);
or U9759 (N_9759,N_9587,N_9528);
xnor U9760 (N_9760,N_9521,N_9425);
or U9761 (N_9761,N_9559,N_9594);
nand U9762 (N_9762,N_9555,N_9463);
nor U9763 (N_9763,N_9492,N_9457);
or U9764 (N_9764,N_9592,N_9560);
xnor U9765 (N_9765,N_9441,N_9430);
and U9766 (N_9766,N_9506,N_9413);
xnor U9767 (N_9767,N_9542,N_9442);
nand U9768 (N_9768,N_9447,N_9434);
nand U9769 (N_9769,N_9435,N_9535);
xor U9770 (N_9770,N_9508,N_9594);
nor U9771 (N_9771,N_9472,N_9402);
or U9772 (N_9772,N_9479,N_9500);
nand U9773 (N_9773,N_9557,N_9441);
nor U9774 (N_9774,N_9583,N_9548);
xor U9775 (N_9775,N_9413,N_9495);
nand U9776 (N_9776,N_9497,N_9414);
nor U9777 (N_9777,N_9432,N_9464);
or U9778 (N_9778,N_9535,N_9506);
xnor U9779 (N_9779,N_9582,N_9479);
xor U9780 (N_9780,N_9472,N_9572);
or U9781 (N_9781,N_9520,N_9488);
or U9782 (N_9782,N_9400,N_9445);
and U9783 (N_9783,N_9506,N_9455);
nand U9784 (N_9784,N_9501,N_9590);
and U9785 (N_9785,N_9468,N_9504);
xor U9786 (N_9786,N_9435,N_9541);
xnor U9787 (N_9787,N_9464,N_9485);
or U9788 (N_9788,N_9407,N_9426);
nor U9789 (N_9789,N_9537,N_9441);
or U9790 (N_9790,N_9592,N_9400);
nand U9791 (N_9791,N_9516,N_9505);
nand U9792 (N_9792,N_9466,N_9557);
nor U9793 (N_9793,N_9433,N_9507);
nand U9794 (N_9794,N_9417,N_9527);
nand U9795 (N_9795,N_9581,N_9455);
and U9796 (N_9796,N_9400,N_9518);
xnor U9797 (N_9797,N_9560,N_9463);
nor U9798 (N_9798,N_9584,N_9505);
xnor U9799 (N_9799,N_9538,N_9506);
nand U9800 (N_9800,N_9746,N_9726);
xor U9801 (N_9801,N_9635,N_9642);
nor U9802 (N_9802,N_9732,N_9723);
or U9803 (N_9803,N_9651,N_9680);
or U9804 (N_9804,N_9637,N_9631);
and U9805 (N_9805,N_9662,N_9724);
or U9806 (N_9806,N_9793,N_9773);
nand U9807 (N_9807,N_9789,N_9760);
xor U9808 (N_9808,N_9739,N_9627);
xor U9809 (N_9809,N_9671,N_9757);
nor U9810 (N_9810,N_9645,N_9759);
and U9811 (N_9811,N_9738,N_9737);
nand U9812 (N_9812,N_9669,N_9753);
nand U9813 (N_9813,N_9626,N_9649);
nor U9814 (N_9814,N_9703,N_9766);
nand U9815 (N_9815,N_9608,N_9799);
nor U9816 (N_9816,N_9691,N_9657);
nand U9817 (N_9817,N_9707,N_9785);
and U9818 (N_9818,N_9733,N_9767);
nor U9819 (N_9819,N_9603,N_9743);
or U9820 (N_9820,N_9659,N_9718);
or U9821 (N_9821,N_9774,N_9663);
or U9822 (N_9822,N_9758,N_9613);
nor U9823 (N_9823,N_9770,N_9678);
nand U9824 (N_9824,N_9742,N_9639);
nand U9825 (N_9825,N_9648,N_9752);
or U9826 (N_9826,N_9750,N_9735);
and U9827 (N_9827,N_9617,N_9775);
xnor U9828 (N_9828,N_9690,N_9778);
or U9829 (N_9829,N_9683,N_9621);
xor U9830 (N_9830,N_9688,N_9640);
or U9831 (N_9831,N_9708,N_9730);
or U9832 (N_9832,N_9716,N_9780);
and U9833 (N_9833,N_9655,N_9611);
or U9834 (N_9834,N_9777,N_9720);
xnor U9835 (N_9835,N_9646,N_9784);
xnor U9836 (N_9836,N_9692,N_9764);
nor U9837 (N_9837,N_9795,N_9763);
nor U9838 (N_9838,N_9729,N_9634);
nor U9839 (N_9839,N_9628,N_9771);
and U9840 (N_9840,N_9652,N_9694);
nand U9841 (N_9841,N_9790,N_9673);
or U9842 (N_9842,N_9705,N_9765);
xor U9843 (N_9843,N_9674,N_9736);
and U9844 (N_9844,N_9658,N_9769);
nand U9845 (N_9845,N_9792,N_9641);
and U9846 (N_9846,N_9682,N_9786);
nor U9847 (N_9847,N_9689,N_9740);
or U9848 (N_9848,N_9711,N_9679);
nand U9849 (N_9849,N_9699,N_9782);
or U9850 (N_9850,N_9632,N_9653);
nand U9851 (N_9851,N_9706,N_9670);
nand U9852 (N_9852,N_9768,N_9638);
and U9853 (N_9853,N_9664,N_9700);
nand U9854 (N_9854,N_9636,N_9610);
nor U9855 (N_9855,N_9614,N_9693);
or U9856 (N_9856,N_9668,N_9776);
and U9857 (N_9857,N_9791,N_9719);
xor U9858 (N_9858,N_9630,N_9676);
xor U9859 (N_9859,N_9675,N_9715);
xnor U9860 (N_9860,N_9687,N_9747);
nand U9861 (N_9861,N_9697,N_9606);
xnor U9862 (N_9862,N_9686,N_9798);
nor U9863 (N_9863,N_9756,N_9623);
nor U9864 (N_9864,N_9744,N_9788);
nand U9865 (N_9865,N_9787,N_9600);
xnor U9866 (N_9866,N_9619,N_9731);
nor U9867 (N_9867,N_9762,N_9751);
or U9868 (N_9868,N_9712,N_9644);
or U9869 (N_9869,N_9772,N_9710);
xor U9870 (N_9870,N_9761,N_9681);
and U9871 (N_9871,N_9783,N_9695);
nand U9872 (N_9872,N_9755,N_9741);
xnor U9873 (N_9873,N_9615,N_9704);
xor U9874 (N_9874,N_9633,N_9725);
or U9875 (N_9875,N_9666,N_9721);
nand U9876 (N_9876,N_9605,N_9643);
and U9877 (N_9877,N_9650,N_9624);
and U9878 (N_9878,N_9722,N_9647);
nor U9879 (N_9879,N_9714,N_9797);
and U9880 (N_9880,N_9734,N_9698);
and U9881 (N_9881,N_9656,N_9748);
or U9882 (N_9882,N_9749,N_9701);
nand U9883 (N_9883,N_9745,N_9654);
xnor U9884 (N_9884,N_9696,N_9713);
or U9885 (N_9885,N_9684,N_9667);
and U9886 (N_9886,N_9609,N_9604);
or U9887 (N_9887,N_9728,N_9629);
nor U9888 (N_9888,N_9661,N_9622);
or U9889 (N_9889,N_9754,N_9618);
nand U9890 (N_9890,N_9612,N_9781);
xnor U9891 (N_9891,N_9685,N_9602);
and U9892 (N_9892,N_9601,N_9620);
xnor U9893 (N_9893,N_9665,N_9779);
or U9894 (N_9894,N_9672,N_9702);
and U9895 (N_9895,N_9794,N_9616);
and U9896 (N_9896,N_9709,N_9796);
and U9897 (N_9897,N_9625,N_9660);
nor U9898 (N_9898,N_9727,N_9677);
nand U9899 (N_9899,N_9717,N_9607);
nand U9900 (N_9900,N_9656,N_9786);
or U9901 (N_9901,N_9625,N_9771);
nand U9902 (N_9902,N_9656,N_9639);
and U9903 (N_9903,N_9776,N_9655);
xnor U9904 (N_9904,N_9665,N_9663);
or U9905 (N_9905,N_9749,N_9636);
nor U9906 (N_9906,N_9763,N_9751);
xnor U9907 (N_9907,N_9764,N_9699);
or U9908 (N_9908,N_9709,N_9721);
nand U9909 (N_9909,N_9676,N_9677);
nor U9910 (N_9910,N_9720,N_9722);
xnor U9911 (N_9911,N_9696,N_9786);
nor U9912 (N_9912,N_9792,N_9717);
xnor U9913 (N_9913,N_9730,N_9729);
nand U9914 (N_9914,N_9736,N_9672);
nand U9915 (N_9915,N_9765,N_9652);
or U9916 (N_9916,N_9738,N_9774);
xor U9917 (N_9917,N_9632,N_9770);
nor U9918 (N_9918,N_9726,N_9615);
xnor U9919 (N_9919,N_9706,N_9788);
or U9920 (N_9920,N_9636,N_9614);
nand U9921 (N_9921,N_9688,N_9785);
and U9922 (N_9922,N_9697,N_9685);
and U9923 (N_9923,N_9788,N_9668);
nand U9924 (N_9924,N_9761,N_9653);
or U9925 (N_9925,N_9790,N_9669);
nand U9926 (N_9926,N_9748,N_9672);
nand U9927 (N_9927,N_9672,N_9779);
or U9928 (N_9928,N_9673,N_9753);
nor U9929 (N_9929,N_9754,N_9789);
xnor U9930 (N_9930,N_9781,N_9751);
nor U9931 (N_9931,N_9618,N_9605);
nor U9932 (N_9932,N_9653,N_9757);
xor U9933 (N_9933,N_9617,N_9639);
nand U9934 (N_9934,N_9765,N_9618);
or U9935 (N_9935,N_9686,N_9764);
and U9936 (N_9936,N_9646,N_9757);
and U9937 (N_9937,N_9730,N_9704);
xor U9938 (N_9938,N_9643,N_9671);
nor U9939 (N_9939,N_9671,N_9651);
or U9940 (N_9940,N_9778,N_9733);
or U9941 (N_9941,N_9600,N_9739);
and U9942 (N_9942,N_9725,N_9631);
and U9943 (N_9943,N_9756,N_9736);
nor U9944 (N_9944,N_9665,N_9712);
or U9945 (N_9945,N_9648,N_9638);
nand U9946 (N_9946,N_9746,N_9620);
nor U9947 (N_9947,N_9709,N_9749);
and U9948 (N_9948,N_9758,N_9604);
and U9949 (N_9949,N_9776,N_9677);
and U9950 (N_9950,N_9785,N_9646);
xor U9951 (N_9951,N_9692,N_9631);
nor U9952 (N_9952,N_9723,N_9716);
nor U9953 (N_9953,N_9638,N_9601);
nand U9954 (N_9954,N_9710,N_9611);
and U9955 (N_9955,N_9732,N_9649);
xnor U9956 (N_9956,N_9726,N_9734);
or U9957 (N_9957,N_9785,N_9744);
nand U9958 (N_9958,N_9626,N_9655);
or U9959 (N_9959,N_9649,N_9652);
and U9960 (N_9960,N_9763,N_9692);
xor U9961 (N_9961,N_9722,N_9766);
nor U9962 (N_9962,N_9721,N_9674);
xnor U9963 (N_9963,N_9680,N_9620);
nand U9964 (N_9964,N_9798,N_9629);
and U9965 (N_9965,N_9720,N_9698);
xor U9966 (N_9966,N_9701,N_9714);
or U9967 (N_9967,N_9703,N_9608);
xor U9968 (N_9968,N_9754,N_9735);
nand U9969 (N_9969,N_9629,N_9610);
nand U9970 (N_9970,N_9798,N_9662);
nor U9971 (N_9971,N_9687,N_9715);
and U9972 (N_9972,N_9709,N_9791);
xor U9973 (N_9973,N_9657,N_9667);
or U9974 (N_9974,N_9776,N_9741);
nand U9975 (N_9975,N_9625,N_9730);
nor U9976 (N_9976,N_9645,N_9607);
xnor U9977 (N_9977,N_9716,N_9750);
nand U9978 (N_9978,N_9700,N_9790);
xor U9979 (N_9979,N_9751,N_9776);
or U9980 (N_9980,N_9662,N_9634);
and U9981 (N_9981,N_9703,N_9710);
or U9982 (N_9982,N_9735,N_9725);
or U9983 (N_9983,N_9796,N_9723);
nor U9984 (N_9984,N_9777,N_9692);
and U9985 (N_9985,N_9623,N_9687);
nand U9986 (N_9986,N_9648,N_9699);
xor U9987 (N_9987,N_9650,N_9724);
and U9988 (N_9988,N_9785,N_9602);
xnor U9989 (N_9989,N_9631,N_9709);
or U9990 (N_9990,N_9692,N_9693);
nor U9991 (N_9991,N_9711,N_9768);
xnor U9992 (N_9992,N_9761,N_9784);
nor U9993 (N_9993,N_9658,N_9720);
nor U9994 (N_9994,N_9755,N_9672);
nand U9995 (N_9995,N_9725,N_9606);
nor U9996 (N_9996,N_9639,N_9778);
and U9997 (N_9997,N_9741,N_9610);
or U9998 (N_9998,N_9709,N_9794);
or U9999 (N_9999,N_9777,N_9748);
xnor U10000 (N_10000,N_9976,N_9801);
nor U10001 (N_10001,N_9980,N_9878);
nor U10002 (N_10002,N_9897,N_9830);
xor U10003 (N_10003,N_9983,N_9853);
nor U10004 (N_10004,N_9968,N_9925);
nand U10005 (N_10005,N_9867,N_9935);
xnor U10006 (N_10006,N_9871,N_9919);
nor U10007 (N_10007,N_9836,N_9906);
and U10008 (N_10008,N_9900,N_9859);
xnor U10009 (N_10009,N_9842,N_9892);
nor U10010 (N_10010,N_9991,N_9927);
and U10011 (N_10011,N_9889,N_9974);
or U10012 (N_10012,N_9998,N_9813);
and U10013 (N_10013,N_9939,N_9808);
nor U10014 (N_10014,N_9885,N_9929);
or U10015 (N_10015,N_9967,N_9891);
xor U10016 (N_10016,N_9922,N_9958);
nand U10017 (N_10017,N_9961,N_9923);
or U10018 (N_10018,N_9843,N_9916);
nor U10019 (N_10019,N_9896,N_9966);
xnor U10020 (N_10020,N_9821,N_9827);
nand U10021 (N_10021,N_9982,N_9999);
nor U10022 (N_10022,N_9936,N_9815);
nor U10023 (N_10023,N_9819,N_9933);
nor U10024 (N_10024,N_9901,N_9829);
nand U10025 (N_10025,N_9838,N_9873);
nor U10026 (N_10026,N_9818,N_9930);
nand U10027 (N_10027,N_9835,N_9811);
xnor U10028 (N_10028,N_9810,N_9984);
nand U10029 (N_10029,N_9945,N_9806);
xnor U10030 (N_10030,N_9877,N_9911);
xnor U10031 (N_10031,N_9940,N_9937);
and U10032 (N_10032,N_9855,N_9832);
nand U10033 (N_10033,N_9890,N_9826);
nor U10034 (N_10034,N_9860,N_9865);
or U10035 (N_10035,N_9938,N_9975);
or U10036 (N_10036,N_9841,N_9944);
or U10037 (N_10037,N_9977,N_9817);
nor U10038 (N_10038,N_9893,N_9963);
xnor U10039 (N_10039,N_9948,N_9912);
nor U10040 (N_10040,N_9844,N_9972);
xnor U10041 (N_10041,N_9883,N_9899);
nor U10042 (N_10042,N_9803,N_9898);
nand U10043 (N_10043,N_9941,N_9874);
xor U10044 (N_10044,N_9834,N_9852);
xnor U10045 (N_10045,N_9954,N_9887);
nand U10046 (N_10046,N_9971,N_9913);
nand U10047 (N_10047,N_9875,N_9847);
or U10048 (N_10048,N_9840,N_9845);
and U10049 (N_10049,N_9986,N_9942);
xnor U10050 (N_10050,N_9992,N_9869);
and U10051 (N_10051,N_9820,N_9988);
nand U10052 (N_10052,N_9969,N_9850);
and U10053 (N_10053,N_9864,N_9962);
or U10054 (N_10054,N_9802,N_9908);
xnor U10055 (N_10055,N_9851,N_9904);
and U10056 (N_10056,N_9895,N_9965);
and U10057 (N_10057,N_9920,N_9863);
xor U10058 (N_10058,N_9837,N_9989);
nand U10059 (N_10059,N_9914,N_9950);
nand U10060 (N_10060,N_9856,N_9973);
and U10061 (N_10061,N_9943,N_9902);
nor U10062 (N_10062,N_9846,N_9924);
or U10063 (N_10063,N_9814,N_9805);
xnor U10064 (N_10064,N_9993,N_9848);
and U10065 (N_10065,N_9882,N_9928);
xor U10066 (N_10066,N_9921,N_9997);
xnor U10067 (N_10067,N_9833,N_9949);
and U10068 (N_10068,N_9978,N_9800);
or U10069 (N_10069,N_9807,N_9981);
nor U10070 (N_10070,N_9812,N_9951);
and U10071 (N_10071,N_9809,N_9964);
or U10072 (N_10072,N_9831,N_9884);
nor U10073 (N_10073,N_9932,N_9828);
nand U10074 (N_10074,N_9823,N_9876);
xor U10075 (N_10075,N_9822,N_9931);
or U10076 (N_10076,N_9990,N_9953);
xor U10077 (N_10077,N_9952,N_9894);
nand U10078 (N_10078,N_9979,N_9985);
or U10079 (N_10079,N_9994,N_9872);
and U10080 (N_10080,N_9905,N_9854);
nand U10081 (N_10081,N_9946,N_9858);
nor U10082 (N_10082,N_9995,N_9955);
and U10083 (N_10083,N_9824,N_9888);
xnor U10084 (N_10084,N_9804,N_9861);
and U10085 (N_10085,N_9909,N_9970);
nand U10086 (N_10086,N_9956,N_9825);
or U10087 (N_10087,N_9862,N_9849);
nand U10088 (N_10088,N_9816,N_9934);
and U10089 (N_10089,N_9996,N_9957);
nand U10090 (N_10090,N_9907,N_9868);
xnor U10091 (N_10091,N_9915,N_9881);
nor U10092 (N_10092,N_9947,N_9857);
xor U10093 (N_10093,N_9886,N_9903);
nor U10094 (N_10094,N_9870,N_9926);
nand U10095 (N_10095,N_9960,N_9918);
or U10096 (N_10096,N_9839,N_9917);
xnor U10097 (N_10097,N_9880,N_9879);
nand U10098 (N_10098,N_9987,N_9910);
nor U10099 (N_10099,N_9866,N_9959);
and U10100 (N_10100,N_9980,N_9977);
nand U10101 (N_10101,N_9892,N_9997);
or U10102 (N_10102,N_9926,N_9952);
xor U10103 (N_10103,N_9851,N_9894);
xnor U10104 (N_10104,N_9888,N_9977);
or U10105 (N_10105,N_9918,N_9841);
xnor U10106 (N_10106,N_9942,N_9886);
nor U10107 (N_10107,N_9911,N_9852);
xnor U10108 (N_10108,N_9937,N_9967);
xnor U10109 (N_10109,N_9986,N_9889);
nand U10110 (N_10110,N_9973,N_9999);
or U10111 (N_10111,N_9962,N_9929);
nand U10112 (N_10112,N_9844,N_9962);
nor U10113 (N_10113,N_9935,N_9883);
or U10114 (N_10114,N_9998,N_9920);
or U10115 (N_10115,N_9957,N_9893);
or U10116 (N_10116,N_9830,N_9805);
nor U10117 (N_10117,N_9820,N_9952);
or U10118 (N_10118,N_9868,N_9891);
nor U10119 (N_10119,N_9878,N_9962);
nor U10120 (N_10120,N_9835,N_9847);
xnor U10121 (N_10121,N_9887,N_9885);
or U10122 (N_10122,N_9977,N_9820);
or U10123 (N_10123,N_9808,N_9822);
nor U10124 (N_10124,N_9929,N_9923);
xnor U10125 (N_10125,N_9999,N_9959);
xor U10126 (N_10126,N_9908,N_9954);
or U10127 (N_10127,N_9985,N_9883);
xnor U10128 (N_10128,N_9872,N_9926);
nand U10129 (N_10129,N_9872,N_9945);
xor U10130 (N_10130,N_9974,N_9955);
xnor U10131 (N_10131,N_9848,N_9992);
or U10132 (N_10132,N_9816,N_9826);
or U10133 (N_10133,N_9832,N_9866);
nor U10134 (N_10134,N_9996,N_9832);
and U10135 (N_10135,N_9966,N_9952);
and U10136 (N_10136,N_9884,N_9809);
or U10137 (N_10137,N_9817,N_9881);
and U10138 (N_10138,N_9868,N_9997);
and U10139 (N_10139,N_9825,N_9952);
nor U10140 (N_10140,N_9999,N_9921);
xor U10141 (N_10141,N_9822,N_9813);
nor U10142 (N_10142,N_9982,N_9806);
xor U10143 (N_10143,N_9800,N_9859);
xnor U10144 (N_10144,N_9820,N_9813);
xnor U10145 (N_10145,N_9883,N_9940);
nor U10146 (N_10146,N_9999,N_9956);
or U10147 (N_10147,N_9983,N_9921);
nor U10148 (N_10148,N_9921,N_9891);
or U10149 (N_10149,N_9922,N_9961);
nor U10150 (N_10150,N_9880,N_9894);
or U10151 (N_10151,N_9971,N_9912);
and U10152 (N_10152,N_9915,N_9953);
or U10153 (N_10153,N_9960,N_9822);
and U10154 (N_10154,N_9941,N_9980);
xnor U10155 (N_10155,N_9838,N_9943);
nor U10156 (N_10156,N_9813,N_9966);
xor U10157 (N_10157,N_9914,N_9837);
and U10158 (N_10158,N_9874,N_9962);
nand U10159 (N_10159,N_9908,N_9838);
xor U10160 (N_10160,N_9861,N_9824);
nor U10161 (N_10161,N_9971,N_9823);
nor U10162 (N_10162,N_9914,N_9921);
or U10163 (N_10163,N_9894,N_9954);
nor U10164 (N_10164,N_9881,N_9861);
xnor U10165 (N_10165,N_9805,N_9838);
and U10166 (N_10166,N_9810,N_9882);
and U10167 (N_10167,N_9928,N_9913);
nand U10168 (N_10168,N_9827,N_9807);
nand U10169 (N_10169,N_9820,N_9812);
xor U10170 (N_10170,N_9954,N_9929);
or U10171 (N_10171,N_9988,N_9998);
xnor U10172 (N_10172,N_9881,N_9866);
nor U10173 (N_10173,N_9998,N_9839);
xor U10174 (N_10174,N_9872,N_9895);
nand U10175 (N_10175,N_9871,N_9960);
nand U10176 (N_10176,N_9875,N_9802);
and U10177 (N_10177,N_9839,N_9959);
xor U10178 (N_10178,N_9866,N_9885);
and U10179 (N_10179,N_9840,N_9864);
and U10180 (N_10180,N_9885,N_9808);
and U10181 (N_10181,N_9809,N_9914);
nor U10182 (N_10182,N_9826,N_9829);
nor U10183 (N_10183,N_9838,N_9892);
or U10184 (N_10184,N_9905,N_9988);
nand U10185 (N_10185,N_9978,N_9839);
nor U10186 (N_10186,N_9945,N_9899);
and U10187 (N_10187,N_9858,N_9963);
xor U10188 (N_10188,N_9898,N_9946);
xor U10189 (N_10189,N_9960,N_9846);
nor U10190 (N_10190,N_9871,N_9992);
or U10191 (N_10191,N_9821,N_9987);
nor U10192 (N_10192,N_9905,N_9855);
and U10193 (N_10193,N_9911,N_9805);
nor U10194 (N_10194,N_9908,N_9988);
or U10195 (N_10195,N_9944,N_9890);
and U10196 (N_10196,N_9818,N_9819);
xor U10197 (N_10197,N_9934,N_9901);
nand U10198 (N_10198,N_9924,N_9949);
and U10199 (N_10199,N_9860,N_9877);
and U10200 (N_10200,N_10089,N_10171);
and U10201 (N_10201,N_10076,N_10094);
nand U10202 (N_10202,N_10038,N_10197);
nor U10203 (N_10203,N_10077,N_10196);
nor U10204 (N_10204,N_10121,N_10090);
nand U10205 (N_10205,N_10006,N_10075);
xor U10206 (N_10206,N_10116,N_10149);
nand U10207 (N_10207,N_10156,N_10024);
or U10208 (N_10208,N_10135,N_10029);
nand U10209 (N_10209,N_10047,N_10065);
and U10210 (N_10210,N_10097,N_10161);
or U10211 (N_10211,N_10180,N_10034);
nor U10212 (N_10212,N_10157,N_10187);
nand U10213 (N_10213,N_10058,N_10183);
or U10214 (N_10214,N_10199,N_10099);
and U10215 (N_10215,N_10134,N_10186);
and U10216 (N_10216,N_10142,N_10013);
nand U10217 (N_10217,N_10009,N_10128);
and U10218 (N_10218,N_10125,N_10012);
nand U10219 (N_10219,N_10062,N_10092);
nor U10220 (N_10220,N_10074,N_10095);
nor U10221 (N_10221,N_10035,N_10046);
and U10222 (N_10222,N_10179,N_10093);
nor U10223 (N_10223,N_10030,N_10194);
nor U10224 (N_10224,N_10081,N_10131);
nor U10225 (N_10225,N_10079,N_10020);
nand U10226 (N_10226,N_10073,N_10049);
or U10227 (N_10227,N_10140,N_10100);
nor U10228 (N_10228,N_10043,N_10101);
xnor U10229 (N_10229,N_10039,N_10174);
and U10230 (N_10230,N_10045,N_10160);
nand U10231 (N_10231,N_10167,N_10106);
nand U10232 (N_10232,N_10069,N_10071);
or U10233 (N_10233,N_10138,N_10153);
nand U10234 (N_10234,N_10011,N_10178);
xnor U10235 (N_10235,N_10133,N_10064);
nand U10236 (N_10236,N_10072,N_10017);
and U10237 (N_10237,N_10170,N_10123);
and U10238 (N_10238,N_10185,N_10127);
and U10239 (N_10239,N_10091,N_10117);
or U10240 (N_10240,N_10018,N_10023);
xnor U10241 (N_10241,N_10086,N_10056);
nor U10242 (N_10242,N_10118,N_10036);
nand U10243 (N_10243,N_10147,N_10145);
nand U10244 (N_10244,N_10002,N_10155);
and U10245 (N_10245,N_10028,N_10141);
xnor U10246 (N_10246,N_10007,N_10022);
nor U10247 (N_10247,N_10126,N_10082);
xnor U10248 (N_10248,N_10098,N_10190);
and U10249 (N_10249,N_10198,N_10003);
nand U10250 (N_10250,N_10087,N_10120);
nor U10251 (N_10251,N_10025,N_10109);
nor U10252 (N_10252,N_10041,N_10172);
xnor U10253 (N_10253,N_10026,N_10068);
nand U10254 (N_10254,N_10195,N_10188);
nand U10255 (N_10255,N_10139,N_10189);
nand U10256 (N_10256,N_10061,N_10132);
nor U10257 (N_10257,N_10021,N_10163);
nand U10258 (N_10258,N_10129,N_10137);
nand U10259 (N_10259,N_10184,N_10169);
and U10260 (N_10260,N_10150,N_10067);
xor U10261 (N_10261,N_10143,N_10103);
nand U10262 (N_10262,N_10173,N_10080);
and U10263 (N_10263,N_10044,N_10158);
or U10264 (N_10264,N_10085,N_10000);
xnor U10265 (N_10265,N_10037,N_10001);
nor U10266 (N_10266,N_10159,N_10083);
or U10267 (N_10267,N_10164,N_10193);
nor U10268 (N_10268,N_10078,N_10004);
or U10269 (N_10269,N_10005,N_10027);
nand U10270 (N_10270,N_10019,N_10048);
or U10271 (N_10271,N_10032,N_10059);
or U10272 (N_10272,N_10177,N_10010);
nand U10273 (N_10273,N_10119,N_10136);
or U10274 (N_10274,N_10114,N_10084);
nand U10275 (N_10275,N_10040,N_10107);
nor U10276 (N_10276,N_10096,N_10181);
or U10277 (N_10277,N_10112,N_10088);
xnor U10278 (N_10278,N_10122,N_10033);
nor U10279 (N_10279,N_10104,N_10057);
xnor U10280 (N_10280,N_10111,N_10053);
xnor U10281 (N_10281,N_10031,N_10113);
and U10282 (N_10282,N_10175,N_10130);
nor U10283 (N_10283,N_10063,N_10148);
xnor U10284 (N_10284,N_10008,N_10192);
nor U10285 (N_10285,N_10108,N_10105);
xnor U10286 (N_10286,N_10146,N_10066);
or U10287 (N_10287,N_10102,N_10042);
nor U10288 (N_10288,N_10014,N_10110);
xnor U10289 (N_10289,N_10154,N_10151);
nand U10290 (N_10290,N_10144,N_10052);
xor U10291 (N_10291,N_10055,N_10176);
xor U10292 (N_10292,N_10162,N_10060);
or U10293 (N_10293,N_10124,N_10166);
and U10294 (N_10294,N_10050,N_10070);
xor U10295 (N_10295,N_10165,N_10152);
xnor U10296 (N_10296,N_10054,N_10182);
and U10297 (N_10297,N_10191,N_10051);
xnor U10298 (N_10298,N_10115,N_10016);
nor U10299 (N_10299,N_10168,N_10015);
xor U10300 (N_10300,N_10149,N_10136);
and U10301 (N_10301,N_10144,N_10195);
or U10302 (N_10302,N_10100,N_10177);
and U10303 (N_10303,N_10180,N_10058);
xnor U10304 (N_10304,N_10162,N_10132);
nand U10305 (N_10305,N_10067,N_10077);
nand U10306 (N_10306,N_10008,N_10049);
xnor U10307 (N_10307,N_10124,N_10096);
or U10308 (N_10308,N_10057,N_10127);
nor U10309 (N_10309,N_10049,N_10136);
and U10310 (N_10310,N_10006,N_10004);
xnor U10311 (N_10311,N_10091,N_10145);
nand U10312 (N_10312,N_10157,N_10158);
nand U10313 (N_10313,N_10096,N_10179);
or U10314 (N_10314,N_10026,N_10032);
nor U10315 (N_10315,N_10002,N_10007);
nand U10316 (N_10316,N_10062,N_10028);
and U10317 (N_10317,N_10011,N_10012);
xor U10318 (N_10318,N_10179,N_10095);
or U10319 (N_10319,N_10147,N_10072);
nand U10320 (N_10320,N_10083,N_10111);
and U10321 (N_10321,N_10005,N_10009);
and U10322 (N_10322,N_10061,N_10018);
xor U10323 (N_10323,N_10140,N_10067);
nand U10324 (N_10324,N_10085,N_10166);
nand U10325 (N_10325,N_10025,N_10018);
nand U10326 (N_10326,N_10098,N_10131);
nor U10327 (N_10327,N_10115,N_10053);
nor U10328 (N_10328,N_10107,N_10089);
nor U10329 (N_10329,N_10154,N_10104);
xnor U10330 (N_10330,N_10041,N_10057);
or U10331 (N_10331,N_10140,N_10053);
xor U10332 (N_10332,N_10042,N_10059);
and U10333 (N_10333,N_10047,N_10067);
and U10334 (N_10334,N_10158,N_10183);
nand U10335 (N_10335,N_10028,N_10157);
nor U10336 (N_10336,N_10156,N_10107);
or U10337 (N_10337,N_10071,N_10018);
nor U10338 (N_10338,N_10027,N_10051);
xnor U10339 (N_10339,N_10086,N_10179);
and U10340 (N_10340,N_10121,N_10136);
xnor U10341 (N_10341,N_10154,N_10100);
xnor U10342 (N_10342,N_10058,N_10157);
or U10343 (N_10343,N_10104,N_10011);
nand U10344 (N_10344,N_10113,N_10105);
and U10345 (N_10345,N_10096,N_10156);
and U10346 (N_10346,N_10136,N_10126);
xnor U10347 (N_10347,N_10094,N_10167);
xnor U10348 (N_10348,N_10072,N_10139);
nand U10349 (N_10349,N_10043,N_10026);
xnor U10350 (N_10350,N_10142,N_10186);
and U10351 (N_10351,N_10079,N_10192);
xor U10352 (N_10352,N_10013,N_10107);
nand U10353 (N_10353,N_10006,N_10033);
nor U10354 (N_10354,N_10054,N_10149);
and U10355 (N_10355,N_10097,N_10181);
nor U10356 (N_10356,N_10036,N_10054);
xnor U10357 (N_10357,N_10147,N_10192);
nand U10358 (N_10358,N_10046,N_10063);
or U10359 (N_10359,N_10121,N_10100);
nor U10360 (N_10360,N_10179,N_10078);
xor U10361 (N_10361,N_10098,N_10078);
and U10362 (N_10362,N_10108,N_10136);
and U10363 (N_10363,N_10043,N_10111);
and U10364 (N_10364,N_10028,N_10049);
xor U10365 (N_10365,N_10133,N_10034);
nand U10366 (N_10366,N_10087,N_10022);
nand U10367 (N_10367,N_10086,N_10016);
nor U10368 (N_10368,N_10145,N_10003);
or U10369 (N_10369,N_10120,N_10114);
nand U10370 (N_10370,N_10024,N_10074);
nor U10371 (N_10371,N_10053,N_10052);
nand U10372 (N_10372,N_10161,N_10080);
or U10373 (N_10373,N_10112,N_10013);
or U10374 (N_10374,N_10156,N_10078);
nand U10375 (N_10375,N_10096,N_10178);
xnor U10376 (N_10376,N_10040,N_10101);
xor U10377 (N_10377,N_10195,N_10164);
or U10378 (N_10378,N_10116,N_10156);
nor U10379 (N_10379,N_10050,N_10084);
or U10380 (N_10380,N_10027,N_10041);
nor U10381 (N_10381,N_10055,N_10097);
nor U10382 (N_10382,N_10183,N_10020);
or U10383 (N_10383,N_10004,N_10170);
and U10384 (N_10384,N_10128,N_10147);
or U10385 (N_10385,N_10130,N_10153);
nand U10386 (N_10386,N_10041,N_10121);
or U10387 (N_10387,N_10153,N_10166);
nand U10388 (N_10388,N_10026,N_10191);
or U10389 (N_10389,N_10033,N_10005);
xnor U10390 (N_10390,N_10152,N_10094);
nand U10391 (N_10391,N_10055,N_10003);
or U10392 (N_10392,N_10166,N_10081);
xnor U10393 (N_10393,N_10046,N_10079);
and U10394 (N_10394,N_10146,N_10084);
and U10395 (N_10395,N_10154,N_10159);
nor U10396 (N_10396,N_10150,N_10132);
or U10397 (N_10397,N_10193,N_10014);
nor U10398 (N_10398,N_10116,N_10153);
xnor U10399 (N_10399,N_10192,N_10129);
nand U10400 (N_10400,N_10312,N_10350);
nor U10401 (N_10401,N_10200,N_10275);
and U10402 (N_10402,N_10342,N_10250);
nor U10403 (N_10403,N_10314,N_10245);
nor U10404 (N_10404,N_10257,N_10234);
and U10405 (N_10405,N_10352,N_10349);
or U10406 (N_10406,N_10203,N_10371);
nor U10407 (N_10407,N_10308,N_10344);
nor U10408 (N_10408,N_10309,N_10322);
nor U10409 (N_10409,N_10380,N_10387);
or U10410 (N_10410,N_10272,N_10399);
nor U10411 (N_10411,N_10252,N_10357);
xnor U10412 (N_10412,N_10355,N_10227);
and U10413 (N_10413,N_10249,N_10319);
and U10414 (N_10414,N_10226,N_10341);
nand U10415 (N_10415,N_10222,N_10392);
and U10416 (N_10416,N_10379,N_10369);
nor U10417 (N_10417,N_10280,N_10232);
nand U10418 (N_10418,N_10265,N_10367);
and U10419 (N_10419,N_10286,N_10266);
or U10420 (N_10420,N_10273,N_10316);
or U10421 (N_10421,N_10331,N_10239);
nand U10422 (N_10422,N_10213,N_10261);
xnor U10423 (N_10423,N_10324,N_10201);
xnor U10424 (N_10424,N_10231,N_10304);
nand U10425 (N_10425,N_10277,N_10386);
and U10426 (N_10426,N_10323,N_10356);
nor U10427 (N_10427,N_10313,N_10298);
or U10428 (N_10428,N_10335,N_10268);
nor U10429 (N_10429,N_10393,N_10364);
nor U10430 (N_10430,N_10247,N_10333);
nand U10431 (N_10431,N_10358,N_10376);
nor U10432 (N_10432,N_10220,N_10372);
xnor U10433 (N_10433,N_10398,N_10296);
xnor U10434 (N_10434,N_10353,N_10307);
nand U10435 (N_10435,N_10329,N_10242);
and U10436 (N_10436,N_10260,N_10334);
or U10437 (N_10437,N_10291,N_10288);
and U10438 (N_10438,N_10271,N_10365);
nand U10439 (N_10439,N_10290,N_10303);
or U10440 (N_10440,N_10240,N_10327);
or U10441 (N_10441,N_10306,N_10388);
nor U10442 (N_10442,N_10326,N_10297);
nand U10443 (N_10443,N_10264,N_10255);
and U10444 (N_10444,N_10321,N_10359);
nand U10445 (N_10445,N_10243,N_10208);
nor U10446 (N_10446,N_10241,N_10237);
nor U10447 (N_10447,N_10218,N_10345);
or U10448 (N_10448,N_10251,N_10395);
nor U10449 (N_10449,N_10246,N_10362);
nand U10450 (N_10450,N_10391,N_10211);
xnor U10451 (N_10451,N_10295,N_10366);
and U10452 (N_10452,N_10228,N_10315);
or U10453 (N_10453,N_10206,N_10368);
and U10454 (N_10454,N_10215,N_10336);
xor U10455 (N_10455,N_10385,N_10305);
xnor U10456 (N_10456,N_10236,N_10343);
xor U10457 (N_10457,N_10262,N_10374);
and U10458 (N_10458,N_10209,N_10301);
and U10459 (N_10459,N_10210,N_10259);
or U10460 (N_10460,N_10382,N_10363);
and U10461 (N_10461,N_10383,N_10394);
nor U10462 (N_10462,N_10270,N_10235);
nor U10463 (N_10463,N_10373,N_10225);
or U10464 (N_10464,N_10337,N_10354);
nor U10465 (N_10465,N_10258,N_10294);
or U10466 (N_10466,N_10238,N_10302);
nor U10467 (N_10467,N_10282,N_10330);
and U10468 (N_10468,N_10311,N_10332);
nand U10469 (N_10469,N_10348,N_10339);
and U10470 (N_10470,N_10390,N_10299);
xnor U10471 (N_10471,N_10292,N_10397);
nand U10472 (N_10472,N_10338,N_10293);
nor U10473 (N_10473,N_10221,N_10328);
and U10474 (N_10474,N_10375,N_10205);
nor U10475 (N_10475,N_10285,N_10253);
nand U10476 (N_10476,N_10219,N_10360);
or U10477 (N_10477,N_10233,N_10325);
and U10478 (N_10478,N_10204,N_10310);
or U10479 (N_10479,N_10283,N_10351);
nor U10480 (N_10480,N_10279,N_10384);
nand U10481 (N_10481,N_10256,N_10212);
nor U10482 (N_10482,N_10244,N_10281);
nor U10483 (N_10483,N_10389,N_10317);
nand U10484 (N_10484,N_10202,N_10248);
nor U10485 (N_10485,N_10320,N_10230);
nor U10486 (N_10486,N_10378,N_10267);
or U10487 (N_10487,N_10214,N_10318);
nor U10488 (N_10488,N_10223,N_10347);
nor U10489 (N_10489,N_10229,N_10254);
or U10490 (N_10490,N_10377,N_10396);
nand U10491 (N_10491,N_10263,N_10381);
xor U10492 (N_10492,N_10300,N_10276);
and U10493 (N_10493,N_10278,N_10274);
or U10494 (N_10494,N_10340,N_10224);
nand U10495 (N_10495,N_10370,N_10284);
and U10496 (N_10496,N_10269,N_10289);
or U10497 (N_10497,N_10346,N_10207);
nand U10498 (N_10498,N_10217,N_10216);
or U10499 (N_10499,N_10361,N_10287);
xnor U10500 (N_10500,N_10269,N_10222);
and U10501 (N_10501,N_10304,N_10320);
nand U10502 (N_10502,N_10379,N_10224);
or U10503 (N_10503,N_10258,N_10253);
nor U10504 (N_10504,N_10222,N_10264);
or U10505 (N_10505,N_10290,N_10355);
nand U10506 (N_10506,N_10222,N_10258);
or U10507 (N_10507,N_10308,N_10289);
xnor U10508 (N_10508,N_10251,N_10235);
nand U10509 (N_10509,N_10209,N_10216);
and U10510 (N_10510,N_10320,N_10376);
or U10511 (N_10511,N_10243,N_10371);
xnor U10512 (N_10512,N_10243,N_10232);
xnor U10513 (N_10513,N_10211,N_10382);
or U10514 (N_10514,N_10271,N_10234);
or U10515 (N_10515,N_10355,N_10288);
or U10516 (N_10516,N_10294,N_10352);
or U10517 (N_10517,N_10344,N_10323);
or U10518 (N_10518,N_10243,N_10253);
nor U10519 (N_10519,N_10313,N_10231);
nor U10520 (N_10520,N_10200,N_10264);
nand U10521 (N_10521,N_10207,N_10276);
xor U10522 (N_10522,N_10299,N_10382);
and U10523 (N_10523,N_10397,N_10216);
nand U10524 (N_10524,N_10308,N_10205);
nand U10525 (N_10525,N_10283,N_10294);
nand U10526 (N_10526,N_10378,N_10276);
xor U10527 (N_10527,N_10347,N_10206);
nor U10528 (N_10528,N_10289,N_10332);
and U10529 (N_10529,N_10296,N_10269);
or U10530 (N_10530,N_10345,N_10343);
xor U10531 (N_10531,N_10252,N_10325);
and U10532 (N_10532,N_10328,N_10261);
and U10533 (N_10533,N_10252,N_10244);
nor U10534 (N_10534,N_10302,N_10231);
and U10535 (N_10535,N_10282,N_10249);
nor U10536 (N_10536,N_10291,N_10365);
or U10537 (N_10537,N_10263,N_10369);
xor U10538 (N_10538,N_10296,N_10200);
nor U10539 (N_10539,N_10273,N_10302);
nand U10540 (N_10540,N_10306,N_10322);
or U10541 (N_10541,N_10319,N_10323);
nand U10542 (N_10542,N_10294,N_10217);
nor U10543 (N_10543,N_10246,N_10327);
and U10544 (N_10544,N_10351,N_10235);
or U10545 (N_10545,N_10349,N_10291);
or U10546 (N_10546,N_10209,N_10383);
xnor U10547 (N_10547,N_10275,N_10311);
xor U10548 (N_10548,N_10217,N_10319);
nor U10549 (N_10549,N_10252,N_10344);
xnor U10550 (N_10550,N_10283,N_10378);
xnor U10551 (N_10551,N_10386,N_10243);
or U10552 (N_10552,N_10342,N_10312);
nand U10553 (N_10553,N_10287,N_10224);
nor U10554 (N_10554,N_10291,N_10242);
or U10555 (N_10555,N_10327,N_10259);
nand U10556 (N_10556,N_10244,N_10285);
nor U10557 (N_10557,N_10314,N_10272);
nand U10558 (N_10558,N_10237,N_10390);
or U10559 (N_10559,N_10331,N_10390);
or U10560 (N_10560,N_10239,N_10309);
and U10561 (N_10561,N_10343,N_10309);
or U10562 (N_10562,N_10269,N_10355);
and U10563 (N_10563,N_10289,N_10328);
nand U10564 (N_10564,N_10373,N_10393);
nor U10565 (N_10565,N_10218,N_10395);
and U10566 (N_10566,N_10223,N_10227);
nor U10567 (N_10567,N_10349,N_10276);
nor U10568 (N_10568,N_10306,N_10224);
or U10569 (N_10569,N_10226,N_10239);
or U10570 (N_10570,N_10368,N_10217);
nand U10571 (N_10571,N_10334,N_10218);
or U10572 (N_10572,N_10241,N_10332);
or U10573 (N_10573,N_10267,N_10288);
and U10574 (N_10574,N_10324,N_10316);
xor U10575 (N_10575,N_10394,N_10287);
xor U10576 (N_10576,N_10244,N_10335);
nor U10577 (N_10577,N_10350,N_10275);
xor U10578 (N_10578,N_10336,N_10333);
or U10579 (N_10579,N_10306,N_10246);
nand U10580 (N_10580,N_10330,N_10316);
or U10581 (N_10581,N_10336,N_10361);
nand U10582 (N_10582,N_10202,N_10398);
or U10583 (N_10583,N_10261,N_10324);
xnor U10584 (N_10584,N_10352,N_10282);
nand U10585 (N_10585,N_10392,N_10250);
nor U10586 (N_10586,N_10257,N_10200);
and U10587 (N_10587,N_10226,N_10244);
xnor U10588 (N_10588,N_10374,N_10254);
nand U10589 (N_10589,N_10367,N_10386);
xnor U10590 (N_10590,N_10390,N_10233);
or U10591 (N_10591,N_10333,N_10311);
nand U10592 (N_10592,N_10338,N_10353);
and U10593 (N_10593,N_10360,N_10378);
nand U10594 (N_10594,N_10343,N_10318);
xnor U10595 (N_10595,N_10334,N_10206);
xor U10596 (N_10596,N_10282,N_10229);
and U10597 (N_10597,N_10200,N_10355);
nor U10598 (N_10598,N_10239,N_10351);
xor U10599 (N_10599,N_10301,N_10311);
nor U10600 (N_10600,N_10597,N_10406);
nand U10601 (N_10601,N_10500,N_10538);
xor U10602 (N_10602,N_10579,N_10498);
nand U10603 (N_10603,N_10527,N_10595);
xor U10604 (N_10604,N_10514,N_10484);
nand U10605 (N_10605,N_10561,N_10466);
and U10606 (N_10606,N_10513,N_10435);
nand U10607 (N_10607,N_10508,N_10430);
nor U10608 (N_10608,N_10476,N_10452);
and U10609 (N_10609,N_10402,N_10460);
nor U10610 (N_10610,N_10502,N_10481);
and U10611 (N_10611,N_10506,N_10469);
or U10612 (N_10612,N_10511,N_10468);
xnor U10613 (N_10613,N_10467,N_10571);
xnor U10614 (N_10614,N_10586,N_10507);
nand U10615 (N_10615,N_10545,N_10457);
or U10616 (N_10616,N_10491,N_10518);
or U10617 (N_10617,N_10437,N_10458);
xnor U10618 (N_10618,N_10431,N_10563);
xor U10619 (N_10619,N_10499,N_10540);
xor U10620 (N_10620,N_10543,N_10525);
or U10621 (N_10621,N_10400,N_10429);
or U10622 (N_10622,N_10464,N_10570);
and U10623 (N_10623,N_10454,N_10456);
xor U10624 (N_10624,N_10510,N_10578);
nor U10625 (N_10625,N_10477,N_10504);
and U10626 (N_10626,N_10584,N_10472);
xor U10627 (N_10627,N_10544,N_10580);
nor U10628 (N_10628,N_10588,N_10433);
nor U10629 (N_10629,N_10416,N_10492);
nor U10630 (N_10630,N_10564,N_10451);
and U10631 (N_10631,N_10573,N_10426);
and U10632 (N_10632,N_10488,N_10547);
or U10633 (N_10633,N_10479,N_10592);
nand U10634 (N_10634,N_10443,N_10432);
or U10635 (N_10635,N_10568,N_10418);
xor U10636 (N_10636,N_10408,N_10449);
nor U10637 (N_10637,N_10576,N_10482);
or U10638 (N_10638,N_10594,N_10490);
nor U10639 (N_10639,N_10523,N_10422);
xnor U10640 (N_10640,N_10436,N_10559);
nand U10641 (N_10641,N_10448,N_10515);
and U10642 (N_10642,N_10516,N_10480);
xor U10643 (N_10643,N_10453,N_10483);
nor U10644 (N_10644,N_10572,N_10522);
and U10645 (N_10645,N_10503,N_10462);
nor U10646 (N_10646,N_10565,N_10412);
or U10647 (N_10647,N_10421,N_10419);
xnor U10648 (N_10648,N_10530,N_10444);
nor U10649 (N_10649,N_10420,N_10599);
nand U10650 (N_10650,N_10475,N_10495);
xnor U10651 (N_10651,N_10596,N_10591);
and U10652 (N_10652,N_10567,N_10427);
or U10653 (N_10653,N_10493,N_10486);
or U10654 (N_10654,N_10417,N_10471);
nand U10655 (N_10655,N_10566,N_10470);
xnor U10656 (N_10656,N_10541,N_10455);
nand U10657 (N_10657,N_10465,N_10546);
nor U10658 (N_10658,N_10562,N_10425);
nor U10659 (N_10659,N_10407,N_10519);
nor U10660 (N_10660,N_10528,N_10549);
or U10661 (N_10661,N_10521,N_10555);
nand U10662 (N_10662,N_10590,N_10526);
nor U10663 (N_10663,N_10478,N_10520);
and U10664 (N_10664,N_10405,N_10461);
nand U10665 (N_10665,N_10553,N_10410);
nor U10666 (N_10666,N_10560,N_10554);
nor U10667 (N_10667,N_10533,N_10445);
nor U10668 (N_10668,N_10575,N_10411);
nor U10669 (N_10669,N_10532,N_10574);
or U10670 (N_10670,N_10428,N_10473);
and U10671 (N_10671,N_10524,N_10593);
nand U10672 (N_10672,N_10534,N_10550);
nor U10673 (N_10673,N_10459,N_10434);
xnor U10674 (N_10674,N_10581,N_10577);
nand U10675 (N_10675,N_10404,N_10542);
and U10676 (N_10676,N_10531,N_10529);
nand U10677 (N_10677,N_10474,N_10557);
xor U10678 (N_10678,N_10558,N_10535);
nand U10679 (N_10679,N_10442,N_10413);
nand U10680 (N_10680,N_10536,N_10403);
or U10681 (N_10681,N_10441,N_10585);
and U10682 (N_10682,N_10497,N_10450);
xnor U10683 (N_10683,N_10414,N_10598);
and U10684 (N_10684,N_10496,N_10512);
nor U10685 (N_10685,N_10446,N_10487);
nand U10686 (N_10686,N_10505,N_10501);
nand U10687 (N_10687,N_10439,N_10582);
nand U10688 (N_10688,N_10583,N_10438);
and U10689 (N_10689,N_10548,N_10509);
nor U10690 (N_10690,N_10551,N_10539);
nor U10691 (N_10691,N_10517,N_10440);
and U10692 (N_10692,N_10552,N_10537);
nor U10693 (N_10693,N_10415,N_10485);
nor U10694 (N_10694,N_10447,N_10463);
or U10695 (N_10695,N_10424,N_10556);
nand U10696 (N_10696,N_10423,N_10494);
xor U10697 (N_10697,N_10409,N_10589);
and U10698 (N_10698,N_10587,N_10569);
or U10699 (N_10699,N_10489,N_10401);
xor U10700 (N_10700,N_10424,N_10416);
nand U10701 (N_10701,N_10599,N_10521);
xnor U10702 (N_10702,N_10564,N_10570);
or U10703 (N_10703,N_10437,N_10462);
nor U10704 (N_10704,N_10536,N_10563);
nor U10705 (N_10705,N_10483,N_10575);
and U10706 (N_10706,N_10568,N_10520);
and U10707 (N_10707,N_10443,N_10439);
nand U10708 (N_10708,N_10488,N_10448);
xor U10709 (N_10709,N_10437,N_10444);
nand U10710 (N_10710,N_10533,N_10597);
or U10711 (N_10711,N_10471,N_10556);
and U10712 (N_10712,N_10516,N_10494);
or U10713 (N_10713,N_10573,N_10507);
and U10714 (N_10714,N_10564,N_10590);
nor U10715 (N_10715,N_10536,N_10418);
nor U10716 (N_10716,N_10557,N_10526);
nor U10717 (N_10717,N_10405,N_10475);
nor U10718 (N_10718,N_10598,N_10552);
xnor U10719 (N_10719,N_10490,N_10402);
or U10720 (N_10720,N_10434,N_10427);
xor U10721 (N_10721,N_10552,N_10596);
or U10722 (N_10722,N_10577,N_10516);
xnor U10723 (N_10723,N_10519,N_10567);
and U10724 (N_10724,N_10480,N_10485);
xor U10725 (N_10725,N_10552,N_10479);
nand U10726 (N_10726,N_10580,N_10541);
or U10727 (N_10727,N_10485,N_10490);
nor U10728 (N_10728,N_10537,N_10421);
or U10729 (N_10729,N_10594,N_10576);
or U10730 (N_10730,N_10580,N_10584);
or U10731 (N_10731,N_10434,N_10527);
xor U10732 (N_10732,N_10535,N_10474);
and U10733 (N_10733,N_10453,N_10595);
nand U10734 (N_10734,N_10471,N_10408);
nand U10735 (N_10735,N_10575,N_10443);
and U10736 (N_10736,N_10422,N_10463);
nand U10737 (N_10737,N_10539,N_10553);
and U10738 (N_10738,N_10465,N_10432);
and U10739 (N_10739,N_10550,N_10584);
or U10740 (N_10740,N_10599,N_10430);
nor U10741 (N_10741,N_10485,N_10411);
and U10742 (N_10742,N_10497,N_10476);
and U10743 (N_10743,N_10425,N_10469);
nor U10744 (N_10744,N_10548,N_10431);
or U10745 (N_10745,N_10471,N_10494);
nor U10746 (N_10746,N_10413,N_10597);
and U10747 (N_10747,N_10441,N_10575);
or U10748 (N_10748,N_10518,N_10470);
nand U10749 (N_10749,N_10549,N_10576);
and U10750 (N_10750,N_10508,N_10488);
nor U10751 (N_10751,N_10512,N_10522);
and U10752 (N_10752,N_10597,N_10463);
or U10753 (N_10753,N_10542,N_10403);
nor U10754 (N_10754,N_10439,N_10427);
and U10755 (N_10755,N_10458,N_10472);
and U10756 (N_10756,N_10469,N_10536);
and U10757 (N_10757,N_10407,N_10414);
xor U10758 (N_10758,N_10519,N_10541);
nand U10759 (N_10759,N_10576,N_10567);
nand U10760 (N_10760,N_10590,N_10452);
or U10761 (N_10761,N_10497,N_10548);
or U10762 (N_10762,N_10418,N_10566);
xor U10763 (N_10763,N_10508,N_10477);
nor U10764 (N_10764,N_10540,N_10501);
nor U10765 (N_10765,N_10568,N_10426);
and U10766 (N_10766,N_10506,N_10453);
nand U10767 (N_10767,N_10554,N_10402);
or U10768 (N_10768,N_10578,N_10530);
xnor U10769 (N_10769,N_10463,N_10408);
or U10770 (N_10770,N_10434,N_10584);
or U10771 (N_10771,N_10572,N_10549);
nor U10772 (N_10772,N_10515,N_10537);
nor U10773 (N_10773,N_10472,N_10485);
xor U10774 (N_10774,N_10591,N_10428);
or U10775 (N_10775,N_10574,N_10503);
nor U10776 (N_10776,N_10538,N_10476);
nand U10777 (N_10777,N_10434,N_10543);
nor U10778 (N_10778,N_10521,N_10426);
nor U10779 (N_10779,N_10421,N_10556);
or U10780 (N_10780,N_10476,N_10419);
or U10781 (N_10781,N_10434,N_10426);
nand U10782 (N_10782,N_10435,N_10537);
or U10783 (N_10783,N_10487,N_10520);
xnor U10784 (N_10784,N_10473,N_10452);
nor U10785 (N_10785,N_10501,N_10537);
nand U10786 (N_10786,N_10428,N_10423);
nand U10787 (N_10787,N_10482,N_10557);
or U10788 (N_10788,N_10420,N_10436);
xor U10789 (N_10789,N_10592,N_10451);
xor U10790 (N_10790,N_10446,N_10527);
nor U10791 (N_10791,N_10409,N_10406);
nor U10792 (N_10792,N_10528,N_10570);
and U10793 (N_10793,N_10468,N_10525);
xor U10794 (N_10794,N_10431,N_10493);
xnor U10795 (N_10795,N_10460,N_10420);
nand U10796 (N_10796,N_10507,N_10474);
nand U10797 (N_10797,N_10481,N_10533);
and U10798 (N_10798,N_10561,N_10519);
or U10799 (N_10799,N_10441,N_10553);
or U10800 (N_10800,N_10694,N_10607);
nand U10801 (N_10801,N_10619,N_10782);
nor U10802 (N_10802,N_10676,N_10683);
and U10803 (N_10803,N_10747,N_10774);
or U10804 (N_10804,N_10618,N_10667);
nand U10805 (N_10805,N_10639,N_10692);
nor U10806 (N_10806,N_10605,N_10695);
nor U10807 (N_10807,N_10709,N_10753);
xnor U10808 (N_10808,N_10784,N_10648);
and U10809 (N_10809,N_10733,N_10778);
and U10810 (N_10810,N_10793,N_10609);
and U10811 (N_10811,N_10725,N_10620);
nor U10812 (N_10812,N_10760,N_10689);
or U10813 (N_10813,N_10650,N_10674);
and U10814 (N_10814,N_10697,N_10644);
nand U10815 (N_10815,N_10742,N_10714);
or U10816 (N_10816,N_10617,N_10748);
and U10817 (N_10817,N_10704,N_10628);
or U10818 (N_10818,N_10737,N_10655);
nor U10819 (N_10819,N_10729,N_10791);
xor U10820 (N_10820,N_10771,N_10625);
or U10821 (N_10821,N_10790,N_10608);
nand U10822 (N_10822,N_10719,N_10634);
and U10823 (N_10823,N_10796,N_10632);
nor U10824 (N_10824,N_10757,N_10746);
nand U10825 (N_10825,N_10705,N_10794);
or U10826 (N_10826,N_10602,N_10783);
xnor U10827 (N_10827,N_10651,N_10613);
nand U10828 (N_10828,N_10684,N_10682);
xor U10829 (N_10829,N_10726,N_10781);
and U10830 (N_10830,N_10600,N_10744);
xor U10831 (N_10831,N_10792,N_10763);
nand U10832 (N_10832,N_10691,N_10732);
xor U10833 (N_10833,N_10604,N_10711);
nand U10834 (N_10834,N_10706,N_10647);
nand U10835 (N_10835,N_10755,N_10713);
xnor U10836 (N_10836,N_10717,N_10675);
nand U10837 (N_10837,N_10730,N_10750);
or U10838 (N_10838,N_10669,N_10652);
or U10839 (N_10839,N_10621,N_10795);
nor U10840 (N_10840,N_10601,N_10788);
nor U10841 (N_10841,N_10645,N_10610);
nand U10842 (N_10842,N_10743,N_10649);
or U10843 (N_10843,N_10672,N_10657);
and U10844 (N_10844,N_10700,N_10777);
xnor U10845 (N_10845,N_10720,N_10681);
or U10846 (N_10846,N_10664,N_10615);
or U10847 (N_10847,N_10764,N_10715);
or U10848 (N_10848,N_10773,N_10679);
or U10849 (N_10849,N_10787,N_10756);
nand U10850 (N_10850,N_10626,N_10734);
nand U10851 (N_10851,N_10762,N_10780);
nor U10852 (N_10852,N_10623,N_10779);
nor U10853 (N_10853,N_10761,N_10660);
and U10854 (N_10854,N_10666,N_10712);
and U10855 (N_10855,N_10718,N_10749);
or U10856 (N_10856,N_10637,N_10786);
nor U10857 (N_10857,N_10641,N_10614);
xnor U10858 (N_10858,N_10668,N_10611);
nand U10859 (N_10859,N_10739,N_10693);
nand U10860 (N_10860,N_10708,N_10789);
or U10861 (N_10861,N_10622,N_10797);
xnor U10862 (N_10862,N_10710,N_10665);
and U10863 (N_10863,N_10653,N_10699);
xor U10864 (N_10864,N_10662,N_10661);
or U10865 (N_10865,N_10656,N_10735);
and U10866 (N_10866,N_10636,N_10659);
or U10867 (N_10867,N_10769,N_10736);
or U10868 (N_10868,N_10654,N_10798);
xor U10869 (N_10869,N_10670,N_10752);
and U10870 (N_10870,N_10646,N_10703);
xor U10871 (N_10871,N_10640,N_10616);
or U10872 (N_10872,N_10680,N_10728);
or U10873 (N_10873,N_10627,N_10698);
or U10874 (N_10874,N_10741,N_10673);
or U10875 (N_10875,N_10631,N_10612);
nor U10876 (N_10876,N_10606,N_10688);
xor U10877 (N_10877,N_10716,N_10766);
or U10878 (N_10878,N_10603,N_10635);
nor U10879 (N_10879,N_10642,N_10686);
nor U10880 (N_10880,N_10678,N_10702);
xnor U10881 (N_10881,N_10740,N_10775);
xnor U10882 (N_10882,N_10707,N_10751);
or U10883 (N_10883,N_10727,N_10745);
nor U10884 (N_10884,N_10690,N_10687);
xor U10885 (N_10885,N_10629,N_10677);
or U10886 (N_10886,N_10701,N_10767);
nor U10887 (N_10887,N_10721,N_10663);
nor U10888 (N_10888,N_10770,N_10696);
nor U10889 (N_10889,N_10799,N_10758);
nor U10890 (N_10890,N_10768,N_10624);
nor U10891 (N_10891,N_10638,N_10643);
xnor U10892 (N_10892,N_10685,N_10772);
or U10893 (N_10893,N_10724,N_10754);
nand U10894 (N_10894,N_10722,N_10633);
nor U10895 (N_10895,N_10765,N_10776);
xnor U10896 (N_10896,N_10630,N_10658);
nor U10897 (N_10897,N_10731,N_10671);
xor U10898 (N_10898,N_10738,N_10723);
nand U10899 (N_10899,N_10785,N_10759);
xnor U10900 (N_10900,N_10641,N_10611);
xnor U10901 (N_10901,N_10647,N_10681);
nor U10902 (N_10902,N_10782,N_10760);
and U10903 (N_10903,N_10726,N_10635);
nor U10904 (N_10904,N_10733,N_10643);
nor U10905 (N_10905,N_10719,N_10657);
nor U10906 (N_10906,N_10619,N_10689);
xor U10907 (N_10907,N_10782,N_10719);
xor U10908 (N_10908,N_10752,N_10626);
or U10909 (N_10909,N_10728,N_10606);
or U10910 (N_10910,N_10753,N_10747);
and U10911 (N_10911,N_10605,N_10600);
xor U10912 (N_10912,N_10794,N_10758);
and U10913 (N_10913,N_10630,N_10775);
nor U10914 (N_10914,N_10618,N_10669);
xnor U10915 (N_10915,N_10668,N_10692);
and U10916 (N_10916,N_10786,N_10734);
xnor U10917 (N_10917,N_10799,N_10603);
or U10918 (N_10918,N_10719,N_10766);
nand U10919 (N_10919,N_10750,N_10610);
nor U10920 (N_10920,N_10758,N_10774);
nor U10921 (N_10921,N_10684,N_10734);
nand U10922 (N_10922,N_10709,N_10665);
or U10923 (N_10923,N_10746,N_10661);
or U10924 (N_10924,N_10693,N_10697);
xor U10925 (N_10925,N_10738,N_10638);
and U10926 (N_10926,N_10737,N_10724);
nor U10927 (N_10927,N_10608,N_10723);
xnor U10928 (N_10928,N_10762,N_10759);
nand U10929 (N_10929,N_10649,N_10682);
xnor U10930 (N_10930,N_10748,N_10717);
nor U10931 (N_10931,N_10728,N_10699);
nand U10932 (N_10932,N_10721,N_10644);
nor U10933 (N_10933,N_10742,N_10658);
or U10934 (N_10934,N_10771,N_10727);
or U10935 (N_10935,N_10614,N_10676);
nand U10936 (N_10936,N_10683,N_10781);
xor U10937 (N_10937,N_10704,N_10764);
or U10938 (N_10938,N_10637,N_10741);
or U10939 (N_10939,N_10664,N_10793);
nor U10940 (N_10940,N_10746,N_10726);
and U10941 (N_10941,N_10658,N_10737);
nor U10942 (N_10942,N_10659,N_10603);
nor U10943 (N_10943,N_10663,N_10752);
and U10944 (N_10944,N_10753,N_10793);
nand U10945 (N_10945,N_10742,N_10648);
and U10946 (N_10946,N_10664,N_10653);
nor U10947 (N_10947,N_10772,N_10733);
xnor U10948 (N_10948,N_10787,N_10714);
or U10949 (N_10949,N_10633,N_10710);
nand U10950 (N_10950,N_10670,N_10609);
nand U10951 (N_10951,N_10643,N_10723);
nand U10952 (N_10952,N_10735,N_10797);
nand U10953 (N_10953,N_10677,N_10616);
nand U10954 (N_10954,N_10691,N_10726);
nand U10955 (N_10955,N_10750,N_10766);
xnor U10956 (N_10956,N_10737,N_10755);
xor U10957 (N_10957,N_10767,N_10721);
nor U10958 (N_10958,N_10633,N_10674);
and U10959 (N_10959,N_10660,N_10630);
xnor U10960 (N_10960,N_10672,N_10705);
or U10961 (N_10961,N_10660,N_10698);
nor U10962 (N_10962,N_10756,N_10648);
nor U10963 (N_10963,N_10788,N_10736);
nand U10964 (N_10964,N_10708,N_10668);
nand U10965 (N_10965,N_10736,N_10781);
xnor U10966 (N_10966,N_10711,N_10736);
and U10967 (N_10967,N_10773,N_10657);
and U10968 (N_10968,N_10649,N_10635);
nand U10969 (N_10969,N_10670,N_10707);
xnor U10970 (N_10970,N_10792,N_10677);
nand U10971 (N_10971,N_10728,N_10696);
xnor U10972 (N_10972,N_10767,N_10796);
nor U10973 (N_10973,N_10782,N_10746);
and U10974 (N_10974,N_10621,N_10788);
or U10975 (N_10975,N_10755,N_10602);
or U10976 (N_10976,N_10709,N_10776);
and U10977 (N_10977,N_10739,N_10683);
or U10978 (N_10978,N_10676,N_10607);
xor U10979 (N_10979,N_10772,N_10610);
nand U10980 (N_10980,N_10732,N_10728);
and U10981 (N_10981,N_10798,N_10751);
and U10982 (N_10982,N_10662,N_10766);
and U10983 (N_10983,N_10660,N_10785);
nand U10984 (N_10984,N_10786,N_10701);
and U10985 (N_10985,N_10602,N_10729);
or U10986 (N_10986,N_10649,N_10754);
or U10987 (N_10987,N_10751,N_10720);
or U10988 (N_10988,N_10629,N_10709);
and U10989 (N_10989,N_10750,N_10787);
nor U10990 (N_10990,N_10722,N_10788);
nor U10991 (N_10991,N_10778,N_10679);
nand U10992 (N_10992,N_10707,N_10687);
and U10993 (N_10993,N_10691,N_10760);
and U10994 (N_10994,N_10690,N_10774);
and U10995 (N_10995,N_10648,N_10770);
xor U10996 (N_10996,N_10617,N_10778);
nor U10997 (N_10997,N_10797,N_10730);
nor U10998 (N_10998,N_10793,N_10798);
nand U10999 (N_10999,N_10761,N_10756);
and U11000 (N_11000,N_10832,N_10883);
or U11001 (N_11001,N_10820,N_10941);
nand U11002 (N_11002,N_10942,N_10866);
nor U11003 (N_11003,N_10921,N_10914);
xor U11004 (N_11004,N_10873,N_10976);
xnor U11005 (N_11005,N_10838,N_10959);
nor U11006 (N_11006,N_10835,N_10897);
nand U11007 (N_11007,N_10855,N_10808);
xnor U11008 (N_11008,N_10990,N_10854);
nand U11009 (N_11009,N_10875,N_10915);
or U11010 (N_11010,N_10971,N_10804);
and U11011 (N_11011,N_10895,N_10884);
xor U11012 (N_11012,N_10890,N_10956);
nor U11013 (N_11013,N_10843,N_10944);
or U11014 (N_11014,N_10858,N_10824);
nand U11015 (N_11015,N_10978,N_10817);
and U11016 (N_11016,N_10874,N_10999);
nand U11017 (N_11017,N_10963,N_10821);
and U11018 (N_11018,N_10975,N_10943);
and U11019 (N_11019,N_10870,N_10907);
nand U11020 (N_11020,N_10932,N_10910);
xnor U11021 (N_11021,N_10871,N_10938);
and U11022 (N_11022,N_10853,N_10954);
or U11023 (N_11023,N_10836,N_10960);
nand U11024 (N_11024,N_10830,N_10969);
nand U11025 (N_11025,N_10998,N_10815);
nor U11026 (N_11026,N_10986,N_10894);
nand U11027 (N_11027,N_10893,N_10974);
or U11028 (N_11028,N_10923,N_10906);
nor U11029 (N_11029,N_10947,N_10805);
xor U11030 (N_11030,N_10810,N_10905);
or U11031 (N_11031,N_10869,N_10839);
xor U11032 (N_11032,N_10861,N_10888);
and U11033 (N_11033,N_10939,N_10864);
nor U11034 (N_11034,N_10967,N_10945);
xor U11035 (N_11035,N_10925,N_10826);
xor U11036 (N_11036,N_10879,N_10886);
nand U11037 (N_11037,N_10973,N_10878);
nand U11038 (N_11038,N_10952,N_10936);
and U11039 (N_11039,N_10991,N_10859);
xnor U11040 (N_11040,N_10989,N_10823);
xnor U11041 (N_11041,N_10857,N_10814);
or U11042 (N_11042,N_10995,N_10908);
nand U11043 (N_11043,N_10957,N_10982);
nand U11044 (N_11044,N_10926,N_10845);
and U11045 (N_11045,N_10802,N_10972);
nor U11046 (N_11046,N_10881,N_10951);
nor U11047 (N_11047,N_10961,N_10992);
xnor U11048 (N_11048,N_10968,N_10800);
xor U11049 (N_11049,N_10940,N_10807);
nand U11050 (N_11050,N_10924,N_10816);
and U11051 (N_11051,N_10948,N_10840);
xnor U11052 (N_11052,N_10933,N_10993);
nand U11053 (N_11053,N_10902,N_10977);
and U11054 (N_11054,N_10987,N_10920);
and U11055 (N_11055,N_10896,N_10867);
xor U11056 (N_11056,N_10980,N_10860);
xnor U11057 (N_11057,N_10806,N_10988);
nor U11058 (N_11058,N_10811,N_10842);
nor U11059 (N_11059,N_10825,N_10931);
nand U11060 (N_11060,N_10953,N_10928);
or U11061 (N_11061,N_10912,N_10970);
nand U11062 (N_11062,N_10898,N_10979);
or U11063 (N_11063,N_10872,N_10966);
xnor U11064 (N_11064,N_10801,N_10812);
nor U11065 (N_11065,N_10903,N_10929);
nand U11066 (N_11066,N_10851,N_10809);
and U11067 (N_11067,N_10965,N_10899);
xor U11068 (N_11068,N_10837,N_10891);
xor U11069 (N_11069,N_10919,N_10900);
or U11070 (N_11070,N_10834,N_10850);
nand U11071 (N_11071,N_10934,N_10937);
and U11072 (N_11072,N_10984,N_10913);
and U11073 (N_11073,N_10983,N_10964);
xnor U11074 (N_11074,N_10885,N_10849);
nand U11075 (N_11075,N_10955,N_10927);
and U11076 (N_11076,N_10862,N_10876);
xor U11077 (N_11077,N_10827,N_10997);
or U11078 (N_11078,N_10962,N_10841);
xnor U11079 (N_11079,N_10828,N_10877);
or U11080 (N_11080,N_10848,N_10844);
and U11081 (N_11081,N_10863,N_10918);
or U11082 (N_11082,N_10868,N_10803);
nor U11083 (N_11083,N_10901,N_10846);
nor U11084 (N_11084,N_10996,N_10958);
xnor U11085 (N_11085,N_10930,N_10813);
or U11086 (N_11086,N_10889,N_10831);
and U11087 (N_11087,N_10917,N_10946);
nor U11088 (N_11088,N_10909,N_10847);
nand U11089 (N_11089,N_10981,N_10892);
or U11090 (N_11090,N_10822,N_10865);
and U11091 (N_11091,N_10887,N_10904);
and U11092 (N_11092,N_10829,N_10985);
and U11093 (N_11093,N_10950,N_10949);
nor U11094 (N_11094,N_10833,N_10922);
nand U11095 (N_11095,N_10819,N_10880);
or U11096 (N_11096,N_10911,N_10818);
nor U11097 (N_11097,N_10935,N_10856);
nor U11098 (N_11098,N_10994,N_10916);
and U11099 (N_11099,N_10852,N_10882);
nor U11100 (N_11100,N_10995,N_10975);
nor U11101 (N_11101,N_10899,N_10858);
nor U11102 (N_11102,N_10837,N_10863);
and U11103 (N_11103,N_10919,N_10806);
or U11104 (N_11104,N_10943,N_10997);
nor U11105 (N_11105,N_10972,N_10981);
xor U11106 (N_11106,N_10905,N_10880);
nand U11107 (N_11107,N_10942,N_10973);
nor U11108 (N_11108,N_10859,N_10961);
nor U11109 (N_11109,N_10961,N_10907);
nor U11110 (N_11110,N_10910,N_10891);
xor U11111 (N_11111,N_10940,N_10975);
or U11112 (N_11112,N_10807,N_10816);
xor U11113 (N_11113,N_10873,N_10933);
and U11114 (N_11114,N_10800,N_10955);
and U11115 (N_11115,N_10876,N_10946);
xnor U11116 (N_11116,N_10821,N_10830);
xor U11117 (N_11117,N_10826,N_10997);
or U11118 (N_11118,N_10895,N_10914);
and U11119 (N_11119,N_10995,N_10956);
or U11120 (N_11120,N_10963,N_10985);
and U11121 (N_11121,N_10841,N_10955);
or U11122 (N_11122,N_10888,N_10982);
and U11123 (N_11123,N_10811,N_10859);
nor U11124 (N_11124,N_10908,N_10913);
xnor U11125 (N_11125,N_10904,N_10946);
or U11126 (N_11126,N_10988,N_10926);
and U11127 (N_11127,N_10908,N_10963);
nand U11128 (N_11128,N_10994,N_10933);
and U11129 (N_11129,N_10816,N_10984);
and U11130 (N_11130,N_10915,N_10872);
and U11131 (N_11131,N_10952,N_10804);
nand U11132 (N_11132,N_10932,N_10820);
or U11133 (N_11133,N_10983,N_10846);
nor U11134 (N_11134,N_10919,N_10824);
nand U11135 (N_11135,N_10996,N_10997);
and U11136 (N_11136,N_10825,N_10859);
nor U11137 (N_11137,N_10977,N_10937);
and U11138 (N_11138,N_10897,N_10997);
or U11139 (N_11139,N_10896,N_10802);
or U11140 (N_11140,N_10824,N_10820);
xor U11141 (N_11141,N_10908,N_10915);
nor U11142 (N_11142,N_10815,N_10979);
nor U11143 (N_11143,N_10909,N_10947);
nand U11144 (N_11144,N_10951,N_10927);
xnor U11145 (N_11145,N_10881,N_10930);
nor U11146 (N_11146,N_10931,N_10910);
xnor U11147 (N_11147,N_10946,N_10952);
xnor U11148 (N_11148,N_10950,N_10915);
xor U11149 (N_11149,N_10979,N_10916);
xnor U11150 (N_11150,N_10895,N_10926);
nor U11151 (N_11151,N_10864,N_10861);
and U11152 (N_11152,N_10952,N_10817);
and U11153 (N_11153,N_10806,N_10931);
nand U11154 (N_11154,N_10862,N_10975);
nand U11155 (N_11155,N_10848,N_10900);
xnor U11156 (N_11156,N_10846,N_10892);
nand U11157 (N_11157,N_10985,N_10890);
or U11158 (N_11158,N_10879,N_10866);
and U11159 (N_11159,N_10933,N_10811);
nor U11160 (N_11160,N_10927,N_10809);
xor U11161 (N_11161,N_10864,N_10819);
and U11162 (N_11162,N_10891,N_10843);
xnor U11163 (N_11163,N_10849,N_10829);
or U11164 (N_11164,N_10808,N_10853);
or U11165 (N_11165,N_10986,N_10883);
xor U11166 (N_11166,N_10809,N_10874);
xor U11167 (N_11167,N_10864,N_10888);
or U11168 (N_11168,N_10977,N_10850);
or U11169 (N_11169,N_10967,N_10930);
nor U11170 (N_11170,N_10886,N_10895);
or U11171 (N_11171,N_10940,N_10994);
xor U11172 (N_11172,N_10877,N_10841);
or U11173 (N_11173,N_10968,N_10833);
or U11174 (N_11174,N_10871,N_10847);
xnor U11175 (N_11175,N_10954,N_10905);
nor U11176 (N_11176,N_10936,N_10819);
xnor U11177 (N_11177,N_10858,N_10968);
xnor U11178 (N_11178,N_10977,N_10800);
and U11179 (N_11179,N_10826,N_10914);
nor U11180 (N_11180,N_10999,N_10864);
nand U11181 (N_11181,N_10982,N_10873);
nand U11182 (N_11182,N_10864,N_10837);
nor U11183 (N_11183,N_10927,N_10937);
nand U11184 (N_11184,N_10920,N_10990);
nor U11185 (N_11185,N_10881,N_10802);
xor U11186 (N_11186,N_10992,N_10876);
nor U11187 (N_11187,N_10876,N_10899);
or U11188 (N_11188,N_10887,N_10987);
xor U11189 (N_11189,N_10863,N_10812);
nand U11190 (N_11190,N_10924,N_10840);
nand U11191 (N_11191,N_10958,N_10849);
nor U11192 (N_11192,N_10853,N_10834);
nand U11193 (N_11193,N_10886,N_10936);
and U11194 (N_11194,N_10904,N_10999);
nand U11195 (N_11195,N_10846,N_10935);
nand U11196 (N_11196,N_10914,N_10863);
nand U11197 (N_11197,N_10977,N_10863);
or U11198 (N_11198,N_10902,N_10867);
and U11199 (N_11199,N_10845,N_10871);
nand U11200 (N_11200,N_11114,N_11197);
and U11201 (N_11201,N_11168,N_11064);
xnor U11202 (N_11202,N_11193,N_11015);
or U11203 (N_11203,N_11179,N_11163);
nor U11204 (N_11204,N_11051,N_11127);
and U11205 (N_11205,N_11062,N_11180);
nand U11206 (N_11206,N_11037,N_11014);
nor U11207 (N_11207,N_11134,N_11147);
nor U11208 (N_11208,N_11145,N_11067);
nor U11209 (N_11209,N_11049,N_11059);
nand U11210 (N_11210,N_11189,N_11106);
nor U11211 (N_11211,N_11151,N_11133);
or U11212 (N_11212,N_11146,N_11034);
nand U11213 (N_11213,N_11043,N_11024);
nor U11214 (N_11214,N_11085,N_11105);
or U11215 (N_11215,N_11052,N_11162);
xnor U11216 (N_11216,N_11040,N_11028);
or U11217 (N_11217,N_11108,N_11002);
nand U11218 (N_11218,N_11148,N_11058);
or U11219 (N_11219,N_11131,N_11022);
or U11220 (N_11220,N_11017,N_11082);
or U11221 (N_11221,N_11126,N_11074);
nand U11222 (N_11222,N_11160,N_11141);
and U11223 (N_11223,N_11050,N_11175);
nor U11224 (N_11224,N_11087,N_11035);
nor U11225 (N_11225,N_11054,N_11078);
or U11226 (N_11226,N_11194,N_11166);
nand U11227 (N_11227,N_11096,N_11107);
xnor U11228 (N_11228,N_11068,N_11120);
and U11229 (N_11229,N_11007,N_11188);
nand U11230 (N_11230,N_11029,N_11178);
or U11231 (N_11231,N_11153,N_11123);
nor U11232 (N_11232,N_11046,N_11139);
xnor U11233 (N_11233,N_11116,N_11138);
xor U11234 (N_11234,N_11185,N_11027);
and U11235 (N_11235,N_11083,N_11129);
or U11236 (N_11236,N_11143,N_11170);
nor U11237 (N_11237,N_11060,N_11005);
and U11238 (N_11238,N_11090,N_11113);
and U11239 (N_11239,N_11161,N_11081);
nand U11240 (N_11240,N_11169,N_11122);
xnor U11241 (N_11241,N_11065,N_11155);
xor U11242 (N_11242,N_11048,N_11124);
nand U11243 (N_11243,N_11041,N_11154);
xnor U11244 (N_11244,N_11172,N_11019);
or U11245 (N_11245,N_11073,N_11110);
and U11246 (N_11246,N_11182,N_11056);
nand U11247 (N_11247,N_11196,N_11112);
xnor U11248 (N_11248,N_11199,N_11095);
nand U11249 (N_11249,N_11044,N_11021);
xnor U11250 (N_11250,N_11069,N_11186);
xnor U11251 (N_11251,N_11103,N_11157);
xnor U11252 (N_11252,N_11176,N_11076);
nor U11253 (N_11253,N_11130,N_11158);
xor U11254 (N_11254,N_11000,N_11091);
and U11255 (N_11255,N_11026,N_11006);
nand U11256 (N_11256,N_11140,N_11117);
nor U11257 (N_11257,N_11165,N_11198);
or U11258 (N_11258,N_11063,N_11086);
xnor U11259 (N_11259,N_11047,N_11101);
nand U11260 (N_11260,N_11039,N_11174);
and U11261 (N_11261,N_11012,N_11079);
xor U11262 (N_11262,N_11032,N_11042);
xnor U11263 (N_11263,N_11094,N_11070);
nor U11264 (N_11264,N_11190,N_11077);
nor U11265 (N_11265,N_11115,N_11100);
and U11266 (N_11266,N_11098,N_11066);
or U11267 (N_11267,N_11003,N_11125);
nor U11268 (N_11268,N_11075,N_11033);
or U11269 (N_11269,N_11030,N_11025);
xor U11270 (N_11270,N_11057,N_11121);
or U11271 (N_11271,N_11099,N_11156);
nand U11272 (N_11272,N_11132,N_11159);
and U11273 (N_11273,N_11195,N_11184);
nor U11274 (N_11274,N_11020,N_11038);
or U11275 (N_11275,N_11128,N_11137);
nand U11276 (N_11276,N_11008,N_11055);
nor U11277 (N_11277,N_11009,N_11097);
and U11278 (N_11278,N_11102,N_11152);
and U11279 (N_11279,N_11192,N_11164);
nor U11280 (N_11280,N_11045,N_11088);
and U11281 (N_11281,N_11092,N_11142);
nand U11282 (N_11282,N_11135,N_11013);
and U11283 (N_11283,N_11001,N_11104);
and U11284 (N_11284,N_11053,N_11093);
xor U11285 (N_11285,N_11018,N_11010);
or U11286 (N_11286,N_11187,N_11080);
or U11287 (N_11287,N_11004,N_11089);
nor U11288 (N_11288,N_11061,N_11167);
nor U11289 (N_11289,N_11071,N_11011);
nor U11290 (N_11290,N_11023,N_11036);
or U11291 (N_11291,N_11136,N_11118);
xor U11292 (N_11292,N_11144,N_11177);
nor U11293 (N_11293,N_11119,N_11072);
nand U11294 (N_11294,N_11031,N_11191);
nor U11295 (N_11295,N_11016,N_11173);
nor U11296 (N_11296,N_11149,N_11084);
xnor U11297 (N_11297,N_11183,N_11181);
or U11298 (N_11298,N_11150,N_11171);
nand U11299 (N_11299,N_11111,N_11109);
nor U11300 (N_11300,N_11041,N_11183);
or U11301 (N_11301,N_11119,N_11089);
and U11302 (N_11302,N_11142,N_11178);
xnor U11303 (N_11303,N_11081,N_11130);
nor U11304 (N_11304,N_11166,N_11119);
xor U11305 (N_11305,N_11150,N_11162);
nand U11306 (N_11306,N_11097,N_11181);
nor U11307 (N_11307,N_11007,N_11100);
nor U11308 (N_11308,N_11150,N_11083);
or U11309 (N_11309,N_11156,N_11058);
nor U11310 (N_11310,N_11133,N_11066);
xnor U11311 (N_11311,N_11184,N_11147);
nand U11312 (N_11312,N_11196,N_11085);
xor U11313 (N_11313,N_11017,N_11149);
and U11314 (N_11314,N_11084,N_11073);
nor U11315 (N_11315,N_11050,N_11140);
nand U11316 (N_11316,N_11025,N_11155);
nor U11317 (N_11317,N_11100,N_11096);
nor U11318 (N_11318,N_11008,N_11135);
xor U11319 (N_11319,N_11036,N_11093);
and U11320 (N_11320,N_11034,N_11153);
xnor U11321 (N_11321,N_11164,N_11022);
or U11322 (N_11322,N_11007,N_11019);
nand U11323 (N_11323,N_11109,N_11089);
nor U11324 (N_11324,N_11008,N_11157);
nor U11325 (N_11325,N_11061,N_11194);
or U11326 (N_11326,N_11066,N_11151);
xnor U11327 (N_11327,N_11077,N_11135);
nor U11328 (N_11328,N_11096,N_11050);
nand U11329 (N_11329,N_11015,N_11073);
or U11330 (N_11330,N_11014,N_11160);
nand U11331 (N_11331,N_11142,N_11009);
nor U11332 (N_11332,N_11167,N_11015);
and U11333 (N_11333,N_11149,N_11075);
nor U11334 (N_11334,N_11099,N_11030);
nor U11335 (N_11335,N_11182,N_11133);
nand U11336 (N_11336,N_11175,N_11041);
nor U11337 (N_11337,N_11040,N_11122);
xnor U11338 (N_11338,N_11020,N_11047);
nand U11339 (N_11339,N_11063,N_11037);
xnor U11340 (N_11340,N_11049,N_11153);
nor U11341 (N_11341,N_11137,N_11134);
or U11342 (N_11342,N_11148,N_11064);
nor U11343 (N_11343,N_11068,N_11109);
and U11344 (N_11344,N_11029,N_11034);
and U11345 (N_11345,N_11044,N_11154);
xnor U11346 (N_11346,N_11130,N_11139);
xnor U11347 (N_11347,N_11113,N_11172);
xor U11348 (N_11348,N_11071,N_11053);
or U11349 (N_11349,N_11196,N_11098);
nor U11350 (N_11350,N_11016,N_11139);
and U11351 (N_11351,N_11087,N_11027);
and U11352 (N_11352,N_11025,N_11198);
or U11353 (N_11353,N_11106,N_11129);
nor U11354 (N_11354,N_11002,N_11150);
nand U11355 (N_11355,N_11145,N_11079);
nand U11356 (N_11356,N_11169,N_11179);
and U11357 (N_11357,N_11025,N_11156);
and U11358 (N_11358,N_11001,N_11187);
or U11359 (N_11359,N_11091,N_11020);
xnor U11360 (N_11360,N_11129,N_11107);
and U11361 (N_11361,N_11084,N_11137);
xnor U11362 (N_11362,N_11056,N_11082);
xor U11363 (N_11363,N_11016,N_11155);
or U11364 (N_11364,N_11169,N_11000);
xnor U11365 (N_11365,N_11012,N_11092);
xor U11366 (N_11366,N_11130,N_11104);
and U11367 (N_11367,N_11120,N_11063);
xnor U11368 (N_11368,N_11048,N_11164);
nand U11369 (N_11369,N_11099,N_11184);
xor U11370 (N_11370,N_11019,N_11199);
nand U11371 (N_11371,N_11106,N_11140);
xor U11372 (N_11372,N_11052,N_11083);
xnor U11373 (N_11373,N_11163,N_11032);
nor U11374 (N_11374,N_11060,N_11009);
nand U11375 (N_11375,N_11016,N_11115);
nor U11376 (N_11376,N_11153,N_11091);
xnor U11377 (N_11377,N_11120,N_11019);
and U11378 (N_11378,N_11092,N_11174);
or U11379 (N_11379,N_11033,N_11056);
xnor U11380 (N_11380,N_11092,N_11030);
and U11381 (N_11381,N_11003,N_11047);
nand U11382 (N_11382,N_11127,N_11065);
nor U11383 (N_11383,N_11147,N_11136);
and U11384 (N_11384,N_11069,N_11198);
or U11385 (N_11385,N_11102,N_11150);
nand U11386 (N_11386,N_11131,N_11002);
nand U11387 (N_11387,N_11024,N_11178);
or U11388 (N_11388,N_11088,N_11068);
and U11389 (N_11389,N_11112,N_11107);
or U11390 (N_11390,N_11134,N_11020);
nand U11391 (N_11391,N_11191,N_11197);
xor U11392 (N_11392,N_11023,N_11005);
and U11393 (N_11393,N_11105,N_11130);
xor U11394 (N_11394,N_11151,N_11197);
nor U11395 (N_11395,N_11101,N_11060);
and U11396 (N_11396,N_11029,N_11085);
nor U11397 (N_11397,N_11171,N_11100);
xor U11398 (N_11398,N_11035,N_11089);
and U11399 (N_11399,N_11067,N_11162);
and U11400 (N_11400,N_11379,N_11357);
and U11401 (N_11401,N_11229,N_11276);
or U11402 (N_11402,N_11368,N_11376);
nor U11403 (N_11403,N_11392,N_11299);
nand U11404 (N_11404,N_11297,N_11257);
nor U11405 (N_11405,N_11285,N_11304);
xnor U11406 (N_11406,N_11355,N_11256);
nand U11407 (N_11407,N_11288,N_11317);
and U11408 (N_11408,N_11373,N_11221);
xor U11409 (N_11409,N_11273,N_11303);
nand U11410 (N_11410,N_11371,N_11334);
and U11411 (N_11411,N_11251,N_11301);
xor U11412 (N_11412,N_11397,N_11306);
or U11413 (N_11413,N_11222,N_11252);
nand U11414 (N_11414,N_11321,N_11372);
xor U11415 (N_11415,N_11282,N_11226);
and U11416 (N_11416,N_11289,N_11325);
or U11417 (N_11417,N_11242,N_11202);
or U11418 (N_11418,N_11220,N_11388);
xor U11419 (N_11419,N_11363,N_11227);
nand U11420 (N_11420,N_11342,N_11259);
xnor U11421 (N_11421,N_11309,N_11267);
nor U11422 (N_11422,N_11211,N_11263);
or U11423 (N_11423,N_11340,N_11295);
xor U11424 (N_11424,N_11380,N_11359);
nand U11425 (N_11425,N_11389,N_11294);
and U11426 (N_11426,N_11287,N_11322);
nor U11427 (N_11427,N_11228,N_11208);
or U11428 (N_11428,N_11284,N_11341);
and U11429 (N_11429,N_11270,N_11356);
xor U11430 (N_11430,N_11366,N_11358);
nor U11431 (N_11431,N_11250,N_11328);
or U11432 (N_11432,N_11308,N_11272);
or U11433 (N_11433,N_11315,N_11383);
xnor U11434 (N_11434,N_11277,N_11262);
and U11435 (N_11435,N_11245,N_11378);
nor U11436 (N_11436,N_11348,N_11247);
or U11437 (N_11437,N_11329,N_11236);
nand U11438 (N_11438,N_11332,N_11286);
or U11439 (N_11439,N_11337,N_11339);
nor U11440 (N_11440,N_11291,N_11253);
xor U11441 (N_11441,N_11369,N_11360);
nor U11442 (N_11442,N_11246,N_11324);
nand U11443 (N_11443,N_11201,N_11384);
or U11444 (N_11444,N_11361,N_11223);
nand U11445 (N_11445,N_11393,N_11327);
nor U11446 (N_11446,N_11314,N_11338);
or U11447 (N_11447,N_11258,N_11346);
or U11448 (N_11448,N_11215,N_11311);
xnor U11449 (N_11449,N_11224,N_11362);
or U11450 (N_11450,N_11264,N_11239);
and U11451 (N_11451,N_11231,N_11399);
and U11452 (N_11452,N_11254,N_11290);
or U11453 (N_11453,N_11292,N_11374);
xor U11454 (N_11454,N_11218,N_11232);
nor U11455 (N_11455,N_11278,N_11249);
nor U11456 (N_11456,N_11336,N_11205);
xnor U11457 (N_11457,N_11293,N_11302);
nor U11458 (N_11458,N_11313,N_11310);
nand U11459 (N_11459,N_11330,N_11333);
nand U11460 (N_11460,N_11391,N_11381);
and U11461 (N_11461,N_11386,N_11350);
or U11462 (N_11462,N_11283,N_11300);
xor U11463 (N_11463,N_11279,N_11255);
nand U11464 (N_11464,N_11234,N_11260);
nor U11465 (N_11465,N_11396,N_11209);
and U11466 (N_11466,N_11269,N_11225);
or U11467 (N_11467,N_11206,N_11237);
or U11468 (N_11468,N_11323,N_11244);
nand U11469 (N_11469,N_11354,N_11216);
nor U11470 (N_11470,N_11230,N_11320);
nand U11471 (N_11471,N_11200,N_11387);
nand U11472 (N_11472,N_11265,N_11395);
nand U11473 (N_11473,N_11210,N_11345);
and U11474 (N_11474,N_11207,N_11280);
xor U11475 (N_11475,N_11261,N_11349);
nand U11476 (N_11476,N_11233,N_11275);
nor U11477 (N_11477,N_11312,N_11235);
nor U11478 (N_11478,N_11365,N_11319);
xnor U11479 (N_11479,N_11335,N_11351);
and U11480 (N_11480,N_11347,N_11219);
xor U11481 (N_11481,N_11398,N_11394);
or U11482 (N_11482,N_11377,N_11353);
xnor U11483 (N_11483,N_11241,N_11248);
or U11484 (N_11484,N_11274,N_11214);
nor U11485 (N_11485,N_11217,N_11375);
nand U11486 (N_11486,N_11203,N_11212);
and U11487 (N_11487,N_11213,N_11364);
nor U11488 (N_11488,N_11266,N_11370);
xnor U11489 (N_11489,N_11204,N_11298);
nand U11490 (N_11490,N_11390,N_11382);
xor U11491 (N_11491,N_11316,N_11243);
xnor U11492 (N_11492,N_11305,N_11268);
nand U11493 (N_11493,N_11344,N_11318);
and U11494 (N_11494,N_11385,N_11367);
nand U11495 (N_11495,N_11326,N_11281);
or U11496 (N_11496,N_11352,N_11238);
nor U11497 (N_11497,N_11331,N_11271);
and U11498 (N_11498,N_11296,N_11343);
nor U11499 (N_11499,N_11307,N_11240);
or U11500 (N_11500,N_11291,N_11228);
nand U11501 (N_11501,N_11388,N_11249);
nand U11502 (N_11502,N_11232,N_11287);
xnor U11503 (N_11503,N_11333,N_11249);
or U11504 (N_11504,N_11269,N_11306);
or U11505 (N_11505,N_11304,N_11214);
or U11506 (N_11506,N_11339,N_11277);
nand U11507 (N_11507,N_11395,N_11372);
nand U11508 (N_11508,N_11251,N_11246);
or U11509 (N_11509,N_11334,N_11391);
nor U11510 (N_11510,N_11217,N_11371);
nand U11511 (N_11511,N_11211,N_11373);
xnor U11512 (N_11512,N_11226,N_11365);
nand U11513 (N_11513,N_11240,N_11335);
xor U11514 (N_11514,N_11320,N_11317);
nand U11515 (N_11515,N_11378,N_11381);
and U11516 (N_11516,N_11375,N_11352);
nand U11517 (N_11517,N_11357,N_11300);
nor U11518 (N_11518,N_11323,N_11377);
nand U11519 (N_11519,N_11292,N_11343);
and U11520 (N_11520,N_11218,N_11282);
xnor U11521 (N_11521,N_11320,N_11234);
xnor U11522 (N_11522,N_11272,N_11393);
nor U11523 (N_11523,N_11244,N_11269);
xnor U11524 (N_11524,N_11369,N_11336);
nand U11525 (N_11525,N_11358,N_11331);
xnor U11526 (N_11526,N_11312,N_11256);
xnor U11527 (N_11527,N_11297,N_11393);
nor U11528 (N_11528,N_11222,N_11375);
nand U11529 (N_11529,N_11396,N_11299);
nand U11530 (N_11530,N_11379,N_11226);
nor U11531 (N_11531,N_11205,N_11375);
or U11532 (N_11532,N_11362,N_11313);
or U11533 (N_11533,N_11256,N_11284);
and U11534 (N_11534,N_11216,N_11384);
and U11535 (N_11535,N_11200,N_11228);
and U11536 (N_11536,N_11312,N_11265);
xnor U11537 (N_11537,N_11365,N_11204);
xor U11538 (N_11538,N_11283,N_11261);
xor U11539 (N_11539,N_11366,N_11372);
nor U11540 (N_11540,N_11282,N_11275);
xnor U11541 (N_11541,N_11215,N_11392);
or U11542 (N_11542,N_11388,N_11290);
or U11543 (N_11543,N_11231,N_11220);
or U11544 (N_11544,N_11249,N_11253);
or U11545 (N_11545,N_11304,N_11257);
and U11546 (N_11546,N_11346,N_11382);
xor U11547 (N_11547,N_11314,N_11356);
or U11548 (N_11548,N_11218,N_11222);
and U11549 (N_11549,N_11395,N_11212);
nand U11550 (N_11550,N_11386,N_11395);
and U11551 (N_11551,N_11206,N_11207);
xnor U11552 (N_11552,N_11326,N_11355);
nor U11553 (N_11553,N_11219,N_11244);
or U11554 (N_11554,N_11230,N_11202);
nor U11555 (N_11555,N_11389,N_11233);
or U11556 (N_11556,N_11340,N_11213);
xor U11557 (N_11557,N_11308,N_11219);
nor U11558 (N_11558,N_11207,N_11224);
nand U11559 (N_11559,N_11228,N_11272);
nand U11560 (N_11560,N_11380,N_11247);
xor U11561 (N_11561,N_11393,N_11396);
nand U11562 (N_11562,N_11247,N_11261);
and U11563 (N_11563,N_11317,N_11269);
and U11564 (N_11564,N_11365,N_11387);
nor U11565 (N_11565,N_11339,N_11363);
xnor U11566 (N_11566,N_11347,N_11306);
nand U11567 (N_11567,N_11319,N_11353);
and U11568 (N_11568,N_11251,N_11382);
and U11569 (N_11569,N_11276,N_11240);
xor U11570 (N_11570,N_11216,N_11206);
nand U11571 (N_11571,N_11263,N_11249);
nand U11572 (N_11572,N_11367,N_11326);
nor U11573 (N_11573,N_11225,N_11307);
nor U11574 (N_11574,N_11311,N_11352);
xor U11575 (N_11575,N_11209,N_11285);
or U11576 (N_11576,N_11377,N_11389);
or U11577 (N_11577,N_11261,N_11222);
xnor U11578 (N_11578,N_11205,N_11341);
nand U11579 (N_11579,N_11217,N_11311);
or U11580 (N_11580,N_11322,N_11237);
nor U11581 (N_11581,N_11210,N_11387);
xnor U11582 (N_11582,N_11332,N_11212);
nand U11583 (N_11583,N_11327,N_11229);
or U11584 (N_11584,N_11392,N_11264);
xnor U11585 (N_11585,N_11310,N_11226);
nand U11586 (N_11586,N_11294,N_11282);
nor U11587 (N_11587,N_11260,N_11277);
xor U11588 (N_11588,N_11263,N_11288);
nand U11589 (N_11589,N_11222,N_11339);
nand U11590 (N_11590,N_11368,N_11253);
xnor U11591 (N_11591,N_11271,N_11318);
and U11592 (N_11592,N_11225,N_11251);
nand U11593 (N_11593,N_11243,N_11378);
nand U11594 (N_11594,N_11219,N_11273);
or U11595 (N_11595,N_11374,N_11250);
nor U11596 (N_11596,N_11214,N_11213);
nor U11597 (N_11597,N_11360,N_11213);
nand U11598 (N_11598,N_11399,N_11362);
or U11599 (N_11599,N_11293,N_11261);
xor U11600 (N_11600,N_11487,N_11559);
nor U11601 (N_11601,N_11585,N_11531);
and U11602 (N_11602,N_11533,N_11513);
xor U11603 (N_11603,N_11411,N_11481);
xnor U11604 (N_11604,N_11410,N_11518);
or U11605 (N_11605,N_11550,N_11443);
xor U11606 (N_11606,N_11579,N_11477);
and U11607 (N_11607,N_11425,N_11407);
or U11608 (N_11608,N_11509,N_11595);
xor U11609 (N_11609,N_11512,N_11575);
nand U11610 (N_11610,N_11536,N_11416);
or U11611 (N_11611,N_11534,N_11440);
nor U11612 (N_11612,N_11406,N_11590);
xor U11613 (N_11613,N_11572,N_11432);
nor U11614 (N_11614,N_11540,N_11589);
xnor U11615 (N_11615,N_11484,N_11593);
nor U11616 (N_11616,N_11529,N_11498);
nor U11617 (N_11617,N_11507,N_11598);
or U11618 (N_11618,N_11458,N_11420);
nand U11619 (N_11619,N_11426,N_11417);
xnor U11620 (N_11620,N_11453,N_11421);
and U11621 (N_11621,N_11478,N_11558);
and U11622 (N_11622,N_11496,N_11403);
xnor U11623 (N_11623,N_11448,N_11427);
nor U11624 (N_11624,N_11497,N_11402);
nor U11625 (N_11625,N_11409,N_11599);
and U11626 (N_11626,N_11460,N_11506);
xor U11627 (N_11627,N_11510,N_11490);
or U11628 (N_11628,N_11455,N_11560);
nor U11629 (N_11629,N_11594,N_11523);
or U11630 (N_11630,N_11555,N_11414);
nor U11631 (N_11631,N_11419,N_11588);
nor U11632 (N_11632,N_11582,N_11461);
or U11633 (N_11633,N_11517,N_11493);
and U11634 (N_11634,N_11538,N_11545);
nand U11635 (N_11635,N_11467,N_11505);
and U11636 (N_11636,N_11591,N_11544);
nand U11637 (N_11637,N_11501,N_11504);
nand U11638 (N_11638,N_11483,N_11454);
xnor U11639 (N_11639,N_11469,N_11479);
and U11640 (N_11640,N_11436,N_11489);
xnor U11641 (N_11641,N_11445,N_11462);
nand U11642 (N_11642,N_11400,N_11530);
or U11643 (N_11643,N_11564,N_11401);
xnor U11644 (N_11644,N_11480,N_11576);
and U11645 (N_11645,N_11514,N_11495);
nor U11646 (N_11646,N_11423,N_11566);
nor U11647 (N_11647,N_11474,N_11541);
and U11648 (N_11648,N_11553,N_11446);
or U11649 (N_11649,N_11431,N_11444);
nor U11650 (N_11650,N_11561,N_11494);
or U11651 (N_11651,N_11537,N_11568);
or U11652 (N_11652,N_11596,N_11449);
xnor U11653 (N_11653,N_11565,N_11442);
xor U11654 (N_11654,N_11503,N_11516);
xor U11655 (N_11655,N_11597,N_11557);
xor U11656 (N_11656,N_11580,N_11567);
xnor U11657 (N_11657,N_11476,N_11571);
and U11658 (N_11658,N_11468,N_11429);
nor U11659 (N_11659,N_11515,N_11470);
or U11660 (N_11660,N_11464,N_11511);
and U11661 (N_11661,N_11551,N_11570);
nand U11662 (N_11662,N_11422,N_11413);
nand U11663 (N_11663,N_11539,N_11578);
or U11664 (N_11664,N_11405,N_11592);
nand U11665 (N_11665,N_11428,N_11433);
xor U11666 (N_11666,N_11408,N_11430);
and U11667 (N_11667,N_11522,N_11418);
nand U11668 (N_11668,N_11577,N_11502);
xnor U11669 (N_11669,N_11482,N_11524);
or U11670 (N_11670,N_11486,N_11404);
xnor U11671 (N_11671,N_11535,N_11434);
and U11672 (N_11672,N_11532,N_11451);
nor U11673 (N_11673,N_11447,N_11439);
nand U11674 (N_11674,N_11528,N_11463);
nor U11675 (N_11675,N_11586,N_11475);
and U11676 (N_11676,N_11456,N_11508);
nand U11677 (N_11677,N_11548,N_11471);
nand U11678 (N_11678,N_11459,N_11581);
nor U11679 (N_11679,N_11525,N_11452);
or U11680 (N_11680,N_11527,N_11519);
nor U11681 (N_11681,N_11549,N_11450);
or U11682 (N_11682,N_11547,N_11546);
xor U11683 (N_11683,N_11554,N_11491);
nor U11684 (N_11684,N_11466,N_11520);
nor U11685 (N_11685,N_11500,N_11556);
xnor U11686 (N_11686,N_11499,N_11521);
xnor U11687 (N_11687,N_11587,N_11412);
and U11688 (N_11688,N_11424,N_11573);
nor U11689 (N_11689,N_11437,N_11526);
or U11690 (N_11690,N_11457,N_11574);
and U11691 (N_11691,N_11563,N_11415);
or U11692 (N_11692,N_11542,N_11488);
and U11693 (N_11693,N_11465,N_11543);
and U11694 (N_11694,N_11562,N_11441);
and U11695 (N_11695,N_11492,N_11435);
nand U11696 (N_11696,N_11552,N_11584);
xor U11697 (N_11697,N_11485,N_11583);
or U11698 (N_11698,N_11438,N_11472);
nand U11699 (N_11699,N_11473,N_11569);
nor U11700 (N_11700,N_11462,N_11470);
nor U11701 (N_11701,N_11550,N_11427);
or U11702 (N_11702,N_11498,N_11537);
nor U11703 (N_11703,N_11431,N_11461);
nand U11704 (N_11704,N_11538,N_11513);
or U11705 (N_11705,N_11423,N_11483);
or U11706 (N_11706,N_11561,N_11546);
nand U11707 (N_11707,N_11592,N_11515);
or U11708 (N_11708,N_11570,N_11444);
nor U11709 (N_11709,N_11567,N_11483);
or U11710 (N_11710,N_11450,N_11464);
or U11711 (N_11711,N_11526,N_11486);
or U11712 (N_11712,N_11580,N_11462);
nor U11713 (N_11713,N_11495,N_11560);
xor U11714 (N_11714,N_11450,N_11462);
nand U11715 (N_11715,N_11599,N_11434);
nor U11716 (N_11716,N_11418,N_11439);
or U11717 (N_11717,N_11552,N_11507);
xnor U11718 (N_11718,N_11541,N_11507);
nand U11719 (N_11719,N_11507,N_11480);
xor U11720 (N_11720,N_11512,N_11480);
xnor U11721 (N_11721,N_11439,N_11489);
xor U11722 (N_11722,N_11433,N_11445);
nor U11723 (N_11723,N_11509,N_11468);
nor U11724 (N_11724,N_11534,N_11491);
nand U11725 (N_11725,N_11424,N_11498);
nor U11726 (N_11726,N_11524,N_11467);
and U11727 (N_11727,N_11586,N_11479);
xor U11728 (N_11728,N_11535,N_11598);
xnor U11729 (N_11729,N_11525,N_11458);
nor U11730 (N_11730,N_11417,N_11485);
xor U11731 (N_11731,N_11526,N_11513);
xnor U11732 (N_11732,N_11563,N_11417);
nand U11733 (N_11733,N_11415,N_11542);
xnor U11734 (N_11734,N_11509,N_11574);
and U11735 (N_11735,N_11446,N_11537);
nand U11736 (N_11736,N_11592,N_11537);
and U11737 (N_11737,N_11519,N_11549);
or U11738 (N_11738,N_11418,N_11502);
nor U11739 (N_11739,N_11518,N_11478);
and U11740 (N_11740,N_11530,N_11422);
or U11741 (N_11741,N_11404,N_11439);
nand U11742 (N_11742,N_11462,N_11501);
and U11743 (N_11743,N_11590,N_11400);
or U11744 (N_11744,N_11516,N_11480);
nor U11745 (N_11745,N_11542,N_11418);
nand U11746 (N_11746,N_11449,N_11506);
nor U11747 (N_11747,N_11595,N_11542);
or U11748 (N_11748,N_11433,N_11522);
or U11749 (N_11749,N_11571,N_11418);
nand U11750 (N_11750,N_11551,N_11542);
or U11751 (N_11751,N_11493,N_11524);
nand U11752 (N_11752,N_11583,N_11435);
xnor U11753 (N_11753,N_11468,N_11425);
and U11754 (N_11754,N_11457,N_11418);
nand U11755 (N_11755,N_11405,N_11535);
nor U11756 (N_11756,N_11560,N_11491);
nor U11757 (N_11757,N_11424,N_11515);
xnor U11758 (N_11758,N_11498,N_11555);
nor U11759 (N_11759,N_11451,N_11445);
nor U11760 (N_11760,N_11561,N_11418);
and U11761 (N_11761,N_11544,N_11493);
or U11762 (N_11762,N_11427,N_11487);
nor U11763 (N_11763,N_11416,N_11455);
or U11764 (N_11764,N_11545,N_11544);
nor U11765 (N_11765,N_11578,N_11483);
nor U11766 (N_11766,N_11462,N_11463);
nand U11767 (N_11767,N_11516,N_11499);
nand U11768 (N_11768,N_11413,N_11411);
nor U11769 (N_11769,N_11579,N_11439);
nand U11770 (N_11770,N_11436,N_11534);
nor U11771 (N_11771,N_11575,N_11447);
and U11772 (N_11772,N_11537,N_11493);
or U11773 (N_11773,N_11564,N_11431);
or U11774 (N_11774,N_11451,N_11597);
xnor U11775 (N_11775,N_11462,N_11440);
nand U11776 (N_11776,N_11485,N_11423);
xor U11777 (N_11777,N_11551,N_11400);
or U11778 (N_11778,N_11490,N_11461);
and U11779 (N_11779,N_11541,N_11471);
and U11780 (N_11780,N_11442,N_11570);
nand U11781 (N_11781,N_11556,N_11433);
and U11782 (N_11782,N_11593,N_11571);
or U11783 (N_11783,N_11538,N_11430);
nand U11784 (N_11784,N_11571,N_11444);
nor U11785 (N_11785,N_11415,N_11580);
nand U11786 (N_11786,N_11555,N_11464);
nand U11787 (N_11787,N_11584,N_11538);
or U11788 (N_11788,N_11418,N_11402);
nand U11789 (N_11789,N_11537,N_11589);
and U11790 (N_11790,N_11597,N_11545);
nor U11791 (N_11791,N_11437,N_11565);
and U11792 (N_11792,N_11456,N_11436);
nor U11793 (N_11793,N_11498,N_11503);
and U11794 (N_11794,N_11485,N_11524);
nand U11795 (N_11795,N_11592,N_11508);
nand U11796 (N_11796,N_11472,N_11433);
and U11797 (N_11797,N_11505,N_11439);
and U11798 (N_11798,N_11403,N_11549);
nand U11799 (N_11799,N_11439,N_11477);
xnor U11800 (N_11800,N_11677,N_11634);
xor U11801 (N_11801,N_11608,N_11694);
nor U11802 (N_11802,N_11788,N_11739);
nand U11803 (N_11803,N_11751,N_11779);
or U11804 (N_11804,N_11697,N_11723);
xnor U11805 (N_11805,N_11733,N_11729);
xnor U11806 (N_11806,N_11609,N_11686);
and U11807 (N_11807,N_11753,N_11630);
or U11808 (N_11808,N_11656,N_11737);
xnor U11809 (N_11809,N_11654,N_11773);
nor U11810 (N_11810,N_11695,N_11628);
and U11811 (N_11811,N_11727,N_11681);
and U11812 (N_11812,N_11692,N_11704);
or U11813 (N_11813,N_11642,N_11775);
or U11814 (N_11814,N_11719,N_11708);
and U11815 (N_11815,N_11669,N_11764);
or U11816 (N_11816,N_11629,N_11663);
nand U11817 (N_11817,N_11740,N_11760);
nand U11818 (N_11818,N_11651,N_11696);
xor U11819 (N_11819,N_11710,N_11678);
nand U11820 (N_11820,N_11780,N_11784);
and U11821 (N_11821,N_11635,N_11799);
and U11822 (N_11822,N_11641,N_11741);
nand U11823 (N_11823,N_11626,N_11755);
nor U11824 (N_11824,N_11643,N_11653);
nor U11825 (N_11825,N_11660,N_11665);
nor U11826 (N_11826,N_11790,N_11683);
xnor U11827 (N_11827,N_11690,N_11624);
and U11828 (N_11828,N_11722,N_11758);
nor U11829 (N_11829,N_11781,N_11794);
nor U11830 (N_11830,N_11714,N_11783);
or U11831 (N_11831,N_11752,N_11796);
nor U11832 (N_11832,N_11633,N_11770);
nor U11833 (N_11833,N_11750,N_11795);
nand U11834 (N_11834,N_11786,N_11668);
xnor U11835 (N_11835,N_11789,N_11709);
and U11836 (N_11836,N_11602,N_11646);
xor U11837 (N_11837,N_11620,N_11610);
nor U11838 (N_11838,N_11787,N_11728);
nor U11839 (N_11839,N_11615,N_11682);
xor U11840 (N_11840,N_11652,N_11631);
nor U11841 (N_11841,N_11691,N_11765);
xor U11842 (N_11842,N_11672,N_11685);
xor U11843 (N_11843,N_11711,N_11797);
nand U11844 (N_11844,N_11661,N_11618);
nor U11845 (N_11845,N_11613,N_11734);
xor U11846 (N_11846,N_11712,N_11627);
and U11847 (N_11847,N_11689,N_11724);
and U11848 (N_11848,N_11623,N_11607);
nor U11849 (N_11849,N_11720,N_11743);
xnor U11850 (N_11850,N_11707,N_11785);
or U11851 (N_11851,N_11671,N_11718);
or U11852 (N_11852,N_11745,N_11744);
or U11853 (N_11853,N_11670,N_11605);
or U11854 (N_11854,N_11732,N_11622);
nor U11855 (N_11855,N_11748,N_11679);
or U11856 (N_11856,N_11657,N_11636);
and U11857 (N_11857,N_11700,N_11638);
nor U11858 (N_11858,N_11747,N_11680);
or U11859 (N_11859,N_11778,N_11650);
xnor U11860 (N_11860,N_11791,N_11759);
nor U11861 (N_11861,N_11721,N_11632);
nand U11862 (N_11862,N_11767,N_11762);
nand U11863 (N_11863,N_11662,N_11798);
nand U11864 (N_11864,N_11617,N_11757);
xnor U11865 (N_11865,N_11639,N_11645);
nand U11866 (N_11866,N_11606,N_11738);
or U11867 (N_11867,N_11725,N_11731);
or U11868 (N_11868,N_11792,N_11612);
or U11869 (N_11869,N_11756,N_11676);
or U11870 (N_11870,N_11693,N_11674);
nor U11871 (N_11871,N_11619,N_11769);
or U11872 (N_11872,N_11621,N_11782);
and U11873 (N_11873,N_11649,N_11776);
or U11874 (N_11874,N_11614,N_11754);
and U11875 (N_11875,N_11648,N_11726);
nor U11876 (N_11876,N_11664,N_11735);
nor U11877 (N_11877,N_11698,N_11768);
xor U11878 (N_11878,N_11611,N_11713);
or U11879 (N_11879,N_11746,N_11640);
or U11880 (N_11880,N_11715,N_11699);
or U11881 (N_11881,N_11675,N_11644);
or U11882 (N_11882,N_11717,N_11742);
and U11883 (N_11883,N_11703,N_11774);
nor U11884 (N_11884,N_11777,N_11667);
and U11885 (N_11885,N_11655,N_11701);
or U11886 (N_11886,N_11730,N_11601);
nand U11887 (N_11887,N_11702,N_11684);
or U11888 (N_11888,N_11736,N_11604);
nor U11889 (N_11889,N_11688,N_11637);
and U11890 (N_11890,N_11749,N_11761);
xor U11891 (N_11891,N_11793,N_11705);
or U11892 (N_11892,N_11716,N_11771);
xnor U11893 (N_11893,N_11600,N_11659);
and U11894 (N_11894,N_11625,N_11603);
xnor U11895 (N_11895,N_11616,N_11766);
xor U11896 (N_11896,N_11706,N_11763);
nand U11897 (N_11897,N_11772,N_11666);
and U11898 (N_11898,N_11673,N_11647);
xnor U11899 (N_11899,N_11658,N_11687);
nor U11900 (N_11900,N_11667,N_11783);
nor U11901 (N_11901,N_11752,N_11640);
nor U11902 (N_11902,N_11782,N_11724);
xor U11903 (N_11903,N_11615,N_11611);
xnor U11904 (N_11904,N_11646,N_11777);
or U11905 (N_11905,N_11774,N_11672);
xnor U11906 (N_11906,N_11765,N_11698);
and U11907 (N_11907,N_11793,N_11678);
and U11908 (N_11908,N_11654,N_11661);
nor U11909 (N_11909,N_11693,N_11794);
and U11910 (N_11910,N_11613,N_11649);
or U11911 (N_11911,N_11708,N_11665);
and U11912 (N_11912,N_11619,N_11732);
and U11913 (N_11913,N_11745,N_11649);
nand U11914 (N_11914,N_11676,N_11788);
nor U11915 (N_11915,N_11626,N_11748);
or U11916 (N_11916,N_11699,N_11712);
nand U11917 (N_11917,N_11765,N_11769);
and U11918 (N_11918,N_11727,N_11756);
and U11919 (N_11919,N_11770,N_11686);
and U11920 (N_11920,N_11769,N_11789);
nor U11921 (N_11921,N_11718,N_11705);
nand U11922 (N_11922,N_11747,N_11714);
or U11923 (N_11923,N_11625,N_11787);
and U11924 (N_11924,N_11712,N_11784);
nor U11925 (N_11925,N_11602,N_11606);
or U11926 (N_11926,N_11617,N_11602);
nand U11927 (N_11927,N_11632,N_11783);
or U11928 (N_11928,N_11634,N_11757);
xnor U11929 (N_11929,N_11698,N_11612);
or U11930 (N_11930,N_11671,N_11676);
or U11931 (N_11931,N_11643,N_11673);
xor U11932 (N_11932,N_11680,N_11789);
nor U11933 (N_11933,N_11734,N_11704);
nand U11934 (N_11934,N_11761,N_11671);
and U11935 (N_11935,N_11729,N_11787);
nor U11936 (N_11936,N_11772,N_11775);
xor U11937 (N_11937,N_11691,N_11753);
xnor U11938 (N_11938,N_11752,N_11671);
xor U11939 (N_11939,N_11750,N_11646);
nor U11940 (N_11940,N_11753,N_11644);
and U11941 (N_11941,N_11679,N_11758);
nand U11942 (N_11942,N_11639,N_11682);
and U11943 (N_11943,N_11691,N_11693);
and U11944 (N_11944,N_11627,N_11769);
xor U11945 (N_11945,N_11701,N_11724);
or U11946 (N_11946,N_11717,N_11605);
and U11947 (N_11947,N_11681,N_11730);
nand U11948 (N_11948,N_11619,N_11765);
or U11949 (N_11949,N_11769,N_11680);
nand U11950 (N_11950,N_11756,N_11628);
nand U11951 (N_11951,N_11654,N_11754);
nor U11952 (N_11952,N_11709,N_11708);
xor U11953 (N_11953,N_11750,N_11660);
and U11954 (N_11954,N_11683,N_11727);
and U11955 (N_11955,N_11621,N_11709);
xnor U11956 (N_11956,N_11686,N_11683);
nand U11957 (N_11957,N_11672,N_11601);
nor U11958 (N_11958,N_11632,N_11647);
nor U11959 (N_11959,N_11669,N_11779);
nand U11960 (N_11960,N_11637,N_11639);
xnor U11961 (N_11961,N_11685,N_11706);
nor U11962 (N_11962,N_11699,N_11688);
nor U11963 (N_11963,N_11757,N_11774);
and U11964 (N_11964,N_11660,N_11794);
nand U11965 (N_11965,N_11648,N_11797);
nand U11966 (N_11966,N_11687,N_11701);
or U11967 (N_11967,N_11675,N_11681);
xnor U11968 (N_11968,N_11660,N_11657);
xor U11969 (N_11969,N_11772,N_11691);
xnor U11970 (N_11970,N_11763,N_11655);
nor U11971 (N_11971,N_11669,N_11777);
nor U11972 (N_11972,N_11755,N_11713);
nand U11973 (N_11973,N_11780,N_11745);
nand U11974 (N_11974,N_11746,N_11718);
nand U11975 (N_11975,N_11687,N_11674);
and U11976 (N_11976,N_11729,N_11707);
or U11977 (N_11977,N_11628,N_11747);
or U11978 (N_11978,N_11765,N_11662);
or U11979 (N_11979,N_11710,N_11729);
nand U11980 (N_11980,N_11758,N_11716);
and U11981 (N_11981,N_11761,N_11678);
nand U11982 (N_11982,N_11741,N_11746);
nand U11983 (N_11983,N_11716,N_11699);
and U11984 (N_11984,N_11797,N_11745);
nand U11985 (N_11985,N_11630,N_11759);
nor U11986 (N_11986,N_11716,N_11626);
nand U11987 (N_11987,N_11670,N_11687);
xnor U11988 (N_11988,N_11734,N_11611);
nor U11989 (N_11989,N_11777,N_11709);
and U11990 (N_11990,N_11719,N_11798);
and U11991 (N_11991,N_11794,N_11796);
and U11992 (N_11992,N_11611,N_11660);
xor U11993 (N_11993,N_11651,N_11756);
nand U11994 (N_11994,N_11724,N_11785);
and U11995 (N_11995,N_11750,N_11648);
xor U11996 (N_11996,N_11660,N_11744);
xnor U11997 (N_11997,N_11645,N_11731);
xor U11998 (N_11998,N_11608,N_11669);
and U11999 (N_11999,N_11714,N_11620);
xnor U12000 (N_12000,N_11979,N_11847);
and U12001 (N_12001,N_11951,N_11973);
nand U12002 (N_12002,N_11833,N_11867);
or U12003 (N_12003,N_11898,N_11976);
and U12004 (N_12004,N_11904,N_11994);
and U12005 (N_12005,N_11881,N_11888);
nor U12006 (N_12006,N_11877,N_11942);
and U12007 (N_12007,N_11985,N_11910);
nor U12008 (N_12008,N_11990,N_11997);
nor U12009 (N_12009,N_11981,N_11883);
nand U12010 (N_12010,N_11882,N_11943);
xor U12011 (N_12011,N_11952,N_11978);
nand U12012 (N_12012,N_11862,N_11961);
and U12013 (N_12013,N_11955,N_11921);
and U12014 (N_12014,N_11966,N_11860);
nor U12015 (N_12015,N_11930,N_11894);
or U12016 (N_12016,N_11923,N_11892);
and U12017 (N_12017,N_11809,N_11907);
or U12018 (N_12018,N_11989,N_11854);
nand U12019 (N_12019,N_11852,N_11840);
nor U12020 (N_12020,N_11993,N_11969);
nor U12021 (N_12021,N_11869,N_11836);
or U12022 (N_12022,N_11992,N_11940);
and U12023 (N_12023,N_11916,N_11948);
and U12024 (N_12024,N_11876,N_11900);
xnor U12025 (N_12025,N_11954,N_11807);
nor U12026 (N_12026,N_11846,N_11866);
nor U12027 (N_12027,N_11855,N_11804);
or U12028 (N_12028,N_11914,N_11863);
or U12029 (N_12029,N_11885,N_11988);
and U12030 (N_12030,N_11825,N_11822);
or U12031 (N_12031,N_11845,N_11811);
nor U12032 (N_12032,N_11972,N_11991);
nand U12033 (N_12033,N_11868,N_11995);
and U12034 (N_12034,N_11920,N_11896);
xor U12035 (N_12035,N_11927,N_11941);
xor U12036 (N_12036,N_11826,N_11932);
nor U12037 (N_12037,N_11899,N_11931);
xnor U12038 (N_12038,N_11873,N_11912);
and U12039 (N_12039,N_11949,N_11977);
and U12040 (N_12040,N_11837,N_11982);
nor U12041 (N_12041,N_11805,N_11925);
nand U12042 (N_12042,N_11959,N_11945);
and U12043 (N_12043,N_11851,N_11859);
and U12044 (N_12044,N_11929,N_11835);
and U12045 (N_12045,N_11820,N_11975);
xor U12046 (N_12046,N_11964,N_11938);
nand U12047 (N_12047,N_11908,N_11953);
xnor U12048 (N_12048,N_11950,N_11838);
and U12049 (N_12049,N_11830,N_11834);
and U12050 (N_12050,N_11870,N_11963);
and U12051 (N_12051,N_11816,N_11880);
xnor U12052 (N_12052,N_11824,N_11819);
nor U12053 (N_12053,N_11903,N_11817);
or U12054 (N_12054,N_11831,N_11909);
nor U12055 (N_12055,N_11874,N_11918);
nand U12056 (N_12056,N_11970,N_11803);
or U12057 (N_12057,N_11984,N_11968);
xor U12058 (N_12058,N_11893,N_11806);
nand U12059 (N_12059,N_11818,N_11810);
and U12060 (N_12060,N_11937,N_11857);
and U12061 (N_12061,N_11808,N_11839);
nor U12062 (N_12062,N_11983,N_11935);
nand U12063 (N_12063,N_11895,N_11971);
and U12064 (N_12064,N_11936,N_11832);
or U12065 (N_12065,N_11884,N_11957);
or U12066 (N_12066,N_11926,N_11865);
or U12067 (N_12067,N_11924,N_11815);
and U12068 (N_12068,N_11919,N_11889);
and U12069 (N_12069,N_11821,N_11879);
xnor U12070 (N_12070,N_11902,N_11913);
xor U12071 (N_12071,N_11823,N_11890);
nor U12072 (N_12072,N_11911,N_11917);
nand U12073 (N_12073,N_11843,N_11946);
or U12074 (N_12074,N_11986,N_11850);
or U12075 (N_12075,N_11956,N_11841);
nor U12076 (N_12076,N_11800,N_11887);
xor U12077 (N_12077,N_11934,N_11939);
nor U12078 (N_12078,N_11974,N_11965);
nand U12079 (N_12079,N_11897,N_11848);
xor U12080 (N_12080,N_11928,N_11858);
nand U12081 (N_12081,N_11844,N_11829);
nand U12082 (N_12082,N_11886,N_11996);
xnor U12083 (N_12083,N_11853,N_11891);
and U12084 (N_12084,N_11958,N_11813);
or U12085 (N_12085,N_11827,N_11814);
nand U12086 (N_12086,N_11861,N_11901);
or U12087 (N_12087,N_11801,N_11842);
and U12088 (N_12088,N_11802,N_11906);
nand U12089 (N_12089,N_11915,N_11987);
nor U12090 (N_12090,N_11967,N_11878);
or U12091 (N_12091,N_11998,N_11947);
and U12092 (N_12092,N_11905,N_11849);
and U12093 (N_12093,N_11933,N_11960);
and U12094 (N_12094,N_11872,N_11962);
or U12095 (N_12095,N_11812,N_11999);
nor U12096 (N_12096,N_11828,N_11864);
nand U12097 (N_12097,N_11980,N_11871);
or U12098 (N_12098,N_11922,N_11944);
xor U12099 (N_12099,N_11875,N_11856);
nand U12100 (N_12100,N_11879,N_11854);
or U12101 (N_12101,N_11937,N_11963);
xnor U12102 (N_12102,N_11803,N_11992);
and U12103 (N_12103,N_11930,N_11803);
or U12104 (N_12104,N_11899,N_11871);
nand U12105 (N_12105,N_11942,N_11858);
xor U12106 (N_12106,N_11813,N_11843);
and U12107 (N_12107,N_11857,N_11977);
or U12108 (N_12108,N_11965,N_11871);
xor U12109 (N_12109,N_11889,N_11964);
nor U12110 (N_12110,N_11847,N_11922);
xnor U12111 (N_12111,N_11919,N_11812);
nor U12112 (N_12112,N_11894,N_11882);
nor U12113 (N_12113,N_11858,N_11897);
nand U12114 (N_12114,N_11859,N_11818);
xnor U12115 (N_12115,N_11945,N_11835);
nor U12116 (N_12116,N_11804,N_11936);
or U12117 (N_12117,N_11945,N_11838);
nand U12118 (N_12118,N_11871,N_11862);
nand U12119 (N_12119,N_11905,N_11921);
and U12120 (N_12120,N_11816,N_11936);
or U12121 (N_12121,N_11990,N_11810);
nor U12122 (N_12122,N_11936,N_11898);
and U12123 (N_12123,N_11975,N_11862);
or U12124 (N_12124,N_11989,N_11922);
or U12125 (N_12125,N_11880,N_11967);
or U12126 (N_12126,N_11949,N_11995);
nor U12127 (N_12127,N_11806,N_11957);
nand U12128 (N_12128,N_11978,N_11881);
and U12129 (N_12129,N_11893,N_11928);
xor U12130 (N_12130,N_11915,N_11896);
or U12131 (N_12131,N_11953,N_11850);
nand U12132 (N_12132,N_11871,N_11935);
nor U12133 (N_12133,N_11924,N_11928);
and U12134 (N_12134,N_11890,N_11853);
xnor U12135 (N_12135,N_11969,N_11856);
nor U12136 (N_12136,N_11807,N_11815);
or U12137 (N_12137,N_11862,N_11818);
and U12138 (N_12138,N_11941,N_11851);
and U12139 (N_12139,N_11904,N_11883);
nor U12140 (N_12140,N_11911,N_11876);
xor U12141 (N_12141,N_11996,N_11942);
or U12142 (N_12142,N_11960,N_11983);
or U12143 (N_12143,N_11815,N_11893);
xor U12144 (N_12144,N_11824,N_11826);
and U12145 (N_12145,N_11839,N_11988);
nor U12146 (N_12146,N_11990,N_11867);
or U12147 (N_12147,N_11892,N_11861);
xnor U12148 (N_12148,N_11899,N_11940);
and U12149 (N_12149,N_11897,N_11947);
nand U12150 (N_12150,N_11840,N_11877);
nand U12151 (N_12151,N_11805,N_11958);
nand U12152 (N_12152,N_11958,N_11850);
nor U12153 (N_12153,N_11932,N_11994);
or U12154 (N_12154,N_11950,N_11911);
xor U12155 (N_12155,N_11949,N_11886);
xor U12156 (N_12156,N_11885,N_11877);
nand U12157 (N_12157,N_11962,N_11864);
nand U12158 (N_12158,N_11968,N_11857);
nor U12159 (N_12159,N_11817,N_11901);
nor U12160 (N_12160,N_11965,N_11932);
or U12161 (N_12161,N_11900,N_11951);
nand U12162 (N_12162,N_11913,N_11877);
and U12163 (N_12163,N_11801,N_11993);
xnor U12164 (N_12164,N_11888,N_11926);
nand U12165 (N_12165,N_11802,N_11988);
and U12166 (N_12166,N_11911,N_11947);
nand U12167 (N_12167,N_11903,N_11915);
and U12168 (N_12168,N_11975,N_11970);
nand U12169 (N_12169,N_11979,N_11939);
or U12170 (N_12170,N_11917,N_11943);
nor U12171 (N_12171,N_11901,N_11920);
nand U12172 (N_12172,N_11918,N_11973);
nor U12173 (N_12173,N_11806,N_11955);
nand U12174 (N_12174,N_11876,N_11935);
nand U12175 (N_12175,N_11882,N_11949);
and U12176 (N_12176,N_11837,N_11920);
xor U12177 (N_12177,N_11944,N_11986);
xnor U12178 (N_12178,N_11825,N_11860);
nor U12179 (N_12179,N_11935,N_11995);
or U12180 (N_12180,N_11923,N_11916);
nor U12181 (N_12181,N_11916,N_11904);
nand U12182 (N_12182,N_11870,N_11912);
or U12183 (N_12183,N_11989,N_11809);
xor U12184 (N_12184,N_11877,N_11821);
and U12185 (N_12185,N_11907,N_11990);
and U12186 (N_12186,N_11946,N_11918);
and U12187 (N_12187,N_11957,N_11843);
and U12188 (N_12188,N_11916,N_11819);
or U12189 (N_12189,N_11951,N_11911);
xnor U12190 (N_12190,N_11976,N_11924);
nand U12191 (N_12191,N_11917,N_11958);
and U12192 (N_12192,N_11955,N_11984);
nand U12193 (N_12193,N_11932,N_11908);
nand U12194 (N_12194,N_11901,N_11857);
nor U12195 (N_12195,N_11881,N_11829);
and U12196 (N_12196,N_11876,N_11848);
or U12197 (N_12197,N_11904,N_11964);
and U12198 (N_12198,N_11957,N_11852);
nor U12199 (N_12199,N_11857,N_11996);
and U12200 (N_12200,N_12065,N_12024);
or U12201 (N_12201,N_12197,N_12171);
or U12202 (N_12202,N_12051,N_12049);
nor U12203 (N_12203,N_12000,N_12156);
nand U12204 (N_12204,N_12083,N_12189);
xnor U12205 (N_12205,N_12195,N_12035);
xor U12206 (N_12206,N_12084,N_12145);
nor U12207 (N_12207,N_12080,N_12126);
nor U12208 (N_12208,N_12002,N_12079);
nand U12209 (N_12209,N_12069,N_12188);
xor U12210 (N_12210,N_12177,N_12157);
nor U12211 (N_12211,N_12064,N_12030);
nand U12212 (N_12212,N_12076,N_12068);
nor U12213 (N_12213,N_12120,N_12115);
or U12214 (N_12214,N_12181,N_12004);
xor U12215 (N_12215,N_12165,N_12057);
xnor U12216 (N_12216,N_12182,N_12152);
nor U12217 (N_12217,N_12167,N_12173);
and U12218 (N_12218,N_12164,N_12070);
and U12219 (N_12219,N_12021,N_12141);
xnor U12220 (N_12220,N_12031,N_12025);
xor U12221 (N_12221,N_12113,N_12135);
nor U12222 (N_12222,N_12052,N_12110);
and U12223 (N_12223,N_12108,N_12046);
or U12224 (N_12224,N_12194,N_12198);
nand U12225 (N_12225,N_12066,N_12101);
nor U12226 (N_12226,N_12158,N_12151);
nand U12227 (N_12227,N_12116,N_12047);
and U12228 (N_12228,N_12143,N_12096);
xor U12229 (N_12229,N_12043,N_12174);
nand U12230 (N_12230,N_12100,N_12048);
xor U12231 (N_12231,N_12040,N_12095);
nor U12232 (N_12232,N_12038,N_12137);
or U12233 (N_12233,N_12099,N_12027);
or U12234 (N_12234,N_12092,N_12082);
nand U12235 (N_12235,N_12187,N_12078);
nor U12236 (N_12236,N_12153,N_12148);
or U12237 (N_12237,N_12125,N_12150);
xnor U12238 (N_12238,N_12106,N_12107);
or U12239 (N_12239,N_12013,N_12199);
and U12240 (N_12240,N_12018,N_12063);
xor U12241 (N_12241,N_12022,N_12073);
xor U12242 (N_12242,N_12044,N_12142);
xor U12243 (N_12243,N_12196,N_12020);
xor U12244 (N_12244,N_12118,N_12178);
or U12245 (N_12245,N_12071,N_12124);
nor U12246 (N_12246,N_12131,N_12132);
and U12247 (N_12247,N_12041,N_12159);
or U12248 (N_12248,N_12146,N_12098);
and U12249 (N_12249,N_12036,N_12185);
or U12250 (N_12250,N_12033,N_12128);
xor U12251 (N_12251,N_12190,N_12161);
nand U12252 (N_12252,N_12179,N_12121);
xnor U12253 (N_12253,N_12055,N_12169);
or U12254 (N_12254,N_12147,N_12129);
and U12255 (N_12255,N_12184,N_12193);
xor U12256 (N_12256,N_12077,N_12001);
and U12257 (N_12257,N_12087,N_12006);
and U12258 (N_12258,N_12176,N_12103);
nor U12259 (N_12259,N_12058,N_12054);
nor U12260 (N_12260,N_12032,N_12061);
xor U12261 (N_12261,N_12136,N_12160);
nand U12262 (N_12262,N_12130,N_12149);
nand U12263 (N_12263,N_12138,N_12155);
nor U12264 (N_12264,N_12028,N_12093);
xor U12265 (N_12265,N_12045,N_12042);
nor U12266 (N_12266,N_12060,N_12029);
or U12267 (N_12267,N_12140,N_12191);
or U12268 (N_12268,N_12162,N_12056);
and U12269 (N_12269,N_12163,N_12019);
xor U12270 (N_12270,N_12117,N_12088);
and U12271 (N_12271,N_12123,N_12183);
and U12272 (N_12272,N_12144,N_12015);
xnor U12273 (N_12273,N_12166,N_12114);
and U12274 (N_12274,N_12005,N_12111);
or U12275 (N_12275,N_12012,N_12172);
or U12276 (N_12276,N_12139,N_12180);
xor U12277 (N_12277,N_12089,N_12094);
nor U12278 (N_12278,N_12085,N_12026);
and U12279 (N_12279,N_12081,N_12011);
or U12280 (N_12280,N_12109,N_12039);
nor U12281 (N_12281,N_12127,N_12010);
and U12282 (N_12282,N_12014,N_12168);
or U12283 (N_12283,N_12023,N_12072);
xor U12284 (N_12284,N_12090,N_12009);
or U12285 (N_12285,N_12053,N_12122);
and U12286 (N_12286,N_12016,N_12104);
xnor U12287 (N_12287,N_12175,N_12037);
or U12288 (N_12288,N_12050,N_12097);
xnor U12289 (N_12289,N_12186,N_12075);
and U12290 (N_12290,N_12059,N_12086);
nor U12291 (N_12291,N_12119,N_12003);
xnor U12292 (N_12292,N_12062,N_12102);
or U12293 (N_12293,N_12008,N_12034);
xnor U12294 (N_12294,N_12074,N_12112);
xor U12295 (N_12295,N_12091,N_12067);
nor U12296 (N_12296,N_12154,N_12192);
xnor U12297 (N_12297,N_12133,N_12007);
and U12298 (N_12298,N_12105,N_12017);
nand U12299 (N_12299,N_12134,N_12170);
or U12300 (N_12300,N_12030,N_12193);
nor U12301 (N_12301,N_12104,N_12152);
and U12302 (N_12302,N_12050,N_12079);
or U12303 (N_12303,N_12034,N_12043);
or U12304 (N_12304,N_12083,N_12041);
and U12305 (N_12305,N_12066,N_12031);
and U12306 (N_12306,N_12156,N_12108);
and U12307 (N_12307,N_12002,N_12123);
nand U12308 (N_12308,N_12077,N_12063);
or U12309 (N_12309,N_12065,N_12146);
or U12310 (N_12310,N_12052,N_12164);
nand U12311 (N_12311,N_12047,N_12049);
or U12312 (N_12312,N_12014,N_12146);
xnor U12313 (N_12313,N_12096,N_12168);
xnor U12314 (N_12314,N_12072,N_12187);
xor U12315 (N_12315,N_12041,N_12192);
xnor U12316 (N_12316,N_12121,N_12074);
or U12317 (N_12317,N_12024,N_12082);
nand U12318 (N_12318,N_12093,N_12140);
nor U12319 (N_12319,N_12153,N_12156);
or U12320 (N_12320,N_12130,N_12116);
xor U12321 (N_12321,N_12110,N_12095);
or U12322 (N_12322,N_12181,N_12095);
and U12323 (N_12323,N_12132,N_12019);
and U12324 (N_12324,N_12038,N_12192);
nand U12325 (N_12325,N_12049,N_12058);
and U12326 (N_12326,N_12108,N_12163);
nand U12327 (N_12327,N_12070,N_12198);
and U12328 (N_12328,N_12102,N_12035);
xnor U12329 (N_12329,N_12123,N_12001);
and U12330 (N_12330,N_12185,N_12137);
or U12331 (N_12331,N_12072,N_12018);
nand U12332 (N_12332,N_12168,N_12197);
xnor U12333 (N_12333,N_12190,N_12023);
or U12334 (N_12334,N_12142,N_12063);
nand U12335 (N_12335,N_12115,N_12125);
xnor U12336 (N_12336,N_12146,N_12164);
or U12337 (N_12337,N_12174,N_12070);
or U12338 (N_12338,N_12103,N_12014);
xor U12339 (N_12339,N_12196,N_12072);
nor U12340 (N_12340,N_12048,N_12196);
nor U12341 (N_12341,N_12022,N_12083);
xnor U12342 (N_12342,N_12007,N_12124);
nand U12343 (N_12343,N_12036,N_12161);
or U12344 (N_12344,N_12120,N_12060);
nand U12345 (N_12345,N_12002,N_12033);
or U12346 (N_12346,N_12091,N_12079);
and U12347 (N_12347,N_12018,N_12013);
nand U12348 (N_12348,N_12035,N_12018);
and U12349 (N_12349,N_12182,N_12001);
nor U12350 (N_12350,N_12044,N_12066);
xor U12351 (N_12351,N_12158,N_12107);
or U12352 (N_12352,N_12187,N_12025);
nor U12353 (N_12353,N_12033,N_12126);
nor U12354 (N_12354,N_12105,N_12004);
or U12355 (N_12355,N_12116,N_12140);
and U12356 (N_12356,N_12126,N_12140);
xor U12357 (N_12357,N_12150,N_12138);
nand U12358 (N_12358,N_12009,N_12196);
and U12359 (N_12359,N_12004,N_12026);
nor U12360 (N_12360,N_12193,N_12099);
and U12361 (N_12361,N_12144,N_12084);
or U12362 (N_12362,N_12117,N_12095);
or U12363 (N_12363,N_12074,N_12095);
nand U12364 (N_12364,N_12028,N_12102);
xnor U12365 (N_12365,N_12113,N_12000);
nand U12366 (N_12366,N_12183,N_12125);
nand U12367 (N_12367,N_12030,N_12075);
and U12368 (N_12368,N_12101,N_12035);
or U12369 (N_12369,N_12169,N_12085);
xor U12370 (N_12370,N_12049,N_12026);
or U12371 (N_12371,N_12045,N_12114);
nand U12372 (N_12372,N_12183,N_12058);
or U12373 (N_12373,N_12018,N_12009);
or U12374 (N_12374,N_12016,N_12134);
and U12375 (N_12375,N_12106,N_12167);
nor U12376 (N_12376,N_12097,N_12182);
xor U12377 (N_12377,N_12036,N_12195);
xnor U12378 (N_12378,N_12025,N_12075);
or U12379 (N_12379,N_12164,N_12192);
or U12380 (N_12380,N_12178,N_12192);
xnor U12381 (N_12381,N_12016,N_12014);
nand U12382 (N_12382,N_12054,N_12001);
xor U12383 (N_12383,N_12005,N_12192);
nand U12384 (N_12384,N_12142,N_12148);
and U12385 (N_12385,N_12138,N_12179);
nor U12386 (N_12386,N_12075,N_12113);
xnor U12387 (N_12387,N_12072,N_12065);
or U12388 (N_12388,N_12161,N_12089);
nand U12389 (N_12389,N_12168,N_12116);
or U12390 (N_12390,N_12152,N_12057);
and U12391 (N_12391,N_12005,N_12084);
nand U12392 (N_12392,N_12070,N_12125);
and U12393 (N_12393,N_12194,N_12167);
xnor U12394 (N_12394,N_12173,N_12055);
and U12395 (N_12395,N_12113,N_12167);
or U12396 (N_12396,N_12188,N_12110);
and U12397 (N_12397,N_12036,N_12140);
nor U12398 (N_12398,N_12142,N_12159);
nor U12399 (N_12399,N_12110,N_12181);
or U12400 (N_12400,N_12296,N_12297);
nand U12401 (N_12401,N_12224,N_12288);
xnor U12402 (N_12402,N_12393,N_12289);
and U12403 (N_12403,N_12353,N_12348);
and U12404 (N_12404,N_12314,N_12385);
nand U12405 (N_12405,N_12293,N_12213);
and U12406 (N_12406,N_12392,N_12240);
nand U12407 (N_12407,N_12202,N_12276);
nand U12408 (N_12408,N_12390,N_12265);
or U12409 (N_12409,N_12238,N_12247);
xnor U12410 (N_12410,N_12342,N_12271);
or U12411 (N_12411,N_12275,N_12231);
nand U12412 (N_12412,N_12267,N_12260);
or U12413 (N_12413,N_12388,N_12264);
and U12414 (N_12414,N_12220,N_12233);
xor U12415 (N_12415,N_12363,N_12345);
xnor U12416 (N_12416,N_12333,N_12237);
xor U12417 (N_12417,N_12295,N_12331);
or U12418 (N_12418,N_12281,N_12208);
nor U12419 (N_12419,N_12355,N_12382);
and U12420 (N_12420,N_12338,N_12313);
and U12421 (N_12421,N_12350,N_12266);
xnor U12422 (N_12422,N_12361,N_12327);
nand U12423 (N_12423,N_12322,N_12334);
nor U12424 (N_12424,N_12210,N_12349);
or U12425 (N_12425,N_12255,N_12308);
nor U12426 (N_12426,N_12230,N_12248);
and U12427 (N_12427,N_12311,N_12206);
nor U12428 (N_12428,N_12274,N_12364);
nand U12429 (N_12429,N_12228,N_12223);
and U12430 (N_12430,N_12347,N_12215);
nor U12431 (N_12431,N_12253,N_12239);
nand U12432 (N_12432,N_12212,N_12387);
nor U12433 (N_12433,N_12242,N_12346);
xnor U12434 (N_12434,N_12324,N_12398);
nor U12435 (N_12435,N_12243,N_12356);
xnor U12436 (N_12436,N_12203,N_12284);
and U12437 (N_12437,N_12290,N_12286);
nand U12438 (N_12438,N_12339,N_12298);
or U12439 (N_12439,N_12234,N_12357);
nand U12440 (N_12440,N_12383,N_12244);
nand U12441 (N_12441,N_12303,N_12258);
or U12442 (N_12442,N_12272,N_12365);
xnor U12443 (N_12443,N_12221,N_12323);
nor U12444 (N_12444,N_12367,N_12249);
xor U12445 (N_12445,N_12270,N_12378);
xnor U12446 (N_12446,N_12326,N_12257);
and U12447 (N_12447,N_12379,N_12394);
xor U12448 (N_12448,N_12211,N_12214);
xor U12449 (N_12449,N_12217,N_12321);
xnor U12450 (N_12450,N_12381,N_12374);
or U12451 (N_12451,N_12373,N_12307);
and U12452 (N_12452,N_12245,N_12225);
and U12453 (N_12453,N_12384,N_12268);
or U12454 (N_12454,N_12261,N_12391);
nand U12455 (N_12455,N_12287,N_12259);
nor U12456 (N_12456,N_12341,N_12377);
or U12457 (N_12457,N_12386,N_12252);
or U12458 (N_12458,N_12319,N_12344);
or U12459 (N_12459,N_12317,N_12219);
or U12460 (N_12460,N_12318,N_12285);
nand U12461 (N_12461,N_12320,N_12222);
and U12462 (N_12462,N_12335,N_12227);
and U12463 (N_12463,N_12325,N_12294);
nor U12464 (N_12464,N_12246,N_12269);
or U12465 (N_12465,N_12305,N_12336);
nand U12466 (N_12466,N_12304,N_12302);
nand U12467 (N_12467,N_12372,N_12280);
nor U12468 (N_12468,N_12209,N_12263);
xnor U12469 (N_12469,N_12236,N_12309);
and U12470 (N_12470,N_12358,N_12329);
or U12471 (N_12471,N_12312,N_12250);
and U12472 (N_12472,N_12337,N_12396);
or U12473 (N_12473,N_12397,N_12291);
xor U12474 (N_12474,N_12360,N_12254);
and U12475 (N_12475,N_12366,N_12251);
nor U12476 (N_12476,N_12389,N_12201);
or U12477 (N_12477,N_12399,N_12226);
or U12478 (N_12478,N_12256,N_12368);
nand U12479 (N_12479,N_12370,N_12310);
nor U12480 (N_12480,N_12205,N_12343);
nor U12481 (N_12481,N_12204,N_12300);
and U12482 (N_12482,N_12273,N_12316);
xnor U12483 (N_12483,N_12207,N_12229);
and U12484 (N_12484,N_12376,N_12315);
nor U12485 (N_12485,N_12301,N_12235);
nand U12486 (N_12486,N_12359,N_12218);
or U12487 (N_12487,N_12278,N_12283);
xor U12488 (N_12488,N_12216,N_12279);
xor U12489 (N_12489,N_12352,N_12375);
nor U12490 (N_12490,N_12369,N_12380);
or U12491 (N_12491,N_12371,N_12232);
xor U12492 (N_12492,N_12351,N_12328);
nor U12493 (N_12493,N_12395,N_12299);
nor U12494 (N_12494,N_12262,N_12332);
nor U12495 (N_12495,N_12200,N_12282);
nor U12496 (N_12496,N_12340,N_12277);
nor U12497 (N_12497,N_12292,N_12362);
or U12498 (N_12498,N_12330,N_12241);
and U12499 (N_12499,N_12354,N_12306);
nand U12500 (N_12500,N_12366,N_12340);
nor U12501 (N_12501,N_12261,N_12347);
xor U12502 (N_12502,N_12356,N_12221);
and U12503 (N_12503,N_12248,N_12345);
nand U12504 (N_12504,N_12226,N_12340);
nand U12505 (N_12505,N_12375,N_12290);
and U12506 (N_12506,N_12342,N_12276);
nor U12507 (N_12507,N_12288,N_12240);
xnor U12508 (N_12508,N_12365,N_12294);
xnor U12509 (N_12509,N_12313,N_12217);
or U12510 (N_12510,N_12275,N_12380);
or U12511 (N_12511,N_12215,N_12325);
nand U12512 (N_12512,N_12296,N_12202);
and U12513 (N_12513,N_12272,N_12345);
xnor U12514 (N_12514,N_12202,N_12292);
nand U12515 (N_12515,N_12279,N_12264);
and U12516 (N_12516,N_12211,N_12364);
or U12517 (N_12517,N_12204,N_12318);
nand U12518 (N_12518,N_12221,N_12392);
nand U12519 (N_12519,N_12363,N_12285);
and U12520 (N_12520,N_12298,N_12327);
and U12521 (N_12521,N_12256,N_12220);
or U12522 (N_12522,N_12342,N_12372);
nand U12523 (N_12523,N_12259,N_12222);
xnor U12524 (N_12524,N_12204,N_12351);
xor U12525 (N_12525,N_12252,N_12313);
nor U12526 (N_12526,N_12372,N_12338);
or U12527 (N_12527,N_12216,N_12290);
xnor U12528 (N_12528,N_12213,N_12233);
nor U12529 (N_12529,N_12397,N_12243);
or U12530 (N_12530,N_12219,N_12214);
and U12531 (N_12531,N_12217,N_12252);
nand U12532 (N_12532,N_12387,N_12296);
nor U12533 (N_12533,N_12227,N_12250);
xor U12534 (N_12534,N_12272,N_12210);
nor U12535 (N_12535,N_12376,N_12254);
or U12536 (N_12536,N_12308,N_12243);
nor U12537 (N_12537,N_12337,N_12299);
xor U12538 (N_12538,N_12399,N_12314);
nor U12539 (N_12539,N_12294,N_12364);
and U12540 (N_12540,N_12259,N_12211);
and U12541 (N_12541,N_12367,N_12371);
and U12542 (N_12542,N_12271,N_12359);
or U12543 (N_12543,N_12394,N_12348);
and U12544 (N_12544,N_12200,N_12299);
or U12545 (N_12545,N_12218,N_12273);
and U12546 (N_12546,N_12269,N_12308);
nand U12547 (N_12547,N_12313,N_12226);
xnor U12548 (N_12548,N_12394,N_12296);
and U12549 (N_12549,N_12236,N_12315);
nand U12550 (N_12550,N_12342,N_12287);
nand U12551 (N_12551,N_12368,N_12283);
xnor U12552 (N_12552,N_12395,N_12319);
nand U12553 (N_12553,N_12236,N_12372);
nand U12554 (N_12554,N_12372,N_12273);
or U12555 (N_12555,N_12220,N_12247);
nand U12556 (N_12556,N_12226,N_12347);
or U12557 (N_12557,N_12316,N_12201);
or U12558 (N_12558,N_12223,N_12268);
and U12559 (N_12559,N_12344,N_12283);
nor U12560 (N_12560,N_12224,N_12349);
or U12561 (N_12561,N_12265,N_12297);
xnor U12562 (N_12562,N_12296,N_12367);
or U12563 (N_12563,N_12233,N_12203);
nand U12564 (N_12564,N_12258,N_12269);
nand U12565 (N_12565,N_12372,N_12245);
xnor U12566 (N_12566,N_12273,N_12301);
or U12567 (N_12567,N_12229,N_12242);
xor U12568 (N_12568,N_12384,N_12295);
and U12569 (N_12569,N_12317,N_12232);
or U12570 (N_12570,N_12374,N_12280);
or U12571 (N_12571,N_12397,N_12310);
nand U12572 (N_12572,N_12251,N_12213);
xor U12573 (N_12573,N_12337,N_12255);
xor U12574 (N_12574,N_12260,N_12357);
and U12575 (N_12575,N_12218,N_12308);
and U12576 (N_12576,N_12371,N_12214);
and U12577 (N_12577,N_12201,N_12317);
nor U12578 (N_12578,N_12357,N_12334);
or U12579 (N_12579,N_12355,N_12270);
nand U12580 (N_12580,N_12216,N_12325);
nand U12581 (N_12581,N_12281,N_12261);
or U12582 (N_12582,N_12345,N_12214);
nor U12583 (N_12583,N_12226,N_12326);
xor U12584 (N_12584,N_12284,N_12292);
xnor U12585 (N_12585,N_12270,N_12265);
or U12586 (N_12586,N_12310,N_12323);
nor U12587 (N_12587,N_12243,N_12354);
and U12588 (N_12588,N_12240,N_12215);
nor U12589 (N_12589,N_12256,N_12230);
nand U12590 (N_12590,N_12315,N_12344);
nand U12591 (N_12591,N_12321,N_12392);
nor U12592 (N_12592,N_12241,N_12368);
nand U12593 (N_12593,N_12311,N_12277);
and U12594 (N_12594,N_12246,N_12337);
nor U12595 (N_12595,N_12252,N_12219);
xnor U12596 (N_12596,N_12261,N_12334);
nand U12597 (N_12597,N_12357,N_12329);
or U12598 (N_12598,N_12288,N_12209);
or U12599 (N_12599,N_12286,N_12259);
and U12600 (N_12600,N_12402,N_12488);
and U12601 (N_12601,N_12516,N_12520);
nand U12602 (N_12602,N_12599,N_12475);
or U12603 (N_12603,N_12597,N_12587);
xor U12604 (N_12604,N_12550,N_12498);
nand U12605 (N_12605,N_12427,N_12552);
xor U12606 (N_12606,N_12580,N_12466);
and U12607 (N_12607,N_12561,N_12583);
or U12608 (N_12608,N_12543,N_12508);
and U12609 (N_12609,N_12577,N_12514);
or U12610 (N_12610,N_12598,N_12525);
nand U12611 (N_12611,N_12503,N_12556);
and U12612 (N_12612,N_12570,N_12581);
and U12613 (N_12613,N_12428,N_12496);
nor U12614 (N_12614,N_12476,N_12578);
nor U12615 (N_12615,N_12575,N_12462);
nor U12616 (N_12616,N_12405,N_12491);
and U12617 (N_12617,N_12432,N_12574);
xor U12618 (N_12618,N_12419,N_12544);
nor U12619 (N_12619,N_12564,N_12468);
nand U12620 (N_12620,N_12499,N_12490);
or U12621 (N_12621,N_12426,N_12584);
and U12622 (N_12622,N_12569,N_12459);
nand U12623 (N_12623,N_12533,N_12545);
xor U12624 (N_12624,N_12589,N_12454);
nor U12625 (N_12625,N_12492,N_12591);
nor U12626 (N_12626,N_12495,N_12524);
or U12627 (N_12627,N_12481,N_12560);
or U12628 (N_12628,N_12504,N_12507);
or U12629 (N_12629,N_12415,N_12472);
or U12630 (N_12630,N_12412,N_12439);
nor U12631 (N_12631,N_12500,N_12450);
or U12632 (N_12632,N_12517,N_12537);
nor U12633 (N_12633,N_12538,N_12562);
and U12634 (N_12634,N_12400,N_12567);
nand U12635 (N_12635,N_12518,N_12565);
and U12636 (N_12636,N_12484,N_12505);
or U12637 (N_12637,N_12557,N_12451);
xor U12638 (N_12638,N_12532,N_12528);
and U12639 (N_12639,N_12407,N_12527);
and U12640 (N_12640,N_12485,N_12573);
xnor U12641 (N_12641,N_12547,N_12494);
or U12642 (N_12642,N_12555,N_12506);
xor U12643 (N_12643,N_12471,N_12596);
or U12644 (N_12644,N_12582,N_12430);
and U12645 (N_12645,N_12420,N_12449);
and U12646 (N_12646,N_12438,N_12452);
nand U12647 (N_12647,N_12572,N_12440);
or U12648 (N_12648,N_12477,N_12534);
and U12649 (N_12649,N_12559,N_12435);
nand U12650 (N_12650,N_12408,N_12447);
xnor U12651 (N_12651,N_12502,N_12425);
or U12652 (N_12652,N_12523,N_12409);
or U12653 (N_12653,N_12474,N_12592);
nand U12654 (N_12654,N_12480,N_12458);
nor U12655 (N_12655,N_12553,N_12585);
and U12656 (N_12656,N_12571,N_12483);
xnor U12657 (N_12657,N_12486,N_12469);
and U12658 (N_12658,N_12539,N_12501);
nand U12659 (N_12659,N_12512,N_12576);
nor U12660 (N_12660,N_12457,N_12411);
and U12661 (N_12661,N_12551,N_12593);
and U12662 (N_12662,N_12563,N_12437);
or U12663 (N_12663,N_12519,N_12414);
and U12664 (N_12664,N_12590,N_12548);
nor U12665 (N_12665,N_12417,N_12406);
or U12666 (N_12666,N_12442,N_12586);
nand U12667 (N_12667,N_12554,N_12515);
or U12668 (N_12668,N_12463,N_12464);
xnor U12669 (N_12669,N_12410,N_12433);
nand U12670 (N_12670,N_12448,N_12588);
and U12671 (N_12671,N_12421,N_12510);
or U12672 (N_12672,N_12436,N_12429);
nand U12673 (N_12673,N_12482,N_12424);
nand U12674 (N_12674,N_12418,N_12441);
and U12675 (N_12675,N_12509,N_12456);
and U12676 (N_12676,N_12540,N_12530);
and U12677 (N_12677,N_12493,N_12558);
and U12678 (N_12678,N_12536,N_12526);
nor U12679 (N_12679,N_12541,N_12542);
nor U12680 (N_12680,N_12529,N_12434);
or U12681 (N_12681,N_12535,N_12473);
nand U12682 (N_12682,N_12453,N_12401);
nand U12683 (N_12683,N_12594,N_12489);
nand U12684 (N_12684,N_12566,N_12479);
nand U12685 (N_12685,N_12595,N_12522);
nor U12686 (N_12686,N_12404,N_12467);
xnor U12687 (N_12687,N_12446,N_12478);
xnor U12688 (N_12688,N_12497,N_12513);
nor U12689 (N_12689,N_12455,N_12549);
nand U12690 (N_12690,N_12531,N_12431);
xnor U12691 (N_12691,N_12422,N_12443);
or U12692 (N_12692,N_12465,N_12413);
or U12693 (N_12693,N_12416,N_12568);
xnor U12694 (N_12694,N_12460,N_12470);
nand U12695 (N_12695,N_12546,N_12487);
and U12696 (N_12696,N_12521,N_12511);
and U12697 (N_12697,N_12444,N_12579);
nand U12698 (N_12698,N_12423,N_12445);
nand U12699 (N_12699,N_12461,N_12403);
nor U12700 (N_12700,N_12524,N_12571);
or U12701 (N_12701,N_12555,N_12493);
nor U12702 (N_12702,N_12454,N_12490);
and U12703 (N_12703,N_12576,N_12525);
nand U12704 (N_12704,N_12465,N_12532);
and U12705 (N_12705,N_12596,N_12571);
xnor U12706 (N_12706,N_12538,N_12461);
nand U12707 (N_12707,N_12428,N_12506);
or U12708 (N_12708,N_12445,N_12480);
xor U12709 (N_12709,N_12409,N_12559);
or U12710 (N_12710,N_12566,N_12436);
and U12711 (N_12711,N_12500,N_12599);
nand U12712 (N_12712,N_12518,N_12590);
nand U12713 (N_12713,N_12588,N_12485);
xnor U12714 (N_12714,N_12508,N_12563);
nor U12715 (N_12715,N_12411,N_12482);
and U12716 (N_12716,N_12480,N_12451);
or U12717 (N_12717,N_12558,N_12582);
nand U12718 (N_12718,N_12453,N_12491);
nor U12719 (N_12719,N_12415,N_12559);
xor U12720 (N_12720,N_12535,N_12520);
nor U12721 (N_12721,N_12401,N_12599);
or U12722 (N_12722,N_12543,N_12460);
and U12723 (N_12723,N_12471,N_12538);
and U12724 (N_12724,N_12496,N_12575);
or U12725 (N_12725,N_12503,N_12509);
xor U12726 (N_12726,N_12563,N_12435);
nor U12727 (N_12727,N_12511,N_12551);
or U12728 (N_12728,N_12537,N_12528);
or U12729 (N_12729,N_12549,N_12470);
or U12730 (N_12730,N_12478,N_12442);
xnor U12731 (N_12731,N_12421,N_12453);
nand U12732 (N_12732,N_12481,N_12592);
and U12733 (N_12733,N_12582,N_12474);
nand U12734 (N_12734,N_12550,N_12434);
nor U12735 (N_12735,N_12493,N_12538);
and U12736 (N_12736,N_12440,N_12590);
or U12737 (N_12737,N_12580,N_12591);
and U12738 (N_12738,N_12562,N_12542);
or U12739 (N_12739,N_12436,N_12571);
nand U12740 (N_12740,N_12528,N_12429);
and U12741 (N_12741,N_12564,N_12488);
nand U12742 (N_12742,N_12427,N_12472);
xnor U12743 (N_12743,N_12562,N_12470);
nand U12744 (N_12744,N_12513,N_12450);
and U12745 (N_12745,N_12442,N_12441);
nand U12746 (N_12746,N_12404,N_12407);
and U12747 (N_12747,N_12537,N_12589);
or U12748 (N_12748,N_12574,N_12462);
nand U12749 (N_12749,N_12596,N_12470);
nand U12750 (N_12750,N_12556,N_12530);
and U12751 (N_12751,N_12519,N_12582);
nor U12752 (N_12752,N_12450,N_12464);
nand U12753 (N_12753,N_12421,N_12476);
nor U12754 (N_12754,N_12564,N_12546);
or U12755 (N_12755,N_12432,N_12572);
nor U12756 (N_12756,N_12559,N_12597);
nor U12757 (N_12757,N_12564,N_12429);
nor U12758 (N_12758,N_12528,N_12502);
xnor U12759 (N_12759,N_12508,N_12545);
xor U12760 (N_12760,N_12431,N_12447);
xor U12761 (N_12761,N_12476,N_12471);
and U12762 (N_12762,N_12479,N_12492);
or U12763 (N_12763,N_12484,N_12593);
or U12764 (N_12764,N_12561,N_12492);
or U12765 (N_12765,N_12470,N_12453);
nor U12766 (N_12766,N_12495,N_12522);
and U12767 (N_12767,N_12401,N_12569);
xor U12768 (N_12768,N_12501,N_12591);
xnor U12769 (N_12769,N_12566,N_12401);
nor U12770 (N_12770,N_12454,N_12562);
nor U12771 (N_12771,N_12446,N_12439);
and U12772 (N_12772,N_12482,N_12573);
nor U12773 (N_12773,N_12545,N_12479);
and U12774 (N_12774,N_12481,N_12464);
and U12775 (N_12775,N_12512,N_12413);
xor U12776 (N_12776,N_12458,N_12451);
or U12777 (N_12777,N_12455,N_12566);
or U12778 (N_12778,N_12424,N_12400);
nand U12779 (N_12779,N_12598,N_12559);
or U12780 (N_12780,N_12576,N_12521);
xor U12781 (N_12781,N_12597,N_12528);
nor U12782 (N_12782,N_12574,N_12431);
or U12783 (N_12783,N_12526,N_12550);
nand U12784 (N_12784,N_12548,N_12445);
and U12785 (N_12785,N_12516,N_12563);
or U12786 (N_12786,N_12451,N_12503);
or U12787 (N_12787,N_12471,N_12464);
xnor U12788 (N_12788,N_12596,N_12508);
nand U12789 (N_12789,N_12430,N_12470);
xor U12790 (N_12790,N_12483,N_12554);
xor U12791 (N_12791,N_12487,N_12580);
and U12792 (N_12792,N_12453,N_12528);
nand U12793 (N_12793,N_12533,N_12569);
xnor U12794 (N_12794,N_12522,N_12535);
xnor U12795 (N_12795,N_12514,N_12594);
xnor U12796 (N_12796,N_12575,N_12550);
and U12797 (N_12797,N_12585,N_12549);
xor U12798 (N_12798,N_12564,N_12545);
or U12799 (N_12799,N_12430,N_12531);
nor U12800 (N_12800,N_12704,N_12796);
nand U12801 (N_12801,N_12724,N_12606);
and U12802 (N_12802,N_12797,N_12771);
nor U12803 (N_12803,N_12696,N_12748);
xor U12804 (N_12804,N_12607,N_12756);
or U12805 (N_12805,N_12776,N_12755);
nor U12806 (N_12806,N_12778,N_12643);
or U12807 (N_12807,N_12630,N_12705);
nand U12808 (N_12808,N_12626,N_12785);
xnor U12809 (N_12809,N_12799,N_12651);
xnor U12810 (N_12810,N_12689,N_12760);
and U12811 (N_12811,N_12610,N_12775);
xnor U12812 (N_12812,N_12611,N_12660);
or U12813 (N_12813,N_12763,N_12674);
nand U12814 (N_12814,N_12642,N_12620);
xor U12815 (N_12815,N_12625,N_12730);
and U12816 (N_12816,N_12713,N_12740);
and U12817 (N_12817,N_12698,N_12742);
nor U12818 (N_12818,N_12703,N_12744);
or U12819 (N_12819,N_12602,N_12685);
nand U12820 (N_12820,N_12684,N_12735);
or U12821 (N_12821,N_12693,N_12787);
nand U12822 (N_12822,N_12732,N_12757);
or U12823 (N_12823,N_12690,N_12792);
xnor U12824 (N_12824,N_12627,N_12761);
or U12825 (N_12825,N_12728,N_12741);
nand U12826 (N_12826,N_12769,N_12609);
xor U12827 (N_12827,N_12716,N_12672);
xor U12828 (N_12828,N_12657,N_12798);
or U12829 (N_12829,N_12782,N_12681);
xnor U12830 (N_12830,N_12658,N_12750);
or U12831 (N_12831,N_12665,N_12624);
xnor U12832 (N_12832,N_12720,N_12712);
nand U12833 (N_12833,N_12613,N_12746);
xor U12834 (N_12834,N_12634,N_12633);
nor U12835 (N_12835,N_12726,N_12710);
and U12836 (N_12836,N_12723,N_12622);
xnor U12837 (N_12837,N_12668,N_12675);
nor U12838 (N_12838,N_12608,N_12768);
nor U12839 (N_12839,N_12629,N_12733);
and U12840 (N_12840,N_12667,N_12784);
and U12841 (N_12841,N_12781,N_12641);
xnor U12842 (N_12842,N_12673,N_12765);
nor U12843 (N_12843,N_12789,N_12655);
and U12844 (N_12844,N_12745,N_12767);
or U12845 (N_12845,N_12692,N_12709);
nand U12846 (N_12846,N_12715,N_12734);
nand U12847 (N_12847,N_12718,N_12616);
xnor U12848 (N_12848,N_12650,N_12614);
xor U12849 (N_12849,N_12680,N_12795);
xor U12850 (N_12850,N_12679,N_12671);
and U12851 (N_12851,N_12661,N_12682);
nand U12852 (N_12852,N_12707,N_12688);
nand U12853 (N_12853,N_12749,N_12617);
nand U12854 (N_12854,N_12612,N_12640);
xnor U12855 (N_12855,N_12645,N_12773);
xor U12856 (N_12856,N_12722,N_12751);
xor U12857 (N_12857,N_12697,N_12701);
and U12858 (N_12858,N_12636,N_12619);
and U12859 (N_12859,N_12621,N_12666);
or U12860 (N_12860,N_12662,N_12711);
nor U12861 (N_12861,N_12601,N_12646);
and U12862 (N_12862,N_12779,N_12649);
and U12863 (N_12863,N_12780,N_12714);
xor U12864 (N_12864,N_12793,N_12706);
nor U12865 (N_12865,N_12727,N_12752);
and U12866 (N_12866,N_12632,N_12788);
xnor U12867 (N_12867,N_12729,N_12770);
nor U12868 (N_12868,N_12754,N_12638);
nor U12869 (N_12869,N_12717,N_12637);
and U12870 (N_12870,N_12766,N_12694);
nor U12871 (N_12871,N_12708,N_12623);
and U12872 (N_12872,N_12656,N_12631);
xor U12873 (N_12873,N_12639,N_12753);
and U12874 (N_12874,N_12615,N_12794);
nand U12875 (N_12875,N_12603,N_12791);
or U12876 (N_12876,N_12669,N_12683);
nand U12877 (N_12877,N_12758,N_12725);
or U12878 (N_12878,N_12764,N_12652);
and U12879 (N_12879,N_12663,N_12686);
and U12880 (N_12880,N_12654,N_12777);
or U12881 (N_12881,N_12635,N_12600);
nand U12882 (N_12882,N_12731,N_12628);
and U12883 (N_12883,N_12772,N_12790);
or U12884 (N_12884,N_12605,N_12774);
xnor U12885 (N_12885,N_12783,N_12699);
xor U12886 (N_12886,N_12678,N_12691);
xor U12887 (N_12887,N_12700,N_12687);
or U12888 (N_12888,N_12647,N_12743);
and U12889 (N_12889,N_12664,N_12719);
or U12890 (N_12890,N_12644,N_12702);
and U12891 (N_12891,N_12659,N_12676);
xnor U12892 (N_12892,N_12653,N_12721);
or U12893 (N_12893,N_12747,N_12604);
nor U12894 (N_12894,N_12737,N_12677);
nor U12895 (N_12895,N_12759,N_12618);
xnor U12896 (N_12896,N_12739,N_12762);
or U12897 (N_12897,N_12786,N_12736);
or U12898 (N_12898,N_12738,N_12648);
or U12899 (N_12899,N_12695,N_12670);
nor U12900 (N_12900,N_12711,N_12704);
and U12901 (N_12901,N_12623,N_12651);
xnor U12902 (N_12902,N_12783,N_12720);
and U12903 (N_12903,N_12728,N_12796);
nor U12904 (N_12904,N_12727,N_12683);
xor U12905 (N_12905,N_12672,N_12751);
or U12906 (N_12906,N_12622,N_12789);
nor U12907 (N_12907,N_12636,N_12760);
or U12908 (N_12908,N_12731,N_12659);
nand U12909 (N_12909,N_12639,N_12657);
nor U12910 (N_12910,N_12647,N_12769);
nor U12911 (N_12911,N_12682,N_12770);
or U12912 (N_12912,N_12639,N_12625);
nor U12913 (N_12913,N_12672,N_12728);
and U12914 (N_12914,N_12693,N_12706);
and U12915 (N_12915,N_12627,N_12690);
and U12916 (N_12916,N_12708,N_12710);
nand U12917 (N_12917,N_12670,N_12747);
or U12918 (N_12918,N_12757,N_12685);
and U12919 (N_12919,N_12687,N_12704);
xnor U12920 (N_12920,N_12639,N_12701);
nand U12921 (N_12921,N_12745,N_12657);
xnor U12922 (N_12922,N_12699,N_12672);
nor U12923 (N_12923,N_12684,N_12783);
nand U12924 (N_12924,N_12623,N_12664);
nand U12925 (N_12925,N_12748,N_12775);
xor U12926 (N_12926,N_12763,N_12656);
or U12927 (N_12927,N_12786,N_12612);
and U12928 (N_12928,N_12684,N_12600);
nand U12929 (N_12929,N_12726,N_12687);
xnor U12930 (N_12930,N_12684,N_12656);
xnor U12931 (N_12931,N_12675,N_12677);
xor U12932 (N_12932,N_12694,N_12683);
xnor U12933 (N_12933,N_12795,N_12652);
and U12934 (N_12934,N_12719,N_12786);
nand U12935 (N_12935,N_12623,N_12746);
and U12936 (N_12936,N_12796,N_12712);
or U12937 (N_12937,N_12790,N_12664);
xnor U12938 (N_12938,N_12601,N_12659);
nand U12939 (N_12939,N_12729,N_12683);
or U12940 (N_12940,N_12615,N_12702);
nand U12941 (N_12941,N_12627,N_12718);
nor U12942 (N_12942,N_12692,N_12681);
nor U12943 (N_12943,N_12623,N_12710);
nand U12944 (N_12944,N_12795,N_12610);
xor U12945 (N_12945,N_12750,N_12713);
nand U12946 (N_12946,N_12676,N_12686);
and U12947 (N_12947,N_12768,N_12711);
or U12948 (N_12948,N_12759,N_12626);
nand U12949 (N_12949,N_12601,N_12784);
nor U12950 (N_12950,N_12645,N_12670);
nor U12951 (N_12951,N_12663,N_12693);
nand U12952 (N_12952,N_12768,N_12688);
nor U12953 (N_12953,N_12661,N_12608);
and U12954 (N_12954,N_12773,N_12633);
nand U12955 (N_12955,N_12773,N_12607);
or U12956 (N_12956,N_12793,N_12676);
nand U12957 (N_12957,N_12607,N_12617);
nor U12958 (N_12958,N_12619,N_12755);
or U12959 (N_12959,N_12633,N_12770);
xnor U12960 (N_12960,N_12730,N_12654);
nor U12961 (N_12961,N_12799,N_12603);
nor U12962 (N_12962,N_12752,N_12655);
nor U12963 (N_12963,N_12620,N_12732);
nand U12964 (N_12964,N_12665,N_12768);
and U12965 (N_12965,N_12764,N_12785);
xor U12966 (N_12966,N_12713,N_12766);
or U12967 (N_12967,N_12726,N_12640);
nand U12968 (N_12968,N_12743,N_12796);
xnor U12969 (N_12969,N_12711,N_12608);
xor U12970 (N_12970,N_12618,N_12653);
and U12971 (N_12971,N_12666,N_12792);
nor U12972 (N_12972,N_12730,N_12708);
nor U12973 (N_12973,N_12675,N_12700);
nor U12974 (N_12974,N_12656,N_12665);
or U12975 (N_12975,N_12625,N_12670);
or U12976 (N_12976,N_12700,N_12614);
nor U12977 (N_12977,N_12652,N_12634);
and U12978 (N_12978,N_12655,N_12609);
or U12979 (N_12979,N_12616,N_12765);
or U12980 (N_12980,N_12703,N_12631);
nor U12981 (N_12981,N_12643,N_12708);
nand U12982 (N_12982,N_12748,N_12626);
or U12983 (N_12983,N_12765,N_12763);
nor U12984 (N_12984,N_12628,N_12784);
and U12985 (N_12985,N_12759,N_12610);
xor U12986 (N_12986,N_12781,N_12666);
xor U12987 (N_12987,N_12739,N_12773);
nor U12988 (N_12988,N_12623,N_12771);
nand U12989 (N_12989,N_12750,N_12759);
and U12990 (N_12990,N_12656,N_12774);
or U12991 (N_12991,N_12613,N_12761);
nor U12992 (N_12992,N_12749,N_12767);
nand U12993 (N_12993,N_12667,N_12654);
or U12994 (N_12994,N_12638,N_12712);
or U12995 (N_12995,N_12725,N_12770);
and U12996 (N_12996,N_12749,N_12784);
xnor U12997 (N_12997,N_12783,N_12765);
or U12998 (N_12998,N_12671,N_12690);
nor U12999 (N_12999,N_12770,N_12688);
and U13000 (N_13000,N_12997,N_12869);
or U13001 (N_13001,N_12870,N_12961);
xor U13002 (N_13002,N_12847,N_12827);
or U13003 (N_13003,N_12916,N_12861);
nor U13004 (N_13004,N_12824,N_12834);
xor U13005 (N_13005,N_12936,N_12904);
and U13006 (N_13006,N_12971,N_12866);
nand U13007 (N_13007,N_12977,N_12946);
nand U13008 (N_13008,N_12811,N_12800);
and U13009 (N_13009,N_12966,N_12846);
nand U13010 (N_13010,N_12973,N_12844);
nand U13011 (N_13011,N_12828,N_12945);
or U13012 (N_13012,N_12931,N_12823);
nor U13013 (N_13013,N_12801,N_12963);
xor U13014 (N_13014,N_12804,N_12842);
nor U13015 (N_13015,N_12814,N_12981);
nor U13016 (N_13016,N_12809,N_12886);
or U13017 (N_13017,N_12903,N_12968);
nand U13018 (N_13018,N_12893,N_12805);
nor U13019 (N_13019,N_12980,N_12826);
and U13020 (N_13020,N_12972,N_12984);
nor U13021 (N_13021,N_12864,N_12908);
nor U13022 (N_13022,N_12987,N_12881);
and U13023 (N_13023,N_12999,N_12810);
nor U13024 (N_13024,N_12806,N_12924);
or U13025 (N_13025,N_12982,N_12803);
nor U13026 (N_13026,N_12871,N_12979);
nor U13027 (N_13027,N_12992,N_12854);
and U13028 (N_13028,N_12900,N_12888);
nand U13029 (N_13029,N_12911,N_12874);
or U13030 (N_13030,N_12855,N_12856);
and U13031 (N_13031,N_12901,N_12905);
or U13032 (N_13032,N_12892,N_12944);
nand U13033 (N_13033,N_12849,N_12995);
nand U13034 (N_13034,N_12830,N_12899);
nand U13035 (N_13035,N_12959,N_12816);
and U13036 (N_13036,N_12838,N_12843);
xor U13037 (N_13037,N_12906,N_12942);
nand U13038 (N_13038,N_12990,N_12926);
or U13039 (N_13039,N_12952,N_12928);
and U13040 (N_13040,N_12807,N_12833);
nand U13041 (N_13041,N_12913,N_12851);
nand U13042 (N_13042,N_12878,N_12895);
or U13043 (N_13043,N_12853,N_12820);
or U13044 (N_13044,N_12883,N_12859);
xor U13045 (N_13045,N_12836,N_12994);
nand U13046 (N_13046,N_12934,N_12974);
and U13047 (N_13047,N_12957,N_12884);
or U13048 (N_13048,N_12887,N_12907);
xor U13049 (N_13049,N_12955,N_12812);
nand U13050 (N_13050,N_12967,N_12845);
or U13051 (N_13051,N_12919,N_12872);
or U13052 (N_13052,N_12948,N_12839);
or U13053 (N_13053,N_12896,N_12985);
and U13054 (N_13054,N_12929,N_12868);
nor U13055 (N_13055,N_12815,N_12802);
or U13056 (N_13056,N_12993,N_12909);
nand U13057 (N_13057,N_12852,N_12947);
and U13058 (N_13058,N_12876,N_12922);
xor U13059 (N_13059,N_12848,N_12877);
nand U13060 (N_13060,N_12943,N_12954);
and U13061 (N_13061,N_12923,N_12910);
nor U13062 (N_13062,N_12912,N_12817);
nand U13063 (N_13063,N_12858,N_12920);
and U13064 (N_13064,N_12918,N_12988);
nand U13065 (N_13065,N_12937,N_12965);
nand U13066 (N_13066,N_12950,N_12819);
or U13067 (N_13067,N_12841,N_12879);
and U13068 (N_13068,N_12921,N_12989);
or U13069 (N_13069,N_12850,N_12986);
xor U13070 (N_13070,N_12970,N_12835);
or U13071 (N_13071,N_12960,N_12938);
nor U13072 (N_13072,N_12953,N_12880);
nand U13073 (N_13073,N_12831,N_12840);
nand U13074 (N_13074,N_12894,N_12935);
nor U13075 (N_13075,N_12939,N_12885);
xnor U13076 (N_13076,N_12962,N_12951);
and U13077 (N_13077,N_12821,N_12991);
and U13078 (N_13078,N_12832,N_12873);
and U13079 (N_13079,N_12857,N_12818);
and U13080 (N_13080,N_12933,N_12829);
nor U13081 (N_13081,N_12976,N_12808);
or U13082 (N_13082,N_12925,N_12964);
xnor U13083 (N_13083,N_12975,N_12956);
or U13084 (N_13084,N_12915,N_12890);
xnor U13085 (N_13085,N_12958,N_12825);
xnor U13086 (N_13086,N_12978,N_12996);
and U13087 (N_13087,N_12875,N_12940);
nand U13088 (N_13088,N_12897,N_12983);
and U13089 (N_13089,N_12932,N_12863);
or U13090 (N_13090,N_12914,N_12927);
nand U13091 (N_13091,N_12969,N_12889);
or U13092 (N_13092,N_12867,N_12917);
and U13093 (N_13093,N_12860,N_12930);
or U13094 (N_13094,N_12837,N_12813);
and U13095 (N_13095,N_12862,N_12865);
xnor U13096 (N_13096,N_12949,N_12891);
or U13097 (N_13097,N_12882,N_12822);
nand U13098 (N_13098,N_12941,N_12998);
and U13099 (N_13099,N_12902,N_12898);
xnor U13100 (N_13100,N_12889,N_12847);
and U13101 (N_13101,N_12843,N_12847);
nand U13102 (N_13102,N_12972,N_12930);
nand U13103 (N_13103,N_12831,N_12936);
xnor U13104 (N_13104,N_12806,N_12822);
xor U13105 (N_13105,N_12959,N_12802);
and U13106 (N_13106,N_12933,N_12954);
nand U13107 (N_13107,N_12820,N_12856);
xnor U13108 (N_13108,N_12991,N_12814);
and U13109 (N_13109,N_12990,N_12979);
and U13110 (N_13110,N_12827,N_12819);
nor U13111 (N_13111,N_12965,N_12802);
xor U13112 (N_13112,N_12947,N_12893);
and U13113 (N_13113,N_12918,N_12972);
or U13114 (N_13114,N_12842,N_12880);
or U13115 (N_13115,N_12875,N_12812);
nor U13116 (N_13116,N_12806,N_12953);
nand U13117 (N_13117,N_12971,N_12973);
and U13118 (N_13118,N_12842,N_12853);
nor U13119 (N_13119,N_12916,N_12960);
nor U13120 (N_13120,N_12974,N_12815);
and U13121 (N_13121,N_12996,N_12972);
nor U13122 (N_13122,N_12945,N_12814);
nor U13123 (N_13123,N_12996,N_12881);
or U13124 (N_13124,N_12994,N_12972);
and U13125 (N_13125,N_12822,N_12812);
xnor U13126 (N_13126,N_12828,N_12938);
xor U13127 (N_13127,N_12813,N_12905);
nand U13128 (N_13128,N_12971,N_12978);
or U13129 (N_13129,N_12991,N_12837);
xor U13130 (N_13130,N_12933,N_12893);
and U13131 (N_13131,N_12846,N_12891);
nor U13132 (N_13132,N_12915,N_12877);
and U13133 (N_13133,N_12962,N_12821);
and U13134 (N_13134,N_12963,N_12885);
nor U13135 (N_13135,N_12834,N_12823);
nand U13136 (N_13136,N_12874,N_12883);
and U13137 (N_13137,N_12992,N_12845);
xor U13138 (N_13138,N_12824,N_12937);
xor U13139 (N_13139,N_12882,N_12888);
nor U13140 (N_13140,N_12937,N_12924);
nand U13141 (N_13141,N_12960,N_12918);
xor U13142 (N_13142,N_12959,N_12844);
xnor U13143 (N_13143,N_12956,N_12974);
nand U13144 (N_13144,N_12898,N_12964);
nor U13145 (N_13145,N_12831,N_12869);
nand U13146 (N_13146,N_12886,N_12949);
and U13147 (N_13147,N_12826,N_12979);
or U13148 (N_13148,N_12858,N_12950);
and U13149 (N_13149,N_12919,N_12840);
xor U13150 (N_13150,N_12983,N_12989);
xor U13151 (N_13151,N_12872,N_12957);
nand U13152 (N_13152,N_12912,N_12922);
or U13153 (N_13153,N_12908,N_12951);
and U13154 (N_13154,N_12813,N_12861);
xor U13155 (N_13155,N_12813,N_12887);
and U13156 (N_13156,N_12800,N_12882);
nand U13157 (N_13157,N_12905,N_12828);
and U13158 (N_13158,N_12916,N_12869);
nand U13159 (N_13159,N_12824,N_12961);
and U13160 (N_13160,N_12884,N_12966);
and U13161 (N_13161,N_12892,N_12912);
xor U13162 (N_13162,N_12980,N_12862);
or U13163 (N_13163,N_12910,N_12936);
and U13164 (N_13164,N_12928,N_12990);
or U13165 (N_13165,N_12851,N_12964);
nor U13166 (N_13166,N_12806,N_12849);
and U13167 (N_13167,N_12923,N_12848);
nand U13168 (N_13168,N_12904,N_12837);
nand U13169 (N_13169,N_12853,N_12843);
nor U13170 (N_13170,N_12944,N_12917);
nand U13171 (N_13171,N_12861,N_12918);
nand U13172 (N_13172,N_12989,N_12869);
and U13173 (N_13173,N_12841,N_12886);
xnor U13174 (N_13174,N_12820,N_12850);
and U13175 (N_13175,N_12929,N_12915);
or U13176 (N_13176,N_12993,N_12873);
nand U13177 (N_13177,N_12917,N_12965);
or U13178 (N_13178,N_12832,N_12820);
xnor U13179 (N_13179,N_12826,N_12861);
xor U13180 (N_13180,N_12959,N_12941);
or U13181 (N_13181,N_12867,N_12878);
or U13182 (N_13182,N_12930,N_12878);
nand U13183 (N_13183,N_12993,N_12862);
or U13184 (N_13184,N_12936,N_12886);
nor U13185 (N_13185,N_12999,N_12965);
xor U13186 (N_13186,N_12906,N_12875);
xor U13187 (N_13187,N_12946,N_12965);
and U13188 (N_13188,N_12861,N_12808);
or U13189 (N_13189,N_12816,N_12829);
or U13190 (N_13190,N_12832,N_12996);
xor U13191 (N_13191,N_12879,N_12872);
xor U13192 (N_13192,N_12961,N_12839);
nand U13193 (N_13193,N_12897,N_12900);
nor U13194 (N_13194,N_12893,N_12925);
nor U13195 (N_13195,N_12996,N_12903);
and U13196 (N_13196,N_12809,N_12814);
xor U13197 (N_13197,N_12805,N_12878);
and U13198 (N_13198,N_12913,N_12942);
and U13199 (N_13199,N_12962,N_12830);
nor U13200 (N_13200,N_13116,N_13145);
nand U13201 (N_13201,N_13037,N_13086);
nor U13202 (N_13202,N_13061,N_13074);
or U13203 (N_13203,N_13080,N_13165);
or U13204 (N_13204,N_13129,N_13007);
nor U13205 (N_13205,N_13142,N_13054);
nor U13206 (N_13206,N_13015,N_13112);
and U13207 (N_13207,N_13032,N_13174);
xor U13208 (N_13208,N_13069,N_13192);
nand U13209 (N_13209,N_13191,N_13138);
or U13210 (N_13210,N_13095,N_13081);
or U13211 (N_13211,N_13092,N_13177);
nor U13212 (N_13212,N_13034,N_13001);
and U13213 (N_13213,N_13070,N_13144);
nand U13214 (N_13214,N_13068,N_13194);
or U13215 (N_13215,N_13052,N_13183);
xnor U13216 (N_13216,N_13009,N_13022);
or U13217 (N_13217,N_13172,N_13004);
xnor U13218 (N_13218,N_13023,N_13018);
nor U13219 (N_13219,N_13132,N_13136);
or U13220 (N_13220,N_13135,N_13100);
nand U13221 (N_13221,N_13117,N_13053);
nand U13222 (N_13222,N_13083,N_13180);
or U13223 (N_13223,N_13048,N_13137);
xnor U13224 (N_13224,N_13064,N_13171);
nand U13225 (N_13225,N_13079,N_13058);
nor U13226 (N_13226,N_13012,N_13031);
nor U13227 (N_13227,N_13188,N_13168);
nand U13228 (N_13228,N_13161,N_13005);
and U13229 (N_13229,N_13152,N_13186);
and U13230 (N_13230,N_13041,N_13082);
nor U13231 (N_13231,N_13110,N_13140);
or U13232 (N_13232,N_13159,N_13045);
nand U13233 (N_13233,N_13000,N_13028);
and U13234 (N_13234,N_13077,N_13162);
nand U13235 (N_13235,N_13169,N_13121);
or U13236 (N_13236,N_13065,N_13198);
nand U13237 (N_13237,N_13067,N_13043);
nor U13238 (N_13238,N_13049,N_13050);
or U13239 (N_13239,N_13127,N_13099);
or U13240 (N_13240,N_13063,N_13090);
or U13241 (N_13241,N_13170,N_13109);
nand U13242 (N_13242,N_13150,N_13060);
and U13243 (N_13243,N_13057,N_13184);
and U13244 (N_13244,N_13014,N_13185);
and U13245 (N_13245,N_13098,N_13062);
xnor U13246 (N_13246,N_13003,N_13181);
nand U13247 (N_13247,N_13106,N_13118);
and U13248 (N_13248,N_13055,N_13143);
and U13249 (N_13249,N_13024,N_13056);
nor U13250 (N_13250,N_13088,N_13036);
or U13251 (N_13251,N_13097,N_13124);
or U13252 (N_13252,N_13158,N_13094);
nand U13253 (N_13253,N_13073,N_13167);
xor U13254 (N_13254,N_13101,N_13146);
and U13255 (N_13255,N_13017,N_13075);
and U13256 (N_13256,N_13039,N_13008);
xnor U13257 (N_13257,N_13160,N_13016);
or U13258 (N_13258,N_13153,N_13115);
xnor U13259 (N_13259,N_13038,N_13199);
and U13260 (N_13260,N_13130,N_13087);
nand U13261 (N_13261,N_13104,N_13187);
nand U13262 (N_13262,N_13030,N_13126);
xor U13263 (N_13263,N_13119,N_13076);
xnor U13264 (N_13264,N_13020,N_13006);
xnor U13265 (N_13265,N_13078,N_13021);
nor U13266 (N_13266,N_13047,N_13046);
or U13267 (N_13267,N_13147,N_13071);
nand U13268 (N_13268,N_13084,N_13089);
nor U13269 (N_13269,N_13085,N_13033);
or U13270 (N_13270,N_13131,N_13107);
nand U13271 (N_13271,N_13040,N_13011);
nand U13272 (N_13272,N_13190,N_13042);
nand U13273 (N_13273,N_13163,N_13013);
and U13274 (N_13274,N_13103,N_13113);
nand U13275 (N_13275,N_13066,N_13179);
or U13276 (N_13276,N_13134,N_13141);
or U13277 (N_13277,N_13108,N_13010);
or U13278 (N_13278,N_13051,N_13133);
nor U13279 (N_13279,N_13157,N_13193);
or U13280 (N_13280,N_13125,N_13019);
xor U13281 (N_13281,N_13105,N_13197);
nor U13282 (N_13282,N_13026,N_13128);
nor U13283 (N_13283,N_13072,N_13155);
xnor U13284 (N_13284,N_13151,N_13120);
nor U13285 (N_13285,N_13027,N_13164);
or U13286 (N_13286,N_13122,N_13196);
and U13287 (N_13287,N_13148,N_13029);
nand U13288 (N_13288,N_13182,N_13166);
or U13289 (N_13289,N_13096,N_13189);
or U13290 (N_13290,N_13123,N_13156);
and U13291 (N_13291,N_13035,N_13044);
or U13292 (N_13292,N_13102,N_13139);
nor U13293 (N_13293,N_13176,N_13173);
and U13294 (N_13294,N_13154,N_13114);
nor U13295 (N_13295,N_13002,N_13149);
or U13296 (N_13296,N_13111,N_13093);
and U13297 (N_13297,N_13195,N_13091);
or U13298 (N_13298,N_13059,N_13175);
xnor U13299 (N_13299,N_13025,N_13178);
nand U13300 (N_13300,N_13068,N_13069);
or U13301 (N_13301,N_13071,N_13054);
xnor U13302 (N_13302,N_13006,N_13026);
xor U13303 (N_13303,N_13148,N_13007);
nand U13304 (N_13304,N_13091,N_13051);
nand U13305 (N_13305,N_13123,N_13069);
nor U13306 (N_13306,N_13077,N_13015);
nor U13307 (N_13307,N_13003,N_13023);
and U13308 (N_13308,N_13149,N_13043);
nand U13309 (N_13309,N_13076,N_13083);
and U13310 (N_13310,N_13059,N_13196);
and U13311 (N_13311,N_13118,N_13071);
nor U13312 (N_13312,N_13001,N_13108);
or U13313 (N_13313,N_13079,N_13174);
xnor U13314 (N_13314,N_13062,N_13165);
or U13315 (N_13315,N_13107,N_13166);
or U13316 (N_13316,N_13045,N_13077);
nand U13317 (N_13317,N_13152,N_13164);
or U13318 (N_13318,N_13096,N_13039);
nand U13319 (N_13319,N_13078,N_13112);
or U13320 (N_13320,N_13175,N_13067);
nand U13321 (N_13321,N_13087,N_13117);
or U13322 (N_13322,N_13033,N_13002);
nor U13323 (N_13323,N_13055,N_13038);
nor U13324 (N_13324,N_13009,N_13068);
nand U13325 (N_13325,N_13005,N_13001);
and U13326 (N_13326,N_13130,N_13006);
or U13327 (N_13327,N_13197,N_13025);
nor U13328 (N_13328,N_13075,N_13003);
nor U13329 (N_13329,N_13113,N_13127);
or U13330 (N_13330,N_13172,N_13035);
and U13331 (N_13331,N_13047,N_13014);
and U13332 (N_13332,N_13048,N_13085);
xor U13333 (N_13333,N_13121,N_13197);
and U13334 (N_13334,N_13020,N_13045);
xor U13335 (N_13335,N_13180,N_13052);
and U13336 (N_13336,N_13040,N_13157);
nor U13337 (N_13337,N_13179,N_13165);
and U13338 (N_13338,N_13067,N_13015);
nor U13339 (N_13339,N_13057,N_13004);
or U13340 (N_13340,N_13017,N_13092);
or U13341 (N_13341,N_13081,N_13014);
xnor U13342 (N_13342,N_13081,N_13142);
or U13343 (N_13343,N_13050,N_13003);
or U13344 (N_13344,N_13188,N_13129);
and U13345 (N_13345,N_13066,N_13181);
or U13346 (N_13346,N_13060,N_13005);
xor U13347 (N_13347,N_13065,N_13168);
nand U13348 (N_13348,N_13067,N_13190);
xor U13349 (N_13349,N_13013,N_13063);
nand U13350 (N_13350,N_13122,N_13026);
xor U13351 (N_13351,N_13147,N_13159);
and U13352 (N_13352,N_13199,N_13113);
and U13353 (N_13353,N_13034,N_13005);
nand U13354 (N_13354,N_13111,N_13144);
nand U13355 (N_13355,N_13196,N_13116);
or U13356 (N_13356,N_13079,N_13096);
nand U13357 (N_13357,N_13074,N_13112);
xnor U13358 (N_13358,N_13198,N_13110);
xnor U13359 (N_13359,N_13147,N_13130);
or U13360 (N_13360,N_13164,N_13110);
nand U13361 (N_13361,N_13192,N_13191);
xor U13362 (N_13362,N_13086,N_13167);
or U13363 (N_13363,N_13081,N_13002);
xnor U13364 (N_13364,N_13195,N_13061);
and U13365 (N_13365,N_13062,N_13054);
or U13366 (N_13366,N_13076,N_13135);
xnor U13367 (N_13367,N_13128,N_13042);
xor U13368 (N_13368,N_13117,N_13132);
nand U13369 (N_13369,N_13010,N_13173);
nand U13370 (N_13370,N_13137,N_13086);
nor U13371 (N_13371,N_13130,N_13052);
nand U13372 (N_13372,N_13030,N_13125);
or U13373 (N_13373,N_13096,N_13148);
or U13374 (N_13374,N_13045,N_13170);
or U13375 (N_13375,N_13133,N_13153);
nand U13376 (N_13376,N_13060,N_13180);
xnor U13377 (N_13377,N_13005,N_13186);
or U13378 (N_13378,N_13166,N_13106);
and U13379 (N_13379,N_13053,N_13068);
nor U13380 (N_13380,N_13030,N_13057);
xor U13381 (N_13381,N_13198,N_13074);
xor U13382 (N_13382,N_13116,N_13154);
or U13383 (N_13383,N_13040,N_13174);
nand U13384 (N_13384,N_13137,N_13131);
nand U13385 (N_13385,N_13190,N_13003);
or U13386 (N_13386,N_13106,N_13103);
xnor U13387 (N_13387,N_13033,N_13107);
nand U13388 (N_13388,N_13022,N_13185);
and U13389 (N_13389,N_13069,N_13025);
nand U13390 (N_13390,N_13136,N_13066);
xnor U13391 (N_13391,N_13091,N_13108);
nor U13392 (N_13392,N_13074,N_13073);
nor U13393 (N_13393,N_13046,N_13012);
xnor U13394 (N_13394,N_13095,N_13196);
nand U13395 (N_13395,N_13175,N_13190);
nand U13396 (N_13396,N_13048,N_13131);
nor U13397 (N_13397,N_13041,N_13152);
and U13398 (N_13398,N_13094,N_13181);
xor U13399 (N_13399,N_13170,N_13026);
xnor U13400 (N_13400,N_13288,N_13201);
xor U13401 (N_13401,N_13260,N_13265);
nand U13402 (N_13402,N_13350,N_13305);
or U13403 (N_13403,N_13285,N_13250);
nand U13404 (N_13404,N_13258,N_13303);
and U13405 (N_13405,N_13280,N_13311);
nor U13406 (N_13406,N_13375,N_13371);
or U13407 (N_13407,N_13242,N_13262);
nand U13408 (N_13408,N_13306,N_13214);
and U13409 (N_13409,N_13398,N_13388);
nor U13410 (N_13410,N_13297,N_13391);
and U13411 (N_13411,N_13358,N_13268);
or U13412 (N_13412,N_13319,N_13218);
xnor U13413 (N_13413,N_13246,N_13219);
and U13414 (N_13414,N_13253,N_13396);
or U13415 (N_13415,N_13333,N_13314);
or U13416 (N_13416,N_13317,N_13393);
nand U13417 (N_13417,N_13276,N_13251);
nor U13418 (N_13418,N_13300,N_13216);
and U13419 (N_13419,N_13349,N_13243);
and U13420 (N_13420,N_13325,N_13362);
nor U13421 (N_13421,N_13222,N_13245);
or U13422 (N_13422,N_13345,N_13360);
nor U13423 (N_13423,N_13205,N_13378);
nor U13424 (N_13424,N_13323,N_13292);
nand U13425 (N_13425,N_13346,N_13359);
nand U13426 (N_13426,N_13293,N_13357);
or U13427 (N_13427,N_13389,N_13334);
xor U13428 (N_13428,N_13225,N_13263);
nor U13429 (N_13429,N_13229,N_13208);
xor U13430 (N_13430,N_13213,N_13384);
and U13431 (N_13431,N_13365,N_13215);
nor U13432 (N_13432,N_13284,N_13249);
nor U13433 (N_13433,N_13294,N_13271);
nor U13434 (N_13434,N_13383,N_13301);
nand U13435 (N_13435,N_13316,N_13361);
nand U13436 (N_13436,N_13283,N_13264);
or U13437 (N_13437,N_13237,N_13256);
and U13438 (N_13438,N_13296,N_13312);
and U13439 (N_13439,N_13254,N_13318);
or U13440 (N_13440,N_13341,N_13255);
and U13441 (N_13441,N_13313,N_13373);
and U13442 (N_13442,N_13269,N_13347);
xnor U13443 (N_13443,N_13340,N_13364);
or U13444 (N_13444,N_13230,N_13370);
or U13445 (N_13445,N_13377,N_13363);
xnor U13446 (N_13446,N_13392,N_13381);
xnor U13447 (N_13447,N_13202,N_13307);
and U13448 (N_13448,N_13295,N_13374);
xor U13449 (N_13449,N_13287,N_13308);
xnor U13450 (N_13450,N_13239,N_13261);
and U13451 (N_13451,N_13210,N_13372);
or U13452 (N_13452,N_13231,N_13257);
nand U13453 (N_13453,N_13366,N_13228);
and U13454 (N_13454,N_13220,N_13356);
nor U13455 (N_13455,N_13326,N_13273);
and U13456 (N_13456,N_13304,N_13277);
or U13457 (N_13457,N_13338,N_13353);
or U13458 (N_13458,N_13328,N_13380);
xnor U13459 (N_13459,N_13227,N_13248);
nand U13460 (N_13460,N_13339,N_13235);
or U13461 (N_13461,N_13233,N_13200);
and U13462 (N_13462,N_13320,N_13289);
and U13463 (N_13463,N_13206,N_13386);
nand U13464 (N_13464,N_13259,N_13309);
and U13465 (N_13465,N_13234,N_13342);
nand U13466 (N_13466,N_13337,N_13315);
nor U13467 (N_13467,N_13212,N_13291);
nand U13468 (N_13468,N_13369,N_13355);
nor U13469 (N_13469,N_13274,N_13322);
and U13470 (N_13470,N_13298,N_13379);
nor U13471 (N_13471,N_13266,N_13387);
xor U13472 (N_13472,N_13221,N_13390);
and U13473 (N_13473,N_13332,N_13209);
nand U13474 (N_13474,N_13330,N_13367);
and U13475 (N_13475,N_13207,N_13211);
nand U13476 (N_13476,N_13335,N_13281);
and U13477 (N_13477,N_13244,N_13336);
xor U13478 (N_13478,N_13290,N_13232);
or U13479 (N_13479,N_13352,N_13310);
or U13480 (N_13480,N_13240,N_13286);
nand U13481 (N_13481,N_13302,N_13376);
and U13482 (N_13482,N_13321,N_13278);
xor U13483 (N_13483,N_13203,N_13368);
nor U13484 (N_13484,N_13299,N_13351);
xnor U13485 (N_13485,N_13343,N_13354);
nand U13486 (N_13486,N_13238,N_13224);
xor U13487 (N_13487,N_13385,N_13247);
and U13488 (N_13488,N_13252,N_13204);
nand U13489 (N_13489,N_13226,N_13327);
nor U13490 (N_13490,N_13344,N_13382);
or U13491 (N_13491,N_13217,N_13236);
or U13492 (N_13492,N_13331,N_13324);
nand U13493 (N_13493,N_13267,N_13282);
nand U13494 (N_13494,N_13395,N_13270);
xnor U13495 (N_13495,N_13241,N_13397);
xor U13496 (N_13496,N_13399,N_13223);
and U13497 (N_13497,N_13348,N_13394);
nand U13498 (N_13498,N_13279,N_13275);
xor U13499 (N_13499,N_13329,N_13272);
or U13500 (N_13500,N_13346,N_13301);
or U13501 (N_13501,N_13338,N_13203);
and U13502 (N_13502,N_13238,N_13303);
nand U13503 (N_13503,N_13275,N_13361);
xor U13504 (N_13504,N_13243,N_13327);
nand U13505 (N_13505,N_13314,N_13216);
nand U13506 (N_13506,N_13335,N_13343);
or U13507 (N_13507,N_13298,N_13227);
xor U13508 (N_13508,N_13246,N_13368);
and U13509 (N_13509,N_13294,N_13207);
nor U13510 (N_13510,N_13227,N_13229);
xnor U13511 (N_13511,N_13253,N_13262);
or U13512 (N_13512,N_13334,N_13238);
nand U13513 (N_13513,N_13274,N_13240);
nor U13514 (N_13514,N_13225,N_13275);
nand U13515 (N_13515,N_13230,N_13302);
or U13516 (N_13516,N_13206,N_13253);
and U13517 (N_13517,N_13337,N_13232);
xnor U13518 (N_13518,N_13353,N_13203);
nor U13519 (N_13519,N_13344,N_13264);
xor U13520 (N_13520,N_13213,N_13396);
nand U13521 (N_13521,N_13321,N_13274);
xor U13522 (N_13522,N_13217,N_13330);
nor U13523 (N_13523,N_13248,N_13253);
and U13524 (N_13524,N_13237,N_13258);
and U13525 (N_13525,N_13301,N_13216);
nand U13526 (N_13526,N_13200,N_13393);
nand U13527 (N_13527,N_13332,N_13325);
or U13528 (N_13528,N_13212,N_13346);
xnor U13529 (N_13529,N_13211,N_13286);
nor U13530 (N_13530,N_13297,N_13203);
nand U13531 (N_13531,N_13383,N_13345);
or U13532 (N_13532,N_13211,N_13321);
or U13533 (N_13533,N_13234,N_13255);
nor U13534 (N_13534,N_13206,N_13323);
nand U13535 (N_13535,N_13263,N_13234);
nand U13536 (N_13536,N_13253,N_13200);
and U13537 (N_13537,N_13229,N_13271);
nand U13538 (N_13538,N_13303,N_13353);
nand U13539 (N_13539,N_13225,N_13243);
nor U13540 (N_13540,N_13382,N_13356);
or U13541 (N_13541,N_13270,N_13279);
nor U13542 (N_13542,N_13380,N_13341);
xor U13543 (N_13543,N_13336,N_13273);
xnor U13544 (N_13544,N_13332,N_13254);
and U13545 (N_13545,N_13285,N_13373);
nand U13546 (N_13546,N_13312,N_13220);
nor U13547 (N_13547,N_13369,N_13232);
xnor U13548 (N_13548,N_13285,N_13319);
and U13549 (N_13549,N_13293,N_13278);
or U13550 (N_13550,N_13202,N_13323);
xor U13551 (N_13551,N_13354,N_13268);
nand U13552 (N_13552,N_13382,N_13222);
xnor U13553 (N_13553,N_13323,N_13213);
nor U13554 (N_13554,N_13272,N_13270);
nand U13555 (N_13555,N_13246,N_13249);
or U13556 (N_13556,N_13235,N_13246);
nor U13557 (N_13557,N_13305,N_13264);
or U13558 (N_13558,N_13379,N_13327);
nor U13559 (N_13559,N_13365,N_13216);
and U13560 (N_13560,N_13224,N_13324);
and U13561 (N_13561,N_13357,N_13266);
nor U13562 (N_13562,N_13350,N_13280);
xor U13563 (N_13563,N_13369,N_13329);
nor U13564 (N_13564,N_13210,N_13233);
and U13565 (N_13565,N_13353,N_13275);
xnor U13566 (N_13566,N_13361,N_13314);
xnor U13567 (N_13567,N_13249,N_13383);
xnor U13568 (N_13568,N_13390,N_13371);
nor U13569 (N_13569,N_13298,N_13334);
nor U13570 (N_13570,N_13390,N_13288);
nor U13571 (N_13571,N_13320,N_13351);
nand U13572 (N_13572,N_13342,N_13218);
and U13573 (N_13573,N_13255,N_13230);
and U13574 (N_13574,N_13396,N_13363);
or U13575 (N_13575,N_13329,N_13333);
xnor U13576 (N_13576,N_13366,N_13350);
xnor U13577 (N_13577,N_13346,N_13214);
nand U13578 (N_13578,N_13246,N_13262);
and U13579 (N_13579,N_13388,N_13288);
or U13580 (N_13580,N_13391,N_13284);
nand U13581 (N_13581,N_13310,N_13351);
or U13582 (N_13582,N_13392,N_13271);
nor U13583 (N_13583,N_13329,N_13239);
nand U13584 (N_13584,N_13395,N_13242);
xnor U13585 (N_13585,N_13285,N_13368);
xor U13586 (N_13586,N_13359,N_13397);
nand U13587 (N_13587,N_13350,N_13337);
or U13588 (N_13588,N_13250,N_13321);
xnor U13589 (N_13589,N_13302,N_13222);
nor U13590 (N_13590,N_13257,N_13342);
or U13591 (N_13591,N_13206,N_13302);
nand U13592 (N_13592,N_13234,N_13311);
xor U13593 (N_13593,N_13361,N_13371);
nor U13594 (N_13594,N_13292,N_13205);
or U13595 (N_13595,N_13364,N_13394);
or U13596 (N_13596,N_13213,N_13205);
or U13597 (N_13597,N_13298,N_13220);
and U13598 (N_13598,N_13251,N_13248);
or U13599 (N_13599,N_13331,N_13387);
xnor U13600 (N_13600,N_13592,N_13531);
or U13601 (N_13601,N_13572,N_13599);
xnor U13602 (N_13602,N_13541,N_13464);
nor U13603 (N_13603,N_13462,N_13578);
nor U13604 (N_13604,N_13480,N_13551);
or U13605 (N_13605,N_13453,N_13526);
xor U13606 (N_13606,N_13476,N_13477);
xor U13607 (N_13607,N_13485,N_13412);
or U13608 (N_13608,N_13594,N_13493);
or U13609 (N_13609,N_13545,N_13590);
nor U13610 (N_13610,N_13484,N_13593);
nand U13611 (N_13611,N_13556,N_13536);
nand U13612 (N_13612,N_13499,N_13549);
nor U13613 (N_13613,N_13431,N_13447);
or U13614 (N_13614,N_13442,N_13420);
and U13615 (N_13615,N_13587,N_13538);
or U13616 (N_13616,N_13466,N_13577);
nor U13617 (N_13617,N_13405,N_13438);
and U13618 (N_13618,N_13585,N_13422);
xor U13619 (N_13619,N_13570,N_13562);
and U13620 (N_13620,N_13471,N_13535);
or U13621 (N_13621,N_13403,N_13576);
nand U13622 (N_13622,N_13546,N_13441);
nor U13623 (N_13623,N_13463,N_13514);
and U13624 (N_13624,N_13490,N_13415);
xnor U13625 (N_13625,N_13452,N_13418);
nand U13626 (N_13626,N_13513,N_13448);
xnor U13627 (N_13627,N_13457,N_13487);
or U13628 (N_13628,N_13416,N_13410);
nor U13629 (N_13629,N_13524,N_13512);
and U13630 (N_13630,N_13552,N_13501);
or U13631 (N_13631,N_13472,N_13433);
nand U13632 (N_13632,N_13543,N_13517);
xnor U13633 (N_13633,N_13561,N_13586);
nand U13634 (N_13634,N_13522,N_13423);
and U13635 (N_13635,N_13525,N_13451);
nor U13636 (N_13636,N_13529,N_13483);
nand U13637 (N_13637,N_13569,N_13437);
nor U13638 (N_13638,N_13467,N_13443);
nor U13639 (N_13639,N_13439,N_13488);
xor U13640 (N_13640,N_13571,N_13544);
nor U13641 (N_13641,N_13589,N_13559);
nor U13642 (N_13642,N_13547,N_13436);
or U13643 (N_13643,N_13555,N_13530);
nor U13644 (N_13644,N_13478,N_13429);
nand U13645 (N_13645,N_13475,N_13519);
or U13646 (N_13646,N_13591,N_13579);
or U13647 (N_13647,N_13406,N_13596);
or U13648 (N_13648,N_13520,N_13409);
nand U13649 (N_13649,N_13560,N_13533);
nand U13650 (N_13650,N_13421,N_13516);
xnor U13651 (N_13651,N_13446,N_13563);
and U13652 (N_13652,N_13414,N_13540);
nand U13653 (N_13653,N_13491,N_13504);
nand U13654 (N_13654,N_13408,N_13444);
nor U13655 (N_13655,N_13427,N_13510);
nor U13656 (N_13656,N_13404,N_13469);
xor U13657 (N_13657,N_13402,N_13567);
nor U13658 (N_13658,N_13494,N_13509);
or U13659 (N_13659,N_13479,N_13550);
xnor U13660 (N_13660,N_13445,N_13511);
nand U13661 (N_13661,N_13458,N_13532);
nand U13662 (N_13662,N_13450,N_13580);
nand U13663 (N_13663,N_13548,N_13523);
xnor U13664 (N_13664,N_13507,N_13461);
nand U13665 (N_13665,N_13468,N_13582);
and U13666 (N_13666,N_13503,N_13474);
and U13667 (N_13667,N_13500,N_13449);
xor U13668 (N_13668,N_13425,N_13481);
or U13669 (N_13669,N_13595,N_13539);
nand U13670 (N_13670,N_13465,N_13534);
or U13671 (N_13671,N_13489,N_13424);
nor U13672 (N_13672,N_13558,N_13455);
nor U13673 (N_13673,N_13454,N_13417);
nand U13674 (N_13674,N_13413,N_13473);
nor U13675 (N_13675,N_13498,N_13515);
and U13676 (N_13676,N_13568,N_13432);
nand U13677 (N_13677,N_13574,N_13518);
xnor U13678 (N_13678,N_13456,N_13581);
or U13679 (N_13679,N_13400,N_13527);
and U13680 (N_13680,N_13573,N_13537);
nor U13681 (N_13681,N_13459,N_13486);
and U13682 (N_13682,N_13553,N_13460);
or U13683 (N_13683,N_13506,N_13508);
nand U13684 (N_13684,N_13554,N_13435);
and U13685 (N_13685,N_13428,N_13411);
xor U13686 (N_13686,N_13542,N_13583);
and U13687 (N_13687,N_13575,N_13401);
xnor U13688 (N_13688,N_13495,N_13588);
or U13689 (N_13689,N_13565,N_13528);
nor U13690 (N_13690,N_13564,N_13597);
nor U13691 (N_13691,N_13470,N_13505);
nand U13692 (N_13692,N_13434,N_13502);
nand U13693 (N_13693,N_13430,N_13426);
or U13694 (N_13694,N_13557,N_13566);
nor U13695 (N_13695,N_13482,N_13419);
or U13696 (N_13696,N_13492,N_13521);
xor U13697 (N_13697,N_13497,N_13584);
and U13698 (N_13698,N_13496,N_13440);
nor U13699 (N_13699,N_13407,N_13598);
nor U13700 (N_13700,N_13409,N_13554);
xnor U13701 (N_13701,N_13436,N_13541);
and U13702 (N_13702,N_13450,N_13477);
xor U13703 (N_13703,N_13512,N_13534);
xor U13704 (N_13704,N_13492,N_13510);
or U13705 (N_13705,N_13441,N_13582);
or U13706 (N_13706,N_13504,N_13454);
nor U13707 (N_13707,N_13427,N_13566);
or U13708 (N_13708,N_13491,N_13424);
nand U13709 (N_13709,N_13451,N_13560);
xnor U13710 (N_13710,N_13517,N_13496);
nand U13711 (N_13711,N_13513,N_13484);
and U13712 (N_13712,N_13444,N_13478);
or U13713 (N_13713,N_13596,N_13508);
nor U13714 (N_13714,N_13587,N_13409);
xnor U13715 (N_13715,N_13495,N_13461);
or U13716 (N_13716,N_13583,N_13531);
nor U13717 (N_13717,N_13472,N_13477);
nand U13718 (N_13718,N_13414,N_13403);
nor U13719 (N_13719,N_13426,N_13572);
nor U13720 (N_13720,N_13565,N_13453);
nor U13721 (N_13721,N_13527,N_13517);
nor U13722 (N_13722,N_13573,N_13472);
xor U13723 (N_13723,N_13497,N_13562);
xor U13724 (N_13724,N_13414,N_13400);
and U13725 (N_13725,N_13533,N_13504);
nand U13726 (N_13726,N_13574,N_13553);
nand U13727 (N_13727,N_13578,N_13565);
and U13728 (N_13728,N_13505,N_13431);
xor U13729 (N_13729,N_13539,N_13449);
or U13730 (N_13730,N_13408,N_13468);
nor U13731 (N_13731,N_13433,N_13419);
or U13732 (N_13732,N_13597,N_13465);
or U13733 (N_13733,N_13415,N_13564);
or U13734 (N_13734,N_13598,N_13477);
nor U13735 (N_13735,N_13547,N_13577);
xnor U13736 (N_13736,N_13599,N_13433);
nor U13737 (N_13737,N_13519,N_13529);
xor U13738 (N_13738,N_13483,N_13433);
xor U13739 (N_13739,N_13468,N_13433);
and U13740 (N_13740,N_13556,N_13433);
nand U13741 (N_13741,N_13492,N_13422);
nand U13742 (N_13742,N_13469,N_13546);
or U13743 (N_13743,N_13413,N_13444);
nor U13744 (N_13744,N_13599,N_13446);
or U13745 (N_13745,N_13563,N_13426);
or U13746 (N_13746,N_13593,N_13569);
xnor U13747 (N_13747,N_13412,N_13526);
nor U13748 (N_13748,N_13583,N_13470);
nor U13749 (N_13749,N_13468,N_13544);
xor U13750 (N_13750,N_13553,N_13538);
nand U13751 (N_13751,N_13425,N_13553);
xnor U13752 (N_13752,N_13405,N_13501);
xnor U13753 (N_13753,N_13419,N_13560);
or U13754 (N_13754,N_13487,N_13476);
xor U13755 (N_13755,N_13426,N_13544);
nor U13756 (N_13756,N_13443,N_13531);
xor U13757 (N_13757,N_13485,N_13486);
and U13758 (N_13758,N_13441,N_13530);
nand U13759 (N_13759,N_13460,N_13418);
xnor U13760 (N_13760,N_13472,N_13507);
xor U13761 (N_13761,N_13553,N_13572);
xnor U13762 (N_13762,N_13590,N_13501);
xnor U13763 (N_13763,N_13583,N_13530);
nor U13764 (N_13764,N_13415,N_13587);
nor U13765 (N_13765,N_13475,N_13527);
nor U13766 (N_13766,N_13425,N_13558);
and U13767 (N_13767,N_13470,N_13558);
and U13768 (N_13768,N_13475,N_13562);
nand U13769 (N_13769,N_13574,N_13577);
nand U13770 (N_13770,N_13419,N_13583);
nand U13771 (N_13771,N_13415,N_13449);
nand U13772 (N_13772,N_13556,N_13439);
and U13773 (N_13773,N_13454,N_13470);
xnor U13774 (N_13774,N_13501,N_13441);
xnor U13775 (N_13775,N_13417,N_13495);
nand U13776 (N_13776,N_13447,N_13515);
or U13777 (N_13777,N_13480,N_13540);
xnor U13778 (N_13778,N_13409,N_13572);
nor U13779 (N_13779,N_13512,N_13437);
nor U13780 (N_13780,N_13452,N_13510);
nor U13781 (N_13781,N_13475,N_13575);
nor U13782 (N_13782,N_13403,N_13581);
nor U13783 (N_13783,N_13548,N_13514);
and U13784 (N_13784,N_13506,N_13443);
or U13785 (N_13785,N_13543,N_13538);
or U13786 (N_13786,N_13462,N_13553);
xnor U13787 (N_13787,N_13535,N_13528);
xnor U13788 (N_13788,N_13513,N_13511);
or U13789 (N_13789,N_13492,N_13478);
nor U13790 (N_13790,N_13498,N_13575);
xnor U13791 (N_13791,N_13531,N_13581);
and U13792 (N_13792,N_13475,N_13427);
and U13793 (N_13793,N_13452,N_13497);
nand U13794 (N_13794,N_13402,N_13551);
xor U13795 (N_13795,N_13529,N_13586);
nand U13796 (N_13796,N_13549,N_13460);
or U13797 (N_13797,N_13454,N_13543);
nor U13798 (N_13798,N_13560,N_13589);
or U13799 (N_13799,N_13539,N_13557);
nor U13800 (N_13800,N_13678,N_13719);
and U13801 (N_13801,N_13662,N_13640);
nand U13802 (N_13802,N_13780,N_13675);
nor U13803 (N_13803,N_13623,N_13771);
nand U13804 (N_13804,N_13611,N_13657);
nor U13805 (N_13805,N_13783,N_13762);
and U13806 (N_13806,N_13788,N_13751);
and U13807 (N_13807,N_13679,N_13641);
or U13808 (N_13808,N_13778,N_13682);
nor U13809 (N_13809,N_13749,N_13646);
xnor U13810 (N_13810,N_13633,N_13631);
or U13811 (N_13811,N_13745,N_13777);
or U13812 (N_13812,N_13651,N_13645);
or U13813 (N_13813,N_13764,N_13725);
or U13814 (N_13814,N_13715,N_13655);
xor U13815 (N_13815,N_13667,N_13659);
and U13816 (N_13816,N_13643,N_13644);
nand U13817 (N_13817,N_13779,N_13602);
or U13818 (N_13818,N_13648,N_13731);
and U13819 (N_13819,N_13649,N_13743);
and U13820 (N_13820,N_13639,N_13609);
xnor U13821 (N_13821,N_13632,N_13683);
nand U13822 (N_13822,N_13753,N_13693);
or U13823 (N_13823,N_13757,N_13746);
or U13824 (N_13824,N_13617,N_13653);
xor U13825 (N_13825,N_13752,N_13766);
nor U13826 (N_13826,N_13716,N_13626);
xor U13827 (N_13827,N_13625,N_13692);
nor U13828 (N_13828,N_13671,N_13768);
xor U13829 (N_13829,N_13786,N_13728);
nor U13830 (N_13830,N_13724,N_13629);
nor U13831 (N_13831,N_13704,N_13736);
nand U13832 (N_13832,N_13707,N_13785);
xor U13833 (N_13833,N_13795,N_13636);
nor U13834 (N_13834,N_13672,N_13601);
nor U13835 (N_13835,N_13723,N_13787);
nand U13836 (N_13836,N_13697,N_13620);
nand U13837 (N_13837,N_13621,N_13790);
or U13838 (N_13838,N_13739,N_13773);
nand U13839 (N_13839,N_13767,N_13690);
nor U13840 (N_13840,N_13726,N_13742);
and U13841 (N_13841,N_13684,N_13670);
nor U13842 (N_13842,N_13732,N_13776);
xor U13843 (N_13843,N_13676,N_13694);
xnor U13844 (N_13844,N_13734,N_13763);
nand U13845 (N_13845,N_13748,N_13661);
nand U13846 (N_13846,N_13614,N_13769);
or U13847 (N_13847,N_13663,N_13691);
nor U13848 (N_13848,N_13666,N_13656);
nand U13849 (N_13849,N_13782,N_13624);
nor U13850 (N_13850,N_13792,N_13754);
nor U13851 (N_13851,N_13711,N_13673);
or U13852 (N_13852,N_13789,N_13775);
or U13853 (N_13853,N_13760,N_13647);
xor U13854 (N_13854,N_13689,N_13721);
xnor U13855 (N_13855,N_13628,N_13607);
xor U13856 (N_13856,N_13677,N_13613);
xnor U13857 (N_13857,N_13695,N_13705);
nor U13858 (N_13858,N_13722,N_13703);
or U13859 (N_13859,N_13619,N_13637);
or U13860 (N_13860,N_13714,N_13627);
and U13861 (N_13861,N_13712,N_13658);
and U13862 (N_13862,N_13793,N_13616);
or U13863 (N_13863,N_13781,N_13744);
xor U13864 (N_13864,N_13688,N_13765);
nor U13865 (N_13865,N_13727,N_13750);
xor U13866 (N_13866,N_13713,N_13642);
and U13867 (N_13867,N_13733,N_13615);
nand U13868 (N_13868,N_13730,N_13741);
or U13869 (N_13869,N_13604,N_13791);
and U13870 (N_13870,N_13696,N_13664);
and U13871 (N_13871,N_13608,N_13710);
nor U13872 (N_13872,N_13622,N_13700);
or U13873 (N_13873,N_13669,N_13794);
nand U13874 (N_13874,N_13654,N_13799);
nand U13875 (N_13875,N_13702,N_13685);
nand U13876 (N_13876,N_13761,N_13606);
and U13877 (N_13877,N_13660,N_13701);
and U13878 (N_13878,N_13796,N_13755);
xnor U13879 (N_13879,N_13729,N_13699);
and U13880 (N_13880,N_13709,N_13797);
nand U13881 (N_13881,N_13770,N_13610);
or U13882 (N_13882,N_13668,N_13612);
nor U13883 (N_13883,N_13740,N_13650);
nor U13884 (N_13884,N_13708,N_13784);
xnor U13885 (N_13885,N_13717,N_13774);
and U13886 (N_13886,N_13665,N_13735);
xor U13887 (N_13887,N_13687,N_13720);
nor U13888 (N_13888,N_13674,N_13634);
xnor U13889 (N_13889,N_13681,N_13756);
nand U13890 (N_13890,N_13635,N_13638);
and U13891 (N_13891,N_13759,N_13630);
xnor U13892 (N_13892,N_13772,N_13603);
and U13893 (N_13893,N_13680,N_13718);
or U13894 (N_13894,N_13798,N_13698);
and U13895 (N_13895,N_13686,N_13738);
nor U13896 (N_13896,N_13758,N_13605);
or U13897 (N_13897,N_13618,N_13600);
or U13898 (N_13898,N_13706,N_13747);
and U13899 (N_13899,N_13737,N_13652);
nor U13900 (N_13900,N_13795,N_13768);
nand U13901 (N_13901,N_13604,N_13735);
nand U13902 (N_13902,N_13795,N_13732);
nand U13903 (N_13903,N_13639,N_13668);
or U13904 (N_13904,N_13788,N_13615);
and U13905 (N_13905,N_13639,N_13775);
or U13906 (N_13906,N_13630,N_13723);
xor U13907 (N_13907,N_13755,N_13622);
nor U13908 (N_13908,N_13790,N_13684);
nor U13909 (N_13909,N_13605,N_13795);
or U13910 (N_13910,N_13642,N_13683);
xnor U13911 (N_13911,N_13657,N_13779);
and U13912 (N_13912,N_13741,N_13761);
or U13913 (N_13913,N_13689,N_13639);
and U13914 (N_13914,N_13709,N_13619);
nor U13915 (N_13915,N_13698,N_13753);
xor U13916 (N_13916,N_13794,N_13682);
nand U13917 (N_13917,N_13710,N_13717);
and U13918 (N_13918,N_13678,N_13761);
nand U13919 (N_13919,N_13634,N_13708);
nor U13920 (N_13920,N_13789,N_13666);
nor U13921 (N_13921,N_13795,N_13682);
xnor U13922 (N_13922,N_13760,N_13632);
nand U13923 (N_13923,N_13600,N_13711);
or U13924 (N_13924,N_13763,N_13712);
nor U13925 (N_13925,N_13756,N_13783);
and U13926 (N_13926,N_13695,N_13694);
xor U13927 (N_13927,N_13725,N_13762);
and U13928 (N_13928,N_13705,N_13637);
and U13929 (N_13929,N_13764,N_13743);
or U13930 (N_13930,N_13674,N_13775);
nor U13931 (N_13931,N_13608,N_13603);
nand U13932 (N_13932,N_13632,N_13628);
nor U13933 (N_13933,N_13669,N_13697);
nor U13934 (N_13934,N_13762,N_13613);
nor U13935 (N_13935,N_13676,N_13753);
xor U13936 (N_13936,N_13687,N_13778);
nand U13937 (N_13937,N_13756,N_13706);
xor U13938 (N_13938,N_13733,N_13777);
xnor U13939 (N_13939,N_13711,N_13704);
nor U13940 (N_13940,N_13682,N_13790);
nand U13941 (N_13941,N_13646,N_13687);
or U13942 (N_13942,N_13674,N_13779);
or U13943 (N_13943,N_13617,N_13601);
and U13944 (N_13944,N_13660,N_13751);
nor U13945 (N_13945,N_13720,N_13646);
nor U13946 (N_13946,N_13645,N_13627);
or U13947 (N_13947,N_13709,N_13799);
xor U13948 (N_13948,N_13741,N_13760);
or U13949 (N_13949,N_13705,N_13647);
nor U13950 (N_13950,N_13688,N_13739);
nand U13951 (N_13951,N_13622,N_13626);
or U13952 (N_13952,N_13649,N_13786);
xnor U13953 (N_13953,N_13618,N_13708);
or U13954 (N_13954,N_13608,N_13672);
or U13955 (N_13955,N_13747,N_13664);
xnor U13956 (N_13956,N_13623,N_13789);
and U13957 (N_13957,N_13775,N_13641);
nand U13958 (N_13958,N_13774,N_13678);
and U13959 (N_13959,N_13606,N_13664);
nand U13960 (N_13960,N_13635,N_13795);
nor U13961 (N_13961,N_13664,N_13771);
and U13962 (N_13962,N_13712,N_13725);
or U13963 (N_13963,N_13631,N_13704);
or U13964 (N_13964,N_13615,N_13637);
or U13965 (N_13965,N_13663,N_13638);
and U13966 (N_13966,N_13652,N_13760);
and U13967 (N_13967,N_13769,N_13722);
or U13968 (N_13968,N_13749,N_13763);
xnor U13969 (N_13969,N_13660,N_13619);
nand U13970 (N_13970,N_13614,N_13704);
and U13971 (N_13971,N_13677,N_13602);
xor U13972 (N_13972,N_13685,N_13727);
or U13973 (N_13973,N_13687,N_13741);
and U13974 (N_13974,N_13705,N_13783);
nor U13975 (N_13975,N_13739,N_13658);
xnor U13976 (N_13976,N_13624,N_13718);
nand U13977 (N_13977,N_13616,N_13779);
xnor U13978 (N_13978,N_13719,N_13629);
nor U13979 (N_13979,N_13736,N_13611);
and U13980 (N_13980,N_13759,N_13726);
xor U13981 (N_13981,N_13674,N_13680);
xor U13982 (N_13982,N_13631,N_13628);
and U13983 (N_13983,N_13629,N_13778);
or U13984 (N_13984,N_13794,N_13603);
nor U13985 (N_13985,N_13705,N_13764);
or U13986 (N_13986,N_13783,N_13601);
nand U13987 (N_13987,N_13700,N_13617);
nand U13988 (N_13988,N_13660,N_13739);
xor U13989 (N_13989,N_13799,N_13774);
or U13990 (N_13990,N_13682,N_13659);
or U13991 (N_13991,N_13637,N_13648);
xor U13992 (N_13992,N_13744,N_13608);
xnor U13993 (N_13993,N_13745,N_13722);
nor U13994 (N_13994,N_13752,N_13666);
or U13995 (N_13995,N_13651,N_13631);
nor U13996 (N_13996,N_13664,N_13626);
xnor U13997 (N_13997,N_13604,N_13719);
or U13998 (N_13998,N_13620,N_13676);
and U13999 (N_13999,N_13718,N_13671);
or U14000 (N_14000,N_13980,N_13907);
nor U14001 (N_14001,N_13892,N_13997);
xnor U14002 (N_14002,N_13861,N_13939);
nand U14003 (N_14003,N_13996,N_13933);
nor U14004 (N_14004,N_13972,N_13986);
nand U14005 (N_14005,N_13800,N_13920);
xnor U14006 (N_14006,N_13949,N_13864);
and U14007 (N_14007,N_13801,N_13914);
xnor U14008 (N_14008,N_13802,N_13957);
nand U14009 (N_14009,N_13875,N_13956);
nor U14010 (N_14010,N_13821,N_13873);
nand U14011 (N_14011,N_13947,N_13898);
xor U14012 (N_14012,N_13926,N_13896);
nand U14013 (N_14013,N_13825,N_13908);
nand U14014 (N_14014,N_13839,N_13915);
and U14015 (N_14015,N_13882,N_13835);
nand U14016 (N_14016,N_13814,N_13921);
nor U14017 (N_14017,N_13970,N_13943);
nand U14018 (N_14018,N_13874,N_13832);
and U14019 (N_14019,N_13923,N_13909);
nor U14020 (N_14020,N_13955,N_13824);
xnor U14021 (N_14021,N_13971,N_13884);
xnor U14022 (N_14022,N_13891,N_13853);
nor U14023 (N_14023,N_13890,N_13885);
or U14024 (N_14024,N_13992,N_13975);
nor U14025 (N_14025,N_13940,N_13831);
or U14026 (N_14026,N_13981,N_13846);
nor U14027 (N_14027,N_13925,N_13974);
or U14028 (N_14028,N_13807,N_13993);
xor U14029 (N_14029,N_13944,N_13912);
nand U14030 (N_14030,N_13911,N_13966);
or U14031 (N_14031,N_13936,N_13952);
or U14032 (N_14032,N_13968,N_13994);
nor U14033 (N_14033,N_13872,N_13880);
or U14034 (N_14034,N_13836,N_13870);
nor U14035 (N_14035,N_13827,N_13929);
or U14036 (N_14036,N_13964,N_13894);
nand U14037 (N_14037,N_13951,N_13806);
or U14038 (N_14038,N_13878,N_13843);
or U14039 (N_14039,N_13906,N_13987);
and U14040 (N_14040,N_13818,N_13830);
nor U14041 (N_14041,N_13938,N_13905);
xnor U14042 (N_14042,N_13927,N_13833);
xor U14043 (N_14043,N_13893,N_13983);
xnor U14044 (N_14044,N_13871,N_13904);
and U14045 (N_14045,N_13946,N_13811);
and U14046 (N_14046,N_13865,N_13916);
and U14047 (N_14047,N_13889,N_13937);
nand U14048 (N_14048,N_13854,N_13919);
nand U14049 (N_14049,N_13813,N_13834);
and U14050 (N_14050,N_13950,N_13913);
xor U14051 (N_14051,N_13895,N_13809);
nor U14052 (N_14052,N_13858,N_13852);
xor U14053 (N_14053,N_13804,N_13859);
and U14054 (N_14054,N_13901,N_13953);
nand U14055 (N_14055,N_13828,N_13999);
nand U14056 (N_14056,N_13841,N_13805);
xnor U14057 (N_14057,N_13899,N_13977);
xnor U14058 (N_14058,N_13822,N_13991);
nand U14059 (N_14059,N_13902,N_13917);
xnor U14060 (N_14060,N_13851,N_13945);
or U14061 (N_14061,N_13823,N_13948);
nor U14062 (N_14062,N_13876,N_13862);
nor U14063 (N_14063,N_13829,N_13935);
nor U14064 (N_14064,N_13808,N_13886);
or U14065 (N_14065,N_13815,N_13842);
and U14066 (N_14066,N_13963,N_13863);
nor U14067 (N_14067,N_13988,N_13810);
or U14068 (N_14068,N_13840,N_13934);
nand U14069 (N_14069,N_13989,N_13837);
nor U14070 (N_14070,N_13803,N_13982);
nor U14071 (N_14071,N_13931,N_13887);
or U14072 (N_14072,N_13826,N_13941);
or U14073 (N_14073,N_13942,N_13869);
xor U14074 (N_14074,N_13866,N_13817);
xnor U14075 (N_14075,N_13812,N_13847);
nand U14076 (N_14076,N_13845,N_13900);
or U14077 (N_14077,N_13918,N_13961);
nand U14078 (N_14078,N_13978,N_13820);
and U14079 (N_14079,N_13969,N_13868);
or U14080 (N_14080,N_13848,N_13838);
nor U14081 (N_14081,N_13960,N_13877);
nand U14082 (N_14082,N_13958,N_13967);
nor U14083 (N_14083,N_13879,N_13850);
and U14084 (N_14084,N_13883,N_13984);
nor U14085 (N_14085,N_13998,N_13849);
nor U14086 (N_14086,N_13897,N_13932);
nand U14087 (N_14087,N_13959,N_13985);
nor U14088 (N_14088,N_13855,N_13965);
nor U14089 (N_14089,N_13857,N_13888);
and U14090 (N_14090,N_13976,N_13903);
nor U14091 (N_14091,N_13816,N_13928);
or U14092 (N_14092,N_13979,N_13867);
xnor U14093 (N_14093,N_13962,N_13924);
nor U14094 (N_14094,N_13973,N_13881);
nand U14095 (N_14095,N_13990,N_13910);
nor U14096 (N_14096,N_13844,N_13860);
and U14097 (N_14097,N_13930,N_13995);
or U14098 (N_14098,N_13922,N_13856);
and U14099 (N_14099,N_13819,N_13954);
nand U14100 (N_14100,N_13819,N_13917);
or U14101 (N_14101,N_13839,N_13814);
nand U14102 (N_14102,N_13995,N_13877);
xnor U14103 (N_14103,N_13965,N_13936);
xor U14104 (N_14104,N_13970,N_13882);
or U14105 (N_14105,N_13823,N_13875);
or U14106 (N_14106,N_13881,N_13852);
and U14107 (N_14107,N_13865,N_13821);
and U14108 (N_14108,N_13873,N_13932);
or U14109 (N_14109,N_13900,N_13918);
xor U14110 (N_14110,N_13883,N_13886);
or U14111 (N_14111,N_13916,N_13962);
xor U14112 (N_14112,N_13946,N_13827);
or U14113 (N_14113,N_13801,N_13882);
nand U14114 (N_14114,N_13892,N_13901);
nand U14115 (N_14115,N_13907,N_13995);
nand U14116 (N_14116,N_13877,N_13965);
nand U14117 (N_14117,N_13866,N_13810);
or U14118 (N_14118,N_13828,N_13818);
or U14119 (N_14119,N_13853,N_13864);
nand U14120 (N_14120,N_13828,N_13834);
xor U14121 (N_14121,N_13978,N_13918);
or U14122 (N_14122,N_13945,N_13913);
nor U14123 (N_14123,N_13821,N_13851);
nor U14124 (N_14124,N_13957,N_13972);
or U14125 (N_14125,N_13979,N_13849);
nand U14126 (N_14126,N_13906,N_13913);
and U14127 (N_14127,N_13947,N_13861);
nand U14128 (N_14128,N_13889,N_13925);
or U14129 (N_14129,N_13851,N_13899);
and U14130 (N_14130,N_13858,N_13996);
and U14131 (N_14131,N_13913,N_13875);
nor U14132 (N_14132,N_13979,N_13914);
nand U14133 (N_14133,N_13856,N_13996);
or U14134 (N_14134,N_13949,N_13901);
nor U14135 (N_14135,N_13809,N_13976);
and U14136 (N_14136,N_13853,N_13801);
nor U14137 (N_14137,N_13872,N_13904);
and U14138 (N_14138,N_13843,N_13879);
or U14139 (N_14139,N_13976,N_13906);
and U14140 (N_14140,N_13901,N_13850);
and U14141 (N_14141,N_13969,N_13850);
xor U14142 (N_14142,N_13818,N_13894);
or U14143 (N_14143,N_13963,N_13890);
and U14144 (N_14144,N_13924,N_13880);
and U14145 (N_14145,N_13838,N_13857);
nor U14146 (N_14146,N_13992,N_13803);
and U14147 (N_14147,N_13917,N_13803);
xor U14148 (N_14148,N_13916,N_13800);
xor U14149 (N_14149,N_13826,N_13981);
nor U14150 (N_14150,N_13979,N_13908);
or U14151 (N_14151,N_13914,N_13971);
xnor U14152 (N_14152,N_13930,N_13833);
and U14153 (N_14153,N_13862,N_13900);
xor U14154 (N_14154,N_13827,N_13870);
xnor U14155 (N_14155,N_13818,N_13985);
and U14156 (N_14156,N_13951,N_13946);
xnor U14157 (N_14157,N_13802,N_13838);
or U14158 (N_14158,N_13898,N_13998);
xnor U14159 (N_14159,N_13818,N_13942);
nor U14160 (N_14160,N_13886,N_13837);
nand U14161 (N_14161,N_13905,N_13820);
xnor U14162 (N_14162,N_13841,N_13968);
and U14163 (N_14163,N_13987,N_13943);
xnor U14164 (N_14164,N_13819,N_13945);
xnor U14165 (N_14165,N_13833,N_13906);
xor U14166 (N_14166,N_13979,N_13935);
and U14167 (N_14167,N_13983,N_13964);
nand U14168 (N_14168,N_13960,N_13993);
nor U14169 (N_14169,N_13905,N_13947);
and U14170 (N_14170,N_13885,N_13915);
nor U14171 (N_14171,N_13927,N_13814);
xor U14172 (N_14172,N_13954,N_13993);
xor U14173 (N_14173,N_13807,N_13811);
or U14174 (N_14174,N_13823,N_13925);
nand U14175 (N_14175,N_13962,N_13982);
and U14176 (N_14176,N_13867,N_13965);
nor U14177 (N_14177,N_13839,N_13875);
nand U14178 (N_14178,N_13835,N_13811);
and U14179 (N_14179,N_13940,N_13955);
xnor U14180 (N_14180,N_13929,N_13810);
and U14181 (N_14181,N_13879,N_13973);
nor U14182 (N_14182,N_13887,N_13886);
and U14183 (N_14183,N_13854,N_13827);
xnor U14184 (N_14184,N_13851,N_13853);
or U14185 (N_14185,N_13969,N_13878);
nand U14186 (N_14186,N_13857,N_13982);
nor U14187 (N_14187,N_13998,N_13945);
and U14188 (N_14188,N_13851,N_13837);
nor U14189 (N_14189,N_13922,N_13962);
nand U14190 (N_14190,N_13805,N_13909);
nand U14191 (N_14191,N_13899,N_13895);
nor U14192 (N_14192,N_13900,N_13836);
nand U14193 (N_14193,N_13900,N_13978);
or U14194 (N_14194,N_13864,N_13918);
nand U14195 (N_14195,N_13879,N_13917);
nand U14196 (N_14196,N_13919,N_13977);
and U14197 (N_14197,N_13905,N_13850);
nand U14198 (N_14198,N_13899,N_13843);
nor U14199 (N_14199,N_13837,N_13968);
or U14200 (N_14200,N_14072,N_14114);
nand U14201 (N_14201,N_14158,N_14075);
or U14202 (N_14202,N_14156,N_14070);
xnor U14203 (N_14203,N_14199,N_14111);
or U14204 (N_14204,N_14018,N_14097);
xnor U14205 (N_14205,N_14115,N_14146);
nor U14206 (N_14206,N_14128,N_14129);
nor U14207 (N_14207,N_14173,N_14047);
xnor U14208 (N_14208,N_14184,N_14071);
xor U14209 (N_14209,N_14085,N_14139);
and U14210 (N_14210,N_14068,N_14086);
or U14211 (N_14211,N_14135,N_14095);
xnor U14212 (N_14212,N_14077,N_14121);
nor U14213 (N_14213,N_14137,N_14040);
nand U14214 (N_14214,N_14175,N_14059);
nor U14215 (N_14215,N_14000,N_14110);
or U14216 (N_14216,N_14002,N_14113);
nand U14217 (N_14217,N_14078,N_14163);
nand U14218 (N_14218,N_14092,N_14025);
and U14219 (N_14219,N_14019,N_14145);
nor U14220 (N_14220,N_14023,N_14049);
nand U14221 (N_14221,N_14159,N_14054);
xor U14222 (N_14222,N_14160,N_14037);
nand U14223 (N_14223,N_14031,N_14117);
xor U14224 (N_14224,N_14043,N_14044);
and U14225 (N_14225,N_14141,N_14197);
or U14226 (N_14226,N_14076,N_14039);
and U14227 (N_14227,N_14195,N_14028);
or U14228 (N_14228,N_14051,N_14073);
and U14229 (N_14229,N_14120,N_14127);
or U14230 (N_14230,N_14003,N_14152);
or U14231 (N_14231,N_14066,N_14100);
nor U14232 (N_14232,N_14150,N_14020);
nor U14233 (N_14233,N_14053,N_14157);
xnor U14234 (N_14234,N_14062,N_14074);
nand U14235 (N_14235,N_14119,N_14176);
or U14236 (N_14236,N_14082,N_14172);
nand U14237 (N_14237,N_14001,N_14084);
or U14238 (N_14238,N_14132,N_14107);
nand U14239 (N_14239,N_14058,N_14178);
and U14240 (N_14240,N_14103,N_14016);
nor U14241 (N_14241,N_14108,N_14013);
nor U14242 (N_14242,N_14151,N_14098);
nand U14243 (N_14243,N_14069,N_14056);
or U14244 (N_14244,N_14138,N_14055);
nor U14245 (N_14245,N_14182,N_14142);
nand U14246 (N_14246,N_14006,N_14034);
nor U14247 (N_14247,N_14079,N_14190);
and U14248 (N_14248,N_14196,N_14126);
or U14249 (N_14249,N_14148,N_14015);
xnor U14250 (N_14250,N_14094,N_14143);
xnor U14251 (N_14251,N_14012,N_14014);
or U14252 (N_14252,N_14166,N_14131);
nand U14253 (N_14253,N_14179,N_14161);
or U14254 (N_14254,N_14189,N_14045);
or U14255 (N_14255,N_14118,N_14004);
and U14256 (N_14256,N_14089,N_14090);
xor U14257 (N_14257,N_14167,N_14191);
nor U14258 (N_14258,N_14099,N_14124);
or U14259 (N_14259,N_14029,N_14093);
xnor U14260 (N_14260,N_14198,N_14130);
xor U14261 (N_14261,N_14183,N_14005);
and U14262 (N_14262,N_14104,N_14109);
xnor U14263 (N_14263,N_14116,N_14033);
and U14264 (N_14264,N_14181,N_14154);
xnor U14265 (N_14265,N_14032,N_14186);
and U14266 (N_14266,N_14180,N_14165);
and U14267 (N_14267,N_14050,N_14106);
and U14268 (N_14268,N_14112,N_14011);
and U14269 (N_14269,N_14088,N_14188);
or U14270 (N_14270,N_14192,N_14164);
xor U14271 (N_14271,N_14194,N_14133);
xor U14272 (N_14272,N_14083,N_14010);
xnor U14273 (N_14273,N_14147,N_14134);
xor U14274 (N_14274,N_14105,N_14060);
xor U14275 (N_14275,N_14169,N_14081);
nor U14276 (N_14276,N_14008,N_14102);
nor U14277 (N_14277,N_14125,N_14168);
nor U14278 (N_14278,N_14162,N_14046);
xor U14279 (N_14279,N_14144,N_14022);
nand U14280 (N_14280,N_14038,N_14026);
nor U14281 (N_14281,N_14171,N_14041);
or U14282 (N_14282,N_14035,N_14007);
nor U14283 (N_14283,N_14027,N_14091);
and U14284 (N_14284,N_14153,N_14174);
nor U14285 (N_14285,N_14048,N_14149);
or U14286 (N_14286,N_14021,N_14065);
and U14287 (N_14287,N_14017,N_14193);
xor U14288 (N_14288,N_14030,N_14185);
or U14289 (N_14289,N_14052,N_14096);
nor U14290 (N_14290,N_14155,N_14177);
xor U14291 (N_14291,N_14063,N_14140);
xnor U14292 (N_14292,N_14122,N_14042);
nand U14293 (N_14293,N_14080,N_14009);
xor U14294 (N_14294,N_14087,N_14024);
or U14295 (N_14295,N_14170,N_14123);
and U14296 (N_14296,N_14064,N_14057);
and U14297 (N_14297,N_14187,N_14136);
and U14298 (N_14298,N_14067,N_14101);
and U14299 (N_14299,N_14061,N_14036);
or U14300 (N_14300,N_14049,N_14089);
nand U14301 (N_14301,N_14040,N_14167);
and U14302 (N_14302,N_14182,N_14096);
xnor U14303 (N_14303,N_14011,N_14007);
nor U14304 (N_14304,N_14168,N_14046);
xnor U14305 (N_14305,N_14024,N_14028);
and U14306 (N_14306,N_14061,N_14067);
nor U14307 (N_14307,N_14185,N_14062);
nand U14308 (N_14308,N_14155,N_14119);
xnor U14309 (N_14309,N_14042,N_14135);
nor U14310 (N_14310,N_14145,N_14170);
and U14311 (N_14311,N_14074,N_14129);
nand U14312 (N_14312,N_14077,N_14066);
nand U14313 (N_14313,N_14059,N_14030);
nor U14314 (N_14314,N_14149,N_14137);
nand U14315 (N_14315,N_14097,N_14113);
nand U14316 (N_14316,N_14161,N_14055);
nor U14317 (N_14317,N_14014,N_14016);
nand U14318 (N_14318,N_14005,N_14056);
xor U14319 (N_14319,N_14174,N_14177);
nor U14320 (N_14320,N_14137,N_14018);
or U14321 (N_14321,N_14157,N_14179);
xnor U14322 (N_14322,N_14050,N_14119);
nand U14323 (N_14323,N_14106,N_14194);
nor U14324 (N_14324,N_14149,N_14178);
nand U14325 (N_14325,N_14145,N_14147);
or U14326 (N_14326,N_14144,N_14158);
and U14327 (N_14327,N_14128,N_14164);
nand U14328 (N_14328,N_14050,N_14080);
or U14329 (N_14329,N_14024,N_14129);
or U14330 (N_14330,N_14008,N_14147);
and U14331 (N_14331,N_14091,N_14162);
and U14332 (N_14332,N_14155,N_14064);
nor U14333 (N_14333,N_14006,N_14174);
nand U14334 (N_14334,N_14119,N_14052);
or U14335 (N_14335,N_14161,N_14154);
and U14336 (N_14336,N_14093,N_14196);
nor U14337 (N_14337,N_14073,N_14193);
or U14338 (N_14338,N_14115,N_14051);
xnor U14339 (N_14339,N_14089,N_14174);
nor U14340 (N_14340,N_14052,N_14047);
and U14341 (N_14341,N_14110,N_14045);
nor U14342 (N_14342,N_14050,N_14040);
or U14343 (N_14343,N_14165,N_14155);
nor U14344 (N_14344,N_14152,N_14002);
and U14345 (N_14345,N_14172,N_14125);
or U14346 (N_14346,N_14002,N_14062);
nor U14347 (N_14347,N_14058,N_14162);
nor U14348 (N_14348,N_14093,N_14045);
and U14349 (N_14349,N_14101,N_14181);
or U14350 (N_14350,N_14171,N_14146);
xnor U14351 (N_14351,N_14197,N_14159);
nor U14352 (N_14352,N_14150,N_14091);
and U14353 (N_14353,N_14150,N_14199);
or U14354 (N_14354,N_14098,N_14056);
nor U14355 (N_14355,N_14098,N_14133);
and U14356 (N_14356,N_14031,N_14032);
nor U14357 (N_14357,N_14162,N_14016);
nand U14358 (N_14358,N_14180,N_14002);
nor U14359 (N_14359,N_14104,N_14063);
and U14360 (N_14360,N_14072,N_14088);
and U14361 (N_14361,N_14122,N_14143);
or U14362 (N_14362,N_14002,N_14006);
or U14363 (N_14363,N_14052,N_14147);
nor U14364 (N_14364,N_14080,N_14063);
xor U14365 (N_14365,N_14198,N_14032);
and U14366 (N_14366,N_14077,N_14100);
and U14367 (N_14367,N_14150,N_14122);
and U14368 (N_14368,N_14080,N_14127);
nor U14369 (N_14369,N_14182,N_14102);
and U14370 (N_14370,N_14129,N_14019);
or U14371 (N_14371,N_14015,N_14160);
or U14372 (N_14372,N_14003,N_14067);
and U14373 (N_14373,N_14027,N_14154);
xor U14374 (N_14374,N_14168,N_14195);
and U14375 (N_14375,N_14022,N_14076);
nand U14376 (N_14376,N_14193,N_14116);
or U14377 (N_14377,N_14116,N_14102);
or U14378 (N_14378,N_14105,N_14199);
nand U14379 (N_14379,N_14175,N_14041);
or U14380 (N_14380,N_14139,N_14190);
xnor U14381 (N_14381,N_14018,N_14142);
or U14382 (N_14382,N_14064,N_14080);
and U14383 (N_14383,N_14115,N_14044);
and U14384 (N_14384,N_14136,N_14013);
or U14385 (N_14385,N_14062,N_14161);
nor U14386 (N_14386,N_14099,N_14173);
and U14387 (N_14387,N_14121,N_14087);
nor U14388 (N_14388,N_14163,N_14017);
nor U14389 (N_14389,N_14100,N_14042);
or U14390 (N_14390,N_14191,N_14086);
xnor U14391 (N_14391,N_14135,N_14191);
and U14392 (N_14392,N_14148,N_14072);
xor U14393 (N_14393,N_14048,N_14083);
or U14394 (N_14394,N_14160,N_14191);
nand U14395 (N_14395,N_14041,N_14006);
xnor U14396 (N_14396,N_14124,N_14180);
or U14397 (N_14397,N_14150,N_14177);
and U14398 (N_14398,N_14049,N_14043);
nand U14399 (N_14399,N_14029,N_14106);
or U14400 (N_14400,N_14351,N_14223);
nand U14401 (N_14401,N_14346,N_14255);
or U14402 (N_14402,N_14243,N_14298);
and U14403 (N_14403,N_14284,N_14214);
and U14404 (N_14404,N_14312,N_14337);
and U14405 (N_14405,N_14279,N_14354);
and U14406 (N_14406,N_14221,N_14265);
or U14407 (N_14407,N_14382,N_14249);
nand U14408 (N_14408,N_14299,N_14210);
xor U14409 (N_14409,N_14252,N_14352);
and U14410 (N_14410,N_14256,N_14291);
nand U14411 (N_14411,N_14209,N_14343);
and U14412 (N_14412,N_14292,N_14368);
or U14413 (N_14413,N_14355,N_14363);
and U14414 (N_14414,N_14331,N_14395);
nand U14415 (N_14415,N_14272,N_14311);
nand U14416 (N_14416,N_14332,N_14396);
nor U14417 (N_14417,N_14371,N_14274);
and U14418 (N_14418,N_14342,N_14226);
xor U14419 (N_14419,N_14372,N_14309);
nor U14420 (N_14420,N_14222,N_14387);
or U14421 (N_14421,N_14360,N_14315);
or U14422 (N_14422,N_14287,N_14306);
and U14423 (N_14423,N_14217,N_14228);
or U14424 (N_14424,N_14200,N_14224);
or U14425 (N_14425,N_14348,N_14376);
and U14426 (N_14426,N_14394,N_14361);
nor U14427 (N_14427,N_14225,N_14379);
xor U14428 (N_14428,N_14257,N_14300);
nor U14429 (N_14429,N_14365,N_14369);
nor U14430 (N_14430,N_14364,N_14324);
xnor U14431 (N_14431,N_14322,N_14208);
and U14432 (N_14432,N_14310,N_14276);
xnor U14433 (N_14433,N_14325,N_14211);
and U14434 (N_14434,N_14207,N_14313);
and U14435 (N_14435,N_14233,N_14201);
xnor U14436 (N_14436,N_14218,N_14353);
nor U14437 (N_14437,N_14202,N_14333);
nor U14438 (N_14438,N_14283,N_14335);
nor U14439 (N_14439,N_14264,N_14319);
and U14440 (N_14440,N_14231,N_14307);
or U14441 (N_14441,N_14340,N_14240);
xnor U14442 (N_14442,N_14349,N_14384);
nand U14443 (N_14443,N_14334,N_14294);
or U14444 (N_14444,N_14383,N_14267);
or U14445 (N_14445,N_14273,N_14268);
xor U14446 (N_14446,N_14341,N_14316);
nand U14447 (N_14447,N_14290,N_14254);
nand U14448 (N_14448,N_14318,N_14356);
nand U14449 (N_14449,N_14280,N_14263);
xor U14450 (N_14450,N_14358,N_14362);
or U14451 (N_14451,N_14314,N_14339);
or U14452 (N_14452,N_14288,N_14237);
nor U14453 (N_14453,N_14326,N_14238);
nand U14454 (N_14454,N_14370,N_14212);
nand U14455 (N_14455,N_14293,N_14388);
and U14456 (N_14456,N_14245,N_14282);
xor U14457 (N_14457,N_14269,N_14305);
and U14458 (N_14458,N_14251,N_14385);
xor U14459 (N_14459,N_14328,N_14205);
xor U14460 (N_14460,N_14236,N_14277);
nor U14461 (N_14461,N_14390,N_14247);
and U14462 (N_14462,N_14206,N_14248);
nor U14463 (N_14463,N_14330,N_14345);
xor U14464 (N_14464,N_14239,N_14281);
and U14465 (N_14465,N_14278,N_14304);
nand U14466 (N_14466,N_14344,N_14338);
xor U14467 (N_14467,N_14232,N_14301);
xor U14468 (N_14468,N_14297,N_14270);
xor U14469 (N_14469,N_14289,N_14253);
and U14470 (N_14470,N_14359,N_14317);
and U14471 (N_14471,N_14374,N_14302);
and U14472 (N_14472,N_14398,N_14320);
nor U14473 (N_14473,N_14336,N_14286);
xor U14474 (N_14474,N_14327,N_14399);
nand U14475 (N_14475,N_14242,N_14392);
nand U14476 (N_14476,N_14244,N_14380);
or U14477 (N_14477,N_14381,N_14308);
nor U14478 (N_14478,N_14227,N_14261);
or U14479 (N_14479,N_14258,N_14295);
xor U14480 (N_14480,N_14389,N_14241);
nand U14481 (N_14481,N_14235,N_14397);
or U14482 (N_14482,N_14321,N_14323);
and U14483 (N_14483,N_14377,N_14250);
nor U14484 (N_14484,N_14220,N_14386);
xor U14485 (N_14485,N_14391,N_14234);
or U14486 (N_14486,N_14204,N_14229);
nor U14487 (N_14487,N_14275,N_14329);
nand U14488 (N_14488,N_14285,N_14259);
nand U14489 (N_14489,N_14271,N_14213);
nand U14490 (N_14490,N_14215,N_14393);
and U14491 (N_14491,N_14246,N_14366);
nand U14492 (N_14492,N_14367,N_14230);
and U14493 (N_14493,N_14216,N_14203);
xnor U14494 (N_14494,N_14262,N_14219);
and U14495 (N_14495,N_14350,N_14303);
and U14496 (N_14496,N_14373,N_14347);
xor U14497 (N_14497,N_14296,N_14260);
or U14498 (N_14498,N_14266,N_14357);
nor U14499 (N_14499,N_14378,N_14375);
nor U14500 (N_14500,N_14216,N_14362);
nor U14501 (N_14501,N_14253,N_14329);
xor U14502 (N_14502,N_14254,N_14245);
xnor U14503 (N_14503,N_14229,N_14395);
nor U14504 (N_14504,N_14363,N_14368);
nand U14505 (N_14505,N_14253,N_14255);
nor U14506 (N_14506,N_14220,N_14383);
xnor U14507 (N_14507,N_14389,N_14311);
or U14508 (N_14508,N_14249,N_14318);
or U14509 (N_14509,N_14308,N_14296);
nor U14510 (N_14510,N_14293,N_14228);
xor U14511 (N_14511,N_14229,N_14383);
nor U14512 (N_14512,N_14256,N_14255);
nand U14513 (N_14513,N_14355,N_14362);
xnor U14514 (N_14514,N_14265,N_14370);
xnor U14515 (N_14515,N_14211,N_14379);
or U14516 (N_14516,N_14371,N_14318);
and U14517 (N_14517,N_14303,N_14300);
nand U14518 (N_14518,N_14298,N_14333);
nand U14519 (N_14519,N_14240,N_14343);
and U14520 (N_14520,N_14266,N_14202);
or U14521 (N_14521,N_14313,N_14375);
nor U14522 (N_14522,N_14270,N_14203);
and U14523 (N_14523,N_14215,N_14354);
and U14524 (N_14524,N_14222,N_14258);
or U14525 (N_14525,N_14362,N_14340);
nor U14526 (N_14526,N_14215,N_14371);
nand U14527 (N_14527,N_14332,N_14261);
and U14528 (N_14528,N_14349,N_14253);
and U14529 (N_14529,N_14223,N_14230);
and U14530 (N_14530,N_14368,N_14295);
or U14531 (N_14531,N_14285,N_14228);
nor U14532 (N_14532,N_14263,N_14348);
nor U14533 (N_14533,N_14363,N_14212);
nor U14534 (N_14534,N_14373,N_14314);
nor U14535 (N_14535,N_14206,N_14294);
xor U14536 (N_14536,N_14308,N_14392);
or U14537 (N_14537,N_14308,N_14333);
or U14538 (N_14538,N_14369,N_14213);
xnor U14539 (N_14539,N_14391,N_14225);
and U14540 (N_14540,N_14214,N_14234);
xor U14541 (N_14541,N_14250,N_14331);
xnor U14542 (N_14542,N_14377,N_14399);
nor U14543 (N_14543,N_14296,N_14207);
xnor U14544 (N_14544,N_14248,N_14242);
or U14545 (N_14545,N_14357,N_14272);
nor U14546 (N_14546,N_14218,N_14204);
xnor U14547 (N_14547,N_14280,N_14232);
and U14548 (N_14548,N_14332,N_14212);
nor U14549 (N_14549,N_14295,N_14220);
xnor U14550 (N_14550,N_14354,N_14200);
and U14551 (N_14551,N_14362,N_14238);
or U14552 (N_14552,N_14334,N_14386);
nor U14553 (N_14553,N_14253,N_14241);
nor U14554 (N_14554,N_14342,N_14370);
xor U14555 (N_14555,N_14396,N_14388);
or U14556 (N_14556,N_14274,N_14395);
nor U14557 (N_14557,N_14278,N_14392);
nand U14558 (N_14558,N_14236,N_14256);
nand U14559 (N_14559,N_14393,N_14291);
or U14560 (N_14560,N_14272,N_14253);
nand U14561 (N_14561,N_14315,N_14326);
nand U14562 (N_14562,N_14292,N_14383);
xor U14563 (N_14563,N_14309,N_14277);
or U14564 (N_14564,N_14299,N_14231);
or U14565 (N_14565,N_14261,N_14247);
or U14566 (N_14566,N_14341,N_14327);
nand U14567 (N_14567,N_14311,N_14262);
xnor U14568 (N_14568,N_14335,N_14242);
xor U14569 (N_14569,N_14344,N_14326);
xnor U14570 (N_14570,N_14397,N_14341);
and U14571 (N_14571,N_14239,N_14290);
xnor U14572 (N_14572,N_14346,N_14328);
and U14573 (N_14573,N_14360,N_14393);
and U14574 (N_14574,N_14322,N_14261);
xor U14575 (N_14575,N_14265,N_14301);
xor U14576 (N_14576,N_14295,N_14354);
or U14577 (N_14577,N_14383,N_14299);
nand U14578 (N_14578,N_14276,N_14381);
or U14579 (N_14579,N_14383,N_14302);
or U14580 (N_14580,N_14248,N_14352);
nand U14581 (N_14581,N_14324,N_14367);
and U14582 (N_14582,N_14294,N_14273);
nand U14583 (N_14583,N_14394,N_14260);
nor U14584 (N_14584,N_14338,N_14316);
nor U14585 (N_14585,N_14338,N_14278);
xor U14586 (N_14586,N_14379,N_14314);
xnor U14587 (N_14587,N_14236,N_14233);
or U14588 (N_14588,N_14357,N_14244);
and U14589 (N_14589,N_14360,N_14213);
and U14590 (N_14590,N_14252,N_14254);
and U14591 (N_14591,N_14247,N_14338);
or U14592 (N_14592,N_14392,N_14399);
nor U14593 (N_14593,N_14380,N_14267);
and U14594 (N_14594,N_14214,N_14296);
xor U14595 (N_14595,N_14370,N_14363);
xnor U14596 (N_14596,N_14208,N_14366);
or U14597 (N_14597,N_14352,N_14282);
or U14598 (N_14598,N_14355,N_14341);
nor U14599 (N_14599,N_14362,N_14351);
nand U14600 (N_14600,N_14426,N_14488);
xor U14601 (N_14601,N_14535,N_14441);
nor U14602 (N_14602,N_14533,N_14512);
xor U14603 (N_14603,N_14517,N_14569);
nor U14604 (N_14604,N_14582,N_14553);
nor U14605 (N_14605,N_14585,N_14438);
or U14606 (N_14606,N_14450,N_14508);
nor U14607 (N_14607,N_14509,N_14490);
nand U14608 (N_14608,N_14458,N_14527);
xnor U14609 (N_14609,N_14465,N_14574);
xor U14610 (N_14610,N_14522,N_14462);
nand U14611 (N_14611,N_14595,N_14597);
nand U14612 (N_14612,N_14514,N_14579);
nand U14613 (N_14613,N_14416,N_14472);
nand U14614 (N_14614,N_14466,N_14463);
and U14615 (N_14615,N_14593,N_14468);
or U14616 (N_14616,N_14564,N_14496);
and U14617 (N_14617,N_14449,N_14523);
nand U14618 (N_14618,N_14550,N_14409);
or U14619 (N_14619,N_14526,N_14495);
or U14620 (N_14620,N_14407,N_14427);
and U14621 (N_14621,N_14411,N_14548);
xor U14622 (N_14622,N_14573,N_14530);
nand U14623 (N_14623,N_14413,N_14539);
nor U14624 (N_14624,N_14544,N_14455);
xnor U14625 (N_14625,N_14570,N_14581);
nand U14626 (N_14626,N_14516,N_14580);
or U14627 (N_14627,N_14474,N_14493);
or U14628 (N_14628,N_14506,N_14439);
or U14629 (N_14629,N_14524,N_14547);
or U14630 (N_14630,N_14489,N_14492);
nor U14631 (N_14631,N_14500,N_14505);
or U14632 (N_14632,N_14470,N_14446);
xor U14633 (N_14633,N_14476,N_14586);
and U14634 (N_14634,N_14520,N_14433);
and U14635 (N_14635,N_14461,N_14454);
and U14636 (N_14636,N_14442,N_14536);
or U14637 (N_14637,N_14437,N_14404);
or U14638 (N_14638,N_14546,N_14475);
nand U14639 (N_14639,N_14419,N_14594);
xor U14640 (N_14640,N_14552,N_14588);
nor U14641 (N_14641,N_14555,N_14507);
or U14642 (N_14642,N_14415,N_14567);
and U14643 (N_14643,N_14557,N_14560);
nand U14644 (N_14644,N_14592,N_14534);
xnor U14645 (N_14645,N_14525,N_14425);
nor U14646 (N_14646,N_14482,N_14484);
or U14647 (N_14647,N_14423,N_14487);
and U14648 (N_14648,N_14444,N_14478);
xnor U14649 (N_14649,N_14542,N_14518);
xnor U14650 (N_14650,N_14485,N_14531);
nand U14651 (N_14651,N_14451,N_14563);
nor U14652 (N_14652,N_14559,N_14429);
xor U14653 (N_14653,N_14504,N_14436);
nor U14654 (N_14654,N_14554,N_14453);
nand U14655 (N_14655,N_14499,N_14578);
nand U14656 (N_14656,N_14480,N_14543);
and U14657 (N_14657,N_14408,N_14587);
xnor U14658 (N_14658,N_14591,N_14410);
and U14659 (N_14659,N_14412,N_14571);
nor U14660 (N_14660,N_14558,N_14452);
xnor U14661 (N_14661,N_14448,N_14471);
xor U14662 (N_14662,N_14540,N_14417);
and U14663 (N_14663,N_14501,N_14549);
xor U14664 (N_14664,N_14434,N_14494);
nand U14665 (N_14665,N_14464,N_14460);
xnor U14666 (N_14666,N_14590,N_14421);
nor U14667 (N_14667,N_14519,N_14447);
and U14668 (N_14668,N_14503,N_14562);
and U14669 (N_14669,N_14467,N_14479);
or U14670 (N_14670,N_14575,N_14583);
and U14671 (N_14671,N_14568,N_14424);
nor U14672 (N_14672,N_14443,N_14589);
or U14673 (N_14673,N_14491,N_14406);
and U14674 (N_14674,N_14486,N_14402);
or U14675 (N_14675,N_14576,N_14561);
nor U14676 (N_14676,N_14545,N_14565);
xnor U14677 (N_14677,N_14577,N_14599);
nand U14678 (N_14678,N_14469,N_14515);
nor U14679 (N_14679,N_14498,N_14405);
or U14680 (N_14680,N_14551,N_14566);
or U14681 (N_14681,N_14529,N_14584);
or U14682 (N_14682,N_14401,N_14422);
or U14683 (N_14683,N_14414,N_14596);
nor U14684 (N_14684,N_14538,N_14420);
or U14685 (N_14685,N_14510,N_14513);
nand U14686 (N_14686,N_14477,N_14440);
xnor U14687 (N_14687,N_14456,N_14598);
xor U14688 (N_14688,N_14431,N_14572);
or U14689 (N_14689,N_14435,N_14528);
nand U14690 (N_14690,N_14483,N_14541);
or U14691 (N_14691,N_14532,N_14502);
and U14692 (N_14692,N_14497,N_14459);
or U14693 (N_14693,N_14418,N_14432);
and U14694 (N_14694,N_14445,N_14521);
nor U14695 (N_14695,N_14428,N_14556);
nand U14696 (N_14696,N_14473,N_14481);
or U14697 (N_14697,N_14511,N_14430);
nand U14698 (N_14698,N_14403,N_14457);
and U14699 (N_14699,N_14400,N_14537);
and U14700 (N_14700,N_14400,N_14547);
nand U14701 (N_14701,N_14529,N_14450);
and U14702 (N_14702,N_14584,N_14590);
nand U14703 (N_14703,N_14454,N_14550);
or U14704 (N_14704,N_14473,N_14408);
nor U14705 (N_14705,N_14585,N_14425);
xor U14706 (N_14706,N_14484,N_14458);
xnor U14707 (N_14707,N_14464,N_14417);
nor U14708 (N_14708,N_14479,N_14506);
and U14709 (N_14709,N_14494,N_14539);
nand U14710 (N_14710,N_14539,N_14553);
and U14711 (N_14711,N_14521,N_14547);
nor U14712 (N_14712,N_14498,N_14573);
or U14713 (N_14713,N_14436,N_14499);
nand U14714 (N_14714,N_14422,N_14499);
nor U14715 (N_14715,N_14448,N_14540);
and U14716 (N_14716,N_14446,N_14461);
nor U14717 (N_14717,N_14531,N_14425);
and U14718 (N_14718,N_14472,N_14482);
and U14719 (N_14719,N_14485,N_14502);
nand U14720 (N_14720,N_14548,N_14520);
or U14721 (N_14721,N_14414,N_14446);
and U14722 (N_14722,N_14443,N_14533);
or U14723 (N_14723,N_14553,N_14517);
or U14724 (N_14724,N_14404,N_14526);
nor U14725 (N_14725,N_14539,N_14569);
xor U14726 (N_14726,N_14402,N_14444);
and U14727 (N_14727,N_14409,N_14474);
and U14728 (N_14728,N_14561,N_14423);
or U14729 (N_14729,N_14460,N_14436);
or U14730 (N_14730,N_14521,N_14517);
or U14731 (N_14731,N_14587,N_14438);
nor U14732 (N_14732,N_14452,N_14531);
and U14733 (N_14733,N_14520,N_14537);
nand U14734 (N_14734,N_14451,N_14502);
nor U14735 (N_14735,N_14571,N_14595);
or U14736 (N_14736,N_14444,N_14559);
nor U14737 (N_14737,N_14481,N_14500);
nor U14738 (N_14738,N_14454,N_14539);
nand U14739 (N_14739,N_14401,N_14565);
xor U14740 (N_14740,N_14447,N_14435);
and U14741 (N_14741,N_14452,N_14453);
xor U14742 (N_14742,N_14504,N_14537);
nor U14743 (N_14743,N_14452,N_14420);
and U14744 (N_14744,N_14488,N_14445);
and U14745 (N_14745,N_14574,N_14540);
nor U14746 (N_14746,N_14408,N_14402);
xor U14747 (N_14747,N_14480,N_14577);
nand U14748 (N_14748,N_14517,N_14501);
nand U14749 (N_14749,N_14555,N_14515);
xnor U14750 (N_14750,N_14569,N_14409);
nor U14751 (N_14751,N_14569,N_14555);
or U14752 (N_14752,N_14434,N_14472);
or U14753 (N_14753,N_14443,N_14474);
nand U14754 (N_14754,N_14424,N_14531);
and U14755 (N_14755,N_14437,N_14453);
xnor U14756 (N_14756,N_14545,N_14598);
nand U14757 (N_14757,N_14438,N_14515);
nand U14758 (N_14758,N_14524,N_14563);
nand U14759 (N_14759,N_14550,N_14536);
nor U14760 (N_14760,N_14537,N_14560);
and U14761 (N_14761,N_14574,N_14412);
nand U14762 (N_14762,N_14517,N_14500);
nand U14763 (N_14763,N_14523,N_14572);
nand U14764 (N_14764,N_14472,N_14510);
nor U14765 (N_14765,N_14561,N_14441);
nor U14766 (N_14766,N_14555,N_14547);
nand U14767 (N_14767,N_14474,N_14404);
nand U14768 (N_14768,N_14564,N_14434);
nor U14769 (N_14769,N_14415,N_14420);
nor U14770 (N_14770,N_14422,N_14545);
and U14771 (N_14771,N_14464,N_14527);
and U14772 (N_14772,N_14423,N_14598);
and U14773 (N_14773,N_14558,N_14568);
or U14774 (N_14774,N_14483,N_14512);
nand U14775 (N_14775,N_14568,N_14546);
xor U14776 (N_14776,N_14585,N_14494);
and U14777 (N_14777,N_14474,N_14581);
nor U14778 (N_14778,N_14465,N_14477);
and U14779 (N_14779,N_14538,N_14500);
or U14780 (N_14780,N_14551,N_14495);
nand U14781 (N_14781,N_14537,N_14442);
nor U14782 (N_14782,N_14521,N_14422);
xor U14783 (N_14783,N_14436,N_14589);
nand U14784 (N_14784,N_14484,N_14583);
nor U14785 (N_14785,N_14472,N_14418);
nor U14786 (N_14786,N_14510,N_14543);
or U14787 (N_14787,N_14403,N_14442);
nor U14788 (N_14788,N_14598,N_14532);
nand U14789 (N_14789,N_14419,N_14447);
and U14790 (N_14790,N_14482,N_14580);
or U14791 (N_14791,N_14463,N_14584);
xnor U14792 (N_14792,N_14461,N_14425);
nand U14793 (N_14793,N_14494,N_14527);
nor U14794 (N_14794,N_14406,N_14526);
and U14795 (N_14795,N_14422,N_14546);
xnor U14796 (N_14796,N_14408,N_14462);
and U14797 (N_14797,N_14431,N_14539);
and U14798 (N_14798,N_14497,N_14509);
nand U14799 (N_14799,N_14466,N_14520);
or U14800 (N_14800,N_14674,N_14600);
or U14801 (N_14801,N_14777,N_14744);
xnor U14802 (N_14802,N_14618,N_14783);
xor U14803 (N_14803,N_14773,N_14703);
nand U14804 (N_14804,N_14766,N_14743);
nor U14805 (N_14805,N_14697,N_14790);
or U14806 (N_14806,N_14740,N_14724);
or U14807 (N_14807,N_14727,N_14616);
nand U14808 (N_14808,N_14612,N_14632);
or U14809 (N_14809,N_14648,N_14673);
xor U14810 (N_14810,N_14621,N_14689);
or U14811 (N_14811,N_14643,N_14719);
nand U14812 (N_14812,N_14650,N_14736);
or U14813 (N_14813,N_14786,N_14679);
xor U14814 (N_14814,N_14717,N_14644);
nor U14815 (N_14815,N_14726,N_14631);
xor U14816 (N_14816,N_14720,N_14760);
xor U14817 (N_14817,N_14658,N_14628);
xnor U14818 (N_14818,N_14706,N_14780);
nand U14819 (N_14819,N_14793,N_14685);
and U14820 (N_14820,N_14601,N_14660);
xor U14821 (N_14821,N_14610,N_14645);
xnor U14822 (N_14822,N_14733,N_14797);
or U14823 (N_14823,N_14732,N_14707);
nand U14824 (N_14824,N_14785,N_14763);
or U14825 (N_14825,N_14620,N_14664);
nor U14826 (N_14826,N_14624,N_14655);
or U14827 (N_14827,N_14634,N_14614);
nand U14828 (N_14828,N_14756,N_14723);
xnor U14829 (N_14829,N_14782,N_14711);
or U14830 (N_14830,N_14626,N_14640);
nand U14831 (N_14831,N_14758,N_14794);
xor U14832 (N_14832,N_14677,N_14653);
xnor U14833 (N_14833,N_14613,N_14730);
nand U14834 (N_14834,N_14642,N_14770);
xor U14835 (N_14835,N_14615,N_14608);
nor U14836 (N_14836,N_14734,N_14798);
and U14837 (N_14837,N_14725,N_14622);
or U14838 (N_14838,N_14665,N_14779);
or U14839 (N_14839,N_14792,N_14709);
or U14840 (N_14840,N_14796,N_14774);
or U14841 (N_14841,N_14729,N_14752);
or U14842 (N_14842,N_14668,N_14764);
and U14843 (N_14843,N_14772,N_14789);
and U14844 (N_14844,N_14684,N_14604);
or U14845 (N_14845,N_14765,N_14741);
and U14846 (N_14846,N_14647,N_14661);
and U14847 (N_14847,N_14769,N_14676);
or U14848 (N_14848,N_14715,N_14619);
xor U14849 (N_14849,N_14651,N_14791);
nor U14850 (N_14850,N_14680,N_14635);
or U14851 (N_14851,N_14775,N_14731);
nand U14852 (N_14852,N_14605,N_14746);
xor U14853 (N_14853,N_14737,N_14754);
nor U14854 (N_14854,N_14670,N_14735);
and U14855 (N_14855,N_14639,N_14784);
or U14856 (N_14856,N_14761,N_14748);
nand U14857 (N_14857,N_14657,N_14712);
nor U14858 (N_14858,N_14662,N_14637);
or U14859 (N_14859,N_14671,N_14759);
and U14860 (N_14860,N_14700,N_14611);
and U14861 (N_14861,N_14795,N_14667);
and U14862 (N_14862,N_14698,N_14623);
nand U14863 (N_14863,N_14776,N_14630);
or U14864 (N_14864,N_14738,N_14739);
and U14865 (N_14865,N_14767,N_14755);
or U14866 (N_14866,N_14659,N_14714);
nand U14867 (N_14867,N_14708,N_14753);
xnor U14868 (N_14868,N_14778,N_14721);
nand U14869 (N_14869,N_14690,N_14749);
nor U14870 (N_14870,N_14688,N_14666);
and U14871 (N_14871,N_14636,N_14705);
and U14872 (N_14872,N_14633,N_14656);
xnor U14873 (N_14873,N_14646,N_14713);
or U14874 (N_14874,N_14602,N_14799);
and U14875 (N_14875,N_14751,N_14771);
nand U14876 (N_14876,N_14757,N_14750);
nand U14877 (N_14877,N_14625,N_14693);
nor U14878 (N_14878,N_14704,N_14694);
nand U14879 (N_14879,N_14641,N_14678);
and U14880 (N_14880,N_14728,N_14687);
nor U14881 (N_14881,N_14695,N_14669);
and U14882 (N_14882,N_14663,N_14699);
xnor U14883 (N_14883,N_14627,N_14654);
nor U14884 (N_14884,N_14617,N_14718);
or U14885 (N_14885,N_14781,N_14696);
xnor U14886 (N_14886,N_14609,N_14710);
or U14887 (N_14887,N_14603,N_14652);
nand U14888 (N_14888,N_14681,N_14691);
and U14889 (N_14889,N_14747,N_14745);
or U14890 (N_14890,N_14787,N_14606);
or U14891 (N_14891,N_14682,N_14788);
and U14892 (N_14892,N_14768,N_14638);
nand U14893 (N_14893,N_14686,N_14722);
xor U14894 (N_14894,N_14629,N_14649);
xnor U14895 (N_14895,N_14672,N_14742);
nor U14896 (N_14896,N_14675,N_14702);
nor U14897 (N_14897,N_14607,N_14683);
nor U14898 (N_14898,N_14762,N_14716);
xor U14899 (N_14899,N_14692,N_14701);
and U14900 (N_14900,N_14613,N_14621);
nor U14901 (N_14901,N_14771,N_14785);
or U14902 (N_14902,N_14715,N_14775);
and U14903 (N_14903,N_14613,N_14746);
and U14904 (N_14904,N_14785,N_14758);
nor U14905 (N_14905,N_14633,N_14626);
and U14906 (N_14906,N_14629,N_14698);
xnor U14907 (N_14907,N_14762,N_14797);
and U14908 (N_14908,N_14641,N_14675);
nand U14909 (N_14909,N_14797,N_14767);
and U14910 (N_14910,N_14643,N_14723);
or U14911 (N_14911,N_14791,N_14754);
nor U14912 (N_14912,N_14703,N_14719);
xor U14913 (N_14913,N_14725,N_14790);
nand U14914 (N_14914,N_14724,N_14692);
nand U14915 (N_14915,N_14699,N_14723);
xnor U14916 (N_14916,N_14744,N_14706);
xnor U14917 (N_14917,N_14694,N_14789);
nor U14918 (N_14918,N_14721,N_14609);
or U14919 (N_14919,N_14656,N_14622);
and U14920 (N_14920,N_14735,N_14713);
nor U14921 (N_14921,N_14709,N_14610);
xnor U14922 (N_14922,N_14788,N_14719);
xnor U14923 (N_14923,N_14734,N_14607);
nor U14924 (N_14924,N_14712,N_14771);
xnor U14925 (N_14925,N_14724,N_14664);
nand U14926 (N_14926,N_14782,N_14700);
or U14927 (N_14927,N_14609,N_14654);
or U14928 (N_14928,N_14687,N_14754);
xnor U14929 (N_14929,N_14775,N_14761);
nand U14930 (N_14930,N_14788,N_14632);
and U14931 (N_14931,N_14757,N_14615);
or U14932 (N_14932,N_14633,N_14679);
nor U14933 (N_14933,N_14709,N_14707);
and U14934 (N_14934,N_14733,N_14643);
or U14935 (N_14935,N_14753,N_14733);
and U14936 (N_14936,N_14692,N_14796);
xor U14937 (N_14937,N_14660,N_14797);
and U14938 (N_14938,N_14688,N_14761);
and U14939 (N_14939,N_14682,N_14641);
and U14940 (N_14940,N_14695,N_14658);
or U14941 (N_14941,N_14761,N_14755);
or U14942 (N_14942,N_14709,N_14680);
nor U14943 (N_14943,N_14674,N_14761);
xnor U14944 (N_14944,N_14657,N_14776);
and U14945 (N_14945,N_14702,N_14689);
nor U14946 (N_14946,N_14677,N_14691);
xor U14947 (N_14947,N_14606,N_14751);
xnor U14948 (N_14948,N_14734,N_14729);
xnor U14949 (N_14949,N_14659,N_14613);
nor U14950 (N_14950,N_14782,N_14648);
nand U14951 (N_14951,N_14627,N_14747);
nor U14952 (N_14952,N_14758,N_14698);
nor U14953 (N_14953,N_14781,N_14799);
nor U14954 (N_14954,N_14729,N_14660);
xor U14955 (N_14955,N_14696,N_14767);
nand U14956 (N_14956,N_14608,N_14673);
and U14957 (N_14957,N_14780,N_14711);
nand U14958 (N_14958,N_14759,N_14649);
and U14959 (N_14959,N_14761,N_14776);
or U14960 (N_14960,N_14764,N_14678);
or U14961 (N_14961,N_14642,N_14759);
nand U14962 (N_14962,N_14744,N_14750);
xnor U14963 (N_14963,N_14659,N_14706);
nand U14964 (N_14964,N_14669,N_14709);
nor U14965 (N_14965,N_14763,N_14639);
nand U14966 (N_14966,N_14788,N_14614);
nor U14967 (N_14967,N_14670,N_14799);
or U14968 (N_14968,N_14622,N_14713);
and U14969 (N_14969,N_14647,N_14740);
nor U14970 (N_14970,N_14749,N_14683);
xor U14971 (N_14971,N_14617,N_14662);
xnor U14972 (N_14972,N_14758,N_14632);
and U14973 (N_14973,N_14709,N_14762);
or U14974 (N_14974,N_14643,N_14710);
xor U14975 (N_14975,N_14666,N_14658);
nor U14976 (N_14976,N_14665,N_14663);
nor U14977 (N_14977,N_14669,N_14676);
nor U14978 (N_14978,N_14797,N_14684);
and U14979 (N_14979,N_14717,N_14729);
and U14980 (N_14980,N_14725,N_14779);
or U14981 (N_14981,N_14797,N_14609);
xor U14982 (N_14982,N_14699,N_14764);
and U14983 (N_14983,N_14680,N_14628);
or U14984 (N_14984,N_14713,N_14636);
xnor U14985 (N_14985,N_14675,N_14627);
and U14986 (N_14986,N_14618,N_14785);
xnor U14987 (N_14987,N_14632,N_14647);
or U14988 (N_14988,N_14712,N_14754);
nand U14989 (N_14989,N_14721,N_14668);
and U14990 (N_14990,N_14610,N_14739);
nand U14991 (N_14991,N_14680,N_14747);
xor U14992 (N_14992,N_14631,N_14759);
xnor U14993 (N_14993,N_14792,N_14670);
nor U14994 (N_14994,N_14796,N_14758);
and U14995 (N_14995,N_14674,N_14665);
nor U14996 (N_14996,N_14656,N_14729);
and U14997 (N_14997,N_14602,N_14739);
xor U14998 (N_14998,N_14727,N_14778);
and U14999 (N_14999,N_14756,N_14720);
xor UO_0 (O_0,N_14998,N_14829);
nor UO_1 (O_1,N_14802,N_14863);
and UO_2 (O_2,N_14959,N_14817);
nand UO_3 (O_3,N_14947,N_14885);
xnor UO_4 (O_4,N_14831,N_14994);
and UO_5 (O_5,N_14974,N_14826);
or UO_6 (O_6,N_14950,N_14939);
nor UO_7 (O_7,N_14805,N_14940);
or UO_8 (O_8,N_14920,N_14929);
or UO_9 (O_9,N_14874,N_14941);
and UO_10 (O_10,N_14870,N_14913);
or UO_11 (O_11,N_14978,N_14850);
xnor UO_12 (O_12,N_14967,N_14897);
nand UO_13 (O_13,N_14835,N_14993);
xor UO_14 (O_14,N_14804,N_14979);
nand UO_15 (O_15,N_14926,N_14873);
or UO_16 (O_16,N_14875,N_14975);
xor UO_17 (O_17,N_14828,N_14987);
xnor UO_18 (O_18,N_14883,N_14942);
nand UO_19 (O_19,N_14868,N_14955);
or UO_20 (O_20,N_14964,N_14958);
or UO_21 (O_21,N_14934,N_14857);
nor UO_22 (O_22,N_14945,N_14907);
nor UO_23 (O_23,N_14815,N_14818);
nor UO_24 (O_24,N_14900,N_14968);
and UO_25 (O_25,N_14984,N_14930);
nand UO_26 (O_26,N_14944,N_14887);
nand UO_27 (O_27,N_14905,N_14886);
nor UO_28 (O_28,N_14812,N_14903);
xor UO_29 (O_29,N_14898,N_14865);
xnor UO_30 (O_30,N_14827,N_14948);
nand UO_31 (O_31,N_14953,N_14973);
xnor UO_32 (O_32,N_14837,N_14952);
nor UO_33 (O_33,N_14824,N_14935);
or UO_34 (O_34,N_14919,N_14871);
or UO_35 (O_35,N_14925,N_14936);
nand UO_36 (O_36,N_14969,N_14854);
or UO_37 (O_37,N_14816,N_14943);
xor UO_38 (O_38,N_14981,N_14949);
nor UO_39 (O_39,N_14962,N_14972);
nand UO_40 (O_40,N_14983,N_14911);
and UO_41 (O_41,N_14841,N_14836);
or UO_42 (O_42,N_14877,N_14823);
and UO_43 (O_43,N_14916,N_14956);
and UO_44 (O_44,N_14808,N_14970);
nor UO_45 (O_45,N_14806,N_14932);
nor UO_46 (O_46,N_14988,N_14985);
and UO_47 (O_47,N_14928,N_14864);
xnor UO_48 (O_48,N_14996,N_14844);
and UO_49 (O_49,N_14915,N_14847);
xor UO_50 (O_50,N_14820,N_14888);
or UO_51 (O_51,N_14891,N_14822);
nor UO_52 (O_52,N_14912,N_14899);
or UO_53 (O_53,N_14963,N_14884);
nand UO_54 (O_54,N_14961,N_14980);
or UO_55 (O_55,N_14861,N_14856);
or UO_56 (O_56,N_14914,N_14890);
or UO_57 (O_57,N_14893,N_14894);
nand UO_58 (O_58,N_14990,N_14896);
nor UO_59 (O_59,N_14937,N_14908);
nor UO_60 (O_60,N_14852,N_14825);
xor UO_61 (O_61,N_14992,N_14855);
or UO_62 (O_62,N_14921,N_14946);
or UO_63 (O_63,N_14851,N_14878);
and UO_64 (O_64,N_14879,N_14830);
nor UO_65 (O_65,N_14848,N_14846);
or UO_66 (O_66,N_14923,N_14845);
or UO_67 (O_67,N_14876,N_14977);
xor UO_68 (O_68,N_14904,N_14869);
or UO_69 (O_69,N_14866,N_14811);
or UO_70 (O_70,N_14842,N_14954);
nand UO_71 (O_71,N_14976,N_14892);
nor UO_72 (O_72,N_14982,N_14924);
nand UO_73 (O_73,N_14819,N_14999);
xor UO_74 (O_74,N_14853,N_14801);
or UO_75 (O_75,N_14995,N_14849);
nand UO_76 (O_76,N_14803,N_14960);
or UO_77 (O_77,N_14991,N_14840);
nand UO_78 (O_78,N_14917,N_14989);
or UO_79 (O_79,N_14833,N_14834);
nand UO_80 (O_80,N_14927,N_14862);
or UO_81 (O_81,N_14889,N_14966);
xor UO_82 (O_82,N_14860,N_14965);
and UO_83 (O_83,N_14814,N_14843);
xnor UO_84 (O_84,N_14971,N_14902);
nand UO_85 (O_85,N_14901,N_14909);
and UO_86 (O_86,N_14986,N_14872);
or UO_87 (O_87,N_14882,N_14895);
and UO_88 (O_88,N_14957,N_14931);
or UO_89 (O_89,N_14821,N_14832);
xnor UO_90 (O_90,N_14910,N_14933);
or UO_91 (O_91,N_14810,N_14838);
nor UO_92 (O_92,N_14800,N_14922);
xor UO_93 (O_93,N_14997,N_14867);
nor UO_94 (O_94,N_14918,N_14951);
or UO_95 (O_95,N_14881,N_14858);
and UO_96 (O_96,N_14807,N_14839);
nor UO_97 (O_97,N_14938,N_14813);
xnor UO_98 (O_98,N_14906,N_14880);
nand UO_99 (O_99,N_14809,N_14859);
or UO_100 (O_100,N_14889,N_14927);
or UO_101 (O_101,N_14946,N_14977);
nand UO_102 (O_102,N_14815,N_14839);
nor UO_103 (O_103,N_14865,N_14871);
and UO_104 (O_104,N_14956,N_14989);
xnor UO_105 (O_105,N_14945,N_14802);
and UO_106 (O_106,N_14874,N_14900);
nor UO_107 (O_107,N_14814,N_14917);
nand UO_108 (O_108,N_14906,N_14951);
xor UO_109 (O_109,N_14843,N_14905);
and UO_110 (O_110,N_14863,N_14820);
nor UO_111 (O_111,N_14820,N_14887);
and UO_112 (O_112,N_14879,N_14895);
xor UO_113 (O_113,N_14819,N_14967);
or UO_114 (O_114,N_14991,N_14963);
xnor UO_115 (O_115,N_14964,N_14908);
nor UO_116 (O_116,N_14972,N_14863);
nor UO_117 (O_117,N_14995,N_14924);
nand UO_118 (O_118,N_14928,N_14965);
or UO_119 (O_119,N_14871,N_14847);
or UO_120 (O_120,N_14803,N_14846);
and UO_121 (O_121,N_14803,N_14913);
nand UO_122 (O_122,N_14804,N_14867);
nor UO_123 (O_123,N_14944,N_14980);
nand UO_124 (O_124,N_14808,N_14911);
and UO_125 (O_125,N_14979,N_14912);
nor UO_126 (O_126,N_14959,N_14857);
xnor UO_127 (O_127,N_14833,N_14826);
xor UO_128 (O_128,N_14954,N_14924);
nand UO_129 (O_129,N_14895,N_14975);
nand UO_130 (O_130,N_14977,N_14890);
nand UO_131 (O_131,N_14911,N_14849);
nor UO_132 (O_132,N_14905,N_14993);
xnor UO_133 (O_133,N_14980,N_14873);
and UO_134 (O_134,N_14862,N_14892);
xnor UO_135 (O_135,N_14895,N_14839);
nor UO_136 (O_136,N_14873,N_14936);
nand UO_137 (O_137,N_14910,N_14809);
xnor UO_138 (O_138,N_14870,N_14800);
xor UO_139 (O_139,N_14943,N_14916);
and UO_140 (O_140,N_14803,N_14897);
xor UO_141 (O_141,N_14948,N_14993);
and UO_142 (O_142,N_14853,N_14870);
or UO_143 (O_143,N_14816,N_14974);
nor UO_144 (O_144,N_14949,N_14879);
or UO_145 (O_145,N_14965,N_14951);
or UO_146 (O_146,N_14864,N_14865);
or UO_147 (O_147,N_14862,N_14934);
xor UO_148 (O_148,N_14876,N_14806);
and UO_149 (O_149,N_14952,N_14977);
nand UO_150 (O_150,N_14884,N_14920);
nand UO_151 (O_151,N_14808,N_14859);
or UO_152 (O_152,N_14881,N_14834);
or UO_153 (O_153,N_14931,N_14916);
xnor UO_154 (O_154,N_14823,N_14800);
and UO_155 (O_155,N_14917,N_14910);
xnor UO_156 (O_156,N_14882,N_14960);
nand UO_157 (O_157,N_14977,N_14879);
and UO_158 (O_158,N_14982,N_14875);
nor UO_159 (O_159,N_14891,N_14818);
and UO_160 (O_160,N_14918,N_14826);
and UO_161 (O_161,N_14834,N_14904);
and UO_162 (O_162,N_14885,N_14938);
xor UO_163 (O_163,N_14940,N_14935);
xnor UO_164 (O_164,N_14845,N_14803);
xnor UO_165 (O_165,N_14938,N_14995);
and UO_166 (O_166,N_14820,N_14912);
or UO_167 (O_167,N_14869,N_14960);
or UO_168 (O_168,N_14965,N_14840);
and UO_169 (O_169,N_14837,N_14908);
nand UO_170 (O_170,N_14954,N_14848);
nor UO_171 (O_171,N_14901,N_14867);
nor UO_172 (O_172,N_14851,N_14901);
and UO_173 (O_173,N_14946,N_14905);
nand UO_174 (O_174,N_14806,N_14990);
xnor UO_175 (O_175,N_14877,N_14863);
nor UO_176 (O_176,N_14922,N_14908);
or UO_177 (O_177,N_14887,N_14934);
xnor UO_178 (O_178,N_14809,N_14941);
xnor UO_179 (O_179,N_14907,N_14908);
and UO_180 (O_180,N_14874,N_14819);
nand UO_181 (O_181,N_14876,N_14929);
nor UO_182 (O_182,N_14953,N_14836);
nor UO_183 (O_183,N_14988,N_14948);
and UO_184 (O_184,N_14974,N_14822);
and UO_185 (O_185,N_14816,N_14991);
nor UO_186 (O_186,N_14965,N_14920);
and UO_187 (O_187,N_14897,N_14932);
nor UO_188 (O_188,N_14836,N_14939);
nor UO_189 (O_189,N_14834,N_14832);
and UO_190 (O_190,N_14920,N_14869);
xnor UO_191 (O_191,N_14994,N_14880);
nor UO_192 (O_192,N_14964,N_14894);
or UO_193 (O_193,N_14930,N_14841);
nor UO_194 (O_194,N_14836,N_14969);
xnor UO_195 (O_195,N_14871,N_14928);
and UO_196 (O_196,N_14887,N_14812);
and UO_197 (O_197,N_14827,N_14931);
nor UO_198 (O_198,N_14950,N_14853);
nor UO_199 (O_199,N_14970,N_14889);
nand UO_200 (O_200,N_14935,N_14922);
nand UO_201 (O_201,N_14807,N_14826);
or UO_202 (O_202,N_14999,N_14835);
and UO_203 (O_203,N_14867,N_14900);
and UO_204 (O_204,N_14981,N_14950);
nand UO_205 (O_205,N_14919,N_14870);
nor UO_206 (O_206,N_14971,N_14949);
or UO_207 (O_207,N_14927,N_14978);
nand UO_208 (O_208,N_14954,N_14912);
nand UO_209 (O_209,N_14963,N_14836);
nand UO_210 (O_210,N_14953,N_14965);
or UO_211 (O_211,N_14833,N_14902);
nand UO_212 (O_212,N_14988,N_14939);
or UO_213 (O_213,N_14865,N_14958);
or UO_214 (O_214,N_14855,N_14895);
xor UO_215 (O_215,N_14848,N_14975);
nor UO_216 (O_216,N_14943,N_14901);
or UO_217 (O_217,N_14949,N_14888);
nor UO_218 (O_218,N_14943,N_14893);
xnor UO_219 (O_219,N_14945,N_14884);
or UO_220 (O_220,N_14953,N_14837);
xor UO_221 (O_221,N_14928,N_14812);
and UO_222 (O_222,N_14826,N_14933);
nor UO_223 (O_223,N_14951,N_14994);
nand UO_224 (O_224,N_14952,N_14883);
xor UO_225 (O_225,N_14843,N_14946);
xor UO_226 (O_226,N_14848,N_14872);
xor UO_227 (O_227,N_14851,N_14954);
nor UO_228 (O_228,N_14897,N_14936);
nor UO_229 (O_229,N_14981,N_14935);
or UO_230 (O_230,N_14964,N_14974);
nand UO_231 (O_231,N_14812,N_14919);
and UO_232 (O_232,N_14883,N_14976);
and UO_233 (O_233,N_14854,N_14869);
and UO_234 (O_234,N_14916,N_14832);
xor UO_235 (O_235,N_14850,N_14820);
nor UO_236 (O_236,N_14800,N_14971);
xnor UO_237 (O_237,N_14848,N_14838);
nor UO_238 (O_238,N_14864,N_14953);
xor UO_239 (O_239,N_14946,N_14962);
or UO_240 (O_240,N_14959,N_14848);
or UO_241 (O_241,N_14953,N_14847);
or UO_242 (O_242,N_14874,N_14817);
nor UO_243 (O_243,N_14950,N_14847);
or UO_244 (O_244,N_14868,N_14893);
or UO_245 (O_245,N_14833,N_14866);
xor UO_246 (O_246,N_14824,N_14979);
nor UO_247 (O_247,N_14827,N_14986);
or UO_248 (O_248,N_14805,N_14806);
nand UO_249 (O_249,N_14884,N_14809);
and UO_250 (O_250,N_14858,N_14926);
xor UO_251 (O_251,N_14836,N_14993);
and UO_252 (O_252,N_14842,N_14967);
xnor UO_253 (O_253,N_14960,N_14880);
xnor UO_254 (O_254,N_14807,N_14883);
xnor UO_255 (O_255,N_14860,N_14956);
and UO_256 (O_256,N_14861,N_14901);
nand UO_257 (O_257,N_14994,N_14890);
xnor UO_258 (O_258,N_14920,N_14852);
or UO_259 (O_259,N_14843,N_14803);
xor UO_260 (O_260,N_14994,N_14910);
or UO_261 (O_261,N_14893,N_14957);
or UO_262 (O_262,N_14861,N_14911);
or UO_263 (O_263,N_14956,N_14900);
nor UO_264 (O_264,N_14819,N_14886);
or UO_265 (O_265,N_14939,N_14978);
or UO_266 (O_266,N_14876,N_14956);
and UO_267 (O_267,N_14810,N_14854);
nand UO_268 (O_268,N_14836,N_14984);
xor UO_269 (O_269,N_14992,N_14953);
and UO_270 (O_270,N_14857,N_14870);
nor UO_271 (O_271,N_14898,N_14860);
xnor UO_272 (O_272,N_14985,N_14939);
and UO_273 (O_273,N_14917,N_14859);
nand UO_274 (O_274,N_14998,N_14958);
and UO_275 (O_275,N_14988,N_14995);
nand UO_276 (O_276,N_14804,N_14987);
nand UO_277 (O_277,N_14850,N_14930);
nor UO_278 (O_278,N_14881,N_14806);
nand UO_279 (O_279,N_14871,N_14897);
nand UO_280 (O_280,N_14946,N_14901);
xnor UO_281 (O_281,N_14915,N_14813);
nor UO_282 (O_282,N_14947,N_14875);
nand UO_283 (O_283,N_14891,N_14916);
xnor UO_284 (O_284,N_14991,N_14813);
nor UO_285 (O_285,N_14886,N_14937);
or UO_286 (O_286,N_14892,N_14888);
or UO_287 (O_287,N_14830,N_14969);
xnor UO_288 (O_288,N_14830,N_14806);
xor UO_289 (O_289,N_14987,N_14884);
and UO_290 (O_290,N_14870,N_14910);
xnor UO_291 (O_291,N_14841,N_14824);
xnor UO_292 (O_292,N_14936,N_14877);
nand UO_293 (O_293,N_14883,N_14814);
xnor UO_294 (O_294,N_14922,N_14984);
or UO_295 (O_295,N_14824,N_14998);
xnor UO_296 (O_296,N_14805,N_14916);
and UO_297 (O_297,N_14883,N_14902);
xor UO_298 (O_298,N_14868,N_14947);
nand UO_299 (O_299,N_14853,N_14840);
or UO_300 (O_300,N_14974,N_14812);
or UO_301 (O_301,N_14887,N_14957);
and UO_302 (O_302,N_14853,N_14999);
nand UO_303 (O_303,N_14960,N_14949);
and UO_304 (O_304,N_14922,N_14879);
nand UO_305 (O_305,N_14938,N_14918);
nor UO_306 (O_306,N_14829,N_14830);
nand UO_307 (O_307,N_14949,N_14896);
nand UO_308 (O_308,N_14945,N_14843);
or UO_309 (O_309,N_14902,N_14932);
nand UO_310 (O_310,N_14834,N_14836);
nand UO_311 (O_311,N_14850,N_14875);
xor UO_312 (O_312,N_14969,N_14951);
or UO_313 (O_313,N_14935,N_14977);
xnor UO_314 (O_314,N_14893,N_14933);
or UO_315 (O_315,N_14885,N_14848);
nand UO_316 (O_316,N_14834,N_14988);
xor UO_317 (O_317,N_14940,N_14807);
or UO_318 (O_318,N_14865,N_14980);
or UO_319 (O_319,N_14961,N_14989);
nor UO_320 (O_320,N_14925,N_14859);
or UO_321 (O_321,N_14884,N_14867);
xor UO_322 (O_322,N_14897,N_14920);
nand UO_323 (O_323,N_14931,N_14917);
nand UO_324 (O_324,N_14859,N_14982);
xor UO_325 (O_325,N_14952,N_14894);
and UO_326 (O_326,N_14872,N_14915);
or UO_327 (O_327,N_14914,N_14897);
nor UO_328 (O_328,N_14979,N_14950);
and UO_329 (O_329,N_14852,N_14936);
or UO_330 (O_330,N_14905,N_14987);
xor UO_331 (O_331,N_14953,N_14842);
nand UO_332 (O_332,N_14815,N_14973);
nand UO_333 (O_333,N_14955,N_14968);
nor UO_334 (O_334,N_14969,N_14806);
or UO_335 (O_335,N_14878,N_14978);
nand UO_336 (O_336,N_14891,N_14957);
xnor UO_337 (O_337,N_14958,N_14876);
nor UO_338 (O_338,N_14819,N_14806);
and UO_339 (O_339,N_14864,N_14917);
or UO_340 (O_340,N_14863,N_14801);
xor UO_341 (O_341,N_14944,N_14886);
and UO_342 (O_342,N_14974,N_14830);
xor UO_343 (O_343,N_14803,N_14837);
or UO_344 (O_344,N_14920,N_14874);
and UO_345 (O_345,N_14959,N_14926);
nor UO_346 (O_346,N_14867,N_14976);
nand UO_347 (O_347,N_14830,N_14912);
or UO_348 (O_348,N_14945,N_14881);
and UO_349 (O_349,N_14809,N_14866);
or UO_350 (O_350,N_14859,N_14942);
xor UO_351 (O_351,N_14914,N_14830);
or UO_352 (O_352,N_14993,N_14808);
and UO_353 (O_353,N_14822,N_14857);
and UO_354 (O_354,N_14824,N_14969);
nor UO_355 (O_355,N_14907,N_14836);
nand UO_356 (O_356,N_14882,N_14857);
and UO_357 (O_357,N_14993,N_14887);
or UO_358 (O_358,N_14968,N_14920);
or UO_359 (O_359,N_14928,N_14866);
xnor UO_360 (O_360,N_14817,N_14989);
nand UO_361 (O_361,N_14978,N_14962);
nor UO_362 (O_362,N_14976,N_14814);
or UO_363 (O_363,N_14994,N_14940);
nand UO_364 (O_364,N_14909,N_14919);
xor UO_365 (O_365,N_14953,N_14885);
xnor UO_366 (O_366,N_14992,N_14834);
nor UO_367 (O_367,N_14908,N_14880);
or UO_368 (O_368,N_14881,N_14949);
nand UO_369 (O_369,N_14892,N_14856);
nor UO_370 (O_370,N_14803,N_14860);
and UO_371 (O_371,N_14918,N_14973);
nor UO_372 (O_372,N_14815,N_14989);
and UO_373 (O_373,N_14851,N_14875);
xnor UO_374 (O_374,N_14811,N_14809);
nor UO_375 (O_375,N_14920,N_14934);
or UO_376 (O_376,N_14855,N_14982);
nor UO_377 (O_377,N_14910,N_14970);
xnor UO_378 (O_378,N_14829,N_14844);
nor UO_379 (O_379,N_14918,N_14908);
nand UO_380 (O_380,N_14883,N_14802);
and UO_381 (O_381,N_14903,N_14908);
xnor UO_382 (O_382,N_14958,N_14881);
nor UO_383 (O_383,N_14821,N_14871);
or UO_384 (O_384,N_14974,N_14859);
xnor UO_385 (O_385,N_14997,N_14946);
nand UO_386 (O_386,N_14988,N_14805);
and UO_387 (O_387,N_14814,N_14953);
xor UO_388 (O_388,N_14870,N_14824);
xor UO_389 (O_389,N_14901,N_14912);
and UO_390 (O_390,N_14965,N_14992);
or UO_391 (O_391,N_14880,N_14883);
nor UO_392 (O_392,N_14831,N_14960);
nor UO_393 (O_393,N_14969,N_14985);
nand UO_394 (O_394,N_14829,N_14988);
or UO_395 (O_395,N_14852,N_14861);
nor UO_396 (O_396,N_14836,N_14947);
or UO_397 (O_397,N_14801,N_14891);
nor UO_398 (O_398,N_14819,N_14987);
xnor UO_399 (O_399,N_14941,N_14858);
or UO_400 (O_400,N_14970,N_14842);
and UO_401 (O_401,N_14918,N_14840);
xor UO_402 (O_402,N_14841,N_14972);
nand UO_403 (O_403,N_14931,N_14818);
or UO_404 (O_404,N_14860,N_14933);
or UO_405 (O_405,N_14925,N_14894);
and UO_406 (O_406,N_14896,N_14974);
xnor UO_407 (O_407,N_14809,N_14985);
nor UO_408 (O_408,N_14992,N_14907);
xnor UO_409 (O_409,N_14988,N_14872);
nand UO_410 (O_410,N_14964,N_14981);
nor UO_411 (O_411,N_14899,N_14914);
nor UO_412 (O_412,N_14970,N_14844);
and UO_413 (O_413,N_14922,N_14824);
xor UO_414 (O_414,N_14939,N_14918);
or UO_415 (O_415,N_14812,N_14973);
nand UO_416 (O_416,N_14949,N_14959);
xor UO_417 (O_417,N_14968,N_14858);
xor UO_418 (O_418,N_14968,N_14845);
or UO_419 (O_419,N_14982,N_14936);
nand UO_420 (O_420,N_14819,N_14801);
or UO_421 (O_421,N_14994,N_14987);
nor UO_422 (O_422,N_14920,N_14961);
nor UO_423 (O_423,N_14943,N_14910);
nor UO_424 (O_424,N_14835,N_14854);
nand UO_425 (O_425,N_14975,N_14920);
xor UO_426 (O_426,N_14985,N_14927);
and UO_427 (O_427,N_14939,N_14993);
nor UO_428 (O_428,N_14800,N_14871);
xor UO_429 (O_429,N_14887,N_14866);
or UO_430 (O_430,N_14827,N_14993);
or UO_431 (O_431,N_14953,N_14987);
and UO_432 (O_432,N_14840,N_14896);
xnor UO_433 (O_433,N_14853,N_14841);
and UO_434 (O_434,N_14968,N_14936);
nand UO_435 (O_435,N_14855,N_14872);
nand UO_436 (O_436,N_14966,N_14926);
nand UO_437 (O_437,N_14898,N_14803);
nor UO_438 (O_438,N_14869,N_14998);
or UO_439 (O_439,N_14865,N_14901);
and UO_440 (O_440,N_14867,N_14934);
nand UO_441 (O_441,N_14904,N_14814);
or UO_442 (O_442,N_14994,N_14805);
xor UO_443 (O_443,N_14974,N_14951);
or UO_444 (O_444,N_14968,N_14987);
and UO_445 (O_445,N_14944,N_14851);
or UO_446 (O_446,N_14920,N_14802);
nand UO_447 (O_447,N_14959,N_14888);
or UO_448 (O_448,N_14814,N_14871);
nand UO_449 (O_449,N_14911,N_14870);
and UO_450 (O_450,N_14807,N_14987);
xor UO_451 (O_451,N_14830,N_14900);
nor UO_452 (O_452,N_14853,N_14814);
xor UO_453 (O_453,N_14904,N_14821);
nor UO_454 (O_454,N_14920,N_14989);
nand UO_455 (O_455,N_14990,N_14960);
or UO_456 (O_456,N_14903,N_14907);
and UO_457 (O_457,N_14943,N_14869);
nand UO_458 (O_458,N_14855,N_14957);
and UO_459 (O_459,N_14861,N_14971);
xor UO_460 (O_460,N_14981,N_14903);
nand UO_461 (O_461,N_14827,N_14807);
xor UO_462 (O_462,N_14898,N_14919);
nor UO_463 (O_463,N_14973,N_14986);
nor UO_464 (O_464,N_14831,N_14903);
or UO_465 (O_465,N_14820,N_14804);
nor UO_466 (O_466,N_14862,N_14818);
xnor UO_467 (O_467,N_14889,N_14900);
nor UO_468 (O_468,N_14887,N_14922);
xnor UO_469 (O_469,N_14921,N_14817);
or UO_470 (O_470,N_14841,N_14919);
nand UO_471 (O_471,N_14801,N_14945);
and UO_472 (O_472,N_14988,N_14931);
xnor UO_473 (O_473,N_14894,N_14880);
and UO_474 (O_474,N_14857,N_14864);
nand UO_475 (O_475,N_14966,N_14955);
nor UO_476 (O_476,N_14866,N_14942);
or UO_477 (O_477,N_14831,N_14969);
nor UO_478 (O_478,N_14806,N_14895);
nand UO_479 (O_479,N_14906,N_14893);
nor UO_480 (O_480,N_14845,N_14870);
nand UO_481 (O_481,N_14818,N_14804);
nor UO_482 (O_482,N_14943,N_14830);
or UO_483 (O_483,N_14910,N_14978);
and UO_484 (O_484,N_14800,N_14911);
nor UO_485 (O_485,N_14914,N_14800);
or UO_486 (O_486,N_14840,N_14852);
nand UO_487 (O_487,N_14896,N_14857);
xor UO_488 (O_488,N_14874,N_14978);
xor UO_489 (O_489,N_14933,N_14959);
xor UO_490 (O_490,N_14810,N_14900);
or UO_491 (O_491,N_14804,N_14980);
xor UO_492 (O_492,N_14961,N_14936);
nand UO_493 (O_493,N_14827,N_14884);
and UO_494 (O_494,N_14910,N_14810);
or UO_495 (O_495,N_14992,N_14806);
nor UO_496 (O_496,N_14974,N_14972);
and UO_497 (O_497,N_14960,N_14929);
or UO_498 (O_498,N_14906,N_14984);
xor UO_499 (O_499,N_14919,N_14982);
xnor UO_500 (O_500,N_14874,N_14936);
xnor UO_501 (O_501,N_14887,N_14933);
nor UO_502 (O_502,N_14836,N_14912);
or UO_503 (O_503,N_14874,N_14965);
nor UO_504 (O_504,N_14909,N_14828);
nand UO_505 (O_505,N_14821,N_14839);
or UO_506 (O_506,N_14982,N_14837);
or UO_507 (O_507,N_14869,N_14906);
or UO_508 (O_508,N_14841,N_14944);
nor UO_509 (O_509,N_14853,N_14928);
nor UO_510 (O_510,N_14819,N_14944);
xor UO_511 (O_511,N_14889,N_14934);
nor UO_512 (O_512,N_14982,N_14953);
or UO_513 (O_513,N_14905,N_14825);
xnor UO_514 (O_514,N_14833,N_14889);
and UO_515 (O_515,N_14936,N_14926);
or UO_516 (O_516,N_14891,N_14800);
nand UO_517 (O_517,N_14968,N_14977);
and UO_518 (O_518,N_14903,N_14993);
nor UO_519 (O_519,N_14848,N_14819);
nand UO_520 (O_520,N_14881,N_14857);
nand UO_521 (O_521,N_14933,N_14880);
nor UO_522 (O_522,N_14901,N_14870);
or UO_523 (O_523,N_14870,N_14947);
xnor UO_524 (O_524,N_14960,N_14847);
nand UO_525 (O_525,N_14847,N_14906);
and UO_526 (O_526,N_14805,N_14823);
and UO_527 (O_527,N_14848,N_14916);
nand UO_528 (O_528,N_14922,N_14942);
nand UO_529 (O_529,N_14840,N_14920);
nand UO_530 (O_530,N_14865,N_14881);
nor UO_531 (O_531,N_14923,N_14868);
nor UO_532 (O_532,N_14885,N_14859);
nand UO_533 (O_533,N_14857,N_14968);
nor UO_534 (O_534,N_14931,N_14987);
and UO_535 (O_535,N_14827,N_14829);
or UO_536 (O_536,N_14884,N_14847);
and UO_537 (O_537,N_14904,N_14958);
nand UO_538 (O_538,N_14872,N_14866);
xor UO_539 (O_539,N_14820,N_14962);
nand UO_540 (O_540,N_14969,N_14827);
nor UO_541 (O_541,N_14904,N_14827);
or UO_542 (O_542,N_14882,N_14896);
xor UO_543 (O_543,N_14823,N_14980);
and UO_544 (O_544,N_14905,N_14827);
nor UO_545 (O_545,N_14800,N_14903);
xnor UO_546 (O_546,N_14840,N_14960);
or UO_547 (O_547,N_14974,N_14988);
xor UO_548 (O_548,N_14945,N_14806);
xnor UO_549 (O_549,N_14851,N_14961);
or UO_550 (O_550,N_14993,N_14977);
and UO_551 (O_551,N_14916,N_14804);
or UO_552 (O_552,N_14883,N_14924);
xnor UO_553 (O_553,N_14824,N_14901);
xnor UO_554 (O_554,N_14807,N_14948);
nor UO_555 (O_555,N_14808,N_14860);
xor UO_556 (O_556,N_14822,N_14858);
or UO_557 (O_557,N_14844,N_14809);
xnor UO_558 (O_558,N_14954,N_14800);
and UO_559 (O_559,N_14895,N_14949);
xnor UO_560 (O_560,N_14809,N_14990);
xor UO_561 (O_561,N_14962,N_14981);
nor UO_562 (O_562,N_14903,N_14803);
and UO_563 (O_563,N_14839,N_14940);
xnor UO_564 (O_564,N_14884,N_14996);
or UO_565 (O_565,N_14960,N_14837);
and UO_566 (O_566,N_14933,N_14804);
or UO_567 (O_567,N_14937,N_14868);
nand UO_568 (O_568,N_14971,N_14983);
xor UO_569 (O_569,N_14866,N_14912);
and UO_570 (O_570,N_14999,N_14800);
or UO_571 (O_571,N_14814,N_14824);
or UO_572 (O_572,N_14886,N_14907);
xor UO_573 (O_573,N_14966,N_14859);
nand UO_574 (O_574,N_14818,N_14995);
or UO_575 (O_575,N_14856,N_14936);
and UO_576 (O_576,N_14949,N_14884);
nand UO_577 (O_577,N_14839,N_14992);
nand UO_578 (O_578,N_14932,N_14802);
nand UO_579 (O_579,N_14898,N_14808);
nand UO_580 (O_580,N_14882,N_14934);
nor UO_581 (O_581,N_14983,N_14845);
or UO_582 (O_582,N_14822,N_14958);
nor UO_583 (O_583,N_14869,N_14863);
or UO_584 (O_584,N_14952,N_14947);
nand UO_585 (O_585,N_14917,N_14962);
or UO_586 (O_586,N_14893,N_14854);
or UO_587 (O_587,N_14933,N_14955);
or UO_588 (O_588,N_14975,N_14829);
or UO_589 (O_589,N_14830,N_14857);
or UO_590 (O_590,N_14860,N_14901);
xnor UO_591 (O_591,N_14882,N_14863);
or UO_592 (O_592,N_14827,N_14854);
or UO_593 (O_593,N_14824,N_14990);
or UO_594 (O_594,N_14852,N_14890);
xnor UO_595 (O_595,N_14853,N_14990);
or UO_596 (O_596,N_14948,N_14931);
nor UO_597 (O_597,N_14822,N_14871);
xor UO_598 (O_598,N_14901,N_14833);
xnor UO_599 (O_599,N_14840,N_14949);
or UO_600 (O_600,N_14862,N_14842);
xnor UO_601 (O_601,N_14993,N_14838);
or UO_602 (O_602,N_14976,N_14873);
nand UO_603 (O_603,N_14950,N_14851);
xnor UO_604 (O_604,N_14880,N_14803);
nor UO_605 (O_605,N_14881,N_14911);
nor UO_606 (O_606,N_14978,N_14842);
xor UO_607 (O_607,N_14946,N_14961);
nand UO_608 (O_608,N_14845,N_14868);
xnor UO_609 (O_609,N_14990,N_14986);
and UO_610 (O_610,N_14879,N_14862);
and UO_611 (O_611,N_14874,N_14808);
nor UO_612 (O_612,N_14816,N_14970);
or UO_613 (O_613,N_14803,N_14874);
and UO_614 (O_614,N_14888,N_14925);
or UO_615 (O_615,N_14838,N_14817);
or UO_616 (O_616,N_14935,N_14840);
or UO_617 (O_617,N_14857,N_14852);
or UO_618 (O_618,N_14837,N_14914);
and UO_619 (O_619,N_14919,N_14875);
nand UO_620 (O_620,N_14856,N_14815);
and UO_621 (O_621,N_14883,N_14936);
xnor UO_622 (O_622,N_14984,N_14926);
and UO_623 (O_623,N_14918,N_14911);
or UO_624 (O_624,N_14939,N_14801);
or UO_625 (O_625,N_14830,N_14972);
nor UO_626 (O_626,N_14842,N_14876);
nor UO_627 (O_627,N_14884,N_14960);
nor UO_628 (O_628,N_14968,N_14892);
nand UO_629 (O_629,N_14981,N_14879);
xor UO_630 (O_630,N_14873,N_14823);
nand UO_631 (O_631,N_14959,N_14952);
or UO_632 (O_632,N_14955,N_14927);
nor UO_633 (O_633,N_14902,N_14929);
and UO_634 (O_634,N_14846,N_14874);
and UO_635 (O_635,N_14963,N_14934);
xnor UO_636 (O_636,N_14826,N_14970);
and UO_637 (O_637,N_14804,N_14911);
xor UO_638 (O_638,N_14925,N_14965);
or UO_639 (O_639,N_14934,N_14838);
and UO_640 (O_640,N_14961,N_14901);
nand UO_641 (O_641,N_14822,N_14925);
nor UO_642 (O_642,N_14859,N_14889);
nor UO_643 (O_643,N_14898,N_14825);
or UO_644 (O_644,N_14961,N_14810);
xnor UO_645 (O_645,N_14969,N_14929);
or UO_646 (O_646,N_14834,N_14855);
or UO_647 (O_647,N_14971,N_14814);
nand UO_648 (O_648,N_14801,N_14988);
xor UO_649 (O_649,N_14948,N_14842);
nor UO_650 (O_650,N_14937,N_14954);
xor UO_651 (O_651,N_14952,N_14826);
or UO_652 (O_652,N_14868,N_14997);
and UO_653 (O_653,N_14964,N_14944);
and UO_654 (O_654,N_14813,N_14914);
nand UO_655 (O_655,N_14994,N_14944);
and UO_656 (O_656,N_14849,N_14945);
or UO_657 (O_657,N_14839,N_14855);
xor UO_658 (O_658,N_14925,N_14968);
xor UO_659 (O_659,N_14920,N_14837);
xnor UO_660 (O_660,N_14890,N_14896);
nand UO_661 (O_661,N_14822,N_14988);
and UO_662 (O_662,N_14945,N_14992);
nand UO_663 (O_663,N_14944,N_14892);
and UO_664 (O_664,N_14877,N_14858);
or UO_665 (O_665,N_14980,N_14853);
nor UO_666 (O_666,N_14975,N_14909);
xor UO_667 (O_667,N_14925,N_14992);
and UO_668 (O_668,N_14898,N_14953);
or UO_669 (O_669,N_14935,N_14801);
nand UO_670 (O_670,N_14889,N_14837);
or UO_671 (O_671,N_14915,N_14851);
xnor UO_672 (O_672,N_14896,N_14997);
and UO_673 (O_673,N_14806,N_14943);
nor UO_674 (O_674,N_14963,N_14954);
xor UO_675 (O_675,N_14957,N_14825);
xor UO_676 (O_676,N_14895,N_14978);
nand UO_677 (O_677,N_14881,N_14925);
and UO_678 (O_678,N_14915,N_14929);
nor UO_679 (O_679,N_14901,N_14897);
xor UO_680 (O_680,N_14818,N_14855);
and UO_681 (O_681,N_14996,N_14864);
nor UO_682 (O_682,N_14892,N_14955);
or UO_683 (O_683,N_14813,N_14872);
nor UO_684 (O_684,N_14808,N_14842);
xor UO_685 (O_685,N_14885,N_14869);
or UO_686 (O_686,N_14840,N_14928);
or UO_687 (O_687,N_14858,N_14947);
xnor UO_688 (O_688,N_14821,N_14819);
and UO_689 (O_689,N_14872,N_14807);
or UO_690 (O_690,N_14826,N_14961);
and UO_691 (O_691,N_14977,N_14874);
xnor UO_692 (O_692,N_14856,N_14972);
nor UO_693 (O_693,N_14964,N_14848);
and UO_694 (O_694,N_14856,N_14998);
nor UO_695 (O_695,N_14921,N_14865);
and UO_696 (O_696,N_14974,N_14997);
nor UO_697 (O_697,N_14834,N_14847);
nor UO_698 (O_698,N_14880,N_14812);
xor UO_699 (O_699,N_14801,N_14949);
and UO_700 (O_700,N_14958,N_14885);
and UO_701 (O_701,N_14833,N_14809);
nand UO_702 (O_702,N_14822,N_14800);
and UO_703 (O_703,N_14895,N_14876);
or UO_704 (O_704,N_14991,N_14979);
and UO_705 (O_705,N_14988,N_14841);
nand UO_706 (O_706,N_14887,N_14825);
nand UO_707 (O_707,N_14911,N_14894);
nor UO_708 (O_708,N_14888,N_14874);
nor UO_709 (O_709,N_14922,N_14889);
nand UO_710 (O_710,N_14995,N_14983);
nor UO_711 (O_711,N_14871,N_14812);
nand UO_712 (O_712,N_14888,N_14868);
nand UO_713 (O_713,N_14820,N_14924);
nor UO_714 (O_714,N_14992,N_14899);
and UO_715 (O_715,N_14881,N_14933);
xnor UO_716 (O_716,N_14856,N_14826);
nand UO_717 (O_717,N_14885,N_14927);
and UO_718 (O_718,N_14943,N_14917);
or UO_719 (O_719,N_14927,N_14899);
nor UO_720 (O_720,N_14853,N_14874);
xor UO_721 (O_721,N_14979,N_14990);
and UO_722 (O_722,N_14929,N_14807);
or UO_723 (O_723,N_14877,N_14912);
and UO_724 (O_724,N_14865,N_14999);
and UO_725 (O_725,N_14848,N_14851);
or UO_726 (O_726,N_14924,N_14970);
nand UO_727 (O_727,N_14957,N_14831);
or UO_728 (O_728,N_14951,N_14907);
or UO_729 (O_729,N_14872,N_14970);
and UO_730 (O_730,N_14940,N_14825);
nor UO_731 (O_731,N_14811,N_14835);
xnor UO_732 (O_732,N_14917,N_14827);
or UO_733 (O_733,N_14844,N_14948);
nand UO_734 (O_734,N_14873,N_14818);
nor UO_735 (O_735,N_14801,N_14940);
and UO_736 (O_736,N_14858,N_14884);
nand UO_737 (O_737,N_14828,N_14930);
or UO_738 (O_738,N_14967,N_14862);
and UO_739 (O_739,N_14825,N_14846);
nor UO_740 (O_740,N_14847,N_14831);
nor UO_741 (O_741,N_14832,N_14809);
nand UO_742 (O_742,N_14875,N_14865);
nor UO_743 (O_743,N_14837,N_14925);
nor UO_744 (O_744,N_14901,N_14919);
nand UO_745 (O_745,N_14993,N_14829);
xor UO_746 (O_746,N_14903,N_14864);
and UO_747 (O_747,N_14886,N_14924);
and UO_748 (O_748,N_14806,N_14952);
nand UO_749 (O_749,N_14972,N_14904);
nor UO_750 (O_750,N_14946,N_14814);
nand UO_751 (O_751,N_14822,N_14830);
or UO_752 (O_752,N_14884,N_14966);
or UO_753 (O_753,N_14837,N_14831);
nand UO_754 (O_754,N_14957,N_14946);
xor UO_755 (O_755,N_14920,N_14867);
or UO_756 (O_756,N_14836,N_14858);
and UO_757 (O_757,N_14984,N_14925);
xnor UO_758 (O_758,N_14936,N_14957);
or UO_759 (O_759,N_14968,N_14846);
xnor UO_760 (O_760,N_14822,N_14850);
nor UO_761 (O_761,N_14978,N_14930);
nand UO_762 (O_762,N_14801,N_14929);
and UO_763 (O_763,N_14915,N_14805);
and UO_764 (O_764,N_14996,N_14829);
or UO_765 (O_765,N_14844,N_14937);
nand UO_766 (O_766,N_14952,N_14845);
nand UO_767 (O_767,N_14834,N_14806);
or UO_768 (O_768,N_14938,N_14896);
xnor UO_769 (O_769,N_14949,N_14923);
nor UO_770 (O_770,N_14828,N_14912);
nand UO_771 (O_771,N_14898,N_14908);
xor UO_772 (O_772,N_14964,N_14851);
nand UO_773 (O_773,N_14949,N_14931);
nand UO_774 (O_774,N_14854,N_14953);
and UO_775 (O_775,N_14916,N_14901);
or UO_776 (O_776,N_14945,N_14915);
and UO_777 (O_777,N_14917,N_14887);
and UO_778 (O_778,N_14999,N_14816);
and UO_779 (O_779,N_14842,N_14975);
nor UO_780 (O_780,N_14955,N_14981);
nor UO_781 (O_781,N_14922,N_14832);
nor UO_782 (O_782,N_14951,N_14880);
or UO_783 (O_783,N_14892,N_14909);
and UO_784 (O_784,N_14985,N_14847);
and UO_785 (O_785,N_14972,N_14959);
nor UO_786 (O_786,N_14924,N_14969);
nor UO_787 (O_787,N_14824,N_14970);
or UO_788 (O_788,N_14832,N_14823);
and UO_789 (O_789,N_14832,N_14947);
xnor UO_790 (O_790,N_14985,N_14966);
or UO_791 (O_791,N_14877,N_14845);
or UO_792 (O_792,N_14946,N_14994);
nor UO_793 (O_793,N_14908,N_14842);
and UO_794 (O_794,N_14916,N_14864);
nor UO_795 (O_795,N_14807,N_14901);
xor UO_796 (O_796,N_14865,N_14955);
and UO_797 (O_797,N_14909,N_14861);
or UO_798 (O_798,N_14957,N_14848);
nand UO_799 (O_799,N_14881,N_14953);
xnor UO_800 (O_800,N_14887,N_14999);
xor UO_801 (O_801,N_14951,N_14890);
xor UO_802 (O_802,N_14828,N_14823);
nor UO_803 (O_803,N_14828,N_14861);
xor UO_804 (O_804,N_14819,N_14842);
nor UO_805 (O_805,N_14930,N_14866);
nand UO_806 (O_806,N_14930,N_14971);
xor UO_807 (O_807,N_14859,N_14922);
and UO_808 (O_808,N_14861,N_14831);
nand UO_809 (O_809,N_14938,N_14894);
xor UO_810 (O_810,N_14810,N_14824);
and UO_811 (O_811,N_14811,N_14970);
and UO_812 (O_812,N_14888,N_14956);
and UO_813 (O_813,N_14935,N_14886);
xnor UO_814 (O_814,N_14943,N_14968);
nor UO_815 (O_815,N_14862,N_14941);
nor UO_816 (O_816,N_14880,N_14997);
and UO_817 (O_817,N_14847,N_14974);
or UO_818 (O_818,N_14865,N_14910);
and UO_819 (O_819,N_14940,N_14972);
nor UO_820 (O_820,N_14819,N_14831);
and UO_821 (O_821,N_14867,N_14818);
and UO_822 (O_822,N_14994,N_14896);
xor UO_823 (O_823,N_14861,N_14884);
and UO_824 (O_824,N_14990,N_14888);
nor UO_825 (O_825,N_14881,N_14936);
and UO_826 (O_826,N_14968,N_14833);
xnor UO_827 (O_827,N_14832,N_14828);
xor UO_828 (O_828,N_14878,N_14893);
and UO_829 (O_829,N_14999,N_14954);
or UO_830 (O_830,N_14964,N_14895);
and UO_831 (O_831,N_14816,N_14862);
xnor UO_832 (O_832,N_14824,N_14994);
xnor UO_833 (O_833,N_14821,N_14997);
nor UO_834 (O_834,N_14837,N_14840);
or UO_835 (O_835,N_14995,N_14826);
and UO_836 (O_836,N_14907,N_14862);
or UO_837 (O_837,N_14829,N_14992);
xnor UO_838 (O_838,N_14891,N_14821);
and UO_839 (O_839,N_14824,N_14852);
or UO_840 (O_840,N_14901,N_14844);
or UO_841 (O_841,N_14834,N_14891);
nor UO_842 (O_842,N_14930,N_14988);
and UO_843 (O_843,N_14806,N_14907);
nor UO_844 (O_844,N_14950,N_14856);
nor UO_845 (O_845,N_14810,N_14985);
nor UO_846 (O_846,N_14968,N_14924);
nor UO_847 (O_847,N_14853,N_14831);
nor UO_848 (O_848,N_14893,N_14962);
or UO_849 (O_849,N_14850,N_14819);
xor UO_850 (O_850,N_14802,N_14934);
or UO_851 (O_851,N_14809,N_14852);
and UO_852 (O_852,N_14955,N_14992);
and UO_853 (O_853,N_14823,N_14875);
and UO_854 (O_854,N_14839,N_14949);
and UO_855 (O_855,N_14824,N_14820);
or UO_856 (O_856,N_14926,N_14806);
nand UO_857 (O_857,N_14900,N_14806);
nor UO_858 (O_858,N_14964,N_14917);
nand UO_859 (O_859,N_14868,N_14935);
and UO_860 (O_860,N_14874,N_14966);
xor UO_861 (O_861,N_14974,N_14983);
or UO_862 (O_862,N_14997,N_14872);
xor UO_863 (O_863,N_14810,N_14948);
nor UO_864 (O_864,N_14900,N_14925);
or UO_865 (O_865,N_14991,N_14874);
and UO_866 (O_866,N_14859,N_14860);
nand UO_867 (O_867,N_14928,N_14993);
nor UO_868 (O_868,N_14972,N_14903);
nor UO_869 (O_869,N_14890,N_14834);
xnor UO_870 (O_870,N_14977,N_14979);
nand UO_871 (O_871,N_14840,N_14819);
and UO_872 (O_872,N_14978,N_14966);
or UO_873 (O_873,N_14977,N_14831);
xnor UO_874 (O_874,N_14884,N_14946);
and UO_875 (O_875,N_14979,N_14833);
nor UO_876 (O_876,N_14801,N_14845);
nor UO_877 (O_877,N_14865,N_14959);
and UO_878 (O_878,N_14835,N_14998);
xnor UO_879 (O_879,N_14902,N_14916);
nand UO_880 (O_880,N_14916,N_14978);
nand UO_881 (O_881,N_14803,N_14926);
xor UO_882 (O_882,N_14863,N_14883);
or UO_883 (O_883,N_14934,N_14803);
and UO_884 (O_884,N_14990,N_14924);
or UO_885 (O_885,N_14985,N_14874);
nor UO_886 (O_886,N_14832,N_14950);
nand UO_887 (O_887,N_14928,N_14960);
xor UO_888 (O_888,N_14858,N_14928);
and UO_889 (O_889,N_14872,N_14965);
nor UO_890 (O_890,N_14856,N_14840);
nand UO_891 (O_891,N_14976,N_14812);
nor UO_892 (O_892,N_14862,N_14918);
nand UO_893 (O_893,N_14819,N_14876);
nand UO_894 (O_894,N_14835,N_14966);
xor UO_895 (O_895,N_14979,N_14825);
xnor UO_896 (O_896,N_14982,N_14963);
nand UO_897 (O_897,N_14866,N_14905);
nor UO_898 (O_898,N_14803,N_14850);
xor UO_899 (O_899,N_14976,N_14831);
nand UO_900 (O_900,N_14831,N_14921);
or UO_901 (O_901,N_14990,N_14883);
xnor UO_902 (O_902,N_14932,N_14998);
or UO_903 (O_903,N_14927,N_14877);
or UO_904 (O_904,N_14867,N_14835);
nand UO_905 (O_905,N_14897,N_14808);
nor UO_906 (O_906,N_14801,N_14859);
or UO_907 (O_907,N_14973,N_14808);
or UO_908 (O_908,N_14827,N_14805);
nand UO_909 (O_909,N_14833,N_14950);
or UO_910 (O_910,N_14846,N_14932);
xor UO_911 (O_911,N_14806,N_14974);
and UO_912 (O_912,N_14842,N_14806);
or UO_913 (O_913,N_14880,N_14862);
and UO_914 (O_914,N_14841,N_14960);
nand UO_915 (O_915,N_14837,N_14897);
xnor UO_916 (O_916,N_14809,N_14962);
xnor UO_917 (O_917,N_14973,N_14904);
xor UO_918 (O_918,N_14981,N_14833);
and UO_919 (O_919,N_14844,N_14961);
or UO_920 (O_920,N_14988,N_14924);
or UO_921 (O_921,N_14994,N_14806);
or UO_922 (O_922,N_14821,N_14959);
nand UO_923 (O_923,N_14947,N_14929);
and UO_924 (O_924,N_14933,N_14849);
xor UO_925 (O_925,N_14931,N_14955);
or UO_926 (O_926,N_14957,N_14939);
nor UO_927 (O_927,N_14992,N_14994);
and UO_928 (O_928,N_14960,N_14877);
and UO_929 (O_929,N_14961,N_14962);
nor UO_930 (O_930,N_14901,N_14973);
nand UO_931 (O_931,N_14884,N_14954);
nor UO_932 (O_932,N_14834,N_14903);
or UO_933 (O_933,N_14893,N_14876);
nor UO_934 (O_934,N_14913,N_14834);
nor UO_935 (O_935,N_14976,N_14846);
nand UO_936 (O_936,N_14991,N_14926);
and UO_937 (O_937,N_14956,N_14931);
and UO_938 (O_938,N_14817,N_14944);
nand UO_939 (O_939,N_14954,N_14959);
and UO_940 (O_940,N_14908,N_14818);
xor UO_941 (O_941,N_14809,N_14840);
nand UO_942 (O_942,N_14905,N_14970);
nand UO_943 (O_943,N_14974,N_14963);
nor UO_944 (O_944,N_14831,N_14965);
or UO_945 (O_945,N_14901,N_14942);
or UO_946 (O_946,N_14932,N_14820);
nand UO_947 (O_947,N_14976,N_14903);
or UO_948 (O_948,N_14912,N_14853);
nor UO_949 (O_949,N_14986,N_14968);
or UO_950 (O_950,N_14845,N_14915);
nor UO_951 (O_951,N_14829,N_14857);
nor UO_952 (O_952,N_14842,N_14919);
and UO_953 (O_953,N_14892,N_14895);
xnor UO_954 (O_954,N_14850,N_14981);
and UO_955 (O_955,N_14887,N_14880);
and UO_956 (O_956,N_14872,N_14919);
and UO_957 (O_957,N_14807,N_14860);
or UO_958 (O_958,N_14947,N_14969);
xnor UO_959 (O_959,N_14835,N_14859);
nor UO_960 (O_960,N_14995,N_14879);
or UO_961 (O_961,N_14856,N_14870);
or UO_962 (O_962,N_14974,N_14889);
nand UO_963 (O_963,N_14941,N_14900);
nand UO_964 (O_964,N_14962,N_14936);
nand UO_965 (O_965,N_14867,N_14980);
nand UO_966 (O_966,N_14917,N_14825);
or UO_967 (O_967,N_14896,N_14889);
nand UO_968 (O_968,N_14840,N_14871);
nand UO_969 (O_969,N_14845,N_14863);
nor UO_970 (O_970,N_14879,N_14811);
nor UO_971 (O_971,N_14984,N_14903);
nand UO_972 (O_972,N_14815,N_14884);
xor UO_973 (O_973,N_14845,N_14961);
nand UO_974 (O_974,N_14957,N_14802);
nor UO_975 (O_975,N_14874,N_14918);
xor UO_976 (O_976,N_14857,N_14961);
and UO_977 (O_977,N_14844,N_14853);
and UO_978 (O_978,N_14987,N_14922);
or UO_979 (O_979,N_14815,N_14881);
nand UO_980 (O_980,N_14982,N_14968);
xnor UO_981 (O_981,N_14971,N_14992);
xnor UO_982 (O_982,N_14883,N_14900);
nor UO_983 (O_983,N_14941,N_14853);
nor UO_984 (O_984,N_14992,N_14973);
and UO_985 (O_985,N_14884,N_14883);
nor UO_986 (O_986,N_14884,N_14952);
or UO_987 (O_987,N_14939,N_14967);
xnor UO_988 (O_988,N_14948,N_14815);
and UO_989 (O_989,N_14903,N_14935);
nand UO_990 (O_990,N_14919,N_14972);
nand UO_991 (O_991,N_14963,N_14808);
nand UO_992 (O_992,N_14822,N_14978);
and UO_993 (O_993,N_14946,N_14830);
nor UO_994 (O_994,N_14976,N_14943);
nor UO_995 (O_995,N_14999,N_14857);
xor UO_996 (O_996,N_14802,N_14820);
and UO_997 (O_997,N_14860,N_14904);
or UO_998 (O_998,N_14881,N_14853);
xnor UO_999 (O_999,N_14984,N_14936);
or UO_1000 (O_1000,N_14929,N_14816);
nand UO_1001 (O_1001,N_14961,N_14922);
nor UO_1002 (O_1002,N_14885,N_14892);
nand UO_1003 (O_1003,N_14968,N_14822);
or UO_1004 (O_1004,N_14815,N_14813);
nor UO_1005 (O_1005,N_14862,N_14821);
nand UO_1006 (O_1006,N_14925,N_14912);
or UO_1007 (O_1007,N_14908,N_14888);
and UO_1008 (O_1008,N_14861,N_14800);
or UO_1009 (O_1009,N_14984,N_14848);
nand UO_1010 (O_1010,N_14942,N_14819);
nor UO_1011 (O_1011,N_14999,N_14823);
xor UO_1012 (O_1012,N_14823,N_14939);
nor UO_1013 (O_1013,N_14982,N_14900);
xnor UO_1014 (O_1014,N_14910,N_14962);
nand UO_1015 (O_1015,N_14942,N_14924);
nor UO_1016 (O_1016,N_14803,N_14910);
or UO_1017 (O_1017,N_14951,N_14810);
and UO_1018 (O_1018,N_14941,N_14927);
and UO_1019 (O_1019,N_14962,N_14878);
xnor UO_1020 (O_1020,N_14834,N_14885);
and UO_1021 (O_1021,N_14984,N_14972);
nand UO_1022 (O_1022,N_14930,N_14865);
nor UO_1023 (O_1023,N_14904,N_14852);
or UO_1024 (O_1024,N_14901,N_14983);
and UO_1025 (O_1025,N_14912,N_14846);
nand UO_1026 (O_1026,N_14900,N_14923);
nand UO_1027 (O_1027,N_14996,N_14833);
nand UO_1028 (O_1028,N_14966,N_14830);
nor UO_1029 (O_1029,N_14850,N_14965);
and UO_1030 (O_1030,N_14907,N_14921);
nand UO_1031 (O_1031,N_14960,N_14926);
and UO_1032 (O_1032,N_14984,N_14941);
or UO_1033 (O_1033,N_14974,N_14858);
nand UO_1034 (O_1034,N_14896,N_14846);
xnor UO_1035 (O_1035,N_14938,N_14886);
or UO_1036 (O_1036,N_14938,N_14905);
and UO_1037 (O_1037,N_14994,N_14882);
xor UO_1038 (O_1038,N_14996,N_14983);
nor UO_1039 (O_1039,N_14820,N_14981);
nor UO_1040 (O_1040,N_14910,N_14924);
and UO_1041 (O_1041,N_14832,N_14857);
nor UO_1042 (O_1042,N_14926,N_14979);
or UO_1043 (O_1043,N_14993,N_14911);
and UO_1044 (O_1044,N_14838,N_14880);
xor UO_1045 (O_1045,N_14953,N_14861);
or UO_1046 (O_1046,N_14928,N_14956);
and UO_1047 (O_1047,N_14898,N_14922);
and UO_1048 (O_1048,N_14938,N_14971);
nand UO_1049 (O_1049,N_14956,N_14893);
and UO_1050 (O_1050,N_14935,N_14919);
xnor UO_1051 (O_1051,N_14976,N_14918);
or UO_1052 (O_1052,N_14811,N_14854);
nor UO_1053 (O_1053,N_14884,N_14956);
nor UO_1054 (O_1054,N_14962,N_14955);
or UO_1055 (O_1055,N_14932,N_14936);
nor UO_1056 (O_1056,N_14903,N_14938);
and UO_1057 (O_1057,N_14845,N_14939);
or UO_1058 (O_1058,N_14827,N_14925);
and UO_1059 (O_1059,N_14862,N_14928);
xor UO_1060 (O_1060,N_14997,N_14822);
nor UO_1061 (O_1061,N_14869,N_14884);
nand UO_1062 (O_1062,N_14972,N_14969);
xor UO_1063 (O_1063,N_14806,N_14925);
nor UO_1064 (O_1064,N_14805,N_14976);
nand UO_1065 (O_1065,N_14847,N_14817);
or UO_1066 (O_1066,N_14885,N_14997);
nor UO_1067 (O_1067,N_14879,N_14863);
nand UO_1068 (O_1068,N_14802,N_14950);
nor UO_1069 (O_1069,N_14890,N_14867);
nor UO_1070 (O_1070,N_14891,N_14995);
xnor UO_1071 (O_1071,N_14832,N_14915);
xor UO_1072 (O_1072,N_14901,N_14985);
nand UO_1073 (O_1073,N_14943,N_14948);
nand UO_1074 (O_1074,N_14836,N_14849);
and UO_1075 (O_1075,N_14844,N_14842);
nor UO_1076 (O_1076,N_14848,N_14988);
or UO_1077 (O_1077,N_14882,N_14900);
nand UO_1078 (O_1078,N_14875,N_14833);
nand UO_1079 (O_1079,N_14889,N_14800);
or UO_1080 (O_1080,N_14820,N_14868);
nand UO_1081 (O_1081,N_14890,N_14878);
nor UO_1082 (O_1082,N_14882,N_14892);
and UO_1083 (O_1083,N_14969,N_14996);
nor UO_1084 (O_1084,N_14940,N_14879);
xnor UO_1085 (O_1085,N_14912,N_14871);
and UO_1086 (O_1086,N_14869,N_14908);
or UO_1087 (O_1087,N_14876,N_14832);
xor UO_1088 (O_1088,N_14882,N_14849);
and UO_1089 (O_1089,N_14838,N_14994);
or UO_1090 (O_1090,N_14906,N_14868);
and UO_1091 (O_1091,N_14810,N_14836);
and UO_1092 (O_1092,N_14945,N_14999);
or UO_1093 (O_1093,N_14833,N_14906);
nor UO_1094 (O_1094,N_14971,N_14960);
and UO_1095 (O_1095,N_14858,N_14995);
nor UO_1096 (O_1096,N_14899,N_14806);
nor UO_1097 (O_1097,N_14922,N_14982);
nor UO_1098 (O_1098,N_14841,N_14998);
nor UO_1099 (O_1099,N_14834,N_14820);
and UO_1100 (O_1100,N_14818,N_14924);
nor UO_1101 (O_1101,N_14991,N_14896);
nor UO_1102 (O_1102,N_14811,N_14873);
nand UO_1103 (O_1103,N_14923,N_14836);
nand UO_1104 (O_1104,N_14825,N_14949);
xnor UO_1105 (O_1105,N_14819,N_14927);
or UO_1106 (O_1106,N_14822,N_14918);
xnor UO_1107 (O_1107,N_14972,N_14851);
and UO_1108 (O_1108,N_14827,N_14851);
or UO_1109 (O_1109,N_14957,N_14983);
and UO_1110 (O_1110,N_14845,N_14900);
and UO_1111 (O_1111,N_14919,N_14928);
nor UO_1112 (O_1112,N_14876,N_14847);
or UO_1113 (O_1113,N_14914,N_14848);
nor UO_1114 (O_1114,N_14858,N_14841);
xor UO_1115 (O_1115,N_14932,N_14946);
nand UO_1116 (O_1116,N_14997,N_14939);
nor UO_1117 (O_1117,N_14948,N_14859);
or UO_1118 (O_1118,N_14851,N_14899);
or UO_1119 (O_1119,N_14926,N_14983);
and UO_1120 (O_1120,N_14879,N_14963);
and UO_1121 (O_1121,N_14952,N_14925);
xnor UO_1122 (O_1122,N_14844,N_14934);
nor UO_1123 (O_1123,N_14960,N_14807);
xnor UO_1124 (O_1124,N_14947,N_14923);
xnor UO_1125 (O_1125,N_14837,N_14895);
nand UO_1126 (O_1126,N_14977,N_14943);
or UO_1127 (O_1127,N_14825,N_14858);
nor UO_1128 (O_1128,N_14932,N_14886);
nor UO_1129 (O_1129,N_14945,N_14942);
nand UO_1130 (O_1130,N_14888,N_14934);
or UO_1131 (O_1131,N_14827,N_14860);
xnor UO_1132 (O_1132,N_14880,N_14996);
nand UO_1133 (O_1133,N_14863,N_14977);
xor UO_1134 (O_1134,N_14941,N_14865);
or UO_1135 (O_1135,N_14942,N_14979);
and UO_1136 (O_1136,N_14836,N_14812);
nand UO_1137 (O_1137,N_14802,N_14933);
xnor UO_1138 (O_1138,N_14854,N_14825);
nor UO_1139 (O_1139,N_14960,N_14985);
or UO_1140 (O_1140,N_14960,N_14843);
xnor UO_1141 (O_1141,N_14812,N_14905);
or UO_1142 (O_1142,N_14987,N_14938);
xor UO_1143 (O_1143,N_14823,N_14926);
and UO_1144 (O_1144,N_14856,N_14948);
and UO_1145 (O_1145,N_14818,N_14859);
nor UO_1146 (O_1146,N_14878,N_14840);
and UO_1147 (O_1147,N_14918,N_14992);
or UO_1148 (O_1148,N_14839,N_14980);
and UO_1149 (O_1149,N_14900,N_14811);
nand UO_1150 (O_1150,N_14999,N_14858);
nand UO_1151 (O_1151,N_14941,N_14806);
and UO_1152 (O_1152,N_14860,N_14833);
nor UO_1153 (O_1153,N_14945,N_14830);
nand UO_1154 (O_1154,N_14961,N_14893);
or UO_1155 (O_1155,N_14986,N_14881);
or UO_1156 (O_1156,N_14869,N_14868);
and UO_1157 (O_1157,N_14863,N_14940);
nand UO_1158 (O_1158,N_14917,N_14861);
nand UO_1159 (O_1159,N_14978,N_14902);
xor UO_1160 (O_1160,N_14839,N_14947);
nand UO_1161 (O_1161,N_14866,N_14973);
xnor UO_1162 (O_1162,N_14988,N_14869);
nand UO_1163 (O_1163,N_14911,N_14818);
and UO_1164 (O_1164,N_14830,N_14965);
and UO_1165 (O_1165,N_14909,N_14925);
nor UO_1166 (O_1166,N_14977,N_14817);
nor UO_1167 (O_1167,N_14943,N_14889);
and UO_1168 (O_1168,N_14958,N_14875);
xor UO_1169 (O_1169,N_14887,N_14938);
and UO_1170 (O_1170,N_14859,N_14849);
and UO_1171 (O_1171,N_14876,N_14898);
nor UO_1172 (O_1172,N_14953,N_14930);
xnor UO_1173 (O_1173,N_14829,N_14927);
nor UO_1174 (O_1174,N_14973,N_14922);
xor UO_1175 (O_1175,N_14901,N_14918);
and UO_1176 (O_1176,N_14840,N_14944);
xor UO_1177 (O_1177,N_14918,N_14845);
and UO_1178 (O_1178,N_14958,N_14802);
xor UO_1179 (O_1179,N_14864,N_14808);
nor UO_1180 (O_1180,N_14881,N_14831);
and UO_1181 (O_1181,N_14991,N_14968);
nand UO_1182 (O_1182,N_14914,N_14978);
xnor UO_1183 (O_1183,N_14928,N_14804);
xnor UO_1184 (O_1184,N_14969,N_14865);
or UO_1185 (O_1185,N_14843,N_14831);
or UO_1186 (O_1186,N_14930,N_14812);
or UO_1187 (O_1187,N_14968,N_14983);
and UO_1188 (O_1188,N_14845,N_14982);
nor UO_1189 (O_1189,N_14875,N_14992);
nand UO_1190 (O_1190,N_14962,N_14862);
xnor UO_1191 (O_1191,N_14805,N_14992);
nand UO_1192 (O_1192,N_14919,N_14860);
and UO_1193 (O_1193,N_14829,N_14837);
and UO_1194 (O_1194,N_14981,N_14871);
and UO_1195 (O_1195,N_14876,N_14851);
and UO_1196 (O_1196,N_14802,N_14884);
xor UO_1197 (O_1197,N_14918,N_14813);
nor UO_1198 (O_1198,N_14837,N_14808);
or UO_1199 (O_1199,N_14801,N_14898);
xor UO_1200 (O_1200,N_14997,N_14996);
xor UO_1201 (O_1201,N_14963,N_14924);
or UO_1202 (O_1202,N_14984,N_14863);
or UO_1203 (O_1203,N_14809,N_14824);
nor UO_1204 (O_1204,N_14906,N_14908);
or UO_1205 (O_1205,N_14947,N_14895);
xnor UO_1206 (O_1206,N_14830,N_14964);
and UO_1207 (O_1207,N_14884,N_14983);
nand UO_1208 (O_1208,N_14893,N_14989);
nor UO_1209 (O_1209,N_14834,N_14980);
or UO_1210 (O_1210,N_14888,N_14932);
nor UO_1211 (O_1211,N_14896,N_14828);
and UO_1212 (O_1212,N_14929,N_14883);
nand UO_1213 (O_1213,N_14996,N_14854);
nand UO_1214 (O_1214,N_14896,N_14978);
xor UO_1215 (O_1215,N_14864,N_14968);
xnor UO_1216 (O_1216,N_14806,N_14935);
or UO_1217 (O_1217,N_14841,N_14990);
or UO_1218 (O_1218,N_14907,N_14875);
and UO_1219 (O_1219,N_14982,N_14965);
nand UO_1220 (O_1220,N_14882,N_14904);
or UO_1221 (O_1221,N_14838,N_14976);
nand UO_1222 (O_1222,N_14812,N_14897);
nor UO_1223 (O_1223,N_14861,N_14830);
or UO_1224 (O_1224,N_14827,N_14880);
or UO_1225 (O_1225,N_14932,N_14933);
nor UO_1226 (O_1226,N_14807,N_14937);
and UO_1227 (O_1227,N_14810,N_14813);
xor UO_1228 (O_1228,N_14880,N_14934);
and UO_1229 (O_1229,N_14983,N_14925);
nand UO_1230 (O_1230,N_14850,N_14945);
and UO_1231 (O_1231,N_14956,N_14817);
or UO_1232 (O_1232,N_14886,N_14828);
or UO_1233 (O_1233,N_14861,N_14976);
and UO_1234 (O_1234,N_14966,N_14829);
xnor UO_1235 (O_1235,N_14979,N_14849);
and UO_1236 (O_1236,N_14973,N_14859);
and UO_1237 (O_1237,N_14879,N_14857);
nor UO_1238 (O_1238,N_14879,N_14913);
nand UO_1239 (O_1239,N_14954,N_14895);
nor UO_1240 (O_1240,N_14901,N_14826);
and UO_1241 (O_1241,N_14919,N_14857);
nand UO_1242 (O_1242,N_14876,N_14807);
xnor UO_1243 (O_1243,N_14912,N_14913);
nor UO_1244 (O_1244,N_14826,N_14917);
or UO_1245 (O_1245,N_14862,N_14887);
xnor UO_1246 (O_1246,N_14930,N_14952);
xnor UO_1247 (O_1247,N_14873,N_14805);
or UO_1248 (O_1248,N_14907,N_14895);
nor UO_1249 (O_1249,N_14918,N_14946);
or UO_1250 (O_1250,N_14877,N_14822);
and UO_1251 (O_1251,N_14996,N_14971);
and UO_1252 (O_1252,N_14941,N_14895);
xor UO_1253 (O_1253,N_14876,N_14939);
xor UO_1254 (O_1254,N_14900,N_14816);
xnor UO_1255 (O_1255,N_14993,N_14964);
nor UO_1256 (O_1256,N_14971,N_14936);
or UO_1257 (O_1257,N_14925,N_14819);
and UO_1258 (O_1258,N_14925,N_14999);
xor UO_1259 (O_1259,N_14940,N_14859);
nand UO_1260 (O_1260,N_14835,N_14996);
and UO_1261 (O_1261,N_14817,N_14820);
or UO_1262 (O_1262,N_14873,N_14942);
xor UO_1263 (O_1263,N_14899,N_14810);
nor UO_1264 (O_1264,N_14878,N_14967);
and UO_1265 (O_1265,N_14866,N_14853);
nand UO_1266 (O_1266,N_14886,N_14823);
and UO_1267 (O_1267,N_14996,N_14963);
and UO_1268 (O_1268,N_14941,N_14916);
nand UO_1269 (O_1269,N_14886,N_14837);
or UO_1270 (O_1270,N_14967,N_14810);
and UO_1271 (O_1271,N_14875,N_14824);
xnor UO_1272 (O_1272,N_14834,N_14967);
xor UO_1273 (O_1273,N_14825,N_14958);
or UO_1274 (O_1274,N_14882,N_14983);
and UO_1275 (O_1275,N_14968,N_14835);
nand UO_1276 (O_1276,N_14975,N_14922);
nor UO_1277 (O_1277,N_14915,N_14879);
nand UO_1278 (O_1278,N_14980,N_14941);
nand UO_1279 (O_1279,N_14942,N_14947);
nand UO_1280 (O_1280,N_14879,N_14907);
nand UO_1281 (O_1281,N_14831,N_14968);
nor UO_1282 (O_1282,N_14805,N_14836);
xnor UO_1283 (O_1283,N_14914,N_14918);
nand UO_1284 (O_1284,N_14884,N_14957);
nor UO_1285 (O_1285,N_14801,N_14967);
nor UO_1286 (O_1286,N_14833,N_14891);
xor UO_1287 (O_1287,N_14933,N_14859);
nand UO_1288 (O_1288,N_14944,N_14990);
nand UO_1289 (O_1289,N_14812,N_14902);
and UO_1290 (O_1290,N_14856,N_14858);
nor UO_1291 (O_1291,N_14909,N_14903);
or UO_1292 (O_1292,N_14934,N_14859);
nand UO_1293 (O_1293,N_14979,N_14886);
and UO_1294 (O_1294,N_14995,N_14906);
nor UO_1295 (O_1295,N_14857,N_14861);
or UO_1296 (O_1296,N_14901,N_14955);
nor UO_1297 (O_1297,N_14840,N_14851);
and UO_1298 (O_1298,N_14806,N_14891);
nor UO_1299 (O_1299,N_14887,N_14953);
nand UO_1300 (O_1300,N_14960,N_14852);
or UO_1301 (O_1301,N_14821,N_14828);
or UO_1302 (O_1302,N_14944,N_14811);
and UO_1303 (O_1303,N_14850,N_14931);
nor UO_1304 (O_1304,N_14885,N_14955);
and UO_1305 (O_1305,N_14810,N_14950);
and UO_1306 (O_1306,N_14981,N_14869);
nor UO_1307 (O_1307,N_14925,N_14893);
or UO_1308 (O_1308,N_14958,N_14871);
xor UO_1309 (O_1309,N_14993,N_14946);
and UO_1310 (O_1310,N_14807,N_14809);
xor UO_1311 (O_1311,N_14896,N_14838);
and UO_1312 (O_1312,N_14945,N_14941);
nand UO_1313 (O_1313,N_14998,N_14863);
nor UO_1314 (O_1314,N_14893,N_14971);
or UO_1315 (O_1315,N_14954,N_14984);
nand UO_1316 (O_1316,N_14942,N_14990);
xor UO_1317 (O_1317,N_14800,N_14868);
xor UO_1318 (O_1318,N_14816,N_14852);
nor UO_1319 (O_1319,N_14977,N_14926);
and UO_1320 (O_1320,N_14847,N_14852);
or UO_1321 (O_1321,N_14931,N_14970);
and UO_1322 (O_1322,N_14855,N_14977);
nor UO_1323 (O_1323,N_14927,N_14935);
or UO_1324 (O_1324,N_14909,N_14880);
or UO_1325 (O_1325,N_14986,N_14802);
nor UO_1326 (O_1326,N_14847,N_14815);
nor UO_1327 (O_1327,N_14802,N_14903);
nor UO_1328 (O_1328,N_14854,N_14957);
or UO_1329 (O_1329,N_14874,N_14946);
and UO_1330 (O_1330,N_14801,N_14901);
nand UO_1331 (O_1331,N_14907,N_14844);
nor UO_1332 (O_1332,N_14916,N_14860);
or UO_1333 (O_1333,N_14896,N_14850);
xor UO_1334 (O_1334,N_14865,N_14931);
nor UO_1335 (O_1335,N_14970,N_14977);
or UO_1336 (O_1336,N_14824,N_14808);
nand UO_1337 (O_1337,N_14934,N_14915);
and UO_1338 (O_1338,N_14847,N_14982);
xor UO_1339 (O_1339,N_14999,N_14926);
and UO_1340 (O_1340,N_14964,N_14947);
or UO_1341 (O_1341,N_14932,N_14876);
nand UO_1342 (O_1342,N_14956,N_14891);
nand UO_1343 (O_1343,N_14810,N_14857);
nand UO_1344 (O_1344,N_14827,N_14846);
nor UO_1345 (O_1345,N_14863,N_14926);
nand UO_1346 (O_1346,N_14850,N_14885);
nand UO_1347 (O_1347,N_14840,N_14910);
xnor UO_1348 (O_1348,N_14834,N_14837);
and UO_1349 (O_1349,N_14858,N_14986);
xnor UO_1350 (O_1350,N_14938,N_14864);
and UO_1351 (O_1351,N_14966,N_14810);
xnor UO_1352 (O_1352,N_14822,N_14860);
xnor UO_1353 (O_1353,N_14938,N_14811);
and UO_1354 (O_1354,N_14801,N_14804);
and UO_1355 (O_1355,N_14851,N_14817);
nor UO_1356 (O_1356,N_14883,N_14882);
and UO_1357 (O_1357,N_14867,N_14837);
nand UO_1358 (O_1358,N_14929,N_14923);
or UO_1359 (O_1359,N_14896,N_14879);
and UO_1360 (O_1360,N_14952,N_14885);
nor UO_1361 (O_1361,N_14985,N_14956);
nor UO_1362 (O_1362,N_14834,N_14945);
nor UO_1363 (O_1363,N_14892,N_14891);
and UO_1364 (O_1364,N_14890,N_14963);
nand UO_1365 (O_1365,N_14811,N_14833);
and UO_1366 (O_1366,N_14954,N_14962);
nor UO_1367 (O_1367,N_14955,N_14965);
nor UO_1368 (O_1368,N_14853,N_14810);
and UO_1369 (O_1369,N_14845,N_14912);
nand UO_1370 (O_1370,N_14981,N_14849);
nand UO_1371 (O_1371,N_14818,N_14965);
or UO_1372 (O_1372,N_14992,N_14943);
or UO_1373 (O_1373,N_14971,N_14887);
and UO_1374 (O_1374,N_14992,N_14935);
or UO_1375 (O_1375,N_14845,N_14988);
nand UO_1376 (O_1376,N_14865,N_14821);
nor UO_1377 (O_1377,N_14803,N_14892);
nand UO_1378 (O_1378,N_14811,N_14877);
nand UO_1379 (O_1379,N_14880,N_14911);
nand UO_1380 (O_1380,N_14809,N_14820);
nor UO_1381 (O_1381,N_14893,N_14995);
or UO_1382 (O_1382,N_14903,N_14986);
and UO_1383 (O_1383,N_14984,N_14878);
nor UO_1384 (O_1384,N_14996,N_14988);
or UO_1385 (O_1385,N_14842,N_14937);
or UO_1386 (O_1386,N_14831,N_14991);
xnor UO_1387 (O_1387,N_14964,N_14919);
and UO_1388 (O_1388,N_14876,N_14853);
nor UO_1389 (O_1389,N_14869,N_14836);
and UO_1390 (O_1390,N_14839,N_14805);
nor UO_1391 (O_1391,N_14891,N_14910);
and UO_1392 (O_1392,N_14870,N_14973);
nand UO_1393 (O_1393,N_14878,N_14831);
or UO_1394 (O_1394,N_14963,N_14817);
nor UO_1395 (O_1395,N_14862,N_14925);
nor UO_1396 (O_1396,N_14918,N_14834);
xor UO_1397 (O_1397,N_14943,N_14851);
nor UO_1398 (O_1398,N_14920,N_14935);
nor UO_1399 (O_1399,N_14897,N_14876);
xnor UO_1400 (O_1400,N_14817,N_14939);
nand UO_1401 (O_1401,N_14958,N_14898);
nor UO_1402 (O_1402,N_14941,N_14819);
and UO_1403 (O_1403,N_14834,N_14822);
nor UO_1404 (O_1404,N_14810,N_14937);
and UO_1405 (O_1405,N_14940,N_14874);
or UO_1406 (O_1406,N_14870,N_14869);
or UO_1407 (O_1407,N_14907,N_14955);
and UO_1408 (O_1408,N_14866,N_14852);
or UO_1409 (O_1409,N_14840,N_14961);
xor UO_1410 (O_1410,N_14822,N_14980);
nand UO_1411 (O_1411,N_14819,N_14851);
and UO_1412 (O_1412,N_14896,N_14945);
xnor UO_1413 (O_1413,N_14997,N_14883);
xor UO_1414 (O_1414,N_14811,N_14838);
or UO_1415 (O_1415,N_14918,N_14814);
and UO_1416 (O_1416,N_14935,N_14936);
nand UO_1417 (O_1417,N_14904,N_14859);
or UO_1418 (O_1418,N_14976,N_14877);
and UO_1419 (O_1419,N_14980,N_14886);
nor UO_1420 (O_1420,N_14886,N_14802);
nand UO_1421 (O_1421,N_14877,N_14883);
and UO_1422 (O_1422,N_14833,N_14924);
nor UO_1423 (O_1423,N_14820,N_14988);
xnor UO_1424 (O_1424,N_14957,N_14814);
xor UO_1425 (O_1425,N_14831,N_14848);
or UO_1426 (O_1426,N_14901,N_14923);
and UO_1427 (O_1427,N_14941,N_14870);
or UO_1428 (O_1428,N_14860,N_14851);
or UO_1429 (O_1429,N_14977,N_14962);
xor UO_1430 (O_1430,N_14975,N_14933);
or UO_1431 (O_1431,N_14825,N_14921);
and UO_1432 (O_1432,N_14966,N_14933);
and UO_1433 (O_1433,N_14852,N_14962);
xor UO_1434 (O_1434,N_14992,N_14970);
nand UO_1435 (O_1435,N_14818,N_14936);
xnor UO_1436 (O_1436,N_14851,N_14890);
and UO_1437 (O_1437,N_14845,N_14916);
and UO_1438 (O_1438,N_14942,N_14958);
nor UO_1439 (O_1439,N_14955,N_14813);
and UO_1440 (O_1440,N_14923,N_14803);
and UO_1441 (O_1441,N_14974,N_14828);
nand UO_1442 (O_1442,N_14812,N_14862);
xnor UO_1443 (O_1443,N_14856,N_14963);
xnor UO_1444 (O_1444,N_14827,N_14831);
or UO_1445 (O_1445,N_14801,N_14822);
nor UO_1446 (O_1446,N_14846,N_14852);
xor UO_1447 (O_1447,N_14868,N_14864);
and UO_1448 (O_1448,N_14969,N_14801);
and UO_1449 (O_1449,N_14931,N_14857);
nor UO_1450 (O_1450,N_14873,N_14820);
or UO_1451 (O_1451,N_14940,N_14957);
or UO_1452 (O_1452,N_14964,N_14909);
and UO_1453 (O_1453,N_14915,N_14883);
and UO_1454 (O_1454,N_14842,N_14846);
or UO_1455 (O_1455,N_14998,N_14860);
nor UO_1456 (O_1456,N_14808,N_14895);
and UO_1457 (O_1457,N_14949,N_14988);
nor UO_1458 (O_1458,N_14872,N_14973);
and UO_1459 (O_1459,N_14928,N_14842);
nand UO_1460 (O_1460,N_14823,N_14820);
and UO_1461 (O_1461,N_14804,N_14937);
or UO_1462 (O_1462,N_14832,N_14964);
xor UO_1463 (O_1463,N_14928,N_14988);
nor UO_1464 (O_1464,N_14815,N_14817);
or UO_1465 (O_1465,N_14884,N_14803);
nand UO_1466 (O_1466,N_14979,N_14948);
and UO_1467 (O_1467,N_14822,N_14983);
and UO_1468 (O_1468,N_14945,N_14982);
xor UO_1469 (O_1469,N_14915,N_14904);
nor UO_1470 (O_1470,N_14947,N_14807);
or UO_1471 (O_1471,N_14950,N_14917);
or UO_1472 (O_1472,N_14806,N_14843);
and UO_1473 (O_1473,N_14912,N_14841);
nor UO_1474 (O_1474,N_14977,N_14981);
xor UO_1475 (O_1475,N_14951,N_14959);
or UO_1476 (O_1476,N_14969,N_14887);
and UO_1477 (O_1477,N_14978,N_14981);
xor UO_1478 (O_1478,N_14922,N_14891);
xor UO_1479 (O_1479,N_14861,N_14968);
and UO_1480 (O_1480,N_14805,N_14886);
or UO_1481 (O_1481,N_14908,N_14931);
xor UO_1482 (O_1482,N_14867,N_14979);
or UO_1483 (O_1483,N_14904,N_14939);
nor UO_1484 (O_1484,N_14818,N_14807);
and UO_1485 (O_1485,N_14996,N_14872);
nand UO_1486 (O_1486,N_14861,N_14863);
nand UO_1487 (O_1487,N_14848,N_14981);
nand UO_1488 (O_1488,N_14870,N_14872);
nand UO_1489 (O_1489,N_14950,N_14952);
or UO_1490 (O_1490,N_14904,N_14822);
nand UO_1491 (O_1491,N_14921,N_14944);
nand UO_1492 (O_1492,N_14821,N_14981);
and UO_1493 (O_1493,N_14957,N_14929);
nand UO_1494 (O_1494,N_14960,N_14966);
or UO_1495 (O_1495,N_14983,N_14998);
and UO_1496 (O_1496,N_14894,N_14921);
nor UO_1497 (O_1497,N_14885,N_14835);
or UO_1498 (O_1498,N_14846,N_14944);
or UO_1499 (O_1499,N_14889,N_14989);
xor UO_1500 (O_1500,N_14887,N_14921);
nor UO_1501 (O_1501,N_14953,N_14883);
xnor UO_1502 (O_1502,N_14820,N_14954);
or UO_1503 (O_1503,N_14841,N_14862);
or UO_1504 (O_1504,N_14970,N_14832);
nand UO_1505 (O_1505,N_14839,N_14847);
nor UO_1506 (O_1506,N_14867,N_14990);
or UO_1507 (O_1507,N_14976,N_14991);
or UO_1508 (O_1508,N_14857,N_14835);
nand UO_1509 (O_1509,N_14876,N_14927);
xnor UO_1510 (O_1510,N_14824,N_14906);
nand UO_1511 (O_1511,N_14896,N_14820);
xnor UO_1512 (O_1512,N_14984,N_14801);
or UO_1513 (O_1513,N_14920,N_14811);
nand UO_1514 (O_1514,N_14963,N_14854);
nand UO_1515 (O_1515,N_14869,N_14952);
nand UO_1516 (O_1516,N_14991,N_14938);
nor UO_1517 (O_1517,N_14853,N_14953);
nor UO_1518 (O_1518,N_14867,N_14811);
nor UO_1519 (O_1519,N_14985,N_14819);
or UO_1520 (O_1520,N_14958,N_14897);
nor UO_1521 (O_1521,N_14802,N_14800);
or UO_1522 (O_1522,N_14992,N_14862);
xor UO_1523 (O_1523,N_14967,N_14879);
or UO_1524 (O_1524,N_14800,N_14962);
xor UO_1525 (O_1525,N_14812,N_14918);
and UO_1526 (O_1526,N_14987,N_14989);
xor UO_1527 (O_1527,N_14893,N_14910);
xnor UO_1528 (O_1528,N_14880,N_14982);
nor UO_1529 (O_1529,N_14990,N_14919);
nand UO_1530 (O_1530,N_14959,N_14878);
xnor UO_1531 (O_1531,N_14810,N_14971);
xor UO_1532 (O_1532,N_14926,N_14935);
nand UO_1533 (O_1533,N_14808,N_14829);
nand UO_1534 (O_1534,N_14866,N_14955);
nand UO_1535 (O_1535,N_14976,N_14821);
nand UO_1536 (O_1536,N_14965,N_14964);
or UO_1537 (O_1537,N_14923,N_14938);
and UO_1538 (O_1538,N_14823,N_14810);
and UO_1539 (O_1539,N_14874,N_14887);
or UO_1540 (O_1540,N_14808,N_14949);
nand UO_1541 (O_1541,N_14831,N_14816);
xnor UO_1542 (O_1542,N_14940,N_14892);
or UO_1543 (O_1543,N_14919,N_14818);
xor UO_1544 (O_1544,N_14988,N_14978);
nor UO_1545 (O_1545,N_14928,N_14838);
and UO_1546 (O_1546,N_14894,N_14966);
or UO_1547 (O_1547,N_14858,N_14958);
and UO_1548 (O_1548,N_14941,N_14956);
nand UO_1549 (O_1549,N_14883,N_14845);
and UO_1550 (O_1550,N_14886,N_14976);
or UO_1551 (O_1551,N_14885,N_14932);
and UO_1552 (O_1552,N_14834,N_14850);
and UO_1553 (O_1553,N_14996,N_14973);
nor UO_1554 (O_1554,N_14994,N_14945);
xor UO_1555 (O_1555,N_14981,N_14918);
nor UO_1556 (O_1556,N_14921,N_14830);
nand UO_1557 (O_1557,N_14901,N_14914);
and UO_1558 (O_1558,N_14944,N_14895);
or UO_1559 (O_1559,N_14960,N_14912);
or UO_1560 (O_1560,N_14800,N_14872);
xor UO_1561 (O_1561,N_14849,N_14941);
nor UO_1562 (O_1562,N_14907,N_14861);
or UO_1563 (O_1563,N_14863,N_14955);
nand UO_1564 (O_1564,N_14965,N_14967);
xor UO_1565 (O_1565,N_14943,N_14932);
xnor UO_1566 (O_1566,N_14975,N_14849);
and UO_1567 (O_1567,N_14842,N_14882);
and UO_1568 (O_1568,N_14879,N_14831);
nor UO_1569 (O_1569,N_14909,N_14887);
xor UO_1570 (O_1570,N_14827,N_14995);
nor UO_1571 (O_1571,N_14864,N_14948);
nor UO_1572 (O_1572,N_14905,N_14864);
xnor UO_1573 (O_1573,N_14955,N_14977);
xor UO_1574 (O_1574,N_14927,N_14917);
nand UO_1575 (O_1575,N_14844,N_14827);
and UO_1576 (O_1576,N_14813,N_14954);
or UO_1577 (O_1577,N_14899,N_14976);
nand UO_1578 (O_1578,N_14852,N_14995);
xor UO_1579 (O_1579,N_14989,N_14932);
nor UO_1580 (O_1580,N_14818,N_14846);
nand UO_1581 (O_1581,N_14950,N_14983);
nor UO_1582 (O_1582,N_14885,N_14994);
and UO_1583 (O_1583,N_14976,N_14998);
xor UO_1584 (O_1584,N_14900,N_14832);
nand UO_1585 (O_1585,N_14878,N_14988);
or UO_1586 (O_1586,N_14838,N_14895);
or UO_1587 (O_1587,N_14800,N_14998);
or UO_1588 (O_1588,N_14952,N_14811);
nor UO_1589 (O_1589,N_14833,N_14940);
or UO_1590 (O_1590,N_14816,N_14849);
nor UO_1591 (O_1591,N_14987,N_14890);
xor UO_1592 (O_1592,N_14822,N_14990);
xor UO_1593 (O_1593,N_14892,N_14851);
nand UO_1594 (O_1594,N_14857,N_14840);
or UO_1595 (O_1595,N_14916,N_14982);
and UO_1596 (O_1596,N_14925,N_14874);
nor UO_1597 (O_1597,N_14817,N_14945);
nand UO_1598 (O_1598,N_14931,N_14973);
or UO_1599 (O_1599,N_14803,N_14801);
nand UO_1600 (O_1600,N_14891,N_14802);
and UO_1601 (O_1601,N_14951,N_14855);
or UO_1602 (O_1602,N_14851,N_14845);
nor UO_1603 (O_1603,N_14896,N_14969);
and UO_1604 (O_1604,N_14840,N_14957);
xor UO_1605 (O_1605,N_14935,N_14883);
nand UO_1606 (O_1606,N_14977,N_14920);
xnor UO_1607 (O_1607,N_14926,N_14940);
nand UO_1608 (O_1608,N_14827,N_14954);
nand UO_1609 (O_1609,N_14993,N_14916);
and UO_1610 (O_1610,N_14830,N_14870);
nor UO_1611 (O_1611,N_14811,N_14976);
or UO_1612 (O_1612,N_14958,N_14931);
nand UO_1613 (O_1613,N_14915,N_14931);
and UO_1614 (O_1614,N_14910,N_14909);
nor UO_1615 (O_1615,N_14831,N_14986);
xor UO_1616 (O_1616,N_14879,N_14832);
nor UO_1617 (O_1617,N_14988,N_14827);
xnor UO_1618 (O_1618,N_14910,N_14887);
nor UO_1619 (O_1619,N_14811,N_14943);
xor UO_1620 (O_1620,N_14844,N_14811);
or UO_1621 (O_1621,N_14895,N_14972);
and UO_1622 (O_1622,N_14916,N_14862);
and UO_1623 (O_1623,N_14876,N_14821);
nor UO_1624 (O_1624,N_14983,N_14993);
or UO_1625 (O_1625,N_14970,N_14936);
xor UO_1626 (O_1626,N_14852,N_14988);
and UO_1627 (O_1627,N_14998,N_14802);
xnor UO_1628 (O_1628,N_14883,N_14907);
nor UO_1629 (O_1629,N_14904,N_14802);
or UO_1630 (O_1630,N_14994,N_14852);
or UO_1631 (O_1631,N_14936,N_14954);
nor UO_1632 (O_1632,N_14895,N_14835);
nor UO_1633 (O_1633,N_14967,N_14898);
and UO_1634 (O_1634,N_14810,N_14990);
and UO_1635 (O_1635,N_14877,N_14916);
nor UO_1636 (O_1636,N_14944,N_14970);
or UO_1637 (O_1637,N_14873,N_14961);
or UO_1638 (O_1638,N_14923,N_14942);
nor UO_1639 (O_1639,N_14825,N_14847);
nand UO_1640 (O_1640,N_14982,N_14828);
nand UO_1641 (O_1641,N_14997,N_14832);
and UO_1642 (O_1642,N_14919,N_14853);
xnor UO_1643 (O_1643,N_14911,N_14934);
xnor UO_1644 (O_1644,N_14966,N_14841);
or UO_1645 (O_1645,N_14963,N_14832);
xnor UO_1646 (O_1646,N_14891,N_14816);
and UO_1647 (O_1647,N_14947,N_14837);
xor UO_1648 (O_1648,N_14847,N_14948);
xor UO_1649 (O_1649,N_14890,N_14905);
xor UO_1650 (O_1650,N_14912,N_14874);
and UO_1651 (O_1651,N_14893,N_14804);
and UO_1652 (O_1652,N_14907,N_14850);
xor UO_1653 (O_1653,N_14882,N_14954);
nand UO_1654 (O_1654,N_14839,N_14814);
or UO_1655 (O_1655,N_14884,N_14848);
xor UO_1656 (O_1656,N_14966,N_14840);
nand UO_1657 (O_1657,N_14852,N_14930);
xnor UO_1658 (O_1658,N_14808,N_14964);
xor UO_1659 (O_1659,N_14854,N_14983);
nand UO_1660 (O_1660,N_14941,N_14937);
and UO_1661 (O_1661,N_14918,N_14889);
or UO_1662 (O_1662,N_14968,N_14938);
and UO_1663 (O_1663,N_14992,N_14883);
xor UO_1664 (O_1664,N_14804,N_14917);
xor UO_1665 (O_1665,N_14960,N_14997);
nor UO_1666 (O_1666,N_14986,N_14876);
and UO_1667 (O_1667,N_14819,N_14958);
and UO_1668 (O_1668,N_14934,N_14863);
or UO_1669 (O_1669,N_14940,N_14997);
xor UO_1670 (O_1670,N_14804,N_14997);
and UO_1671 (O_1671,N_14990,N_14863);
or UO_1672 (O_1672,N_14944,N_14969);
xnor UO_1673 (O_1673,N_14927,N_14969);
and UO_1674 (O_1674,N_14900,N_14807);
nand UO_1675 (O_1675,N_14817,N_14802);
xnor UO_1676 (O_1676,N_14862,N_14834);
nor UO_1677 (O_1677,N_14879,N_14919);
and UO_1678 (O_1678,N_14867,N_14985);
nor UO_1679 (O_1679,N_14986,N_14996);
and UO_1680 (O_1680,N_14865,N_14800);
and UO_1681 (O_1681,N_14971,N_14913);
xnor UO_1682 (O_1682,N_14873,N_14968);
xor UO_1683 (O_1683,N_14967,N_14807);
nor UO_1684 (O_1684,N_14956,N_14920);
nand UO_1685 (O_1685,N_14906,N_14844);
xor UO_1686 (O_1686,N_14945,N_14853);
nand UO_1687 (O_1687,N_14838,N_14927);
and UO_1688 (O_1688,N_14898,N_14916);
and UO_1689 (O_1689,N_14825,N_14993);
nand UO_1690 (O_1690,N_14850,N_14846);
or UO_1691 (O_1691,N_14839,N_14837);
xor UO_1692 (O_1692,N_14805,N_14950);
or UO_1693 (O_1693,N_14837,N_14904);
nor UO_1694 (O_1694,N_14918,N_14871);
or UO_1695 (O_1695,N_14956,N_14909);
xor UO_1696 (O_1696,N_14955,N_14818);
nand UO_1697 (O_1697,N_14805,N_14891);
xor UO_1698 (O_1698,N_14848,N_14841);
xnor UO_1699 (O_1699,N_14801,N_14968);
and UO_1700 (O_1700,N_14857,N_14951);
or UO_1701 (O_1701,N_14949,N_14942);
nand UO_1702 (O_1702,N_14947,N_14883);
nor UO_1703 (O_1703,N_14964,N_14906);
nand UO_1704 (O_1704,N_14980,N_14905);
xnor UO_1705 (O_1705,N_14831,N_14852);
xnor UO_1706 (O_1706,N_14854,N_14855);
nand UO_1707 (O_1707,N_14803,N_14855);
or UO_1708 (O_1708,N_14806,N_14946);
nor UO_1709 (O_1709,N_14943,N_14963);
or UO_1710 (O_1710,N_14815,N_14997);
and UO_1711 (O_1711,N_14866,N_14831);
or UO_1712 (O_1712,N_14913,N_14901);
nor UO_1713 (O_1713,N_14993,N_14847);
nor UO_1714 (O_1714,N_14833,N_14971);
nor UO_1715 (O_1715,N_14879,N_14817);
nand UO_1716 (O_1716,N_14836,N_14894);
xnor UO_1717 (O_1717,N_14988,N_14885);
xnor UO_1718 (O_1718,N_14867,N_14820);
nor UO_1719 (O_1719,N_14962,N_14857);
and UO_1720 (O_1720,N_14916,N_14921);
nor UO_1721 (O_1721,N_14894,N_14878);
nor UO_1722 (O_1722,N_14837,N_14997);
and UO_1723 (O_1723,N_14886,N_14899);
nand UO_1724 (O_1724,N_14866,N_14864);
xnor UO_1725 (O_1725,N_14886,N_14955);
and UO_1726 (O_1726,N_14995,N_14864);
nand UO_1727 (O_1727,N_14834,N_14846);
nor UO_1728 (O_1728,N_14932,N_14835);
xnor UO_1729 (O_1729,N_14978,N_14856);
nand UO_1730 (O_1730,N_14840,N_14958);
or UO_1731 (O_1731,N_14919,N_14806);
nor UO_1732 (O_1732,N_14822,N_14856);
xnor UO_1733 (O_1733,N_14866,N_14914);
nand UO_1734 (O_1734,N_14994,N_14905);
nor UO_1735 (O_1735,N_14969,N_14803);
and UO_1736 (O_1736,N_14885,N_14996);
xnor UO_1737 (O_1737,N_14873,N_14958);
and UO_1738 (O_1738,N_14916,N_14834);
xor UO_1739 (O_1739,N_14908,N_14896);
and UO_1740 (O_1740,N_14904,N_14883);
or UO_1741 (O_1741,N_14946,N_14956);
xnor UO_1742 (O_1742,N_14937,N_14841);
or UO_1743 (O_1743,N_14854,N_14842);
nand UO_1744 (O_1744,N_14814,N_14995);
xnor UO_1745 (O_1745,N_14891,N_14902);
nor UO_1746 (O_1746,N_14969,N_14848);
nand UO_1747 (O_1747,N_14917,N_14991);
nor UO_1748 (O_1748,N_14906,N_14878);
xor UO_1749 (O_1749,N_14901,N_14940);
nor UO_1750 (O_1750,N_14865,N_14802);
nor UO_1751 (O_1751,N_14853,N_14846);
or UO_1752 (O_1752,N_14808,N_14972);
nor UO_1753 (O_1753,N_14835,N_14924);
nor UO_1754 (O_1754,N_14974,N_14990);
nor UO_1755 (O_1755,N_14999,N_14854);
nor UO_1756 (O_1756,N_14869,N_14819);
nand UO_1757 (O_1757,N_14978,N_14852);
and UO_1758 (O_1758,N_14921,N_14897);
or UO_1759 (O_1759,N_14865,N_14883);
nand UO_1760 (O_1760,N_14827,N_14909);
nand UO_1761 (O_1761,N_14836,N_14940);
or UO_1762 (O_1762,N_14805,N_14830);
nor UO_1763 (O_1763,N_14856,N_14951);
nand UO_1764 (O_1764,N_14865,N_14829);
and UO_1765 (O_1765,N_14928,N_14848);
and UO_1766 (O_1766,N_14892,N_14990);
nor UO_1767 (O_1767,N_14842,N_14941);
nor UO_1768 (O_1768,N_14840,N_14828);
or UO_1769 (O_1769,N_14912,N_14977);
nand UO_1770 (O_1770,N_14921,N_14977);
nor UO_1771 (O_1771,N_14893,N_14888);
nor UO_1772 (O_1772,N_14918,N_14937);
and UO_1773 (O_1773,N_14909,N_14998);
and UO_1774 (O_1774,N_14822,N_14826);
and UO_1775 (O_1775,N_14984,N_14855);
or UO_1776 (O_1776,N_14991,N_14806);
xnor UO_1777 (O_1777,N_14838,N_14826);
and UO_1778 (O_1778,N_14945,N_14968);
xnor UO_1779 (O_1779,N_14832,N_14841);
nand UO_1780 (O_1780,N_14967,N_14863);
nand UO_1781 (O_1781,N_14888,N_14972);
xnor UO_1782 (O_1782,N_14874,N_14908);
and UO_1783 (O_1783,N_14961,N_14822);
and UO_1784 (O_1784,N_14912,N_14908);
or UO_1785 (O_1785,N_14956,N_14940);
nand UO_1786 (O_1786,N_14921,N_14885);
nor UO_1787 (O_1787,N_14879,N_14824);
and UO_1788 (O_1788,N_14849,N_14893);
xor UO_1789 (O_1789,N_14997,N_14977);
or UO_1790 (O_1790,N_14904,N_14854);
or UO_1791 (O_1791,N_14992,N_14893);
xnor UO_1792 (O_1792,N_14946,N_14968);
xnor UO_1793 (O_1793,N_14971,N_14932);
and UO_1794 (O_1794,N_14888,N_14899);
or UO_1795 (O_1795,N_14825,N_14892);
or UO_1796 (O_1796,N_14913,N_14884);
nand UO_1797 (O_1797,N_14800,N_14940);
and UO_1798 (O_1798,N_14846,N_14922);
nor UO_1799 (O_1799,N_14854,N_14945);
and UO_1800 (O_1800,N_14892,N_14922);
xnor UO_1801 (O_1801,N_14818,N_14932);
nor UO_1802 (O_1802,N_14830,N_14983);
xor UO_1803 (O_1803,N_14812,N_14820);
or UO_1804 (O_1804,N_14839,N_14957);
nand UO_1805 (O_1805,N_14888,N_14906);
or UO_1806 (O_1806,N_14873,N_14846);
and UO_1807 (O_1807,N_14945,N_14815);
nand UO_1808 (O_1808,N_14859,N_14819);
nor UO_1809 (O_1809,N_14981,N_14967);
xnor UO_1810 (O_1810,N_14809,N_14928);
and UO_1811 (O_1811,N_14809,N_14912);
xor UO_1812 (O_1812,N_14875,N_14916);
nor UO_1813 (O_1813,N_14875,N_14815);
nand UO_1814 (O_1814,N_14847,N_14943);
nor UO_1815 (O_1815,N_14914,N_14851);
nor UO_1816 (O_1816,N_14853,N_14828);
nand UO_1817 (O_1817,N_14829,N_14852);
and UO_1818 (O_1818,N_14966,N_14990);
or UO_1819 (O_1819,N_14995,N_14978);
xor UO_1820 (O_1820,N_14809,N_14922);
nor UO_1821 (O_1821,N_14802,N_14949);
nor UO_1822 (O_1822,N_14809,N_14980);
nor UO_1823 (O_1823,N_14880,N_14925);
xnor UO_1824 (O_1824,N_14993,N_14839);
and UO_1825 (O_1825,N_14995,N_14897);
xnor UO_1826 (O_1826,N_14941,N_14827);
and UO_1827 (O_1827,N_14936,N_14822);
xnor UO_1828 (O_1828,N_14975,N_14955);
nor UO_1829 (O_1829,N_14986,N_14871);
xnor UO_1830 (O_1830,N_14956,N_14834);
nand UO_1831 (O_1831,N_14878,N_14879);
nand UO_1832 (O_1832,N_14838,N_14933);
and UO_1833 (O_1833,N_14951,N_14867);
or UO_1834 (O_1834,N_14803,N_14821);
or UO_1835 (O_1835,N_14820,N_14903);
nor UO_1836 (O_1836,N_14997,N_14803);
nand UO_1837 (O_1837,N_14900,N_14898);
and UO_1838 (O_1838,N_14909,N_14895);
or UO_1839 (O_1839,N_14942,N_14892);
and UO_1840 (O_1840,N_14953,N_14961);
nor UO_1841 (O_1841,N_14866,N_14983);
or UO_1842 (O_1842,N_14932,N_14844);
or UO_1843 (O_1843,N_14950,N_14966);
nor UO_1844 (O_1844,N_14800,N_14885);
and UO_1845 (O_1845,N_14990,N_14826);
and UO_1846 (O_1846,N_14869,N_14961);
or UO_1847 (O_1847,N_14810,N_14996);
or UO_1848 (O_1848,N_14926,N_14963);
nand UO_1849 (O_1849,N_14917,N_14949);
nor UO_1850 (O_1850,N_14957,N_14947);
nand UO_1851 (O_1851,N_14964,N_14883);
and UO_1852 (O_1852,N_14847,N_14921);
nor UO_1853 (O_1853,N_14987,N_14954);
nand UO_1854 (O_1854,N_14842,N_14840);
nor UO_1855 (O_1855,N_14975,N_14807);
nand UO_1856 (O_1856,N_14815,N_14891);
nand UO_1857 (O_1857,N_14998,N_14857);
nor UO_1858 (O_1858,N_14978,N_14843);
and UO_1859 (O_1859,N_14843,N_14943);
or UO_1860 (O_1860,N_14952,N_14995);
and UO_1861 (O_1861,N_14858,N_14893);
or UO_1862 (O_1862,N_14846,N_14919);
xnor UO_1863 (O_1863,N_14827,N_14804);
nand UO_1864 (O_1864,N_14856,N_14816);
xnor UO_1865 (O_1865,N_14842,N_14851);
nor UO_1866 (O_1866,N_14860,N_14853);
nand UO_1867 (O_1867,N_14953,N_14845);
and UO_1868 (O_1868,N_14958,N_14903);
xnor UO_1869 (O_1869,N_14823,N_14957);
or UO_1870 (O_1870,N_14806,N_14934);
or UO_1871 (O_1871,N_14902,N_14970);
nor UO_1872 (O_1872,N_14894,N_14932);
or UO_1873 (O_1873,N_14977,N_14885);
or UO_1874 (O_1874,N_14958,N_14801);
xnor UO_1875 (O_1875,N_14901,N_14830);
and UO_1876 (O_1876,N_14962,N_14883);
nand UO_1877 (O_1877,N_14904,N_14984);
xor UO_1878 (O_1878,N_14888,N_14819);
or UO_1879 (O_1879,N_14966,N_14809);
nand UO_1880 (O_1880,N_14831,N_14909);
and UO_1881 (O_1881,N_14913,N_14931);
or UO_1882 (O_1882,N_14805,N_14951);
or UO_1883 (O_1883,N_14884,N_14887);
nor UO_1884 (O_1884,N_14825,N_14920);
or UO_1885 (O_1885,N_14944,N_14914);
and UO_1886 (O_1886,N_14909,N_14872);
and UO_1887 (O_1887,N_14951,N_14840);
and UO_1888 (O_1888,N_14925,N_14991);
or UO_1889 (O_1889,N_14865,N_14902);
xor UO_1890 (O_1890,N_14873,N_14884);
xor UO_1891 (O_1891,N_14966,N_14938);
and UO_1892 (O_1892,N_14970,N_14981);
or UO_1893 (O_1893,N_14935,N_14871);
and UO_1894 (O_1894,N_14898,N_14986);
nand UO_1895 (O_1895,N_14936,N_14886);
nand UO_1896 (O_1896,N_14953,N_14827);
nor UO_1897 (O_1897,N_14937,N_14877);
nor UO_1898 (O_1898,N_14800,N_14852);
nand UO_1899 (O_1899,N_14934,N_14861);
nand UO_1900 (O_1900,N_14988,N_14873);
nand UO_1901 (O_1901,N_14837,N_14864);
and UO_1902 (O_1902,N_14805,N_14943);
nor UO_1903 (O_1903,N_14889,N_14994);
or UO_1904 (O_1904,N_14844,N_14893);
nand UO_1905 (O_1905,N_14972,N_14882);
or UO_1906 (O_1906,N_14800,N_14902);
nor UO_1907 (O_1907,N_14907,N_14853);
xor UO_1908 (O_1908,N_14829,N_14861);
and UO_1909 (O_1909,N_14932,N_14903);
or UO_1910 (O_1910,N_14918,N_14944);
and UO_1911 (O_1911,N_14824,N_14865);
nand UO_1912 (O_1912,N_14886,N_14985);
xor UO_1913 (O_1913,N_14999,N_14864);
nand UO_1914 (O_1914,N_14847,N_14875);
and UO_1915 (O_1915,N_14917,N_14816);
and UO_1916 (O_1916,N_14869,N_14916);
nand UO_1917 (O_1917,N_14815,N_14840);
or UO_1918 (O_1918,N_14843,N_14949);
nand UO_1919 (O_1919,N_14903,N_14871);
or UO_1920 (O_1920,N_14810,N_14945);
or UO_1921 (O_1921,N_14931,N_14909);
or UO_1922 (O_1922,N_14954,N_14885);
nand UO_1923 (O_1923,N_14949,N_14993);
or UO_1924 (O_1924,N_14826,N_14857);
xnor UO_1925 (O_1925,N_14846,N_14813);
xnor UO_1926 (O_1926,N_14948,N_14874);
or UO_1927 (O_1927,N_14999,N_14911);
or UO_1928 (O_1928,N_14813,N_14906);
nor UO_1929 (O_1929,N_14968,N_14872);
or UO_1930 (O_1930,N_14943,N_14982);
nor UO_1931 (O_1931,N_14978,N_14948);
or UO_1932 (O_1932,N_14943,N_14933);
nand UO_1933 (O_1933,N_14958,N_14905);
or UO_1934 (O_1934,N_14833,N_14808);
or UO_1935 (O_1935,N_14816,N_14867);
nand UO_1936 (O_1936,N_14871,N_14936);
xor UO_1937 (O_1937,N_14853,N_14897);
or UO_1938 (O_1938,N_14983,N_14813);
xnor UO_1939 (O_1939,N_14988,N_14955);
and UO_1940 (O_1940,N_14899,N_14903);
xor UO_1941 (O_1941,N_14855,N_14902);
nor UO_1942 (O_1942,N_14952,N_14829);
and UO_1943 (O_1943,N_14918,N_14898);
and UO_1944 (O_1944,N_14997,N_14843);
nor UO_1945 (O_1945,N_14970,N_14834);
or UO_1946 (O_1946,N_14955,N_14994);
and UO_1947 (O_1947,N_14876,N_14849);
or UO_1948 (O_1948,N_14818,N_14917);
nor UO_1949 (O_1949,N_14991,N_14939);
or UO_1950 (O_1950,N_14933,N_14993);
nand UO_1951 (O_1951,N_14867,N_14974);
nor UO_1952 (O_1952,N_14848,N_14847);
and UO_1953 (O_1953,N_14832,N_14816);
nand UO_1954 (O_1954,N_14881,N_14972);
or UO_1955 (O_1955,N_14845,N_14937);
xnor UO_1956 (O_1956,N_14801,N_14974);
nand UO_1957 (O_1957,N_14879,N_14947);
or UO_1958 (O_1958,N_14956,N_14921);
nor UO_1959 (O_1959,N_14835,N_14959);
nand UO_1960 (O_1960,N_14894,N_14998);
xor UO_1961 (O_1961,N_14930,N_14862);
nand UO_1962 (O_1962,N_14984,N_14905);
nor UO_1963 (O_1963,N_14831,N_14828);
and UO_1964 (O_1964,N_14807,N_14941);
nor UO_1965 (O_1965,N_14948,N_14846);
nand UO_1966 (O_1966,N_14857,N_14846);
and UO_1967 (O_1967,N_14996,N_14915);
nand UO_1968 (O_1968,N_14872,N_14806);
nand UO_1969 (O_1969,N_14943,N_14988);
nand UO_1970 (O_1970,N_14882,N_14862);
xor UO_1971 (O_1971,N_14822,N_14862);
and UO_1972 (O_1972,N_14954,N_14817);
nand UO_1973 (O_1973,N_14808,N_14855);
nand UO_1974 (O_1974,N_14959,N_14965);
or UO_1975 (O_1975,N_14964,N_14959);
or UO_1976 (O_1976,N_14860,N_14831);
nor UO_1977 (O_1977,N_14941,N_14999);
or UO_1978 (O_1978,N_14952,N_14896);
and UO_1979 (O_1979,N_14875,N_14929);
or UO_1980 (O_1980,N_14965,N_14854);
or UO_1981 (O_1981,N_14963,N_14875);
nor UO_1982 (O_1982,N_14865,N_14890);
xnor UO_1983 (O_1983,N_14920,N_14992);
nor UO_1984 (O_1984,N_14900,N_14906);
nor UO_1985 (O_1985,N_14929,N_14823);
nor UO_1986 (O_1986,N_14964,N_14900);
or UO_1987 (O_1987,N_14896,N_14957);
or UO_1988 (O_1988,N_14893,N_14814);
or UO_1989 (O_1989,N_14815,N_14885);
nor UO_1990 (O_1990,N_14944,N_14831);
nand UO_1991 (O_1991,N_14930,N_14945);
or UO_1992 (O_1992,N_14855,N_14877);
and UO_1993 (O_1993,N_14843,N_14941);
or UO_1994 (O_1994,N_14975,N_14904);
and UO_1995 (O_1995,N_14815,N_14878);
xnor UO_1996 (O_1996,N_14802,N_14829);
xnor UO_1997 (O_1997,N_14929,N_14903);
or UO_1998 (O_1998,N_14965,N_14849);
nor UO_1999 (O_1999,N_14840,N_14830);
endmodule