module basic_500_3000_500_15_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_44,In_294);
nor U1 (N_1,In_280,In_398);
nor U2 (N_2,In_490,In_354);
nand U3 (N_3,In_136,In_360);
and U4 (N_4,In_271,In_24);
nand U5 (N_5,In_9,In_172);
nand U6 (N_6,In_141,In_473);
nor U7 (N_7,In_322,In_69);
nand U8 (N_8,In_98,In_5);
nand U9 (N_9,In_279,In_284);
and U10 (N_10,In_337,In_492);
nor U11 (N_11,In_80,In_140);
nand U12 (N_12,In_265,In_139);
nand U13 (N_13,In_92,In_198);
nand U14 (N_14,In_157,In_384);
nor U15 (N_15,In_481,In_435);
nor U16 (N_16,In_397,In_462);
or U17 (N_17,In_361,In_247);
nand U18 (N_18,In_143,In_177);
and U19 (N_19,In_463,In_224);
nand U20 (N_20,In_132,In_425);
and U21 (N_21,In_221,In_412);
nand U22 (N_22,In_467,In_445);
nor U23 (N_23,In_328,In_63);
nor U24 (N_24,In_450,In_448);
nor U25 (N_25,In_357,In_129);
nor U26 (N_26,In_378,In_166);
or U27 (N_27,In_119,In_223);
and U28 (N_28,In_454,In_13);
nand U29 (N_29,In_417,In_308);
or U30 (N_30,In_188,In_465);
nor U31 (N_31,In_428,In_321);
nand U32 (N_32,In_174,In_444);
nor U33 (N_33,In_372,In_493);
nor U34 (N_34,In_53,In_281);
nor U35 (N_35,In_186,In_56);
nor U36 (N_36,In_408,In_289);
nand U37 (N_37,In_103,In_386);
nand U38 (N_38,In_209,In_402);
or U39 (N_39,In_31,In_218);
nand U40 (N_40,In_96,In_429);
nor U41 (N_41,In_306,In_230);
nand U42 (N_42,In_373,In_347);
or U43 (N_43,In_14,In_393);
or U44 (N_44,In_86,In_73);
and U45 (N_45,In_227,In_318);
nor U46 (N_46,In_127,In_311);
nand U47 (N_47,In_187,In_236);
or U48 (N_48,In_154,In_447);
or U49 (N_49,In_90,In_195);
nand U50 (N_50,In_210,In_240);
or U51 (N_51,In_253,In_309);
and U52 (N_52,In_11,In_142);
nand U53 (N_53,In_111,In_67);
and U54 (N_54,In_367,In_411);
nor U55 (N_55,In_81,In_72);
and U56 (N_56,In_107,In_315);
nand U57 (N_57,In_12,In_285);
or U58 (N_58,In_213,In_248);
and U59 (N_59,In_160,In_162);
nand U60 (N_60,In_304,In_194);
nand U61 (N_61,In_399,In_460);
and U62 (N_62,In_87,In_33);
nand U63 (N_63,In_388,In_28);
nor U64 (N_64,In_474,In_250);
nand U65 (N_65,In_349,In_35);
or U66 (N_66,In_327,In_482);
or U67 (N_67,In_396,In_233);
and U68 (N_68,In_257,In_254);
and U69 (N_69,In_291,In_256);
nand U70 (N_70,In_344,In_179);
or U71 (N_71,In_216,In_206);
and U72 (N_72,In_430,In_379);
and U73 (N_73,In_22,In_458);
nor U74 (N_74,In_190,In_491);
nor U75 (N_75,In_380,In_274);
and U76 (N_76,In_365,In_93);
nor U77 (N_77,In_20,In_62);
xor U78 (N_78,In_49,In_359);
and U79 (N_79,In_434,In_363);
or U80 (N_80,In_426,In_97);
nor U81 (N_81,In_243,In_152);
or U82 (N_82,In_339,In_244);
or U83 (N_83,In_32,In_150);
or U84 (N_84,In_60,In_219);
nor U85 (N_85,In_488,In_483);
or U86 (N_86,In_212,In_124);
and U87 (N_87,In_235,In_374);
nor U88 (N_88,In_25,In_433);
or U89 (N_89,In_178,In_27);
or U90 (N_90,In_346,In_217);
nand U91 (N_91,In_249,In_335);
or U92 (N_92,In_468,In_261);
or U93 (N_93,In_452,In_287);
and U94 (N_94,In_118,In_406);
nor U95 (N_95,In_196,In_76);
nor U96 (N_96,In_277,In_484);
and U97 (N_97,In_381,In_290);
or U98 (N_98,In_2,In_138);
or U99 (N_99,In_102,In_436);
nor U100 (N_100,In_211,In_158);
nor U101 (N_101,In_260,In_151);
or U102 (N_102,In_222,In_312);
xnor U103 (N_103,In_364,In_479);
and U104 (N_104,In_446,In_376);
nand U105 (N_105,In_193,In_17);
nand U106 (N_106,In_275,In_123);
and U107 (N_107,In_99,In_153);
or U108 (N_108,In_15,In_295);
nor U109 (N_109,In_342,In_299);
nor U110 (N_110,In_431,In_204);
and U111 (N_111,In_348,In_16);
or U112 (N_112,In_182,In_115);
or U113 (N_113,In_496,In_207);
nand U114 (N_114,In_173,In_355);
nand U115 (N_115,In_457,In_47);
and U116 (N_116,In_316,In_55);
and U117 (N_117,In_246,In_245);
or U118 (N_118,In_18,In_499);
or U119 (N_119,In_110,In_453);
and U120 (N_120,In_165,In_89);
nor U121 (N_121,In_34,In_241);
and U122 (N_122,In_181,In_438);
and U123 (N_123,In_4,In_362);
or U124 (N_124,In_121,In_68);
and U125 (N_125,In_470,In_325);
and U126 (N_126,In_215,In_421);
nor U127 (N_127,In_466,In_146);
nand U128 (N_128,In_113,In_175);
nor U129 (N_129,In_251,In_371);
nand U130 (N_130,In_497,In_258);
or U131 (N_131,In_8,In_432);
and U132 (N_132,In_353,In_427);
and U133 (N_133,In_148,In_391);
and U134 (N_134,In_268,In_440);
and U135 (N_135,In_341,In_390);
and U136 (N_136,In_84,In_352);
or U137 (N_137,In_338,In_155);
and U138 (N_138,In_85,In_266);
nand U139 (N_139,In_122,In_145);
nand U140 (N_140,In_486,In_487);
nand U141 (N_141,In_310,In_120);
or U142 (N_142,In_21,In_79);
nand U143 (N_143,In_292,In_133);
or U144 (N_144,In_38,In_326);
nor U145 (N_145,In_0,In_461);
nand U146 (N_146,In_340,In_65);
nor U147 (N_147,In_313,In_125);
nor U148 (N_148,In_6,In_405);
or U149 (N_149,In_377,In_104);
or U150 (N_150,In_203,In_7);
or U151 (N_151,In_392,In_305);
and U152 (N_152,In_319,In_343);
nand U153 (N_153,In_416,In_382);
and U154 (N_154,In_495,In_226);
and U155 (N_155,In_423,In_41);
and U156 (N_156,In_234,In_95);
or U157 (N_157,In_114,In_3);
and U158 (N_158,In_282,In_40);
or U159 (N_159,In_403,In_52);
nor U160 (N_160,In_419,In_191);
xnor U161 (N_161,In_54,In_51);
nand U162 (N_162,In_314,In_176);
nand U163 (N_163,In_137,In_189);
or U164 (N_164,In_164,In_451);
nor U165 (N_165,In_331,In_231);
xor U166 (N_166,In_385,In_336);
or U167 (N_167,In_37,In_401);
and U168 (N_168,In_201,In_442);
nand U169 (N_169,In_135,In_116);
and U170 (N_170,In_167,In_46);
nand U171 (N_171,In_61,In_200);
or U172 (N_172,In_267,In_498);
nand U173 (N_173,In_296,In_101);
nor U174 (N_174,In_414,In_297);
nor U175 (N_175,In_356,In_202);
nand U176 (N_176,In_131,In_420);
or U177 (N_177,In_147,In_1);
nor U178 (N_178,In_263,In_464);
nand U179 (N_179,In_43,In_437);
nand U180 (N_180,In_409,In_395);
nand U181 (N_181,In_333,In_288);
and U182 (N_182,In_273,In_170);
or U183 (N_183,In_171,In_272);
nor U184 (N_184,In_106,In_109);
and U185 (N_185,In_205,In_300);
and U186 (N_186,In_161,In_149);
and U187 (N_187,In_413,In_323);
or U188 (N_188,In_259,In_82);
and U189 (N_189,In_130,In_330);
nand U190 (N_190,In_262,In_472);
or U191 (N_191,In_30,In_293);
and U192 (N_192,In_39,In_441);
or U193 (N_193,In_459,In_220);
and U194 (N_194,In_480,In_48);
and U195 (N_195,In_485,In_302);
or U196 (N_196,In_71,In_23);
or U197 (N_197,In_94,In_351);
or U198 (N_198,In_74,In_350);
and U199 (N_199,In_475,In_208);
and U200 (N_200,N_167,N_85);
and U201 (N_201,N_13,N_173);
and U202 (N_202,N_38,N_148);
nand U203 (N_203,N_177,N_51);
nand U204 (N_204,N_46,N_144);
and U205 (N_205,In_415,N_82);
nand U206 (N_206,In_183,In_494);
or U207 (N_207,N_63,In_77);
nand U208 (N_208,In_45,In_418);
nand U209 (N_209,N_110,In_478);
and U210 (N_210,In_185,N_151);
nor U211 (N_211,In_455,N_152);
or U212 (N_212,N_59,In_232);
nor U213 (N_213,N_43,In_184);
nor U214 (N_214,N_25,In_237);
or U215 (N_215,N_37,N_27);
or U216 (N_216,N_116,In_242);
nor U217 (N_217,N_123,N_163);
nand U218 (N_218,N_128,N_5);
or U219 (N_219,In_229,N_113);
nand U220 (N_220,N_141,In_255);
nor U221 (N_221,N_90,In_320);
or U222 (N_222,N_69,N_115);
nand U223 (N_223,N_49,N_83);
or U224 (N_224,N_105,N_60);
nor U225 (N_225,In_471,In_298);
or U226 (N_226,In_78,N_181);
and U227 (N_227,In_59,N_58);
and U228 (N_228,N_176,In_180);
nor U229 (N_229,N_89,N_126);
and U230 (N_230,In_368,In_449);
and U231 (N_231,In_301,N_186);
nor U232 (N_232,N_179,In_36);
nand U233 (N_233,N_134,N_145);
nor U234 (N_234,In_307,In_57);
nand U235 (N_235,In_358,N_103);
or U236 (N_236,N_30,In_128);
and U237 (N_237,In_422,In_424);
or U238 (N_238,In_332,N_199);
nand U239 (N_239,N_54,In_88);
and U240 (N_240,N_122,N_66);
nor U241 (N_241,N_45,N_80);
nor U242 (N_242,In_394,N_107);
and U243 (N_243,In_387,In_370);
or U244 (N_244,N_157,In_375);
nor U245 (N_245,In_192,N_187);
or U246 (N_246,N_31,N_153);
nand U247 (N_247,N_11,N_93);
nand U248 (N_248,In_64,In_58);
xor U249 (N_249,N_2,N_168);
and U250 (N_250,N_92,N_53);
and U251 (N_251,N_70,In_214);
nor U252 (N_252,In_383,N_188);
nand U253 (N_253,In_70,N_74);
nand U254 (N_254,N_81,N_171);
nand U255 (N_255,In_345,N_109);
nand U256 (N_256,In_404,N_149);
nor U257 (N_257,In_197,N_102);
xor U258 (N_258,In_169,N_64);
nor U259 (N_259,N_120,N_68);
or U260 (N_260,N_195,N_147);
and U261 (N_261,N_86,In_477);
and U262 (N_262,In_476,N_142);
nor U263 (N_263,N_165,N_47);
nor U264 (N_264,N_197,In_156);
xor U265 (N_265,In_66,N_169);
nand U266 (N_266,N_26,N_158);
nand U267 (N_267,N_184,In_283);
and U268 (N_268,In_19,N_79);
nand U269 (N_269,N_124,In_443);
and U270 (N_270,In_400,In_83);
or U271 (N_271,In_324,In_366);
nand U272 (N_272,N_35,N_3);
nor U273 (N_273,N_191,In_269);
nor U274 (N_274,In_439,In_369);
nand U275 (N_275,N_52,N_155);
nor U276 (N_276,N_4,N_32);
and U277 (N_277,N_6,N_99);
and U278 (N_278,In_407,N_170);
nand U279 (N_279,N_159,N_174);
nor U280 (N_280,N_192,In_239);
and U281 (N_281,N_19,N_160);
nor U282 (N_282,N_182,N_8);
nor U283 (N_283,N_71,In_159);
and U284 (N_284,N_34,N_178);
nor U285 (N_285,N_22,N_73);
and U286 (N_286,In_91,N_156);
nor U287 (N_287,N_114,N_161);
nor U288 (N_288,N_91,N_61);
nor U289 (N_289,N_136,N_57);
nor U290 (N_290,N_190,In_252);
nand U291 (N_291,N_97,N_189);
nor U292 (N_292,N_137,N_98);
nor U293 (N_293,N_175,N_138);
and U294 (N_294,N_40,N_84);
nand U295 (N_295,N_9,N_28);
and U296 (N_296,N_48,N_55);
nand U297 (N_297,N_106,In_26);
and U298 (N_298,N_75,N_0);
and U299 (N_299,N_125,N_16);
xnor U300 (N_300,In_199,In_286);
nor U301 (N_301,N_14,N_108);
or U302 (N_302,In_163,In_264);
nand U303 (N_303,N_119,In_238);
or U304 (N_304,N_94,N_78);
and U305 (N_305,N_185,In_75);
or U306 (N_306,N_24,In_144);
or U307 (N_307,N_121,N_101);
nand U308 (N_308,In_303,N_146);
and U309 (N_309,N_194,N_7);
xnor U310 (N_310,N_65,N_62);
and U311 (N_311,N_72,N_135);
and U312 (N_312,In_276,N_118);
nor U313 (N_313,In_134,In_410);
nand U314 (N_314,N_15,N_87);
or U315 (N_315,N_164,In_108);
nor U316 (N_316,N_183,N_198);
and U317 (N_317,N_33,N_139);
nand U318 (N_318,N_127,In_100);
nand U319 (N_319,N_150,N_117);
or U320 (N_320,N_96,N_95);
nand U321 (N_321,In_270,N_50);
nor U322 (N_322,In_228,In_389);
nand U323 (N_323,In_317,N_17);
or U324 (N_324,In_126,N_140);
nor U325 (N_325,N_20,In_329);
and U326 (N_326,N_36,N_196);
and U327 (N_327,N_21,N_77);
and U328 (N_328,N_67,N_39);
and U329 (N_329,N_154,N_112);
nor U330 (N_330,N_41,In_334);
nor U331 (N_331,N_29,In_225);
nor U332 (N_332,N_23,N_88);
nor U333 (N_333,N_12,N_162);
or U334 (N_334,N_130,In_117);
nand U335 (N_335,N_10,N_180);
nor U336 (N_336,N_131,N_111);
and U337 (N_337,In_168,N_143);
nand U338 (N_338,In_105,In_278);
nand U339 (N_339,N_129,In_50);
and U340 (N_340,N_104,N_42);
nor U341 (N_341,In_469,In_10);
nor U342 (N_342,N_56,In_29);
and U343 (N_343,In_489,In_42);
nor U344 (N_344,In_456,N_166);
nor U345 (N_345,N_100,N_133);
and U346 (N_346,N_193,N_76);
and U347 (N_347,N_172,N_1);
nand U348 (N_348,N_132,In_112);
nand U349 (N_349,N_18,N_44);
nand U350 (N_350,N_41,N_172);
nor U351 (N_351,N_120,In_489);
or U352 (N_352,N_22,N_169);
or U353 (N_353,N_30,N_179);
and U354 (N_354,N_181,In_168);
nand U355 (N_355,In_36,In_383);
xor U356 (N_356,N_96,N_113);
xnor U357 (N_357,In_163,N_174);
nor U358 (N_358,N_29,In_232);
nand U359 (N_359,N_32,N_199);
nand U360 (N_360,N_5,N_150);
nor U361 (N_361,N_14,N_130);
nor U362 (N_362,N_66,In_199);
and U363 (N_363,N_5,In_108);
or U364 (N_364,N_135,N_114);
and U365 (N_365,In_404,In_400);
or U366 (N_366,In_407,N_124);
and U367 (N_367,N_149,N_30);
nand U368 (N_368,In_303,N_26);
and U369 (N_369,N_24,N_64);
and U370 (N_370,N_27,N_128);
and U371 (N_371,N_147,N_160);
nor U372 (N_372,N_71,N_92);
or U373 (N_373,N_132,In_283);
nor U374 (N_374,N_72,N_35);
and U375 (N_375,N_165,N_137);
and U376 (N_376,N_182,N_183);
nor U377 (N_377,N_126,N_136);
nand U378 (N_378,In_29,In_278);
and U379 (N_379,N_186,In_264);
or U380 (N_380,N_187,N_194);
xnor U381 (N_381,N_78,N_132);
nor U382 (N_382,In_410,N_98);
nor U383 (N_383,N_54,N_112);
and U384 (N_384,N_155,N_170);
nand U385 (N_385,N_180,In_237);
nor U386 (N_386,In_332,N_59);
nor U387 (N_387,In_276,N_123);
nor U388 (N_388,N_148,N_151);
nor U389 (N_389,N_41,N_63);
and U390 (N_390,In_383,N_119);
xor U391 (N_391,In_375,N_58);
nand U392 (N_392,In_83,In_264);
nand U393 (N_393,In_443,N_10);
and U394 (N_394,In_64,N_25);
or U395 (N_395,N_93,N_43);
nand U396 (N_396,In_422,N_147);
or U397 (N_397,N_173,In_242);
nand U398 (N_398,N_48,N_119);
nor U399 (N_399,In_404,In_26);
nor U400 (N_400,N_207,N_273);
or U401 (N_401,N_219,N_250);
nand U402 (N_402,N_259,N_300);
nor U403 (N_403,N_397,N_233);
nor U404 (N_404,N_387,N_241);
nand U405 (N_405,N_323,N_344);
and U406 (N_406,N_216,N_339);
and U407 (N_407,N_265,N_292);
nand U408 (N_408,N_340,N_261);
and U409 (N_409,N_303,N_368);
and U410 (N_410,N_230,N_364);
nand U411 (N_411,N_346,N_285);
xnor U412 (N_412,N_232,N_394);
nand U413 (N_413,N_386,N_319);
nand U414 (N_414,N_399,N_272);
nor U415 (N_415,N_375,N_389);
or U416 (N_416,N_200,N_353);
or U417 (N_417,N_263,N_248);
or U418 (N_418,N_298,N_302);
nand U419 (N_419,N_356,N_251);
or U420 (N_420,N_286,N_209);
xnor U421 (N_421,N_225,N_226);
nor U422 (N_422,N_279,N_260);
xnor U423 (N_423,N_244,N_224);
nand U424 (N_424,N_218,N_258);
nand U425 (N_425,N_213,N_235);
and U426 (N_426,N_229,N_270);
or U427 (N_427,N_307,N_212);
nand U428 (N_428,N_347,N_374);
nand U429 (N_429,N_255,N_227);
nor U430 (N_430,N_236,N_327);
xor U431 (N_431,N_379,N_243);
nand U432 (N_432,N_335,N_317);
and U433 (N_433,N_211,N_361);
and U434 (N_434,N_349,N_357);
and U435 (N_435,N_281,N_332);
nor U436 (N_436,N_383,N_322);
and U437 (N_437,N_294,N_311);
or U438 (N_438,N_382,N_264);
nor U439 (N_439,N_378,N_358);
nor U440 (N_440,N_262,N_352);
or U441 (N_441,N_398,N_329);
nand U442 (N_442,N_284,N_308);
or U443 (N_443,N_377,N_336);
or U444 (N_444,N_245,N_202);
and U445 (N_445,N_291,N_337);
nand U446 (N_446,N_393,N_201);
and U447 (N_447,N_277,N_326);
nor U448 (N_448,N_275,N_328);
nor U449 (N_449,N_363,N_391);
or U450 (N_450,N_214,N_256);
nor U451 (N_451,N_350,N_316);
and U452 (N_452,N_208,N_289);
nand U453 (N_453,N_370,N_305);
xor U454 (N_454,N_396,N_280);
nor U455 (N_455,N_367,N_333);
nor U456 (N_456,N_372,N_206);
and U457 (N_457,N_274,N_269);
nor U458 (N_458,N_282,N_309);
and U459 (N_459,N_334,N_238);
and U460 (N_460,N_257,N_310);
and U461 (N_461,N_321,N_355);
or U462 (N_462,N_395,N_295);
nor U463 (N_463,N_249,N_228);
and U464 (N_464,N_267,N_371);
or U465 (N_465,N_252,N_297);
nand U466 (N_466,N_296,N_242);
nand U467 (N_467,N_385,N_221);
nand U468 (N_468,N_345,N_354);
nand U469 (N_469,N_287,N_278);
nand U470 (N_470,N_390,N_343);
or U471 (N_471,N_290,N_373);
or U472 (N_472,N_223,N_366);
nand U473 (N_473,N_359,N_348);
nor U474 (N_474,N_362,N_380);
or U475 (N_475,N_301,N_239);
and U476 (N_476,N_217,N_320);
xor U477 (N_477,N_253,N_324);
and U478 (N_478,N_222,N_276);
and U479 (N_479,N_234,N_231);
nand U480 (N_480,N_288,N_351);
nor U481 (N_481,N_203,N_299);
and U482 (N_482,N_215,N_268);
or U483 (N_483,N_312,N_314);
or U484 (N_484,N_388,N_271);
or U485 (N_485,N_204,N_246);
or U486 (N_486,N_325,N_304);
nor U487 (N_487,N_293,N_369);
and U488 (N_488,N_331,N_306);
or U489 (N_489,N_205,N_237);
nor U490 (N_490,N_266,N_330);
or U491 (N_491,N_254,N_381);
and U492 (N_492,N_247,N_283);
or U493 (N_493,N_392,N_376);
nor U494 (N_494,N_338,N_365);
or U495 (N_495,N_341,N_360);
or U496 (N_496,N_315,N_210);
or U497 (N_497,N_384,N_240);
and U498 (N_498,N_313,N_342);
and U499 (N_499,N_220,N_318);
nor U500 (N_500,N_366,N_312);
and U501 (N_501,N_309,N_228);
nand U502 (N_502,N_330,N_314);
or U503 (N_503,N_234,N_263);
or U504 (N_504,N_332,N_272);
and U505 (N_505,N_318,N_271);
and U506 (N_506,N_211,N_213);
or U507 (N_507,N_253,N_330);
nand U508 (N_508,N_338,N_375);
or U509 (N_509,N_375,N_245);
and U510 (N_510,N_293,N_206);
nor U511 (N_511,N_241,N_239);
and U512 (N_512,N_296,N_352);
or U513 (N_513,N_313,N_248);
nand U514 (N_514,N_290,N_271);
or U515 (N_515,N_270,N_386);
nor U516 (N_516,N_277,N_360);
and U517 (N_517,N_358,N_375);
and U518 (N_518,N_295,N_352);
xnor U519 (N_519,N_211,N_229);
nor U520 (N_520,N_207,N_254);
and U521 (N_521,N_334,N_392);
and U522 (N_522,N_283,N_225);
nor U523 (N_523,N_279,N_295);
and U524 (N_524,N_202,N_341);
or U525 (N_525,N_332,N_361);
nor U526 (N_526,N_371,N_205);
nor U527 (N_527,N_206,N_324);
nand U528 (N_528,N_256,N_272);
or U529 (N_529,N_379,N_222);
nor U530 (N_530,N_347,N_248);
nor U531 (N_531,N_241,N_219);
and U532 (N_532,N_296,N_297);
or U533 (N_533,N_203,N_363);
xnor U534 (N_534,N_209,N_307);
nand U535 (N_535,N_363,N_336);
or U536 (N_536,N_243,N_249);
and U537 (N_537,N_335,N_337);
or U538 (N_538,N_240,N_386);
or U539 (N_539,N_226,N_204);
or U540 (N_540,N_314,N_245);
nand U541 (N_541,N_349,N_227);
nor U542 (N_542,N_252,N_276);
and U543 (N_543,N_258,N_270);
nand U544 (N_544,N_232,N_327);
nor U545 (N_545,N_360,N_225);
nand U546 (N_546,N_372,N_375);
and U547 (N_547,N_277,N_241);
or U548 (N_548,N_300,N_313);
nand U549 (N_549,N_269,N_372);
nor U550 (N_550,N_346,N_239);
nand U551 (N_551,N_322,N_329);
and U552 (N_552,N_366,N_235);
nand U553 (N_553,N_394,N_238);
or U554 (N_554,N_259,N_357);
or U555 (N_555,N_380,N_356);
and U556 (N_556,N_370,N_315);
or U557 (N_557,N_246,N_264);
and U558 (N_558,N_204,N_326);
nand U559 (N_559,N_330,N_208);
or U560 (N_560,N_375,N_315);
nor U561 (N_561,N_237,N_340);
nor U562 (N_562,N_215,N_388);
nand U563 (N_563,N_292,N_232);
or U564 (N_564,N_268,N_244);
or U565 (N_565,N_292,N_244);
or U566 (N_566,N_371,N_375);
and U567 (N_567,N_233,N_245);
or U568 (N_568,N_310,N_326);
nor U569 (N_569,N_384,N_216);
and U570 (N_570,N_384,N_283);
nor U571 (N_571,N_295,N_249);
or U572 (N_572,N_225,N_391);
and U573 (N_573,N_202,N_241);
and U574 (N_574,N_252,N_298);
nor U575 (N_575,N_292,N_351);
nor U576 (N_576,N_381,N_221);
nand U577 (N_577,N_264,N_279);
or U578 (N_578,N_268,N_389);
and U579 (N_579,N_228,N_269);
nor U580 (N_580,N_279,N_290);
or U581 (N_581,N_283,N_226);
or U582 (N_582,N_270,N_344);
nand U583 (N_583,N_302,N_238);
or U584 (N_584,N_335,N_353);
or U585 (N_585,N_375,N_234);
and U586 (N_586,N_301,N_235);
nand U587 (N_587,N_382,N_216);
and U588 (N_588,N_251,N_217);
or U589 (N_589,N_283,N_219);
or U590 (N_590,N_398,N_200);
and U591 (N_591,N_249,N_230);
nand U592 (N_592,N_249,N_263);
or U593 (N_593,N_278,N_347);
and U594 (N_594,N_363,N_376);
and U595 (N_595,N_352,N_395);
nor U596 (N_596,N_381,N_219);
and U597 (N_597,N_204,N_278);
or U598 (N_598,N_223,N_343);
nand U599 (N_599,N_311,N_319);
nor U600 (N_600,N_461,N_468);
nand U601 (N_601,N_491,N_504);
and U602 (N_602,N_446,N_456);
nand U603 (N_603,N_583,N_598);
nand U604 (N_604,N_453,N_594);
nor U605 (N_605,N_506,N_514);
and U606 (N_606,N_557,N_499);
or U607 (N_607,N_459,N_497);
and U608 (N_608,N_515,N_512);
nand U609 (N_609,N_546,N_571);
nand U610 (N_610,N_490,N_457);
nor U611 (N_611,N_418,N_413);
or U612 (N_612,N_467,N_484);
nor U613 (N_613,N_523,N_486);
or U614 (N_614,N_581,N_465);
and U615 (N_615,N_590,N_508);
or U616 (N_616,N_405,N_529);
or U617 (N_617,N_547,N_574);
nand U618 (N_618,N_430,N_445);
nor U619 (N_619,N_509,N_427);
xnor U620 (N_620,N_584,N_537);
and U621 (N_621,N_488,N_409);
or U622 (N_622,N_558,N_522);
xor U623 (N_623,N_585,N_441);
nor U624 (N_624,N_443,N_551);
and U625 (N_625,N_505,N_424);
nand U626 (N_626,N_544,N_552);
and U627 (N_627,N_483,N_404);
nor U628 (N_628,N_464,N_421);
or U629 (N_629,N_535,N_554);
nand U630 (N_630,N_451,N_543);
nand U631 (N_631,N_586,N_530);
or U632 (N_632,N_423,N_496);
nor U633 (N_633,N_489,N_526);
nand U634 (N_634,N_481,N_541);
and U635 (N_635,N_596,N_498);
and U636 (N_636,N_563,N_435);
or U637 (N_637,N_479,N_533);
or U638 (N_638,N_415,N_428);
nor U639 (N_639,N_532,N_476);
nor U640 (N_640,N_438,N_475);
or U641 (N_641,N_442,N_434);
or U642 (N_642,N_556,N_559);
or U643 (N_643,N_507,N_545);
nor U644 (N_644,N_444,N_576);
nor U645 (N_645,N_494,N_539);
xor U646 (N_646,N_538,N_450);
xnor U647 (N_647,N_495,N_500);
nand U648 (N_648,N_448,N_471);
and U649 (N_649,N_401,N_536);
nand U650 (N_650,N_580,N_587);
nand U651 (N_651,N_542,N_567);
nor U652 (N_652,N_597,N_540);
or U653 (N_653,N_501,N_439);
nand U654 (N_654,N_452,N_503);
and U655 (N_655,N_518,N_449);
or U656 (N_656,N_455,N_429);
or U657 (N_657,N_454,N_589);
nor U658 (N_658,N_458,N_520);
and U659 (N_659,N_473,N_466);
or U660 (N_660,N_564,N_569);
nand U661 (N_661,N_517,N_548);
or U662 (N_662,N_521,N_422);
xnor U663 (N_663,N_433,N_407);
nor U664 (N_664,N_555,N_534);
and U665 (N_665,N_437,N_560);
nor U666 (N_666,N_578,N_412);
and U667 (N_667,N_414,N_474);
nor U668 (N_668,N_469,N_463);
or U669 (N_669,N_527,N_595);
or U670 (N_670,N_516,N_524);
and U671 (N_671,N_493,N_565);
nor U672 (N_672,N_416,N_408);
and U673 (N_673,N_440,N_410);
nand U674 (N_674,N_502,N_492);
or U675 (N_675,N_513,N_572);
xnor U676 (N_676,N_553,N_591);
and U677 (N_677,N_519,N_432);
nand U678 (N_678,N_550,N_588);
nand U679 (N_679,N_447,N_561);
nand U680 (N_680,N_593,N_549);
and U681 (N_681,N_480,N_470);
and U682 (N_682,N_406,N_570);
or U683 (N_683,N_419,N_525);
and U684 (N_684,N_426,N_592);
or U685 (N_685,N_460,N_472);
and U686 (N_686,N_575,N_577);
nand U687 (N_687,N_511,N_573);
and U688 (N_688,N_411,N_510);
or U689 (N_689,N_478,N_417);
xor U690 (N_690,N_400,N_425);
xnor U691 (N_691,N_568,N_402);
nand U692 (N_692,N_531,N_436);
or U693 (N_693,N_579,N_482);
and U694 (N_694,N_487,N_477);
nor U695 (N_695,N_403,N_566);
nand U696 (N_696,N_462,N_528);
or U697 (N_697,N_582,N_562);
or U698 (N_698,N_599,N_431);
or U699 (N_699,N_420,N_485);
nor U700 (N_700,N_527,N_423);
and U701 (N_701,N_534,N_466);
nand U702 (N_702,N_469,N_483);
nand U703 (N_703,N_453,N_591);
nor U704 (N_704,N_551,N_470);
nand U705 (N_705,N_572,N_509);
or U706 (N_706,N_504,N_409);
nor U707 (N_707,N_559,N_565);
nand U708 (N_708,N_465,N_449);
and U709 (N_709,N_593,N_489);
nor U710 (N_710,N_415,N_591);
or U711 (N_711,N_462,N_483);
and U712 (N_712,N_506,N_408);
or U713 (N_713,N_475,N_538);
and U714 (N_714,N_595,N_576);
nand U715 (N_715,N_541,N_434);
or U716 (N_716,N_414,N_584);
or U717 (N_717,N_595,N_512);
nor U718 (N_718,N_475,N_546);
nor U719 (N_719,N_451,N_412);
nand U720 (N_720,N_564,N_426);
or U721 (N_721,N_465,N_476);
nand U722 (N_722,N_470,N_499);
nand U723 (N_723,N_527,N_460);
nor U724 (N_724,N_530,N_410);
nand U725 (N_725,N_412,N_508);
or U726 (N_726,N_485,N_570);
nor U727 (N_727,N_558,N_495);
nand U728 (N_728,N_539,N_552);
and U729 (N_729,N_457,N_496);
nor U730 (N_730,N_520,N_528);
and U731 (N_731,N_575,N_544);
or U732 (N_732,N_508,N_446);
or U733 (N_733,N_541,N_546);
nor U734 (N_734,N_542,N_460);
or U735 (N_735,N_478,N_574);
or U736 (N_736,N_481,N_550);
nand U737 (N_737,N_402,N_487);
and U738 (N_738,N_525,N_530);
nand U739 (N_739,N_439,N_498);
nor U740 (N_740,N_516,N_483);
and U741 (N_741,N_510,N_401);
or U742 (N_742,N_478,N_452);
nand U743 (N_743,N_436,N_473);
or U744 (N_744,N_503,N_414);
nor U745 (N_745,N_495,N_468);
nor U746 (N_746,N_580,N_496);
and U747 (N_747,N_427,N_445);
or U748 (N_748,N_415,N_504);
or U749 (N_749,N_468,N_401);
and U750 (N_750,N_534,N_473);
nor U751 (N_751,N_496,N_484);
and U752 (N_752,N_411,N_431);
nand U753 (N_753,N_410,N_434);
or U754 (N_754,N_523,N_531);
nand U755 (N_755,N_561,N_495);
and U756 (N_756,N_426,N_494);
nand U757 (N_757,N_429,N_582);
or U758 (N_758,N_585,N_491);
or U759 (N_759,N_488,N_588);
nor U760 (N_760,N_543,N_565);
or U761 (N_761,N_588,N_551);
or U762 (N_762,N_407,N_501);
and U763 (N_763,N_515,N_449);
or U764 (N_764,N_597,N_458);
nand U765 (N_765,N_443,N_476);
or U766 (N_766,N_563,N_532);
and U767 (N_767,N_471,N_495);
and U768 (N_768,N_454,N_582);
nor U769 (N_769,N_433,N_591);
nor U770 (N_770,N_525,N_499);
nor U771 (N_771,N_512,N_470);
or U772 (N_772,N_588,N_443);
nor U773 (N_773,N_543,N_497);
and U774 (N_774,N_440,N_547);
nor U775 (N_775,N_568,N_410);
nor U776 (N_776,N_531,N_545);
and U777 (N_777,N_492,N_416);
or U778 (N_778,N_454,N_413);
or U779 (N_779,N_526,N_442);
nor U780 (N_780,N_590,N_548);
nand U781 (N_781,N_555,N_466);
xnor U782 (N_782,N_509,N_580);
nor U783 (N_783,N_413,N_538);
nand U784 (N_784,N_547,N_576);
or U785 (N_785,N_413,N_455);
and U786 (N_786,N_484,N_516);
xor U787 (N_787,N_405,N_429);
nand U788 (N_788,N_404,N_592);
nor U789 (N_789,N_467,N_595);
nor U790 (N_790,N_428,N_456);
and U791 (N_791,N_420,N_560);
nor U792 (N_792,N_494,N_469);
or U793 (N_793,N_404,N_578);
or U794 (N_794,N_594,N_470);
nor U795 (N_795,N_441,N_577);
and U796 (N_796,N_468,N_402);
nand U797 (N_797,N_540,N_551);
nor U798 (N_798,N_521,N_513);
nand U799 (N_799,N_447,N_469);
and U800 (N_800,N_660,N_796);
and U801 (N_801,N_630,N_685);
nand U802 (N_802,N_674,N_643);
and U803 (N_803,N_797,N_669);
and U804 (N_804,N_746,N_725);
nor U805 (N_805,N_614,N_753);
xor U806 (N_806,N_784,N_772);
or U807 (N_807,N_798,N_728);
nand U808 (N_808,N_686,N_778);
nand U809 (N_809,N_737,N_745);
nand U810 (N_810,N_601,N_622);
nand U811 (N_811,N_717,N_793);
or U812 (N_812,N_786,N_767);
and U813 (N_813,N_758,N_649);
xnor U814 (N_814,N_641,N_678);
and U815 (N_815,N_713,N_705);
nand U816 (N_816,N_799,N_756);
or U817 (N_817,N_739,N_671);
nand U818 (N_818,N_629,N_761);
nand U819 (N_819,N_723,N_646);
nand U820 (N_820,N_600,N_736);
or U821 (N_821,N_738,N_779);
nor U822 (N_822,N_608,N_611);
and U823 (N_823,N_644,N_710);
nor U824 (N_824,N_700,N_744);
nor U825 (N_825,N_691,N_607);
or U826 (N_826,N_795,N_742);
and U827 (N_827,N_708,N_662);
nor U828 (N_828,N_677,N_659);
and U829 (N_829,N_731,N_690);
and U830 (N_830,N_768,N_626);
or U831 (N_831,N_670,N_760);
or U832 (N_832,N_610,N_722);
nand U833 (N_833,N_785,N_763);
nand U834 (N_834,N_667,N_730);
nand U835 (N_835,N_766,N_762);
or U836 (N_836,N_656,N_675);
or U837 (N_837,N_698,N_651);
nor U838 (N_838,N_620,N_765);
nor U839 (N_839,N_773,N_748);
and U840 (N_840,N_769,N_618);
and U841 (N_841,N_615,N_645);
nand U842 (N_842,N_719,N_639);
and U843 (N_843,N_788,N_774);
and U844 (N_844,N_775,N_628);
and U845 (N_845,N_636,N_634);
nand U846 (N_846,N_612,N_602);
nand U847 (N_847,N_695,N_653);
xor U848 (N_848,N_782,N_791);
and U849 (N_849,N_684,N_790);
or U850 (N_850,N_741,N_687);
and U851 (N_851,N_661,N_633);
and U852 (N_852,N_640,N_740);
or U853 (N_853,N_727,N_642);
and U854 (N_854,N_676,N_777);
nor U855 (N_855,N_781,N_755);
or U856 (N_856,N_603,N_616);
or U857 (N_857,N_759,N_693);
nor U858 (N_858,N_624,N_711);
nor U859 (N_859,N_694,N_697);
nor U860 (N_860,N_702,N_679);
nor U861 (N_861,N_625,N_726);
or U862 (N_862,N_672,N_680);
or U863 (N_863,N_701,N_637);
and U864 (N_864,N_735,N_689);
and U865 (N_865,N_709,N_605);
nand U866 (N_866,N_668,N_655);
or U867 (N_867,N_609,N_658);
and U868 (N_868,N_617,N_771);
nand U869 (N_869,N_794,N_619);
nor U870 (N_870,N_692,N_673);
nand U871 (N_871,N_757,N_652);
and U872 (N_872,N_627,N_783);
and U873 (N_873,N_776,N_654);
nand U874 (N_874,N_699,N_704);
nand U875 (N_875,N_706,N_703);
nor U876 (N_876,N_712,N_666);
and U877 (N_877,N_635,N_683);
nand U878 (N_878,N_650,N_707);
and U879 (N_879,N_754,N_664);
or U880 (N_880,N_688,N_604);
nor U881 (N_881,N_792,N_613);
nor U882 (N_882,N_657,N_638);
nor U883 (N_883,N_789,N_787);
nand U884 (N_884,N_732,N_696);
nor U885 (N_885,N_682,N_665);
and U886 (N_886,N_749,N_663);
or U887 (N_887,N_632,N_752);
nor U888 (N_888,N_747,N_720);
nand U889 (N_889,N_764,N_621);
and U890 (N_890,N_724,N_716);
nor U891 (N_891,N_623,N_729);
or U892 (N_892,N_733,N_715);
nand U893 (N_893,N_751,N_631);
nor U894 (N_894,N_718,N_770);
nor U895 (N_895,N_780,N_721);
and U896 (N_896,N_714,N_606);
nand U897 (N_897,N_648,N_681);
and U898 (N_898,N_743,N_734);
nor U899 (N_899,N_750,N_647);
nand U900 (N_900,N_745,N_738);
nand U901 (N_901,N_606,N_671);
xnor U902 (N_902,N_728,N_654);
nor U903 (N_903,N_750,N_781);
and U904 (N_904,N_642,N_684);
and U905 (N_905,N_716,N_645);
nand U906 (N_906,N_758,N_789);
xor U907 (N_907,N_648,N_625);
and U908 (N_908,N_695,N_706);
nand U909 (N_909,N_635,N_609);
nand U910 (N_910,N_750,N_658);
and U911 (N_911,N_696,N_662);
nand U912 (N_912,N_745,N_720);
and U913 (N_913,N_764,N_741);
and U914 (N_914,N_701,N_723);
nand U915 (N_915,N_708,N_692);
or U916 (N_916,N_639,N_794);
and U917 (N_917,N_701,N_725);
and U918 (N_918,N_691,N_606);
and U919 (N_919,N_683,N_760);
nand U920 (N_920,N_780,N_689);
and U921 (N_921,N_659,N_703);
xnor U922 (N_922,N_684,N_625);
nor U923 (N_923,N_617,N_778);
and U924 (N_924,N_625,N_615);
nor U925 (N_925,N_690,N_663);
or U926 (N_926,N_698,N_600);
nand U927 (N_927,N_771,N_629);
or U928 (N_928,N_722,N_746);
xnor U929 (N_929,N_662,N_778);
nor U930 (N_930,N_798,N_663);
and U931 (N_931,N_718,N_739);
or U932 (N_932,N_659,N_784);
nor U933 (N_933,N_661,N_686);
nor U934 (N_934,N_619,N_779);
or U935 (N_935,N_749,N_606);
and U936 (N_936,N_626,N_690);
nand U937 (N_937,N_693,N_726);
or U938 (N_938,N_779,N_773);
or U939 (N_939,N_622,N_687);
or U940 (N_940,N_645,N_776);
and U941 (N_941,N_640,N_754);
and U942 (N_942,N_692,N_731);
nand U943 (N_943,N_712,N_622);
nor U944 (N_944,N_738,N_771);
or U945 (N_945,N_698,N_763);
or U946 (N_946,N_728,N_702);
or U947 (N_947,N_739,N_767);
or U948 (N_948,N_778,N_612);
nor U949 (N_949,N_743,N_776);
nor U950 (N_950,N_623,N_616);
or U951 (N_951,N_695,N_783);
or U952 (N_952,N_718,N_629);
nand U953 (N_953,N_728,N_675);
nor U954 (N_954,N_761,N_752);
nor U955 (N_955,N_714,N_650);
nor U956 (N_956,N_692,N_679);
nor U957 (N_957,N_787,N_603);
and U958 (N_958,N_671,N_605);
or U959 (N_959,N_623,N_706);
nor U960 (N_960,N_731,N_606);
nand U961 (N_961,N_629,N_627);
nor U962 (N_962,N_796,N_601);
nor U963 (N_963,N_725,N_704);
nor U964 (N_964,N_770,N_608);
or U965 (N_965,N_731,N_623);
and U966 (N_966,N_703,N_760);
and U967 (N_967,N_661,N_733);
and U968 (N_968,N_640,N_786);
and U969 (N_969,N_723,N_633);
nor U970 (N_970,N_668,N_787);
nor U971 (N_971,N_637,N_707);
and U972 (N_972,N_741,N_607);
or U973 (N_973,N_706,N_629);
or U974 (N_974,N_786,N_709);
xnor U975 (N_975,N_735,N_639);
nor U976 (N_976,N_660,N_791);
or U977 (N_977,N_620,N_763);
nand U978 (N_978,N_754,N_728);
or U979 (N_979,N_773,N_754);
and U980 (N_980,N_604,N_637);
nand U981 (N_981,N_731,N_750);
nor U982 (N_982,N_639,N_795);
or U983 (N_983,N_748,N_797);
nand U984 (N_984,N_792,N_606);
nor U985 (N_985,N_722,N_644);
nand U986 (N_986,N_787,N_642);
nand U987 (N_987,N_741,N_720);
nor U988 (N_988,N_792,N_616);
nor U989 (N_989,N_630,N_678);
or U990 (N_990,N_759,N_743);
nand U991 (N_991,N_749,N_629);
or U992 (N_992,N_609,N_679);
nand U993 (N_993,N_675,N_607);
nor U994 (N_994,N_665,N_684);
nor U995 (N_995,N_669,N_671);
nand U996 (N_996,N_731,N_621);
nand U997 (N_997,N_770,N_783);
or U998 (N_998,N_685,N_728);
or U999 (N_999,N_690,N_782);
xnor U1000 (N_1000,N_939,N_943);
or U1001 (N_1001,N_880,N_819);
and U1002 (N_1002,N_987,N_917);
or U1003 (N_1003,N_849,N_936);
nor U1004 (N_1004,N_850,N_892);
nor U1005 (N_1005,N_967,N_928);
and U1006 (N_1006,N_813,N_888);
nor U1007 (N_1007,N_872,N_840);
or U1008 (N_1008,N_983,N_916);
nand U1009 (N_1009,N_816,N_870);
nand U1010 (N_1010,N_864,N_860);
or U1011 (N_1011,N_809,N_823);
and U1012 (N_1012,N_838,N_893);
nor U1013 (N_1013,N_990,N_802);
nor U1014 (N_1014,N_821,N_854);
nor U1015 (N_1015,N_918,N_830);
nor U1016 (N_1016,N_997,N_826);
and U1017 (N_1017,N_906,N_904);
nor U1018 (N_1018,N_804,N_898);
nor U1019 (N_1019,N_811,N_933);
and U1020 (N_1020,N_922,N_837);
nor U1021 (N_1021,N_889,N_969);
or U1022 (N_1022,N_896,N_842);
nor U1023 (N_1023,N_964,N_881);
or U1024 (N_1024,N_828,N_911);
or U1025 (N_1025,N_859,N_873);
or U1026 (N_1026,N_940,N_993);
or U1027 (N_1027,N_952,N_865);
or U1028 (N_1028,N_812,N_862);
or U1029 (N_1029,N_942,N_808);
or U1030 (N_1030,N_947,N_908);
and U1031 (N_1031,N_937,N_920);
nand U1032 (N_1032,N_944,N_978);
and U1033 (N_1033,N_949,N_836);
and U1034 (N_1034,N_847,N_962);
or U1035 (N_1035,N_909,N_930);
or U1036 (N_1036,N_806,N_878);
or U1037 (N_1037,N_955,N_883);
and U1038 (N_1038,N_975,N_886);
nand U1039 (N_1039,N_844,N_998);
nor U1040 (N_1040,N_891,N_919);
nand U1041 (N_1041,N_950,N_938);
nand U1042 (N_1042,N_985,N_807);
nor U1043 (N_1043,N_925,N_877);
nor U1044 (N_1044,N_900,N_853);
or U1045 (N_1045,N_984,N_994);
nor U1046 (N_1046,N_824,N_981);
nor U1047 (N_1047,N_946,N_831);
nand U1048 (N_1048,N_801,N_833);
nand U1049 (N_1049,N_982,N_827);
nor U1050 (N_1050,N_958,N_810);
and U1051 (N_1051,N_834,N_858);
or U1052 (N_1052,N_926,N_868);
nor U1053 (N_1053,N_825,N_876);
nor U1054 (N_1054,N_961,N_992);
nand U1055 (N_1055,N_913,N_832);
and U1056 (N_1056,N_866,N_829);
nand U1057 (N_1057,N_959,N_966);
and U1058 (N_1058,N_910,N_848);
and U1059 (N_1059,N_945,N_934);
nand U1060 (N_1060,N_953,N_935);
or U1061 (N_1061,N_820,N_863);
nand U1062 (N_1062,N_931,N_960);
nand U1063 (N_1063,N_815,N_852);
and U1064 (N_1064,N_805,N_897);
and U1065 (N_1065,N_875,N_991);
nor U1066 (N_1066,N_869,N_914);
nor U1067 (N_1067,N_856,N_927);
and U1068 (N_1068,N_890,N_841);
nor U1069 (N_1069,N_843,N_970);
nand U1070 (N_1070,N_867,N_932);
and U1071 (N_1071,N_979,N_839);
nor U1072 (N_1072,N_973,N_887);
nand U1073 (N_1073,N_874,N_996);
nand U1074 (N_1074,N_905,N_907);
or U1075 (N_1075,N_956,N_915);
and U1076 (N_1076,N_976,N_954);
and U1077 (N_1077,N_965,N_971);
or U1078 (N_1078,N_871,N_885);
nor U1079 (N_1079,N_803,N_846);
or U1080 (N_1080,N_980,N_968);
and U1081 (N_1081,N_951,N_963);
xor U1082 (N_1082,N_855,N_924);
or U1083 (N_1083,N_921,N_857);
nor U1084 (N_1084,N_845,N_948);
nor U1085 (N_1085,N_986,N_822);
and U1086 (N_1086,N_818,N_974);
nor U1087 (N_1087,N_817,N_912);
nand U1088 (N_1088,N_895,N_879);
nand U1089 (N_1089,N_972,N_899);
or U1090 (N_1090,N_884,N_882);
nand U1091 (N_1091,N_929,N_989);
and U1092 (N_1092,N_977,N_894);
nand U1093 (N_1093,N_941,N_902);
or U1094 (N_1094,N_800,N_835);
or U1095 (N_1095,N_995,N_923);
nor U1096 (N_1096,N_957,N_988);
nor U1097 (N_1097,N_999,N_814);
and U1098 (N_1098,N_851,N_901);
nor U1099 (N_1099,N_903,N_861);
or U1100 (N_1100,N_844,N_863);
nand U1101 (N_1101,N_896,N_983);
nand U1102 (N_1102,N_996,N_962);
and U1103 (N_1103,N_904,N_896);
nand U1104 (N_1104,N_808,N_852);
nand U1105 (N_1105,N_958,N_945);
nand U1106 (N_1106,N_955,N_839);
nor U1107 (N_1107,N_906,N_865);
nor U1108 (N_1108,N_840,N_915);
or U1109 (N_1109,N_814,N_896);
xnor U1110 (N_1110,N_914,N_899);
or U1111 (N_1111,N_938,N_888);
nor U1112 (N_1112,N_961,N_850);
nor U1113 (N_1113,N_967,N_989);
and U1114 (N_1114,N_943,N_932);
and U1115 (N_1115,N_812,N_882);
nor U1116 (N_1116,N_867,N_970);
or U1117 (N_1117,N_939,N_824);
xnor U1118 (N_1118,N_967,N_877);
nand U1119 (N_1119,N_935,N_872);
or U1120 (N_1120,N_980,N_933);
nand U1121 (N_1121,N_834,N_880);
nand U1122 (N_1122,N_900,N_874);
nor U1123 (N_1123,N_870,N_843);
nor U1124 (N_1124,N_946,N_882);
and U1125 (N_1125,N_834,N_954);
nand U1126 (N_1126,N_874,N_965);
and U1127 (N_1127,N_946,N_988);
and U1128 (N_1128,N_959,N_876);
and U1129 (N_1129,N_887,N_932);
nor U1130 (N_1130,N_956,N_911);
or U1131 (N_1131,N_935,N_983);
nand U1132 (N_1132,N_944,N_981);
nor U1133 (N_1133,N_849,N_982);
nand U1134 (N_1134,N_869,N_938);
and U1135 (N_1135,N_888,N_892);
and U1136 (N_1136,N_987,N_928);
and U1137 (N_1137,N_964,N_928);
xor U1138 (N_1138,N_983,N_949);
nor U1139 (N_1139,N_948,N_848);
nor U1140 (N_1140,N_820,N_964);
nand U1141 (N_1141,N_847,N_911);
or U1142 (N_1142,N_964,N_925);
and U1143 (N_1143,N_990,N_807);
and U1144 (N_1144,N_819,N_823);
nand U1145 (N_1145,N_832,N_916);
nor U1146 (N_1146,N_935,N_869);
and U1147 (N_1147,N_827,N_804);
or U1148 (N_1148,N_856,N_979);
nand U1149 (N_1149,N_944,N_895);
nand U1150 (N_1150,N_905,N_991);
nor U1151 (N_1151,N_812,N_980);
and U1152 (N_1152,N_891,N_840);
nor U1153 (N_1153,N_985,N_817);
nor U1154 (N_1154,N_837,N_959);
nand U1155 (N_1155,N_851,N_931);
nand U1156 (N_1156,N_894,N_805);
nand U1157 (N_1157,N_844,N_971);
nand U1158 (N_1158,N_829,N_884);
or U1159 (N_1159,N_871,N_955);
nand U1160 (N_1160,N_944,N_974);
nor U1161 (N_1161,N_855,N_827);
and U1162 (N_1162,N_893,N_830);
or U1163 (N_1163,N_956,N_818);
nor U1164 (N_1164,N_845,N_879);
nand U1165 (N_1165,N_920,N_930);
xnor U1166 (N_1166,N_886,N_938);
nor U1167 (N_1167,N_875,N_862);
or U1168 (N_1168,N_828,N_999);
or U1169 (N_1169,N_959,N_905);
or U1170 (N_1170,N_821,N_815);
nor U1171 (N_1171,N_968,N_955);
nand U1172 (N_1172,N_986,N_945);
nand U1173 (N_1173,N_900,N_812);
or U1174 (N_1174,N_848,N_991);
or U1175 (N_1175,N_886,N_839);
or U1176 (N_1176,N_828,N_885);
or U1177 (N_1177,N_855,N_818);
or U1178 (N_1178,N_947,N_852);
nand U1179 (N_1179,N_938,N_868);
and U1180 (N_1180,N_828,N_997);
nor U1181 (N_1181,N_808,N_927);
nand U1182 (N_1182,N_821,N_939);
nand U1183 (N_1183,N_916,N_981);
and U1184 (N_1184,N_998,N_918);
nand U1185 (N_1185,N_833,N_921);
nand U1186 (N_1186,N_848,N_939);
nor U1187 (N_1187,N_859,N_894);
and U1188 (N_1188,N_894,N_934);
and U1189 (N_1189,N_898,N_841);
nor U1190 (N_1190,N_899,N_905);
or U1191 (N_1191,N_825,N_927);
nor U1192 (N_1192,N_869,N_936);
or U1193 (N_1193,N_999,N_869);
or U1194 (N_1194,N_818,N_854);
nor U1195 (N_1195,N_873,N_900);
or U1196 (N_1196,N_883,N_834);
nor U1197 (N_1197,N_927,N_828);
or U1198 (N_1198,N_885,N_930);
or U1199 (N_1199,N_880,N_953);
and U1200 (N_1200,N_1003,N_1140);
and U1201 (N_1201,N_1009,N_1085);
nor U1202 (N_1202,N_1192,N_1118);
and U1203 (N_1203,N_1083,N_1036);
or U1204 (N_1204,N_1099,N_1107);
and U1205 (N_1205,N_1135,N_1053);
or U1206 (N_1206,N_1178,N_1113);
xor U1207 (N_1207,N_1055,N_1082);
nor U1208 (N_1208,N_1195,N_1026);
nand U1209 (N_1209,N_1191,N_1148);
xnor U1210 (N_1210,N_1045,N_1087);
nor U1211 (N_1211,N_1096,N_1056);
and U1212 (N_1212,N_1095,N_1090);
or U1213 (N_1213,N_1180,N_1170);
nor U1214 (N_1214,N_1164,N_1077);
or U1215 (N_1215,N_1187,N_1112);
and U1216 (N_1216,N_1144,N_1182);
nor U1217 (N_1217,N_1080,N_1198);
nand U1218 (N_1218,N_1196,N_1151);
and U1219 (N_1219,N_1158,N_1162);
nand U1220 (N_1220,N_1066,N_1146);
nand U1221 (N_1221,N_1021,N_1044);
nor U1222 (N_1222,N_1027,N_1068);
and U1223 (N_1223,N_1069,N_1150);
and U1224 (N_1224,N_1011,N_1037);
xor U1225 (N_1225,N_1124,N_1015);
and U1226 (N_1226,N_1172,N_1032);
and U1227 (N_1227,N_1040,N_1183);
nor U1228 (N_1228,N_1057,N_1020);
and U1229 (N_1229,N_1154,N_1089);
xor U1230 (N_1230,N_1052,N_1078);
nor U1231 (N_1231,N_1049,N_1145);
nand U1232 (N_1232,N_1035,N_1104);
and U1233 (N_1233,N_1159,N_1122);
xor U1234 (N_1234,N_1119,N_1141);
nor U1235 (N_1235,N_1058,N_1163);
xnor U1236 (N_1236,N_1152,N_1093);
nor U1237 (N_1237,N_1102,N_1184);
nand U1238 (N_1238,N_1063,N_1060);
and U1239 (N_1239,N_1153,N_1006);
and U1240 (N_1240,N_1030,N_1149);
and U1241 (N_1241,N_1092,N_1130);
nor U1242 (N_1242,N_1174,N_1143);
and U1243 (N_1243,N_1034,N_1016);
nor U1244 (N_1244,N_1022,N_1156);
nor U1245 (N_1245,N_1038,N_1181);
or U1246 (N_1246,N_1199,N_1160);
nor U1247 (N_1247,N_1074,N_1046);
or U1248 (N_1248,N_1007,N_1147);
and U1249 (N_1249,N_1193,N_1041);
nor U1250 (N_1250,N_1125,N_1039);
or U1251 (N_1251,N_1098,N_1079);
and U1252 (N_1252,N_1194,N_1111);
or U1253 (N_1253,N_1029,N_1012);
nand U1254 (N_1254,N_1185,N_1086);
nand U1255 (N_1255,N_1000,N_1008);
and U1256 (N_1256,N_1103,N_1142);
nand U1257 (N_1257,N_1167,N_1054);
nor U1258 (N_1258,N_1128,N_1127);
nor U1259 (N_1259,N_1065,N_1101);
nand U1260 (N_1260,N_1166,N_1100);
and U1261 (N_1261,N_1070,N_1123);
xor U1262 (N_1262,N_1088,N_1018);
or U1263 (N_1263,N_1108,N_1121);
nor U1264 (N_1264,N_1097,N_1050);
nor U1265 (N_1265,N_1106,N_1179);
xor U1266 (N_1266,N_1043,N_1042);
xnor U1267 (N_1267,N_1134,N_1173);
or U1268 (N_1268,N_1129,N_1189);
and U1269 (N_1269,N_1132,N_1117);
and U1270 (N_1270,N_1025,N_1155);
nand U1271 (N_1271,N_1062,N_1126);
nand U1272 (N_1272,N_1168,N_1019);
nand U1273 (N_1273,N_1013,N_1033);
or U1274 (N_1274,N_1169,N_1071);
xnor U1275 (N_1275,N_1105,N_1115);
or U1276 (N_1276,N_1190,N_1005);
or U1277 (N_1277,N_1137,N_1076);
nand U1278 (N_1278,N_1175,N_1028);
and U1279 (N_1279,N_1059,N_1064);
nand U1280 (N_1280,N_1010,N_1084);
or U1281 (N_1281,N_1120,N_1061);
nor U1282 (N_1282,N_1136,N_1072);
or U1283 (N_1283,N_1014,N_1001);
nand U1284 (N_1284,N_1023,N_1109);
nor U1285 (N_1285,N_1133,N_1067);
or U1286 (N_1286,N_1114,N_1188);
nand U1287 (N_1287,N_1073,N_1116);
nor U1288 (N_1288,N_1048,N_1139);
nor U1289 (N_1289,N_1051,N_1177);
nand U1290 (N_1290,N_1017,N_1024);
nand U1291 (N_1291,N_1165,N_1138);
xnor U1292 (N_1292,N_1157,N_1094);
xnor U1293 (N_1293,N_1171,N_1176);
nand U1294 (N_1294,N_1004,N_1161);
and U1295 (N_1295,N_1131,N_1110);
and U1296 (N_1296,N_1075,N_1047);
nand U1297 (N_1297,N_1002,N_1081);
nand U1298 (N_1298,N_1186,N_1091);
nand U1299 (N_1299,N_1031,N_1197);
and U1300 (N_1300,N_1058,N_1105);
and U1301 (N_1301,N_1014,N_1152);
and U1302 (N_1302,N_1031,N_1141);
or U1303 (N_1303,N_1135,N_1046);
nand U1304 (N_1304,N_1166,N_1154);
and U1305 (N_1305,N_1155,N_1117);
or U1306 (N_1306,N_1046,N_1036);
nor U1307 (N_1307,N_1059,N_1159);
or U1308 (N_1308,N_1099,N_1114);
nor U1309 (N_1309,N_1163,N_1067);
and U1310 (N_1310,N_1109,N_1002);
nor U1311 (N_1311,N_1064,N_1068);
or U1312 (N_1312,N_1013,N_1119);
nor U1313 (N_1313,N_1158,N_1147);
nor U1314 (N_1314,N_1042,N_1017);
and U1315 (N_1315,N_1096,N_1145);
or U1316 (N_1316,N_1064,N_1115);
or U1317 (N_1317,N_1061,N_1064);
nand U1318 (N_1318,N_1166,N_1034);
and U1319 (N_1319,N_1182,N_1105);
or U1320 (N_1320,N_1141,N_1160);
and U1321 (N_1321,N_1037,N_1128);
nand U1322 (N_1322,N_1178,N_1025);
and U1323 (N_1323,N_1091,N_1143);
nor U1324 (N_1324,N_1001,N_1101);
nor U1325 (N_1325,N_1087,N_1140);
or U1326 (N_1326,N_1112,N_1149);
nor U1327 (N_1327,N_1032,N_1002);
nand U1328 (N_1328,N_1174,N_1042);
nor U1329 (N_1329,N_1141,N_1066);
or U1330 (N_1330,N_1181,N_1097);
or U1331 (N_1331,N_1191,N_1094);
and U1332 (N_1332,N_1115,N_1198);
nor U1333 (N_1333,N_1050,N_1192);
nor U1334 (N_1334,N_1088,N_1184);
nand U1335 (N_1335,N_1138,N_1073);
or U1336 (N_1336,N_1073,N_1081);
or U1337 (N_1337,N_1058,N_1010);
or U1338 (N_1338,N_1186,N_1077);
and U1339 (N_1339,N_1153,N_1044);
nand U1340 (N_1340,N_1195,N_1079);
nand U1341 (N_1341,N_1169,N_1094);
xor U1342 (N_1342,N_1171,N_1010);
nor U1343 (N_1343,N_1181,N_1087);
or U1344 (N_1344,N_1174,N_1062);
or U1345 (N_1345,N_1161,N_1088);
or U1346 (N_1346,N_1094,N_1168);
nand U1347 (N_1347,N_1152,N_1121);
nand U1348 (N_1348,N_1101,N_1156);
nand U1349 (N_1349,N_1052,N_1083);
nand U1350 (N_1350,N_1179,N_1134);
nor U1351 (N_1351,N_1103,N_1030);
nor U1352 (N_1352,N_1109,N_1106);
nor U1353 (N_1353,N_1141,N_1001);
and U1354 (N_1354,N_1124,N_1121);
or U1355 (N_1355,N_1011,N_1158);
and U1356 (N_1356,N_1068,N_1020);
nand U1357 (N_1357,N_1026,N_1122);
and U1358 (N_1358,N_1094,N_1060);
or U1359 (N_1359,N_1164,N_1001);
nor U1360 (N_1360,N_1185,N_1131);
and U1361 (N_1361,N_1001,N_1011);
nand U1362 (N_1362,N_1090,N_1061);
or U1363 (N_1363,N_1063,N_1074);
nor U1364 (N_1364,N_1133,N_1046);
or U1365 (N_1365,N_1126,N_1058);
nand U1366 (N_1366,N_1199,N_1070);
or U1367 (N_1367,N_1070,N_1149);
or U1368 (N_1368,N_1147,N_1020);
xor U1369 (N_1369,N_1068,N_1190);
or U1370 (N_1370,N_1080,N_1108);
nor U1371 (N_1371,N_1140,N_1062);
and U1372 (N_1372,N_1030,N_1037);
and U1373 (N_1373,N_1153,N_1081);
or U1374 (N_1374,N_1149,N_1175);
nand U1375 (N_1375,N_1139,N_1069);
nor U1376 (N_1376,N_1041,N_1169);
nor U1377 (N_1377,N_1009,N_1003);
and U1378 (N_1378,N_1111,N_1029);
and U1379 (N_1379,N_1151,N_1109);
nand U1380 (N_1380,N_1091,N_1073);
nor U1381 (N_1381,N_1060,N_1109);
or U1382 (N_1382,N_1135,N_1198);
or U1383 (N_1383,N_1172,N_1074);
or U1384 (N_1384,N_1005,N_1089);
or U1385 (N_1385,N_1042,N_1119);
and U1386 (N_1386,N_1130,N_1108);
nor U1387 (N_1387,N_1070,N_1090);
and U1388 (N_1388,N_1068,N_1039);
or U1389 (N_1389,N_1079,N_1017);
or U1390 (N_1390,N_1137,N_1096);
or U1391 (N_1391,N_1031,N_1026);
xnor U1392 (N_1392,N_1189,N_1012);
and U1393 (N_1393,N_1155,N_1191);
and U1394 (N_1394,N_1036,N_1128);
xor U1395 (N_1395,N_1161,N_1182);
nand U1396 (N_1396,N_1192,N_1153);
and U1397 (N_1397,N_1143,N_1119);
nand U1398 (N_1398,N_1137,N_1129);
or U1399 (N_1399,N_1192,N_1021);
and U1400 (N_1400,N_1294,N_1221);
or U1401 (N_1401,N_1325,N_1244);
xor U1402 (N_1402,N_1211,N_1274);
and U1403 (N_1403,N_1375,N_1347);
nand U1404 (N_1404,N_1355,N_1239);
and U1405 (N_1405,N_1372,N_1389);
nand U1406 (N_1406,N_1218,N_1309);
nor U1407 (N_1407,N_1227,N_1205);
or U1408 (N_1408,N_1271,N_1292);
nand U1409 (N_1409,N_1288,N_1395);
nand U1410 (N_1410,N_1224,N_1301);
and U1411 (N_1411,N_1258,N_1350);
nand U1412 (N_1412,N_1353,N_1393);
or U1413 (N_1413,N_1287,N_1275);
or U1414 (N_1414,N_1206,N_1201);
or U1415 (N_1415,N_1212,N_1380);
nand U1416 (N_1416,N_1366,N_1264);
and U1417 (N_1417,N_1386,N_1253);
nand U1418 (N_1418,N_1367,N_1270);
nor U1419 (N_1419,N_1236,N_1210);
or U1420 (N_1420,N_1250,N_1234);
or U1421 (N_1421,N_1373,N_1223);
nand U1422 (N_1422,N_1334,N_1396);
and U1423 (N_1423,N_1360,N_1310);
or U1424 (N_1424,N_1217,N_1313);
and U1425 (N_1425,N_1207,N_1352);
nor U1426 (N_1426,N_1315,N_1384);
or U1427 (N_1427,N_1241,N_1317);
and U1428 (N_1428,N_1358,N_1340);
and U1429 (N_1429,N_1243,N_1300);
and U1430 (N_1430,N_1220,N_1260);
nor U1431 (N_1431,N_1204,N_1302);
or U1432 (N_1432,N_1256,N_1346);
or U1433 (N_1433,N_1327,N_1262);
and U1434 (N_1434,N_1251,N_1277);
or U1435 (N_1435,N_1359,N_1318);
nor U1436 (N_1436,N_1216,N_1249);
and U1437 (N_1437,N_1208,N_1361);
xnor U1438 (N_1438,N_1235,N_1279);
nor U1439 (N_1439,N_1276,N_1293);
and U1440 (N_1440,N_1322,N_1265);
or U1441 (N_1441,N_1349,N_1338);
nand U1442 (N_1442,N_1398,N_1392);
nor U1443 (N_1443,N_1222,N_1383);
nand U1444 (N_1444,N_1286,N_1344);
and U1445 (N_1445,N_1328,N_1343);
nand U1446 (N_1446,N_1374,N_1291);
or U1447 (N_1447,N_1306,N_1254);
nand U1448 (N_1448,N_1336,N_1261);
nand U1449 (N_1449,N_1278,N_1378);
or U1450 (N_1450,N_1399,N_1385);
xnor U1451 (N_1451,N_1273,N_1297);
and U1452 (N_1452,N_1242,N_1363);
or U1453 (N_1453,N_1268,N_1345);
nand U1454 (N_1454,N_1357,N_1321);
nor U1455 (N_1455,N_1368,N_1365);
nand U1456 (N_1456,N_1226,N_1280);
and U1457 (N_1457,N_1296,N_1284);
and U1458 (N_1458,N_1305,N_1331);
or U1459 (N_1459,N_1298,N_1283);
nand U1460 (N_1460,N_1299,N_1289);
nor U1461 (N_1461,N_1219,N_1339);
xor U1462 (N_1462,N_1307,N_1387);
and U1463 (N_1463,N_1209,N_1379);
nand U1464 (N_1464,N_1203,N_1214);
nor U1465 (N_1465,N_1232,N_1285);
nor U1466 (N_1466,N_1319,N_1245);
nor U1467 (N_1467,N_1351,N_1369);
xor U1468 (N_1468,N_1337,N_1335);
nand U1469 (N_1469,N_1326,N_1202);
or U1470 (N_1470,N_1281,N_1213);
and U1471 (N_1471,N_1330,N_1238);
nor U1472 (N_1472,N_1370,N_1371);
or U1473 (N_1473,N_1329,N_1324);
and U1474 (N_1474,N_1377,N_1314);
and U1475 (N_1475,N_1381,N_1311);
nand U1476 (N_1476,N_1255,N_1397);
nand U1477 (N_1477,N_1303,N_1252);
or U1478 (N_1478,N_1229,N_1391);
nor U1479 (N_1479,N_1316,N_1290);
or U1480 (N_1480,N_1240,N_1247);
nand U1481 (N_1481,N_1354,N_1356);
or U1482 (N_1482,N_1257,N_1341);
or U1483 (N_1483,N_1332,N_1308);
nand U1484 (N_1484,N_1230,N_1233);
and U1485 (N_1485,N_1388,N_1342);
nand U1486 (N_1486,N_1362,N_1215);
nor U1487 (N_1487,N_1259,N_1246);
and U1488 (N_1488,N_1295,N_1320);
and U1489 (N_1489,N_1382,N_1228);
nand U1490 (N_1490,N_1231,N_1323);
or U1491 (N_1491,N_1282,N_1225);
or U1492 (N_1492,N_1267,N_1304);
and U1493 (N_1493,N_1376,N_1272);
or U1494 (N_1494,N_1237,N_1263);
or U1495 (N_1495,N_1364,N_1200);
nor U1496 (N_1496,N_1248,N_1266);
or U1497 (N_1497,N_1394,N_1348);
nor U1498 (N_1498,N_1312,N_1390);
nor U1499 (N_1499,N_1333,N_1269);
and U1500 (N_1500,N_1280,N_1370);
nand U1501 (N_1501,N_1326,N_1278);
or U1502 (N_1502,N_1287,N_1364);
or U1503 (N_1503,N_1380,N_1354);
and U1504 (N_1504,N_1331,N_1221);
or U1505 (N_1505,N_1208,N_1270);
nor U1506 (N_1506,N_1212,N_1228);
and U1507 (N_1507,N_1387,N_1393);
and U1508 (N_1508,N_1253,N_1362);
and U1509 (N_1509,N_1391,N_1219);
nand U1510 (N_1510,N_1282,N_1271);
nor U1511 (N_1511,N_1308,N_1333);
nor U1512 (N_1512,N_1394,N_1203);
nor U1513 (N_1513,N_1206,N_1308);
or U1514 (N_1514,N_1310,N_1353);
or U1515 (N_1515,N_1277,N_1362);
nand U1516 (N_1516,N_1301,N_1245);
and U1517 (N_1517,N_1240,N_1326);
nor U1518 (N_1518,N_1210,N_1311);
nand U1519 (N_1519,N_1382,N_1387);
nor U1520 (N_1520,N_1214,N_1264);
and U1521 (N_1521,N_1333,N_1354);
nor U1522 (N_1522,N_1304,N_1262);
nor U1523 (N_1523,N_1305,N_1217);
nand U1524 (N_1524,N_1386,N_1238);
nor U1525 (N_1525,N_1258,N_1333);
or U1526 (N_1526,N_1233,N_1245);
or U1527 (N_1527,N_1253,N_1214);
and U1528 (N_1528,N_1228,N_1276);
or U1529 (N_1529,N_1251,N_1261);
nor U1530 (N_1530,N_1377,N_1288);
nand U1531 (N_1531,N_1225,N_1258);
nor U1532 (N_1532,N_1370,N_1260);
nand U1533 (N_1533,N_1343,N_1322);
nor U1534 (N_1534,N_1368,N_1394);
nor U1535 (N_1535,N_1310,N_1279);
nor U1536 (N_1536,N_1346,N_1324);
nand U1537 (N_1537,N_1270,N_1330);
nor U1538 (N_1538,N_1228,N_1302);
or U1539 (N_1539,N_1359,N_1253);
and U1540 (N_1540,N_1241,N_1272);
or U1541 (N_1541,N_1236,N_1204);
xnor U1542 (N_1542,N_1289,N_1260);
nor U1543 (N_1543,N_1277,N_1208);
or U1544 (N_1544,N_1268,N_1373);
or U1545 (N_1545,N_1273,N_1359);
nand U1546 (N_1546,N_1242,N_1354);
or U1547 (N_1547,N_1207,N_1224);
xnor U1548 (N_1548,N_1267,N_1363);
and U1549 (N_1549,N_1248,N_1346);
nand U1550 (N_1550,N_1226,N_1233);
and U1551 (N_1551,N_1231,N_1318);
nand U1552 (N_1552,N_1203,N_1266);
nor U1553 (N_1553,N_1242,N_1323);
nand U1554 (N_1554,N_1258,N_1365);
or U1555 (N_1555,N_1362,N_1317);
and U1556 (N_1556,N_1281,N_1222);
or U1557 (N_1557,N_1389,N_1370);
nand U1558 (N_1558,N_1282,N_1248);
nor U1559 (N_1559,N_1352,N_1312);
and U1560 (N_1560,N_1384,N_1216);
and U1561 (N_1561,N_1329,N_1249);
and U1562 (N_1562,N_1337,N_1250);
or U1563 (N_1563,N_1261,N_1314);
nand U1564 (N_1564,N_1211,N_1243);
nor U1565 (N_1565,N_1296,N_1324);
and U1566 (N_1566,N_1299,N_1277);
nand U1567 (N_1567,N_1258,N_1251);
nand U1568 (N_1568,N_1371,N_1249);
nor U1569 (N_1569,N_1397,N_1211);
or U1570 (N_1570,N_1311,N_1382);
nor U1571 (N_1571,N_1209,N_1271);
and U1572 (N_1572,N_1354,N_1217);
nor U1573 (N_1573,N_1387,N_1319);
nor U1574 (N_1574,N_1234,N_1330);
and U1575 (N_1575,N_1377,N_1275);
nor U1576 (N_1576,N_1236,N_1263);
nand U1577 (N_1577,N_1223,N_1367);
or U1578 (N_1578,N_1303,N_1344);
or U1579 (N_1579,N_1308,N_1220);
nand U1580 (N_1580,N_1258,N_1257);
and U1581 (N_1581,N_1345,N_1323);
and U1582 (N_1582,N_1243,N_1293);
or U1583 (N_1583,N_1211,N_1363);
nor U1584 (N_1584,N_1311,N_1399);
and U1585 (N_1585,N_1249,N_1326);
xor U1586 (N_1586,N_1289,N_1348);
nand U1587 (N_1587,N_1382,N_1214);
nand U1588 (N_1588,N_1381,N_1286);
nand U1589 (N_1589,N_1398,N_1240);
nand U1590 (N_1590,N_1281,N_1214);
nor U1591 (N_1591,N_1336,N_1294);
or U1592 (N_1592,N_1321,N_1308);
or U1593 (N_1593,N_1213,N_1255);
nand U1594 (N_1594,N_1343,N_1281);
or U1595 (N_1595,N_1345,N_1364);
or U1596 (N_1596,N_1200,N_1385);
and U1597 (N_1597,N_1283,N_1263);
xnor U1598 (N_1598,N_1306,N_1379);
nand U1599 (N_1599,N_1281,N_1375);
and U1600 (N_1600,N_1481,N_1567);
nor U1601 (N_1601,N_1571,N_1591);
and U1602 (N_1602,N_1524,N_1553);
nor U1603 (N_1603,N_1476,N_1549);
nor U1604 (N_1604,N_1415,N_1435);
nand U1605 (N_1605,N_1523,N_1551);
nor U1606 (N_1606,N_1425,N_1426);
and U1607 (N_1607,N_1564,N_1525);
nand U1608 (N_1608,N_1593,N_1510);
nand U1609 (N_1609,N_1483,N_1474);
nor U1610 (N_1610,N_1556,N_1516);
nor U1611 (N_1611,N_1491,N_1460);
and U1612 (N_1612,N_1541,N_1423);
nor U1613 (N_1613,N_1503,N_1507);
or U1614 (N_1614,N_1436,N_1496);
xor U1615 (N_1615,N_1585,N_1506);
or U1616 (N_1616,N_1433,N_1440);
nor U1617 (N_1617,N_1498,N_1451);
and U1618 (N_1618,N_1467,N_1413);
or U1619 (N_1619,N_1478,N_1545);
xnor U1620 (N_1620,N_1522,N_1566);
and U1621 (N_1621,N_1400,N_1490);
nand U1622 (N_1622,N_1419,N_1495);
xnor U1623 (N_1623,N_1497,N_1493);
nor U1624 (N_1624,N_1530,N_1461);
or U1625 (N_1625,N_1442,N_1458);
nand U1626 (N_1626,N_1544,N_1464);
nor U1627 (N_1627,N_1465,N_1597);
nor U1628 (N_1628,N_1521,N_1534);
nor U1629 (N_1629,N_1470,N_1412);
nand U1630 (N_1630,N_1587,N_1552);
or U1631 (N_1631,N_1502,N_1573);
nor U1632 (N_1632,N_1428,N_1526);
nor U1633 (N_1633,N_1579,N_1456);
xor U1634 (N_1634,N_1529,N_1431);
or U1635 (N_1635,N_1462,N_1590);
nand U1636 (N_1636,N_1559,N_1475);
or U1637 (N_1637,N_1580,N_1518);
xnor U1638 (N_1638,N_1505,N_1535);
and U1639 (N_1639,N_1565,N_1404);
or U1640 (N_1640,N_1487,N_1512);
and U1641 (N_1641,N_1469,N_1560);
nor U1642 (N_1642,N_1595,N_1468);
nor U1643 (N_1643,N_1520,N_1517);
and U1644 (N_1644,N_1504,N_1427);
nand U1645 (N_1645,N_1546,N_1463);
nand U1646 (N_1646,N_1443,N_1508);
nand U1647 (N_1647,N_1482,N_1547);
and U1648 (N_1648,N_1448,N_1557);
nor U1649 (N_1649,N_1539,N_1537);
and U1650 (N_1650,N_1414,N_1485);
or U1651 (N_1651,N_1471,N_1430);
or U1652 (N_1652,N_1574,N_1411);
and U1653 (N_1653,N_1441,N_1527);
xor U1654 (N_1654,N_1501,N_1432);
nor U1655 (N_1655,N_1540,N_1420);
or U1656 (N_1656,N_1446,N_1429);
nor U1657 (N_1657,N_1438,N_1445);
nand U1658 (N_1658,N_1407,N_1548);
nand U1659 (N_1659,N_1437,N_1492);
nor U1660 (N_1660,N_1416,N_1554);
and U1661 (N_1661,N_1596,N_1499);
nand U1662 (N_1662,N_1582,N_1409);
and U1663 (N_1663,N_1577,N_1405);
nor U1664 (N_1664,N_1408,N_1439);
nor U1665 (N_1665,N_1533,N_1569);
nor U1666 (N_1666,N_1401,N_1417);
or U1667 (N_1667,N_1454,N_1570);
nor U1668 (N_1668,N_1418,N_1466);
or U1669 (N_1669,N_1459,N_1480);
nand U1670 (N_1670,N_1576,N_1402);
nand U1671 (N_1671,N_1403,N_1575);
nand U1672 (N_1672,N_1421,N_1538);
xor U1673 (N_1673,N_1449,N_1543);
or U1674 (N_1674,N_1588,N_1568);
nand U1675 (N_1675,N_1455,N_1584);
nand U1676 (N_1676,N_1477,N_1484);
and U1677 (N_1677,N_1550,N_1472);
and U1678 (N_1678,N_1558,N_1489);
and U1679 (N_1679,N_1542,N_1599);
nand U1680 (N_1680,N_1488,N_1422);
or U1681 (N_1681,N_1598,N_1594);
nor U1682 (N_1682,N_1447,N_1592);
nor U1683 (N_1683,N_1513,N_1452);
or U1684 (N_1684,N_1562,N_1532);
or U1685 (N_1685,N_1450,N_1434);
xnor U1686 (N_1686,N_1424,N_1457);
or U1687 (N_1687,N_1563,N_1486);
nor U1688 (N_1688,N_1586,N_1479);
nand U1689 (N_1689,N_1536,N_1519);
nand U1690 (N_1690,N_1531,N_1589);
and U1691 (N_1691,N_1453,N_1500);
and U1692 (N_1692,N_1572,N_1555);
nor U1693 (N_1693,N_1406,N_1444);
nor U1694 (N_1694,N_1494,N_1528);
nor U1695 (N_1695,N_1410,N_1511);
or U1696 (N_1696,N_1514,N_1581);
nor U1697 (N_1697,N_1515,N_1578);
and U1698 (N_1698,N_1561,N_1473);
nor U1699 (N_1699,N_1509,N_1583);
or U1700 (N_1700,N_1593,N_1514);
nand U1701 (N_1701,N_1516,N_1430);
or U1702 (N_1702,N_1403,N_1486);
or U1703 (N_1703,N_1449,N_1538);
nor U1704 (N_1704,N_1487,N_1547);
nand U1705 (N_1705,N_1431,N_1414);
and U1706 (N_1706,N_1440,N_1511);
or U1707 (N_1707,N_1539,N_1400);
nand U1708 (N_1708,N_1568,N_1489);
and U1709 (N_1709,N_1545,N_1537);
nor U1710 (N_1710,N_1409,N_1558);
nand U1711 (N_1711,N_1560,N_1503);
nand U1712 (N_1712,N_1555,N_1598);
nor U1713 (N_1713,N_1513,N_1563);
nor U1714 (N_1714,N_1582,N_1487);
or U1715 (N_1715,N_1400,N_1465);
and U1716 (N_1716,N_1539,N_1526);
or U1717 (N_1717,N_1456,N_1589);
or U1718 (N_1718,N_1447,N_1590);
or U1719 (N_1719,N_1584,N_1599);
nand U1720 (N_1720,N_1569,N_1424);
and U1721 (N_1721,N_1532,N_1498);
nor U1722 (N_1722,N_1569,N_1449);
or U1723 (N_1723,N_1432,N_1519);
nand U1724 (N_1724,N_1548,N_1523);
or U1725 (N_1725,N_1574,N_1433);
nor U1726 (N_1726,N_1406,N_1516);
nor U1727 (N_1727,N_1429,N_1416);
nand U1728 (N_1728,N_1564,N_1405);
or U1729 (N_1729,N_1550,N_1514);
or U1730 (N_1730,N_1537,N_1408);
nor U1731 (N_1731,N_1434,N_1574);
and U1732 (N_1732,N_1509,N_1494);
and U1733 (N_1733,N_1475,N_1508);
or U1734 (N_1734,N_1530,N_1455);
xor U1735 (N_1735,N_1423,N_1400);
nor U1736 (N_1736,N_1423,N_1586);
nor U1737 (N_1737,N_1574,N_1481);
and U1738 (N_1738,N_1556,N_1455);
nor U1739 (N_1739,N_1415,N_1462);
nand U1740 (N_1740,N_1451,N_1415);
and U1741 (N_1741,N_1480,N_1537);
xor U1742 (N_1742,N_1551,N_1449);
nand U1743 (N_1743,N_1440,N_1578);
or U1744 (N_1744,N_1440,N_1586);
and U1745 (N_1745,N_1514,N_1482);
nor U1746 (N_1746,N_1516,N_1415);
or U1747 (N_1747,N_1575,N_1471);
and U1748 (N_1748,N_1451,N_1540);
and U1749 (N_1749,N_1445,N_1467);
or U1750 (N_1750,N_1475,N_1565);
nor U1751 (N_1751,N_1403,N_1416);
nor U1752 (N_1752,N_1435,N_1527);
nand U1753 (N_1753,N_1437,N_1536);
nor U1754 (N_1754,N_1491,N_1572);
and U1755 (N_1755,N_1556,N_1401);
nand U1756 (N_1756,N_1482,N_1495);
and U1757 (N_1757,N_1405,N_1409);
and U1758 (N_1758,N_1584,N_1494);
nor U1759 (N_1759,N_1455,N_1462);
and U1760 (N_1760,N_1575,N_1596);
nand U1761 (N_1761,N_1528,N_1442);
nand U1762 (N_1762,N_1450,N_1565);
nand U1763 (N_1763,N_1517,N_1455);
nor U1764 (N_1764,N_1479,N_1560);
nor U1765 (N_1765,N_1493,N_1475);
or U1766 (N_1766,N_1451,N_1468);
nor U1767 (N_1767,N_1406,N_1421);
nand U1768 (N_1768,N_1553,N_1443);
or U1769 (N_1769,N_1510,N_1480);
nand U1770 (N_1770,N_1437,N_1561);
or U1771 (N_1771,N_1524,N_1456);
nand U1772 (N_1772,N_1438,N_1595);
nand U1773 (N_1773,N_1436,N_1585);
and U1774 (N_1774,N_1413,N_1526);
nor U1775 (N_1775,N_1457,N_1484);
or U1776 (N_1776,N_1469,N_1509);
and U1777 (N_1777,N_1448,N_1555);
nor U1778 (N_1778,N_1407,N_1554);
nand U1779 (N_1779,N_1442,N_1426);
nor U1780 (N_1780,N_1515,N_1583);
or U1781 (N_1781,N_1503,N_1578);
or U1782 (N_1782,N_1414,N_1481);
nor U1783 (N_1783,N_1429,N_1505);
or U1784 (N_1784,N_1458,N_1523);
and U1785 (N_1785,N_1593,N_1437);
and U1786 (N_1786,N_1563,N_1521);
nor U1787 (N_1787,N_1563,N_1588);
nand U1788 (N_1788,N_1437,N_1541);
nand U1789 (N_1789,N_1562,N_1534);
nor U1790 (N_1790,N_1458,N_1422);
nor U1791 (N_1791,N_1506,N_1556);
and U1792 (N_1792,N_1411,N_1450);
or U1793 (N_1793,N_1543,N_1478);
nand U1794 (N_1794,N_1449,N_1411);
nand U1795 (N_1795,N_1532,N_1507);
xor U1796 (N_1796,N_1587,N_1585);
nand U1797 (N_1797,N_1566,N_1467);
nand U1798 (N_1798,N_1456,N_1583);
nor U1799 (N_1799,N_1514,N_1568);
nor U1800 (N_1800,N_1758,N_1725);
or U1801 (N_1801,N_1666,N_1770);
or U1802 (N_1802,N_1647,N_1696);
nand U1803 (N_1803,N_1756,N_1761);
or U1804 (N_1804,N_1798,N_1730);
nand U1805 (N_1805,N_1786,N_1695);
and U1806 (N_1806,N_1659,N_1767);
and U1807 (N_1807,N_1775,N_1631);
nor U1808 (N_1808,N_1711,N_1755);
or U1809 (N_1809,N_1684,N_1637);
nor U1810 (N_1810,N_1656,N_1774);
nor U1811 (N_1811,N_1669,N_1621);
nor U1812 (N_1812,N_1672,N_1632);
nor U1813 (N_1813,N_1629,N_1752);
nand U1814 (N_1814,N_1733,N_1754);
nand U1815 (N_1815,N_1636,N_1705);
or U1816 (N_1816,N_1640,N_1764);
nand U1817 (N_1817,N_1757,N_1694);
and U1818 (N_1818,N_1735,N_1744);
nor U1819 (N_1819,N_1792,N_1617);
and U1820 (N_1820,N_1707,N_1793);
nand U1821 (N_1821,N_1759,N_1720);
nor U1822 (N_1822,N_1794,N_1797);
or U1823 (N_1823,N_1686,N_1700);
or U1824 (N_1824,N_1762,N_1748);
nor U1825 (N_1825,N_1788,N_1665);
nor U1826 (N_1826,N_1716,N_1655);
and U1827 (N_1827,N_1766,N_1677);
and U1828 (N_1828,N_1690,N_1732);
nor U1829 (N_1829,N_1685,N_1625);
nor U1830 (N_1830,N_1709,N_1602);
or U1831 (N_1831,N_1741,N_1615);
nand U1832 (N_1832,N_1646,N_1605);
or U1833 (N_1833,N_1664,N_1638);
or U1834 (N_1834,N_1708,N_1639);
or U1835 (N_1835,N_1603,N_1783);
and U1836 (N_1836,N_1739,N_1692);
nand U1837 (N_1837,N_1727,N_1723);
nand U1838 (N_1838,N_1743,N_1777);
and U1839 (N_1839,N_1791,N_1795);
or U1840 (N_1840,N_1628,N_1765);
nand U1841 (N_1841,N_1620,N_1771);
nand U1842 (N_1842,N_1643,N_1719);
or U1843 (N_1843,N_1648,N_1718);
nor U1844 (N_1844,N_1654,N_1616);
nor U1845 (N_1845,N_1769,N_1623);
nand U1846 (N_1846,N_1763,N_1658);
nor U1847 (N_1847,N_1633,N_1630);
nand U1848 (N_1848,N_1697,N_1751);
nand U1849 (N_1849,N_1745,N_1750);
or U1850 (N_1850,N_1731,N_1649);
or U1851 (N_1851,N_1657,N_1760);
or U1852 (N_1852,N_1671,N_1740);
nand U1853 (N_1853,N_1789,N_1753);
or U1854 (N_1854,N_1728,N_1737);
or U1855 (N_1855,N_1681,N_1699);
nor U1856 (N_1856,N_1679,N_1749);
or U1857 (N_1857,N_1722,N_1784);
or U1858 (N_1858,N_1676,N_1670);
nand U1859 (N_1859,N_1680,N_1703);
and U1860 (N_1860,N_1609,N_1641);
or U1861 (N_1861,N_1645,N_1683);
xnor U1862 (N_1862,N_1714,N_1606);
nor U1863 (N_1863,N_1607,N_1799);
nand U1864 (N_1864,N_1668,N_1611);
nand U1865 (N_1865,N_1678,N_1742);
and U1866 (N_1866,N_1702,N_1772);
or U1867 (N_1867,N_1626,N_1717);
or U1868 (N_1868,N_1776,N_1721);
or U1869 (N_1869,N_1673,N_1687);
or U1870 (N_1870,N_1601,N_1779);
and U1871 (N_1871,N_1701,N_1667);
nand U1872 (N_1872,N_1619,N_1746);
or U1873 (N_1873,N_1738,N_1693);
and U1874 (N_1874,N_1642,N_1780);
and U1875 (N_1875,N_1747,N_1773);
and U1876 (N_1876,N_1651,N_1663);
and U1877 (N_1877,N_1782,N_1618);
or U1878 (N_1878,N_1624,N_1614);
or U1879 (N_1879,N_1653,N_1644);
or U1880 (N_1880,N_1634,N_1710);
nand U1881 (N_1881,N_1787,N_1674);
nor U1882 (N_1882,N_1781,N_1778);
nor U1883 (N_1883,N_1712,N_1652);
or U1884 (N_1884,N_1698,N_1661);
and U1885 (N_1885,N_1662,N_1682);
nor U1886 (N_1886,N_1713,N_1715);
and U1887 (N_1887,N_1600,N_1688);
nand U1888 (N_1888,N_1724,N_1785);
or U1889 (N_1889,N_1691,N_1608);
nor U1890 (N_1890,N_1729,N_1768);
nor U1891 (N_1891,N_1704,N_1622);
nand U1892 (N_1892,N_1610,N_1627);
or U1893 (N_1893,N_1612,N_1613);
nand U1894 (N_1894,N_1736,N_1604);
and U1895 (N_1895,N_1796,N_1726);
or U1896 (N_1896,N_1689,N_1734);
and U1897 (N_1897,N_1706,N_1675);
or U1898 (N_1898,N_1790,N_1650);
or U1899 (N_1899,N_1635,N_1660);
and U1900 (N_1900,N_1622,N_1694);
nand U1901 (N_1901,N_1711,N_1703);
or U1902 (N_1902,N_1618,N_1683);
and U1903 (N_1903,N_1654,N_1799);
or U1904 (N_1904,N_1664,N_1735);
and U1905 (N_1905,N_1712,N_1772);
xor U1906 (N_1906,N_1631,N_1652);
and U1907 (N_1907,N_1611,N_1602);
nor U1908 (N_1908,N_1668,N_1616);
nand U1909 (N_1909,N_1754,N_1734);
and U1910 (N_1910,N_1749,N_1644);
and U1911 (N_1911,N_1736,N_1781);
nand U1912 (N_1912,N_1736,N_1724);
nand U1913 (N_1913,N_1730,N_1683);
nor U1914 (N_1914,N_1670,N_1602);
and U1915 (N_1915,N_1660,N_1676);
xor U1916 (N_1916,N_1783,N_1758);
and U1917 (N_1917,N_1735,N_1713);
or U1918 (N_1918,N_1608,N_1769);
nor U1919 (N_1919,N_1692,N_1751);
nor U1920 (N_1920,N_1748,N_1611);
and U1921 (N_1921,N_1694,N_1716);
or U1922 (N_1922,N_1677,N_1693);
or U1923 (N_1923,N_1792,N_1754);
nand U1924 (N_1924,N_1646,N_1708);
or U1925 (N_1925,N_1707,N_1686);
nor U1926 (N_1926,N_1704,N_1647);
and U1927 (N_1927,N_1691,N_1796);
xor U1928 (N_1928,N_1694,N_1639);
or U1929 (N_1929,N_1682,N_1702);
nand U1930 (N_1930,N_1644,N_1646);
or U1931 (N_1931,N_1686,N_1628);
or U1932 (N_1932,N_1797,N_1626);
nor U1933 (N_1933,N_1664,N_1665);
and U1934 (N_1934,N_1748,N_1775);
nand U1935 (N_1935,N_1711,N_1653);
and U1936 (N_1936,N_1763,N_1798);
and U1937 (N_1937,N_1701,N_1608);
or U1938 (N_1938,N_1737,N_1745);
nand U1939 (N_1939,N_1709,N_1771);
or U1940 (N_1940,N_1790,N_1609);
nor U1941 (N_1941,N_1721,N_1648);
and U1942 (N_1942,N_1772,N_1776);
xnor U1943 (N_1943,N_1691,N_1791);
nand U1944 (N_1944,N_1611,N_1793);
and U1945 (N_1945,N_1798,N_1771);
and U1946 (N_1946,N_1691,N_1609);
nor U1947 (N_1947,N_1707,N_1709);
xnor U1948 (N_1948,N_1615,N_1755);
nand U1949 (N_1949,N_1751,N_1672);
or U1950 (N_1950,N_1799,N_1636);
nand U1951 (N_1951,N_1659,N_1746);
or U1952 (N_1952,N_1729,N_1629);
or U1953 (N_1953,N_1627,N_1715);
or U1954 (N_1954,N_1787,N_1634);
nand U1955 (N_1955,N_1672,N_1699);
nand U1956 (N_1956,N_1643,N_1775);
xnor U1957 (N_1957,N_1700,N_1748);
and U1958 (N_1958,N_1646,N_1642);
nand U1959 (N_1959,N_1629,N_1686);
nand U1960 (N_1960,N_1758,N_1665);
or U1961 (N_1961,N_1730,N_1765);
nand U1962 (N_1962,N_1741,N_1749);
nand U1963 (N_1963,N_1637,N_1735);
or U1964 (N_1964,N_1726,N_1612);
nor U1965 (N_1965,N_1745,N_1680);
nand U1966 (N_1966,N_1728,N_1794);
or U1967 (N_1967,N_1761,N_1622);
and U1968 (N_1968,N_1674,N_1761);
or U1969 (N_1969,N_1743,N_1717);
and U1970 (N_1970,N_1640,N_1753);
nor U1971 (N_1971,N_1694,N_1671);
or U1972 (N_1972,N_1759,N_1794);
nor U1973 (N_1973,N_1790,N_1692);
nor U1974 (N_1974,N_1719,N_1623);
or U1975 (N_1975,N_1701,N_1653);
nand U1976 (N_1976,N_1653,N_1739);
nor U1977 (N_1977,N_1634,N_1677);
nor U1978 (N_1978,N_1646,N_1687);
and U1979 (N_1979,N_1727,N_1701);
nor U1980 (N_1980,N_1673,N_1757);
or U1981 (N_1981,N_1755,N_1771);
nor U1982 (N_1982,N_1744,N_1734);
or U1983 (N_1983,N_1720,N_1753);
and U1984 (N_1984,N_1611,N_1653);
nor U1985 (N_1985,N_1652,N_1743);
and U1986 (N_1986,N_1693,N_1782);
nor U1987 (N_1987,N_1610,N_1616);
and U1988 (N_1988,N_1626,N_1632);
or U1989 (N_1989,N_1676,N_1702);
and U1990 (N_1990,N_1732,N_1677);
nand U1991 (N_1991,N_1655,N_1615);
and U1992 (N_1992,N_1643,N_1705);
nor U1993 (N_1993,N_1701,N_1744);
nand U1994 (N_1994,N_1737,N_1668);
nor U1995 (N_1995,N_1788,N_1631);
or U1996 (N_1996,N_1636,N_1675);
nand U1997 (N_1997,N_1709,N_1740);
nand U1998 (N_1998,N_1770,N_1791);
or U1999 (N_1999,N_1671,N_1661);
nor U2000 (N_2000,N_1834,N_1852);
or U2001 (N_2001,N_1906,N_1871);
nor U2002 (N_2002,N_1987,N_1998);
or U2003 (N_2003,N_1831,N_1887);
nand U2004 (N_2004,N_1911,N_1919);
or U2005 (N_2005,N_1847,N_1805);
nor U2006 (N_2006,N_1809,N_1803);
or U2007 (N_2007,N_1974,N_1886);
or U2008 (N_2008,N_1840,N_1829);
nand U2009 (N_2009,N_1827,N_1913);
nor U2010 (N_2010,N_1877,N_1898);
or U2011 (N_2011,N_1873,N_1843);
nand U2012 (N_2012,N_1901,N_1930);
or U2013 (N_2013,N_1958,N_1909);
nand U2014 (N_2014,N_1836,N_1975);
nand U2015 (N_2015,N_1815,N_1949);
nor U2016 (N_2016,N_1994,N_1870);
nand U2017 (N_2017,N_1972,N_1957);
nand U2018 (N_2018,N_1828,N_1977);
nor U2019 (N_2019,N_1825,N_1981);
nand U2020 (N_2020,N_1948,N_1863);
or U2021 (N_2021,N_1874,N_1989);
nand U2022 (N_2022,N_1826,N_1850);
nand U2023 (N_2023,N_1893,N_1867);
nand U2024 (N_2024,N_1882,N_1967);
or U2025 (N_2025,N_1813,N_1978);
nand U2026 (N_2026,N_1822,N_1844);
xor U2027 (N_2027,N_1859,N_1858);
nor U2028 (N_2028,N_1985,N_1979);
nor U2029 (N_2029,N_1976,N_1854);
and U2030 (N_2030,N_1996,N_1971);
nand U2031 (N_2031,N_1885,N_1997);
or U2032 (N_2032,N_1936,N_1904);
nor U2033 (N_2033,N_1897,N_1889);
nand U2034 (N_2034,N_1969,N_1944);
and U2035 (N_2035,N_1865,N_1970);
and U2036 (N_2036,N_1895,N_1862);
and U2037 (N_2037,N_1954,N_1864);
and U2038 (N_2038,N_1907,N_1816);
nor U2039 (N_2039,N_1807,N_1992);
xnor U2040 (N_2040,N_1848,N_1851);
nand U2041 (N_2041,N_1879,N_1802);
or U2042 (N_2042,N_1888,N_1963);
and U2043 (N_2043,N_1892,N_1896);
nor U2044 (N_2044,N_1951,N_1835);
nor U2045 (N_2045,N_1926,N_1868);
or U2046 (N_2046,N_1960,N_1962);
or U2047 (N_2047,N_1925,N_1812);
nor U2048 (N_2048,N_1806,N_1853);
nand U2049 (N_2049,N_1929,N_1961);
and U2050 (N_2050,N_1839,N_1928);
and U2051 (N_2051,N_1846,N_1823);
nand U2052 (N_2052,N_1866,N_1821);
nand U2053 (N_2053,N_1938,N_1902);
or U2054 (N_2054,N_1855,N_1956);
and U2055 (N_2055,N_1966,N_1912);
or U2056 (N_2056,N_1965,N_1917);
or U2057 (N_2057,N_1861,N_1869);
nor U2058 (N_2058,N_1884,N_1991);
or U2059 (N_2059,N_1986,N_1801);
xor U2060 (N_2060,N_1933,N_1837);
xnor U2061 (N_2061,N_1832,N_1808);
nor U2062 (N_2062,N_1946,N_1817);
nor U2063 (N_2063,N_1814,N_1943);
nand U2064 (N_2064,N_1937,N_1953);
nand U2065 (N_2065,N_1939,N_1990);
or U2066 (N_2066,N_1924,N_1935);
and U2067 (N_2067,N_1880,N_1824);
nor U2068 (N_2068,N_1860,N_1940);
and U2069 (N_2069,N_1890,N_1915);
nor U2070 (N_2070,N_1804,N_1838);
or U2071 (N_2071,N_1820,N_1900);
nor U2072 (N_2072,N_1830,N_1841);
nor U2073 (N_2073,N_1811,N_1945);
nand U2074 (N_2074,N_1941,N_1983);
or U2075 (N_2075,N_1950,N_1923);
nor U2076 (N_2076,N_1947,N_1955);
or U2077 (N_2077,N_1968,N_1980);
and U2078 (N_2078,N_1856,N_1833);
and U2079 (N_2079,N_1927,N_1921);
nor U2080 (N_2080,N_1899,N_1872);
nand U2081 (N_2081,N_1800,N_1842);
and U2082 (N_2082,N_1932,N_1819);
or U2083 (N_2083,N_1875,N_1964);
and U2084 (N_2084,N_1952,N_1876);
nor U2085 (N_2085,N_1849,N_1883);
and U2086 (N_2086,N_1999,N_1995);
nor U2087 (N_2087,N_1903,N_1920);
and U2088 (N_2088,N_1905,N_1934);
or U2089 (N_2089,N_1973,N_1982);
and U2090 (N_2090,N_1931,N_1942);
and U2091 (N_2091,N_1894,N_1914);
nor U2092 (N_2092,N_1918,N_1845);
and U2093 (N_2093,N_1818,N_1891);
nand U2094 (N_2094,N_1878,N_1908);
nand U2095 (N_2095,N_1916,N_1810);
or U2096 (N_2096,N_1993,N_1959);
nor U2097 (N_2097,N_1984,N_1910);
and U2098 (N_2098,N_1922,N_1988);
and U2099 (N_2099,N_1881,N_1857);
and U2100 (N_2100,N_1943,N_1868);
and U2101 (N_2101,N_1982,N_1989);
nor U2102 (N_2102,N_1839,N_1822);
nand U2103 (N_2103,N_1994,N_1959);
nand U2104 (N_2104,N_1866,N_1898);
xor U2105 (N_2105,N_1822,N_1836);
and U2106 (N_2106,N_1873,N_1814);
or U2107 (N_2107,N_1998,N_1967);
and U2108 (N_2108,N_1993,N_1916);
nor U2109 (N_2109,N_1889,N_1998);
and U2110 (N_2110,N_1947,N_1894);
xnor U2111 (N_2111,N_1914,N_1877);
or U2112 (N_2112,N_1979,N_1852);
nand U2113 (N_2113,N_1943,N_1981);
nor U2114 (N_2114,N_1990,N_1996);
nor U2115 (N_2115,N_1996,N_1905);
or U2116 (N_2116,N_1957,N_1884);
nor U2117 (N_2117,N_1882,N_1975);
nand U2118 (N_2118,N_1895,N_1981);
or U2119 (N_2119,N_1803,N_1800);
nand U2120 (N_2120,N_1887,N_1911);
xnor U2121 (N_2121,N_1814,N_1827);
and U2122 (N_2122,N_1977,N_1946);
and U2123 (N_2123,N_1805,N_1862);
nand U2124 (N_2124,N_1802,N_1853);
xor U2125 (N_2125,N_1859,N_1930);
or U2126 (N_2126,N_1866,N_1801);
or U2127 (N_2127,N_1944,N_1978);
and U2128 (N_2128,N_1901,N_1892);
or U2129 (N_2129,N_1883,N_1854);
nor U2130 (N_2130,N_1890,N_1980);
xnor U2131 (N_2131,N_1853,N_1988);
nor U2132 (N_2132,N_1831,N_1926);
nand U2133 (N_2133,N_1823,N_1835);
nand U2134 (N_2134,N_1805,N_1879);
or U2135 (N_2135,N_1972,N_1898);
and U2136 (N_2136,N_1857,N_1847);
or U2137 (N_2137,N_1935,N_1954);
nor U2138 (N_2138,N_1857,N_1928);
or U2139 (N_2139,N_1880,N_1802);
and U2140 (N_2140,N_1937,N_1811);
nor U2141 (N_2141,N_1996,N_1980);
nor U2142 (N_2142,N_1977,N_1825);
nand U2143 (N_2143,N_1970,N_1851);
or U2144 (N_2144,N_1880,N_1957);
and U2145 (N_2145,N_1851,N_1961);
or U2146 (N_2146,N_1857,N_1905);
nand U2147 (N_2147,N_1891,N_1942);
or U2148 (N_2148,N_1950,N_1916);
or U2149 (N_2149,N_1839,N_1918);
nand U2150 (N_2150,N_1964,N_1916);
or U2151 (N_2151,N_1897,N_1904);
nor U2152 (N_2152,N_1852,N_1898);
and U2153 (N_2153,N_1854,N_1840);
or U2154 (N_2154,N_1906,N_1917);
or U2155 (N_2155,N_1905,N_1853);
nand U2156 (N_2156,N_1887,N_1823);
and U2157 (N_2157,N_1955,N_1923);
nor U2158 (N_2158,N_1990,N_1927);
and U2159 (N_2159,N_1858,N_1887);
and U2160 (N_2160,N_1893,N_1814);
nand U2161 (N_2161,N_1912,N_1885);
or U2162 (N_2162,N_1957,N_1873);
and U2163 (N_2163,N_1876,N_1811);
or U2164 (N_2164,N_1878,N_1987);
or U2165 (N_2165,N_1980,N_1835);
or U2166 (N_2166,N_1915,N_1844);
nand U2167 (N_2167,N_1863,N_1861);
nor U2168 (N_2168,N_1945,N_1998);
and U2169 (N_2169,N_1952,N_1860);
nand U2170 (N_2170,N_1821,N_1933);
xnor U2171 (N_2171,N_1829,N_1937);
nor U2172 (N_2172,N_1833,N_1844);
or U2173 (N_2173,N_1950,N_1867);
or U2174 (N_2174,N_1861,N_1828);
and U2175 (N_2175,N_1992,N_1877);
nor U2176 (N_2176,N_1921,N_1825);
nor U2177 (N_2177,N_1810,N_1975);
nand U2178 (N_2178,N_1907,N_1857);
nor U2179 (N_2179,N_1925,N_1936);
nand U2180 (N_2180,N_1983,N_1856);
nor U2181 (N_2181,N_1999,N_1861);
and U2182 (N_2182,N_1848,N_1991);
and U2183 (N_2183,N_1923,N_1825);
and U2184 (N_2184,N_1892,N_1990);
nor U2185 (N_2185,N_1902,N_1890);
nor U2186 (N_2186,N_1835,N_1981);
and U2187 (N_2187,N_1939,N_1804);
and U2188 (N_2188,N_1817,N_1935);
nand U2189 (N_2189,N_1937,N_1899);
nor U2190 (N_2190,N_1964,N_1913);
nand U2191 (N_2191,N_1948,N_1864);
or U2192 (N_2192,N_1880,N_1823);
or U2193 (N_2193,N_1885,N_1874);
nand U2194 (N_2194,N_1907,N_1908);
nand U2195 (N_2195,N_1886,N_1828);
and U2196 (N_2196,N_1801,N_1913);
or U2197 (N_2197,N_1834,N_1950);
nand U2198 (N_2198,N_1816,N_1831);
nor U2199 (N_2199,N_1949,N_1933);
nor U2200 (N_2200,N_2160,N_2031);
and U2201 (N_2201,N_2147,N_2073);
nor U2202 (N_2202,N_2064,N_2018);
or U2203 (N_2203,N_2047,N_2174);
or U2204 (N_2204,N_2187,N_2097);
nand U2205 (N_2205,N_2177,N_2185);
and U2206 (N_2206,N_2171,N_2036);
nand U2207 (N_2207,N_2077,N_2149);
nand U2208 (N_2208,N_2133,N_2045);
nor U2209 (N_2209,N_2119,N_2144);
or U2210 (N_2210,N_2078,N_2146);
nor U2211 (N_2211,N_2101,N_2090);
or U2212 (N_2212,N_2027,N_2014);
or U2213 (N_2213,N_2015,N_2143);
and U2214 (N_2214,N_2161,N_2030);
or U2215 (N_2215,N_2115,N_2121);
and U2216 (N_2216,N_2009,N_2085);
and U2217 (N_2217,N_2021,N_2059);
nor U2218 (N_2218,N_2100,N_2139);
nand U2219 (N_2219,N_2158,N_2175);
nand U2220 (N_2220,N_2191,N_2125);
or U2221 (N_2221,N_2098,N_2196);
and U2222 (N_2222,N_2010,N_2197);
or U2223 (N_2223,N_2041,N_2130);
or U2224 (N_2224,N_2103,N_2105);
nor U2225 (N_2225,N_2190,N_2000);
or U2226 (N_2226,N_2020,N_2194);
nor U2227 (N_2227,N_2028,N_2050);
or U2228 (N_2228,N_2019,N_2142);
and U2229 (N_2229,N_2003,N_2043);
nand U2230 (N_2230,N_2135,N_2172);
nand U2231 (N_2231,N_2181,N_2168);
nand U2232 (N_2232,N_2183,N_2094);
and U2233 (N_2233,N_2195,N_2192);
nand U2234 (N_2234,N_2163,N_2122);
and U2235 (N_2235,N_2040,N_2012);
or U2236 (N_2236,N_2092,N_2060);
xnor U2237 (N_2237,N_2004,N_2044);
and U2238 (N_2238,N_2046,N_2072);
and U2239 (N_2239,N_2083,N_2176);
nand U2240 (N_2240,N_2173,N_2082);
or U2241 (N_2241,N_2055,N_2076);
and U2242 (N_2242,N_2066,N_2179);
or U2243 (N_2243,N_2029,N_2091);
nor U2244 (N_2244,N_2025,N_2096);
nand U2245 (N_2245,N_2141,N_2071);
or U2246 (N_2246,N_2167,N_2129);
and U2247 (N_2247,N_2053,N_2153);
nand U2248 (N_2248,N_2049,N_2033);
nor U2249 (N_2249,N_2007,N_2169);
nand U2250 (N_2250,N_2037,N_2118);
or U2251 (N_2251,N_2107,N_2198);
and U2252 (N_2252,N_2013,N_2166);
and U2253 (N_2253,N_2038,N_2156);
nand U2254 (N_2254,N_2112,N_2017);
nand U2255 (N_2255,N_2126,N_2102);
nand U2256 (N_2256,N_2113,N_2128);
xor U2257 (N_2257,N_2095,N_2093);
nor U2258 (N_2258,N_2109,N_2131);
nand U2259 (N_2259,N_2032,N_2048);
xor U2260 (N_2260,N_2116,N_2150);
xor U2261 (N_2261,N_2088,N_2016);
xnor U2262 (N_2262,N_2188,N_2068);
and U2263 (N_2263,N_2123,N_2111);
and U2264 (N_2264,N_2124,N_2023);
and U2265 (N_2265,N_2104,N_2193);
nand U2266 (N_2266,N_2110,N_2106);
and U2267 (N_2267,N_2099,N_2070);
nor U2268 (N_2268,N_2054,N_2145);
nor U2269 (N_2269,N_2022,N_2108);
nand U2270 (N_2270,N_2001,N_2164);
nand U2271 (N_2271,N_2155,N_2136);
and U2272 (N_2272,N_2199,N_2127);
and U2273 (N_2273,N_2154,N_2114);
nand U2274 (N_2274,N_2006,N_2079);
and U2275 (N_2275,N_2042,N_2008);
or U2276 (N_2276,N_2165,N_2159);
nand U2277 (N_2277,N_2061,N_2157);
nor U2278 (N_2278,N_2180,N_2186);
nand U2279 (N_2279,N_2080,N_2069);
nor U2280 (N_2280,N_2184,N_2152);
and U2281 (N_2281,N_2002,N_2132);
and U2282 (N_2282,N_2034,N_2074);
and U2283 (N_2283,N_2067,N_2057);
or U2284 (N_2284,N_2035,N_2162);
or U2285 (N_2285,N_2065,N_2084);
or U2286 (N_2286,N_2170,N_2062);
or U2287 (N_2287,N_2140,N_2058);
nor U2288 (N_2288,N_2120,N_2051);
and U2289 (N_2289,N_2039,N_2117);
nand U2290 (N_2290,N_2011,N_2024);
and U2291 (N_2291,N_2134,N_2189);
nor U2292 (N_2292,N_2178,N_2087);
or U2293 (N_2293,N_2089,N_2182);
or U2294 (N_2294,N_2052,N_2075);
xor U2295 (N_2295,N_2137,N_2063);
or U2296 (N_2296,N_2151,N_2056);
nor U2297 (N_2297,N_2081,N_2026);
and U2298 (N_2298,N_2148,N_2005);
nand U2299 (N_2299,N_2086,N_2138);
nor U2300 (N_2300,N_2086,N_2011);
or U2301 (N_2301,N_2003,N_2041);
nor U2302 (N_2302,N_2066,N_2119);
and U2303 (N_2303,N_2197,N_2154);
xor U2304 (N_2304,N_2003,N_2088);
nand U2305 (N_2305,N_2178,N_2144);
nand U2306 (N_2306,N_2182,N_2129);
nor U2307 (N_2307,N_2051,N_2052);
nor U2308 (N_2308,N_2067,N_2029);
and U2309 (N_2309,N_2098,N_2174);
and U2310 (N_2310,N_2036,N_2099);
and U2311 (N_2311,N_2154,N_2138);
or U2312 (N_2312,N_2113,N_2041);
nor U2313 (N_2313,N_2162,N_2059);
and U2314 (N_2314,N_2021,N_2014);
nand U2315 (N_2315,N_2034,N_2190);
nor U2316 (N_2316,N_2177,N_2171);
nand U2317 (N_2317,N_2114,N_2182);
nand U2318 (N_2318,N_2114,N_2111);
nand U2319 (N_2319,N_2024,N_2018);
or U2320 (N_2320,N_2042,N_2047);
and U2321 (N_2321,N_2160,N_2155);
nand U2322 (N_2322,N_2052,N_2037);
nor U2323 (N_2323,N_2130,N_2002);
and U2324 (N_2324,N_2001,N_2093);
nor U2325 (N_2325,N_2026,N_2017);
nor U2326 (N_2326,N_2036,N_2192);
nand U2327 (N_2327,N_2195,N_2173);
and U2328 (N_2328,N_2087,N_2069);
and U2329 (N_2329,N_2044,N_2154);
nand U2330 (N_2330,N_2029,N_2083);
nand U2331 (N_2331,N_2133,N_2174);
or U2332 (N_2332,N_2102,N_2032);
or U2333 (N_2333,N_2150,N_2037);
nor U2334 (N_2334,N_2146,N_2162);
nor U2335 (N_2335,N_2134,N_2084);
nor U2336 (N_2336,N_2165,N_2095);
nor U2337 (N_2337,N_2122,N_2034);
nand U2338 (N_2338,N_2173,N_2152);
and U2339 (N_2339,N_2050,N_2052);
or U2340 (N_2340,N_2157,N_2103);
or U2341 (N_2341,N_2114,N_2136);
nor U2342 (N_2342,N_2137,N_2053);
nand U2343 (N_2343,N_2086,N_2161);
nor U2344 (N_2344,N_2101,N_2144);
nand U2345 (N_2345,N_2143,N_2041);
and U2346 (N_2346,N_2026,N_2181);
and U2347 (N_2347,N_2165,N_2005);
nand U2348 (N_2348,N_2055,N_2156);
and U2349 (N_2349,N_2136,N_2195);
or U2350 (N_2350,N_2020,N_2170);
nor U2351 (N_2351,N_2105,N_2017);
nor U2352 (N_2352,N_2032,N_2110);
and U2353 (N_2353,N_2178,N_2018);
nor U2354 (N_2354,N_2083,N_2136);
or U2355 (N_2355,N_2030,N_2005);
nor U2356 (N_2356,N_2129,N_2004);
xnor U2357 (N_2357,N_2122,N_2193);
nand U2358 (N_2358,N_2131,N_2047);
or U2359 (N_2359,N_2036,N_2176);
nand U2360 (N_2360,N_2000,N_2050);
and U2361 (N_2361,N_2199,N_2062);
nand U2362 (N_2362,N_2180,N_2028);
nor U2363 (N_2363,N_2161,N_2058);
or U2364 (N_2364,N_2057,N_2148);
or U2365 (N_2365,N_2199,N_2026);
or U2366 (N_2366,N_2052,N_2058);
nand U2367 (N_2367,N_2158,N_2019);
nor U2368 (N_2368,N_2170,N_2187);
or U2369 (N_2369,N_2018,N_2182);
or U2370 (N_2370,N_2172,N_2034);
nand U2371 (N_2371,N_2114,N_2088);
and U2372 (N_2372,N_2157,N_2092);
nand U2373 (N_2373,N_2054,N_2107);
or U2374 (N_2374,N_2075,N_2078);
nor U2375 (N_2375,N_2196,N_2198);
nand U2376 (N_2376,N_2169,N_2118);
or U2377 (N_2377,N_2129,N_2005);
and U2378 (N_2378,N_2151,N_2069);
or U2379 (N_2379,N_2078,N_2147);
nand U2380 (N_2380,N_2016,N_2118);
nor U2381 (N_2381,N_2023,N_2006);
and U2382 (N_2382,N_2160,N_2132);
nand U2383 (N_2383,N_2115,N_2168);
nand U2384 (N_2384,N_2157,N_2046);
or U2385 (N_2385,N_2058,N_2095);
nor U2386 (N_2386,N_2004,N_2144);
nor U2387 (N_2387,N_2152,N_2169);
or U2388 (N_2388,N_2024,N_2115);
nor U2389 (N_2389,N_2187,N_2089);
or U2390 (N_2390,N_2091,N_2060);
nor U2391 (N_2391,N_2128,N_2029);
or U2392 (N_2392,N_2147,N_2065);
nand U2393 (N_2393,N_2104,N_2163);
nor U2394 (N_2394,N_2178,N_2172);
nand U2395 (N_2395,N_2197,N_2013);
and U2396 (N_2396,N_2141,N_2131);
nand U2397 (N_2397,N_2007,N_2173);
nor U2398 (N_2398,N_2047,N_2121);
nand U2399 (N_2399,N_2010,N_2147);
nand U2400 (N_2400,N_2249,N_2312);
xor U2401 (N_2401,N_2376,N_2340);
nor U2402 (N_2402,N_2306,N_2203);
nor U2403 (N_2403,N_2315,N_2231);
nor U2404 (N_2404,N_2354,N_2360);
or U2405 (N_2405,N_2365,N_2269);
nand U2406 (N_2406,N_2343,N_2396);
and U2407 (N_2407,N_2273,N_2251);
or U2408 (N_2408,N_2261,N_2355);
nand U2409 (N_2409,N_2311,N_2244);
and U2410 (N_2410,N_2295,N_2260);
or U2411 (N_2411,N_2236,N_2363);
nor U2412 (N_2412,N_2252,N_2209);
nor U2413 (N_2413,N_2377,N_2243);
nand U2414 (N_2414,N_2335,N_2397);
or U2415 (N_2415,N_2290,N_2389);
nor U2416 (N_2416,N_2215,N_2283);
and U2417 (N_2417,N_2382,N_2374);
or U2418 (N_2418,N_2358,N_2264);
or U2419 (N_2419,N_2320,N_2324);
and U2420 (N_2420,N_2334,N_2395);
nor U2421 (N_2421,N_2388,N_2292);
and U2422 (N_2422,N_2341,N_2278);
or U2423 (N_2423,N_2275,N_2375);
nand U2424 (N_2424,N_2279,N_2228);
or U2425 (N_2425,N_2255,N_2351);
nor U2426 (N_2426,N_2391,N_2346);
and U2427 (N_2427,N_2232,N_2282);
and U2428 (N_2428,N_2366,N_2218);
and U2429 (N_2429,N_2336,N_2298);
nor U2430 (N_2430,N_2247,N_2380);
or U2431 (N_2431,N_2221,N_2390);
or U2432 (N_2432,N_2245,N_2299);
nand U2433 (N_2433,N_2222,N_2370);
or U2434 (N_2434,N_2270,N_2208);
and U2435 (N_2435,N_2263,N_2259);
nor U2436 (N_2436,N_2289,N_2210);
and U2437 (N_2437,N_2394,N_2268);
nand U2438 (N_2438,N_2226,N_2250);
nand U2439 (N_2439,N_2239,N_2300);
and U2440 (N_2440,N_2317,N_2265);
xnor U2441 (N_2441,N_2202,N_2297);
or U2442 (N_2442,N_2381,N_2353);
nor U2443 (N_2443,N_2308,N_2288);
nand U2444 (N_2444,N_2281,N_2387);
nor U2445 (N_2445,N_2213,N_2293);
nand U2446 (N_2446,N_2223,N_2371);
or U2447 (N_2447,N_2284,N_2227);
nand U2448 (N_2448,N_2313,N_2328);
nand U2449 (N_2449,N_2201,N_2330);
or U2450 (N_2450,N_2253,N_2305);
nor U2451 (N_2451,N_2323,N_2206);
nor U2452 (N_2452,N_2224,N_2230);
and U2453 (N_2453,N_2373,N_2339);
nand U2454 (N_2454,N_2383,N_2348);
xor U2455 (N_2455,N_2214,N_2256);
nor U2456 (N_2456,N_2307,N_2241);
and U2457 (N_2457,N_2296,N_2337);
and U2458 (N_2458,N_2258,N_2229);
or U2459 (N_2459,N_2357,N_2399);
nor U2460 (N_2460,N_2386,N_2310);
or U2461 (N_2461,N_2220,N_2359);
and U2462 (N_2462,N_2361,N_2217);
and U2463 (N_2463,N_2276,N_2302);
or U2464 (N_2464,N_2257,N_2267);
nor U2465 (N_2465,N_2356,N_2322);
nand U2466 (N_2466,N_2344,N_2392);
and U2467 (N_2467,N_2393,N_2338);
nand U2468 (N_2468,N_2368,N_2238);
and U2469 (N_2469,N_2347,N_2235);
or U2470 (N_2470,N_2325,N_2274);
nor U2471 (N_2471,N_2277,N_2364);
nor U2472 (N_2472,N_2205,N_2352);
and U2473 (N_2473,N_2349,N_2319);
or U2474 (N_2474,N_2372,N_2398);
nand U2475 (N_2475,N_2280,N_2384);
nor U2476 (N_2476,N_2329,N_2327);
nand U2477 (N_2477,N_2309,N_2291);
nor U2478 (N_2478,N_2219,N_2242);
nor U2479 (N_2479,N_2369,N_2240);
nor U2480 (N_2480,N_2204,N_2237);
nand U2481 (N_2481,N_2272,N_2379);
or U2482 (N_2482,N_2285,N_2314);
nand U2483 (N_2483,N_2316,N_2212);
and U2484 (N_2484,N_2378,N_2262);
nand U2485 (N_2485,N_2287,N_2233);
nor U2486 (N_2486,N_2207,N_2333);
or U2487 (N_2487,N_2286,N_2211);
nor U2488 (N_2488,N_2294,N_2304);
and U2489 (N_2489,N_2254,N_2321);
and U2490 (N_2490,N_2362,N_2350);
nor U2491 (N_2491,N_2342,N_2234);
or U2492 (N_2492,N_2200,N_2367);
and U2493 (N_2493,N_2266,N_2248);
nand U2494 (N_2494,N_2225,N_2326);
or U2495 (N_2495,N_2303,N_2385);
nand U2496 (N_2496,N_2345,N_2318);
and U2497 (N_2497,N_2246,N_2332);
or U2498 (N_2498,N_2271,N_2331);
nand U2499 (N_2499,N_2216,N_2301);
and U2500 (N_2500,N_2345,N_2272);
xor U2501 (N_2501,N_2309,N_2358);
nor U2502 (N_2502,N_2343,N_2381);
nor U2503 (N_2503,N_2365,N_2398);
or U2504 (N_2504,N_2255,N_2282);
and U2505 (N_2505,N_2279,N_2395);
xor U2506 (N_2506,N_2218,N_2283);
or U2507 (N_2507,N_2213,N_2359);
nand U2508 (N_2508,N_2329,N_2217);
or U2509 (N_2509,N_2358,N_2321);
nand U2510 (N_2510,N_2239,N_2291);
nor U2511 (N_2511,N_2289,N_2226);
or U2512 (N_2512,N_2392,N_2211);
or U2513 (N_2513,N_2352,N_2257);
or U2514 (N_2514,N_2260,N_2322);
nand U2515 (N_2515,N_2319,N_2397);
nand U2516 (N_2516,N_2366,N_2391);
and U2517 (N_2517,N_2223,N_2272);
nor U2518 (N_2518,N_2343,N_2304);
or U2519 (N_2519,N_2246,N_2346);
nand U2520 (N_2520,N_2368,N_2266);
or U2521 (N_2521,N_2392,N_2224);
nand U2522 (N_2522,N_2229,N_2204);
and U2523 (N_2523,N_2333,N_2234);
nor U2524 (N_2524,N_2294,N_2397);
or U2525 (N_2525,N_2294,N_2217);
nor U2526 (N_2526,N_2318,N_2326);
nor U2527 (N_2527,N_2208,N_2229);
nor U2528 (N_2528,N_2355,N_2310);
and U2529 (N_2529,N_2300,N_2286);
xnor U2530 (N_2530,N_2292,N_2399);
nor U2531 (N_2531,N_2213,N_2316);
and U2532 (N_2532,N_2273,N_2355);
or U2533 (N_2533,N_2309,N_2303);
nand U2534 (N_2534,N_2219,N_2277);
nand U2535 (N_2535,N_2386,N_2367);
or U2536 (N_2536,N_2269,N_2268);
nor U2537 (N_2537,N_2271,N_2356);
and U2538 (N_2538,N_2310,N_2229);
and U2539 (N_2539,N_2307,N_2231);
nor U2540 (N_2540,N_2347,N_2203);
or U2541 (N_2541,N_2307,N_2235);
nand U2542 (N_2542,N_2369,N_2345);
and U2543 (N_2543,N_2234,N_2313);
or U2544 (N_2544,N_2253,N_2306);
nor U2545 (N_2545,N_2233,N_2289);
nand U2546 (N_2546,N_2256,N_2227);
nor U2547 (N_2547,N_2246,N_2207);
or U2548 (N_2548,N_2279,N_2254);
nand U2549 (N_2549,N_2366,N_2359);
xnor U2550 (N_2550,N_2326,N_2204);
nor U2551 (N_2551,N_2366,N_2224);
nand U2552 (N_2552,N_2257,N_2322);
or U2553 (N_2553,N_2201,N_2283);
and U2554 (N_2554,N_2254,N_2269);
and U2555 (N_2555,N_2394,N_2250);
or U2556 (N_2556,N_2390,N_2281);
or U2557 (N_2557,N_2279,N_2262);
nand U2558 (N_2558,N_2285,N_2350);
nor U2559 (N_2559,N_2293,N_2223);
and U2560 (N_2560,N_2380,N_2342);
or U2561 (N_2561,N_2298,N_2288);
and U2562 (N_2562,N_2287,N_2384);
nor U2563 (N_2563,N_2242,N_2278);
nor U2564 (N_2564,N_2272,N_2385);
nor U2565 (N_2565,N_2298,N_2273);
or U2566 (N_2566,N_2375,N_2382);
and U2567 (N_2567,N_2276,N_2303);
and U2568 (N_2568,N_2245,N_2342);
or U2569 (N_2569,N_2243,N_2226);
nor U2570 (N_2570,N_2227,N_2207);
and U2571 (N_2571,N_2392,N_2383);
and U2572 (N_2572,N_2384,N_2274);
or U2573 (N_2573,N_2321,N_2310);
and U2574 (N_2574,N_2390,N_2238);
or U2575 (N_2575,N_2207,N_2284);
nor U2576 (N_2576,N_2261,N_2280);
and U2577 (N_2577,N_2337,N_2397);
and U2578 (N_2578,N_2293,N_2288);
xor U2579 (N_2579,N_2331,N_2246);
and U2580 (N_2580,N_2342,N_2239);
or U2581 (N_2581,N_2287,N_2302);
nand U2582 (N_2582,N_2345,N_2284);
and U2583 (N_2583,N_2252,N_2288);
nor U2584 (N_2584,N_2252,N_2254);
nand U2585 (N_2585,N_2324,N_2335);
nand U2586 (N_2586,N_2207,N_2362);
nand U2587 (N_2587,N_2293,N_2238);
and U2588 (N_2588,N_2223,N_2262);
nor U2589 (N_2589,N_2217,N_2385);
nand U2590 (N_2590,N_2353,N_2319);
or U2591 (N_2591,N_2250,N_2380);
or U2592 (N_2592,N_2264,N_2238);
or U2593 (N_2593,N_2284,N_2384);
nor U2594 (N_2594,N_2356,N_2249);
and U2595 (N_2595,N_2335,N_2280);
nor U2596 (N_2596,N_2398,N_2380);
or U2597 (N_2597,N_2316,N_2245);
or U2598 (N_2598,N_2242,N_2282);
and U2599 (N_2599,N_2263,N_2371);
nand U2600 (N_2600,N_2517,N_2452);
nor U2601 (N_2601,N_2453,N_2559);
or U2602 (N_2602,N_2518,N_2488);
and U2603 (N_2603,N_2465,N_2587);
nand U2604 (N_2604,N_2526,N_2525);
and U2605 (N_2605,N_2433,N_2573);
nor U2606 (N_2606,N_2532,N_2427);
nor U2607 (N_2607,N_2406,N_2473);
nor U2608 (N_2608,N_2597,N_2482);
nor U2609 (N_2609,N_2572,N_2520);
or U2610 (N_2610,N_2466,N_2591);
and U2611 (N_2611,N_2413,N_2435);
nand U2612 (N_2612,N_2451,N_2458);
or U2613 (N_2613,N_2567,N_2495);
or U2614 (N_2614,N_2471,N_2514);
and U2615 (N_2615,N_2533,N_2568);
nor U2616 (N_2616,N_2456,N_2483);
nand U2617 (N_2617,N_2565,N_2404);
nand U2618 (N_2618,N_2407,N_2580);
or U2619 (N_2619,N_2444,N_2554);
nand U2620 (N_2620,N_2599,N_2434);
nand U2621 (N_2621,N_2418,N_2592);
nor U2622 (N_2622,N_2472,N_2497);
and U2623 (N_2623,N_2474,N_2539);
or U2624 (N_2624,N_2460,N_2432);
nor U2625 (N_2625,N_2414,N_2566);
nor U2626 (N_2626,N_2551,N_2596);
and U2627 (N_2627,N_2498,N_2475);
nand U2628 (N_2628,N_2534,N_2513);
and U2629 (N_2629,N_2405,N_2535);
nand U2630 (N_2630,N_2457,N_2512);
or U2631 (N_2631,N_2503,N_2586);
nand U2632 (N_2632,N_2582,N_2481);
and U2633 (N_2633,N_2486,N_2505);
or U2634 (N_2634,N_2555,N_2529);
nor U2635 (N_2635,N_2410,N_2543);
and U2636 (N_2636,N_2480,N_2511);
nand U2637 (N_2637,N_2455,N_2593);
and U2638 (N_2638,N_2490,N_2544);
nor U2639 (N_2639,N_2504,N_2575);
xnor U2640 (N_2640,N_2428,N_2516);
or U2641 (N_2641,N_2564,N_2494);
nor U2642 (N_2642,N_2493,N_2485);
or U2643 (N_2643,N_2492,N_2546);
and U2644 (N_2644,N_2468,N_2469);
or U2645 (N_2645,N_2579,N_2524);
nand U2646 (N_2646,N_2430,N_2470);
nor U2647 (N_2647,N_2562,N_2431);
nor U2648 (N_2648,N_2550,N_2589);
nor U2649 (N_2649,N_2585,N_2416);
or U2650 (N_2650,N_2527,N_2522);
nand U2651 (N_2651,N_2436,N_2446);
nand U2652 (N_2652,N_2558,N_2496);
or U2653 (N_2653,N_2467,N_2426);
nor U2654 (N_2654,N_2438,N_2560);
nand U2655 (N_2655,N_2442,N_2561);
nand U2656 (N_2656,N_2464,N_2425);
and U2657 (N_2657,N_2443,N_2519);
and U2658 (N_2658,N_2508,N_2423);
or U2659 (N_2659,N_2581,N_2549);
nor U2660 (N_2660,N_2515,N_2584);
nand U2661 (N_2661,N_2487,N_2540);
and U2662 (N_2662,N_2429,N_2440);
and U2663 (N_2663,N_2548,N_2400);
or U2664 (N_2664,N_2476,N_2574);
and U2665 (N_2665,N_2437,N_2547);
or U2666 (N_2666,N_2403,N_2530);
or U2667 (N_2667,N_2552,N_2577);
xnor U2668 (N_2668,N_2510,N_2402);
xnor U2669 (N_2669,N_2594,N_2536);
or U2670 (N_2670,N_2588,N_2422);
and U2671 (N_2671,N_2528,N_2563);
nand U2672 (N_2672,N_2479,N_2509);
xnor U2673 (N_2673,N_2448,N_2598);
nor U2674 (N_2674,N_2489,N_2545);
and U2675 (N_2675,N_2478,N_2531);
and U2676 (N_2676,N_2537,N_2570);
or U2677 (N_2677,N_2409,N_2454);
nand U2678 (N_2678,N_2417,N_2556);
or U2679 (N_2679,N_2449,N_2507);
or U2680 (N_2680,N_2415,N_2459);
nand U2681 (N_2681,N_2500,N_2445);
or U2682 (N_2682,N_2408,N_2501);
nand U2683 (N_2683,N_2590,N_2424);
nor U2684 (N_2684,N_2595,N_2491);
nor U2685 (N_2685,N_2441,N_2502);
and U2686 (N_2686,N_2450,N_2553);
nor U2687 (N_2687,N_2484,N_2542);
or U2688 (N_2688,N_2538,N_2421);
nand U2689 (N_2689,N_2583,N_2569);
or U2690 (N_2690,N_2461,N_2477);
nor U2691 (N_2691,N_2521,N_2401);
nand U2692 (N_2692,N_2447,N_2419);
nand U2693 (N_2693,N_2506,N_2412);
or U2694 (N_2694,N_2499,N_2411);
or U2695 (N_2695,N_2571,N_2463);
nor U2696 (N_2696,N_2576,N_2541);
nor U2697 (N_2697,N_2523,N_2557);
nor U2698 (N_2698,N_2462,N_2439);
nor U2699 (N_2699,N_2578,N_2420);
nand U2700 (N_2700,N_2552,N_2587);
and U2701 (N_2701,N_2483,N_2513);
and U2702 (N_2702,N_2504,N_2570);
and U2703 (N_2703,N_2574,N_2412);
or U2704 (N_2704,N_2494,N_2451);
nand U2705 (N_2705,N_2404,N_2436);
or U2706 (N_2706,N_2507,N_2592);
or U2707 (N_2707,N_2520,N_2504);
nand U2708 (N_2708,N_2453,N_2502);
or U2709 (N_2709,N_2468,N_2493);
and U2710 (N_2710,N_2500,N_2588);
or U2711 (N_2711,N_2437,N_2471);
or U2712 (N_2712,N_2584,N_2433);
nand U2713 (N_2713,N_2418,N_2479);
nor U2714 (N_2714,N_2422,N_2480);
nand U2715 (N_2715,N_2459,N_2499);
or U2716 (N_2716,N_2490,N_2555);
or U2717 (N_2717,N_2412,N_2508);
nand U2718 (N_2718,N_2503,N_2594);
xor U2719 (N_2719,N_2529,N_2530);
or U2720 (N_2720,N_2450,N_2480);
nand U2721 (N_2721,N_2466,N_2479);
nor U2722 (N_2722,N_2465,N_2461);
and U2723 (N_2723,N_2481,N_2560);
nor U2724 (N_2724,N_2542,N_2482);
nand U2725 (N_2725,N_2404,N_2514);
and U2726 (N_2726,N_2421,N_2556);
nor U2727 (N_2727,N_2486,N_2430);
nand U2728 (N_2728,N_2591,N_2423);
and U2729 (N_2729,N_2480,N_2456);
and U2730 (N_2730,N_2469,N_2544);
or U2731 (N_2731,N_2527,N_2426);
nand U2732 (N_2732,N_2433,N_2557);
and U2733 (N_2733,N_2594,N_2466);
and U2734 (N_2734,N_2433,N_2477);
or U2735 (N_2735,N_2419,N_2450);
and U2736 (N_2736,N_2446,N_2503);
and U2737 (N_2737,N_2435,N_2426);
or U2738 (N_2738,N_2491,N_2417);
nand U2739 (N_2739,N_2588,N_2517);
and U2740 (N_2740,N_2485,N_2589);
and U2741 (N_2741,N_2479,N_2576);
nand U2742 (N_2742,N_2587,N_2507);
nor U2743 (N_2743,N_2470,N_2552);
and U2744 (N_2744,N_2519,N_2408);
nor U2745 (N_2745,N_2529,N_2518);
or U2746 (N_2746,N_2419,N_2515);
and U2747 (N_2747,N_2587,N_2563);
nand U2748 (N_2748,N_2544,N_2525);
nand U2749 (N_2749,N_2575,N_2437);
nor U2750 (N_2750,N_2418,N_2414);
or U2751 (N_2751,N_2563,N_2571);
nand U2752 (N_2752,N_2494,N_2421);
or U2753 (N_2753,N_2461,N_2578);
nand U2754 (N_2754,N_2581,N_2472);
nand U2755 (N_2755,N_2406,N_2534);
or U2756 (N_2756,N_2520,N_2481);
and U2757 (N_2757,N_2429,N_2546);
and U2758 (N_2758,N_2511,N_2561);
nand U2759 (N_2759,N_2484,N_2493);
or U2760 (N_2760,N_2452,N_2515);
and U2761 (N_2761,N_2411,N_2565);
and U2762 (N_2762,N_2580,N_2565);
and U2763 (N_2763,N_2580,N_2596);
nor U2764 (N_2764,N_2596,N_2427);
or U2765 (N_2765,N_2467,N_2451);
or U2766 (N_2766,N_2419,N_2467);
nor U2767 (N_2767,N_2579,N_2549);
and U2768 (N_2768,N_2572,N_2549);
or U2769 (N_2769,N_2426,N_2575);
nand U2770 (N_2770,N_2418,N_2445);
nand U2771 (N_2771,N_2463,N_2464);
and U2772 (N_2772,N_2566,N_2484);
nand U2773 (N_2773,N_2404,N_2500);
nand U2774 (N_2774,N_2407,N_2517);
nand U2775 (N_2775,N_2443,N_2457);
and U2776 (N_2776,N_2576,N_2484);
nand U2777 (N_2777,N_2578,N_2501);
nor U2778 (N_2778,N_2498,N_2456);
or U2779 (N_2779,N_2508,N_2450);
nand U2780 (N_2780,N_2581,N_2483);
or U2781 (N_2781,N_2529,N_2557);
or U2782 (N_2782,N_2536,N_2550);
or U2783 (N_2783,N_2494,N_2423);
and U2784 (N_2784,N_2508,N_2488);
nor U2785 (N_2785,N_2511,N_2578);
nor U2786 (N_2786,N_2567,N_2420);
nor U2787 (N_2787,N_2466,N_2434);
nor U2788 (N_2788,N_2575,N_2497);
nor U2789 (N_2789,N_2520,N_2424);
nand U2790 (N_2790,N_2574,N_2499);
and U2791 (N_2791,N_2518,N_2539);
xnor U2792 (N_2792,N_2540,N_2433);
nand U2793 (N_2793,N_2559,N_2546);
nor U2794 (N_2794,N_2459,N_2509);
nor U2795 (N_2795,N_2495,N_2528);
or U2796 (N_2796,N_2584,N_2496);
xor U2797 (N_2797,N_2593,N_2539);
nand U2798 (N_2798,N_2541,N_2480);
or U2799 (N_2799,N_2555,N_2444);
nand U2800 (N_2800,N_2661,N_2738);
nand U2801 (N_2801,N_2745,N_2788);
nor U2802 (N_2802,N_2743,N_2754);
and U2803 (N_2803,N_2773,N_2688);
nand U2804 (N_2804,N_2669,N_2622);
nor U2805 (N_2805,N_2652,N_2769);
or U2806 (N_2806,N_2741,N_2796);
and U2807 (N_2807,N_2670,N_2713);
nand U2808 (N_2808,N_2641,N_2785);
and U2809 (N_2809,N_2680,N_2799);
or U2810 (N_2810,N_2730,N_2763);
nand U2811 (N_2811,N_2710,N_2623);
or U2812 (N_2812,N_2752,N_2677);
nand U2813 (N_2813,N_2604,N_2748);
or U2814 (N_2814,N_2779,N_2697);
and U2815 (N_2815,N_2747,N_2784);
nor U2816 (N_2816,N_2735,N_2795);
and U2817 (N_2817,N_2750,N_2667);
and U2818 (N_2818,N_2665,N_2625);
and U2819 (N_2819,N_2690,N_2771);
or U2820 (N_2820,N_2718,N_2668);
nor U2821 (N_2821,N_2774,N_2689);
and U2822 (N_2822,N_2659,N_2644);
nor U2823 (N_2823,N_2778,N_2706);
nor U2824 (N_2824,N_2708,N_2662);
and U2825 (N_2825,N_2768,N_2603);
and U2826 (N_2826,N_2681,N_2618);
nor U2827 (N_2827,N_2602,N_2759);
or U2828 (N_2828,N_2649,N_2628);
nand U2829 (N_2829,N_2715,N_2617);
or U2830 (N_2830,N_2650,N_2627);
or U2831 (N_2831,N_2700,N_2631);
and U2832 (N_2832,N_2709,N_2639);
or U2833 (N_2833,N_2675,N_2701);
and U2834 (N_2834,N_2722,N_2762);
or U2835 (N_2835,N_2682,N_2655);
and U2836 (N_2836,N_2605,N_2653);
nand U2837 (N_2837,N_2601,N_2792);
or U2838 (N_2838,N_2736,N_2726);
and U2839 (N_2839,N_2698,N_2629);
nor U2840 (N_2840,N_2751,N_2685);
and U2841 (N_2841,N_2711,N_2787);
nor U2842 (N_2842,N_2699,N_2634);
or U2843 (N_2843,N_2610,N_2776);
or U2844 (N_2844,N_2672,N_2797);
nor U2845 (N_2845,N_2728,N_2648);
xor U2846 (N_2846,N_2615,N_2764);
nor U2847 (N_2847,N_2614,N_2737);
and U2848 (N_2848,N_2739,N_2782);
nor U2849 (N_2849,N_2758,N_2723);
nor U2850 (N_2850,N_2767,N_2645);
nor U2851 (N_2851,N_2635,N_2724);
nor U2852 (N_2852,N_2626,N_2714);
or U2853 (N_2853,N_2676,N_2760);
nand U2854 (N_2854,N_2798,N_2775);
nor U2855 (N_2855,N_2646,N_2766);
nand U2856 (N_2856,N_2679,N_2611);
nor U2857 (N_2857,N_2756,N_2647);
nand U2858 (N_2858,N_2633,N_2632);
nor U2859 (N_2859,N_2656,N_2664);
nand U2860 (N_2860,N_2640,N_2753);
and U2861 (N_2861,N_2624,N_2777);
and U2862 (N_2862,N_2761,N_2673);
nand U2863 (N_2863,N_2636,N_2686);
and U2864 (N_2864,N_2702,N_2732);
and U2865 (N_2865,N_2719,N_2794);
and U2866 (N_2866,N_2717,N_2733);
or U2867 (N_2867,N_2731,N_2740);
or U2868 (N_2868,N_2783,N_2674);
and U2869 (N_2869,N_2729,N_2654);
and U2870 (N_2870,N_2608,N_2630);
nor U2871 (N_2871,N_2660,N_2609);
nand U2872 (N_2872,N_2712,N_2725);
or U2873 (N_2873,N_2651,N_2613);
nand U2874 (N_2874,N_2720,N_2643);
nand U2875 (N_2875,N_2757,N_2683);
or U2876 (N_2876,N_2692,N_2791);
or U2877 (N_2877,N_2694,N_2642);
nor U2878 (N_2878,N_2606,N_2789);
or U2879 (N_2879,N_2707,N_2696);
nor U2880 (N_2880,N_2678,N_2607);
or U2881 (N_2881,N_2704,N_2727);
nor U2882 (N_2882,N_2620,N_2755);
nand U2883 (N_2883,N_2693,N_2721);
or U2884 (N_2884,N_2793,N_2781);
nor U2885 (N_2885,N_2749,N_2770);
nor U2886 (N_2886,N_2616,N_2612);
or U2887 (N_2887,N_2666,N_2684);
nor U2888 (N_2888,N_2742,N_2671);
nor U2889 (N_2889,N_2705,N_2687);
or U2890 (N_2890,N_2637,N_2786);
nand U2891 (N_2891,N_2600,N_2619);
and U2892 (N_2892,N_2772,N_2734);
nand U2893 (N_2893,N_2658,N_2638);
and U2894 (N_2894,N_2695,N_2703);
nor U2895 (N_2895,N_2716,N_2744);
or U2896 (N_2896,N_2691,N_2790);
and U2897 (N_2897,N_2621,N_2780);
or U2898 (N_2898,N_2663,N_2765);
nand U2899 (N_2899,N_2746,N_2657);
or U2900 (N_2900,N_2640,N_2618);
nor U2901 (N_2901,N_2639,N_2642);
or U2902 (N_2902,N_2660,N_2745);
nand U2903 (N_2903,N_2603,N_2695);
or U2904 (N_2904,N_2649,N_2721);
nand U2905 (N_2905,N_2670,N_2657);
or U2906 (N_2906,N_2609,N_2770);
and U2907 (N_2907,N_2756,N_2721);
and U2908 (N_2908,N_2622,N_2723);
and U2909 (N_2909,N_2643,N_2628);
and U2910 (N_2910,N_2635,N_2691);
or U2911 (N_2911,N_2608,N_2720);
xor U2912 (N_2912,N_2667,N_2681);
or U2913 (N_2913,N_2691,N_2641);
or U2914 (N_2914,N_2653,N_2780);
nor U2915 (N_2915,N_2609,N_2732);
nand U2916 (N_2916,N_2728,N_2714);
nand U2917 (N_2917,N_2729,N_2721);
nand U2918 (N_2918,N_2754,N_2742);
and U2919 (N_2919,N_2679,N_2608);
or U2920 (N_2920,N_2686,N_2668);
nand U2921 (N_2921,N_2724,N_2713);
and U2922 (N_2922,N_2654,N_2621);
nor U2923 (N_2923,N_2663,N_2716);
nor U2924 (N_2924,N_2634,N_2787);
and U2925 (N_2925,N_2745,N_2799);
nor U2926 (N_2926,N_2635,N_2799);
nor U2927 (N_2927,N_2685,N_2625);
nand U2928 (N_2928,N_2797,N_2612);
and U2929 (N_2929,N_2681,N_2727);
and U2930 (N_2930,N_2613,N_2654);
nand U2931 (N_2931,N_2620,N_2788);
and U2932 (N_2932,N_2614,N_2615);
nand U2933 (N_2933,N_2783,N_2799);
or U2934 (N_2934,N_2697,N_2683);
or U2935 (N_2935,N_2668,N_2779);
nor U2936 (N_2936,N_2743,N_2745);
or U2937 (N_2937,N_2729,N_2639);
nand U2938 (N_2938,N_2772,N_2690);
nand U2939 (N_2939,N_2708,N_2752);
nand U2940 (N_2940,N_2647,N_2678);
or U2941 (N_2941,N_2753,N_2627);
nor U2942 (N_2942,N_2652,N_2794);
and U2943 (N_2943,N_2714,N_2648);
or U2944 (N_2944,N_2736,N_2728);
and U2945 (N_2945,N_2786,N_2797);
nor U2946 (N_2946,N_2787,N_2705);
nand U2947 (N_2947,N_2647,N_2652);
or U2948 (N_2948,N_2692,N_2637);
nand U2949 (N_2949,N_2618,N_2788);
nor U2950 (N_2950,N_2787,N_2715);
nand U2951 (N_2951,N_2645,N_2623);
nor U2952 (N_2952,N_2611,N_2649);
xnor U2953 (N_2953,N_2742,N_2702);
or U2954 (N_2954,N_2619,N_2656);
or U2955 (N_2955,N_2642,N_2728);
nor U2956 (N_2956,N_2789,N_2779);
and U2957 (N_2957,N_2767,N_2631);
nand U2958 (N_2958,N_2633,N_2637);
nor U2959 (N_2959,N_2629,N_2745);
and U2960 (N_2960,N_2772,N_2610);
nor U2961 (N_2961,N_2760,N_2792);
nand U2962 (N_2962,N_2673,N_2785);
nor U2963 (N_2963,N_2620,N_2612);
nand U2964 (N_2964,N_2738,N_2784);
and U2965 (N_2965,N_2793,N_2617);
xnor U2966 (N_2966,N_2775,N_2779);
nor U2967 (N_2967,N_2787,N_2618);
nand U2968 (N_2968,N_2629,N_2797);
nor U2969 (N_2969,N_2754,N_2724);
and U2970 (N_2970,N_2764,N_2722);
nand U2971 (N_2971,N_2710,N_2618);
or U2972 (N_2972,N_2703,N_2681);
nor U2973 (N_2973,N_2721,N_2724);
or U2974 (N_2974,N_2609,N_2672);
nor U2975 (N_2975,N_2746,N_2768);
nand U2976 (N_2976,N_2718,N_2742);
nor U2977 (N_2977,N_2688,N_2798);
and U2978 (N_2978,N_2781,N_2644);
or U2979 (N_2979,N_2795,N_2779);
or U2980 (N_2980,N_2638,N_2722);
and U2981 (N_2981,N_2772,N_2641);
and U2982 (N_2982,N_2618,N_2778);
or U2983 (N_2983,N_2799,N_2632);
and U2984 (N_2984,N_2721,N_2688);
nand U2985 (N_2985,N_2701,N_2671);
nand U2986 (N_2986,N_2787,N_2636);
nand U2987 (N_2987,N_2704,N_2725);
or U2988 (N_2988,N_2644,N_2723);
or U2989 (N_2989,N_2741,N_2756);
nor U2990 (N_2990,N_2606,N_2652);
nor U2991 (N_2991,N_2767,N_2618);
nand U2992 (N_2992,N_2732,N_2630);
and U2993 (N_2993,N_2626,N_2758);
nor U2994 (N_2994,N_2786,N_2750);
nand U2995 (N_2995,N_2757,N_2705);
or U2996 (N_2996,N_2716,N_2781);
nor U2997 (N_2997,N_2719,N_2658);
and U2998 (N_2998,N_2620,N_2618);
nand U2999 (N_2999,N_2633,N_2636);
nor UO_0 (O_0,N_2957,N_2916);
nor UO_1 (O_1,N_2923,N_2959);
nor UO_2 (O_2,N_2911,N_2875);
nor UO_3 (O_3,N_2980,N_2895);
and UO_4 (O_4,N_2843,N_2878);
or UO_5 (O_5,N_2941,N_2823);
nor UO_6 (O_6,N_2931,N_2915);
nor UO_7 (O_7,N_2995,N_2889);
or UO_8 (O_8,N_2836,N_2805);
nand UO_9 (O_9,N_2954,N_2934);
nand UO_10 (O_10,N_2953,N_2863);
nand UO_11 (O_11,N_2929,N_2835);
nand UO_12 (O_12,N_2832,N_2833);
or UO_13 (O_13,N_2872,N_2873);
nand UO_14 (O_14,N_2879,N_2815);
nand UO_15 (O_15,N_2821,N_2838);
and UO_16 (O_16,N_2845,N_2985);
nor UO_17 (O_17,N_2860,N_2861);
xor UO_18 (O_18,N_2983,N_2856);
nand UO_19 (O_19,N_2877,N_2882);
and UO_20 (O_20,N_2884,N_2935);
nor UO_21 (O_21,N_2842,N_2822);
or UO_22 (O_22,N_2810,N_2930);
nand UO_23 (O_23,N_2939,N_2994);
or UO_24 (O_24,N_2853,N_2936);
nor UO_25 (O_25,N_2806,N_2852);
nor UO_26 (O_26,N_2865,N_2801);
and UO_27 (O_27,N_2909,N_2971);
and UO_28 (O_28,N_2844,N_2849);
nand UO_29 (O_29,N_2947,N_2892);
or UO_30 (O_30,N_2855,N_2904);
nor UO_31 (O_31,N_2829,N_2964);
xor UO_32 (O_32,N_2982,N_2928);
or UO_33 (O_33,N_2919,N_2898);
nand UO_34 (O_34,N_2816,N_2820);
nor UO_35 (O_35,N_2914,N_2968);
or UO_36 (O_36,N_2926,N_2803);
nor UO_37 (O_37,N_2808,N_2946);
and UO_38 (O_38,N_2937,N_2874);
and UO_39 (O_39,N_2961,N_2933);
nand UO_40 (O_40,N_2924,N_2812);
or UO_41 (O_41,N_2825,N_2988);
nand UO_42 (O_42,N_2973,N_2885);
and UO_43 (O_43,N_2862,N_2886);
and UO_44 (O_44,N_2893,N_2948);
nor UO_45 (O_45,N_2958,N_2920);
nor UO_46 (O_46,N_2972,N_2876);
nor UO_47 (O_47,N_2817,N_2918);
and UO_48 (O_48,N_2917,N_2827);
nand UO_49 (O_49,N_2925,N_2858);
nand UO_50 (O_50,N_2955,N_2999);
nor UO_51 (O_51,N_2970,N_2945);
and UO_52 (O_52,N_2870,N_2802);
and UO_53 (O_53,N_2976,N_2977);
nand UO_54 (O_54,N_2975,N_2819);
nor UO_55 (O_55,N_2901,N_2996);
nor UO_56 (O_56,N_2859,N_2997);
nand UO_57 (O_57,N_2944,N_2991);
xnor UO_58 (O_58,N_2866,N_2960);
or UO_59 (O_59,N_2981,N_2830);
nor UO_60 (O_60,N_2824,N_2956);
nor UO_61 (O_61,N_2967,N_2962);
nand UO_62 (O_62,N_2927,N_2834);
nand UO_63 (O_63,N_2902,N_2807);
nor UO_64 (O_64,N_2912,N_2896);
xor UO_65 (O_65,N_2891,N_2940);
or UO_66 (O_66,N_2813,N_2921);
or UO_67 (O_67,N_2831,N_2951);
or UO_68 (O_68,N_2890,N_2992);
nand UO_69 (O_69,N_2894,N_2974);
nor UO_70 (O_70,N_2857,N_2809);
or UO_71 (O_71,N_2989,N_2905);
and UO_72 (O_72,N_2839,N_2867);
or UO_73 (O_73,N_2932,N_2811);
nand UO_74 (O_74,N_2906,N_2984);
nor UO_75 (O_75,N_2850,N_2847);
nand UO_76 (O_76,N_2979,N_2907);
and UO_77 (O_77,N_2851,N_2903);
and UO_78 (O_78,N_2881,N_2804);
and UO_79 (O_79,N_2900,N_2952);
or UO_80 (O_80,N_2883,N_2887);
nand UO_81 (O_81,N_2826,N_2854);
nand UO_82 (O_82,N_2942,N_2897);
nor UO_83 (O_83,N_2943,N_2965);
or UO_84 (O_84,N_2828,N_2913);
and UO_85 (O_85,N_2969,N_2990);
or UO_86 (O_86,N_2922,N_2910);
nand UO_87 (O_87,N_2868,N_2848);
nor UO_88 (O_88,N_2841,N_2880);
and UO_89 (O_89,N_2993,N_2949);
nand UO_90 (O_90,N_2978,N_2986);
nand UO_91 (O_91,N_2963,N_2950);
and UO_92 (O_92,N_2871,N_2846);
nand UO_93 (O_93,N_2998,N_2837);
xnor UO_94 (O_94,N_2869,N_2888);
nor UO_95 (O_95,N_2818,N_2864);
nor UO_96 (O_96,N_2987,N_2899);
nand UO_97 (O_97,N_2966,N_2840);
nand UO_98 (O_98,N_2814,N_2800);
or UO_99 (O_99,N_2938,N_2908);
or UO_100 (O_100,N_2848,N_2881);
nor UO_101 (O_101,N_2856,N_2891);
nor UO_102 (O_102,N_2880,N_2901);
or UO_103 (O_103,N_2826,N_2990);
or UO_104 (O_104,N_2879,N_2974);
and UO_105 (O_105,N_2994,N_2997);
nor UO_106 (O_106,N_2867,N_2950);
nand UO_107 (O_107,N_2974,N_2979);
xnor UO_108 (O_108,N_2824,N_2892);
nor UO_109 (O_109,N_2880,N_2871);
and UO_110 (O_110,N_2930,N_2856);
xnor UO_111 (O_111,N_2935,N_2832);
or UO_112 (O_112,N_2803,N_2964);
xnor UO_113 (O_113,N_2874,N_2876);
and UO_114 (O_114,N_2922,N_2858);
nor UO_115 (O_115,N_2828,N_2839);
nand UO_116 (O_116,N_2802,N_2857);
or UO_117 (O_117,N_2953,N_2948);
and UO_118 (O_118,N_2983,N_2973);
and UO_119 (O_119,N_2985,N_2926);
nand UO_120 (O_120,N_2900,N_2995);
and UO_121 (O_121,N_2822,N_2833);
and UO_122 (O_122,N_2956,N_2911);
nor UO_123 (O_123,N_2835,N_2871);
or UO_124 (O_124,N_2855,N_2928);
and UO_125 (O_125,N_2920,N_2961);
nand UO_126 (O_126,N_2956,N_2866);
nor UO_127 (O_127,N_2978,N_2812);
nand UO_128 (O_128,N_2860,N_2864);
nand UO_129 (O_129,N_2962,N_2802);
or UO_130 (O_130,N_2926,N_2999);
nor UO_131 (O_131,N_2985,N_2916);
nand UO_132 (O_132,N_2833,N_2852);
nor UO_133 (O_133,N_2892,N_2911);
nor UO_134 (O_134,N_2995,N_2929);
and UO_135 (O_135,N_2878,N_2830);
or UO_136 (O_136,N_2826,N_2981);
or UO_137 (O_137,N_2940,N_2862);
or UO_138 (O_138,N_2858,N_2894);
or UO_139 (O_139,N_2950,N_2946);
and UO_140 (O_140,N_2978,N_2975);
nand UO_141 (O_141,N_2847,N_2887);
nor UO_142 (O_142,N_2918,N_2880);
nor UO_143 (O_143,N_2883,N_2856);
xor UO_144 (O_144,N_2906,N_2998);
or UO_145 (O_145,N_2918,N_2977);
and UO_146 (O_146,N_2943,N_2958);
nand UO_147 (O_147,N_2919,N_2999);
or UO_148 (O_148,N_2956,N_2980);
nor UO_149 (O_149,N_2957,N_2891);
nor UO_150 (O_150,N_2979,N_2842);
nor UO_151 (O_151,N_2922,N_2948);
and UO_152 (O_152,N_2864,N_2902);
nand UO_153 (O_153,N_2910,N_2801);
nor UO_154 (O_154,N_2857,N_2896);
and UO_155 (O_155,N_2906,N_2860);
and UO_156 (O_156,N_2806,N_2860);
or UO_157 (O_157,N_2861,N_2978);
or UO_158 (O_158,N_2905,N_2803);
and UO_159 (O_159,N_2890,N_2842);
or UO_160 (O_160,N_2858,N_2935);
nor UO_161 (O_161,N_2972,N_2978);
or UO_162 (O_162,N_2889,N_2819);
nor UO_163 (O_163,N_2821,N_2860);
nor UO_164 (O_164,N_2884,N_2817);
xnor UO_165 (O_165,N_2819,N_2988);
nand UO_166 (O_166,N_2841,N_2930);
xor UO_167 (O_167,N_2919,N_2904);
nand UO_168 (O_168,N_2926,N_2907);
or UO_169 (O_169,N_2884,N_2824);
nand UO_170 (O_170,N_2929,N_2990);
nand UO_171 (O_171,N_2957,N_2856);
or UO_172 (O_172,N_2855,N_2937);
nand UO_173 (O_173,N_2987,N_2893);
and UO_174 (O_174,N_2869,N_2921);
nand UO_175 (O_175,N_2847,N_2899);
or UO_176 (O_176,N_2908,N_2884);
and UO_177 (O_177,N_2922,N_2944);
nor UO_178 (O_178,N_2946,N_2949);
nor UO_179 (O_179,N_2824,N_2987);
and UO_180 (O_180,N_2981,N_2934);
and UO_181 (O_181,N_2930,N_2802);
nand UO_182 (O_182,N_2921,N_2965);
and UO_183 (O_183,N_2951,N_2936);
nor UO_184 (O_184,N_2974,N_2969);
nor UO_185 (O_185,N_2877,N_2939);
nand UO_186 (O_186,N_2918,N_2888);
nand UO_187 (O_187,N_2851,N_2834);
xor UO_188 (O_188,N_2910,N_2928);
or UO_189 (O_189,N_2956,N_2900);
nand UO_190 (O_190,N_2891,N_2824);
or UO_191 (O_191,N_2856,N_2892);
nand UO_192 (O_192,N_2839,N_2832);
and UO_193 (O_193,N_2842,N_2874);
or UO_194 (O_194,N_2882,N_2815);
and UO_195 (O_195,N_2843,N_2976);
nand UO_196 (O_196,N_2892,N_2842);
or UO_197 (O_197,N_2817,N_2827);
and UO_198 (O_198,N_2906,N_2963);
nor UO_199 (O_199,N_2822,N_2884);
and UO_200 (O_200,N_2925,N_2834);
nand UO_201 (O_201,N_2938,N_2910);
nand UO_202 (O_202,N_2978,N_2858);
or UO_203 (O_203,N_2885,N_2955);
nor UO_204 (O_204,N_2810,N_2968);
xor UO_205 (O_205,N_2933,N_2944);
nand UO_206 (O_206,N_2858,N_2860);
nor UO_207 (O_207,N_2968,N_2969);
nand UO_208 (O_208,N_2887,N_2858);
nor UO_209 (O_209,N_2914,N_2996);
xor UO_210 (O_210,N_2951,N_2983);
and UO_211 (O_211,N_2879,N_2919);
nor UO_212 (O_212,N_2957,N_2966);
and UO_213 (O_213,N_2816,N_2980);
and UO_214 (O_214,N_2918,N_2898);
or UO_215 (O_215,N_2808,N_2832);
and UO_216 (O_216,N_2857,N_2806);
and UO_217 (O_217,N_2848,N_2867);
xor UO_218 (O_218,N_2895,N_2914);
nor UO_219 (O_219,N_2804,N_2942);
nand UO_220 (O_220,N_2819,N_2849);
or UO_221 (O_221,N_2874,N_2873);
and UO_222 (O_222,N_2952,N_2997);
or UO_223 (O_223,N_2982,N_2824);
nand UO_224 (O_224,N_2931,N_2807);
and UO_225 (O_225,N_2814,N_2953);
nand UO_226 (O_226,N_2959,N_2965);
and UO_227 (O_227,N_2804,N_2938);
or UO_228 (O_228,N_2950,N_2888);
nand UO_229 (O_229,N_2964,N_2872);
or UO_230 (O_230,N_2828,N_2943);
and UO_231 (O_231,N_2822,N_2958);
and UO_232 (O_232,N_2942,N_2992);
and UO_233 (O_233,N_2893,N_2894);
xnor UO_234 (O_234,N_2859,N_2950);
nor UO_235 (O_235,N_2956,N_2860);
xnor UO_236 (O_236,N_2851,N_2873);
nand UO_237 (O_237,N_2916,N_2832);
nand UO_238 (O_238,N_2992,N_2948);
and UO_239 (O_239,N_2811,N_2871);
nand UO_240 (O_240,N_2988,N_2975);
or UO_241 (O_241,N_2803,N_2987);
nand UO_242 (O_242,N_2861,N_2825);
and UO_243 (O_243,N_2983,N_2869);
nand UO_244 (O_244,N_2955,N_2974);
nor UO_245 (O_245,N_2886,N_2879);
or UO_246 (O_246,N_2897,N_2855);
and UO_247 (O_247,N_2978,N_2955);
nand UO_248 (O_248,N_2847,N_2870);
nor UO_249 (O_249,N_2917,N_2844);
or UO_250 (O_250,N_2917,N_2936);
nand UO_251 (O_251,N_2966,N_2842);
or UO_252 (O_252,N_2897,N_2910);
and UO_253 (O_253,N_2960,N_2905);
xnor UO_254 (O_254,N_2874,N_2995);
nand UO_255 (O_255,N_2942,N_2959);
or UO_256 (O_256,N_2973,N_2988);
nor UO_257 (O_257,N_2821,N_2949);
xnor UO_258 (O_258,N_2816,N_2981);
nand UO_259 (O_259,N_2807,N_2894);
or UO_260 (O_260,N_2914,N_2995);
or UO_261 (O_261,N_2871,N_2980);
nand UO_262 (O_262,N_2923,N_2850);
and UO_263 (O_263,N_2929,N_2824);
nor UO_264 (O_264,N_2924,N_2988);
nand UO_265 (O_265,N_2963,N_2816);
nand UO_266 (O_266,N_2886,N_2875);
nand UO_267 (O_267,N_2906,N_2897);
or UO_268 (O_268,N_2986,N_2829);
nor UO_269 (O_269,N_2877,N_2983);
nor UO_270 (O_270,N_2999,N_2997);
or UO_271 (O_271,N_2930,N_2986);
and UO_272 (O_272,N_2961,N_2899);
nand UO_273 (O_273,N_2817,N_2984);
and UO_274 (O_274,N_2986,N_2849);
or UO_275 (O_275,N_2994,N_2918);
or UO_276 (O_276,N_2849,N_2880);
and UO_277 (O_277,N_2839,N_2897);
and UO_278 (O_278,N_2918,N_2945);
nand UO_279 (O_279,N_2957,N_2890);
nor UO_280 (O_280,N_2801,N_2905);
nor UO_281 (O_281,N_2818,N_2909);
and UO_282 (O_282,N_2958,N_2947);
nor UO_283 (O_283,N_2867,N_2925);
nor UO_284 (O_284,N_2981,N_2896);
and UO_285 (O_285,N_2854,N_2902);
and UO_286 (O_286,N_2863,N_2835);
and UO_287 (O_287,N_2955,N_2891);
nor UO_288 (O_288,N_2980,N_2869);
nor UO_289 (O_289,N_2999,N_2911);
and UO_290 (O_290,N_2967,N_2934);
or UO_291 (O_291,N_2919,N_2810);
nor UO_292 (O_292,N_2866,N_2992);
or UO_293 (O_293,N_2801,N_2915);
or UO_294 (O_294,N_2974,N_2902);
nor UO_295 (O_295,N_2885,N_2968);
nand UO_296 (O_296,N_2945,N_2968);
nor UO_297 (O_297,N_2882,N_2896);
and UO_298 (O_298,N_2835,N_2866);
nand UO_299 (O_299,N_2821,N_2867);
nor UO_300 (O_300,N_2882,N_2917);
or UO_301 (O_301,N_2922,N_2896);
nor UO_302 (O_302,N_2966,N_2905);
or UO_303 (O_303,N_2905,N_2808);
and UO_304 (O_304,N_2949,N_2858);
or UO_305 (O_305,N_2883,N_2898);
and UO_306 (O_306,N_2945,N_2859);
nand UO_307 (O_307,N_2835,N_2839);
and UO_308 (O_308,N_2983,N_2985);
nor UO_309 (O_309,N_2857,N_2943);
or UO_310 (O_310,N_2861,N_2911);
and UO_311 (O_311,N_2810,N_2887);
nand UO_312 (O_312,N_2987,N_2815);
nand UO_313 (O_313,N_2945,N_2949);
and UO_314 (O_314,N_2917,N_2855);
or UO_315 (O_315,N_2864,N_2947);
nand UO_316 (O_316,N_2882,N_2800);
nand UO_317 (O_317,N_2952,N_2912);
nand UO_318 (O_318,N_2868,N_2936);
or UO_319 (O_319,N_2809,N_2933);
xor UO_320 (O_320,N_2986,N_2917);
nand UO_321 (O_321,N_2876,N_2925);
or UO_322 (O_322,N_2864,N_2823);
xnor UO_323 (O_323,N_2906,N_2802);
or UO_324 (O_324,N_2951,N_2913);
or UO_325 (O_325,N_2832,N_2813);
nor UO_326 (O_326,N_2844,N_2897);
nor UO_327 (O_327,N_2838,N_2855);
or UO_328 (O_328,N_2869,N_2949);
nor UO_329 (O_329,N_2942,N_2812);
and UO_330 (O_330,N_2996,N_2984);
or UO_331 (O_331,N_2913,N_2999);
or UO_332 (O_332,N_2947,N_2878);
nand UO_333 (O_333,N_2895,N_2849);
nor UO_334 (O_334,N_2997,N_2906);
or UO_335 (O_335,N_2857,N_2963);
nor UO_336 (O_336,N_2806,N_2921);
or UO_337 (O_337,N_2837,N_2871);
nand UO_338 (O_338,N_2922,N_2981);
or UO_339 (O_339,N_2832,N_2941);
nand UO_340 (O_340,N_2980,N_2859);
and UO_341 (O_341,N_2804,N_2852);
nand UO_342 (O_342,N_2928,N_2806);
nand UO_343 (O_343,N_2809,N_2938);
nor UO_344 (O_344,N_2984,N_2942);
and UO_345 (O_345,N_2901,N_2832);
nor UO_346 (O_346,N_2888,N_2861);
nor UO_347 (O_347,N_2877,N_2819);
nand UO_348 (O_348,N_2869,N_2909);
or UO_349 (O_349,N_2810,N_2844);
nand UO_350 (O_350,N_2876,N_2835);
or UO_351 (O_351,N_2805,N_2849);
or UO_352 (O_352,N_2822,N_2974);
and UO_353 (O_353,N_2871,N_2869);
nor UO_354 (O_354,N_2834,N_2972);
nand UO_355 (O_355,N_2843,N_2983);
nor UO_356 (O_356,N_2953,N_2932);
or UO_357 (O_357,N_2933,N_2887);
nand UO_358 (O_358,N_2987,N_2921);
or UO_359 (O_359,N_2904,N_2936);
and UO_360 (O_360,N_2875,N_2927);
nor UO_361 (O_361,N_2938,N_2848);
xor UO_362 (O_362,N_2927,N_2867);
or UO_363 (O_363,N_2941,N_2967);
nand UO_364 (O_364,N_2993,N_2862);
or UO_365 (O_365,N_2840,N_2932);
and UO_366 (O_366,N_2887,N_2812);
nor UO_367 (O_367,N_2888,N_2914);
nand UO_368 (O_368,N_2995,N_2808);
nor UO_369 (O_369,N_2996,N_2909);
nor UO_370 (O_370,N_2834,N_2828);
or UO_371 (O_371,N_2942,N_2836);
nor UO_372 (O_372,N_2983,N_2977);
nand UO_373 (O_373,N_2929,N_2811);
and UO_374 (O_374,N_2992,N_2954);
and UO_375 (O_375,N_2823,N_2909);
and UO_376 (O_376,N_2930,N_2832);
and UO_377 (O_377,N_2871,N_2899);
nand UO_378 (O_378,N_2996,N_2845);
nand UO_379 (O_379,N_2943,N_2833);
nor UO_380 (O_380,N_2893,N_2962);
nand UO_381 (O_381,N_2826,N_2985);
and UO_382 (O_382,N_2979,N_2977);
or UO_383 (O_383,N_2866,N_2865);
nand UO_384 (O_384,N_2838,N_2926);
nor UO_385 (O_385,N_2877,N_2911);
nand UO_386 (O_386,N_2922,N_2998);
nor UO_387 (O_387,N_2858,N_2951);
and UO_388 (O_388,N_2804,N_2901);
nand UO_389 (O_389,N_2888,N_2854);
nor UO_390 (O_390,N_2866,N_2890);
and UO_391 (O_391,N_2874,N_2825);
nor UO_392 (O_392,N_2957,N_2886);
and UO_393 (O_393,N_2902,N_2917);
nor UO_394 (O_394,N_2978,N_2841);
nor UO_395 (O_395,N_2996,N_2994);
or UO_396 (O_396,N_2864,N_2870);
and UO_397 (O_397,N_2918,N_2961);
nand UO_398 (O_398,N_2802,N_2807);
and UO_399 (O_399,N_2809,N_2855);
nor UO_400 (O_400,N_2901,N_2936);
or UO_401 (O_401,N_2807,N_2850);
nor UO_402 (O_402,N_2897,N_2931);
nor UO_403 (O_403,N_2918,N_2811);
nand UO_404 (O_404,N_2990,N_2978);
nand UO_405 (O_405,N_2972,N_2870);
and UO_406 (O_406,N_2949,N_2847);
nand UO_407 (O_407,N_2965,N_2983);
nor UO_408 (O_408,N_2859,N_2959);
and UO_409 (O_409,N_2847,N_2934);
nor UO_410 (O_410,N_2852,N_2801);
xnor UO_411 (O_411,N_2942,N_2951);
and UO_412 (O_412,N_2863,N_2939);
nor UO_413 (O_413,N_2946,N_2983);
and UO_414 (O_414,N_2919,N_2859);
nand UO_415 (O_415,N_2999,N_2855);
or UO_416 (O_416,N_2954,N_2817);
nand UO_417 (O_417,N_2843,N_2861);
and UO_418 (O_418,N_2848,N_2927);
nor UO_419 (O_419,N_2810,N_2806);
nor UO_420 (O_420,N_2905,N_2825);
nor UO_421 (O_421,N_2826,N_2917);
or UO_422 (O_422,N_2904,N_2979);
or UO_423 (O_423,N_2971,N_2951);
nand UO_424 (O_424,N_2812,N_2973);
nand UO_425 (O_425,N_2972,N_2857);
nor UO_426 (O_426,N_2822,N_2855);
nand UO_427 (O_427,N_2959,N_2986);
and UO_428 (O_428,N_2840,N_2950);
and UO_429 (O_429,N_2981,N_2953);
nor UO_430 (O_430,N_2980,N_2951);
nand UO_431 (O_431,N_2852,N_2932);
and UO_432 (O_432,N_2926,N_2983);
nor UO_433 (O_433,N_2944,N_2813);
and UO_434 (O_434,N_2882,N_2837);
or UO_435 (O_435,N_2869,N_2995);
nand UO_436 (O_436,N_2847,N_2834);
and UO_437 (O_437,N_2932,N_2931);
and UO_438 (O_438,N_2982,N_2884);
nor UO_439 (O_439,N_2838,N_2852);
nand UO_440 (O_440,N_2946,N_2836);
nor UO_441 (O_441,N_2829,N_2887);
and UO_442 (O_442,N_2865,N_2974);
or UO_443 (O_443,N_2820,N_2984);
nor UO_444 (O_444,N_2990,N_2859);
or UO_445 (O_445,N_2860,N_2835);
and UO_446 (O_446,N_2965,N_2859);
and UO_447 (O_447,N_2825,N_2922);
and UO_448 (O_448,N_2933,N_2996);
nand UO_449 (O_449,N_2942,N_2912);
nand UO_450 (O_450,N_2995,N_2926);
nor UO_451 (O_451,N_2913,N_2858);
nand UO_452 (O_452,N_2949,N_2865);
or UO_453 (O_453,N_2804,N_2808);
nand UO_454 (O_454,N_2818,N_2955);
or UO_455 (O_455,N_2862,N_2835);
nor UO_456 (O_456,N_2872,N_2939);
nor UO_457 (O_457,N_2928,N_2942);
nand UO_458 (O_458,N_2976,N_2889);
nand UO_459 (O_459,N_2933,N_2829);
or UO_460 (O_460,N_2993,N_2912);
nand UO_461 (O_461,N_2939,N_2985);
nand UO_462 (O_462,N_2855,N_2987);
and UO_463 (O_463,N_2889,N_2932);
nor UO_464 (O_464,N_2967,N_2909);
nor UO_465 (O_465,N_2843,N_2923);
nand UO_466 (O_466,N_2980,N_2836);
nand UO_467 (O_467,N_2934,N_2900);
or UO_468 (O_468,N_2848,N_2933);
and UO_469 (O_469,N_2904,N_2809);
or UO_470 (O_470,N_2939,N_2915);
nor UO_471 (O_471,N_2963,N_2949);
and UO_472 (O_472,N_2846,N_2963);
nand UO_473 (O_473,N_2823,N_2938);
or UO_474 (O_474,N_2894,N_2988);
nand UO_475 (O_475,N_2960,N_2974);
or UO_476 (O_476,N_2866,N_2979);
and UO_477 (O_477,N_2970,N_2915);
nand UO_478 (O_478,N_2936,N_2964);
or UO_479 (O_479,N_2800,N_2937);
and UO_480 (O_480,N_2810,N_2993);
nand UO_481 (O_481,N_2860,N_2886);
nor UO_482 (O_482,N_2830,N_2816);
or UO_483 (O_483,N_2960,N_2977);
nand UO_484 (O_484,N_2859,N_2928);
or UO_485 (O_485,N_2840,N_2842);
or UO_486 (O_486,N_2972,N_2929);
nor UO_487 (O_487,N_2832,N_2855);
nand UO_488 (O_488,N_2902,N_2945);
nor UO_489 (O_489,N_2970,N_2932);
nor UO_490 (O_490,N_2970,N_2999);
and UO_491 (O_491,N_2811,N_2801);
or UO_492 (O_492,N_2947,N_2896);
nor UO_493 (O_493,N_2975,N_2930);
nor UO_494 (O_494,N_2973,N_2840);
or UO_495 (O_495,N_2966,N_2833);
nand UO_496 (O_496,N_2949,N_2897);
and UO_497 (O_497,N_2824,N_2974);
nor UO_498 (O_498,N_2832,N_2806);
and UO_499 (O_499,N_2988,N_2940);
endmodule