module basic_2000_20000_2500_5_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1804,In_758);
or U1 (N_1,In_1915,In_1101);
nor U2 (N_2,In_178,In_856);
and U3 (N_3,In_1218,In_904);
nor U4 (N_4,In_215,In_1470);
nor U5 (N_5,In_1515,In_1333);
nor U6 (N_6,In_366,In_297);
nor U7 (N_7,In_888,In_770);
or U8 (N_8,In_1388,In_145);
or U9 (N_9,In_112,In_59);
nor U10 (N_10,In_1638,In_263);
or U11 (N_11,In_1625,In_572);
xor U12 (N_12,In_532,In_1053);
or U13 (N_13,In_325,In_910);
and U14 (N_14,In_1921,In_703);
nand U15 (N_15,In_1807,In_933);
nor U16 (N_16,In_642,In_1773);
or U17 (N_17,In_1262,In_1257);
xnor U18 (N_18,In_378,In_1203);
and U19 (N_19,In_1310,In_818);
nand U20 (N_20,In_460,In_1635);
nand U21 (N_21,In_1761,In_1661);
and U22 (N_22,In_567,In_622);
nand U23 (N_23,In_508,In_260);
or U24 (N_24,In_339,In_1819);
nand U25 (N_25,In_1327,In_1621);
and U26 (N_26,In_1589,In_1489);
or U27 (N_27,In_810,In_1681);
or U28 (N_28,In_182,In_1545);
nor U29 (N_29,In_1579,In_323);
and U30 (N_30,In_1781,In_531);
nand U31 (N_31,In_1837,In_1948);
or U32 (N_32,In_39,In_38);
xor U33 (N_33,In_1528,In_1085);
and U34 (N_34,In_851,In_95);
nor U35 (N_35,In_1194,In_461);
nand U36 (N_36,In_1147,In_1021);
and U37 (N_37,In_1757,In_43);
nor U38 (N_38,In_1318,In_432);
and U39 (N_39,In_1936,In_1389);
and U40 (N_40,In_1994,In_1288);
or U41 (N_41,In_1825,In_1441);
or U42 (N_42,In_1302,In_131);
and U43 (N_43,In_1364,In_418);
and U44 (N_44,In_354,In_393);
or U45 (N_45,In_1598,In_887);
and U46 (N_46,In_189,In_971);
xor U47 (N_47,In_1970,In_850);
nand U48 (N_48,In_1393,In_1444);
or U49 (N_49,In_1006,In_1407);
or U50 (N_50,In_1971,In_1743);
or U51 (N_51,In_1356,In_53);
nor U52 (N_52,In_363,In_493);
xnor U53 (N_53,In_1337,In_1093);
or U54 (N_54,In_1365,In_561);
nand U55 (N_55,In_1496,In_753);
nand U56 (N_56,In_1843,In_190);
or U57 (N_57,In_1069,In_1602);
nor U58 (N_58,In_292,In_1737);
nand U59 (N_59,In_945,In_184);
and U60 (N_60,In_458,In_1062);
or U61 (N_61,In_259,In_161);
xor U62 (N_62,In_605,In_246);
xor U63 (N_63,In_601,In_64);
nor U64 (N_64,In_1520,In_1749);
and U65 (N_65,In_149,In_1325);
or U66 (N_66,In_1672,In_1537);
or U67 (N_67,In_333,In_537);
and U68 (N_68,In_1692,In_1111);
nor U69 (N_69,In_1308,In_1228);
and U70 (N_70,In_592,In_1173);
or U71 (N_71,In_1135,In_828);
and U72 (N_72,In_673,In_1384);
nor U73 (N_73,In_84,In_750);
or U74 (N_74,In_1840,In_879);
nand U75 (N_75,In_29,In_1964);
nand U76 (N_76,In_1078,In_594);
or U77 (N_77,In_1096,In_580);
or U78 (N_78,In_421,In_1392);
nand U79 (N_79,In_1829,In_152);
or U80 (N_80,In_132,In_1774);
nand U81 (N_81,In_1720,In_1335);
nor U82 (N_82,In_1517,In_586);
nor U83 (N_83,In_637,In_644);
or U84 (N_84,In_610,In_1400);
and U85 (N_85,In_502,In_1801);
and U86 (N_86,In_1766,In_369);
nor U87 (N_87,In_1883,In_443);
nand U88 (N_88,In_1614,In_898);
nor U89 (N_89,In_1273,In_1090);
nor U90 (N_90,In_880,In_1243);
nor U91 (N_91,In_1726,In_1500);
nor U92 (N_92,In_1097,In_1495);
nand U93 (N_93,In_869,In_852);
xor U94 (N_94,In_1009,In_1282);
and U95 (N_95,In_1949,In_1490);
nand U96 (N_96,In_72,In_788);
or U97 (N_97,In_66,In_547);
and U98 (N_98,In_221,In_1331);
or U99 (N_99,In_353,In_1468);
xnor U100 (N_100,In_490,In_652);
xor U101 (N_101,In_1751,In_1975);
or U102 (N_102,In_1982,In_1769);
nor U103 (N_103,In_1787,In_831);
and U104 (N_104,In_1080,In_1952);
xnor U105 (N_105,In_1362,In_1212);
xnor U106 (N_106,In_96,In_1951);
xnor U107 (N_107,In_714,In_1865);
nor U108 (N_108,In_1013,In_992);
nor U109 (N_109,In_1172,In_188);
and U110 (N_110,In_1906,In_1011);
nand U111 (N_111,In_650,In_437);
nand U112 (N_112,In_1518,In_370);
or U113 (N_113,In_481,In_157);
nand U114 (N_114,In_839,In_118);
nor U115 (N_115,In_206,In_338);
nand U116 (N_116,In_842,In_272);
nand U117 (N_117,In_1633,In_1597);
or U118 (N_118,In_204,In_247);
nor U119 (N_119,In_902,In_1986);
nand U120 (N_120,In_12,In_543);
nor U121 (N_121,In_924,In_294);
nor U122 (N_122,In_81,In_1667);
and U123 (N_123,In_242,In_829);
or U124 (N_124,In_1358,In_577);
or U125 (N_125,In_290,In_239);
xor U126 (N_126,In_1455,In_168);
nand U127 (N_127,In_1121,In_1143);
xor U128 (N_128,In_14,In_1838);
nand U129 (N_129,In_316,In_931);
or U130 (N_130,In_1103,In_628);
xnor U131 (N_131,In_611,In_466);
or U132 (N_132,In_1245,In_558);
nor U133 (N_133,In_684,In_1059);
or U134 (N_134,In_1999,In_254);
nand U135 (N_135,In_185,In_997);
or U136 (N_136,In_1516,In_312);
and U137 (N_137,In_1151,In_863);
and U138 (N_138,In_1776,In_546);
or U139 (N_139,In_698,In_730);
xor U140 (N_140,In_49,In_1313);
and U141 (N_141,In_394,In_1467);
and U142 (N_142,In_146,In_1759);
or U143 (N_143,In_1442,In_1736);
nand U144 (N_144,In_667,In_262);
and U145 (N_145,In_494,In_1847);
and U146 (N_146,In_1217,In_225);
nor U147 (N_147,In_1409,In_860);
or U148 (N_148,In_1966,In_467);
nor U149 (N_149,In_1158,In_1108);
or U150 (N_150,In_1839,In_666);
or U151 (N_151,In_659,In_76);
nor U152 (N_152,In_1593,In_1312);
nand U153 (N_153,In_731,In_1521);
or U154 (N_154,In_1000,In_177);
or U155 (N_155,In_1895,In_1943);
or U156 (N_156,In_1694,In_791);
or U157 (N_157,In_47,In_1463);
xnor U158 (N_158,In_173,In_1664);
nand U159 (N_159,In_1872,In_471);
and U160 (N_160,In_1081,In_680);
and U161 (N_161,In_1146,In_1691);
and U162 (N_162,In_195,In_1709);
nor U163 (N_163,In_261,In_885);
and U164 (N_164,In_1535,In_520);
and U165 (N_165,In_193,In_1512);
nand U166 (N_166,In_1131,In_656);
nand U167 (N_167,In_1969,In_277);
and U168 (N_168,In_1904,In_562);
nand U169 (N_169,In_1042,In_1268);
nor U170 (N_170,In_1411,In_317);
nor U171 (N_171,In_1957,In_91);
nand U172 (N_172,In_83,In_187);
or U173 (N_173,In_395,In_115);
nand U174 (N_174,In_687,In_1821);
xor U175 (N_175,In_1511,In_958);
nor U176 (N_176,In_535,In_506);
and U177 (N_177,In_1946,In_1645);
or U178 (N_178,In_462,In_1192);
nand U179 (N_179,In_1197,In_1580);
xnor U180 (N_180,In_351,In_745);
or U181 (N_181,In_1811,In_1035);
nand U182 (N_182,In_1875,In_20);
or U183 (N_183,In_1486,In_1693);
or U184 (N_184,In_111,In_1247);
and U185 (N_185,In_1647,In_526);
nor U186 (N_186,In_889,In_534);
and U187 (N_187,In_275,In_1064);
or U188 (N_188,In_1808,In_805);
nand U189 (N_189,In_1851,In_1695);
or U190 (N_190,In_1261,In_1809);
and U191 (N_191,In_1513,In_1834);
nand U192 (N_192,In_1762,In_415);
xnor U193 (N_193,In_915,In_191);
nor U194 (N_194,In_991,In_138);
nand U195 (N_195,In_1287,In_383);
or U196 (N_196,In_1134,In_1507);
nor U197 (N_197,In_1534,In_942);
and U198 (N_198,In_1935,In_947);
nor U199 (N_199,In_1629,In_1918);
or U200 (N_200,In_253,In_1188);
and U201 (N_201,In_151,In_1576);
xor U202 (N_202,In_1290,In_9);
and U203 (N_203,In_960,In_278);
or U204 (N_204,In_1316,In_241);
and U205 (N_205,In_1213,In_454);
or U206 (N_206,In_160,In_1706);
nand U207 (N_207,In_783,In_304);
and U208 (N_208,In_1497,In_607);
nor U209 (N_209,In_1219,In_307);
or U210 (N_210,In_273,In_735);
nand U211 (N_211,In_796,In_1690);
nor U212 (N_212,In_1399,In_1697);
or U213 (N_213,In_205,In_308);
and U214 (N_214,In_1403,In_268);
xor U215 (N_215,In_1896,In_930);
and U216 (N_216,In_1648,In_597);
xnor U217 (N_217,In_1958,In_1433);
xor U218 (N_218,In_781,In_736);
nor U219 (N_219,In_1230,In_614);
and U220 (N_220,In_983,In_104);
and U221 (N_221,In_86,In_1586);
xor U222 (N_222,In_1169,In_1996);
nor U223 (N_223,In_231,In_596);
xor U224 (N_224,In_590,In_1443);
or U225 (N_225,In_1562,In_1917);
or U226 (N_226,In_374,In_1014);
xnor U227 (N_227,In_925,In_1723);
or U228 (N_228,In_1123,In_105);
or U229 (N_229,In_192,In_1307);
or U230 (N_230,In_229,In_1270);
and U231 (N_231,In_625,In_1742);
xor U232 (N_232,In_61,In_202);
or U233 (N_233,In_858,In_1439);
or U234 (N_234,In_385,In_1300);
nor U235 (N_235,In_384,In_1272);
or U236 (N_236,In_1233,In_1833);
nor U237 (N_237,In_566,In_1007);
and U238 (N_238,In_517,In_1005);
or U239 (N_239,In_1799,In_1201);
xnor U240 (N_240,In_1551,In_1832);
nand U241 (N_241,In_1630,In_1073);
and U242 (N_242,In_1494,In_1022);
or U243 (N_243,In_1155,In_778);
or U244 (N_244,In_1481,In_1133);
and U245 (N_245,In_1378,In_108);
or U246 (N_246,In_34,In_1395);
nand U247 (N_247,In_1920,In_961);
or U248 (N_248,In_1698,In_1279);
or U249 (N_249,In_761,In_99);
xnor U250 (N_250,In_1871,In_677);
and U251 (N_251,In_413,In_1050);
or U252 (N_252,In_347,In_470);
nor U253 (N_253,In_1772,In_134);
nand U254 (N_254,In_1755,In_1499);
and U255 (N_255,In_1707,In_1588);
and U256 (N_256,In_13,In_1447);
or U257 (N_257,In_609,In_1449);
or U258 (N_258,In_1379,In_514);
and U259 (N_259,In_1747,In_1207);
nor U260 (N_260,In_792,In_1074);
xor U261 (N_261,In_515,In_1296);
nand U262 (N_262,In_156,In_1940);
nor U263 (N_263,In_722,In_1571);
or U264 (N_264,In_744,In_237);
and U265 (N_265,In_314,In_1857);
nor U266 (N_266,In_916,In_843);
and U267 (N_267,In_1700,In_912);
xor U268 (N_268,In_318,In_895);
or U269 (N_269,In_1510,In_1374);
nand U270 (N_270,In_846,In_1705);
or U271 (N_271,In_342,In_199);
and U272 (N_272,In_1063,In_1342);
and U273 (N_273,In_1675,In_696);
nand U274 (N_274,In_1202,In_620);
nand U275 (N_275,In_1289,In_1619);
xnor U276 (N_276,In_35,In_545);
nor U277 (N_277,In_281,In_1129);
and U278 (N_278,In_1031,In_416);
nor U279 (N_279,In_721,In_657);
or U280 (N_280,In_377,In_1983);
and U281 (N_281,In_1898,In_893);
and U282 (N_282,In_1298,In_840);
nand U283 (N_283,In_806,In_946);
nand U284 (N_284,In_172,In_1753);
and U285 (N_285,In_1263,In_1354);
or U286 (N_286,In_1352,In_1546);
and U287 (N_287,In_1204,In_560);
nor U288 (N_288,In_953,In_1456);
or U289 (N_289,In_60,In_1842);
or U290 (N_290,In_1028,In_1460);
and U291 (N_291,In_1817,In_1828);
or U292 (N_292,In_1137,In_1265);
nor U293 (N_293,In_774,In_58);
or U294 (N_294,In_1109,In_295);
xnor U295 (N_295,In_940,In_807);
or U296 (N_296,In_465,In_1223);
nor U297 (N_297,In_1886,In_1822);
or U298 (N_298,In_8,In_1531);
nand U299 (N_299,In_1884,In_170);
nand U300 (N_300,In_557,In_1873);
xor U301 (N_301,In_1730,In_144);
nor U302 (N_302,In_668,In_581);
nor U303 (N_303,In_1894,In_235);
and U304 (N_304,In_801,In_1285);
nor U305 (N_305,In_536,In_727);
or U306 (N_306,In_1475,In_444);
and U307 (N_307,In_116,In_1974);
or U308 (N_308,In_1396,In_569);
xnor U309 (N_309,In_407,In_1798);
nor U310 (N_310,In_1424,In_604);
nand U311 (N_311,In_503,In_1890);
nor U312 (N_312,In_986,In_1315);
xor U313 (N_313,In_1544,In_709);
or U314 (N_314,In_1122,In_1345);
or U315 (N_315,In_1859,In_408);
nand U316 (N_316,In_403,In_1160);
or U317 (N_317,In_688,In_1408);
and U318 (N_318,In_1320,In_361);
nor U319 (N_319,In_10,In_1934);
or U320 (N_320,In_1989,In_1532);
xnor U321 (N_321,In_1955,In_1665);
or U322 (N_322,In_186,In_908);
and U323 (N_323,In_1435,In_387);
or U324 (N_324,In_866,In_1277);
or U325 (N_325,In_1925,In_564);
nand U326 (N_326,In_950,In_541);
nor U327 (N_327,In_1371,In_1274);
nor U328 (N_328,In_1412,In_250);
nand U329 (N_329,In_1972,In_627);
or U330 (N_330,In_158,In_1870);
nand U331 (N_331,In_349,In_738);
and U332 (N_332,In_1613,In_1330);
nor U333 (N_333,In_1015,In_686);
or U334 (N_334,In_282,In_1208);
and U335 (N_335,In_398,In_271);
nor U336 (N_336,In_274,In_1182);
and U337 (N_337,In_814,In_615);
and U338 (N_338,In_1627,In_1605);
and U339 (N_339,In_926,In_400);
or U340 (N_340,In_1476,In_1479);
nor U341 (N_341,In_1901,In_1548);
and U342 (N_342,In_1542,In_1603);
nand U343 (N_343,In_1234,In_240);
nor U344 (N_344,In_1116,In_857);
and U345 (N_345,In_321,In_1721);
or U346 (N_346,In_1067,In_340);
nand U347 (N_347,In_1823,In_1419);
or U348 (N_348,In_1954,In_420);
xor U349 (N_349,In_951,In_219);
xnor U350 (N_350,In_837,In_1679);
and U351 (N_351,In_1852,In_1193);
and U352 (N_352,In_1729,In_344);
and U353 (N_353,In_1309,In_1750);
nor U354 (N_354,In_1696,In_1657);
or U355 (N_355,In_468,In_68);
and U356 (N_356,In_1939,In_1127);
or U357 (N_357,In_1323,In_1522);
nand U358 (N_358,In_1083,In_447);
nand U359 (N_359,In_1926,In_870);
and U360 (N_360,In_101,In_1734);
nand U361 (N_361,In_327,In_1459);
or U362 (N_362,In_148,In_1054);
nor U363 (N_363,In_1812,In_1237);
or U364 (N_364,In_396,In_1487);
nand U365 (N_365,In_117,In_85);
and U366 (N_366,In_871,In_602);
and U367 (N_367,In_772,In_683);
nor U368 (N_368,In_426,In_1682);
nor U369 (N_369,In_252,In_1557);
nor U370 (N_370,In_643,In_201);
nand U371 (N_371,In_948,In_966);
nor U372 (N_372,In_1195,In_1631);
nor U373 (N_373,In_701,In_1764);
and U374 (N_374,In_886,In_1348);
or U375 (N_375,In_923,In_1584);
nand U376 (N_376,In_65,In_1908);
xnor U377 (N_377,In_1306,In_332);
nand U378 (N_378,In_1278,In_474);
or U379 (N_379,In_341,In_795);
or U380 (N_380,In_1866,In_631);
and U381 (N_381,In_563,In_1818);
nand U382 (N_382,In_516,In_1610);
or U383 (N_383,In_519,In_207);
and U384 (N_384,In_1592,In_1530);
nand U385 (N_385,In_1716,In_1235);
or U386 (N_386,In_386,In_1225);
xor U387 (N_387,In_573,In_174);
nor U388 (N_388,In_909,In_1209);
or U389 (N_389,In_220,In_1024);
and U390 (N_390,In_763,In_1797);
nor U391 (N_391,In_626,In_238);
nand U392 (N_392,In_1091,In_1538);
nand U393 (N_393,In_1332,In_565);
and U394 (N_394,In_419,In_22);
or U395 (N_395,In_838,In_927);
and U396 (N_396,In_965,In_1733);
and U397 (N_397,In_1683,In_538);
xnor U398 (N_398,In_1071,In_1924);
or U399 (N_399,In_1712,In_1673);
and U400 (N_400,In_1806,In_1432);
and U401 (N_401,In_859,In_1240);
or U402 (N_402,In_1075,In_1991);
and U403 (N_403,In_1159,In_1440);
nor U404 (N_404,In_624,In_422);
nor U405 (N_405,In_1820,In_439);
and U406 (N_406,In_883,In_1008);
or U407 (N_407,In_257,In_410);
nor U408 (N_408,In_276,In_999);
or U409 (N_409,In_1055,In_1880);
nand U410 (N_410,In_734,In_1451);
xnor U411 (N_411,In_613,In_412);
nand U412 (N_412,In_441,In_1641);
nand U413 (N_413,In_1785,In_1196);
and U414 (N_414,In_336,In_1722);
nand U415 (N_415,In_331,In_1504);
and U416 (N_416,In_1555,In_932);
nand U417 (N_417,In_1710,In_1836);
nand U418 (N_418,In_599,In_1919);
nor U419 (N_419,In_1968,In_1858);
or U420 (N_420,In_1303,In_389);
nor U421 (N_421,In_1582,In_654);
or U422 (N_422,In_664,In_759);
xor U423 (N_423,In_1377,In_1452);
or U424 (N_424,In_694,In_1523);
xor U425 (N_425,In_1,In_1375);
or U426 (N_426,In_1783,In_446);
nor U427 (N_427,In_710,In_1790);
nor U428 (N_428,In_179,In_352);
nand U429 (N_429,In_165,In_955);
xor U430 (N_430,In_218,In_1119);
nor U431 (N_431,In_1321,In_1941);
or U432 (N_432,In_1529,In_1699);
and U433 (N_433,In_1577,In_554);
nor U434 (N_434,In_436,In_1397);
or U435 (N_435,In_1607,In_1453);
and U436 (N_436,In_1461,In_855);
and U437 (N_437,In_1187,In_127);
or U438 (N_438,In_348,In_1029);
and U439 (N_439,In_1387,In_962);
xor U440 (N_440,In_1492,In_1560);
and U441 (N_441,In_11,In_1242);
nand U442 (N_442,In_1394,In_793);
nand U443 (N_443,In_1226,In_214);
or U444 (N_444,In_212,In_1869);
and U445 (N_445,In_492,In_1161);
or U446 (N_446,In_894,In_365);
and U447 (N_447,In_1536,In_630);
nor U448 (N_448,In_691,In_230);
or U449 (N_449,In_1087,In_718);
nand U450 (N_450,In_388,In_821);
nand U451 (N_451,In_819,In_1800);
or U452 (N_452,In_1585,In_209);
nand U453 (N_453,In_1864,In_903);
and U454 (N_454,In_1142,In_1253);
nand U455 (N_455,In_171,In_1329);
xor U456 (N_456,In_1148,In_764);
or U457 (N_457,In_919,In_120);
xnor U458 (N_458,In_397,In_357);
or U459 (N_459,In_969,In_456);
xnor U460 (N_460,In_476,In_1259);
nor U461 (N_461,In_1478,In_1961);
and U462 (N_462,In_934,In_897);
nor U463 (N_463,In_1466,In_90);
and U464 (N_464,In_100,In_1136);
nand U465 (N_465,In_1092,In_551);
xor U466 (N_466,In_881,In_300);
or U467 (N_467,In_1628,In_1727);
or U468 (N_468,In_1777,In_1844);
and U469 (N_469,In_1328,In_1417);
nand U470 (N_470,In_1252,In_865);
xor U471 (N_471,In_1036,In_937);
and U472 (N_472,In_1086,In_970);
nor U473 (N_473,In_488,In_1561);
or U474 (N_474,In_509,In_479);
or U475 (N_475,In_1846,In_1297);
or U476 (N_476,In_26,In_540);
nor U477 (N_477,In_1763,In_1185);
xnor U478 (N_478,In_762,In_1003);
or U479 (N_479,In_1385,In_936);
nor U480 (N_480,In_982,In_1286);
xnor U481 (N_481,In_1711,In_1120);
nand U482 (N_482,In_576,In_356);
nand U483 (N_483,In_980,In_500);
and U484 (N_484,In_1406,In_616);
and U485 (N_485,In_1594,In_1636);
nand U486 (N_486,In_1903,In_914);
and U487 (N_487,In_346,In_1214);
nand U488 (N_488,In_704,In_1089);
or U489 (N_489,In_1654,In_1336);
or U490 (N_490,In_651,In_747);
and U491 (N_491,In_80,In_1355);
xor U492 (N_492,In_248,In_1113);
xor U493 (N_493,In_1065,In_175);
xnor U494 (N_494,In_1574,In_1445);
or U495 (N_495,In_973,In_303);
nand U496 (N_496,In_1855,In_102);
nand U497 (N_497,In_1567,In_223);
nor U498 (N_498,In_675,In_1179);
and U499 (N_499,In_635,In_288);
nand U500 (N_500,In_689,In_638);
nand U501 (N_501,In_1639,In_1656);
nor U502 (N_502,In_676,In_1779);
or U503 (N_503,In_1688,In_1905);
nand U504 (N_504,In_1291,In_1596);
or U505 (N_505,In_7,In_293);
or U506 (N_506,In_181,In_972);
or U507 (N_507,In_87,In_724);
and U508 (N_508,In_1519,In_669);
and U509 (N_509,In_106,In_1079);
nand U510 (N_510,In_824,In_1189);
and U511 (N_511,In_789,In_549);
nand U512 (N_512,In_1126,In_529);
nand U513 (N_513,In_1269,In_1125);
or U514 (N_514,In_648,In_1931);
xor U515 (N_515,In_719,In_442);
and U516 (N_516,In_489,In_362);
or U517 (N_517,In_113,In_918);
and U518 (N_518,In_530,In_720);
or U519 (N_519,In_1724,In_1426);
nor U520 (N_520,In_776,In_1341);
and U521 (N_521,In_1210,In_1244);
nand U522 (N_522,In_1474,In_1220);
or U523 (N_523,In_1176,In_1177);
nor U524 (N_524,In_42,In_1043);
nor U525 (N_525,In_25,In_1976);
nor U526 (N_526,In_89,In_457);
nand U527 (N_527,In_737,In_92);
and U528 (N_528,In_485,In_1376);
and U529 (N_529,In_1543,In_981);
nor U530 (N_530,In_921,In_16);
nor U531 (N_531,In_1816,In_1027);
and U532 (N_532,In_1701,In_674);
nand U533 (N_533,In_944,In_608);
and U534 (N_534,In_298,In_1581);
and U535 (N_535,In_123,In_681);
nor U536 (N_536,In_715,In_1524);
or U537 (N_537,In_848,In_533);
nand U538 (N_538,In_1634,In_1186);
or U539 (N_539,In_409,In_343);
nand U540 (N_540,In_1876,In_1980);
or U541 (N_541,In_1326,In_1112);
or U542 (N_542,In_345,In_1367);
or U543 (N_543,In_98,In_287);
and U544 (N_544,In_748,In_1200);
nor U545 (N_545,In_1788,In_280);
and U546 (N_546,In_984,In_834);
xor U547 (N_547,In_1425,In_478);
and U548 (N_548,In_1051,In_717);
nand U549 (N_549,In_1569,In_1735);
and U550 (N_550,In_1482,In_1620);
or U551 (N_551,In_1480,In_451);
nand U552 (N_552,In_319,In_1897);
nor U553 (N_553,In_431,In_328);
nand U554 (N_554,In_841,In_130);
nand U555 (N_555,In_1258,In_1191);
and U556 (N_556,In_1646,In_800);
and U557 (N_557,In_1334,In_1502);
or U558 (N_558,In_1623,In_1359);
xnor U559 (N_559,In_760,In_1264);
nor U560 (N_560,In_1416,In_324);
nand U561 (N_561,In_1752,In_1115);
and U562 (N_562,In_450,In_555);
nand U563 (N_563,In_1423,In_711);
nor U564 (N_564,In_382,In_1280);
or U565 (N_565,In_139,In_641);
nor U566 (N_566,In_1549,In_1708);
nor U567 (N_567,In_1163,In_211);
nor U568 (N_568,In_1640,In_1038);
and U569 (N_569,In_832,In_1012);
or U570 (N_570,In_71,In_699);
or U571 (N_571,In_716,In_1139);
and U572 (N_572,In_1420,In_73);
xnor U573 (N_573,In_2,In_653);
or U574 (N_574,In_1382,In_1663);
and U575 (N_575,In_825,In_1768);
nand U576 (N_576,In_1963,In_826);
xor U577 (N_577,In_162,In_126);
or U578 (N_578,In_6,In_524);
nand U579 (N_579,In_270,In_963);
or U580 (N_580,In_1618,In_335);
and U581 (N_581,In_1767,In_1256);
and U582 (N_582,In_0,In_1786);
nand U583 (N_583,In_469,In_5);
or U584 (N_584,In_706,In_376);
nor U585 (N_585,In_528,In_1140);
and U586 (N_586,In_1427,In_878);
nand U587 (N_587,In_1889,In_1227);
nor U588 (N_588,In_1503,In_1215);
nand U589 (N_589,In_1347,In_1018);
or U590 (N_590,In_775,In_1251);
or U591 (N_591,In_1740,In_1703);
and U592 (N_592,In_1390,In_935);
or U593 (N_593,In_1879,In_1784);
xor U594 (N_594,In_453,In_702);
nor U595 (N_595,In_1680,In_571);
nor U596 (N_596,In_473,In_1715);
and U597 (N_597,In_1659,In_1815);
nand U598 (N_598,In_1758,In_114);
nor U599 (N_599,In_226,In_621);
xor U600 (N_600,In_236,In_768);
nor U601 (N_601,In_729,In_196);
and U602 (N_602,In_1662,In_452);
or U603 (N_603,In_1049,In_1102);
or U604 (N_604,In_1509,In_1653);
and U605 (N_605,In_1756,In_1670);
nor U606 (N_606,In_329,In_1566);
nor U607 (N_607,In_291,In_979);
or U608 (N_608,In_844,In_286);
nor U609 (N_609,In_646,In_1106);
nor U610 (N_610,In_591,In_284);
and U611 (N_611,In_1472,In_234);
and U612 (N_612,In_1853,In_1372);
nand U613 (N_613,In_1174,In_227);
or U614 (N_614,In_1741,In_1739);
nor U615 (N_615,In_1276,In_1850);
nor U616 (N_616,In_256,In_1250);
nor U617 (N_617,In_1343,In_854);
nor U618 (N_618,In_1084,In_97);
nor U619 (N_619,In_48,In_1911);
or U620 (N_620,In_82,In_301);
and U621 (N_621,In_1590,In_368);
nor U622 (N_622,In_425,In_1082);
xor U623 (N_623,In_900,In_194);
and U624 (N_624,In_773,In_1266);
and U625 (N_625,In_1527,In_685);
xnor U626 (N_626,In_1044,In_1344);
or U627 (N_627,In_872,In_875);
and U628 (N_628,In_1231,In_1292);
nor U629 (N_629,In_917,In_978);
or U630 (N_630,In_1626,In_1778);
or U631 (N_631,In_1525,In_1178);
nand U632 (N_632,In_121,In_31);
nand U633 (N_633,In_251,In_1909);
nand U634 (N_634,In_359,In_306);
or U635 (N_635,In_1878,In_827);
nor U636 (N_636,In_1514,In_1072);
nor U637 (N_637,In_1034,In_1248);
nor U638 (N_638,In_1835,In_15);
nand U639 (N_639,In_1360,In_166);
nor U640 (N_640,In_315,In_891);
nor U641 (N_641,In_299,In_1649);
xnor U642 (N_642,In_486,In_896);
xor U643 (N_643,In_892,In_355);
nor U644 (N_644,In_1128,In_1020);
and U645 (N_645,In_833,In_1655);
nor U646 (N_646,In_371,In_1030);
nand U647 (N_647,In_588,In_582);
and U648 (N_648,In_44,In_1141);
nand U649 (N_649,In_1066,In_1493);
nand U650 (N_650,In_107,In_901);
nor U651 (N_651,In_475,In_1912);
nand U652 (N_652,In_1962,In_996);
or U653 (N_653,In_1099,In_1260);
or U654 (N_654,In_55,In_1684);
or U655 (N_655,In_1944,In_911);
xnor U656 (N_656,In_381,In_1154);
nor U657 (N_657,In_1351,In_1923);
or U658 (N_658,In_1554,In_518);
and U659 (N_659,In_584,In_1922);
nor U660 (N_660,In_1937,In_949);
nand U661 (N_661,In_1678,In_1984);
or U662 (N_662,In_1792,In_1484);
or U663 (N_663,In_867,In_1033);
xor U664 (N_664,In_122,In_1563);
and U665 (N_665,In_445,In_1644);
or U666 (N_666,In_662,In_713);
or U667 (N_667,In_1415,In_217);
nand U668 (N_668,In_752,In_56);
xor U669 (N_669,In_1001,In_527);
nor U670 (N_670,In_4,In_405);
and U671 (N_671,In_285,In_1637);
or U672 (N_672,In_749,In_1893);
or U673 (N_673,In_164,In_1095);
nor U674 (N_674,In_1045,In_210);
nand U675 (N_675,In_1945,In_593);
nor U676 (N_676,In_663,In_1181);
and U677 (N_677,In_70,In_1199);
and U678 (N_678,In_544,In_279);
nand U679 (N_679,In_1885,In_133);
or U680 (N_680,In_678,In_367);
and U681 (N_681,In_1322,In_1167);
nor U682 (N_682,In_1041,In_1907);
and U683 (N_683,In_777,In_1275);
or U684 (N_684,In_103,In_682);
nor U685 (N_685,In_1236,In_167);
nand U686 (N_686,In_743,In_1892);
and U687 (N_687,In_1070,In_808);
nand U688 (N_688,In_1601,In_1927);
nand U689 (N_689,In_751,In_399);
nor U690 (N_690,In_1796,In_1650);
nor U691 (N_691,In_1488,In_435);
nor U692 (N_692,In_1803,In_296);
or U693 (N_693,In_1216,In_482);
nand U694 (N_694,In_46,In_129);
and U695 (N_695,In_1913,In_1299);
and U696 (N_696,In_232,In_1793);
xor U697 (N_697,In_1608,In_449);
nand U698 (N_698,In_994,In_1953);
nand U699 (N_699,In_1867,In_1985);
xor U700 (N_700,In_28,In_401);
and U701 (N_701,In_1789,In_1770);
or U702 (N_702,In_1458,In_1023);
nor U703 (N_703,In_334,In_957);
or U704 (N_704,In_1448,In_477);
xor U705 (N_705,In_200,In_690);
nand U706 (N_706,In_402,In_598);
nor U707 (N_707,In_37,In_1831);
xnor U708 (N_708,In_559,In_1040);
xor U709 (N_709,In_1138,In_733);
nand U710 (N_710,In_1473,In_1947);
or U711 (N_711,In_1254,In_1552);
and U712 (N_712,In_40,In_1222);
nor U713 (N_713,In_1959,In_809);
and U714 (N_714,In_1241,In_1979);
and U715 (N_715,In_124,In_1609);
xnor U716 (N_716,In_1583,In_424);
xor U717 (N_717,In_756,In_823);
and U718 (N_718,In_1616,In_633);
xor U719 (N_719,In_150,In_938);
xnor U720 (N_720,In_766,In_1591);
nand U721 (N_721,In_1025,In_977);
or U722 (N_722,In_1052,In_1877);
nor U723 (N_723,In_864,In_1942);
xnor U724 (N_724,In_645,In_1689);
xnor U725 (N_725,In_147,In_1717);
nor U726 (N_726,In_1827,In_1145);
and U727 (N_727,In_1813,In_1998);
and U728 (N_728,In_1246,In_1916);
nand U729 (N_729,In_1606,In_390);
nor U730 (N_730,In_1462,In_94);
or U731 (N_731,In_1746,In_1175);
and U732 (N_732,In_249,In_1541);
or U733 (N_733,In_141,In_125);
nor U734 (N_734,In_57,In_672);
xor U735 (N_735,In_1505,In_665);
nand U736 (N_736,In_216,In_985);
and U737 (N_737,In_23,In_434);
nor U738 (N_738,In_1965,In_1930);
and U739 (N_739,In_36,In_1848);
and U740 (N_740,In_375,In_50);
xor U741 (N_741,In_330,In_929);
xnor U742 (N_742,In_392,In_849);
nor U743 (N_743,In_989,In_640);
nor U744 (N_744,In_1350,In_1149);
or U745 (N_745,In_429,In_1932);
nand U746 (N_746,In_742,In_754);
nand U747 (N_747,In_1293,In_1671);
or U748 (N_748,In_1100,In_1132);
nor U749 (N_749,In_1381,In_797);
or U750 (N_750,In_976,In_337);
nor U751 (N_751,In_203,In_176);
and U752 (N_752,In_1632,In_813);
or U753 (N_753,In_523,In_1600);
nor U754 (N_754,In_1437,In_1599);
nand U755 (N_755,In_1305,In_1431);
and U756 (N_756,In_661,In_862);
nor U757 (N_757,In_228,In_583);
nand U758 (N_758,In_1651,In_1713);
nand U759 (N_759,In_1165,In_1765);
or U760 (N_760,In_265,In_1805);
nand U761 (N_761,In_820,In_922);
xor U762 (N_762,In_510,In_1791);
nand U763 (N_763,In_1284,In_1950);
xor U764 (N_764,In_1981,In_1780);
and U765 (N_765,In_1794,In_1719);
nand U766 (N_766,In_1745,In_1617);
xnor U767 (N_767,In_406,In_404);
nand U768 (N_768,In_438,In_794);
nor U769 (N_769,In_32,In_1224);
or U770 (N_770,In_817,In_1539);
and U771 (N_771,In_876,In_782);
xnor U772 (N_772,In_1311,In_786);
nor U773 (N_773,In_3,In_197);
nand U774 (N_774,In_1206,In_1775);
nand U775 (N_775,In_1995,In_1057);
nor U776 (N_776,In_1992,In_1910);
nand U777 (N_777,In_480,In_1849);
or U778 (N_778,In_411,In_726);
xnor U779 (N_779,In_632,In_1114);
nor U780 (N_780,In_1361,In_326);
or U781 (N_781,In_1587,In_1485);
and U782 (N_782,In_491,In_69);
nand U783 (N_783,In_548,In_440);
nand U784 (N_784,In_815,In_1249);
nor U785 (N_785,In_1369,In_993);
nand U786 (N_786,In_1255,In_21);
or U787 (N_787,In_1032,In_1624);
nor U788 (N_788,In_1611,In_1414);
and U789 (N_789,In_213,In_1068);
and U790 (N_790,In_1391,In_1353);
nor U791 (N_791,In_267,In_623);
nor U792 (N_792,In_1677,In_812);
nand U793 (N_793,In_589,In_1882);
nand U794 (N_794,In_1760,In_1928);
and U795 (N_795,In_1477,In_1221);
or U796 (N_796,In_1471,In_636);
or U797 (N_797,In_1824,In_899);
nor U798 (N_798,In_1418,In_995);
nand U799 (N_799,In_1450,In_845);
or U800 (N_800,In_1026,In_700);
and U801 (N_801,In_1902,In_649);
and U802 (N_802,In_1171,In_1732);
or U803 (N_803,In_522,In_380);
nand U804 (N_804,In_1370,In_804);
or U805 (N_805,In_1380,In_430);
nand U806 (N_806,In_755,In_63);
or U807 (N_807,In_313,In_964);
or U808 (N_808,In_1002,In_990);
and U809 (N_809,In_1498,In_767);
nand U810 (N_810,In_913,In_836);
or U811 (N_811,In_959,In_1402);
nand U812 (N_812,In_119,In_693);
or U813 (N_813,In_1398,In_1997);
nor U814 (N_814,In_1150,In_542);
nand U815 (N_815,In_1612,In_163);
and U816 (N_816,In_1046,In_1744);
nor U817 (N_817,In_697,In_24);
nand U818 (N_818,In_128,In_505);
and U819 (N_819,In_1162,In_487);
or U820 (N_820,In_732,In_1413);
or U821 (N_821,In_618,In_1802);
and U822 (N_822,In_224,In_723);
and U823 (N_823,In_364,In_525);
nor U824 (N_824,In_1281,In_1578);
and U825 (N_825,In_906,In_1211);
and U826 (N_826,In_830,In_579);
nor U827 (N_827,In_350,In_1666);
nand U828 (N_828,In_1118,In_679);
and U829 (N_829,In_433,In_1642);
or U830 (N_830,In_595,In_1814);
or U831 (N_831,In_941,In_1295);
or U832 (N_832,In_692,In_974);
nor U833 (N_833,In_30,In_998);
nor U834 (N_834,In_1565,In_309);
and U835 (N_835,In_255,In_513);
nor U836 (N_836,In_708,In_1061);
nor U837 (N_837,In_785,In_1184);
or U838 (N_838,In_154,In_1198);
nand U839 (N_839,In_483,In_1156);
nor U840 (N_840,In_1283,In_575);
nand U841 (N_841,In_1860,In_1465);
nor U842 (N_842,In_780,In_320);
or U843 (N_843,In_1973,In_521);
and U844 (N_844,In_1368,In_222);
nor U845 (N_845,In_1550,In_17);
nand U846 (N_846,In_305,In_570);
or U847 (N_847,In_707,In_1899);
nand U848 (N_848,In_1685,In_784);
or U849 (N_849,In_1556,In_1314);
and U850 (N_850,In_1868,In_988);
or U851 (N_851,In_1862,In_740);
and U852 (N_852,In_1301,In_1668);
and U853 (N_853,In_874,In_1469);
and U854 (N_854,In_1595,In_1383);
nand U855 (N_855,In_414,In_428);
and U856 (N_856,In_1863,In_1421);
and U857 (N_857,In_1401,In_1088);
nand U858 (N_858,In_1438,In_1267);
nor U859 (N_859,In_504,In_169);
nor U860 (N_860,In_1164,In_1058);
nor U861 (N_861,In_1725,In_1891);
xnor U862 (N_862,In_137,In_498);
nand U863 (N_863,In_712,In_1900);
or U864 (N_864,In_975,In_511);
nor U865 (N_865,In_952,In_1060);
nand U866 (N_866,In_1674,In_1676);
or U867 (N_867,In_391,In_574);
xnor U868 (N_868,In_1319,In_18);
nand U869 (N_869,In_1967,In_155);
or U870 (N_870,In_847,In_1604);
nor U871 (N_871,In_552,In_27);
nor U872 (N_872,In_779,In_1238);
or U873 (N_873,In_1183,In_484);
nand U874 (N_874,In_1410,In_289);
and U875 (N_875,In_512,In_634);
and U876 (N_876,In_1457,In_1960);
nand U877 (N_877,In_373,In_423);
and U878 (N_878,In_1168,In_556);
and U879 (N_879,In_920,In_658);
xor U880 (N_880,In_1294,In_1170);
nand U881 (N_881,In_1553,In_739);
nand U882 (N_882,In_1977,In_244);
nand U883 (N_883,In_1105,In_816);
nor U884 (N_884,In_1076,In_243);
xor U885 (N_885,In_78,In_1731);
nor U886 (N_886,In_417,In_803);
nor U887 (N_887,In_283,In_358);
or U888 (N_888,In_360,In_245);
nand U889 (N_889,In_1357,In_1830);
nand U890 (N_890,In_1881,In_52);
or U891 (N_891,In_1570,In_670);
nor U892 (N_892,In_1491,In_198);
and U893 (N_893,In_1107,In_1810);
or U894 (N_894,In_1748,In_1019);
and U895 (N_895,In_1404,In_600);
nor U896 (N_896,In_798,In_1446);
and U897 (N_897,In_464,In_1430);
xnor U898 (N_898,In_1434,In_1094);
nor U899 (N_899,In_499,In_1338);
xor U900 (N_900,In_550,In_1988);
nor U901 (N_901,In_1568,In_41);
nand U902 (N_902,In_1888,In_463);
or U903 (N_903,In_33,In_1687);
and U904 (N_904,In_1622,In_507);
nor U905 (N_905,In_1117,In_497);
nor U906 (N_906,In_1205,In_1686);
nand U907 (N_907,In_1339,In_1795);
nand U908 (N_908,In_705,In_427);
nand U909 (N_909,In_787,In_877);
and U910 (N_910,In_1929,In_51);
nand U911 (N_911,In_757,In_1239);
xnor U912 (N_912,In_1615,In_1990);
nor U913 (N_913,In_88,In_1317);
and U914 (N_914,In_1153,In_1152);
nor U915 (N_915,In_75,In_1229);
and U916 (N_916,In_19,In_1660);
xnor U917 (N_917,In_77,In_1340);
nor U918 (N_918,In_1454,In_1017);
nand U919 (N_919,In_1669,In_553);
or U920 (N_920,In_1933,In_578);
nand U921 (N_921,In_695,In_1540);
nor U922 (N_922,In_539,In_943);
nand U923 (N_923,In_907,In_1841);
nor U924 (N_924,In_1874,In_501);
or U925 (N_925,In_1658,In_1728);
nor U926 (N_926,In_1016,In_1652);
and U927 (N_927,In_1373,In_1526);
or U928 (N_928,In_1366,In_769);
and U929 (N_929,In_142,In_1098);
xor U930 (N_930,In_143,In_968);
nor U931 (N_931,In_1144,In_617);
or U932 (N_932,In_1956,In_1714);
or U933 (N_933,In_1166,In_233);
nand U934 (N_934,In_79,In_1572);
nor U935 (N_935,In_1643,In_585);
or U936 (N_936,In_1738,In_183);
nor U937 (N_937,In_606,In_1704);
nand U938 (N_938,In_136,In_1464);
nor U939 (N_939,In_765,In_1429);
or U940 (N_940,In_1110,In_496);
nand U941 (N_941,In_603,In_45);
nand U942 (N_942,In_629,In_1130);
nand U943 (N_943,In_322,In_1501);
nand U944 (N_944,In_140,In_1854);
and U945 (N_945,In_802,In_1914);
nor U946 (N_946,In_619,In_790);
nand U947 (N_947,In_495,In_1506);
nor U948 (N_948,In_882,In_835);
or U949 (N_949,In_1573,In_1428);
xnor U950 (N_950,In_956,In_1077);
nor U951 (N_951,In_1861,In_1564);
nor U952 (N_952,In_1887,In_1782);
nor U953 (N_953,In_1436,In_725);
and U954 (N_954,In_853,In_1771);
and U955 (N_955,In_455,In_822);
and U956 (N_956,In_1324,In_379);
and U957 (N_957,In_967,In_1386);
nor U958 (N_958,In_884,In_1558);
nor U959 (N_959,In_159,In_258);
and U960 (N_960,In_266,In_639);
or U961 (N_961,In_310,In_1047);
and U962 (N_962,In_928,In_135);
nor U963 (N_963,In_1190,In_372);
nor U964 (N_964,In_1124,In_868);
or U965 (N_965,In_67,In_1702);
and U966 (N_966,In_987,In_1232);
xnor U967 (N_967,In_1856,In_1056);
and U968 (N_968,In_1010,In_905);
and U969 (N_969,In_671,In_890);
or U970 (N_970,In_1271,In_1104);
or U971 (N_971,In_153,In_741);
and U972 (N_972,In_1483,In_1845);
and U973 (N_973,In_459,In_873);
or U974 (N_974,In_62,In_269);
and U975 (N_975,In_93,In_311);
and U976 (N_976,In_1346,In_1993);
nor U977 (N_977,In_448,In_1826);
nand U978 (N_978,In_1754,In_1304);
nor U979 (N_979,In_728,In_1987);
nand U980 (N_980,In_180,In_1048);
nor U981 (N_981,In_1180,In_587);
or U982 (N_982,In_1559,In_1938);
nor U983 (N_983,In_799,In_811);
or U984 (N_984,In_1157,In_861);
or U985 (N_985,In_568,In_302);
or U986 (N_986,In_472,In_1978);
or U987 (N_987,In_1547,In_208);
nand U988 (N_988,In_1349,In_954);
xor U989 (N_989,In_110,In_1575);
or U990 (N_990,In_771,In_746);
nor U991 (N_991,In_54,In_74);
xnor U992 (N_992,In_264,In_660);
nand U993 (N_993,In_612,In_939);
nor U994 (N_994,In_1508,In_1363);
xor U995 (N_995,In_1004,In_655);
or U996 (N_996,In_1405,In_1039);
or U997 (N_997,In_1533,In_1037);
and U998 (N_998,In_1718,In_109);
nor U999 (N_999,In_647,In_1422);
or U1000 (N_1000,In_1839,In_1101);
and U1001 (N_1001,In_455,In_1524);
or U1002 (N_1002,In_147,In_414);
or U1003 (N_1003,In_1900,In_1068);
xor U1004 (N_1004,In_1336,In_1080);
nand U1005 (N_1005,In_185,In_43);
nor U1006 (N_1006,In_97,In_249);
nor U1007 (N_1007,In_1762,In_462);
and U1008 (N_1008,In_1549,In_451);
xnor U1009 (N_1009,In_827,In_870);
xor U1010 (N_1010,In_1238,In_326);
nand U1011 (N_1011,In_447,In_467);
nor U1012 (N_1012,In_284,In_143);
and U1013 (N_1013,In_1968,In_381);
or U1014 (N_1014,In_1436,In_1960);
and U1015 (N_1015,In_1320,In_1282);
nand U1016 (N_1016,In_1185,In_680);
nor U1017 (N_1017,In_1035,In_1099);
nor U1018 (N_1018,In_1270,In_1676);
xnor U1019 (N_1019,In_1284,In_611);
nand U1020 (N_1020,In_570,In_1978);
nand U1021 (N_1021,In_261,In_1569);
nor U1022 (N_1022,In_520,In_487);
nor U1023 (N_1023,In_1339,In_1499);
or U1024 (N_1024,In_853,In_1150);
nand U1025 (N_1025,In_518,In_1855);
nor U1026 (N_1026,In_1110,In_1797);
nor U1027 (N_1027,In_1725,In_973);
and U1028 (N_1028,In_979,In_894);
nor U1029 (N_1029,In_862,In_33);
nor U1030 (N_1030,In_144,In_70);
xnor U1031 (N_1031,In_241,In_894);
nor U1032 (N_1032,In_1850,In_985);
nor U1033 (N_1033,In_1726,In_344);
nor U1034 (N_1034,In_1645,In_1582);
nor U1035 (N_1035,In_574,In_1077);
or U1036 (N_1036,In_378,In_282);
nor U1037 (N_1037,In_775,In_509);
xnor U1038 (N_1038,In_759,In_1591);
or U1039 (N_1039,In_679,In_1899);
nor U1040 (N_1040,In_1441,In_1682);
and U1041 (N_1041,In_1748,In_600);
nor U1042 (N_1042,In_1023,In_409);
or U1043 (N_1043,In_514,In_43);
or U1044 (N_1044,In_27,In_1501);
and U1045 (N_1045,In_323,In_98);
or U1046 (N_1046,In_1799,In_470);
or U1047 (N_1047,In_1285,In_1736);
xor U1048 (N_1048,In_1327,In_1658);
and U1049 (N_1049,In_1712,In_704);
or U1050 (N_1050,In_1766,In_533);
xor U1051 (N_1051,In_1183,In_990);
nor U1052 (N_1052,In_712,In_700);
xnor U1053 (N_1053,In_1197,In_765);
nand U1054 (N_1054,In_1191,In_115);
or U1055 (N_1055,In_114,In_1517);
or U1056 (N_1056,In_1579,In_1567);
or U1057 (N_1057,In_116,In_1157);
or U1058 (N_1058,In_1333,In_1599);
xnor U1059 (N_1059,In_1554,In_1014);
nor U1060 (N_1060,In_229,In_687);
nand U1061 (N_1061,In_395,In_317);
nor U1062 (N_1062,In_535,In_541);
nor U1063 (N_1063,In_219,In_690);
and U1064 (N_1064,In_1869,In_1547);
nor U1065 (N_1065,In_260,In_908);
nand U1066 (N_1066,In_730,In_1351);
or U1067 (N_1067,In_1013,In_199);
or U1068 (N_1068,In_958,In_1999);
nor U1069 (N_1069,In_87,In_918);
nor U1070 (N_1070,In_662,In_389);
nand U1071 (N_1071,In_1425,In_45);
nor U1072 (N_1072,In_532,In_15);
nor U1073 (N_1073,In_552,In_578);
and U1074 (N_1074,In_1095,In_445);
nand U1075 (N_1075,In_1057,In_746);
nor U1076 (N_1076,In_910,In_1850);
nor U1077 (N_1077,In_1473,In_183);
and U1078 (N_1078,In_1338,In_1407);
or U1079 (N_1079,In_616,In_534);
and U1080 (N_1080,In_1116,In_1005);
nand U1081 (N_1081,In_396,In_139);
or U1082 (N_1082,In_1345,In_412);
xor U1083 (N_1083,In_282,In_1495);
or U1084 (N_1084,In_893,In_256);
or U1085 (N_1085,In_1678,In_540);
or U1086 (N_1086,In_62,In_1640);
or U1087 (N_1087,In_563,In_1212);
or U1088 (N_1088,In_181,In_1811);
or U1089 (N_1089,In_1500,In_288);
or U1090 (N_1090,In_1779,In_1266);
or U1091 (N_1091,In_43,In_1);
and U1092 (N_1092,In_124,In_1024);
or U1093 (N_1093,In_1817,In_319);
nor U1094 (N_1094,In_1723,In_23);
nand U1095 (N_1095,In_1329,In_920);
nand U1096 (N_1096,In_1659,In_448);
and U1097 (N_1097,In_683,In_1989);
nand U1098 (N_1098,In_867,In_745);
nor U1099 (N_1099,In_133,In_1877);
and U1100 (N_1100,In_411,In_730);
or U1101 (N_1101,In_1152,In_183);
nor U1102 (N_1102,In_1223,In_185);
or U1103 (N_1103,In_872,In_1121);
nand U1104 (N_1104,In_186,In_1772);
and U1105 (N_1105,In_1113,In_1634);
or U1106 (N_1106,In_44,In_1693);
nand U1107 (N_1107,In_1658,In_177);
and U1108 (N_1108,In_601,In_1493);
nor U1109 (N_1109,In_1182,In_1628);
nor U1110 (N_1110,In_108,In_75);
nor U1111 (N_1111,In_243,In_251);
xor U1112 (N_1112,In_17,In_1392);
and U1113 (N_1113,In_747,In_1432);
nor U1114 (N_1114,In_519,In_1453);
xnor U1115 (N_1115,In_1225,In_1818);
nand U1116 (N_1116,In_131,In_493);
nand U1117 (N_1117,In_1143,In_339);
nand U1118 (N_1118,In_1502,In_1745);
nor U1119 (N_1119,In_648,In_1224);
nor U1120 (N_1120,In_282,In_206);
or U1121 (N_1121,In_1500,In_498);
or U1122 (N_1122,In_678,In_810);
or U1123 (N_1123,In_563,In_510);
or U1124 (N_1124,In_1755,In_998);
nor U1125 (N_1125,In_847,In_334);
and U1126 (N_1126,In_210,In_1379);
and U1127 (N_1127,In_477,In_1970);
and U1128 (N_1128,In_1669,In_260);
nand U1129 (N_1129,In_1499,In_425);
xor U1130 (N_1130,In_392,In_1585);
and U1131 (N_1131,In_1345,In_799);
nand U1132 (N_1132,In_1151,In_675);
nand U1133 (N_1133,In_1268,In_1357);
or U1134 (N_1134,In_1596,In_382);
xnor U1135 (N_1135,In_1007,In_901);
nor U1136 (N_1136,In_1373,In_1940);
or U1137 (N_1137,In_526,In_283);
xor U1138 (N_1138,In_1054,In_1413);
and U1139 (N_1139,In_121,In_296);
nor U1140 (N_1140,In_154,In_146);
and U1141 (N_1141,In_814,In_1493);
and U1142 (N_1142,In_1764,In_1994);
and U1143 (N_1143,In_1178,In_1);
xnor U1144 (N_1144,In_377,In_678);
nand U1145 (N_1145,In_1431,In_124);
and U1146 (N_1146,In_148,In_28);
and U1147 (N_1147,In_1145,In_424);
nand U1148 (N_1148,In_709,In_1776);
and U1149 (N_1149,In_1428,In_0);
and U1150 (N_1150,In_921,In_1682);
and U1151 (N_1151,In_535,In_573);
nor U1152 (N_1152,In_788,In_1319);
or U1153 (N_1153,In_1272,In_263);
or U1154 (N_1154,In_726,In_872);
and U1155 (N_1155,In_1453,In_367);
nor U1156 (N_1156,In_999,In_1420);
nor U1157 (N_1157,In_1839,In_1757);
or U1158 (N_1158,In_418,In_1131);
nor U1159 (N_1159,In_1593,In_1562);
and U1160 (N_1160,In_291,In_1953);
xnor U1161 (N_1161,In_361,In_578);
xnor U1162 (N_1162,In_779,In_651);
nor U1163 (N_1163,In_1523,In_1618);
xnor U1164 (N_1164,In_754,In_1191);
or U1165 (N_1165,In_1225,In_1578);
nor U1166 (N_1166,In_1311,In_1084);
nand U1167 (N_1167,In_1502,In_514);
or U1168 (N_1168,In_806,In_941);
nand U1169 (N_1169,In_1133,In_351);
nor U1170 (N_1170,In_191,In_1912);
xor U1171 (N_1171,In_1001,In_682);
nand U1172 (N_1172,In_1486,In_0);
or U1173 (N_1173,In_1858,In_270);
nor U1174 (N_1174,In_995,In_966);
or U1175 (N_1175,In_1953,In_927);
or U1176 (N_1176,In_924,In_450);
nor U1177 (N_1177,In_1789,In_1583);
and U1178 (N_1178,In_1915,In_983);
nand U1179 (N_1179,In_1128,In_736);
or U1180 (N_1180,In_1175,In_930);
and U1181 (N_1181,In_1392,In_518);
xnor U1182 (N_1182,In_1812,In_574);
nor U1183 (N_1183,In_1373,In_1641);
nor U1184 (N_1184,In_836,In_1557);
nor U1185 (N_1185,In_216,In_1474);
nor U1186 (N_1186,In_1427,In_1747);
nor U1187 (N_1187,In_1189,In_339);
nor U1188 (N_1188,In_729,In_139);
or U1189 (N_1189,In_1741,In_108);
nor U1190 (N_1190,In_1339,In_513);
and U1191 (N_1191,In_1483,In_1610);
xor U1192 (N_1192,In_716,In_94);
nor U1193 (N_1193,In_490,In_445);
or U1194 (N_1194,In_1997,In_28);
and U1195 (N_1195,In_1457,In_1886);
xnor U1196 (N_1196,In_1027,In_647);
xnor U1197 (N_1197,In_148,In_1285);
nand U1198 (N_1198,In_580,In_1573);
nand U1199 (N_1199,In_848,In_128);
nor U1200 (N_1200,In_980,In_412);
or U1201 (N_1201,In_458,In_1629);
and U1202 (N_1202,In_550,In_117);
and U1203 (N_1203,In_950,In_1018);
xor U1204 (N_1204,In_543,In_1072);
nor U1205 (N_1205,In_1933,In_1376);
or U1206 (N_1206,In_31,In_650);
nor U1207 (N_1207,In_1905,In_1662);
nand U1208 (N_1208,In_499,In_1789);
xnor U1209 (N_1209,In_1028,In_908);
nand U1210 (N_1210,In_436,In_1707);
nand U1211 (N_1211,In_1605,In_1586);
and U1212 (N_1212,In_1236,In_1775);
and U1213 (N_1213,In_1491,In_1303);
and U1214 (N_1214,In_1507,In_703);
nand U1215 (N_1215,In_201,In_528);
nand U1216 (N_1216,In_378,In_1878);
nand U1217 (N_1217,In_65,In_1135);
nor U1218 (N_1218,In_1265,In_1097);
and U1219 (N_1219,In_1484,In_622);
nor U1220 (N_1220,In_601,In_1940);
nand U1221 (N_1221,In_717,In_237);
nand U1222 (N_1222,In_867,In_330);
and U1223 (N_1223,In_1215,In_932);
or U1224 (N_1224,In_1836,In_1738);
nand U1225 (N_1225,In_95,In_963);
xnor U1226 (N_1226,In_1992,In_1638);
and U1227 (N_1227,In_1074,In_1015);
nor U1228 (N_1228,In_483,In_369);
nand U1229 (N_1229,In_720,In_1453);
xor U1230 (N_1230,In_98,In_1401);
nand U1231 (N_1231,In_1805,In_1675);
nand U1232 (N_1232,In_1949,In_1061);
nor U1233 (N_1233,In_1488,In_798);
nand U1234 (N_1234,In_1860,In_1742);
nand U1235 (N_1235,In_436,In_1855);
nand U1236 (N_1236,In_1475,In_929);
nor U1237 (N_1237,In_1906,In_1667);
nor U1238 (N_1238,In_953,In_553);
and U1239 (N_1239,In_1225,In_144);
nand U1240 (N_1240,In_416,In_819);
xnor U1241 (N_1241,In_1954,In_444);
nand U1242 (N_1242,In_12,In_356);
and U1243 (N_1243,In_1012,In_871);
nand U1244 (N_1244,In_261,In_1128);
or U1245 (N_1245,In_214,In_1277);
nor U1246 (N_1246,In_1019,In_1357);
nor U1247 (N_1247,In_563,In_695);
nand U1248 (N_1248,In_338,In_1879);
and U1249 (N_1249,In_444,In_1483);
nand U1250 (N_1250,In_92,In_1731);
or U1251 (N_1251,In_137,In_1881);
or U1252 (N_1252,In_1139,In_264);
or U1253 (N_1253,In_968,In_505);
and U1254 (N_1254,In_1922,In_1218);
nor U1255 (N_1255,In_403,In_1766);
and U1256 (N_1256,In_1456,In_969);
and U1257 (N_1257,In_896,In_720);
or U1258 (N_1258,In_1318,In_583);
nor U1259 (N_1259,In_509,In_309);
nand U1260 (N_1260,In_1036,In_1659);
and U1261 (N_1261,In_1964,In_537);
nand U1262 (N_1262,In_1162,In_29);
and U1263 (N_1263,In_673,In_1049);
nor U1264 (N_1264,In_1296,In_1485);
nand U1265 (N_1265,In_1568,In_502);
nand U1266 (N_1266,In_1041,In_1774);
nor U1267 (N_1267,In_1311,In_687);
or U1268 (N_1268,In_610,In_343);
or U1269 (N_1269,In_303,In_1039);
or U1270 (N_1270,In_1390,In_1331);
or U1271 (N_1271,In_1338,In_1206);
xor U1272 (N_1272,In_1393,In_1337);
nand U1273 (N_1273,In_367,In_1958);
nor U1274 (N_1274,In_758,In_1114);
nor U1275 (N_1275,In_1900,In_1524);
or U1276 (N_1276,In_242,In_1484);
or U1277 (N_1277,In_1930,In_163);
and U1278 (N_1278,In_662,In_1665);
or U1279 (N_1279,In_1745,In_341);
or U1280 (N_1280,In_784,In_832);
xnor U1281 (N_1281,In_1705,In_214);
and U1282 (N_1282,In_684,In_1831);
nor U1283 (N_1283,In_734,In_384);
nand U1284 (N_1284,In_1278,In_1108);
or U1285 (N_1285,In_1455,In_418);
and U1286 (N_1286,In_618,In_1028);
or U1287 (N_1287,In_1873,In_772);
nand U1288 (N_1288,In_1993,In_1495);
nor U1289 (N_1289,In_564,In_681);
and U1290 (N_1290,In_1717,In_235);
nand U1291 (N_1291,In_973,In_1700);
nor U1292 (N_1292,In_168,In_1228);
xor U1293 (N_1293,In_1634,In_1630);
nor U1294 (N_1294,In_191,In_1118);
and U1295 (N_1295,In_623,In_528);
or U1296 (N_1296,In_1622,In_432);
or U1297 (N_1297,In_1159,In_77);
or U1298 (N_1298,In_1682,In_268);
nor U1299 (N_1299,In_89,In_1018);
nand U1300 (N_1300,In_662,In_1125);
nand U1301 (N_1301,In_374,In_1488);
nand U1302 (N_1302,In_218,In_67);
and U1303 (N_1303,In_847,In_576);
and U1304 (N_1304,In_1110,In_1855);
and U1305 (N_1305,In_1997,In_550);
and U1306 (N_1306,In_1298,In_765);
nor U1307 (N_1307,In_1982,In_1864);
nand U1308 (N_1308,In_519,In_235);
and U1309 (N_1309,In_1410,In_249);
nor U1310 (N_1310,In_1875,In_1086);
nand U1311 (N_1311,In_1765,In_1648);
nand U1312 (N_1312,In_616,In_984);
and U1313 (N_1313,In_1011,In_1150);
or U1314 (N_1314,In_737,In_829);
nand U1315 (N_1315,In_1938,In_1993);
and U1316 (N_1316,In_976,In_64);
or U1317 (N_1317,In_512,In_1647);
or U1318 (N_1318,In_876,In_1804);
nand U1319 (N_1319,In_897,In_26);
nor U1320 (N_1320,In_1006,In_1042);
or U1321 (N_1321,In_463,In_771);
xor U1322 (N_1322,In_672,In_347);
or U1323 (N_1323,In_1221,In_1538);
or U1324 (N_1324,In_25,In_997);
nand U1325 (N_1325,In_720,In_60);
nand U1326 (N_1326,In_1670,In_918);
xor U1327 (N_1327,In_1568,In_636);
nand U1328 (N_1328,In_1048,In_502);
or U1329 (N_1329,In_523,In_1589);
or U1330 (N_1330,In_1911,In_1399);
or U1331 (N_1331,In_318,In_956);
or U1332 (N_1332,In_27,In_1911);
nor U1333 (N_1333,In_785,In_591);
nor U1334 (N_1334,In_262,In_1122);
or U1335 (N_1335,In_1040,In_92);
nand U1336 (N_1336,In_226,In_373);
nand U1337 (N_1337,In_339,In_1293);
and U1338 (N_1338,In_1607,In_879);
nand U1339 (N_1339,In_443,In_751);
and U1340 (N_1340,In_832,In_1210);
nor U1341 (N_1341,In_1385,In_566);
and U1342 (N_1342,In_496,In_1300);
nor U1343 (N_1343,In_1840,In_1547);
or U1344 (N_1344,In_996,In_758);
or U1345 (N_1345,In_1922,In_1291);
and U1346 (N_1346,In_82,In_1079);
nor U1347 (N_1347,In_1615,In_1800);
and U1348 (N_1348,In_577,In_838);
nand U1349 (N_1349,In_1475,In_225);
nand U1350 (N_1350,In_727,In_541);
and U1351 (N_1351,In_257,In_57);
nor U1352 (N_1352,In_1237,In_1786);
and U1353 (N_1353,In_1577,In_707);
nand U1354 (N_1354,In_212,In_1297);
or U1355 (N_1355,In_1095,In_1);
nand U1356 (N_1356,In_1122,In_1800);
or U1357 (N_1357,In_1284,In_1191);
or U1358 (N_1358,In_86,In_1432);
nand U1359 (N_1359,In_534,In_1398);
or U1360 (N_1360,In_600,In_1229);
xor U1361 (N_1361,In_520,In_1156);
nor U1362 (N_1362,In_859,In_266);
nor U1363 (N_1363,In_776,In_137);
nor U1364 (N_1364,In_115,In_1700);
nand U1365 (N_1365,In_1268,In_740);
or U1366 (N_1366,In_370,In_1513);
or U1367 (N_1367,In_877,In_1851);
and U1368 (N_1368,In_1240,In_1339);
or U1369 (N_1369,In_772,In_667);
or U1370 (N_1370,In_305,In_1894);
nand U1371 (N_1371,In_1297,In_1393);
xor U1372 (N_1372,In_1649,In_1647);
nand U1373 (N_1373,In_1520,In_1731);
nor U1374 (N_1374,In_332,In_1551);
nor U1375 (N_1375,In_236,In_1627);
nand U1376 (N_1376,In_70,In_1464);
and U1377 (N_1377,In_1885,In_1040);
or U1378 (N_1378,In_1318,In_86);
or U1379 (N_1379,In_1959,In_1912);
nor U1380 (N_1380,In_1066,In_849);
nand U1381 (N_1381,In_1453,In_670);
or U1382 (N_1382,In_11,In_7);
and U1383 (N_1383,In_257,In_996);
or U1384 (N_1384,In_399,In_752);
nor U1385 (N_1385,In_491,In_1771);
or U1386 (N_1386,In_656,In_1700);
and U1387 (N_1387,In_365,In_671);
or U1388 (N_1388,In_1053,In_1664);
nand U1389 (N_1389,In_490,In_1591);
nor U1390 (N_1390,In_1331,In_1441);
or U1391 (N_1391,In_1147,In_422);
nor U1392 (N_1392,In_635,In_886);
nor U1393 (N_1393,In_782,In_594);
xor U1394 (N_1394,In_93,In_790);
or U1395 (N_1395,In_241,In_365);
nand U1396 (N_1396,In_1411,In_1558);
and U1397 (N_1397,In_539,In_378);
and U1398 (N_1398,In_1971,In_1959);
and U1399 (N_1399,In_1705,In_604);
and U1400 (N_1400,In_1218,In_1825);
nand U1401 (N_1401,In_971,In_1665);
xor U1402 (N_1402,In_1775,In_2);
xnor U1403 (N_1403,In_730,In_1781);
and U1404 (N_1404,In_1206,In_1137);
or U1405 (N_1405,In_1601,In_654);
xnor U1406 (N_1406,In_266,In_802);
or U1407 (N_1407,In_983,In_1389);
nor U1408 (N_1408,In_1499,In_62);
and U1409 (N_1409,In_1090,In_1734);
nand U1410 (N_1410,In_1790,In_533);
and U1411 (N_1411,In_1840,In_440);
nor U1412 (N_1412,In_2,In_1598);
and U1413 (N_1413,In_1202,In_1376);
or U1414 (N_1414,In_1667,In_560);
and U1415 (N_1415,In_1631,In_804);
xnor U1416 (N_1416,In_1570,In_1002);
nand U1417 (N_1417,In_879,In_1756);
and U1418 (N_1418,In_8,In_116);
nand U1419 (N_1419,In_955,In_151);
nand U1420 (N_1420,In_512,In_1250);
nor U1421 (N_1421,In_1039,In_842);
nand U1422 (N_1422,In_1233,In_950);
nand U1423 (N_1423,In_1161,In_1470);
nor U1424 (N_1424,In_697,In_1073);
and U1425 (N_1425,In_95,In_18);
xor U1426 (N_1426,In_1689,In_784);
xor U1427 (N_1427,In_1296,In_549);
and U1428 (N_1428,In_1825,In_711);
or U1429 (N_1429,In_561,In_1242);
or U1430 (N_1430,In_1711,In_1128);
nand U1431 (N_1431,In_983,In_690);
nor U1432 (N_1432,In_887,In_1589);
nor U1433 (N_1433,In_1518,In_383);
and U1434 (N_1434,In_1642,In_1574);
and U1435 (N_1435,In_676,In_878);
nor U1436 (N_1436,In_480,In_829);
nand U1437 (N_1437,In_309,In_1954);
nand U1438 (N_1438,In_1680,In_1122);
nand U1439 (N_1439,In_762,In_787);
nor U1440 (N_1440,In_1816,In_795);
and U1441 (N_1441,In_419,In_510);
xor U1442 (N_1442,In_1008,In_1843);
nor U1443 (N_1443,In_669,In_377);
nor U1444 (N_1444,In_1381,In_431);
nand U1445 (N_1445,In_1892,In_1682);
nor U1446 (N_1446,In_1906,In_1578);
xnor U1447 (N_1447,In_823,In_1550);
and U1448 (N_1448,In_1454,In_187);
nor U1449 (N_1449,In_951,In_300);
or U1450 (N_1450,In_737,In_1691);
and U1451 (N_1451,In_1513,In_1687);
or U1452 (N_1452,In_1705,In_1927);
nor U1453 (N_1453,In_1147,In_1354);
and U1454 (N_1454,In_1140,In_975);
or U1455 (N_1455,In_406,In_745);
nor U1456 (N_1456,In_480,In_1833);
and U1457 (N_1457,In_17,In_1703);
nand U1458 (N_1458,In_1598,In_430);
nand U1459 (N_1459,In_1823,In_743);
xnor U1460 (N_1460,In_593,In_188);
nor U1461 (N_1461,In_832,In_1190);
or U1462 (N_1462,In_841,In_1206);
and U1463 (N_1463,In_1368,In_1522);
nand U1464 (N_1464,In_1710,In_1535);
and U1465 (N_1465,In_1413,In_613);
and U1466 (N_1466,In_710,In_1745);
nand U1467 (N_1467,In_567,In_171);
xnor U1468 (N_1468,In_1997,In_705);
nor U1469 (N_1469,In_1231,In_1983);
nand U1470 (N_1470,In_497,In_1842);
or U1471 (N_1471,In_187,In_845);
or U1472 (N_1472,In_425,In_1507);
nand U1473 (N_1473,In_195,In_783);
xor U1474 (N_1474,In_337,In_1453);
nand U1475 (N_1475,In_818,In_1996);
and U1476 (N_1476,In_34,In_589);
or U1477 (N_1477,In_727,In_1656);
or U1478 (N_1478,In_1399,In_1900);
or U1479 (N_1479,In_768,In_462);
or U1480 (N_1480,In_1389,In_1629);
nand U1481 (N_1481,In_1919,In_187);
nor U1482 (N_1482,In_398,In_1281);
nand U1483 (N_1483,In_1084,In_1570);
and U1484 (N_1484,In_1429,In_843);
and U1485 (N_1485,In_283,In_874);
nand U1486 (N_1486,In_625,In_690);
or U1487 (N_1487,In_1359,In_190);
or U1488 (N_1488,In_532,In_643);
and U1489 (N_1489,In_1716,In_1253);
nand U1490 (N_1490,In_1066,In_1021);
and U1491 (N_1491,In_46,In_1112);
and U1492 (N_1492,In_698,In_1343);
and U1493 (N_1493,In_1643,In_1199);
xor U1494 (N_1494,In_1627,In_751);
nand U1495 (N_1495,In_195,In_1592);
nor U1496 (N_1496,In_876,In_740);
and U1497 (N_1497,In_1103,In_1376);
or U1498 (N_1498,In_1249,In_975);
or U1499 (N_1499,In_318,In_1421);
xor U1500 (N_1500,In_1677,In_1120);
or U1501 (N_1501,In_209,In_1449);
or U1502 (N_1502,In_1427,In_700);
or U1503 (N_1503,In_107,In_431);
or U1504 (N_1504,In_1480,In_138);
or U1505 (N_1505,In_1352,In_1754);
and U1506 (N_1506,In_1358,In_1673);
nand U1507 (N_1507,In_752,In_1699);
xor U1508 (N_1508,In_494,In_1037);
xor U1509 (N_1509,In_364,In_1363);
or U1510 (N_1510,In_118,In_1900);
or U1511 (N_1511,In_518,In_1160);
and U1512 (N_1512,In_1072,In_168);
or U1513 (N_1513,In_1244,In_569);
and U1514 (N_1514,In_101,In_1994);
and U1515 (N_1515,In_257,In_1946);
and U1516 (N_1516,In_511,In_1042);
and U1517 (N_1517,In_1872,In_558);
xor U1518 (N_1518,In_963,In_1132);
xnor U1519 (N_1519,In_1506,In_829);
and U1520 (N_1520,In_1729,In_1464);
or U1521 (N_1521,In_1643,In_66);
or U1522 (N_1522,In_180,In_734);
and U1523 (N_1523,In_811,In_264);
nand U1524 (N_1524,In_167,In_1194);
or U1525 (N_1525,In_1736,In_1870);
xnor U1526 (N_1526,In_1459,In_1313);
nor U1527 (N_1527,In_1099,In_106);
nor U1528 (N_1528,In_1868,In_415);
or U1529 (N_1529,In_376,In_571);
and U1530 (N_1530,In_510,In_36);
xor U1531 (N_1531,In_561,In_1035);
and U1532 (N_1532,In_1437,In_1712);
or U1533 (N_1533,In_1222,In_350);
and U1534 (N_1534,In_1162,In_778);
nand U1535 (N_1535,In_1949,In_754);
or U1536 (N_1536,In_330,In_1180);
nor U1537 (N_1537,In_1277,In_208);
nand U1538 (N_1538,In_1717,In_491);
or U1539 (N_1539,In_552,In_1761);
nand U1540 (N_1540,In_1420,In_758);
nor U1541 (N_1541,In_79,In_1835);
or U1542 (N_1542,In_255,In_1140);
nand U1543 (N_1543,In_1911,In_1096);
nor U1544 (N_1544,In_1343,In_1338);
nor U1545 (N_1545,In_45,In_286);
and U1546 (N_1546,In_842,In_1872);
or U1547 (N_1547,In_288,In_404);
nand U1548 (N_1548,In_487,In_1530);
or U1549 (N_1549,In_1120,In_1868);
nor U1550 (N_1550,In_1866,In_1381);
nand U1551 (N_1551,In_1053,In_635);
nand U1552 (N_1552,In_509,In_1226);
or U1553 (N_1553,In_1785,In_651);
nand U1554 (N_1554,In_1822,In_307);
nand U1555 (N_1555,In_1370,In_823);
and U1556 (N_1556,In_528,In_438);
nor U1557 (N_1557,In_1007,In_1340);
nor U1558 (N_1558,In_1738,In_1134);
nor U1559 (N_1559,In_719,In_709);
or U1560 (N_1560,In_547,In_1213);
nand U1561 (N_1561,In_1901,In_453);
nand U1562 (N_1562,In_733,In_929);
nand U1563 (N_1563,In_884,In_593);
and U1564 (N_1564,In_670,In_1945);
xor U1565 (N_1565,In_1755,In_306);
nand U1566 (N_1566,In_1544,In_916);
nand U1567 (N_1567,In_150,In_1190);
nor U1568 (N_1568,In_1182,In_779);
nand U1569 (N_1569,In_519,In_664);
nand U1570 (N_1570,In_1539,In_1573);
nand U1571 (N_1571,In_800,In_1035);
or U1572 (N_1572,In_1406,In_1820);
xnor U1573 (N_1573,In_74,In_1567);
nor U1574 (N_1574,In_661,In_1523);
nand U1575 (N_1575,In_566,In_263);
and U1576 (N_1576,In_888,In_1009);
and U1577 (N_1577,In_857,In_1892);
or U1578 (N_1578,In_897,In_1742);
nor U1579 (N_1579,In_1738,In_1628);
nand U1580 (N_1580,In_1824,In_1652);
and U1581 (N_1581,In_723,In_922);
nand U1582 (N_1582,In_1120,In_691);
nor U1583 (N_1583,In_1573,In_764);
nor U1584 (N_1584,In_964,In_384);
nand U1585 (N_1585,In_1756,In_1440);
nand U1586 (N_1586,In_58,In_1177);
nand U1587 (N_1587,In_1768,In_1512);
and U1588 (N_1588,In_488,In_256);
nor U1589 (N_1589,In_363,In_695);
nand U1590 (N_1590,In_926,In_766);
and U1591 (N_1591,In_428,In_581);
and U1592 (N_1592,In_674,In_1401);
or U1593 (N_1593,In_448,In_1392);
nand U1594 (N_1594,In_1156,In_553);
and U1595 (N_1595,In_445,In_549);
nor U1596 (N_1596,In_65,In_1586);
nand U1597 (N_1597,In_968,In_976);
nor U1598 (N_1598,In_1493,In_480);
and U1599 (N_1599,In_655,In_1986);
nand U1600 (N_1600,In_577,In_1293);
or U1601 (N_1601,In_925,In_1464);
nand U1602 (N_1602,In_26,In_467);
xor U1603 (N_1603,In_1915,In_555);
nor U1604 (N_1604,In_707,In_1641);
nor U1605 (N_1605,In_1547,In_859);
nor U1606 (N_1606,In_903,In_855);
and U1607 (N_1607,In_429,In_1380);
or U1608 (N_1608,In_1780,In_210);
and U1609 (N_1609,In_616,In_682);
and U1610 (N_1610,In_436,In_151);
and U1611 (N_1611,In_1790,In_414);
nor U1612 (N_1612,In_277,In_1275);
and U1613 (N_1613,In_406,In_417);
nand U1614 (N_1614,In_1928,In_1488);
nor U1615 (N_1615,In_1516,In_1901);
or U1616 (N_1616,In_727,In_305);
or U1617 (N_1617,In_1609,In_163);
xor U1618 (N_1618,In_1705,In_409);
nor U1619 (N_1619,In_373,In_769);
nor U1620 (N_1620,In_1549,In_1906);
and U1621 (N_1621,In_356,In_1304);
and U1622 (N_1622,In_1743,In_685);
and U1623 (N_1623,In_1018,In_1589);
nor U1624 (N_1624,In_201,In_840);
nor U1625 (N_1625,In_209,In_939);
xor U1626 (N_1626,In_777,In_76);
or U1627 (N_1627,In_1127,In_998);
and U1628 (N_1628,In_1566,In_1290);
xor U1629 (N_1629,In_912,In_1962);
nand U1630 (N_1630,In_1715,In_1687);
and U1631 (N_1631,In_1747,In_1391);
or U1632 (N_1632,In_1305,In_460);
or U1633 (N_1633,In_1058,In_813);
and U1634 (N_1634,In_917,In_240);
nor U1635 (N_1635,In_201,In_1075);
nand U1636 (N_1636,In_131,In_864);
and U1637 (N_1637,In_1266,In_1933);
or U1638 (N_1638,In_1661,In_402);
nand U1639 (N_1639,In_219,In_1174);
or U1640 (N_1640,In_1898,In_245);
nor U1641 (N_1641,In_369,In_488);
and U1642 (N_1642,In_751,In_1997);
or U1643 (N_1643,In_1455,In_1843);
or U1644 (N_1644,In_1585,In_828);
or U1645 (N_1645,In_698,In_1009);
nor U1646 (N_1646,In_90,In_394);
and U1647 (N_1647,In_64,In_1007);
and U1648 (N_1648,In_1012,In_1730);
nand U1649 (N_1649,In_897,In_328);
nor U1650 (N_1650,In_158,In_1763);
and U1651 (N_1651,In_168,In_247);
or U1652 (N_1652,In_1847,In_476);
nand U1653 (N_1653,In_1468,In_1589);
nand U1654 (N_1654,In_1902,In_1568);
nand U1655 (N_1655,In_1187,In_623);
and U1656 (N_1656,In_1997,In_950);
or U1657 (N_1657,In_1174,In_834);
xnor U1658 (N_1658,In_1282,In_664);
and U1659 (N_1659,In_13,In_43);
or U1660 (N_1660,In_1210,In_1066);
xor U1661 (N_1661,In_1368,In_1307);
or U1662 (N_1662,In_1464,In_1839);
or U1663 (N_1663,In_998,In_1126);
nor U1664 (N_1664,In_392,In_744);
or U1665 (N_1665,In_105,In_1021);
and U1666 (N_1666,In_1265,In_966);
nand U1667 (N_1667,In_1553,In_1881);
xnor U1668 (N_1668,In_1724,In_405);
or U1669 (N_1669,In_276,In_1164);
nand U1670 (N_1670,In_1131,In_848);
nor U1671 (N_1671,In_1770,In_345);
nand U1672 (N_1672,In_524,In_1556);
or U1673 (N_1673,In_611,In_458);
nand U1674 (N_1674,In_129,In_566);
nand U1675 (N_1675,In_1038,In_289);
or U1676 (N_1676,In_1271,In_94);
xnor U1677 (N_1677,In_691,In_1504);
xor U1678 (N_1678,In_477,In_1142);
nor U1679 (N_1679,In_61,In_1947);
and U1680 (N_1680,In_451,In_884);
nand U1681 (N_1681,In_1239,In_470);
nand U1682 (N_1682,In_194,In_950);
and U1683 (N_1683,In_893,In_1464);
nor U1684 (N_1684,In_627,In_245);
nand U1685 (N_1685,In_577,In_588);
and U1686 (N_1686,In_812,In_1700);
nand U1687 (N_1687,In_224,In_763);
and U1688 (N_1688,In_1407,In_1458);
and U1689 (N_1689,In_1073,In_84);
nand U1690 (N_1690,In_705,In_1271);
nand U1691 (N_1691,In_35,In_1212);
nor U1692 (N_1692,In_150,In_1703);
and U1693 (N_1693,In_990,In_1843);
xor U1694 (N_1694,In_1022,In_1961);
nand U1695 (N_1695,In_141,In_164);
or U1696 (N_1696,In_633,In_1564);
or U1697 (N_1697,In_1774,In_817);
nor U1698 (N_1698,In_176,In_1546);
nand U1699 (N_1699,In_1457,In_161);
or U1700 (N_1700,In_129,In_240);
and U1701 (N_1701,In_355,In_1972);
and U1702 (N_1702,In_1793,In_846);
xnor U1703 (N_1703,In_1961,In_1928);
nand U1704 (N_1704,In_1360,In_1555);
nand U1705 (N_1705,In_1850,In_1894);
or U1706 (N_1706,In_1729,In_245);
and U1707 (N_1707,In_640,In_1049);
nand U1708 (N_1708,In_1511,In_153);
nor U1709 (N_1709,In_1641,In_1055);
xor U1710 (N_1710,In_882,In_1870);
and U1711 (N_1711,In_930,In_906);
or U1712 (N_1712,In_252,In_89);
nor U1713 (N_1713,In_1541,In_1795);
nor U1714 (N_1714,In_32,In_953);
nor U1715 (N_1715,In_1603,In_1536);
or U1716 (N_1716,In_1154,In_612);
and U1717 (N_1717,In_712,In_1731);
xor U1718 (N_1718,In_880,In_1795);
nor U1719 (N_1719,In_1715,In_684);
nor U1720 (N_1720,In_1001,In_1643);
or U1721 (N_1721,In_371,In_607);
nand U1722 (N_1722,In_316,In_880);
or U1723 (N_1723,In_19,In_415);
and U1724 (N_1724,In_1539,In_1144);
and U1725 (N_1725,In_948,In_403);
or U1726 (N_1726,In_1004,In_1576);
nand U1727 (N_1727,In_1793,In_58);
nand U1728 (N_1728,In_1865,In_1995);
nand U1729 (N_1729,In_291,In_259);
and U1730 (N_1730,In_508,In_1838);
nor U1731 (N_1731,In_1123,In_1258);
nor U1732 (N_1732,In_697,In_1709);
xor U1733 (N_1733,In_1008,In_2);
and U1734 (N_1734,In_398,In_347);
nor U1735 (N_1735,In_780,In_1495);
nor U1736 (N_1736,In_1446,In_1795);
xnor U1737 (N_1737,In_374,In_1079);
or U1738 (N_1738,In_1496,In_25);
nor U1739 (N_1739,In_205,In_43);
nor U1740 (N_1740,In_237,In_1122);
nand U1741 (N_1741,In_274,In_362);
nor U1742 (N_1742,In_1822,In_1396);
nand U1743 (N_1743,In_1102,In_1679);
or U1744 (N_1744,In_277,In_1511);
nand U1745 (N_1745,In_918,In_1833);
nor U1746 (N_1746,In_1048,In_865);
nand U1747 (N_1747,In_517,In_1147);
nand U1748 (N_1748,In_763,In_713);
nand U1749 (N_1749,In_1131,In_69);
xor U1750 (N_1750,In_92,In_1518);
and U1751 (N_1751,In_698,In_607);
xor U1752 (N_1752,In_455,In_1742);
xnor U1753 (N_1753,In_631,In_1549);
and U1754 (N_1754,In_400,In_1381);
xnor U1755 (N_1755,In_266,In_860);
and U1756 (N_1756,In_1103,In_1039);
nor U1757 (N_1757,In_1484,In_1041);
and U1758 (N_1758,In_820,In_424);
or U1759 (N_1759,In_1252,In_1163);
or U1760 (N_1760,In_1557,In_668);
nor U1761 (N_1761,In_332,In_399);
and U1762 (N_1762,In_724,In_930);
and U1763 (N_1763,In_573,In_1406);
xnor U1764 (N_1764,In_47,In_294);
xor U1765 (N_1765,In_1616,In_720);
xor U1766 (N_1766,In_211,In_287);
nand U1767 (N_1767,In_257,In_186);
nand U1768 (N_1768,In_90,In_867);
or U1769 (N_1769,In_899,In_809);
nor U1770 (N_1770,In_637,In_433);
and U1771 (N_1771,In_1446,In_1922);
or U1772 (N_1772,In_558,In_1938);
or U1773 (N_1773,In_84,In_331);
nand U1774 (N_1774,In_1314,In_833);
nor U1775 (N_1775,In_1658,In_1166);
nand U1776 (N_1776,In_510,In_1511);
nor U1777 (N_1777,In_1720,In_1357);
and U1778 (N_1778,In_1733,In_824);
or U1779 (N_1779,In_1293,In_137);
or U1780 (N_1780,In_1359,In_297);
and U1781 (N_1781,In_974,In_338);
or U1782 (N_1782,In_450,In_1222);
and U1783 (N_1783,In_1810,In_1967);
nor U1784 (N_1784,In_111,In_46);
and U1785 (N_1785,In_304,In_1530);
or U1786 (N_1786,In_1491,In_13);
or U1787 (N_1787,In_206,In_1066);
nor U1788 (N_1788,In_435,In_887);
nand U1789 (N_1789,In_1709,In_936);
or U1790 (N_1790,In_376,In_589);
and U1791 (N_1791,In_1102,In_1464);
nand U1792 (N_1792,In_1144,In_1659);
or U1793 (N_1793,In_363,In_1583);
and U1794 (N_1794,In_979,In_1186);
nand U1795 (N_1795,In_1667,In_1256);
and U1796 (N_1796,In_1195,In_1586);
nand U1797 (N_1797,In_238,In_776);
and U1798 (N_1798,In_1440,In_518);
and U1799 (N_1799,In_141,In_966);
nand U1800 (N_1800,In_367,In_1997);
nand U1801 (N_1801,In_242,In_430);
nand U1802 (N_1802,In_56,In_1878);
or U1803 (N_1803,In_313,In_1160);
or U1804 (N_1804,In_433,In_860);
xnor U1805 (N_1805,In_1018,In_879);
or U1806 (N_1806,In_1897,In_1405);
and U1807 (N_1807,In_1468,In_753);
nand U1808 (N_1808,In_1972,In_1434);
or U1809 (N_1809,In_801,In_1399);
or U1810 (N_1810,In_799,In_1831);
and U1811 (N_1811,In_257,In_982);
nand U1812 (N_1812,In_399,In_287);
nand U1813 (N_1813,In_1394,In_439);
or U1814 (N_1814,In_614,In_783);
nor U1815 (N_1815,In_1216,In_2);
nand U1816 (N_1816,In_149,In_614);
nor U1817 (N_1817,In_1958,In_693);
nand U1818 (N_1818,In_843,In_1124);
and U1819 (N_1819,In_224,In_1131);
nand U1820 (N_1820,In_392,In_824);
nor U1821 (N_1821,In_1979,In_1955);
and U1822 (N_1822,In_1362,In_537);
xnor U1823 (N_1823,In_1836,In_628);
nand U1824 (N_1824,In_671,In_1218);
nor U1825 (N_1825,In_1308,In_1023);
nor U1826 (N_1826,In_1558,In_1523);
and U1827 (N_1827,In_1703,In_806);
nor U1828 (N_1828,In_358,In_653);
nor U1829 (N_1829,In_1870,In_851);
and U1830 (N_1830,In_1552,In_746);
nor U1831 (N_1831,In_1200,In_1268);
and U1832 (N_1832,In_998,In_993);
nor U1833 (N_1833,In_1151,In_1831);
nand U1834 (N_1834,In_1000,In_1170);
xnor U1835 (N_1835,In_691,In_100);
or U1836 (N_1836,In_1521,In_823);
nand U1837 (N_1837,In_959,In_1900);
and U1838 (N_1838,In_763,In_302);
nor U1839 (N_1839,In_682,In_549);
nand U1840 (N_1840,In_1150,In_1831);
or U1841 (N_1841,In_1438,In_1234);
xnor U1842 (N_1842,In_1611,In_182);
nor U1843 (N_1843,In_1414,In_1835);
or U1844 (N_1844,In_463,In_916);
or U1845 (N_1845,In_1864,In_1516);
and U1846 (N_1846,In_1777,In_23);
nand U1847 (N_1847,In_365,In_302);
or U1848 (N_1848,In_296,In_1748);
nand U1849 (N_1849,In_1882,In_1461);
or U1850 (N_1850,In_1531,In_856);
nand U1851 (N_1851,In_837,In_1504);
nand U1852 (N_1852,In_1136,In_1816);
or U1853 (N_1853,In_1274,In_620);
xnor U1854 (N_1854,In_393,In_1836);
nand U1855 (N_1855,In_316,In_1783);
nor U1856 (N_1856,In_1514,In_183);
and U1857 (N_1857,In_768,In_1772);
nand U1858 (N_1858,In_803,In_538);
nor U1859 (N_1859,In_1247,In_428);
and U1860 (N_1860,In_823,In_1392);
nand U1861 (N_1861,In_549,In_1061);
xnor U1862 (N_1862,In_829,In_830);
and U1863 (N_1863,In_1846,In_1704);
and U1864 (N_1864,In_849,In_1441);
xnor U1865 (N_1865,In_562,In_279);
nor U1866 (N_1866,In_1867,In_1560);
xor U1867 (N_1867,In_229,In_23);
nor U1868 (N_1868,In_1446,In_1740);
and U1869 (N_1869,In_1160,In_1548);
and U1870 (N_1870,In_1626,In_126);
nand U1871 (N_1871,In_1844,In_423);
or U1872 (N_1872,In_1313,In_1449);
or U1873 (N_1873,In_700,In_1550);
or U1874 (N_1874,In_1612,In_0);
or U1875 (N_1875,In_837,In_703);
nor U1876 (N_1876,In_97,In_891);
or U1877 (N_1877,In_441,In_1788);
or U1878 (N_1878,In_1486,In_625);
xnor U1879 (N_1879,In_628,In_669);
xor U1880 (N_1880,In_720,In_225);
or U1881 (N_1881,In_1243,In_1928);
or U1882 (N_1882,In_698,In_1236);
nor U1883 (N_1883,In_1364,In_1721);
and U1884 (N_1884,In_1072,In_1500);
and U1885 (N_1885,In_981,In_1229);
or U1886 (N_1886,In_655,In_1330);
nand U1887 (N_1887,In_1833,In_632);
nor U1888 (N_1888,In_43,In_757);
and U1889 (N_1889,In_49,In_847);
nand U1890 (N_1890,In_524,In_750);
nor U1891 (N_1891,In_696,In_892);
nor U1892 (N_1892,In_33,In_664);
nand U1893 (N_1893,In_958,In_1708);
nand U1894 (N_1894,In_1982,In_852);
or U1895 (N_1895,In_682,In_508);
and U1896 (N_1896,In_1396,In_1177);
or U1897 (N_1897,In_912,In_1978);
nand U1898 (N_1898,In_1904,In_1621);
nor U1899 (N_1899,In_176,In_118);
or U1900 (N_1900,In_369,In_891);
and U1901 (N_1901,In_1093,In_1781);
nor U1902 (N_1902,In_5,In_1496);
nand U1903 (N_1903,In_1373,In_515);
xor U1904 (N_1904,In_65,In_301);
and U1905 (N_1905,In_1016,In_137);
and U1906 (N_1906,In_301,In_1292);
or U1907 (N_1907,In_1712,In_318);
and U1908 (N_1908,In_1349,In_1063);
nand U1909 (N_1909,In_961,In_1259);
nor U1910 (N_1910,In_881,In_1899);
nand U1911 (N_1911,In_1879,In_1086);
and U1912 (N_1912,In_681,In_776);
or U1913 (N_1913,In_262,In_1325);
and U1914 (N_1914,In_1794,In_1051);
or U1915 (N_1915,In_361,In_1781);
nor U1916 (N_1916,In_1836,In_1933);
and U1917 (N_1917,In_1712,In_1429);
nand U1918 (N_1918,In_1961,In_608);
or U1919 (N_1919,In_25,In_1657);
and U1920 (N_1920,In_1028,In_1583);
or U1921 (N_1921,In_936,In_1113);
nor U1922 (N_1922,In_1439,In_825);
and U1923 (N_1923,In_1443,In_434);
nand U1924 (N_1924,In_48,In_1585);
or U1925 (N_1925,In_1426,In_108);
or U1926 (N_1926,In_1314,In_856);
and U1927 (N_1927,In_1701,In_1730);
and U1928 (N_1928,In_1732,In_1757);
nor U1929 (N_1929,In_355,In_1072);
and U1930 (N_1930,In_1401,In_354);
nand U1931 (N_1931,In_1810,In_955);
and U1932 (N_1932,In_1858,In_854);
and U1933 (N_1933,In_383,In_1182);
nand U1934 (N_1934,In_1617,In_966);
nor U1935 (N_1935,In_276,In_1955);
nand U1936 (N_1936,In_369,In_548);
or U1937 (N_1937,In_232,In_1484);
xor U1938 (N_1938,In_992,In_545);
nor U1939 (N_1939,In_1458,In_771);
xnor U1940 (N_1940,In_147,In_74);
or U1941 (N_1941,In_204,In_500);
or U1942 (N_1942,In_1961,In_1823);
or U1943 (N_1943,In_1202,In_885);
nor U1944 (N_1944,In_1128,In_403);
nor U1945 (N_1945,In_849,In_67);
nand U1946 (N_1946,In_1439,In_1600);
nor U1947 (N_1947,In_364,In_1933);
nor U1948 (N_1948,In_1066,In_896);
nor U1949 (N_1949,In_1277,In_1854);
and U1950 (N_1950,In_930,In_577);
or U1951 (N_1951,In_335,In_812);
nand U1952 (N_1952,In_287,In_1554);
nor U1953 (N_1953,In_1348,In_376);
xnor U1954 (N_1954,In_874,In_1294);
nor U1955 (N_1955,In_658,In_534);
or U1956 (N_1956,In_436,In_1766);
nor U1957 (N_1957,In_1753,In_1111);
nand U1958 (N_1958,In_191,In_1226);
or U1959 (N_1959,In_363,In_1368);
and U1960 (N_1960,In_813,In_357);
nor U1961 (N_1961,In_1936,In_1468);
and U1962 (N_1962,In_641,In_318);
nand U1963 (N_1963,In_1734,In_613);
nand U1964 (N_1964,In_384,In_1263);
or U1965 (N_1965,In_1615,In_843);
nand U1966 (N_1966,In_1368,In_1544);
and U1967 (N_1967,In_1679,In_1487);
and U1968 (N_1968,In_1124,In_1179);
and U1969 (N_1969,In_302,In_520);
nand U1970 (N_1970,In_341,In_643);
or U1971 (N_1971,In_1845,In_544);
nand U1972 (N_1972,In_672,In_893);
or U1973 (N_1973,In_973,In_684);
nand U1974 (N_1974,In_827,In_675);
nand U1975 (N_1975,In_389,In_1074);
nor U1976 (N_1976,In_86,In_456);
nand U1977 (N_1977,In_1390,In_166);
or U1978 (N_1978,In_1042,In_1021);
xor U1979 (N_1979,In_1985,In_1133);
or U1980 (N_1980,In_1737,In_471);
or U1981 (N_1981,In_319,In_135);
and U1982 (N_1982,In_648,In_1479);
nand U1983 (N_1983,In_1596,In_1788);
nor U1984 (N_1984,In_657,In_1099);
nor U1985 (N_1985,In_706,In_338);
nand U1986 (N_1986,In_467,In_524);
or U1987 (N_1987,In_710,In_384);
or U1988 (N_1988,In_114,In_996);
and U1989 (N_1989,In_1877,In_1712);
and U1990 (N_1990,In_1909,In_1229);
nand U1991 (N_1991,In_567,In_226);
and U1992 (N_1992,In_917,In_1614);
nand U1993 (N_1993,In_1669,In_1636);
xor U1994 (N_1994,In_732,In_1810);
and U1995 (N_1995,In_1367,In_27);
nand U1996 (N_1996,In_361,In_1087);
or U1997 (N_1997,In_1920,In_555);
or U1998 (N_1998,In_1575,In_1678);
and U1999 (N_1999,In_1299,In_1988);
and U2000 (N_2000,In_614,In_346);
nand U2001 (N_2001,In_585,In_88);
nor U2002 (N_2002,In_1509,In_536);
nand U2003 (N_2003,In_1971,In_608);
or U2004 (N_2004,In_1197,In_272);
or U2005 (N_2005,In_172,In_472);
xnor U2006 (N_2006,In_979,In_1395);
nand U2007 (N_2007,In_1323,In_1014);
xor U2008 (N_2008,In_1687,In_1233);
nand U2009 (N_2009,In_1547,In_888);
nand U2010 (N_2010,In_888,In_1704);
or U2011 (N_2011,In_833,In_618);
nand U2012 (N_2012,In_358,In_964);
nand U2013 (N_2013,In_445,In_715);
and U2014 (N_2014,In_144,In_1018);
nor U2015 (N_2015,In_1901,In_95);
nand U2016 (N_2016,In_1356,In_1417);
nand U2017 (N_2017,In_1176,In_1810);
nor U2018 (N_2018,In_1491,In_900);
nand U2019 (N_2019,In_1395,In_1276);
nor U2020 (N_2020,In_1825,In_1199);
and U2021 (N_2021,In_484,In_1595);
nand U2022 (N_2022,In_430,In_1272);
nor U2023 (N_2023,In_1201,In_45);
xnor U2024 (N_2024,In_1104,In_1269);
or U2025 (N_2025,In_1927,In_1892);
xor U2026 (N_2026,In_1984,In_554);
or U2027 (N_2027,In_92,In_901);
nor U2028 (N_2028,In_253,In_1542);
and U2029 (N_2029,In_1934,In_1694);
nand U2030 (N_2030,In_1119,In_1584);
nor U2031 (N_2031,In_920,In_1208);
and U2032 (N_2032,In_1197,In_1617);
and U2033 (N_2033,In_1228,In_1765);
and U2034 (N_2034,In_430,In_426);
and U2035 (N_2035,In_1753,In_1743);
and U2036 (N_2036,In_893,In_1051);
nand U2037 (N_2037,In_89,In_225);
nand U2038 (N_2038,In_1130,In_126);
nor U2039 (N_2039,In_1535,In_1936);
xnor U2040 (N_2040,In_665,In_180);
nor U2041 (N_2041,In_358,In_1679);
or U2042 (N_2042,In_211,In_507);
and U2043 (N_2043,In_1642,In_1264);
and U2044 (N_2044,In_201,In_923);
nand U2045 (N_2045,In_269,In_1970);
nor U2046 (N_2046,In_793,In_1193);
or U2047 (N_2047,In_1852,In_1337);
nand U2048 (N_2048,In_1680,In_1381);
nand U2049 (N_2049,In_225,In_1219);
xor U2050 (N_2050,In_154,In_892);
nand U2051 (N_2051,In_288,In_287);
or U2052 (N_2052,In_105,In_1760);
nor U2053 (N_2053,In_1320,In_1483);
and U2054 (N_2054,In_835,In_513);
nand U2055 (N_2055,In_1483,In_1455);
nor U2056 (N_2056,In_1445,In_774);
or U2057 (N_2057,In_1195,In_1282);
and U2058 (N_2058,In_1343,In_153);
and U2059 (N_2059,In_894,In_1797);
and U2060 (N_2060,In_1092,In_368);
nor U2061 (N_2061,In_1840,In_839);
nor U2062 (N_2062,In_977,In_598);
nand U2063 (N_2063,In_1784,In_122);
and U2064 (N_2064,In_1793,In_1544);
or U2065 (N_2065,In_1005,In_661);
nand U2066 (N_2066,In_1315,In_990);
nor U2067 (N_2067,In_1688,In_1563);
xnor U2068 (N_2068,In_1028,In_1307);
and U2069 (N_2069,In_1853,In_1432);
or U2070 (N_2070,In_334,In_514);
or U2071 (N_2071,In_1739,In_121);
and U2072 (N_2072,In_202,In_1095);
and U2073 (N_2073,In_1065,In_1197);
and U2074 (N_2074,In_1237,In_1425);
and U2075 (N_2075,In_308,In_151);
nor U2076 (N_2076,In_1613,In_789);
and U2077 (N_2077,In_997,In_1410);
nor U2078 (N_2078,In_1724,In_334);
nand U2079 (N_2079,In_1413,In_984);
or U2080 (N_2080,In_556,In_646);
or U2081 (N_2081,In_483,In_427);
nor U2082 (N_2082,In_596,In_1272);
and U2083 (N_2083,In_1111,In_799);
nand U2084 (N_2084,In_903,In_1896);
nand U2085 (N_2085,In_1723,In_1483);
and U2086 (N_2086,In_928,In_756);
and U2087 (N_2087,In_378,In_1491);
or U2088 (N_2088,In_1376,In_1391);
or U2089 (N_2089,In_1602,In_1311);
nand U2090 (N_2090,In_293,In_1230);
nand U2091 (N_2091,In_1596,In_1939);
nor U2092 (N_2092,In_135,In_1199);
nand U2093 (N_2093,In_1965,In_70);
nand U2094 (N_2094,In_258,In_1824);
xor U2095 (N_2095,In_520,In_1784);
nor U2096 (N_2096,In_1005,In_365);
or U2097 (N_2097,In_1813,In_1869);
nand U2098 (N_2098,In_455,In_1672);
nor U2099 (N_2099,In_613,In_1036);
nand U2100 (N_2100,In_677,In_1877);
nand U2101 (N_2101,In_1700,In_139);
nand U2102 (N_2102,In_972,In_729);
nor U2103 (N_2103,In_1874,In_1249);
nor U2104 (N_2104,In_1694,In_1817);
nand U2105 (N_2105,In_161,In_440);
nor U2106 (N_2106,In_1407,In_1700);
xnor U2107 (N_2107,In_1208,In_794);
and U2108 (N_2108,In_814,In_1200);
nand U2109 (N_2109,In_1120,In_1162);
or U2110 (N_2110,In_971,In_1478);
and U2111 (N_2111,In_25,In_472);
nor U2112 (N_2112,In_885,In_529);
and U2113 (N_2113,In_639,In_207);
or U2114 (N_2114,In_189,In_5);
nor U2115 (N_2115,In_768,In_1331);
and U2116 (N_2116,In_1710,In_929);
xnor U2117 (N_2117,In_405,In_1232);
nand U2118 (N_2118,In_993,In_649);
or U2119 (N_2119,In_1444,In_908);
xor U2120 (N_2120,In_191,In_280);
and U2121 (N_2121,In_600,In_1632);
nor U2122 (N_2122,In_388,In_1687);
nor U2123 (N_2123,In_1474,In_1592);
or U2124 (N_2124,In_1317,In_351);
or U2125 (N_2125,In_1790,In_1584);
and U2126 (N_2126,In_1391,In_29);
or U2127 (N_2127,In_595,In_1285);
nor U2128 (N_2128,In_959,In_1705);
and U2129 (N_2129,In_1714,In_650);
nand U2130 (N_2130,In_669,In_102);
or U2131 (N_2131,In_1338,In_1904);
and U2132 (N_2132,In_1712,In_1237);
nand U2133 (N_2133,In_684,In_1406);
or U2134 (N_2134,In_1383,In_694);
nand U2135 (N_2135,In_341,In_132);
nor U2136 (N_2136,In_562,In_323);
nor U2137 (N_2137,In_1110,In_1733);
nand U2138 (N_2138,In_1764,In_22);
nor U2139 (N_2139,In_1411,In_331);
or U2140 (N_2140,In_1019,In_1361);
xor U2141 (N_2141,In_1608,In_155);
and U2142 (N_2142,In_779,In_172);
nand U2143 (N_2143,In_853,In_100);
or U2144 (N_2144,In_328,In_1191);
nor U2145 (N_2145,In_1114,In_1554);
and U2146 (N_2146,In_252,In_624);
xor U2147 (N_2147,In_690,In_1843);
and U2148 (N_2148,In_698,In_434);
nor U2149 (N_2149,In_400,In_479);
and U2150 (N_2150,In_350,In_1377);
or U2151 (N_2151,In_1979,In_1417);
and U2152 (N_2152,In_69,In_1325);
xor U2153 (N_2153,In_584,In_870);
nand U2154 (N_2154,In_1414,In_1405);
nand U2155 (N_2155,In_1287,In_671);
nor U2156 (N_2156,In_1126,In_1832);
or U2157 (N_2157,In_202,In_1891);
xor U2158 (N_2158,In_1453,In_976);
nor U2159 (N_2159,In_1189,In_1282);
or U2160 (N_2160,In_1386,In_970);
or U2161 (N_2161,In_61,In_1981);
and U2162 (N_2162,In_301,In_751);
or U2163 (N_2163,In_368,In_212);
nor U2164 (N_2164,In_1350,In_10);
nor U2165 (N_2165,In_198,In_230);
xor U2166 (N_2166,In_436,In_1730);
xor U2167 (N_2167,In_1053,In_852);
and U2168 (N_2168,In_1229,In_311);
or U2169 (N_2169,In_13,In_1881);
and U2170 (N_2170,In_1784,In_408);
or U2171 (N_2171,In_636,In_1939);
nand U2172 (N_2172,In_1418,In_1357);
nor U2173 (N_2173,In_1268,In_1675);
nand U2174 (N_2174,In_545,In_411);
nor U2175 (N_2175,In_1406,In_1260);
and U2176 (N_2176,In_617,In_945);
nand U2177 (N_2177,In_769,In_323);
nor U2178 (N_2178,In_1235,In_440);
nor U2179 (N_2179,In_1594,In_1114);
nor U2180 (N_2180,In_1217,In_1962);
xnor U2181 (N_2181,In_655,In_317);
nor U2182 (N_2182,In_1654,In_619);
nor U2183 (N_2183,In_1036,In_75);
nand U2184 (N_2184,In_1771,In_436);
nand U2185 (N_2185,In_187,In_1979);
or U2186 (N_2186,In_599,In_1010);
or U2187 (N_2187,In_783,In_1586);
nor U2188 (N_2188,In_1000,In_1603);
nand U2189 (N_2189,In_311,In_1854);
nand U2190 (N_2190,In_1254,In_1909);
nand U2191 (N_2191,In_90,In_1545);
or U2192 (N_2192,In_188,In_1548);
nand U2193 (N_2193,In_1965,In_1958);
and U2194 (N_2194,In_1626,In_27);
nand U2195 (N_2195,In_1015,In_637);
nand U2196 (N_2196,In_418,In_4);
or U2197 (N_2197,In_991,In_938);
nand U2198 (N_2198,In_1531,In_1660);
nand U2199 (N_2199,In_122,In_1441);
or U2200 (N_2200,In_1676,In_563);
xnor U2201 (N_2201,In_120,In_1655);
xor U2202 (N_2202,In_420,In_399);
or U2203 (N_2203,In_471,In_1443);
or U2204 (N_2204,In_703,In_1953);
nor U2205 (N_2205,In_239,In_1095);
nor U2206 (N_2206,In_656,In_37);
nor U2207 (N_2207,In_945,In_874);
nor U2208 (N_2208,In_1644,In_1458);
nand U2209 (N_2209,In_308,In_384);
and U2210 (N_2210,In_1110,In_755);
or U2211 (N_2211,In_737,In_259);
nor U2212 (N_2212,In_1051,In_1232);
nor U2213 (N_2213,In_1648,In_1248);
nor U2214 (N_2214,In_1241,In_1772);
and U2215 (N_2215,In_365,In_316);
nor U2216 (N_2216,In_1213,In_287);
nand U2217 (N_2217,In_470,In_155);
nand U2218 (N_2218,In_1022,In_1684);
and U2219 (N_2219,In_15,In_19);
or U2220 (N_2220,In_1569,In_557);
nand U2221 (N_2221,In_777,In_371);
or U2222 (N_2222,In_112,In_1431);
nand U2223 (N_2223,In_1186,In_52);
and U2224 (N_2224,In_407,In_366);
nor U2225 (N_2225,In_465,In_426);
and U2226 (N_2226,In_1937,In_618);
or U2227 (N_2227,In_536,In_230);
nor U2228 (N_2228,In_59,In_1283);
or U2229 (N_2229,In_1790,In_1023);
xnor U2230 (N_2230,In_1799,In_578);
or U2231 (N_2231,In_1244,In_940);
nor U2232 (N_2232,In_1221,In_402);
nor U2233 (N_2233,In_1358,In_1400);
xnor U2234 (N_2234,In_1543,In_1894);
or U2235 (N_2235,In_1283,In_710);
or U2236 (N_2236,In_147,In_1166);
and U2237 (N_2237,In_1680,In_965);
nor U2238 (N_2238,In_184,In_1110);
or U2239 (N_2239,In_1631,In_1425);
nor U2240 (N_2240,In_35,In_822);
nand U2241 (N_2241,In_735,In_945);
and U2242 (N_2242,In_334,In_1234);
and U2243 (N_2243,In_1798,In_1380);
nand U2244 (N_2244,In_428,In_1764);
or U2245 (N_2245,In_1908,In_1725);
and U2246 (N_2246,In_1388,In_626);
or U2247 (N_2247,In_469,In_273);
and U2248 (N_2248,In_416,In_946);
nor U2249 (N_2249,In_1601,In_1513);
or U2250 (N_2250,In_320,In_133);
nor U2251 (N_2251,In_690,In_1089);
nand U2252 (N_2252,In_1943,In_197);
or U2253 (N_2253,In_1046,In_854);
nand U2254 (N_2254,In_112,In_330);
nand U2255 (N_2255,In_1179,In_1397);
nor U2256 (N_2256,In_180,In_812);
nor U2257 (N_2257,In_247,In_1122);
or U2258 (N_2258,In_1878,In_419);
and U2259 (N_2259,In_542,In_8);
and U2260 (N_2260,In_939,In_1999);
nor U2261 (N_2261,In_807,In_1825);
and U2262 (N_2262,In_1767,In_1419);
and U2263 (N_2263,In_1055,In_147);
or U2264 (N_2264,In_1902,In_1085);
and U2265 (N_2265,In_1614,In_1161);
xnor U2266 (N_2266,In_1880,In_672);
nand U2267 (N_2267,In_849,In_1434);
or U2268 (N_2268,In_293,In_653);
or U2269 (N_2269,In_795,In_997);
xor U2270 (N_2270,In_201,In_1774);
xor U2271 (N_2271,In_1906,In_546);
or U2272 (N_2272,In_1900,In_608);
and U2273 (N_2273,In_238,In_390);
nor U2274 (N_2274,In_355,In_350);
or U2275 (N_2275,In_357,In_1676);
and U2276 (N_2276,In_689,In_572);
nor U2277 (N_2277,In_1122,In_1116);
xor U2278 (N_2278,In_421,In_991);
nand U2279 (N_2279,In_1521,In_1067);
nand U2280 (N_2280,In_425,In_789);
nor U2281 (N_2281,In_1135,In_586);
nand U2282 (N_2282,In_768,In_592);
or U2283 (N_2283,In_643,In_1684);
or U2284 (N_2284,In_1818,In_114);
or U2285 (N_2285,In_1697,In_395);
and U2286 (N_2286,In_218,In_873);
or U2287 (N_2287,In_389,In_1384);
or U2288 (N_2288,In_807,In_193);
nand U2289 (N_2289,In_1449,In_1021);
and U2290 (N_2290,In_11,In_1018);
nand U2291 (N_2291,In_1172,In_1793);
and U2292 (N_2292,In_1353,In_251);
nand U2293 (N_2293,In_1102,In_1460);
nor U2294 (N_2294,In_819,In_539);
and U2295 (N_2295,In_1123,In_405);
and U2296 (N_2296,In_959,In_1578);
nand U2297 (N_2297,In_768,In_717);
or U2298 (N_2298,In_1557,In_599);
and U2299 (N_2299,In_1771,In_1694);
or U2300 (N_2300,In_188,In_486);
or U2301 (N_2301,In_632,In_739);
nor U2302 (N_2302,In_1638,In_295);
or U2303 (N_2303,In_1542,In_360);
nor U2304 (N_2304,In_1343,In_1620);
nor U2305 (N_2305,In_250,In_98);
or U2306 (N_2306,In_403,In_1734);
nor U2307 (N_2307,In_663,In_624);
nor U2308 (N_2308,In_1096,In_1678);
or U2309 (N_2309,In_1935,In_1916);
nor U2310 (N_2310,In_1564,In_737);
nand U2311 (N_2311,In_1568,In_5);
and U2312 (N_2312,In_305,In_545);
and U2313 (N_2313,In_75,In_268);
and U2314 (N_2314,In_1865,In_1651);
or U2315 (N_2315,In_1348,In_1277);
nor U2316 (N_2316,In_70,In_1020);
xnor U2317 (N_2317,In_755,In_1658);
nand U2318 (N_2318,In_1106,In_1107);
and U2319 (N_2319,In_1970,In_271);
and U2320 (N_2320,In_1996,In_1771);
and U2321 (N_2321,In_1420,In_963);
nor U2322 (N_2322,In_1706,In_1705);
and U2323 (N_2323,In_316,In_429);
or U2324 (N_2324,In_758,In_1565);
xnor U2325 (N_2325,In_1132,In_824);
nand U2326 (N_2326,In_338,In_1031);
or U2327 (N_2327,In_430,In_155);
nand U2328 (N_2328,In_1168,In_1686);
and U2329 (N_2329,In_1671,In_1034);
or U2330 (N_2330,In_1115,In_727);
nor U2331 (N_2331,In_1191,In_157);
and U2332 (N_2332,In_30,In_605);
nand U2333 (N_2333,In_569,In_1380);
nand U2334 (N_2334,In_509,In_324);
nand U2335 (N_2335,In_577,In_439);
and U2336 (N_2336,In_1332,In_1268);
xnor U2337 (N_2337,In_1008,In_1136);
nand U2338 (N_2338,In_514,In_1383);
or U2339 (N_2339,In_166,In_1965);
and U2340 (N_2340,In_1829,In_1447);
nor U2341 (N_2341,In_1163,In_1921);
nand U2342 (N_2342,In_1743,In_1694);
xor U2343 (N_2343,In_920,In_1340);
or U2344 (N_2344,In_79,In_1186);
and U2345 (N_2345,In_35,In_1451);
xor U2346 (N_2346,In_627,In_417);
or U2347 (N_2347,In_1826,In_859);
nand U2348 (N_2348,In_1059,In_341);
or U2349 (N_2349,In_1944,In_1368);
and U2350 (N_2350,In_1159,In_1175);
nand U2351 (N_2351,In_1321,In_989);
and U2352 (N_2352,In_1139,In_1909);
and U2353 (N_2353,In_814,In_843);
and U2354 (N_2354,In_1834,In_1374);
nand U2355 (N_2355,In_1466,In_1186);
or U2356 (N_2356,In_1751,In_1033);
and U2357 (N_2357,In_143,In_1757);
or U2358 (N_2358,In_266,In_431);
nor U2359 (N_2359,In_731,In_830);
nand U2360 (N_2360,In_522,In_1957);
nand U2361 (N_2361,In_1028,In_1301);
and U2362 (N_2362,In_1614,In_74);
or U2363 (N_2363,In_243,In_394);
and U2364 (N_2364,In_118,In_623);
nand U2365 (N_2365,In_1938,In_1608);
and U2366 (N_2366,In_1946,In_1870);
or U2367 (N_2367,In_1386,In_1340);
xnor U2368 (N_2368,In_1374,In_1548);
and U2369 (N_2369,In_1012,In_1841);
and U2370 (N_2370,In_570,In_1429);
xor U2371 (N_2371,In_1015,In_1974);
and U2372 (N_2372,In_275,In_1987);
nor U2373 (N_2373,In_499,In_671);
or U2374 (N_2374,In_44,In_1030);
nor U2375 (N_2375,In_600,In_1750);
or U2376 (N_2376,In_904,In_1699);
and U2377 (N_2377,In_1741,In_873);
and U2378 (N_2378,In_523,In_891);
nand U2379 (N_2379,In_1749,In_1272);
or U2380 (N_2380,In_1778,In_1041);
nand U2381 (N_2381,In_366,In_1188);
nor U2382 (N_2382,In_907,In_1546);
nor U2383 (N_2383,In_835,In_888);
nand U2384 (N_2384,In_1488,In_1412);
or U2385 (N_2385,In_519,In_1702);
xnor U2386 (N_2386,In_678,In_297);
nor U2387 (N_2387,In_1528,In_402);
or U2388 (N_2388,In_1023,In_1632);
nor U2389 (N_2389,In_1682,In_701);
and U2390 (N_2390,In_1311,In_1162);
or U2391 (N_2391,In_776,In_1492);
nor U2392 (N_2392,In_732,In_1724);
nand U2393 (N_2393,In_1422,In_966);
or U2394 (N_2394,In_919,In_1396);
xnor U2395 (N_2395,In_101,In_134);
nor U2396 (N_2396,In_694,In_1978);
xnor U2397 (N_2397,In_1149,In_716);
nor U2398 (N_2398,In_97,In_1556);
xor U2399 (N_2399,In_268,In_1217);
or U2400 (N_2400,In_868,In_1223);
nor U2401 (N_2401,In_83,In_1143);
xor U2402 (N_2402,In_1736,In_380);
and U2403 (N_2403,In_1955,In_1307);
and U2404 (N_2404,In_789,In_1734);
nor U2405 (N_2405,In_1112,In_1491);
nand U2406 (N_2406,In_253,In_819);
and U2407 (N_2407,In_1623,In_801);
nand U2408 (N_2408,In_1459,In_1714);
or U2409 (N_2409,In_28,In_1334);
and U2410 (N_2410,In_1184,In_1099);
xnor U2411 (N_2411,In_1388,In_1730);
xor U2412 (N_2412,In_1882,In_1405);
nand U2413 (N_2413,In_1157,In_536);
and U2414 (N_2414,In_653,In_1675);
nand U2415 (N_2415,In_1936,In_791);
nand U2416 (N_2416,In_698,In_758);
xnor U2417 (N_2417,In_1383,In_1298);
or U2418 (N_2418,In_776,In_551);
and U2419 (N_2419,In_748,In_1526);
nor U2420 (N_2420,In_1304,In_1850);
nand U2421 (N_2421,In_864,In_937);
nor U2422 (N_2422,In_1309,In_1400);
or U2423 (N_2423,In_1277,In_1757);
or U2424 (N_2424,In_209,In_1576);
nor U2425 (N_2425,In_1177,In_279);
nor U2426 (N_2426,In_1478,In_1590);
nor U2427 (N_2427,In_592,In_325);
nand U2428 (N_2428,In_1802,In_1117);
and U2429 (N_2429,In_162,In_1920);
nor U2430 (N_2430,In_1171,In_973);
or U2431 (N_2431,In_779,In_1783);
nand U2432 (N_2432,In_1231,In_30);
nor U2433 (N_2433,In_738,In_365);
xnor U2434 (N_2434,In_633,In_1501);
nor U2435 (N_2435,In_1937,In_454);
nor U2436 (N_2436,In_1598,In_213);
and U2437 (N_2437,In_1059,In_1938);
and U2438 (N_2438,In_1309,In_1326);
nand U2439 (N_2439,In_1971,In_1399);
or U2440 (N_2440,In_1487,In_1032);
xnor U2441 (N_2441,In_991,In_696);
nor U2442 (N_2442,In_1487,In_1828);
or U2443 (N_2443,In_1480,In_1503);
or U2444 (N_2444,In_340,In_1210);
nor U2445 (N_2445,In_1744,In_884);
nor U2446 (N_2446,In_1483,In_429);
nor U2447 (N_2447,In_815,In_957);
and U2448 (N_2448,In_323,In_1821);
nor U2449 (N_2449,In_121,In_1171);
nand U2450 (N_2450,In_1665,In_282);
or U2451 (N_2451,In_1132,In_1109);
and U2452 (N_2452,In_27,In_1837);
nand U2453 (N_2453,In_1994,In_637);
and U2454 (N_2454,In_847,In_1272);
nor U2455 (N_2455,In_1100,In_1438);
or U2456 (N_2456,In_1483,In_948);
or U2457 (N_2457,In_582,In_1629);
and U2458 (N_2458,In_1875,In_324);
nand U2459 (N_2459,In_676,In_1114);
or U2460 (N_2460,In_1390,In_1052);
or U2461 (N_2461,In_1811,In_231);
nor U2462 (N_2462,In_198,In_1034);
or U2463 (N_2463,In_1959,In_155);
xnor U2464 (N_2464,In_1692,In_1433);
or U2465 (N_2465,In_824,In_1858);
or U2466 (N_2466,In_1822,In_1342);
and U2467 (N_2467,In_1580,In_1436);
nand U2468 (N_2468,In_1751,In_1015);
nand U2469 (N_2469,In_970,In_1236);
or U2470 (N_2470,In_202,In_651);
and U2471 (N_2471,In_1690,In_254);
or U2472 (N_2472,In_1603,In_1624);
or U2473 (N_2473,In_1475,In_439);
and U2474 (N_2474,In_172,In_252);
and U2475 (N_2475,In_1360,In_1428);
or U2476 (N_2476,In_419,In_808);
nor U2477 (N_2477,In_591,In_524);
or U2478 (N_2478,In_1231,In_1412);
or U2479 (N_2479,In_1836,In_196);
or U2480 (N_2480,In_271,In_1896);
and U2481 (N_2481,In_1466,In_856);
or U2482 (N_2482,In_263,In_1069);
and U2483 (N_2483,In_759,In_1812);
nand U2484 (N_2484,In_178,In_1748);
or U2485 (N_2485,In_550,In_405);
or U2486 (N_2486,In_465,In_1153);
nand U2487 (N_2487,In_559,In_1472);
nor U2488 (N_2488,In_1874,In_1695);
xnor U2489 (N_2489,In_1777,In_495);
and U2490 (N_2490,In_460,In_856);
nand U2491 (N_2491,In_1459,In_1892);
xor U2492 (N_2492,In_1131,In_1407);
or U2493 (N_2493,In_1617,In_835);
and U2494 (N_2494,In_1954,In_1287);
or U2495 (N_2495,In_135,In_1296);
or U2496 (N_2496,In_1404,In_681);
or U2497 (N_2497,In_1344,In_1149);
or U2498 (N_2498,In_1740,In_999);
and U2499 (N_2499,In_1951,In_353);
or U2500 (N_2500,In_783,In_251);
nand U2501 (N_2501,In_447,In_1502);
or U2502 (N_2502,In_1602,In_502);
and U2503 (N_2503,In_1203,In_229);
or U2504 (N_2504,In_1708,In_690);
and U2505 (N_2505,In_1182,In_1300);
or U2506 (N_2506,In_1014,In_1040);
nand U2507 (N_2507,In_1233,In_968);
nor U2508 (N_2508,In_683,In_1371);
nor U2509 (N_2509,In_722,In_850);
and U2510 (N_2510,In_1580,In_1819);
and U2511 (N_2511,In_1183,In_993);
nor U2512 (N_2512,In_1629,In_323);
and U2513 (N_2513,In_365,In_373);
nand U2514 (N_2514,In_176,In_587);
or U2515 (N_2515,In_1604,In_824);
nand U2516 (N_2516,In_1905,In_591);
xnor U2517 (N_2517,In_1495,In_576);
xor U2518 (N_2518,In_1726,In_1059);
nand U2519 (N_2519,In_298,In_315);
nor U2520 (N_2520,In_761,In_1098);
xnor U2521 (N_2521,In_1729,In_1175);
nand U2522 (N_2522,In_939,In_76);
nor U2523 (N_2523,In_1347,In_1859);
and U2524 (N_2524,In_1035,In_939);
nor U2525 (N_2525,In_1705,In_1789);
or U2526 (N_2526,In_773,In_281);
or U2527 (N_2527,In_1154,In_1579);
and U2528 (N_2528,In_847,In_249);
nand U2529 (N_2529,In_340,In_1983);
and U2530 (N_2530,In_1387,In_816);
nor U2531 (N_2531,In_505,In_1163);
or U2532 (N_2532,In_1610,In_718);
nor U2533 (N_2533,In_575,In_360);
and U2534 (N_2534,In_274,In_979);
xor U2535 (N_2535,In_1700,In_284);
nor U2536 (N_2536,In_879,In_1986);
or U2537 (N_2537,In_794,In_402);
or U2538 (N_2538,In_915,In_339);
or U2539 (N_2539,In_1078,In_1402);
and U2540 (N_2540,In_1311,In_1231);
nand U2541 (N_2541,In_1125,In_1080);
and U2542 (N_2542,In_1911,In_1543);
and U2543 (N_2543,In_1901,In_320);
and U2544 (N_2544,In_1993,In_66);
or U2545 (N_2545,In_509,In_364);
nor U2546 (N_2546,In_32,In_683);
or U2547 (N_2547,In_462,In_256);
or U2548 (N_2548,In_826,In_1541);
nor U2549 (N_2549,In_1384,In_1597);
and U2550 (N_2550,In_546,In_1556);
nor U2551 (N_2551,In_313,In_1881);
nor U2552 (N_2552,In_1015,In_218);
nand U2553 (N_2553,In_943,In_1667);
or U2554 (N_2554,In_1786,In_1385);
nand U2555 (N_2555,In_1175,In_339);
nor U2556 (N_2556,In_1686,In_66);
xnor U2557 (N_2557,In_363,In_597);
and U2558 (N_2558,In_1537,In_1936);
nand U2559 (N_2559,In_270,In_1428);
xnor U2560 (N_2560,In_1337,In_1252);
or U2561 (N_2561,In_1263,In_1230);
nand U2562 (N_2562,In_1024,In_759);
and U2563 (N_2563,In_282,In_1703);
and U2564 (N_2564,In_1215,In_1574);
nand U2565 (N_2565,In_912,In_1312);
and U2566 (N_2566,In_1334,In_1703);
nor U2567 (N_2567,In_1182,In_37);
xor U2568 (N_2568,In_1204,In_1731);
nor U2569 (N_2569,In_1148,In_80);
nor U2570 (N_2570,In_623,In_487);
and U2571 (N_2571,In_132,In_123);
nor U2572 (N_2572,In_1991,In_1146);
nand U2573 (N_2573,In_1580,In_657);
nor U2574 (N_2574,In_1563,In_1717);
nand U2575 (N_2575,In_1711,In_1896);
nor U2576 (N_2576,In_940,In_150);
nand U2577 (N_2577,In_649,In_223);
nand U2578 (N_2578,In_1838,In_1972);
or U2579 (N_2579,In_1070,In_239);
nor U2580 (N_2580,In_888,In_1741);
and U2581 (N_2581,In_922,In_476);
and U2582 (N_2582,In_723,In_837);
xnor U2583 (N_2583,In_1685,In_790);
xnor U2584 (N_2584,In_1667,In_1651);
xor U2585 (N_2585,In_1282,In_10);
and U2586 (N_2586,In_80,In_501);
nor U2587 (N_2587,In_524,In_316);
nor U2588 (N_2588,In_1214,In_1987);
nand U2589 (N_2589,In_149,In_1723);
and U2590 (N_2590,In_1335,In_1547);
and U2591 (N_2591,In_1030,In_878);
xnor U2592 (N_2592,In_1087,In_690);
nand U2593 (N_2593,In_1826,In_431);
or U2594 (N_2594,In_1940,In_818);
nand U2595 (N_2595,In_956,In_517);
and U2596 (N_2596,In_1250,In_415);
or U2597 (N_2597,In_1961,In_1043);
nand U2598 (N_2598,In_749,In_376);
xnor U2599 (N_2599,In_986,In_140);
or U2600 (N_2600,In_1451,In_1514);
nor U2601 (N_2601,In_1017,In_326);
nor U2602 (N_2602,In_1064,In_1243);
nor U2603 (N_2603,In_908,In_1524);
xor U2604 (N_2604,In_1000,In_814);
nand U2605 (N_2605,In_346,In_595);
nand U2606 (N_2606,In_1374,In_992);
xnor U2607 (N_2607,In_1849,In_1928);
and U2608 (N_2608,In_310,In_385);
and U2609 (N_2609,In_1614,In_1454);
nor U2610 (N_2610,In_374,In_1165);
or U2611 (N_2611,In_824,In_226);
nand U2612 (N_2612,In_1902,In_588);
nor U2613 (N_2613,In_1483,In_192);
nor U2614 (N_2614,In_1738,In_574);
nor U2615 (N_2615,In_82,In_111);
or U2616 (N_2616,In_534,In_1247);
nand U2617 (N_2617,In_483,In_798);
nor U2618 (N_2618,In_1551,In_761);
or U2619 (N_2619,In_1503,In_786);
nand U2620 (N_2620,In_910,In_82);
and U2621 (N_2621,In_124,In_910);
nand U2622 (N_2622,In_1150,In_1786);
or U2623 (N_2623,In_391,In_677);
or U2624 (N_2624,In_1421,In_953);
nor U2625 (N_2625,In_1918,In_1431);
nand U2626 (N_2626,In_1424,In_1762);
or U2627 (N_2627,In_1042,In_198);
nor U2628 (N_2628,In_1042,In_1004);
and U2629 (N_2629,In_1849,In_1161);
or U2630 (N_2630,In_177,In_1194);
nand U2631 (N_2631,In_1645,In_3);
xor U2632 (N_2632,In_1098,In_1078);
nand U2633 (N_2633,In_957,In_1472);
nand U2634 (N_2634,In_68,In_1630);
nor U2635 (N_2635,In_1795,In_1856);
nand U2636 (N_2636,In_651,In_575);
or U2637 (N_2637,In_1212,In_1611);
xor U2638 (N_2638,In_1938,In_1764);
nor U2639 (N_2639,In_1350,In_1335);
and U2640 (N_2640,In_1125,In_1110);
and U2641 (N_2641,In_1678,In_1288);
and U2642 (N_2642,In_342,In_915);
or U2643 (N_2643,In_937,In_466);
nor U2644 (N_2644,In_1812,In_65);
nor U2645 (N_2645,In_1322,In_26);
or U2646 (N_2646,In_466,In_332);
nor U2647 (N_2647,In_1260,In_746);
or U2648 (N_2648,In_718,In_824);
nor U2649 (N_2649,In_1002,In_563);
nor U2650 (N_2650,In_1525,In_1248);
or U2651 (N_2651,In_534,In_1623);
xnor U2652 (N_2652,In_1741,In_1857);
nor U2653 (N_2653,In_169,In_688);
xor U2654 (N_2654,In_1979,In_196);
or U2655 (N_2655,In_1532,In_843);
nand U2656 (N_2656,In_1524,In_1298);
nor U2657 (N_2657,In_243,In_1099);
xnor U2658 (N_2658,In_474,In_575);
xnor U2659 (N_2659,In_1250,In_549);
nor U2660 (N_2660,In_715,In_1247);
and U2661 (N_2661,In_712,In_806);
nor U2662 (N_2662,In_1528,In_1828);
nor U2663 (N_2663,In_1166,In_1240);
and U2664 (N_2664,In_1457,In_379);
nand U2665 (N_2665,In_771,In_748);
nor U2666 (N_2666,In_683,In_1532);
or U2667 (N_2667,In_1088,In_1498);
xnor U2668 (N_2668,In_265,In_1049);
nor U2669 (N_2669,In_1618,In_1966);
or U2670 (N_2670,In_205,In_705);
or U2671 (N_2671,In_699,In_385);
nor U2672 (N_2672,In_119,In_632);
nor U2673 (N_2673,In_631,In_1449);
and U2674 (N_2674,In_1227,In_1943);
nor U2675 (N_2675,In_213,In_620);
nand U2676 (N_2676,In_1824,In_266);
and U2677 (N_2677,In_1129,In_1971);
and U2678 (N_2678,In_1891,In_181);
nor U2679 (N_2679,In_381,In_1775);
or U2680 (N_2680,In_414,In_1939);
and U2681 (N_2681,In_1441,In_145);
nand U2682 (N_2682,In_826,In_1288);
nand U2683 (N_2683,In_923,In_1896);
and U2684 (N_2684,In_1349,In_348);
xnor U2685 (N_2685,In_1628,In_547);
and U2686 (N_2686,In_683,In_870);
and U2687 (N_2687,In_1075,In_356);
and U2688 (N_2688,In_434,In_1786);
and U2689 (N_2689,In_260,In_186);
xnor U2690 (N_2690,In_607,In_1304);
nand U2691 (N_2691,In_1037,In_915);
nor U2692 (N_2692,In_400,In_1012);
nand U2693 (N_2693,In_838,In_322);
nand U2694 (N_2694,In_312,In_1754);
nand U2695 (N_2695,In_943,In_886);
or U2696 (N_2696,In_1363,In_1947);
nand U2697 (N_2697,In_205,In_1588);
or U2698 (N_2698,In_1241,In_1721);
nor U2699 (N_2699,In_442,In_1321);
and U2700 (N_2700,In_965,In_864);
and U2701 (N_2701,In_552,In_632);
xnor U2702 (N_2702,In_790,In_1432);
nand U2703 (N_2703,In_868,In_626);
and U2704 (N_2704,In_1256,In_625);
or U2705 (N_2705,In_1712,In_1044);
xnor U2706 (N_2706,In_148,In_138);
nand U2707 (N_2707,In_846,In_368);
and U2708 (N_2708,In_891,In_1393);
xnor U2709 (N_2709,In_1699,In_1875);
nand U2710 (N_2710,In_1567,In_149);
or U2711 (N_2711,In_1585,In_1326);
nand U2712 (N_2712,In_1508,In_1114);
nor U2713 (N_2713,In_1978,In_427);
or U2714 (N_2714,In_72,In_1829);
nor U2715 (N_2715,In_1238,In_1222);
or U2716 (N_2716,In_638,In_1012);
nand U2717 (N_2717,In_175,In_376);
nor U2718 (N_2718,In_438,In_267);
nand U2719 (N_2719,In_1769,In_576);
and U2720 (N_2720,In_1474,In_1921);
and U2721 (N_2721,In_181,In_1638);
xor U2722 (N_2722,In_1839,In_405);
nand U2723 (N_2723,In_475,In_737);
xor U2724 (N_2724,In_1828,In_965);
or U2725 (N_2725,In_206,In_179);
or U2726 (N_2726,In_977,In_1878);
nand U2727 (N_2727,In_724,In_1943);
nand U2728 (N_2728,In_1194,In_1865);
xnor U2729 (N_2729,In_815,In_1916);
xor U2730 (N_2730,In_1449,In_1224);
or U2731 (N_2731,In_176,In_309);
or U2732 (N_2732,In_1500,In_11);
nor U2733 (N_2733,In_6,In_490);
nor U2734 (N_2734,In_600,In_1690);
nor U2735 (N_2735,In_1606,In_427);
nand U2736 (N_2736,In_1072,In_716);
and U2737 (N_2737,In_1887,In_1361);
or U2738 (N_2738,In_1948,In_1380);
nor U2739 (N_2739,In_1665,In_1982);
and U2740 (N_2740,In_269,In_1836);
nor U2741 (N_2741,In_1479,In_552);
nand U2742 (N_2742,In_341,In_1123);
and U2743 (N_2743,In_1228,In_111);
and U2744 (N_2744,In_216,In_284);
and U2745 (N_2745,In_917,In_1634);
xor U2746 (N_2746,In_1795,In_1485);
nand U2747 (N_2747,In_1914,In_1630);
nor U2748 (N_2748,In_1482,In_912);
nor U2749 (N_2749,In_818,In_480);
nor U2750 (N_2750,In_1628,In_1421);
and U2751 (N_2751,In_369,In_1456);
and U2752 (N_2752,In_1672,In_821);
nand U2753 (N_2753,In_451,In_1195);
or U2754 (N_2754,In_494,In_281);
nand U2755 (N_2755,In_1307,In_1332);
nor U2756 (N_2756,In_1813,In_941);
nor U2757 (N_2757,In_879,In_129);
nor U2758 (N_2758,In_1810,In_1229);
or U2759 (N_2759,In_1868,In_76);
or U2760 (N_2760,In_1336,In_231);
or U2761 (N_2761,In_1800,In_383);
or U2762 (N_2762,In_1242,In_893);
nand U2763 (N_2763,In_753,In_1628);
nand U2764 (N_2764,In_1329,In_1771);
nor U2765 (N_2765,In_1105,In_1223);
and U2766 (N_2766,In_1198,In_700);
nand U2767 (N_2767,In_481,In_61);
nor U2768 (N_2768,In_984,In_1113);
xnor U2769 (N_2769,In_250,In_1756);
and U2770 (N_2770,In_1019,In_1328);
or U2771 (N_2771,In_489,In_1117);
and U2772 (N_2772,In_1693,In_864);
nor U2773 (N_2773,In_868,In_1873);
or U2774 (N_2774,In_1912,In_1885);
or U2775 (N_2775,In_682,In_1304);
or U2776 (N_2776,In_629,In_14);
nor U2777 (N_2777,In_1654,In_1825);
nor U2778 (N_2778,In_697,In_1742);
nor U2779 (N_2779,In_1121,In_18);
or U2780 (N_2780,In_299,In_1723);
and U2781 (N_2781,In_1500,In_216);
xor U2782 (N_2782,In_813,In_218);
nor U2783 (N_2783,In_453,In_310);
nand U2784 (N_2784,In_1370,In_1080);
and U2785 (N_2785,In_653,In_1904);
nand U2786 (N_2786,In_427,In_900);
and U2787 (N_2787,In_1235,In_1115);
nand U2788 (N_2788,In_1109,In_1067);
and U2789 (N_2789,In_966,In_231);
nor U2790 (N_2790,In_1803,In_1326);
nand U2791 (N_2791,In_1290,In_1675);
xor U2792 (N_2792,In_698,In_660);
xnor U2793 (N_2793,In_1224,In_736);
nand U2794 (N_2794,In_1802,In_50);
or U2795 (N_2795,In_1443,In_1057);
or U2796 (N_2796,In_710,In_1320);
and U2797 (N_2797,In_966,In_1355);
and U2798 (N_2798,In_1433,In_1482);
nor U2799 (N_2799,In_529,In_1578);
nand U2800 (N_2800,In_1564,In_1140);
nor U2801 (N_2801,In_1969,In_1687);
and U2802 (N_2802,In_1297,In_965);
and U2803 (N_2803,In_1680,In_716);
nor U2804 (N_2804,In_545,In_119);
nand U2805 (N_2805,In_1487,In_846);
nand U2806 (N_2806,In_1189,In_507);
nor U2807 (N_2807,In_1692,In_112);
and U2808 (N_2808,In_581,In_20);
nand U2809 (N_2809,In_475,In_996);
nand U2810 (N_2810,In_1237,In_1531);
nand U2811 (N_2811,In_1838,In_1893);
or U2812 (N_2812,In_821,In_146);
nand U2813 (N_2813,In_178,In_573);
nor U2814 (N_2814,In_1448,In_968);
and U2815 (N_2815,In_629,In_1146);
nor U2816 (N_2816,In_765,In_592);
nand U2817 (N_2817,In_551,In_619);
nand U2818 (N_2818,In_1973,In_412);
xnor U2819 (N_2819,In_921,In_1232);
nor U2820 (N_2820,In_1277,In_1397);
and U2821 (N_2821,In_1041,In_1266);
or U2822 (N_2822,In_45,In_323);
nand U2823 (N_2823,In_887,In_190);
xnor U2824 (N_2824,In_1357,In_269);
or U2825 (N_2825,In_1093,In_1458);
and U2826 (N_2826,In_61,In_384);
nand U2827 (N_2827,In_567,In_1356);
or U2828 (N_2828,In_720,In_823);
and U2829 (N_2829,In_1232,In_583);
nor U2830 (N_2830,In_603,In_404);
or U2831 (N_2831,In_1907,In_1469);
nand U2832 (N_2832,In_1825,In_271);
nor U2833 (N_2833,In_1580,In_1732);
and U2834 (N_2834,In_1622,In_1323);
or U2835 (N_2835,In_928,In_350);
xnor U2836 (N_2836,In_324,In_1579);
or U2837 (N_2837,In_1655,In_85);
nand U2838 (N_2838,In_1104,In_837);
nand U2839 (N_2839,In_1162,In_1552);
nand U2840 (N_2840,In_1193,In_1086);
and U2841 (N_2841,In_1530,In_657);
nor U2842 (N_2842,In_595,In_859);
nor U2843 (N_2843,In_1789,In_1041);
and U2844 (N_2844,In_1663,In_1116);
and U2845 (N_2845,In_457,In_666);
and U2846 (N_2846,In_906,In_1218);
or U2847 (N_2847,In_165,In_1988);
nand U2848 (N_2848,In_1133,In_1072);
and U2849 (N_2849,In_1220,In_1330);
and U2850 (N_2850,In_943,In_1992);
and U2851 (N_2851,In_161,In_626);
or U2852 (N_2852,In_1911,In_311);
nand U2853 (N_2853,In_1384,In_1448);
or U2854 (N_2854,In_901,In_1476);
nand U2855 (N_2855,In_1821,In_1990);
or U2856 (N_2856,In_905,In_1676);
or U2857 (N_2857,In_700,In_886);
nor U2858 (N_2858,In_1158,In_1114);
and U2859 (N_2859,In_359,In_728);
and U2860 (N_2860,In_221,In_671);
nor U2861 (N_2861,In_1058,In_982);
and U2862 (N_2862,In_1966,In_829);
nand U2863 (N_2863,In_4,In_1392);
and U2864 (N_2864,In_640,In_1588);
nand U2865 (N_2865,In_793,In_1337);
or U2866 (N_2866,In_54,In_1860);
nand U2867 (N_2867,In_908,In_385);
xor U2868 (N_2868,In_401,In_1138);
or U2869 (N_2869,In_110,In_1711);
and U2870 (N_2870,In_1003,In_1131);
and U2871 (N_2871,In_1002,In_1424);
nor U2872 (N_2872,In_75,In_138);
and U2873 (N_2873,In_3,In_850);
nand U2874 (N_2874,In_1446,In_210);
nor U2875 (N_2875,In_1966,In_1538);
nor U2876 (N_2876,In_455,In_1814);
xor U2877 (N_2877,In_1828,In_499);
nor U2878 (N_2878,In_765,In_1781);
nand U2879 (N_2879,In_603,In_247);
or U2880 (N_2880,In_864,In_796);
nand U2881 (N_2881,In_864,In_1118);
nand U2882 (N_2882,In_1591,In_144);
xor U2883 (N_2883,In_492,In_1181);
or U2884 (N_2884,In_1152,In_1496);
and U2885 (N_2885,In_1174,In_1467);
and U2886 (N_2886,In_1867,In_1872);
nand U2887 (N_2887,In_408,In_1309);
and U2888 (N_2888,In_1863,In_1528);
nor U2889 (N_2889,In_1501,In_1518);
nor U2890 (N_2890,In_1644,In_1117);
xor U2891 (N_2891,In_1827,In_1207);
or U2892 (N_2892,In_1669,In_1352);
xor U2893 (N_2893,In_517,In_1852);
or U2894 (N_2894,In_1046,In_384);
nand U2895 (N_2895,In_790,In_1492);
or U2896 (N_2896,In_1996,In_1871);
nor U2897 (N_2897,In_1827,In_1873);
and U2898 (N_2898,In_1735,In_1805);
or U2899 (N_2899,In_858,In_1083);
and U2900 (N_2900,In_1441,In_1252);
nor U2901 (N_2901,In_634,In_475);
nand U2902 (N_2902,In_559,In_1214);
and U2903 (N_2903,In_1984,In_1098);
xnor U2904 (N_2904,In_537,In_935);
or U2905 (N_2905,In_249,In_1822);
nor U2906 (N_2906,In_1706,In_1758);
or U2907 (N_2907,In_615,In_718);
or U2908 (N_2908,In_1942,In_714);
or U2909 (N_2909,In_875,In_1930);
nor U2910 (N_2910,In_1087,In_1794);
nand U2911 (N_2911,In_366,In_941);
nand U2912 (N_2912,In_1159,In_164);
or U2913 (N_2913,In_932,In_1639);
nor U2914 (N_2914,In_1771,In_274);
and U2915 (N_2915,In_1334,In_1813);
or U2916 (N_2916,In_783,In_1904);
nor U2917 (N_2917,In_1531,In_388);
nor U2918 (N_2918,In_1035,In_1657);
and U2919 (N_2919,In_56,In_754);
nand U2920 (N_2920,In_503,In_261);
nor U2921 (N_2921,In_1947,In_1352);
nand U2922 (N_2922,In_1849,In_775);
nand U2923 (N_2923,In_51,In_1770);
nand U2924 (N_2924,In_165,In_709);
nor U2925 (N_2925,In_323,In_599);
nor U2926 (N_2926,In_1756,In_1764);
or U2927 (N_2927,In_1473,In_894);
and U2928 (N_2928,In_579,In_1956);
or U2929 (N_2929,In_1485,In_1196);
or U2930 (N_2930,In_170,In_404);
xnor U2931 (N_2931,In_264,In_1112);
or U2932 (N_2932,In_1140,In_717);
xor U2933 (N_2933,In_1501,In_1732);
xor U2934 (N_2934,In_626,In_369);
nor U2935 (N_2935,In_999,In_372);
and U2936 (N_2936,In_887,In_543);
or U2937 (N_2937,In_1685,In_1120);
nand U2938 (N_2938,In_6,In_68);
nor U2939 (N_2939,In_1288,In_29);
and U2940 (N_2940,In_1792,In_1073);
and U2941 (N_2941,In_513,In_1246);
or U2942 (N_2942,In_557,In_55);
nor U2943 (N_2943,In_1630,In_1106);
xor U2944 (N_2944,In_1539,In_617);
or U2945 (N_2945,In_203,In_51);
and U2946 (N_2946,In_1860,In_1666);
and U2947 (N_2947,In_1288,In_1199);
and U2948 (N_2948,In_411,In_1264);
nand U2949 (N_2949,In_1624,In_477);
nand U2950 (N_2950,In_1434,In_1944);
or U2951 (N_2951,In_1168,In_901);
nor U2952 (N_2952,In_254,In_1034);
nor U2953 (N_2953,In_970,In_1524);
xor U2954 (N_2954,In_1836,In_1419);
nand U2955 (N_2955,In_1392,In_607);
and U2956 (N_2956,In_697,In_1158);
nor U2957 (N_2957,In_1742,In_1845);
nand U2958 (N_2958,In_24,In_250);
and U2959 (N_2959,In_1129,In_53);
or U2960 (N_2960,In_70,In_465);
nor U2961 (N_2961,In_1964,In_675);
nand U2962 (N_2962,In_1077,In_1269);
nor U2963 (N_2963,In_1366,In_1539);
and U2964 (N_2964,In_299,In_1842);
xnor U2965 (N_2965,In_1796,In_1191);
nor U2966 (N_2966,In_803,In_1533);
and U2967 (N_2967,In_1321,In_1677);
xor U2968 (N_2968,In_1765,In_1281);
or U2969 (N_2969,In_1743,In_1383);
and U2970 (N_2970,In_1004,In_1905);
nor U2971 (N_2971,In_1475,In_1792);
or U2972 (N_2972,In_181,In_26);
nand U2973 (N_2973,In_496,In_708);
nand U2974 (N_2974,In_1103,In_1311);
and U2975 (N_2975,In_311,In_810);
nand U2976 (N_2976,In_1697,In_62);
or U2977 (N_2977,In_1178,In_770);
nor U2978 (N_2978,In_1884,In_541);
xor U2979 (N_2979,In_515,In_514);
nor U2980 (N_2980,In_335,In_863);
xnor U2981 (N_2981,In_1507,In_1115);
nand U2982 (N_2982,In_70,In_1007);
nor U2983 (N_2983,In_1943,In_688);
or U2984 (N_2984,In_404,In_1122);
or U2985 (N_2985,In_1752,In_55);
and U2986 (N_2986,In_1561,In_754);
nor U2987 (N_2987,In_812,In_1158);
and U2988 (N_2988,In_1041,In_557);
and U2989 (N_2989,In_1185,In_340);
nor U2990 (N_2990,In_5,In_1512);
nand U2991 (N_2991,In_1245,In_723);
nand U2992 (N_2992,In_1653,In_283);
nor U2993 (N_2993,In_1535,In_1993);
nor U2994 (N_2994,In_1415,In_259);
xnor U2995 (N_2995,In_912,In_927);
or U2996 (N_2996,In_906,In_845);
and U2997 (N_2997,In_1609,In_1979);
nand U2998 (N_2998,In_1097,In_1150);
nor U2999 (N_2999,In_385,In_1379);
and U3000 (N_3000,In_1195,In_1441);
nor U3001 (N_3001,In_714,In_665);
or U3002 (N_3002,In_1065,In_652);
or U3003 (N_3003,In_1794,In_366);
xor U3004 (N_3004,In_1889,In_1846);
or U3005 (N_3005,In_1262,In_1014);
nor U3006 (N_3006,In_177,In_424);
and U3007 (N_3007,In_635,In_1884);
nand U3008 (N_3008,In_562,In_1808);
and U3009 (N_3009,In_1328,In_917);
and U3010 (N_3010,In_470,In_684);
and U3011 (N_3011,In_1132,In_880);
nand U3012 (N_3012,In_1251,In_528);
nand U3013 (N_3013,In_747,In_952);
and U3014 (N_3014,In_957,In_1379);
nand U3015 (N_3015,In_756,In_123);
and U3016 (N_3016,In_27,In_1182);
or U3017 (N_3017,In_1253,In_375);
or U3018 (N_3018,In_1669,In_11);
and U3019 (N_3019,In_1127,In_456);
nand U3020 (N_3020,In_1127,In_1431);
and U3021 (N_3021,In_1193,In_328);
or U3022 (N_3022,In_1285,In_162);
and U3023 (N_3023,In_593,In_457);
xor U3024 (N_3024,In_1770,In_1516);
and U3025 (N_3025,In_497,In_939);
and U3026 (N_3026,In_190,In_994);
or U3027 (N_3027,In_735,In_1253);
xor U3028 (N_3028,In_47,In_1837);
nor U3029 (N_3029,In_510,In_1834);
or U3030 (N_3030,In_766,In_1865);
or U3031 (N_3031,In_124,In_1940);
or U3032 (N_3032,In_126,In_608);
nand U3033 (N_3033,In_665,In_1937);
nor U3034 (N_3034,In_885,In_1672);
nor U3035 (N_3035,In_1202,In_804);
and U3036 (N_3036,In_40,In_285);
nor U3037 (N_3037,In_1361,In_1592);
or U3038 (N_3038,In_1019,In_1251);
nor U3039 (N_3039,In_217,In_1396);
nor U3040 (N_3040,In_1153,In_1633);
nand U3041 (N_3041,In_1462,In_1953);
and U3042 (N_3042,In_1705,In_1710);
nand U3043 (N_3043,In_432,In_1044);
xnor U3044 (N_3044,In_877,In_641);
nor U3045 (N_3045,In_11,In_1553);
or U3046 (N_3046,In_2,In_939);
nand U3047 (N_3047,In_465,In_191);
or U3048 (N_3048,In_956,In_410);
xnor U3049 (N_3049,In_290,In_1670);
and U3050 (N_3050,In_1317,In_633);
nor U3051 (N_3051,In_297,In_1016);
xnor U3052 (N_3052,In_882,In_334);
xor U3053 (N_3053,In_871,In_246);
nand U3054 (N_3054,In_456,In_1389);
xor U3055 (N_3055,In_1769,In_497);
nor U3056 (N_3056,In_970,In_12);
and U3057 (N_3057,In_336,In_1817);
nand U3058 (N_3058,In_783,In_122);
nand U3059 (N_3059,In_29,In_24);
or U3060 (N_3060,In_708,In_486);
nor U3061 (N_3061,In_441,In_772);
nor U3062 (N_3062,In_412,In_1084);
and U3063 (N_3063,In_409,In_474);
or U3064 (N_3064,In_773,In_982);
xnor U3065 (N_3065,In_752,In_837);
and U3066 (N_3066,In_1088,In_338);
nand U3067 (N_3067,In_1604,In_1509);
or U3068 (N_3068,In_78,In_1590);
xnor U3069 (N_3069,In_821,In_794);
nand U3070 (N_3070,In_1688,In_1116);
nor U3071 (N_3071,In_1906,In_619);
or U3072 (N_3072,In_202,In_982);
or U3073 (N_3073,In_1004,In_128);
and U3074 (N_3074,In_1091,In_1105);
nand U3075 (N_3075,In_137,In_47);
nor U3076 (N_3076,In_1689,In_1742);
and U3077 (N_3077,In_267,In_1292);
and U3078 (N_3078,In_1082,In_644);
or U3079 (N_3079,In_1633,In_1899);
or U3080 (N_3080,In_277,In_145);
and U3081 (N_3081,In_630,In_1671);
and U3082 (N_3082,In_1459,In_1293);
nand U3083 (N_3083,In_555,In_1543);
or U3084 (N_3084,In_1311,In_834);
and U3085 (N_3085,In_988,In_1717);
nand U3086 (N_3086,In_1980,In_712);
nor U3087 (N_3087,In_1192,In_377);
and U3088 (N_3088,In_364,In_422);
and U3089 (N_3089,In_1877,In_37);
nand U3090 (N_3090,In_1629,In_1709);
nand U3091 (N_3091,In_1920,In_1886);
nor U3092 (N_3092,In_1240,In_515);
xnor U3093 (N_3093,In_1147,In_1731);
nor U3094 (N_3094,In_916,In_1439);
nor U3095 (N_3095,In_1965,In_337);
nand U3096 (N_3096,In_1634,In_771);
xnor U3097 (N_3097,In_1997,In_1895);
or U3098 (N_3098,In_741,In_1993);
and U3099 (N_3099,In_920,In_426);
or U3100 (N_3100,In_144,In_1618);
nand U3101 (N_3101,In_1022,In_1223);
or U3102 (N_3102,In_224,In_1665);
or U3103 (N_3103,In_626,In_1774);
or U3104 (N_3104,In_536,In_753);
or U3105 (N_3105,In_1851,In_1458);
or U3106 (N_3106,In_275,In_453);
and U3107 (N_3107,In_1836,In_59);
nor U3108 (N_3108,In_930,In_1718);
or U3109 (N_3109,In_292,In_329);
or U3110 (N_3110,In_731,In_654);
nor U3111 (N_3111,In_1809,In_847);
or U3112 (N_3112,In_1446,In_1575);
and U3113 (N_3113,In_411,In_1335);
nand U3114 (N_3114,In_1318,In_97);
and U3115 (N_3115,In_457,In_1132);
and U3116 (N_3116,In_1116,In_657);
and U3117 (N_3117,In_1167,In_775);
or U3118 (N_3118,In_143,In_1069);
nand U3119 (N_3119,In_821,In_1577);
xnor U3120 (N_3120,In_1957,In_581);
and U3121 (N_3121,In_359,In_384);
and U3122 (N_3122,In_1850,In_1416);
nor U3123 (N_3123,In_804,In_1356);
nor U3124 (N_3124,In_697,In_280);
and U3125 (N_3125,In_986,In_16);
and U3126 (N_3126,In_1137,In_1247);
nand U3127 (N_3127,In_1521,In_231);
and U3128 (N_3128,In_9,In_889);
and U3129 (N_3129,In_1201,In_1260);
or U3130 (N_3130,In_1915,In_369);
xor U3131 (N_3131,In_522,In_314);
nor U3132 (N_3132,In_590,In_1773);
or U3133 (N_3133,In_1742,In_1160);
or U3134 (N_3134,In_811,In_790);
and U3135 (N_3135,In_76,In_1818);
nor U3136 (N_3136,In_1599,In_1202);
nor U3137 (N_3137,In_403,In_1764);
or U3138 (N_3138,In_483,In_980);
nor U3139 (N_3139,In_1850,In_64);
nor U3140 (N_3140,In_27,In_815);
nor U3141 (N_3141,In_135,In_292);
xor U3142 (N_3142,In_534,In_595);
or U3143 (N_3143,In_1467,In_1432);
nor U3144 (N_3144,In_737,In_415);
nor U3145 (N_3145,In_298,In_1506);
nand U3146 (N_3146,In_263,In_1811);
or U3147 (N_3147,In_735,In_1152);
or U3148 (N_3148,In_1376,In_1216);
and U3149 (N_3149,In_470,In_1450);
and U3150 (N_3150,In_1760,In_1287);
or U3151 (N_3151,In_41,In_1196);
nand U3152 (N_3152,In_1269,In_1578);
nor U3153 (N_3153,In_1264,In_56);
or U3154 (N_3154,In_1459,In_1538);
and U3155 (N_3155,In_1951,In_1767);
nor U3156 (N_3156,In_1586,In_1867);
nor U3157 (N_3157,In_331,In_413);
nand U3158 (N_3158,In_1364,In_909);
nor U3159 (N_3159,In_243,In_368);
nand U3160 (N_3160,In_1233,In_470);
or U3161 (N_3161,In_1489,In_1234);
and U3162 (N_3162,In_685,In_1826);
nand U3163 (N_3163,In_411,In_890);
and U3164 (N_3164,In_309,In_1489);
nor U3165 (N_3165,In_930,In_1207);
nand U3166 (N_3166,In_1214,In_763);
nand U3167 (N_3167,In_757,In_476);
nand U3168 (N_3168,In_1164,In_1377);
and U3169 (N_3169,In_1226,In_1862);
or U3170 (N_3170,In_137,In_1222);
nor U3171 (N_3171,In_597,In_1948);
nand U3172 (N_3172,In_1926,In_339);
nand U3173 (N_3173,In_1872,In_413);
or U3174 (N_3174,In_1481,In_290);
nand U3175 (N_3175,In_1691,In_1481);
or U3176 (N_3176,In_1816,In_1510);
nor U3177 (N_3177,In_293,In_720);
nor U3178 (N_3178,In_1407,In_1966);
and U3179 (N_3179,In_1499,In_281);
and U3180 (N_3180,In_1174,In_1943);
nand U3181 (N_3181,In_1692,In_1839);
or U3182 (N_3182,In_637,In_1080);
nor U3183 (N_3183,In_693,In_1486);
xnor U3184 (N_3184,In_44,In_1137);
nand U3185 (N_3185,In_1521,In_1627);
and U3186 (N_3186,In_907,In_1368);
or U3187 (N_3187,In_1845,In_726);
nor U3188 (N_3188,In_1310,In_1142);
nand U3189 (N_3189,In_1135,In_825);
nand U3190 (N_3190,In_45,In_623);
xnor U3191 (N_3191,In_1685,In_1578);
nand U3192 (N_3192,In_870,In_1341);
or U3193 (N_3193,In_1919,In_1653);
or U3194 (N_3194,In_451,In_832);
nand U3195 (N_3195,In_1235,In_680);
xor U3196 (N_3196,In_588,In_767);
nand U3197 (N_3197,In_1633,In_1802);
nor U3198 (N_3198,In_139,In_0);
nor U3199 (N_3199,In_1506,In_550);
nor U3200 (N_3200,In_98,In_1860);
xnor U3201 (N_3201,In_526,In_318);
or U3202 (N_3202,In_668,In_1766);
and U3203 (N_3203,In_1107,In_606);
or U3204 (N_3204,In_1548,In_486);
nand U3205 (N_3205,In_1580,In_1622);
and U3206 (N_3206,In_1544,In_1072);
and U3207 (N_3207,In_591,In_631);
or U3208 (N_3208,In_934,In_469);
and U3209 (N_3209,In_578,In_1640);
or U3210 (N_3210,In_252,In_1464);
and U3211 (N_3211,In_270,In_1860);
and U3212 (N_3212,In_170,In_1407);
xnor U3213 (N_3213,In_1752,In_1663);
nor U3214 (N_3214,In_686,In_1102);
nand U3215 (N_3215,In_1164,In_58);
or U3216 (N_3216,In_1060,In_751);
or U3217 (N_3217,In_705,In_857);
nor U3218 (N_3218,In_308,In_773);
nor U3219 (N_3219,In_1700,In_1372);
nor U3220 (N_3220,In_181,In_976);
nand U3221 (N_3221,In_1591,In_228);
xor U3222 (N_3222,In_1351,In_1985);
nor U3223 (N_3223,In_1821,In_1452);
or U3224 (N_3224,In_317,In_1376);
and U3225 (N_3225,In_492,In_1775);
or U3226 (N_3226,In_1755,In_1157);
or U3227 (N_3227,In_1346,In_36);
nand U3228 (N_3228,In_1729,In_112);
and U3229 (N_3229,In_26,In_714);
xor U3230 (N_3230,In_406,In_245);
nand U3231 (N_3231,In_1140,In_1093);
nand U3232 (N_3232,In_1099,In_131);
or U3233 (N_3233,In_1704,In_1441);
and U3234 (N_3234,In_1493,In_1925);
xnor U3235 (N_3235,In_828,In_1553);
or U3236 (N_3236,In_650,In_1504);
xnor U3237 (N_3237,In_53,In_1375);
nor U3238 (N_3238,In_1615,In_1468);
nor U3239 (N_3239,In_1669,In_1095);
nand U3240 (N_3240,In_14,In_1903);
and U3241 (N_3241,In_961,In_751);
nor U3242 (N_3242,In_1382,In_1980);
nand U3243 (N_3243,In_515,In_162);
xor U3244 (N_3244,In_995,In_912);
xnor U3245 (N_3245,In_370,In_1889);
nor U3246 (N_3246,In_1319,In_566);
or U3247 (N_3247,In_1136,In_526);
or U3248 (N_3248,In_388,In_1049);
or U3249 (N_3249,In_264,In_590);
nand U3250 (N_3250,In_209,In_630);
or U3251 (N_3251,In_1818,In_1530);
or U3252 (N_3252,In_599,In_760);
nand U3253 (N_3253,In_363,In_1917);
nor U3254 (N_3254,In_629,In_455);
nand U3255 (N_3255,In_1933,In_687);
nor U3256 (N_3256,In_870,In_1056);
and U3257 (N_3257,In_913,In_288);
and U3258 (N_3258,In_438,In_1459);
nor U3259 (N_3259,In_1803,In_1562);
nand U3260 (N_3260,In_1142,In_557);
or U3261 (N_3261,In_370,In_991);
nor U3262 (N_3262,In_977,In_1824);
nand U3263 (N_3263,In_1015,In_795);
or U3264 (N_3264,In_1622,In_1179);
nor U3265 (N_3265,In_804,In_253);
and U3266 (N_3266,In_570,In_1893);
nor U3267 (N_3267,In_1301,In_1471);
xnor U3268 (N_3268,In_1598,In_128);
xor U3269 (N_3269,In_1771,In_1864);
nor U3270 (N_3270,In_1107,In_507);
nor U3271 (N_3271,In_406,In_1293);
nand U3272 (N_3272,In_1434,In_875);
or U3273 (N_3273,In_1046,In_109);
or U3274 (N_3274,In_861,In_1215);
nor U3275 (N_3275,In_1729,In_547);
and U3276 (N_3276,In_1552,In_692);
nand U3277 (N_3277,In_1862,In_399);
nor U3278 (N_3278,In_904,In_1631);
and U3279 (N_3279,In_1672,In_725);
nand U3280 (N_3280,In_1703,In_1655);
and U3281 (N_3281,In_1501,In_778);
xnor U3282 (N_3282,In_111,In_103);
xor U3283 (N_3283,In_1455,In_1275);
nand U3284 (N_3284,In_189,In_1176);
or U3285 (N_3285,In_142,In_1682);
nand U3286 (N_3286,In_1300,In_261);
nand U3287 (N_3287,In_1944,In_349);
nor U3288 (N_3288,In_863,In_1565);
xnor U3289 (N_3289,In_1664,In_410);
nor U3290 (N_3290,In_1747,In_855);
nand U3291 (N_3291,In_1422,In_1979);
and U3292 (N_3292,In_929,In_1994);
nor U3293 (N_3293,In_1794,In_952);
xnor U3294 (N_3294,In_1177,In_837);
nand U3295 (N_3295,In_702,In_357);
and U3296 (N_3296,In_489,In_370);
and U3297 (N_3297,In_1558,In_687);
nand U3298 (N_3298,In_489,In_954);
nor U3299 (N_3299,In_258,In_1213);
nor U3300 (N_3300,In_1334,In_1623);
and U3301 (N_3301,In_1160,In_364);
or U3302 (N_3302,In_242,In_56);
or U3303 (N_3303,In_1760,In_1001);
or U3304 (N_3304,In_1235,In_1964);
or U3305 (N_3305,In_1947,In_242);
nor U3306 (N_3306,In_638,In_1459);
or U3307 (N_3307,In_1218,In_588);
and U3308 (N_3308,In_1944,In_1075);
nor U3309 (N_3309,In_940,In_1395);
or U3310 (N_3310,In_499,In_1165);
nor U3311 (N_3311,In_692,In_502);
and U3312 (N_3312,In_1934,In_117);
or U3313 (N_3313,In_310,In_135);
and U3314 (N_3314,In_436,In_716);
or U3315 (N_3315,In_1070,In_1238);
xnor U3316 (N_3316,In_775,In_779);
nor U3317 (N_3317,In_1305,In_73);
nor U3318 (N_3318,In_926,In_170);
nand U3319 (N_3319,In_905,In_922);
nor U3320 (N_3320,In_1600,In_1114);
nor U3321 (N_3321,In_1213,In_1271);
or U3322 (N_3322,In_1207,In_1948);
and U3323 (N_3323,In_265,In_1453);
nand U3324 (N_3324,In_177,In_1014);
and U3325 (N_3325,In_1518,In_437);
and U3326 (N_3326,In_511,In_901);
nor U3327 (N_3327,In_44,In_1873);
xor U3328 (N_3328,In_875,In_855);
nor U3329 (N_3329,In_846,In_504);
nor U3330 (N_3330,In_668,In_132);
and U3331 (N_3331,In_1063,In_270);
or U3332 (N_3332,In_1111,In_753);
and U3333 (N_3333,In_1878,In_1979);
nor U3334 (N_3334,In_1170,In_683);
nor U3335 (N_3335,In_684,In_1706);
nand U3336 (N_3336,In_1060,In_970);
and U3337 (N_3337,In_187,In_259);
and U3338 (N_3338,In_833,In_1724);
nor U3339 (N_3339,In_1432,In_1700);
and U3340 (N_3340,In_1762,In_120);
nand U3341 (N_3341,In_745,In_224);
nor U3342 (N_3342,In_1451,In_45);
xnor U3343 (N_3343,In_112,In_689);
and U3344 (N_3344,In_1830,In_1615);
nor U3345 (N_3345,In_1106,In_1244);
and U3346 (N_3346,In_1039,In_1087);
or U3347 (N_3347,In_544,In_1046);
or U3348 (N_3348,In_398,In_1579);
nor U3349 (N_3349,In_1789,In_1422);
and U3350 (N_3350,In_1456,In_716);
or U3351 (N_3351,In_550,In_764);
and U3352 (N_3352,In_1915,In_210);
or U3353 (N_3353,In_80,In_1534);
nand U3354 (N_3354,In_1455,In_112);
nand U3355 (N_3355,In_791,In_9);
nand U3356 (N_3356,In_1622,In_1277);
and U3357 (N_3357,In_710,In_1141);
nor U3358 (N_3358,In_764,In_1663);
nand U3359 (N_3359,In_81,In_161);
or U3360 (N_3360,In_163,In_900);
nand U3361 (N_3361,In_455,In_484);
and U3362 (N_3362,In_1497,In_1061);
or U3363 (N_3363,In_240,In_555);
and U3364 (N_3364,In_1492,In_1904);
nor U3365 (N_3365,In_1173,In_113);
or U3366 (N_3366,In_398,In_471);
nand U3367 (N_3367,In_1553,In_162);
or U3368 (N_3368,In_1500,In_933);
and U3369 (N_3369,In_1567,In_551);
or U3370 (N_3370,In_616,In_1540);
nor U3371 (N_3371,In_21,In_894);
nor U3372 (N_3372,In_699,In_192);
nor U3373 (N_3373,In_801,In_61);
xnor U3374 (N_3374,In_1736,In_307);
nor U3375 (N_3375,In_355,In_1054);
and U3376 (N_3376,In_288,In_1835);
xor U3377 (N_3377,In_136,In_1052);
or U3378 (N_3378,In_153,In_956);
nor U3379 (N_3379,In_1517,In_943);
and U3380 (N_3380,In_1195,In_1543);
or U3381 (N_3381,In_89,In_216);
nor U3382 (N_3382,In_520,In_1055);
nor U3383 (N_3383,In_1802,In_635);
nand U3384 (N_3384,In_1329,In_587);
xor U3385 (N_3385,In_1840,In_1444);
nor U3386 (N_3386,In_589,In_1028);
xor U3387 (N_3387,In_208,In_777);
nand U3388 (N_3388,In_1792,In_1939);
or U3389 (N_3389,In_783,In_229);
nand U3390 (N_3390,In_946,In_475);
or U3391 (N_3391,In_1447,In_488);
or U3392 (N_3392,In_1045,In_467);
and U3393 (N_3393,In_1494,In_692);
nand U3394 (N_3394,In_1609,In_1362);
nand U3395 (N_3395,In_553,In_1580);
nand U3396 (N_3396,In_1505,In_1212);
nor U3397 (N_3397,In_418,In_1620);
or U3398 (N_3398,In_1491,In_698);
and U3399 (N_3399,In_1278,In_1654);
nand U3400 (N_3400,In_1377,In_1828);
and U3401 (N_3401,In_1054,In_915);
or U3402 (N_3402,In_438,In_200);
xor U3403 (N_3403,In_1916,In_217);
or U3404 (N_3404,In_865,In_1504);
and U3405 (N_3405,In_1228,In_485);
nand U3406 (N_3406,In_1719,In_448);
xor U3407 (N_3407,In_508,In_1322);
nand U3408 (N_3408,In_840,In_1741);
nor U3409 (N_3409,In_1877,In_1519);
or U3410 (N_3410,In_1552,In_512);
nand U3411 (N_3411,In_1664,In_1022);
xor U3412 (N_3412,In_861,In_1218);
nor U3413 (N_3413,In_655,In_1047);
and U3414 (N_3414,In_342,In_862);
nand U3415 (N_3415,In_1932,In_978);
nor U3416 (N_3416,In_1583,In_733);
nand U3417 (N_3417,In_1474,In_1091);
or U3418 (N_3418,In_525,In_1073);
and U3419 (N_3419,In_722,In_1952);
and U3420 (N_3420,In_361,In_308);
or U3421 (N_3421,In_615,In_733);
and U3422 (N_3422,In_591,In_600);
and U3423 (N_3423,In_411,In_669);
nor U3424 (N_3424,In_998,In_726);
and U3425 (N_3425,In_572,In_1800);
and U3426 (N_3426,In_938,In_1078);
nand U3427 (N_3427,In_570,In_1741);
and U3428 (N_3428,In_394,In_1789);
and U3429 (N_3429,In_443,In_1624);
or U3430 (N_3430,In_1709,In_808);
or U3431 (N_3431,In_766,In_985);
nand U3432 (N_3432,In_1713,In_621);
and U3433 (N_3433,In_991,In_1726);
nor U3434 (N_3434,In_739,In_718);
nor U3435 (N_3435,In_1072,In_1553);
xor U3436 (N_3436,In_1918,In_1086);
xor U3437 (N_3437,In_1089,In_595);
or U3438 (N_3438,In_1363,In_1497);
or U3439 (N_3439,In_1068,In_347);
xnor U3440 (N_3440,In_897,In_601);
nand U3441 (N_3441,In_859,In_664);
or U3442 (N_3442,In_1177,In_1590);
and U3443 (N_3443,In_715,In_373);
and U3444 (N_3444,In_1037,In_440);
nand U3445 (N_3445,In_852,In_1663);
and U3446 (N_3446,In_403,In_49);
and U3447 (N_3447,In_1944,In_489);
and U3448 (N_3448,In_194,In_138);
nand U3449 (N_3449,In_1152,In_1678);
xnor U3450 (N_3450,In_324,In_1691);
nor U3451 (N_3451,In_416,In_1001);
nor U3452 (N_3452,In_395,In_567);
or U3453 (N_3453,In_1916,In_1676);
and U3454 (N_3454,In_1344,In_115);
or U3455 (N_3455,In_729,In_1446);
and U3456 (N_3456,In_713,In_1726);
or U3457 (N_3457,In_832,In_660);
nand U3458 (N_3458,In_734,In_1);
and U3459 (N_3459,In_1301,In_1734);
and U3460 (N_3460,In_170,In_893);
and U3461 (N_3461,In_1838,In_605);
nor U3462 (N_3462,In_416,In_580);
nor U3463 (N_3463,In_594,In_1781);
xor U3464 (N_3464,In_1160,In_1156);
nand U3465 (N_3465,In_1335,In_547);
nor U3466 (N_3466,In_465,In_722);
nand U3467 (N_3467,In_572,In_1170);
and U3468 (N_3468,In_1842,In_487);
and U3469 (N_3469,In_1746,In_341);
or U3470 (N_3470,In_788,In_215);
or U3471 (N_3471,In_1049,In_1175);
nand U3472 (N_3472,In_1551,In_1667);
or U3473 (N_3473,In_1420,In_34);
nand U3474 (N_3474,In_595,In_816);
nor U3475 (N_3475,In_882,In_412);
nor U3476 (N_3476,In_798,In_416);
or U3477 (N_3477,In_1092,In_1396);
nor U3478 (N_3478,In_1309,In_1247);
or U3479 (N_3479,In_832,In_223);
and U3480 (N_3480,In_1190,In_92);
nand U3481 (N_3481,In_634,In_1638);
nor U3482 (N_3482,In_1045,In_1183);
nor U3483 (N_3483,In_551,In_540);
nand U3484 (N_3484,In_1644,In_703);
or U3485 (N_3485,In_965,In_1661);
and U3486 (N_3486,In_95,In_299);
nor U3487 (N_3487,In_1472,In_1498);
or U3488 (N_3488,In_241,In_1085);
and U3489 (N_3489,In_926,In_1045);
or U3490 (N_3490,In_1126,In_703);
and U3491 (N_3491,In_1242,In_1703);
nor U3492 (N_3492,In_1546,In_1038);
and U3493 (N_3493,In_38,In_1515);
nand U3494 (N_3494,In_392,In_966);
or U3495 (N_3495,In_1796,In_1443);
and U3496 (N_3496,In_66,In_1650);
and U3497 (N_3497,In_1902,In_62);
and U3498 (N_3498,In_630,In_572);
nand U3499 (N_3499,In_802,In_1460);
nand U3500 (N_3500,In_1128,In_1791);
nor U3501 (N_3501,In_673,In_698);
or U3502 (N_3502,In_1069,In_43);
nor U3503 (N_3503,In_987,In_1860);
xnor U3504 (N_3504,In_30,In_1952);
or U3505 (N_3505,In_1428,In_258);
or U3506 (N_3506,In_1728,In_104);
xor U3507 (N_3507,In_141,In_1599);
nand U3508 (N_3508,In_1113,In_359);
or U3509 (N_3509,In_119,In_509);
and U3510 (N_3510,In_1702,In_58);
nand U3511 (N_3511,In_1541,In_714);
and U3512 (N_3512,In_156,In_150);
or U3513 (N_3513,In_1600,In_853);
nor U3514 (N_3514,In_597,In_672);
nor U3515 (N_3515,In_1290,In_1953);
nand U3516 (N_3516,In_969,In_1711);
or U3517 (N_3517,In_657,In_168);
nor U3518 (N_3518,In_1311,In_98);
or U3519 (N_3519,In_1528,In_909);
and U3520 (N_3520,In_1514,In_1926);
nor U3521 (N_3521,In_452,In_38);
xnor U3522 (N_3522,In_59,In_887);
nand U3523 (N_3523,In_670,In_977);
xor U3524 (N_3524,In_83,In_455);
and U3525 (N_3525,In_339,In_969);
nor U3526 (N_3526,In_1111,In_12);
and U3527 (N_3527,In_1361,In_1012);
nor U3528 (N_3528,In_78,In_1399);
and U3529 (N_3529,In_430,In_1460);
nand U3530 (N_3530,In_1311,In_1791);
nand U3531 (N_3531,In_881,In_753);
and U3532 (N_3532,In_736,In_1389);
nand U3533 (N_3533,In_1098,In_1016);
or U3534 (N_3534,In_1280,In_242);
and U3535 (N_3535,In_446,In_713);
or U3536 (N_3536,In_1830,In_1461);
xor U3537 (N_3537,In_1752,In_844);
or U3538 (N_3538,In_301,In_1797);
nand U3539 (N_3539,In_1469,In_1259);
and U3540 (N_3540,In_1490,In_1227);
nor U3541 (N_3541,In_1146,In_1841);
or U3542 (N_3542,In_1921,In_352);
nand U3543 (N_3543,In_1834,In_1178);
or U3544 (N_3544,In_423,In_1740);
xnor U3545 (N_3545,In_382,In_1377);
nor U3546 (N_3546,In_196,In_261);
or U3547 (N_3547,In_723,In_1677);
and U3548 (N_3548,In_1909,In_1351);
nor U3549 (N_3549,In_147,In_933);
and U3550 (N_3550,In_1161,In_480);
nor U3551 (N_3551,In_1672,In_1766);
or U3552 (N_3552,In_1744,In_3);
or U3553 (N_3553,In_1084,In_1192);
nor U3554 (N_3554,In_197,In_127);
or U3555 (N_3555,In_1364,In_175);
nand U3556 (N_3556,In_116,In_62);
xnor U3557 (N_3557,In_125,In_686);
nor U3558 (N_3558,In_326,In_1677);
or U3559 (N_3559,In_1708,In_1071);
or U3560 (N_3560,In_116,In_1719);
nor U3561 (N_3561,In_1545,In_1436);
or U3562 (N_3562,In_1086,In_949);
and U3563 (N_3563,In_1046,In_1451);
or U3564 (N_3564,In_1736,In_665);
xnor U3565 (N_3565,In_569,In_1070);
xnor U3566 (N_3566,In_1756,In_916);
or U3567 (N_3567,In_1332,In_1321);
nor U3568 (N_3568,In_1314,In_1213);
and U3569 (N_3569,In_1795,In_916);
or U3570 (N_3570,In_452,In_1152);
and U3571 (N_3571,In_762,In_731);
or U3572 (N_3572,In_1924,In_1726);
nand U3573 (N_3573,In_586,In_1458);
nor U3574 (N_3574,In_503,In_1653);
and U3575 (N_3575,In_1867,In_196);
nor U3576 (N_3576,In_1917,In_1446);
or U3577 (N_3577,In_1691,In_669);
nand U3578 (N_3578,In_208,In_674);
nor U3579 (N_3579,In_933,In_1266);
nand U3580 (N_3580,In_851,In_686);
or U3581 (N_3581,In_1658,In_74);
or U3582 (N_3582,In_425,In_1885);
and U3583 (N_3583,In_1217,In_534);
and U3584 (N_3584,In_1759,In_169);
and U3585 (N_3585,In_1070,In_883);
nand U3586 (N_3586,In_1406,In_0);
nand U3587 (N_3587,In_1593,In_538);
or U3588 (N_3588,In_1190,In_987);
and U3589 (N_3589,In_1420,In_1004);
nand U3590 (N_3590,In_1462,In_223);
nor U3591 (N_3591,In_1442,In_1728);
and U3592 (N_3592,In_1791,In_1340);
and U3593 (N_3593,In_1408,In_1713);
xnor U3594 (N_3594,In_418,In_1828);
and U3595 (N_3595,In_1236,In_1694);
nor U3596 (N_3596,In_1093,In_422);
or U3597 (N_3597,In_878,In_1787);
and U3598 (N_3598,In_327,In_494);
nand U3599 (N_3599,In_1831,In_1954);
nor U3600 (N_3600,In_536,In_612);
nand U3601 (N_3601,In_280,In_1229);
nor U3602 (N_3602,In_685,In_151);
and U3603 (N_3603,In_1606,In_1983);
or U3604 (N_3604,In_417,In_915);
nor U3605 (N_3605,In_275,In_918);
and U3606 (N_3606,In_986,In_1276);
nand U3607 (N_3607,In_289,In_1528);
or U3608 (N_3608,In_192,In_1325);
nor U3609 (N_3609,In_1234,In_1292);
nor U3610 (N_3610,In_1727,In_1685);
and U3611 (N_3611,In_1583,In_13);
nand U3612 (N_3612,In_1184,In_11);
and U3613 (N_3613,In_1760,In_1660);
and U3614 (N_3614,In_527,In_1008);
and U3615 (N_3615,In_1463,In_1195);
and U3616 (N_3616,In_158,In_546);
and U3617 (N_3617,In_861,In_1060);
nand U3618 (N_3618,In_213,In_1704);
and U3619 (N_3619,In_475,In_133);
nor U3620 (N_3620,In_1027,In_1264);
and U3621 (N_3621,In_934,In_511);
or U3622 (N_3622,In_203,In_1589);
nand U3623 (N_3623,In_2,In_1889);
or U3624 (N_3624,In_196,In_675);
or U3625 (N_3625,In_1972,In_605);
or U3626 (N_3626,In_690,In_1971);
nand U3627 (N_3627,In_969,In_1296);
or U3628 (N_3628,In_1814,In_643);
nor U3629 (N_3629,In_1063,In_626);
xor U3630 (N_3630,In_800,In_1626);
and U3631 (N_3631,In_1838,In_1432);
nand U3632 (N_3632,In_1881,In_1833);
or U3633 (N_3633,In_1845,In_1112);
nand U3634 (N_3634,In_478,In_114);
nand U3635 (N_3635,In_59,In_1584);
and U3636 (N_3636,In_1055,In_329);
and U3637 (N_3637,In_421,In_1030);
or U3638 (N_3638,In_1939,In_7);
nand U3639 (N_3639,In_621,In_1812);
nor U3640 (N_3640,In_1310,In_479);
nor U3641 (N_3641,In_1439,In_1249);
and U3642 (N_3642,In_94,In_1957);
or U3643 (N_3643,In_452,In_903);
xor U3644 (N_3644,In_268,In_324);
nor U3645 (N_3645,In_755,In_263);
or U3646 (N_3646,In_151,In_176);
nand U3647 (N_3647,In_1905,In_778);
nand U3648 (N_3648,In_1753,In_90);
or U3649 (N_3649,In_1787,In_805);
nand U3650 (N_3650,In_1640,In_1747);
nor U3651 (N_3651,In_1172,In_1402);
or U3652 (N_3652,In_542,In_252);
xnor U3653 (N_3653,In_1528,In_306);
or U3654 (N_3654,In_675,In_1978);
or U3655 (N_3655,In_1624,In_1110);
nand U3656 (N_3656,In_86,In_71);
nand U3657 (N_3657,In_1836,In_1167);
nand U3658 (N_3658,In_491,In_1823);
or U3659 (N_3659,In_127,In_205);
or U3660 (N_3660,In_1456,In_1981);
xor U3661 (N_3661,In_994,In_198);
nor U3662 (N_3662,In_983,In_89);
nand U3663 (N_3663,In_930,In_946);
or U3664 (N_3664,In_1843,In_1835);
and U3665 (N_3665,In_1035,In_699);
or U3666 (N_3666,In_436,In_1608);
nor U3667 (N_3667,In_361,In_1252);
nand U3668 (N_3668,In_1403,In_1480);
xor U3669 (N_3669,In_790,In_1220);
xor U3670 (N_3670,In_385,In_367);
nand U3671 (N_3671,In_1901,In_940);
nand U3672 (N_3672,In_1502,In_1697);
nand U3673 (N_3673,In_1417,In_1502);
and U3674 (N_3674,In_751,In_786);
nor U3675 (N_3675,In_1054,In_1684);
nand U3676 (N_3676,In_1031,In_1919);
nor U3677 (N_3677,In_176,In_945);
nand U3678 (N_3678,In_1063,In_915);
and U3679 (N_3679,In_768,In_917);
nor U3680 (N_3680,In_583,In_944);
xor U3681 (N_3681,In_1772,In_1217);
or U3682 (N_3682,In_188,In_140);
nand U3683 (N_3683,In_694,In_1871);
and U3684 (N_3684,In_129,In_1488);
or U3685 (N_3685,In_667,In_603);
nand U3686 (N_3686,In_630,In_112);
xor U3687 (N_3687,In_504,In_420);
nand U3688 (N_3688,In_7,In_2);
nand U3689 (N_3689,In_1802,In_1295);
nand U3690 (N_3690,In_813,In_993);
nand U3691 (N_3691,In_771,In_1906);
nand U3692 (N_3692,In_1257,In_1580);
nor U3693 (N_3693,In_306,In_1403);
or U3694 (N_3694,In_835,In_1216);
nand U3695 (N_3695,In_905,In_374);
nand U3696 (N_3696,In_1377,In_57);
nand U3697 (N_3697,In_1045,In_1694);
and U3698 (N_3698,In_952,In_690);
or U3699 (N_3699,In_1008,In_1941);
or U3700 (N_3700,In_833,In_873);
nand U3701 (N_3701,In_308,In_542);
or U3702 (N_3702,In_190,In_1442);
nand U3703 (N_3703,In_1123,In_1281);
nand U3704 (N_3704,In_877,In_1271);
and U3705 (N_3705,In_282,In_1868);
or U3706 (N_3706,In_936,In_191);
and U3707 (N_3707,In_1580,In_1037);
nand U3708 (N_3708,In_64,In_1426);
and U3709 (N_3709,In_701,In_1529);
nand U3710 (N_3710,In_1950,In_1306);
or U3711 (N_3711,In_1325,In_1478);
xor U3712 (N_3712,In_75,In_303);
or U3713 (N_3713,In_1713,In_1990);
and U3714 (N_3714,In_878,In_1529);
nand U3715 (N_3715,In_1221,In_1603);
and U3716 (N_3716,In_1708,In_1565);
or U3717 (N_3717,In_551,In_382);
nor U3718 (N_3718,In_612,In_1956);
nor U3719 (N_3719,In_1252,In_944);
and U3720 (N_3720,In_104,In_444);
nor U3721 (N_3721,In_990,In_1864);
nor U3722 (N_3722,In_1651,In_932);
or U3723 (N_3723,In_1928,In_19);
nor U3724 (N_3724,In_1308,In_95);
or U3725 (N_3725,In_1121,In_289);
nor U3726 (N_3726,In_234,In_1962);
or U3727 (N_3727,In_1117,In_766);
xor U3728 (N_3728,In_1026,In_925);
or U3729 (N_3729,In_50,In_777);
nor U3730 (N_3730,In_1949,In_1959);
nor U3731 (N_3731,In_945,In_5);
nand U3732 (N_3732,In_167,In_1046);
and U3733 (N_3733,In_214,In_1534);
nor U3734 (N_3734,In_794,In_1805);
nand U3735 (N_3735,In_1830,In_521);
nand U3736 (N_3736,In_1618,In_254);
or U3737 (N_3737,In_1568,In_1215);
or U3738 (N_3738,In_268,In_259);
and U3739 (N_3739,In_992,In_789);
nand U3740 (N_3740,In_418,In_877);
nand U3741 (N_3741,In_985,In_729);
nand U3742 (N_3742,In_1269,In_1338);
or U3743 (N_3743,In_1921,In_751);
nor U3744 (N_3744,In_1185,In_1572);
and U3745 (N_3745,In_130,In_1668);
or U3746 (N_3746,In_93,In_222);
nand U3747 (N_3747,In_1022,In_391);
nor U3748 (N_3748,In_1224,In_1202);
nor U3749 (N_3749,In_1331,In_487);
nand U3750 (N_3750,In_419,In_1410);
and U3751 (N_3751,In_276,In_1554);
and U3752 (N_3752,In_445,In_791);
nand U3753 (N_3753,In_1867,In_633);
nor U3754 (N_3754,In_187,In_1231);
nor U3755 (N_3755,In_1164,In_673);
nand U3756 (N_3756,In_228,In_290);
and U3757 (N_3757,In_732,In_258);
and U3758 (N_3758,In_1255,In_1375);
nand U3759 (N_3759,In_1912,In_34);
nor U3760 (N_3760,In_1459,In_606);
or U3761 (N_3761,In_274,In_472);
nand U3762 (N_3762,In_173,In_92);
and U3763 (N_3763,In_1749,In_1619);
and U3764 (N_3764,In_90,In_608);
or U3765 (N_3765,In_320,In_392);
nand U3766 (N_3766,In_351,In_588);
and U3767 (N_3767,In_1512,In_1580);
or U3768 (N_3768,In_464,In_1933);
and U3769 (N_3769,In_1521,In_1295);
or U3770 (N_3770,In_1946,In_1484);
xor U3771 (N_3771,In_416,In_812);
nor U3772 (N_3772,In_1477,In_653);
xor U3773 (N_3773,In_218,In_652);
nor U3774 (N_3774,In_30,In_797);
or U3775 (N_3775,In_1664,In_1875);
nand U3776 (N_3776,In_1157,In_1539);
xor U3777 (N_3777,In_16,In_1094);
or U3778 (N_3778,In_1209,In_996);
nand U3779 (N_3779,In_233,In_46);
xnor U3780 (N_3780,In_816,In_1469);
nand U3781 (N_3781,In_102,In_512);
nor U3782 (N_3782,In_472,In_856);
or U3783 (N_3783,In_434,In_1708);
nor U3784 (N_3784,In_370,In_760);
or U3785 (N_3785,In_697,In_1059);
nand U3786 (N_3786,In_79,In_1437);
nor U3787 (N_3787,In_1694,In_705);
nor U3788 (N_3788,In_1259,In_656);
nand U3789 (N_3789,In_1670,In_461);
and U3790 (N_3790,In_115,In_1295);
xor U3791 (N_3791,In_301,In_1955);
and U3792 (N_3792,In_1905,In_106);
nor U3793 (N_3793,In_589,In_1139);
nor U3794 (N_3794,In_1396,In_1778);
nor U3795 (N_3795,In_1149,In_1579);
nand U3796 (N_3796,In_1051,In_1549);
nor U3797 (N_3797,In_1246,In_379);
nor U3798 (N_3798,In_1990,In_549);
and U3799 (N_3799,In_430,In_1759);
nor U3800 (N_3800,In_688,In_1725);
nor U3801 (N_3801,In_1457,In_1780);
nor U3802 (N_3802,In_1651,In_1936);
nor U3803 (N_3803,In_745,In_323);
and U3804 (N_3804,In_601,In_355);
xnor U3805 (N_3805,In_301,In_483);
or U3806 (N_3806,In_27,In_1525);
or U3807 (N_3807,In_204,In_1632);
xnor U3808 (N_3808,In_603,In_1591);
or U3809 (N_3809,In_740,In_1463);
nand U3810 (N_3810,In_390,In_332);
xor U3811 (N_3811,In_210,In_1064);
or U3812 (N_3812,In_669,In_1307);
xnor U3813 (N_3813,In_802,In_733);
and U3814 (N_3814,In_1006,In_1342);
nor U3815 (N_3815,In_1947,In_228);
nor U3816 (N_3816,In_1717,In_1695);
xnor U3817 (N_3817,In_968,In_1272);
xnor U3818 (N_3818,In_1363,In_451);
or U3819 (N_3819,In_597,In_753);
nand U3820 (N_3820,In_1698,In_4);
nor U3821 (N_3821,In_557,In_1789);
or U3822 (N_3822,In_1244,In_1052);
nor U3823 (N_3823,In_733,In_348);
nand U3824 (N_3824,In_313,In_366);
nor U3825 (N_3825,In_1140,In_210);
or U3826 (N_3826,In_1921,In_729);
nor U3827 (N_3827,In_1681,In_1252);
nor U3828 (N_3828,In_1813,In_646);
nand U3829 (N_3829,In_155,In_1762);
and U3830 (N_3830,In_497,In_435);
nand U3831 (N_3831,In_1131,In_801);
and U3832 (N_3832,In_1314,In_550);
or U3833 (N_3833,In_273,In_1288);
nand U3834 (N_3834,In_864,In_202);
nor U3835 (N_3835,In_1051,In_505);
and U3836 (N_3836,In_1721,In_790);
and U3837 (N_3837,In_255,In_1790);
or U3838 (N_3838,In_786,In_1130);
xnor U3839 (N_3839,In_74,In_445);
nor U3840 (N_3840,In_302,In_1402);
or U3841 (N_3841,In_1128,In_51);
nor U3842 (N_3842,In_712,In_848);
nand U3843 (N_3843,In_1003,In_1719);
or U3844 (N_3844,In_1085,In_766);
nor U3845 (N_3845,In_1336,In_1755);
or U3846 (N_3846,In_631,In_457);
nor U3847 (N_3847,In_1924,In_1528);
nor U3848 (N_3848,In_149,In_1140);
or U3849 (N_3849,In_1550,In_691);
and U3850 (N_3850,In_1518,In_567);
nand U3851 (N_3851,In_589,In_1726);
xnor U3852 (N_3852,In_1481,In_1706);
nor U3853 (N_3853,In_1734,In_1718);
and U3854 (N_3854,In_1027,In_1311);
or U3855 (N_3855,In_299,In_1442);
or U3856 (N_3856,In_176,In_777);
and U3857 (N_3857,In_894,In_1697);
nand U3858 (N_3858,In_925,In_1653);
nand U3859 (N_3859,In_844,In_1149);
and U3860 (N_3860,In_1908,In_97);
and U3861 (N_3861,In_641,In_838);
nor U3862 (N_3862,In_1519,In_239);
nand U3863 (N_3863,In_624,In_985);
xnor U3864 (N_3864,In_1222,In_1693);
xnor U3865 (N_3865,In_1033,In_209);
or U3866 (N_3866,In_1625,In_1216);
and U3867 (N_3867,In_740,In_295);
and U3868 (N_3868,In_1458,In_1405);
xnor U3869 (N_3869,In_494,In_1168);
and U3870 (N_3870,In_1767,In_1392);
or U3871 (N_3871,In_416,In_1841);
and U3872 (N_3872,In_1769,In_670);
or U3873 (N_3873,In_837,In_301);
and U3874 (N_3874,In_457,In_533);
xor U3875 (N_3875,In_1261,In_209);
and U3876 (N_3876,In_44,In_405);
nand U3877 (N_3877,In_1371,In_208);
or U3878 (N_3878,In_497,In_1991);
nand U3879 (N_3879,In_1444,In_1020);
or U3880 (N_3880,In_605,In_627);
nand U3881 (N_3881,In_1256,In_1444);
or U3882 (N_3882,In_416,In_883);
and U3883 (N_3883,In_1171,In_1756);
nand U3884 (N_3884,In_1903,In_522);
or U3885 (N_3885,In_250,In_412);
nor U3886 (N_3886,In_1188,In_357);
nor U3887 (N_3887,In_1941,In_486);
nand U3888 (N_3888,In_194,In_1139);
or U3889 (N_3889,In_1596,In_330);
nor U3890 (N_3890,In_484,In_40);
nor U3891 (N_3891,In_826,In_209);
and U3892 (N_3892,In_27,In_1725);
nand U3893 (N_3893,In_1015,In_896);
nor U3894 (N_3894,In_1629,In_1610);
and U3895 (N_3895,In_1644,In_408);
or U3896 (N_3896,In_1413,In_1628);
or U3897 (N_3897,In_460,In_1473);
and U3898 (N_3898,In_1689,In_310);
or U3899 (N_3899,In_1123,In_197);
or U3900 (N_3900,In_560,In_316);
nor U3901 (N_3901,In_1084,In_1552);
nor U3902 (N_3902,In_133,In_1904);
or U3903 (N_3903,In_884,In_1070);
nor U3904 (N_3904,In_704,In_450);
and U3905 (N_3905,In_670,In_1079);
and U3906 (N_3906,In_927,In_1153);
or U3907 (N_3907,In_1249,In_1423);
xnor U3908 (N_3908,In_645,In_1869);
or U3909 (N_3909,In_1337,In_1231);
nand U3910 (N_3910,In_1230,In_1024);
nand U3911 (N_3911,In_988,In_1691);
nor U3912 (N_3912,In_472,In_1138);
nor U3913 (N_3913,In_1249,In_35);
nand U3914 (N_3914,In_1096,In_564);
nor U3915 (N_3915,In_1678,In_1277);
nand U3916 (N_3916,In_269,In_1655);
nand U3917 (N_3917,In_1987,In_1418);
and U3918 (N_3918,In_1230,In_889);
or U3919 (N_3919,In_1362,In_378);
xnor U3920 (N_3920,In_535,In_552);
nor U3921 (N_3921,In_1693,In_572);
and U3922 (N_3922,In_1667,In_1812);
or U3923 (N_3923,In_368,In_431);
or U3924 (N_3924,In_547,In_1094);
nor U3925 (N_3925,In_1661,In_1968);
and U3926 (N_3926,In_938,In_235);
nand U3927 (N_3927,In_794,In_873);
nor U3928 (N_3928,In_1117,In_349);
nor U3929 (N_3929,In_800,In_1431);
nand U3930 (N_3930,In_1828,In_1759);
or U3931 (N_3931,In_903,In_598);
or U3932 (N_3932,In_390,In_1466);
xnor U3933 (N_3933,In_504,In_1939);
or U3934 (N_3934,In_1430,In_847);
and U3935 (N_3935,In_900,In_1518);
and U3936 (N_3936,In_738,In_1574);
or U3937 (N_3937,In_1481,In_1897);
or U3938 (N_3938,In_139,In_1315);
nand U3939 (N_3939,In_1696,In_239);
nand U3940 (N_3940,In_242,In_492);
and U3941 (N_3941,In_1670,In_766);
and U3942 (N_3942,In_1914,In_1710);
and U3943 (N_3943,In_219,In_1715);
and U3944 (N_3944,In_239,In_530);
or U3945 (N_3945,In_1545,In_1174);
nor U3946 (N_3946,In_1964,In_769);
xor U3947 (N_3947,In_1497,In_617);
and U3948 (N_3948,In_1653,In_876);
nor U3949 (N_3949,In_1751,In_1955);
nor U3950 (N_3950,In_1970,In_136);
and U3951 (N_3951,In_1628,In_644);
and U3952 (N_3952,In_1816,In_1043);
nand U3953 (N_3953,In_951,In_1701);
nand U3954 (N_3954,In_902,In_528);
nor U3955 (N_3955,In_258,In_1758);
or U3956 (N_3956,In_556,In_1189);
nand U3957 (N_3957,In_1009,In_365);
nand U3958 (N_3958,In_691,In_1162);
and U3959 (N_3959,In_959,In_1101);
and U3960 (N_3960,In_1869,In_103);
xnor U3961 (N_3961,In_400,In_865);
and U3962 (N_3962,In_767,In_995);
nor U3963 (N_3963,In_1884,In_68);
nor U3964 (N_3964,In_256,In_931);
nor U3965 (N_3965,In_1964,In_1485);
or U3966 (N_3966,In_1080,In_1294);
xnor U3967 (N_3967,In_1730,In_1984);
nor U3968 (N_3968,In_1199,In_988);
nand U3969 (N_3969,In_1020,In_1593);
or U3970 (N_3970,In_82,In_1971);
nor U3971 (N_3971,In_1482,In_1765);
or U3972 (N_3972,In_1708,In_1544);
nand U3973 (N_3973,In_1982,In_1594);
and U3974 (N_3974,In_1876,In_1011);
nor U3975 (N_3975,In_1435,In_751);
or U3976 (N_3976,In_450,In_357);
nor U3977 (N_3977,In_781,In_1094);
or U3978 (N_3978,In_1238,In_341);
nand U3979 (N_3979,In_765,In_1875);
nand U3980 (N_3980,In_1321,In_1310);
or U3981 (N_3981,In_736,In_1277);
nor U3982 (N_3982,In_1770,In_452);
nand U3983 (N_3983,In_574,In_584);
xor U3984 (N_3984,In_1024,In_472);
and U3985 (N_3985,In_1020,In_392);
or U3986 (N_3986,In_1480,In_1488);
or U3987 (N_3987,In_1859,In_1480);
and U3988 (N_3988,In_189,In_1032);
nor U3989 (N_3989,In_1875,In_1481);
nor U3990 (N_3990,In_1645,In_528);
or U3991 (N_3991,In_1391,In_688);
and U3992 (N_3992,In_1356,In_265);
and U3993 (N_3993,In_802,In_1649);
nand U3994 (N_3994,In_1873,In_19);
or U3995 (N_3995,In_1125,In_1879);
and U3996 (N_3996,In_1935,In_1424);
nor U3997 (N_3997,In_698,In_1220);
and U3998 (N_3998,In_70,In_95);
nor U3999 (N_3999,In_1038,In_1116);
and U4000 (N_4000,N_3680,N_3822);
nand U4001 (N_4001,N_3376,N_924);
and U4002 (N_4002,N_2056,N_2184);
nor U4003 (N_4003,N_2813,N_2080);
and U4004 (N_4004,N_3569,N_1733);
and U4005 (N_4005,N_532,N_2958);
nand U4006 (N_4006,N_732,N_486);
or U4007 (N_4007,N_3167,N_2016);
and U4008 (N_4008,N_3848,N_3778);
and U4009 (N_4009,N_1842,N_3929);
nand U4010 (N_4010,N_1208,N_2);
nand U4011 (N_4011,N_3427,N_1136);
or U4012 (N_4012,N_2992,N_3843);
and U4013 (N_4013,N_329,N_1890);
nand U4014 (N_4014,N_3551,N_3650);
or U4015 (N_4015,N_1020,N_1412);
or U4016 (N_4016,N_2158,N_3657);
or U4017 (N_4017,N_2105,N_3531);
nor U4018 (N_4018,N_1717,N_1658);
xnor U4019 (N_4019,N_822,N_1009);
xnor U4020 (N_4020,N_675,N_2096);
nor U4021 (N_4021,N_3597,N_3481);
xor U4022 (N_4022,N_2589,N_3095);
nand U4023 (N_4023,N_2608,N_1268);
nor U4024 (N_4024,N_129,N_811);
nand U4025 (N_4025,N_2546,N_2790);
and U4026 (N_4026,N_896,N_3284);
nand U4027 (N_4027,N_1666,N_3614);
and U4028 (N_4028,N_1444,N_2991);
nor U4029 (N_4029,N_1931,N_2865);
and U4030 (N_4030,N_615,N_661);
nand U4031 (N_4031,N_2462,N_2422);
nor U4032 (N_4032,N_1740,N_3892);
and U4033 (N_4033,N_3156,N_507);
or U4034 (N_4034,N_2383,N_94);
nand U4035 (N_4035,N_3611,N_1430);
nand U4036 (N_4036,N_1448,N_3369);
or U4037 (N_4037,N_1787,N_1005);
and U4038 (N_4038,N_2543,N_3838);
xnor U4039 (N_4039,N_1022,N_442);
nand U4040 (N_4040,N_2671,N_3518);
nor U4041 (N_4041,N_1129,N_3114);
and U4042 (N_4042,N_2092,N_810);
nor U4043 (N_4043,N_3087,N_2504);
nor U4044 (N_4044,N_3283,N_3493);
or U4045 (N_4045,N_626,N_3533);
or U4046 (N_4046,N_2627,N_674);
and U4047 (N_4047,N_1859,N_851);
and U4048 (N_4048,N_1610,N_2057);
and U4049 (N_4049,N_3814,N_2540);
nand U4050 (N_4050,N_3578,N_3863);
nand U4051 (N_4051,N_1767,N_158);
or U4052 (N_4052,N_1607,N_2690);
nor U4053 (N_4053,N_1651,N_999);
and U4054 (N_4054,N_225,N_2493);
nor U4055 (N_4055,N_2325,N_2647);
or U4056 (N_4056,N_448,N_1392);
nor U4057 (N_4057,N_1739,N_359);
nor U4058 (N_4058,N_808,N_2379);
nand U4059 (N_4059,N_2240,N_3761);
nand U4060 (N_4060,N_1612,N_2773);
xor U4061 (N_4061,N_2639,N_3445);
and U4062 (N_4062,N_914,N_3270);
nand U4063 (N_4063,N_743,N_2413);
and U4064 (N_4064,N_3251,N_171);
and U4065 (N_4065,N_93,N_2272);
nor U4066 (N_4066,N_861,N_1528);
nand U4067 (N_4067,N_2837,N_2831);
and U4068 (N_4068,N_2825,N_2220);
or U4069 (N_4069,N_1302,N_2883);
and U4070 (N_4070,N_887,N_3756);
xnor U4071 (N_4071,N_320,N_3277);
nand U4072 (N_4072,N_3046,N_1289);
nor U4073 (N_4073,N_1923,N_3148);
nand U4074 (N_4074,N_1903,N_3220);
nand U4075 (N_4075,N_2094,N_2557);
or U4076 (N_4076,N_513,N_47);
nor U4077 (N_4077,N_3656,N_3997);
nor U4078 (N_4078,N_739,N_3991);
or U4079 (N_4079,N_2547,N_3617);
nand U4080 (N_4080,N_2595,N_3763);
nor U4081 (N_4081,N_3223,N_1635);
xor U4082 (N_4082,N_2154,N_145);
and U4083 (N_4083,N_1569,N_457);
or U4084 (N_4084,N_3951,N_3714);
nor U4085 (N_4085,N_514,N_781);
nor U4086 (N_4086,N_1453,N_809);
and U4087 (N_4087,N_2536,N_1193);
xor U4088 (N_4088,N_2732,N_1535);
nand U4089 (N_4089,N_693,N_1078);
xor U4090 (N_4090,N_1529,N_860);
and U4091 (N_4091,N_3374,N_213);
nor U4092 (N_4092,N_1937,N_1714);
or U4093 (N_4093,N_2053,N_3889);
or U4094 (N_4094,N_3624,N_2706);
xnor U4095 (N_4095,N_3032,N_2606);
nand U4096 (N_4096,N_2443,N_2797);
nor U4097 (N_4097,N_3135,N_900);
and U4098 (N_4098,N_2194,N_3126);
and U4099 (N_4099,N_1347,N_2609);
and U4100 (N_4100,N_819,N_2115);
and U4101 (N_4101,N_107,N_2229);
or U4102 (N_4102,N_2988,N_1017);
and U4103 (N_4103,N_2385,N_2784);
nand U4104 (N_4104,N_519,N_2245);
nor U4105 (N_4105,N_1650,N_836);
or U4106 (N_4106,N_2049,N_3579);
and U4107 (N_4107,N_1500,N_3600);
nand U4108 (N_4108,N_389,N_3887);
and U4109 (N_4109,N_1488,N_2394);
nand U4110 (N_4110,N_3788,N_371);
nor U4111 (N_4111,N_1463,N_3218);
nand U4112 (N_4112,N_535,N_2370);
and U4113 (N_4113,N_3049,N_431);
nand U4114 (N_4114,N_3994,N_3237);
nand U4115 (N_4115,N_3219,N_3820);
or U4116 (N_4116,N_3279,N_2852);
nand U4117 (N_4117,N_1369,N_1396);
and U4118 (N_4118,N_2404,N_2928);
nand U4119 (N_4119,N_3799,N_3988);
or U4120 (N_4120,N_3603,N_908);
or U4121 (N_4121,N_3268,N_2276);
nor U4122 (N_4122,N_1323,N_1883);
nor U4123 (N_4123,N_3366,N_2983);
or U4124 (N_4124,N_2913,N_1209);
or U4125 (N_4125,N_901,N_3652);
nor U4126 (N_4126,N_3409,N_951);
or U4127 (N_4127,N_1655,N_1893);
or U4128 (N_4128,N_2836,N_1509);
nand U4129 (N_4129,N_2938,N_711);
or U4130 (N_4130,N_2399,N_812);
nand U4131 (N_4131,N_1846,N_1382);
or U4132 (N_4132,N_1711,N_501);
and U4133 (N_4133,N_3587,N_3999);
xor U4134 (N_4134,N_2352,N_1605);
and U4135 (N_4135,N_534,N_1844);
nand U4136 (N_4136,N_1068,N_2728);
and U4137 (N_4137,N_2045,N_1913);
nor U4138 (N_4138,N_2658,N_2452);
nor U4139 (N_4139,N_889,N_2727);
or U4140 (N_4140,N_2204,N_3222);
and U4141 (N_4141,N_981,N_545);
nand U4142 (N_4142,N_3361,N_2231);
and U4143 (N_4143,N_3496,N_202);
and U4144 (N_4144,N_3478,N_3598);
and U4145 (N_4145,N_2306,N_1641);
nand U4146 (N_4146,N_2791,N_3082);
or U4147 (N_4147,N_3451,N_622);
and U4148 (N_4148,N_103,N_686);
or U4149 (N_4149,N_2774,N_2844);
and U4150 (N_4150,N_2392,N_3417);
or U4151 (N_4151,N_2261,N_1928);
nand U4152 (N_4152,N_3976,N_655);
nand U4153 (N_4153,N_943,N_2775);
and U4154 (N_4154,N_2283,N_2406);
nand U4155 (N_4155,N_1083,N_1097);
nand U4156 (N_4156,N_2402,N_2042);
nand U4157 (N_4157,N_740,N_3421);
or U4158 (N_4158,N_1737,N_911);
nor U4159 (N_4159,N_789,N_802);
and U4160 (N_4160,N_3819,N_1161);
nor U4161 (N_4161,N_1356,N_2485);
nor U4162 (N_4162,N_3815,N_2280);
and U4163 (N_4163,N_2167,N_2268);
and U4164 (N_4164,N_1979,N_3190);
xnor U4165 (N_4165,N_904,N_3310);
nor U4166 (N_4166,N_2720,N_1592);
or U4167 (N_4167,N_1933,N_299);
xnor U4168 (N_4168,N_800,N_1867);
nor U4169 (N_4169,N_1315,N_1037);
nor U4170 (N_4170,N_363,N_3331);
or U4171 (N_4171,N_3258,N_1755);
or U4172 (N_4172,N_3038,N_3159);
and U4173 (N_4173,N_1627,N_512);
nand U4174 (N_4174,N_584,N_474);
nand U4175 (N_4175,N_2340,N_2177);
nor U4176 (N_4176,N_3048,N_1510);
xnor U4177 (N_4177,N_2926,N_342);
or U4178 (N_4178,N_415,N_3716);
and U4179 (N_4179,N_2253,N_3036);
or U4180 (N_4180,N_2739,N_1874);
or U4181 (N_4181,N_3448,N_197);
nor U4182 (N_4182,N_3945,N_1970);
and U4183 (N_4183,N_1590,N_1858);
or U4184 (N_4184,N_560,N_2564);
nor U4185 (N_4185,N_3910,N_2679);
xnor U4186 (N_4186,N_3912,N_1971);
nand U4187 (N_4187,N_3691,N_2922);
nor U4188 (N_4188,N_365,N_134);
or U4189 (N_4189,N_849,N_3803);
or U4190 (N_4190,N_153,N_1828);
and U4191 (N_4191,N_1667,N_3018);
or U4192 (N_4192,N_1887,N_3468);
or U4193 (N_4193,N_1332,N_72);
and U4194 (N_4194,N_3825,N_1327);
or U4195 (N_4195,N_1433,N_287);
xor U4196 (N_4196,N_1517,N_2886);
and U4197 (N_4197,N_3362,N_2834);
nor U4198 (N_4198,N_587,N_3171);
nand U4199 (N_4199,N_3253,N_3630);
or U4200 (N_4200,N_1993,N_3174);
nand U4201 (N_4201,N_445,N_1987);
xor U4202 (N_4202,N_3970,N_1270);
xor U4203 (N_4203,N_3584,N_2409);
nor U4204 (N_4204,N_2651,N_888);
nand U4205 (N_4205,N_2555,N_189);
nand U4206 (N_4206,N_1511,N_2211);
or U4207 (N_4207,N_1777,N_2709);
and U4208 (N_4208,N_3397,N_3917);
nor U4209 (N_4209,N_3944,N_1324);
nor U4210 (N_4210,N_2190,N_2026);
and U4211 (N_4211,N_2336,N_133);
or U4212 (N_4212,N_2110,N_2420);
or U4213 (N_4213,N_958,N_2722);
nand U4214 (N_4214,N_1969,N_1124);
nand U4215 (N_4215,N_2839,N_151);
and U4216 (N_4216,N_1222,N_1845);
or U4217 (N_4217,N_2697,N_3086);
nor U4218 (N_4218,N_654,N_297);
xor U4219 (N_4219,N_978,N_32);
and U4220 (N_4220,N_88,N_2532);
nor U4221 (N_4221,N_2556,N_2113);
nor U4222 (N_4222,N_1705,N_466);
or U4223 (N_4223,N_1829,N_1484);
nand U4224 (N_4224,N_1772,N_3981);
and U4225 (N_4225,N_1045,N_2685);
nand U4226 (N_4226,N_2902,N_823);
nor U4227 (N_4227,N_1227,N_2971);
and U4228 (N_4228,N_1095,N_3226);
and U4229 (N_4229,N_2475,N_3700);
and U4230 (N_4230,N_3818,N_2391);
or U4231 (N_4231,N_51,N_3107);
or U4232 (N_4232,N_2680,N_1762);
nand U4233 (N_4233,N_379,N_1120);
or U4234 (N_4234,N_3149,N_366);
nor U4235 (N_4235,N_3425,N_1371);
xnor U4236 (N_4236,N_376,N_1113);
or U4237 (N_4237,N_96,N_1905);
nand U4238 (N_4238,N_2318,N_2206);
nand U4239 (N_4239,N_232,N_2172);
nor U4240 (N_4240,N_1404,N_623);
xnor U4241 (N_4241,N_2098,N_3888);
and U4242 (N_4242,N_85,N_3653);
or U4243 (N_4243,N_1431,N_2818);
or U4244 (N_4244,N_877,N_3150);
or U4245 (N_4245,N_1977,N_3278);
nor U4246 (N_4246,N_2994,N_2232);
or U4247 (N_4247,N_912,N_3968);
and U4248 (N_4248,N_1114,N_2754);
nor U4249 (N_4249,N_2386,N_84);
or U4250 (N_4250,N_629,N_2711);
nor U4251 (N_4251,N_1978,N_2866);
and U4252 (N_4252,N_2257,N_1275);
and U4253 (N_4253,N_105,N_3766);
nor U4254 (N_4254,N_1060,N_2918);
and U4255 (N_4255,N_2858,N_1850);
or U4256 (N_4256,N_1902,N_2473);
nor U4257 (N_4257,N_1101,N_2324);
and U4258 (N_4258,N_1831,N_2959);
nand U4259 (N_4259,N_966,N_3249);
xnor U4260 (N_4260,N_2565,N_1881);
or U4261 (N_4261,N_3909,N_483);
and U4262 (N_4262,N_3117,N_2970);
and U4263 (N_4263,N_455,N_182);
nor U4264 (N_4264,N_1443,N_926);
xor U4265 (N_4265,N_3088,N_2932);
nand U4266 (N_4266,N_2884,N_333);
or U4267 (N_4267,N_2648,N_1712);
nor U4268 (N_4268,N_1586,N_2246);
or U4269 (N_4269,N_2695,N_3817);
or U4270 (N_4270,N_2024,N_2981);
nand U4271 (N_4271,N_611,N_2411);
nor U4272 (N_4272,N_1322,N_2795);
and U4273 (N_4273,N_2888,N_75);
or U4274 (N_4274,N_1074,N_2300);
or U4275 (N_4275,N_2949,N_3878);
and U4276 (N_4276,N_3155,N_3660);
and U4277 (N_4277,N_2474,N_458);
or U4278 (N_4278,N_2946,N_405);
nor U4279 (N_4279,N_1056,N_1941);
or U4280 (N_4280,N_1450,N_2762);
and U4281 (N_4281,N_794,N_3798);
nor U4282 (N_4282,N_2696,N_2366);
or U4283 (N_4283,N_2599,N_1819);
or U4284 (N_4284,N_1638,N_757);
nor U4285 (N_4285,N_1219,N_847);
nor U4286 (N_4286,N_73,N_1091);
and U4287 (N_4287,N_1698,N_3883);
and U4288 (N_4288,N_87,N_3835);
nand U4289 (N_4289,N_175,N_268);
nand U4290 (N_4290,N_1361,N_3373);
nand U4291 (N_4291,N_1646,N_3961);
nand U4292 (N_4292,N_357,N_2179);
nand U4293 (N_4293,N_2617,N_1279);
and U4294 (N_4294,N_1104,N_2381);
and U4295 (N_4295,N_1507,N_3552);
and U4296 (N_4296,N_1560,N_3083);
xnor U4297 (N_4297,N_3881,N_211);
nor U4298 (N_4298,N_697,N_1008);
and U4299 (N_4299,N_1898,N_2623);
nor U4300 (N_4300,N_1699,N_1585);
nor U4301 (N_4301,N_1377,N_1052);
nand U4302 (N_4302,N_2665,N_824);
or U4303 (N_4303,N_195,N_3077);
and U4304 (N_4304,N_2315,N_1892);
or U4305 (N_4305,N_497,N_1454);
nand U4306 (N_4306,N_3420,N_2141);
nand U4307 (N_4307,N_1732,N_1836);
or U4308 (N_4308,N_3963,N_3966);
nor U4309 (N_4309,N_1197,N_3539);
nor U4310 (N_4310,N_1873,N_2664);
nand U4311 (N_4311,N_2088,N_893);
or U4312 (N_4312,N_132,N_1564);
nand U4313 (N_4313,N_2718,N_3685);
or U4314 (N_4314,N_2495,N_1589);
and U4315 (N_4315,N_3664,N_662);
xor U4316 (N_4316,N_3172,N_2631);
and U4317 (N_4317,N_2183,N_3248);
nor U4318 (N_4318,N_1326,N_2066);
and U4319 (N_4319,N_2998,N_3252);
nor U4320 (N_4320,N_476,N_3751);
or U4321 (N_4321,N_2840,N_2731);
nand U4322 (N_4322,N_2345,N_2126);
and U4323 (N_4323,N_3859,N_3068);
and U4324 (N_4324,N_1587,N_1662);
or U4325 (N_4325,N_3382,N_2523);
and U4326 (N_4326,N_2770,N_1385);
or U4327 (N_4327,N_1783,N_500);
nand U4328 (N_4328,N_3572,N_2821);
nand U4329 (N_4329,N_1034,N_336);
or U4330 (N_4330,N_2093,N_122);
and U4331 (N_4331,N_3338,N_2657);
nand U4332 (N_4332,N_374,N_60);
and U4333 (N_4333,N_902,N_1687);
nand U4334 (N_4334,N_3666,N_1946);
nor U4335 (N_4335,N_1615,N_637);
and U4336 (N_4336,N_2851,N_2396);
nor U4337 (N_4337,N_1989,N_3341);
and U4338 (N_4338,N_1276,N_716);
nor U4339 (N_4339,N_1678,N_567);
nor U4340 (N_4340,N_45,N_1201);
or U4341 (N_4341,N_2864,N_1421);
nor U4342 (N_4342,N_343,N_2307);
and U4343 (N_4343,N_2186,N_1491);
or U4344 (N_4344,N_115,N_837);
nand U4345 (N_4345,N_3923,N_2103);
and U4346 (N_4346,N_1947,N_3715);
or U4347 (N_4347,N_1644,N_765);
nor U4348 (N_4348,N_3722,N_2330);
nand U4349 (N_4349,N_3677,N_1797);
nor U4350 (N_4350,N_727,N_948);
or U4351 (N_4351,N_987,N_1824);
nor U4352 (N_4352,N_3008,N_309);
and U4353 (N_4353,N_746,N_1288);
or U4354 (N_4354,N_1548,N_438);
and U4355 (N_4355,N_940,N_3105);
nand U4356 (N_4356,N_1985,N_1749);
xor U4357 (N_4357,N_3428,N_2271);
and U4358 (N_4358,N_969,N_563);
and U4359 (N_4359,N_421,N_1487);
nand U4360 (N_4360,N_1127,N_2410);
or U4361 (N_4361,N_2957,N_866);
or U4362 (N_4362,N_3161,N_3683);
nand U4363 (N_4363,N_3244,N_270);
nor U4364 (N_4364,N_2419,N_1178);
and U4365 (N_4365,N_971,N_2581);
and U4366 (N_4366,N_2823,N_506);
and U4367 (N_4367,N_773,N_2051);
and U4368 (N_4368,N_1282,N_3675);
and U4369 (N_4369,N_1494,N_1531);
or U4370 (N_4370,N_3254,N_261);
nand U4371 (N_4371,N_643,N_125);
or U4372 (N_4372,N_3906,N_556);
or U4373 (N_4373,N_1110,N_1281);
nor U4374 (N_4374,N_3595,N_1062);
and U4375 (N_4375,N_1362,N_2202);
nand U4376 (N_4376,N_2193,N_1580);
and U4377 (N_4377,N_8,N_551);
or U4378 (N_4378,N_1794,N_2963);
nor U4379 (N_4379,N_3378,N_710);
and U4380 (N_4380,N_186,N_3467);
and U4381 (N_4381,N_2900,N_355);
and U4382 (N_4382,N_3986,N_792);
or U4383 (N_4383,N_222,N_1861);
or U4384 (N_4384,N_2130,N_853);
nor U4385 (N_4385,N_1550,N_1907);
nor U4386 (N_4386,N_3489,N_1796);
xor U4387 (N_4387,N_1004,N_1939);
and U4388 (N_4388,N_1960,N_161);
or U4389 (N_4389,N_2414,N_2487);
and U4390 (N_4390,N_3011,N_2243);
nor U4391 (N_4391,N_592,N_1776);
or U4392 (N_4392,N_2525,N_2436);
nand U4393 (N_4393,N_2804,N_1770);
and U4394 (N_4394,N_3506,N_3476);
nand U4395 (N_4395,N_1990,N_1827);
nand U4396 (N_4396,N_2353,N_1713);
nand U4397 (N_4397,N_1496,N_1061);
or U4398 (N_4398,N_181,N_1472);
and U4399 (N_4399,N_150,N_467);
and U4400 (N_4400,N_605,N_1233);
or U4401 (N_4401,N_2277,N_3439);
or U4402 (N_4402,N_2252,N_1793);
nand U4403 (N_4403,N_3027,N_2433);
nand U4404 (N_4404,N_2046,N_1109);
xor U4405 (N_4405,N_2986,N_1806);
xnor U4406 (N_4406,N_3354,N_2374);
and U4407 (N_4407,N_2264,N_148);
nor U4408 (N_4408,N_3871,N_1578);
and U4409 (N_4409,N_2012,N_2135);
and U4410 (N_4410,N_2917,N_1389);
nor U4411 (N_4411,N_1912,N_2102);
nand U4412 (N_4412,N_3651,N_2239);
or U4413 (N_4413,N_2314,N_3124);
xor U4414 (N_4414,N_2430,N_3588);
or U4415 (N_4415,N_3127,N_3793);
nor U4416 (N_4416,N_3480,N_1352);
or U4417 (N_4417,N_1452,N_1613);
nand U4418 (N_4418,N_3875,N_2048);
nor U4419 (N_4419,N_2979,N_3522);
nor U4420 (N_4420,N_852,N_425);
nand U4421 (N_4421,N_1121,N_3065);
nand U4422 (N_4422,N_2999,N_2893);
or U4423 (N_4423,N_2757,N_3646);
nor U4424 (N_4424,N_2638,N_2808);
xor U4425 (N_4425,N_1599,N_21);
nand U4426 (N_4426,N_1896,N_3599);
and U4427 (N_4427,N_3402,N_843);
and U4428 (N_4428,N_3564,N_3816);
xor U4429 (N_4429,N_3558,N_216);
and U4430 (N_4430,N_1837,N_1381);
nor U4431 (N_4431,N_3667,N_269);
and U4432 (N_4432,N_388,N_2029);
nand U4433 (N_4433,N_2930,N_250);
and U4434 (N_4434,N_3876,N_1163);
nor U4435 (N_4435,N_3777,N_1403);
nand U4436 (N_4436,N_1130,N_2439);
nor U4437 (N_4437,N_219,N_1616);
xnor U4438 (N_4438,N_1042,N_1349);
and U4439 (N_4439,N_638,N_690);
nand U4440 (N_4440,N_1365,N_785);
and U4441 (N_4441,N_1584,N_2263);
nor U4442 (N_4442,N_116,N_2191);
or U4443 (N_4443,N_2768,N_2673);
or U4444 (N_4444,N_2227,N_214);
or U4445 (N_4445,N_1194,N_3854);
nand U4446 (N_4446,N_360,N_2656);
nor U4447 (N_4447,N_2437,N_3001);
and U4448 (N_4448,N_2490,N_2182);
and U4449 (N_4449,N_639,N_684);
and U4450 (N_4450,N_2329,N_2919);
and U4451 (N_4451,N_2223,N_44);
xor U4452 (N_4452,N_1264,N_373);
nor U4453 (N_4453,N_524,N_3749);
nand U4454 (N_4454,N_286,N_930);
or U4455 (N_4455,N_2855,N_627);
nand U4456 (N_4456,N_3288,N_1050);
or U4457 (N_4457,N_3261,N_2552);
nand U4458 (N_4458,N_3596,N_1891);
nand U4459 (N_4459,N_3760,N_2766);
and U4460 (N_4460,N_1354,N_387);
or U4461 (N_4461,N_3045,N_2961);
or U4462 (N_4462,N_2593,N_3710);
and U4463 (N_4463,N_417,N_1160);
nor U4464 (N_4464,N_672,N_2131);
xor U4465 (N_4465,N_1287,N_1218);
nand U4466 (N_4466,N_2378,N_946);
or U4467 (N_4467,N_2972,N_2514);
nand U4468 (N_4468,N_3509,N_1090);
nor U4469 (N_4469,N_3543,N_3524);
nor U4470 (N_4470,N_2342,N_1563);
or U4471 (N_4471,N_3092,N_3574);
nand U4472 (N_4472,N_3385,N_680);
or U4473 (N_4473,N_2400,N_2729);
and U4474 (N_4474,N_2934,N_330);
nand U4475 (N_4475,N_3381,N_2746);
or U4476 (N_4476,N_3457,N_2134);
and U4477 (N_4477,N_2786,N_2085);
and U4478 (N_4478,N_3673,N_3239);
nor U4479 (N_4479,N_3056,N_191);
and U4480 (N_4480,N_322,N_338);
nand U4481 (N_4481,N_1724,N_1840);
nand U4482 (N_4482,N_588,N_1838);
xor U4483 (N_4483,N_1286,N_679);
or U4484 (N_4484,N_392,N_100);
nand U4485 (N_4485,N_3462,N_980);
nor U4486 (N_4486,N_2175,N_435);
nand U4487 (N_4487,N_2798,N_1930);
and U4488 (N_4488,N_140,N_3739);
nand U4489 (N_4489,N_3300,N_2138);
and U4490 (N_4490,N_3946,N_1583);
xor U4491 (N_4491,N_3037,N_3166);
and U4492 (N_4492,N_2265,N_1555);
nor U4493 (N_4493,N_2987,N_2824);
or U4494 (N_4494,N_2403,N_2682);
nand U4495 (N_4495,N_597,N_209);
nor U4496 (N_4496,N_282,N_2629);
nand U4497 (N_4497,N_1618,N_296);
nand U4498 (N_4498,N_1871,N_3850);
or U4499 (N_4499,N_2666,N_2829);
and U4500 (N_4500,N_2519,N_2921);
or U4501 (N_4501,N_3943,N_1333);
xnor U4502 (N_4502,N_1596,N_1862);
and U4503 (N_4503,N_1379,N_2905);
nand U4504 (N_4504,N_3780,N_3712);
nor U4505 (N_4505,N_1546,N_169);
or U4506 (N_4506,N_3009,N_2426);
and U4507 (N_4507,N_3511,N_576);
and U4508 (N_4508,N_1790,N_3202);
nand U4509 (N_4509,N_3186,N_1682);
or U4510 (N_4510,N_3618,N_273);
nand U4511 (N_4511,N_1458,N_3307);
xor U4512 (N_4512,N_3089,N_3111);
and U4513 (N_4513,N_2524,N_2541);
or U4514 (N_4514,N_1951,N_659);
or U4515 (N_4515,N_2212,N_1927);
nor U4516 (N_4516,N_1417,N_1346);
nand U4517 (N_4517,N_1826,N_776);
nor U4518 (N_4518,N_2445,N_1665);
nand U4519 (N_4519,N_1133,N_3977);
nand U4520 (N_4520,N_257,N_1813);
nand U4521 (N_4521,N_3776,N_27);
and U4522 (N_4522,N_3304,N_3449);
or U4523 (N_4523,N_1521,N_2869);
or U4524 (N_4524,N_596,N_787);
xnor U4525 (N_4525,N_1864,N_783);
or U4526 (N_4526,N_2989,N_3713);
nand U4527 (N_4527,N_65,N_3686);
and U4528 (N_4528,N_3231,N_2794);
and U4529 (N_4529,N_3726,N_992);
nand U4530 (N_4530,N_42,N_1476);
and U4531 (N_4531,N_1805,N_2969);
nor U4532 (N_4532,N_883,N_1808);
nand U4533 (N_4533,N_1936,N_244);
nor U4534 (N_4534,N_2649,N_1547);
nor U4535 (N_4535,N_2692,N_265);
nor U4536 (N_4536,N_985,N_2801);
nor U4537 (N_4537,N_3375,N_828);
nand U4538 (N_4538,N_671,N_472);
or U4539 (N_4539,N_1435,N_807);
and U4540 (N_4540,N_997,N_2501);
nand U4541 (N_4541,N_3631,N_2654);
xnor U4542 (N_4542,N_404,N_2341);
or U4543 (N_4543,N_872,N_223);
nand U4544 (N_4544,N_1809,N_1328);
xor U4545 (N_4545,N_480,N_2037);
or U4546 (N_4546,N_198,N_368);
nor U4547 (N_4547,N_2901,N_1076);
xor U4548 (N_4548,N_2457,N_2259);
nor U4549 (N_4549,N_1621,N_3648);
nand U4550 (N_4550,N_3670,N_2146);
xnor U4551 (N_4551,N_3554,N_1729);
nand U4552 (N_4552,N_1801,N_1111);
and U4553 (N_4553,N_2293,N_1059);
xnor U4554 (N_4554,N_3266,N_3858);
nor U4555 (N_4555,N_3995,N_2713);
and U4556 (N_4556,N_3975,N_1138);
or U4557 (N_4557,N_1290,N_650);
xor U4558 (N_4558,N_2674,N_183);
nor U4559 (N_4559,N_1919,N_1530);
or U4560 (N_4560,N_1058,N_3334);
nor U4561 (N_4561,N_1962,N_3418);
nor U4562 (N_4562,N_2527,N_3494);
and U4563 (N_4563,N_3786,N_3422);
xnor U4564 (N_4564,N_413,N_3952);
or U4565 (N_4565,N_1336,N_1541);
xnor U4566 (N_4566,N_1660,N_972);
and U4567 (N_4567,N_1284,N_3504);
or U4568 (N_4568,N_1703,N_3235);
nor U4569 (N_4569,N_3285,N_2672);
and U4570 (N_4570,N_179,N_2077);
nor U4571 (N_4571,N_2192,N_3163);
xnor U4572 (N_4572,N_504,N_1670);
nand U4573 (N_4573,N_1259,N_2241);
or U4574 (N_4574,N_3787,N_1906);
and U4575 (N_4575,N_2576,N_3575);
xor U4576 (N_4576,N_2973,N_291);
nand U4577 (N_4577,N_720,N_2817);
and U4578 (N_4578,N_2082,N_3781);
nand U4579 (N_4579,N_351,N_2694);
nand U4580 (N_4580,N_2751,N_2575);
or U4581 (N_4581,N_1278,N_1470);
and U4582 (N_4582,N_3571,N_699);
nor U4583 (N_4583,N_2362,N_2297);
and U4584 (N_4584,N_3195,N_1899);
and U4585 (N_4585,N_1986,N_2755);
and U4586 (N_4586,N_390,N_2912);
nand U4587 (N_4587,N_747,N_2974);
and U4588 (N_4588,N_2405,N_2136);
xor U4589 (N_4589,N_1865,N_2633);
and U4590 (N_4590,N_2365,N_1934);
or U4591 (N_4591,N_3510,N_1350);
nor U4592 (N_4592,N_2363,N_2558);
nand U4593 (N_4593,N_280,N_1664);
nand U4594 (N_4594,N_3434,N_2234);
xor U4595 (N_4595,N_2249,N_3993);
and U4596 (N_4596,N_3309,N_1501);
nor U4597 (N_4597,N_63,N_2064);
nor U4598 (N_4598,N_470,N_3865);
xnor U4599 (N_4599,N_1224,N_1321);
nor U4600 (N_4600,N_2164,N_600);
nand U4601 (N_4601,N_3070,N_54);
nor U4602 (N_4602,N_2553,N_1765);
nand U4603 (N_4603,N_2787,N_3639);
or U4604 (N_4604,N_813,N_117);
and U4605 (N_4605,N_2025,N_1967);
nand U4606 (N_4606,N_1524,N_318);
nor U4607 (N_4607,N_1426,N_1774);
nor U4608 (N_4608,N_57,N_1185);
or U4609 (N_4609,N_2067,N_3517);
nand U4610 (N_4610,N_3849,N_1677);
or U4611 (N_4611,N_2478,N_328);
nand U4612 (N_4612,N_395,N_3413);
nor U4613 (N_4613,N_3209,N_217);
nand U4614 (N_4614,N_581,N_3267);
nor U4615 (N_4615,N_400,N_3470);
and U4616 (N_4616,N_3989,N_1786);
and U4617 (N_4617,N_1676,N_226);
or U4618 (N_4618,N_3679,N_3286);
nor U4619 (N_4619,N_3152,N_1976);
nand U4620 (N_4620,N_2014,N_3841);
and U4621 (N_4621,N_964,N_3262);
nor U4622 (N_4622,N_2605,N_3521);
nor U4623 (N_4623,N_1815,N_449);
xnor U4624 (N_4624,N_647,N_2904);
and U4625 (N_4625,N_938,N_256);
and U4626 (N_4626,N_2395,N_3019);
nor U4627 (N_4627,N_432,N_308);
or U4628 (N_4628,N_2091,N_427);
or U4629 (N_4629,N_1600,N_4);
or U4630 (N_4630,N_3151,N_2978);
xor U4631 (N_4631,N_2145,N_1473);
and U4632 (N_4632,N_665,N_3767);
nor U4633 (N_4633,N_3059,N_891);
or U4634 (N_4634,N_1393,N_619);
and U4635 (N_4635,N_2453,N_2127);
or U4636 (N_4636,N_670,N_3965);
nor U4637 (N_4637,N_2712,N_135);
nand U4638 (N_4638,N_3292,N_2856);
or U4639 (N_4639,N_3625,N_170);
xor U4640 (N_4640,N_606,N_3949);
nor U4641 (N_4641,N_3138,N_1540);
nor U4642 (N_4642,N_521,N_1566);
and U4643 (N_4643,N_2346,N_386);
nor U4644 (N_4644,N_1388,N_479);
and U4645 (N_4645,N_3079,N_2559);
nand U4646 (N_4646,N_977,N_446);
nor U4647 (N_4647,N_3932,N_2168);
nor U4648 (N_4648,N_2357,N_1174);
nor U4649 (N_4649,N_3407,N_2686);
or U4650 (N_4650,N_2238,N_74);
nand U4651 (N_4651,N_3210,N_3436);
nor U4652 (N_4652,N_3196,N_3842);
or U4653 (N_4653,N_267,N_712);
nand U4654 (N_4654,N_2539,N_177);
nor U4655 (N_4655,N_3440,N_3523);
nor U4656 (N_4656,N_1910,N_2767);
and U4657 (N_4657,N_3426,N_1345);
and U4658 (N_4658,N_656,N_2566);
xnor U4659 (N_4659,N_2267,N_1571);
or U4660 (N_4660,N_264,N_2388);
nor U4661 (N_4661,N_1439,N_2715);
nor U4662 (N_4662,N_3669,N_3096);
xor U4663 (N_4663,N_3689,N_1598);
or U4664 (N_4664,N_3924,N_3941);
or U4665 (N_4665,N_284,N_242);
nand U4666 (N_4666,N_3622,N_3372);
and U4667 (N_4667,N_2914,N_3905);
and U4668 (N_4668,N_2843,N_1285);
nor U4669 (N_4669,N_1608,N_1897);
nor U4670 (N_4670,N_3931,N_657);
or U4671 (N_4671,N_1123,N_11);
and U4672 (N_4672,N_2653,N_3747);
nor U4673 (N_4673,N_3157,N_3581);
or U4674 (N_4674,N_314,N_2667);
nor U4675 (N_4675,N_2714,N_2322);
xnor U4676 (N_4676,N_886,N_399);
nor U4677 (N_4677,N_3663,N_707);
and U4678 (N_4678,N_1527,N_1447);
or U4679 (N_4679,N_2187,N_1157);
nor U4680 (N_4680,N_3029,N_1788);
and U4681 (N_4681,N_2597,N_304);
and U4682 (N_4682,N_1206,N_867);
nand U4683 (N_4683,N_681,N_1959);
and U4684 (N_4684,N_994,N_1816);
nand U4685 (N_4685,N_3536,N_2213);
nor U4686 (N_4686,N_2181,N_1957);
nor U4687 (N_4687,N_2360,N_1738);
xor U4688 (N_4688,N_1707,N_114);
nor U4689 (N_4689,N_3719,N_1177);
xor U4690 (N_4690,N_2945,N_204);
xor U4691 (N_4691,N_334,N_3594);
nand U4692 (N_4692,N_230,N_354);
nor U4693 (N_4693,N_137,N_3050);
nor U4694 (N_4694,N_1366,N_3168);
nand U4695 (N_4695,N_516,N_3840);
nand U4696 (N_4696,N_3012,N_573);
xor U4697 (N_4697,N_3937,N_2745);
nor U4698 (N_4698,N_570,N_2361);
nor U4699 (N_4699,N_1624,N_3692);
nand U4700 (N_4700,N_682,N_1419);
xnor U4701 (N_4701,N_1982,N_2486);
nand U4702 (N_4702,N_127,N_3123);
nand U4703 (N_4703,N_407,N_3141);
or U4704 (N_4704,N_1066,N_90);
nor U4705 (N_4705,N_1203,N_3112);
nor U4706 (N_4706,N_185,N_3125);
xor U4707 (N_4707,N_208,N_574);
xnor U4708 (N_4708,N_3143,N_2984);
nor U4709 (N_4709,N_1313,N_854);
and U4710 (N_4710,N_2108,N_3484);
or U4711 (N_4711,N_3214,N_3485);
xor U4712 (N_4712,N_3437,N_1779);
xor U4713 (N_4713,N_976,N_3084);
or U4714 (N_4714,N_2890,N_1179);
or U4715 (N_4715,N_3416,N_2614);
or U4716 (N_4716,N_1525,N_3379);
or U4717 (N_4717,N_251,N_1506);
and U4718 (N_4718,N_590,N_1542);
or U4719 (N_4719,N_2894,N_2749);
and U4720 (N_4720,N_2000,N_1102);
and U4721 (N_4721,N_1186,N_3384);
and U4722 (N_4722,N_3313,N_2196);
or U4723 (N_4723,N_2628,N_412);
or U4724 (N_4724,N_666,N_3794);
or U4725 (N_4725,N_2407,N_3796);
or U4726 (N_4726,N_26,N_1309);
or U4727 (N_4727,N_243,N_1981);
and U4728 (N_4728,N_1652,N_1438);
nand U4729 (N_4729,N_30,N_350);
or U4730 (N_4730,N_1734,N_1964);
and U4731 (N_4731,N_316,N_110);
nand U4732 (N_4732,N_1117,N_2740);
and U4733 (N_4733,N_1002,N_3591);
or U4734 (N_4734,N_454,N_91);
nand U4735 (N_4735,N_1576,N_2990);
and U4736 (N_4736,N_1689,N_1158);
or U4737 (N_4737,N_80,N_1088);
or U4738 (N_4738,N_1825,N_1211);
or U4739 (N_4739,N_537,N_3899);
and U4740 (N_4740,N_3211,N_756);
nor U4741 (N_4741,N_1513,N_1230);
or U4742 (N_4742,N_733,N_758);
or U4743 (N_4743,N_406,N_3351);
or U4744 (N_4744,N_3191,N_857);
nor U4745 (N_4745,N_499,N_2531);
and U4746 (N_4746,N_2044,N_302);
nor U4747 (N_4747,N_433,N_3705);
xor U4748 (N_4748,N_2810,N_1462);
nand U4749 (N_4749,N_2954,N_410);
nand U4750 (N_4750,N_3460,N_2748);
xnor U4751 (N_4751,N_1799,N_311);
xor U4752 (N_4752,N_688,N_2663);
nor U4753 (N_4753,N_565,N_3602);
nand U4754 (N_4754,N_3205,N_1429);
or U4755 (N_4755,N_176,N_3321);
or U4756 (N_4756,N_1716,N_3297);
and U4757 (N_4757,N_523,N_2344);
nor U4758 (N_4758,N_3074,N_188);
and U4759 (N_4759,N_995,N_2763);
and U4760 (N_4760,N_3401,N_2140);
or U4761 (N_4761,N_1904,N_312);
or U4762 (N_4762,N_2435,N_508);
nand U4763 (N_4763,N_3142,N_2792);
xor U4764 (N_4764,N_2530,N_2621);
or U4765 (N_4765,N_1115,N_553);
or U4766 (N_4766,N_403,N_936);
and U4767 (N_4767,N_2073,N_2331);
nor U4768 (N_4768,N_698,N_3746);
nor U4769 (N_4769,N_3030,N_734);
xor U4770 (N_4770,N_3386,N_1026);
nand U4771 (N_4771,N_2549,N_1231);
xor U4772 (N_4772,N_420,N_2432);
nand U4773 (N_4773,N_3067,N_1334);
nor U4774 (N_4774,N_1997,N_1360);
and U4775 (N_4775,N_163,N_2178);
nor U4776 (N_4776,N_3532,N_1503);
and U4777 (N_4777,N_2287,N_3298);
xor U4778 (N_4778,N_3729,N_1917);
nand U4779 (N_4779,N_2032,N_3345);
nand U4780 (N_4780,N_644,N_1295);
nor U4781 (N_4781,N_3128,N_1051);
nand U4782 (N_4782,N_3014,N_1759);
and U4783 (N_4783,N_916,N_2169);
and U4784 (N_4784,N_430,N_3200);
or U4785 (N_4785,N_2225,N_2343);
nand U4786 (N_4786,N_136,N_108);
nand U4787 (N_4787,N_2805,N_2909);
nor U4788 (N_4788,N_3182,N_3836);
or U4789 (N_4789,N_1065,N_3545);
or U4790 (N_4790,N_2571,N_2814);
nor U4791 (N_4791,N_2827,N_1411);
nor U4792 (N_4792,N_2545,N_3396);
and U4793 (N_4793,N_2952,N_3140);
or U4794 (N_4794,N_3612,N_3256);
and U4795 (N_4795,N_1155,N_1142);
nand U4796 (N_4796,N_833,N_1182);
nor U4797 (N_4797,N_266,N_3987);
nor U4798 (N_4798,N_2876,N_1107);
or U4799 (N_4799,N_3576,N_2087);
nand U4800 (N_4800,N_1972,N_2570);
nor U4801 (N_4801,N_3742,N_1040);
nor U4802 (N_4802,N_1263,N_1817);
xor U4803 (N_4803,N_456,N_1204);
nor U4804 (N_4804,N_2920,N_705);
or U4805 (N_4805,N_633,N_3274);
xor U4806 (N_4806,N_2668,N_2084);
nor U4807 (N_4807,N_2561,N_925);
or U4808 (N_4808,N_1118,N_651);
xor U4809 (N_4809,N_2678,N_3893);
xnor U4810 (N_4810,N_604,N_935);
nand U4811 (N_4811,N_609,N_3040);
nand U4812 (N_4812,N_2592,N_59);
nor U4813 (N_4813,N_3957,N_2849);
nand U4814 (N_4814,N_2018,N_3983);
or U4815 (N_4815,N_3353,N_3589);
or U4816 (N_4816,N_2425,N_1633);
and U4817 (N_4817,N_778,N_998);
or U4818 (N_4818,N_3590,N_3064);
and U4819 (N_4819,N_1170,N_1172);
and U4820 (N_4820,N_1539,N_3852);
and U4821 (N_4821,N_1722,N_2109);
xnor U4822 (N_4822,N_1241,N_3861);
nor U4823 (N_4823,N_919,N_64);
nor U4824 (N_4824,N_3287,N_1973);
nor U4825 (N_4825,N_301,N_2822);
or U4826 (N_4826,N_2652,N_2148);
xnor U4827 (N_4827,N_298,N_3642);
or U4828 (N_4828,N_353,N_3711);
nand U4829 (N_4829,N_963,N_3021);
nor U4830 (N_4830,N_3508,N_2752);
nor U4831 (N_4831,N_68,N_2328);
nor U4832 (N_4832,N_2659,N_3305);
nand U4833 (N_4833,N_1731,N_3566);
xor U4834 (N_4834,N_3301,N_956);
nand U4835 (N_4835,N_616,N_3110);
and U4836 (N_4836,N_1754,N_2459);
and U4837 (N_4837,N_323,N_2036);
nor U4838 (N_4838,N_3791,N_2924);
and U4839 (N_4839,N_3839,N_221);
or U4840 (N_4840,N_53,N_2398);
nand U4841 (N_4841,N_2221,N_1342);
nand U4842 (N_4842,N_3120,N_2121);
nand U4843 (N_4843,N_3387,N_2055);
and U4844 (N_4844,N_2270,N_3259);
nor U4845 (N_4845,N_1140,N_2472);
nand U4846 (N_4846,N_1337,N_2099);
or U4847 (N_4847,N_1567,N_775);
and U4848 (N_4848,N_3582,N_1376);
nand U4849 (N_4849,N_3627,N_2962);
and U4850 (N_4850,N_1719,N_109);
nor U4851 (N_4851,N_3208,N_2075);
nor U4852 (N_4852,N_2423,N_767);
nand U4853 (N_4853,N_3688,N_1523);
nand U4854 (N_4854,N_1691,N_917);
nand U4855 (N_4855,N_788,N_2777);
and U4856 (N_4856,N_2771,N_3921);
or U4857 (N_4857,N_3880,N_1084);
nand U4858 (N_4858,N_3694,N_86);
nor U4859 (N_4859,N_2584,N_1619);
and U4860 (N_4860,N_3103,N_281);
nand U4861 (N_4861,N_2062,N_2031);
xor U4862 (N_4862,N_2415,N_3179);
and U4863 (N_4863,N_1357,N_939);
nand U4864 (N_4864,N_3444,N_2590);
nor U4865 (N_4865,N_895,N_831);
nor U4866 (N_4866,N_952,N_106);
nor U4867 (N_4867,N_2861,N_1956);
nor U4868 (N_4868,N_1449,N_3907);
nand U4869 (N_4869,N_2898,N_2291);
nor U4870 (N_4870,N_944,N_1192);
or U4871 (N_4871,N_147,N_2704);
and U4872 (N_4872,N_3537,N_3108);
nand U4873 (N_4873,N_1775,N_2997);
or U4874 (N_4874,N_2023,N_3022);
nor U4875 (N_4875,N_239,N_2941);
nand U4876 (N_4876,N_2139,N_1191);
and U4877 (N_4877,N_910,N_3469);
nor U4878 (N_4878,N_502,N_3708);
and U4879 (N_4879,N_591,N_409);
nor U4880 (N_4880,N_838,N_3306);
nand U4881 (N_4881,N_1125,N_3463);
xor U4882 (N_4882,N_1234,N_903);
or U4883 (N_4883,N_1048,N_1686);
nand U4884 (N_4884,N_2228,N_498);
nor U4885 (N_4885,N_719,N_196);
or U4886 (N_4886,N_3939,N_548);
and U4887 (N_4887,N_1266,N_3443);
nor U4888 (N_4888,N_1007,N_2747);
xnor U4889 (N_4889,N_583,N_1884);
or U4890 (N_4890,N_2323,N_3497);
or U4891 (N_4891,N_3942,N_1199);
nand U4892 (N_4892,N_2508,N_1519);
nor U4893 (N_4893,N_2161,N_2943);
nor U4894 (N_4894,N_1694,N_1144);
nor U4895 (N_4895,N_814,N_1940);
xnor U4896 (N_4896,N_3455,N_1437);
nand U4897 (N_4897,N_3640,N_393);
or U4898 (N_4898,N_3956,N_593);
xor U4899 (N_4899,N_3499,N_1159);
nor U4900 (N_4900,N_3349,N_3091);
or U4901 (N_4901,N_272,N_295);
nand U4902 (N_4902,N_2022,N_347);
and U4903 (N_4903,N_1582,N_3184);
or U4904 (N_4904,N_620,N_1071);
nand U4905 (N_4905,N_1081,N_1645);
nand U4906 (N_4906,N_3568,N_375);
nor U4907 (N_4907,N_3515,N_2020);
and U4908 (N_4908,N_1011,N_1671);
nor U4909 (N_4909,N_3687,N_3734);
nor U4910 (N_4910,N_2743,N_2625);
nand U4911 (N_4911,N_3474,N_3033);
nor U4912 (N_4912,N_1137,N_2655);
and U4913 (N_4913,N_2298,N_3604);
nor U4914 (N_4914,N_19,N_2734);
nand U4915 (N_4915,N_3847,N_3754);
nor U4916 (N_4916,N_2013,N_799);
and U4917 (N_4917,N_1246,N_95);
or U4918 (N_4918,N_864,N_2123);
nand U4919 (N_4919,N_2841,N_1147);
and U4920 (N_4920,N_2030,N_1888);
nor U4921 (N_4921,N_1661,N_3831);
and U4922 (N_4922,N_1915,N_3704);
nor U4923 (N_4923,N_536,N_1879);
and U4924 (N_4924,N_3772,N_1165);
and U4925 (N_4925,N_3458,N_2832);
xnor U4926 (N_4926,N_2424,N_2275);
nand U4927 (N_4927,N_1156,N_1152);
and U4928 (N_4928,N_2551,N_1847);
or U4929 (N_4929,N_1625,N_2803);
and U4930 (N_4930,N_1143,N_2977);
nand U4931 (N_4931,N_2850,N_3960);
xor U4932 (N_4932,N_798,N_2936);
nor U4933 (N_4933,N_764,N_696);
nor U4934 (N_4934,N_3557,N_70);
nor U4935 (N_4935,N_2892,N_568);
or U4936 (N_4936,N_2669,N_2925);
or U4937 (N_4937,N_2699,N_3233);
xnor U4938 (N_4938,N_1485,N_3412);
xnor U4939 (N_4939,N_1656,N_1397);
or U4940 (N_4940,N_826,N_1750);
nand U4941 (N_4941,N_2811,N_3433);
or U4942 (N_4942,N_215,N_673);
nor U4943 (N_4943,N_3333,N_3482);
nand U4944 (N_4944,N_2579,N_3055);
nor U4945 (N_4945,N_2573,N_1166);
and U4946 (N_4946,N_1067,N_290);
nand U4947 (N_4947,N_3002,N_2598);
and U4948 (N_4948,N_1486,N_983);
nand U4949 (N_4949,N_2061,N_1911);
nand U4950 (N_4950,N_1307,N_2456);
or U4951 (N_4951,N_1814,N_873);
and U4952 (N_4952,N_3432,N_3851);
xnor U4953 (N_4953,N_397,N_3323);
nand U4954 (N_4954,N_1255,N_3773);
nand U4955 (N_4955,N_2587,N_2373);
nand U4956 (N_4956,N_33,N_2948);
nor U4957 (N_4957,N_3393,N_1340);
nor U4958 (N_4958,N_905,N_3774);
xnor U4959 (N_4959,N_820,N_3188);
and U4960 (N_4960,N_1966,N_362);
nand U4961 (N_4961,N_582,N_634);
nor U4962 (N_4962,N_3213,N_1690);
or U4963 (N_4963,N_3808,N_346);
nand U4964 (N_4964,N_1306,N_3519);
nand U4965 (N_4965,N_2434,N_1436);
nor U4966 (N_4966,N_1961,N_3556);
or U4967 (N_4967,N_178,N_2497);
xor U4968 (N_4968,N_2660,N_3368);
nand U4969 (N_4969,N_2431,N_3882);
nor U4970 (N_4970,N_1316,N_779);
nor U4971 (N_4971,N_1196,N_973);
xor U4972 (N_4972,N_1082,N_2759);
nor U4973 (N_4973,N_2290,N_43);
nor U4974 (N_4974,N_763,N_1766);
or U4975 (N_4975,N_3824,N_3465);
or U4976 (N_4976,N_3178,N_3996);
nor U4977 (N_4977,N_2964,N_1920);
and U4978 (N_4978,N_1769,N_1758);
nor U4979 (N_4979,N_793,N_2993);
or U4980 (N_4980,N_1277,N_715);
xnor U4981 (N_4981,N_2007,N_834);
nor U4982 (N_4982,N_1909,N_1070);
nor U4983 (N_4983,N_3183,N_1010);
nor U4984 (N_4984,N_3661,N_1406);
and U4985 (N_4985,N_101,N_2438);
nand U4986 (N_4986,N_160,N_3644);
and U4987 (N_4987,N_3903,N_2313);
or U4988 (N_4988,N_3833,N_2107);
nand U4989 (N_4989,N_1693,N_2603);
nor U4990 (N_4990,N_3529,N_141);
nor U4991 (N_4991,N_2931,N_2848);
xor U4992 (N_4992,N_2441,N_2873);
and U4993 (N_4993,N_1684,N_1768);
and U4994 (N_4994,N_3380,N_2710);
and U4995 (N_4995,N_3007,N_3199);
and U4996 (N_4996,N_676,N_1673);
or U4997 (N_4997,N_1477,N_307);
nor U4998 (N_4998,N_3389,N_3741);
nor U4999 (N_4999,N_1383,N_3862);
nand U5000 (N_5000,N_870,N_3606);
xnor U5001 (N_5001,N_2200,N_3805);
nand U5002 (N_5002,N_3281,N_1394);
and U5003 (N_5003,N_2489,N_1116);
and U5004 (N_5004,N_3028,N_3102);
nor U5005 (N_5005,N_3229,N_1046);
nand U5006 (N_5006,N_3240,N_1188);
or U5007 (N_5007,N_3453,N_949);
or U5008 (N_5008,N_447,N_1780);
xnor U5009 (N_5009,N_337,N_3853);
nor U5010 (N_5010,N_3350,N_2707);
or U5011 (N_5011,N_3000,N_2165);
nor U5012 (N_5012,N_3212,N_599);
nand U5013 (N_5013,N_3902,N_1000);
xnor U5014 (N_5014,N_1355,N_3980);
or U5015 (N_5015,N_2583,N_2643);
or U5016 (N_5016,N_892,N_1929);
and U5017 (N_5017,N_2302,N_2619);
or U5018 (N_5018,N_2586,N_3868);
nand U5019 (N_5019,N_426,N_941);
nand U5020 (N_5020,N_1833,N_1318);
nor U5021 (N_5021,N_635,N_653);
and U5022 (N_5022,N_28,N_937);
and U5023 (N_5023,N_850,N_3020);
nor U5024 (N_5024,N_3347,N_2479);
nor U5025 (N_5025,N_685,N_652);
nand U5026 (N_5026,N_3737,N_631);
nand U5027 (N_5027,N_2199,N_950);
nor U5028 (N_5028,N_1551,N_3282);
or U5029 (N_5029,N_305,N_3053);
nand U5030 (N_5030,N_3629,N_331);
nor U5031 (N_5031,N_3299,N_1032);
and U5032 (N_5032,N_3263,N_874);
and U5033 (N_5033,N_370,N_2033);
or U5034 (N_5034,N_2491,N_3633);
and U5035 (N_5035,N_2517,N_303);
and U5036 (N_5036,N_871,N_341);
and U5037 (N_5037,N_1803,N_3154);
or U5038 (N_5038,N_2079,N_1339);
or U5039 (N_5039,N_968,N_774);
xnor U5040 (N_5040,N_37,N_385);
or U5041 (N_5041,N_2074,N_3330);
and U5042 (N_5042,N_832,N_2511);
nor U5043 (N_5043,N_3447,N_332);
and U5044 (N_5044,N_3357,N_1565);
nand U5045 (N_5045,N_961,N_3998);
nor U5046 (N_5046,N_667,N_875);
and U5047 (N_5047,N_557,N_48);
or U5048 (N_5048,N_1162,N_2038);
nand U5049 (N_5049,N_2681,N_1659);
nor U5050 (N_5050,N_152,N_277);
xnor U5051 (N_5051,N_2008,N_1611);
nand U5052 (N_5052,N_1023,N_3654);
or U5053 (N_5053,N_2244,N_2601);
xor U5054 (N_5054,N_1080,N_986);
and U5055 (N_5055,N_1335,N_2035);
and U5056 (N_5056,N_2906,N_1900);
nor U5057 (N_5057,N_1425,N_993);
nor U5058 (N_5058,N_3992,N_3886);
and U5059 (N_5059,N_2809,N_3516);
nand U5060 (N_5060,N_3061,N_1781);
and U5061 (N_5061,N_1108,N_2011);
or U5062 (N_5062,N_3492,N_1267);
nand U5063 (N_5063,N_3136,N_1695);
nor U5064 (N_5064,N_1830,N_771);
xor U5065 (N_5065,N_796,N_1581);
or U5066 (N_5066,N_2940,N_1370);
and U5067 (N_5067,N_586,N_982);
nor U5068 (N_5068,N_3934,N_547);
nand U5069 (N_5069,N_3870,N_3225);
and U5070 (N_5070,N_2069,N_510);
xnor U5071 (N_5071,N_3725,N_205);
xor U5072 (N_5072,N_1872,N_2034);
and U5073 (N_5073,N_1495,N_2089);
or U5074 (N_5074,N_481,N_1955);
nor U5075 (N_5075,N_528,N_149);
nand U5076 (N_5076,N_1953,N_1606);
or U5077 (N_5077,N_367,N_2368);
nand U5078 (N_5078,N_2778,N_3335);
nor U5079 (N_5079,N_1105,N_2982);
nor U5080 (N_5080,N_167,N_1949);
and U5081 (N_5081,N_742,N_1505);
nor U5082 (N_5082,N_2009,N_1594);
or U5083 (N_5083,N_2005,N_3145);
or U5084 (N_5084,N_340,N_3230);
and U5085 (N_5085,N_293,N_3723);
xnor U5086 (N_5086,N_2447,N_3967);
and U5087 (N_5087,N_16,N_612);
nand U5088 (N_5088,N_790,N_252);
nor U5089 (N_5089,N_3914,N_1446);
nand U5090 (N_5090,N_2644,N_3562);
nor U5091 (N_5091,N_2017,N_1422);
and U5092 (N_5092,N_3314,N_1869);
or U5093 (N_5093,N_361,N_2857);
or U5094 (N_5094,N_2207,N_3867);
nand U5095 (N_5095,N_1016,N_50);
nand U5096 (N_5096,N_3731,N_3665);
nor U5097 (N_5097,N_2632,N_3823);
xor U5098 (N_5098,N_1053,N_1367);
nand U5099 (N_5099,N_3332,N_2507);
nand U5100 (N_5100,N_3925,N_2124);
nand U5101 (N_5101,N_422,N_2218);
and U5102 (N_5102,N_1715,N_3394);
nor U5103 (N_5103,N_1751,N_2247);
nor U5104 (N_5104,N_2101,N_2451);
or U5105 (N_5105,N_1213,N_3189);
or U5106 (N_5106,N_1308,N_317);
or U5107 (N_5107,N_3275,N_3828);
nand U5108 (N_5108,N_929,N_2705);
nand U5109 (N_5109,N_726,N_1753);
nand U5110 (N_5110,N_3162,N_3800);
and U5111 (N_5111,N_1877,N_428);
or U5112 (N_5112,N_1483,N_3546);
nor U5113 (N_5113,N_1420,N_3860);
or U5114 (N_5114,N_1704,N_744);
or U5115 (N_5115,N_2634,N_3410);
nor U5116 (N_5116,N_3371,N_2670);
and U5117 (N_5117,N_3115,N_3094);
nor U5118 (N_5118,N_1922,N_2482);
or U5119 (N_5119,N_572,N_3885);
and U5120 (N_5120,N_3016,N_3649);
and U5121 (N_5121,N_2157,N_2320);
and U5122 (N_5122,N_624,N_3122);
and U5123 (N_5123,N_1176,N_164);
xnor U5124 (N_5124,N_2887,N_3346);
or U5125 (N_5125,N_2054,N_1718);
nand U5126 (N_5126,N_473,N_1852);
and U5127 (N_5127,N_2895,N_921);
and U5128 (N_5128,N_1039,N_3874);
or U5129 (N_5129,N_460,N_1198);
and U5130 (N_5130,N_2515,N_2397);
nor U5131 (N_5131,N_2305,N_846);
or U5132 (N_5132,N_1629,N_1375);
nor U5133 (N_5133,N_3475,N_2334);
or U5134 (N_5134,N_2041,N_1622);
nor U5135 (N_5135,N_278,N_382);
nand U5136 (N_5136,N_1878,N_1338);
and U5137 (N_5137,N_3834,N_2859);
xnor U5138 (N_5138,N_356,N_3626);
or U5139 (N_5139,N_750,N_762);
xnor U5140 (N_5140,N_3502,N_2367);
nand U5141 (N_5141,N_1597,N_1520);
and U5142 (N_5142,N_184,N_3442);
nor U5143 (N_5143,N_3873,N_249);
nand U5144 (N_5144,N_3486,N_2006);
and U5145 (N_5145,N_496,N_1938);
nor U5146 (N_5146,N_1465,N_2610);
or U5147 (N_5147,N_614,N_3950);
nand U5148 (N_5148,N_424,N_2125);
nand U5149 (N_5149,N_2351,N_2389);
xor U5150 (N_5150,N_2716,N_98);
nand U5151 (N_5151,N_894,N_99);
or U5152 (N_5152,N_2289,N_3607);
nand U5153 (N_5153,N_2477,N_1921);
nor U5154 (N_5154,N_2520,N_2421);
and U5155 (N_5155,N_1924,N_2521);
nor U5156 (N_5156,N_752,N_391);
or U5157 (N_5157,N_2260,N_3783);
and U5158 (N_5158,N_2604,N_996);
nand U5159 (N_5159,N_3908,N_2224);
and U5160 (N_5160,N_817,N_2369);
nand U5161 (N_5161,N_1992,N_1478);
and U5162 (N_5162,N_285,N_1942);
xor U5163 (N_5163,N_2560,N_254);
or U5164 (N_5164,N_3740,N_2111);
and U5165 (N_5165,N_464,N_859);
xor U5166 (N_5166,N_533,N_2284);
nor U5167 (N_5167,N_2845,N_3750);
nand U5168 (N_5168,N_1537,N_3395);
nand U5169 (N_5169,N_212,N_1089);
nand U5170 (N_5170,N_1344,N_3242);
nand U5171 (N_5171,N_1918,N_327);
and U5172 (N_5172,N_79,N_2662);
and U5173 (N_5173,N_1498,N_3585);
and U5174 (N_5174,N_1798,N_2058);
nand U5175 (N_5175,N_1489,N_227);
nor U5176 (N_5176,N_2881,N_2880);
and U5177 (N_5177,N_2753,N_1257);
nand U5178 (N_5178,N_2875,N_2339);
nor U5179 (N_5179,N_1093,N_2563);
nor U5180 (N_5180,N_3701,N_1880);
nor U5181 (N_5181,N_3339,N_801);
or U5182 (N_5182,N_2960,N_2744);
nand U5183 (N_5183,N_979,N_915);
nor U5184 (N_5184,N_3488,N_3466);
and U5185 (N_5185,N_3608,N_2466);
xor U5186 (N_5186,N_2250,N_1908);
or U5187 (N_5187,N_663,N_1310);
nand U5188 (N_5188,N_2891,N_1373);
nand U5189 (N_5189,N_1562,N_1504);
or U5190 (N_5190,N_3869,N_2256);
nor U5191 (N_5191,N_2216,N_83);
and U5192 (N_5192,N_2142,N_1358);
nand U5193 (N_5193,N_2156,N_1445);
nand U5194 (N_5194,N_475,N_41);
or U5195 (N_5195,N_539,N_1041);
nand U5196 (N_5196,N_1493,N_1821);
nor U5197 (N_5197,N_2335,N_3080);
nand U5198 (N_5198,N_82,N_3446);
and U5199 (N_5199,N_1368,N_2789);
or U5200 (N_5200,N_2442,N_1514);
or U5201 (N_5201,N_566,N_1593);
nor U5202 (N_5202,N_3245,N_144);
nand U5203 (N_5203,N_1532,N_3736);
xnor U5204 (N_5204,N_3414,N_970);
nand U5205 (N_5205,N_2635,N_2281);
nor U5206 (N_5206,N_1018,N_3320);
nand U5207 (N_5207,N_955,N_199);
xor U5208 (N_5208,N_3542,N_2208);
or U5209 (N_5209,N_2198,N_2819);
or U5210 (N_5210,N_3844,N_975);
nand U5211 (N_5211,N_3709,N_2273);
nand U5212 (N_5212,N_487,N_1044);
nor U5213 (N_5213,N_3954,N_1843);
nor U5214 (N_5214,N_3634,N_1359);
nand U5215 (N_5215,N_235,N_2698);
nand U5216 (N_5216,N_1648,N_2862);
or U5217 (N_5217,N_138,N_1468);
xnor U5218 (N_5218,N_2815,N_29);
nor U5219 (N_5219,N_564,N_678);
and U5220 (N_5220,N_1013,N_2348);
nor U5221 (N_5221,N_2151,N_2572);
or U5222 (N_5222,N_2544,N_1579);
and U5223 (N_5223,N_1710,N_2481);
or U5224 (N_5224,N_640,N_541);
or U5225 (N_5225,N_1735,N_2996);
and U5226 (N_5226,N_434,N_1402);
nor U5227 (N_5227,N_2684,N_112);
nand U5228 (N_5228,N_2942,N_700);
nor U5229 (N_5229,N_3804,N_2687);
xnor U5230 (N_5230,N_3935,N_321);
nand U5231 (N_5231,N_271,N_1205);
or U5232 (N_5232,N_1508,N_782);
nor U5233 (N_5233,N_602,N_1886);
nor U5234 (N_5234,N_3827,N_3429);
nand U5235 (N_5235,N_1232,N_704);
and U5236 (N_5236,N_3423,N_3678);
nor U5237 (N_5237,N_1782,N_1885);
xor U5238 (N_5238,N_3406,N_1558);
nand U5239 (N_5239,N_2197,N_2310);
xnor U5240 (N_5240,N_2137,N_3658);
nor U5241 (N_5241,N_3768,N_1212);
xnor U5242 (N_5242,N_1240,N_128);
nand U5243 (N_5243,N_3344,N_3728);
or U5244 (N_5244,N_1975,N_3512);
xor U5245 (N_5245,N_3160,N_3236);
and U5246 (N_5246,N_2528,N_841);
nor U5247 (N_5247,N_3547,N_279);
nand U5248 (N_5248,N_2577,N_1006);
xor U5249 (N_5249,N_3388,N_1464);
and U5250 (N_5250,N_3922,N_1720);
xnor U5251 (N_5251,N_1839,N_3308);
nor U5252 (N_5252,N_408,N_554);
or U5253 (N_5253,N_1763,N_1602);
nor U5254 (N_5254,N_56,N_1079);
nand U5255 (N_5255,N_2796,N_3289);
or U5256 (N_5256,N_625,N_3718);
and U5257 (N_5257,N_1085,N_241);
and U5258 (N_5258,N_3400,N_275);
nor U5259 (N_5259,N_3181,N_398);
xor U5260 (N_5260,N_2418,N_2661);
nand U5261 (N_5261,N_2269,N_2708);
nor U5262 (N_5262,N_1854,N_3294);
nand U5263 (N_5263,N_766,N_2449);
nand U5264 (N_5264,N_1249,N_3577);
nor U5265 (N_5265,N_713,N_1189);
and U5266 (N_5266,N_3276,N_1764);
and U5267 (N_5267,N_3328,N_3450);
and U5268 (N_5268,N_2359,N_3153);
nand U5269 (N_5269,N_3192,N_1855);
or U5270 (N_5270,N_283,N_1297);
and U5271 (N_5271,N_121,N_1623);
nor U5272 (N_5272,N_2953,N_1012);
and U5273 (N_5273,N_1653,N_2683);
nor U5274 (N_5274,N_40,N_1643);
nand U5275 (N_5275,N_884,N_1314);
or U5276 (N_5276,N_1434,N_1502);
nor U5277 (N_5277,N_1795,N_2736);
or U5278 (N_5278,N_664,N_3500);
and U5279 (N_5279,N_3752,N_1260);
and U5280 (N_5280,N_3336,N_2826);
xor U5281 (N_5281,N_130,N_2717);
or U5282 (N_5282,N_3553,N_610);
nand U5283 (N_5283,N_2835,N_3173);
nor U5284 (N_5284,N_1320,N_1818);
or U5285 (N_5285,N_1999,N_989);
nand U5286 (N_5286,N_2965,N_118);
nand U5287 (N_5287,N_1169,N_2927);
or U5288 (N_5288,N_1746,N_1654);
nand U5289 (N_5289,N_3933,N_495);
and U5290 (N_5290,N_1771,N_2237);
xor U5291 (N_5291,N_1895,N_1761);
xnor U5292 (N_5292,N_3872,N_1741);
nand U5293 (N_5293,N_503,N_525);
nand U5294 (N_5294,N_1242,N_1784);
nand U5295 (N_5295,N_3472,N_613);
nor U5296 (N_5296,N_2309,N_2112);
nor U5297 (N_5297,N_3228,N_868);
and U5298 (N_5298,N_1948,N_1459);
and U5299 (N_5299,N_2401,N_759);
xor U5300 (N_5300,N_1668,N_2781);
or U5301 (N_5301,N_3203,N_3790);
or U5302 (N_5302,N_515,N_3241);
nand U5303 (N_5303,N_1364,N_2626);
or U5304 (N_5304,N_1054,N_1747);
xnor U5305 (N_5305,N_450,N_3916);
and U5306 (N_5306,N_1331,N_2944);
or U5307 (N_5307,N_2483,N_20);
nor U5308 (N_5308,N_3337,N_630);
nand U5309 (N_5309,N_2779,N_3471);
nor U5310 (N_5310,N_1298,N_111);
nor U5311 (N_5311,N_18,N_2585);
or U5312 (N_5312,N_253,N_1253);
and U5313 (N_5313,N_1663,N_738);
xnor U5314 (N_5314,N_13,N_2640);
and U5315 (N_5315,N_601,N_401);
and U5316 (N_5316,N_839,N_3041);
xor U5317 (N_5317,N_913,N_2382);
and U5318 (N_5318,N_2143,N_703);
or U5319 (N_5319,N_383,N_2299);
and U5320 (N_5320,N_2968,N_3479);
nand U5321 (N_5321,N_384,N_3464);
nor U5322 (N_5322,N_2761,N_3419);
or U5323 (N_5323,N_2128,N_17);
nand U5324 (N_5324,N_729,N_2783);
or U5325 (N_5325,N_3864,N_677);
and U5326 (N_5326,N_3365,N_3408);
and U5327 (N_5327,N_806,N_378);
nand U5328 (N_5328,N_876,N_2676);
nand U5329 (N_5329,N_3784,N_3358);
nor U5330 (N_5330,N_2806,N_377);
or U5331 (N_5331,N_1792,N_1995);
and U5332 (N_5332,N_898,N_2677);
and U5333 (N_5333,N_3487,N_2591);
or U5334 (N_5334,N_66,N_3054);
nor U5335 (N_5335,N_1415,N_3316);
nand U5336 (N_5336,N_1187,N_1991);
nor U5337 (N_5337,N_1812,N_3919);
or U5338 (N_5338,N_1778,N_1440);
or U5339 (N_5339,N_1730,N_529);
nand U5340 (N_5340,N_595,N_2868);
nor U5341 (N_5341,N_1271,N_2063);
xnor U5342 (N_5342,N_288,N_1106);
nor U5343 (N_5343,N_2019,N_2129);
nand U5344 (N_5344,N_3072,N_2153);
and U5345 (N_5345,N_3293,N_1469);
nor U5346 (N_5346,N_3894,N_3758);
or U5347 (N_5347,N_594,N_3137);
nor U5348 (N_5348,N_3550,N_3139);
nor U5349 (N_5349,N_2408,N_3158);
nor U5350 (N_5350,N_3671,N_452);
and U5351 (N_5351,N_1181,N_2226);
and U5352 (N_5352,N_3185,N_3264);
nor U5353 (N_5353,N_3097,N_3744);
nor U5354 (N_5354,N_1723,N_1390);
nor U5355 (N_5355,N_3013,N_1632);
nand U5356 (N_5356,N_3325,N_3175);
nor U5357 (N_5357,N_1003,N_3340);
and U5358 (N_5358,N_3329,N_2117);
nor U5359 (N_5359,N_2209,N_23);
nor U5360 (N_5360,N_2122,N_229);
nor U5361 (N_5361,N_3319,N_3363);
nand U5362 (N_5362,N_3303,N_2702);
xnor U5363 (N_5363,N_3690,N_718);
or U5364 (N_5364,N_1609,N_240);
nand U5365 (N_5365,N_546,N_575);
or U5366 (N_5366,N_1481,N_1804);
and U5367 (N_5367,N_2624,N_562);
xor U5368 (N_5368,N_62,N_1461);
nand U5369 (N_5369,N_0,N_484);
xor U5370 (N_5370,N_1391,N_1148);
xor U5371 (N_5371,N_3620,N_1190);
and U5372 (N_5372,N_723,N_1272);
and U5373 (N_5373,N_1119,N_3250);
nand U5374 (N_5374,N_339,N_714);
nor U5375 (N_5375,N_463,N_1019);
or U5376 (N_5376,N_3681,N_2144);
and U5377 (N_5377,N_2258,N_2003);
xnor U5378 (N_5378,N_2537,N_3170);
nand U5379 (N_5379,N_2282,N_1398);
nor U5380 (N_5380,N_1294,N_3930);
xor U5381 (N_5381,N_3748,N_289);
nand U5382 (N_5382,N_3355,N_2040);
nand U5383 (N_5383,N_1736,N_3081);
and U5384 (N_5384,N_3676,N_3441);
or U5385 (N_5385,N_437,N_1866);
nor U5386 (N_5386,N_3812,N_2650);
and U5387 (N_5387,N_2469,N_2812);
nor U5388 (N_5388,N_1252,N_104);
and U5389 (N_5389,N_2461,N_1171);
and U5390 (N_5390,N_2349,N_1030);
nand U5391 (N_5391,N_2506,N_1998);
nand U5392 (N_5392,N_2780,N_1456);
or U5393 (N_5393,N_3404,N_804);
or U5394 (N_5394,N_918,N_878);
or U5395 (N_5395,N_928,N_2616);
and U5396 (N_5396,N_194,N_3771);
and U5397 (N_5397,N_2937,N_2703);
nor U5398 (N_5398,N_2760,N_2476);
nand U5399 (N_5399,N_2319,N_1015);
or U5400 (N_5400,N_3017,N_2210);
nand U5401 (N_5401,N_247,N_3005);
nand U5402 (N_5402,N_172,N_1466);
nand U5403 (N_5403,N_1418,N_306);
or U5404 (N_5404,N_3129,N_441);
or U5405 (N_5405,N_3031,N_246);
or U5406 (N_5406,N_1180,N_2464);
and U5407 (N_5407,N_394,N_3459);
nand U5408 (N_5408,N_2607,N_1153);
or U5409 (N_5409,N_1994,N_1378);
nor U5410 (N_5410,N_803,N_648);
nor U5411 (N_5411,N_1944,N_3969);
or U5412 (N_5412,N_1791,N_2027);
nand U5413 (N_5413,N_3707,N_3176);
nand U5414 (N_5414,N_1748,N_1851);
and U5415 (N_5415,N_3144,N_9);
and U5416 (N_5416,N_1175,N_3477);
and U5417 (N_5417,N_2975,N_345);
nor U5418 (N_5418,N_2526,N_855);
or U5419 (N_5419,N_1708,N_1029);
nand U5420 (N_5420,N_818,N_1925);
xor U5421 (N_5421,N_660,N_2097);
nor U5422 (N_5422,N_2376,N_1952);
nand U5423 (N_5423,N_3424,N_2882);
nor U5424 (N_5424,N_2793,N_3042);
and U5425 (N_5425,N_2512,N_1575);
or U5426 (N_5426,N_580,N_3984);
xnor U5427 (N_5427,N_2615,N_92);
or U5428 (N_5428,N_641,N_2133);
xnor U5429 (N_5429,N_3377,N_3383);
or U5430 (N_5430,N_1490,N_349);
nor U5431 (N_5431,N_15,N_844);
and U5432 (N_5432,N_2304,N_2980);
or U5433 (N_5433,N_2215,N_1556);
nor U5434 (N_5434,N_380,N_3164);
or U5435 (N_5435,N_1250,N_3724);
nand U5436 (N_5436,N_2100,N_1410);
or U5437 (N_5437,N_3948,N_530);
nand U5438 (N_5438,N_3232,N_3260);
nand U5439 (N_5439,N_1554,N_737);
or U5440 (N_5440,N_2562,N_3507);
or U5441 (N_5441,N_1841,N_2646);
nand U5442 (N_5442,N_443,N_3782);
or U5443 (N_5443,N_1214,N_3955);
nor U5444 (N_5444,N_531,N_1634);
nor U5445 (N_5445,N_2065,N_494);
and U5446 (N_5446,N_1849,N_207);
xnor U5447 (N_5447,N_1296,N_1341);
or U5448 (N_5448,N_2393,N_1280);
or U5449 (N_5449,N_2217,N_768);
or U5450 (N_5450,N_1057,N_3845);
and U5451 (N_5451,N_3900,N_5);
nor U5452 (N_5452,N_1330,N_2620);
nand U5453 (N_5453,N_468,N_1482);
nor U5454 (N_5454,N_3234,N_2001);
xnor U5455 (N_5455,N_1574,N_25);
nor U5456 (N_5456,N_3057,N_3352);
nand U5457 (N_5457,N_3897,N_3390);
xor U5458 (N_5458,N_156,N_2503);
nor U5459 (N_5459,N_3891,N_3326);
nor U5460 (N_5460,N_984,N_493);
and U5461 (N_5461,N_1870,N_1549);
nor U5462 (N_5462,N_2242,N_1980);
nor U5463 (N_5463,N_3503,N_848);
and U5464 (N_5464,N_772,N_1409);
or U5465 (N_5465,N_1238,N_120);
and U5466 (N_5466,N_1604,N_259);
nor U5467 (N_5467,N_735,N_2251);
or U5468 (N_5468,N_1696,N_2039);
or U5469 (N_5469,N_2233,N_3637);
nand U5470 (N_5470,N_3180,N_2800);
and U5471 (N_5471,N_722,N_2149);
or U5472 (N_5472,N_3106,N_190);
nor U5473 (N_5473,N_934,N_372);
xnor U5474 (N_5474,N_1300,N_1164);
and U5475 (N_5475,N_645,N_3563);
or U5476 (N_5476,N_3063,N_1617);
nor U5477 (N_5477,N_418,N_1756);
nand U5478 (N_5478,N_3918,N_396);
nand U5479 (N_5479,N_2076,N_607);
nor U5480 (N_5480,N_569,N_2916);
nand U5481 (N_5481,N_2878,N_1591);
nor U5482 (N_5482,N_736,N_2321);
and U5483 (N_5483,N_1269,N_3044);
nand U5484 (N_5484,N_2535,N_649);
or U5485 (N_5485,N_3615,N_22);
or U5486 (N_5486,N_1832,N_579);
nand U5487 (N_5487,N_2966,N_2807);
nand U5488 (N_5488,N_3010,N_2578);
and U5489 (N_5489,N_3116,N_78);
nand U5490 (N_5490,N_974,N_1860);
or U5491 (N_5491,N_3753,N_1573);
nand U5492 (N_5492,N_1317,N_755);
and U5493 (N_5493,N_2429,N_3898);
nor U5494 (N_5494,N_1274,N_1408);
nand U5495 (N_5495,N_3490,N_1725);
and U5496 (N_5496,N_1773,N_578);
nor U5497 (N_5497,N_3302,N_2955);
or U5498 (N_5498,N_1223,N_1626);
or U5499 (N_5499,N_1311,N_2460);
nand U5500 (N_5500,N_2750,N_1561);
nand U5501 (N_5501,N_1428,N_882);
nor U5502 (N_5502,N_1348,N_1974);
nand U5503 (N_5503,N_1631,N_668);
and U5504 (N_5504,N_2279,N_2950);
or U5505 (N_5505,N_2612,N_728);
nand U5506 (N_5506,N_2602,N_2863);
nor U5507 (N_5507,N_113,N_2059);
and U5508 (N_5508,N_3985,N_3628);
or U5509 (N_5509,N_3247,N_3911);
nand U5510 (N_5510,N_702,N_3896);
or U5511 (N_5511,N_488,N_436);
nand U5512 (N_5512,N_2358,N_960);
nor U5513 (N_5513,N_3024,N_2513);
or U5514 (N_5514,N_1835,N_3555);
and U5515 (N_5515,N_2735,N_3926);
nand U5516 (N_5516,N_1497,N_210);
nand U5517 (N_5517,N_658,N_2637);
and U5518 (N_5518,N_598,N_3573);
nand U5519 (N_5519,N_2338,N_3775);
xnor U5520 (N_5520,N_2538,N_897);
and U5521 (N_5521,N_3327,N_890);
and U5522 (N_5522,N_67,N_3146);
xnor U5523 (N_5523,N_2788,N_2173);
nand U5524 (N_5524,N_1047,N_2467);
and U5525 (N_5525,N_3454,N_2274);
nand U5526 (N_5526,N_3246,N_701);
xor U5527 (N_5527,N_3962,N_1132);
and U5528 (N_5528,N_2455,N_2205);
or U5529 (N_5529,N_967,N_228);
nor U5530 (N_5530,N_3762,N_1200);
nor U5531 (N_5531,N_791,N_1001);
or U5532 (N_5532,N_1914,N_2081);
nand U5533 (N_5533,N_3593,N_2554);
or U5534 (N_5534,N_3177,N_490);
nor U5535 (N_5535,N_957,N_881);
or U5536 (N_5536,N_1432,N_3785);
nand U5537 (N_5537,N_3456,N_3525);
nand U5538 (N_5538,N_3699,N_3364);
or U5539 (N_5539,N_3789,N_224);
nand U5540 (N_5540,N_2611,N_2854);
nand U5541 (N_5541,N_749,N_3730);
and U5542 (N_5542,N_1614,N_2641);
or U5543 (N_5543,N_3561,N_717);
and U5544 (N_5544,N_2496,N_1312);
or U5545 (N_5545,N_3359,N_730);
and U5546 (N_5546,N_3391,N_3227);
nand U5547 (N_5547,N_741,N_1229);
or U5548 (N_5548,N_1374,N_325);
or U5549 (N_5549,N_206,N_3121);
or U5550 (N_5550,N_3877,N_1043);
nand U5551 (N_5551,N_1386,N_165);
nand U5552 (N_5552,N_1261,N_3187);
nand U5553 (N_5553,N_6,N_3324);
nor U5554 (N_5554,N_1351,N_2147);
and U5555 (N_5555,N_2114,N_2412);
or U5556 (N_5556,N_543,N_2842);
and U5557 (N_5557,N_159,N_174);
xnor U5558 (N_5558,N_947,N_3430);
nor U5559 (N_5559,N_2645,N_1451);
nand U5560 (N_5560,N_2470,N_3119);
nor U5561 (N_5561,N_3265,N_2741);
and U5562 (N_5562,N_1848,N_815);
nor U5563 (N_5563,N_233,N_3703);
and U5564 (N_5564,N_725,N_2301);
nor U5565 (N_5565,N_2995,N_2160);
and U5566 (N_5566,N_1588,N_3613);
and U5567 (N_5567,N_751,N_2613);
xor U5568 (N_5568,N_3062,N_2772);
nand U5569 (N_5569,N_1674,N_780);
or U5570 (N_5570,N_646,N_2529);
xor U5571 (N_5571,N_748,N_146);
or U5572 (N_5572,N_2387,N_865);
nand U5573 (N_5573,N_3093,N_2350);
nand U5574 (N_5574,N_3635,N_36);
nand U5575 (N_5575,N_97,N_1304);
nor U5576 (N_5576,N_965,N_3047);
nand U5577 (N_5577,N_3913,N_3026);
nor U5578 (N_5578,N_2730,N_1128);
nor U5579 (N_5579,N_1150,N_344);
nand U5580 (N_5580,N_3695,N_416);
and U5581 (N_5581,N_381,N_1025);
or U5582 (N_5582,N_1064,N_1958);
and U5583 (N_5583,N_1688,N_1228);
and U5584 (N_5584,N_77,N_2879);
nand U5585 (N_5585,N_1480,N_3132);
and U5586 (N_5586,N_3099,N_709);
and U5587 (N_5587,N_2897,N_3035);
and U5588 (N_5588,N_1086,N_1901);
nor U5589 (N_5589,N_168,N_2550);
or U5590 (N_5590,N_3415,N_324);
and U5591 (N_5591,N_3198,N_300);
and U5592 (N_5592,N_2630,N_1526);
nor U5593 (N_5593,N_1963,N_258);
or U5594 (N_5594,N_193,N_3272);
and U5595 (N_5595,N_3197,N_3978);
nand U5596 (N_5596,N_3370,N_2769);
or U5597 (N_5597,N_2356,N_3792);
and U5598 (N_5598,N_2693,N_3356);
nand U5599 (N_5599,N_1283,N_3959);
and U5600 (N_5600,N_3936,N_2816);
nand U5601 (N_5601,N_2326,N_922);
nor U5602 (N_5602,N_3207,N_608);
xor U5603 (N_5603,N_761,N_3501);
and U5604 (N_5604,N_1467,N_1709);
nor U5605 (N_5605,N_2083,N_692);
and U5606 (N_5606,N_3765,N_34);
or U5607 (N_5607,N_1063,N_1299);
xnor U5608 (N_5608,N_2159,N_3583);
and U5609 (N_5609,N_2312,N_2390);
or U5610 (N_5610,N_1460,N_1073);
nor U5611 (N_5611,N_544,N_3290);
and U5612 (N_5612,N_1038,N_2776);
nor U5613 (N_5613,N_2337,N_1305);
and U5614 (N_5614,N_3829,N_292);
nor U5615 (N_5615,N_3857,N_2286);
nand U5616 (N_5616,N_1499,N_319);
nand U5617 (N_5617,N_3940,N_1950);
or U5618 (N_5618,N_2582,N_1697);
and U5619 (N_5619,N_2090,N_81);
and U5620 (N_5620,N_1834,N_220);
and U5621 (N_5621,N_621,N_1414);
nor U5622 (N_5622,N_348,N_2002);
nand U5623 (N_5623,N_550,N_2903);
nor U5624 (N_5624,N_1262,N_1536);
or U5625 (N_5625,N_238,N_731);
or U5626 (N_5626,N_1226,N_1572);
or U5627 (N_5627,N_1675,N_218);
and U5628 (N_5628,N_2372,N_2195);
nor U5629 (N_5629,N_1853,N_2116);
and U5630 (N_5630,N_907,N_3915);
or U5631 (N_5631,N_1823,N_1471);
xnor U5632 (N_5632,N_1033,N_3312);
nor U5633 (N_5633,N_2171,N_618);
nor U5634 (N_5634,N_3904,N_1112);
and U5635 (N_5635,N_3971,N_2596);
nand U5636 (N_5636,N_2733,N_3619);
nand U5637 (N_5637,N_1301,N_3565);
or U5638 (N_5638,N_3360,N_1210);
or U5639 (N_5639,N_3315,N_2580);
or U5640 (N_5640,N_585,N_885);
and U5641 (N_5641,N_2162,N_1868);
or U5642 (N_5642,N_3807,N_694);
nor U5643 (N_5643,N_708,N_276);
nand U5644 (N_5644,N_157,N_3641);
nor U5645 (N_5645,N_263,N_3085);
and U5646 (N_5646,N_2719,N_1752);
nor U5647 (N_5647,N_2700,N_3567);
nor U5648 (N_5648,N_162,N_2021);
nand U5649 (N_5649,N_1533,N_2155);
or U5650 (N_5650,N_1247,N_3801);
or U5651 (N_5651,N_2522,N_2010);
and U5652 (N_5652,N_3034,N_231);
nand U5653 (N_5653,N_491,N_3318);
or U5654 (N_5654,N_2050,N_3342);
nand U5655 (N_5655,N_2292,N_2043);
and U5656 (N_5656,N_173,N_3732);
and U5657 (N_5657,N_1021,N_1036);
or U5658 (N_5658,N_2052,N_414);
nor U5659 (N_5659,N_3733,N_1802);
nor U5660 (N_5660,N_255,N_2166);
nand U5661 (N_5661,N_3411,N_3);
xnor U5662 (N_5662,N_1742,N_1258);
or U5663 (N_5663,N_1630,N_945);
or U5664 (N_5664,N_1512,N_1559);
nand U5665 (N_5665,N_1372,N_760);
and U5666 (N_5666,N_1217,N_3973);
or U5667 (N_5667,N_2758,N_2078);
nor U5668 (N_5668,N_816,N_245);
and U5669 (N_5669,N_2498,N_754);
or U5670 (N_5670,N_1254,N_76);
nand U5671 (N_5671,N_3452,N_3514);
or U5672 (N_5672,N_3483,N_1757);
nor U5673 (N_5673,N_3280,N_2967);
nor U5674 (N_5674,N_2152,N_1245);
nand U5675 (N_5675,N_990,N_2642);
and U5676 (N_5676,N_3846,N_2574);
or U5677 (N_5677,N_558,N_1395);
and U5678 (N_5678,N_1407,N_180);
and U5679 (N_5679,N_517,N_1685);
or U5680 (N_5680,N_603,N_1983);
nor U5681 (N_5681,N_2915,N_2327);
and U5682 (N_5682,N_123,N_1785);
or U5683 (N_5683,N_1882,N_3779);
or U5684 (N_5684,N_2266,N_2377);
or U5685 (N_5685,N_3405,N_1239);
or U5686 (N_5686,N_784,N_453);
nor U5687 (N_5687,N_3586,N_1876);
and U5688 (N_5688,N_1049,N_1413);
nor U5689 (N_5689,N_2618,N_1401);
or U5690 (N_5690,N_3693,N_3745);
or U5691 (N_5691,N_2484,N_1728);
and U5692 (N_5692,N_3645,N_2500);
nor U5693 (N_5693,N_3243,N_2896);
nor U5694 (N_5694,N_1811,N_1807);
or U5695 (N_5695,N_1945,N_1474);
nor U5696 (N_5696,N_840,N_3169);
nor U5697 (N_5697,N_3069,N_2494);
nor U5698 (N_5698,N_1244,N_1479);
nor U5699 (N_5699,N_3826,N_2163);
nand U5700 (N_5700,N_1984,N_1889);
and U5701 (N_5701,N_2427,N_862);
and U5702 (N_5702,N_909,N_2737);
and U5703 (N_5703,N_1293,N_1857);
nor U5704 (N_5704,N_294,N_858);
xnor U5705 (N_5705,N_2908,N_1642);
xnor U5706 (N_5706,N_2417,N_1515);
and U5707 (N_5707,N_505,N_3979);
and U5708 (N_5708,N_3296,N_1399);
nor U5709 (N_5709,N_69,N_769);
nand U5710 (N_5710,N_482,N_642);
and U5711 (N_5711,N_3058,N_1916);
nor U5712 (N_5712,N_440,N_3473);
and U5713 (N_5713,N_1423,N_1820);
and U5714 (N_5714,N_326,N_55);
nand U5715 (N_5715,N_477,N_2458);
and U5716 (N_5716,N_856,N_2569);
nand U5717 (N_5717,N_1014,N_2170);
xor U5718 (N_5718,N_3901,N_1679);
or U5719 (N_5719,N_954,N_35);
and U5720 (N_5720,N_1943,N_3609);
nor U5721 (N_5721,N_2480,N_1094);
nand U5722 (N_5722,N_461,N_1657);
nor U5723 (N_5723,N_3098,N_1207);
nand U5724 (N_5724,N_3075,N_1701);
and U5725 (N_5725,N_3759,N_2688);
nor U5726 (N_5726,N_3498,N_2188);
and U5727 (N_5727,N_2119,N_3696);
or U5728 (N_5728,N_1141,N_451);
nor U5729 (N_5729,N_1680,N_1251);
nor U5730 (N_5730,N_518,N_2254);
and U5731 (N_5731,N_577,N_3855);
nand U5732 (N_5732,N_2047,N_3802);
and U5733 (N_5733,N_2132,N_2499);
nand U5734 (N_5734,N_248,N_991);
nand U5735 (N_5735,N_1256,N_3735);
and U5736 (N_5736,N_2505,N_2176);
nor U5737 (N_5737,N_369,N_3317);
nand U5738 (N_5738,N_2118,N_2465);
nor U5739 (N_5739,N_3623,N_805);
or U5740 (N_5740,N_1225,N_617);
or U5741 (N_5741,N_3764,N_1167);
and U5742 (N_5742,N_1237,N_683);
or U5743 (N_5743,N_797,N_1319);
xor U5744 (N_5744,N_3682,N_1416);
nand U5745 (N_5745,N_927,N_2070);
nor U5746 (N_5746,N_2877,N_2502);
nor U5747 (N_5747,N_1744,N_2723);
nor U5748 (N_5748,N_444,N_2120);
and U5749 (N_5749,N_2870,N_419);
nand U5750 (N_5750,N_1099,N_2214);
nor U5751 (N_5751,N_2236,N_2518);
or U5752 (N_5752,N_1134,N_2853);
nor U5753 (N_5753,N_3221,N_3438);
or U5754 (N_5754,N_1721,N_3255);
or U5755 (N_5755,N_923,N_795);
or U5756 (N_5756,N_2471,N_201);
nand U5757 (N_5757,N_2724,N_234);
nor U5758 (N_5758,N_1184,N_1822);
or U5759 (N_5759,N_2303,N_1092);
or U5760 (N_5760,N_1035,N_126);
nor U5761 (N_5761,N_1522,N_1273);
or U5762 (N_5762,N_52,N_1647);
nor U5763 (N_5763,N_143,N_2488);
or U5764 (N_5764,N_1405,N_3947);
xor U5765 (N_5765,N_3856,N_1363);
and U5766 (N_5766,N_2860,N_471);
or U5767 (N_5767,N_3435,N_3795);
or U5768 (N_5768,N_2516,N_3073);
xor U5769 (N_5769,N_2594,N_1353);
nor U5770 (N_5770,N_706,N_821);
or U5771 (N_5771,N_2371,N_1028);
nand U5772 (N_5772,N_3530,N_920);
nor U5773 (N_5773,N_1195,N_2510);
nor U5774 (N_5774,N_3051,N_3811);
nor U5775 (N_5775,N_3958,N_2675);
or U5776 (N_5776,N_2354,N_1131);
and U5777 (N_5777,N_3431,N_1475);
nor U5778 (N_5778,N_1292,N_2939);
or U5779 (N_5779,N_1343,N_3090);
and U5780 (N_5780,N_2622,N_2203);
nor U5781 (N_5781,N_402,N_1457);
or U5782 (N_5782,N_3025,N_520);
nor U5783 (N_5783,N_3217,N_2568);
nand U5784 (N_5784,N_2333,N_3616);
nand U5785 (N_5785,N_1669,N_46);
xnor U5786 (N_5786,N_933,N_2534);
or U5787 (N_5787,N_2296,N_119);
nand U5788 (N_5788,N_509,N_1727);
xnor U5789 (N_5789,N_1126,N_2222);
or U5790 (N_5790,N_236,N_2509);
or U5791 (N_5791,N_2463,N_155);
or U5792 (N_5792,N_689,N_2830);
nand U5793 (N_5793,N_830,N_1183);
and U5794 (N_5794,N_1031,N_721);
nor U5795 (N_5795,N_478,N_2956);
and U5796 (N_5796,N_3647,N_2285);
or U5797 (N_5797,N_1235,N_835);
nand U5798 (N_5798,N_364,N_3505);
or U5799 (N_5799,N_3541,N_842);
and U5800 (N_5800,N_1384,N_777);
or U5801 (N_5801,N_260,N_3206);
and U5802 (N_5802,N_2947,N_589);
nor U5803 (N_5803,N_1894,N_2907);
and U5804 (N_5804,N_3147,N_1577);
nand U5805 (N_5805,N_469,N_1);
and U5806 (N_5806,N_3535,N_2701);
nand U5807 (N_5807,N_2548,N_3104);
nor U5808 (N_5808,N_3271,N_3060);
nand U5809 (N_5809,N_2450,N_3534);
nor U5810 (N_5810,N_3118,N_2355);
or U5811 (N_5811,N_527,N_2448);
and U5812 (N_5812,N_2201,N_262);
or U5813 (N_5813,N_1620,N_3538);
nand U5814 (N_5814,N_1216,N_1455);
nor U5815 (N_5815,N_1545,N_1543);
and U5816 (N_5816,N_559,N_571);
nor U5817 (N_5817,N_71,N_31);
nor U5818 (N_5818,N_1221,N_1077);
and U5819 (N_5819,N_2015,N_2782);
nand U5820 (N_5820,N_1637,N_1636);
or U5821 (N_5821,N_459,N_3592);
or U5822 (N_5822,N_102,N_7);
nor U5823 (N_5823,N_953,N_1706);
or U5824 (N_5824,N_2086,N_3953);
nor U5825 (N_5825,N_1672,N_1544);
and U5826 (N_5826,N_2185,N_1122);
nand U5827 (N_5827,N_2454,N_3895);
or U5828 (N_5828,N_411,N_1789);
and U5829 (N_5829,N_3837,N_3109);
xor U5830 (N_5830,N_2542,N_3884);
nor U5831 (N_5831,N_1427,N_2871);
and U5832 (N_5832,N_906,N_1683);
and U5833 (N_5833,N_1265,N_1442);
nor U5834 (N_5834,N_538,N_825);
nor U5835 (N_5835,N_3698,N_2885);
or U5836 (N_5836,N_39,N_3133);
or U5837 (N_5837,N_3755,N_3392);
nand U5838 (N_5838,N_2820,N_3322);
and U5839 (N_5839,N_3134,N_2533);
and U5840 (N_5840,N_2294,N_3513);
or U5841 (N_5841,N_3224,N_1329);
nand U5842 (N_5842,N_1926,N_3003);
and U5843 (N_5843,N_489,N_2230);
nand U5844 (N_5844,N_2150,N_1069);
or U5845 (N_5845,N_3920,N_3348);
nor U5846 (N_5846,N_3201,N_49);
or U5847 (N_5847,N_770,N_2838);
and U5848 (N_5848,N_1800,N_2278);
or U5849 (N_5849,N_3052,N_131);
or U5850 (N_5850,N_1726,N_1700);
nor U5851 (N_5851,N_3078,N_3928);
or U5852 (N_5852,N_2874,N_845);
xor U5853 (N_5853,N_3632,N_358);
nor U5854 (N_5854,N_3964,N_3662);
nand U5855 (N_5855,N_187,N_1096);
nand U5856 (N_5856,N_540,N_2976);
xnor U5857 (N_5857,N_3130,N_2828);
xnor U5858 (N_5858,N_2248,N_1380);
and U5859 (N_5859,N_3830,N_1055);
nor U5860 (N_5860,N_2689,N_1932);
xnor U5861 (N_5861,N_745,N_3100);
nand U5862 (N_5862,N_3269,N_2416);
nand U5863 (N_5863,N_1387,N_2923);
nand U5864 (N_5864,N_1024,N_1441);
nand U5865 (N_5865,N_3938,N_10);
nor U5866 (N_5866,N_3697,N_1553);
nand U5867 (N_5867,N_3461,N_12);
xor U5868 (N_5868,N_3813,N_1151);
nand U5869 (N_5869,N_1303,N_2492);
or U5870 (N_5870,N_2867,N_3066);
nor U5871 (N_5871,N_3215,N_628);
or U5872 (N_5872,N_695,N_3668);
xor U5873 (N_5873,N_3738,N_38);
xor U5874 (N_5874,N_2028,N_2468);
xnor U5875 (N_5875,N_3559,N_2911);
nor U5876 (N_5876,N_3990,N_3638);
and U5877 (N_5877,N_3601,N_829);
nor U5878 (N_5878,N_2375,N_3216);
nor U5879 (N_5879,N_1215,N_931);
nand U5880 (N_5880,N_2929,N_3621);
and U5881 (N_5881,N_2691,N_154);
nor U5882 (N_5882,N_492,N_636);
nand U5883 (N_5883,N_2600,N_352);
nor U5884 (N_5884,N_89,N_3821);
nand U5885 (N_5885,N_1027,N_988);
nand U5886 (N_5886,N_1639,N_3636);
nor U5887 (N_5887,N_3548,N_1743);
nor U5888 (N_5888,N_3643,N_3076);
or U5889 (N_5889,N_2235,N_1100);
or U5890 (N_5890,N_3113,N_1692);
xnor U5891 (N_5891,N_2742,N_959);
nor U5892 (N_5892,N_429,N_3727);
or U5893 (N_5893,N_142,N_3015);
or U5894 (N_5894,N_58,N_1291);
and U5895 (N_5895,N_3570,N_3580);
nand U5896 (N_5896,N_3193,N_2756);
nor U5897 (N_5897,N_423,N_3706);
nor U5898 (N_5898,N_1146,N_2833);
nor U5899 (N_5899,N_2316,N_14);
and U5900 (N_5900,N_2725,N_691);
and U5901 (N_5901,N_3194,N_1135);
nand U5902 (N_5902,N_2846,N_2384);
and U5903 (N_5903,N_2588,N_1557);
and U5904 (N_5904,N_2068,N_2446);
and U5905 (N_5905,N_3006,N_3526);
nor U5906 (N_5906,N_1154,N_2262);
nand U5907 (N_5907,N_552,N_3004);
nor U5908 (N_5908,N_3674,N_3023);
nor U5909 (N_5909,N_753,N_3560);
or U5910 (N_5910,N_1954,N_3769);
and U5911 (N_5911,N_2721,N_1492);
nand U5912 (N_5912,N_3367,N_3165);
nor U5913 (N_5913,N_1220,N_1538);
xor U5914 (N_5914,N_2174,N_1139);
and U5915 (N_5915,N_3610,N_932);
nand U5916 (N_5916,N_561,N_2308);
and U5917 (N_5917,N_3343,N_1988);
and U5918 (N_5918,N_1518,N_3655);
nor U5919 (N_5919,N_237,N_1173);
nand U5920 (N_5920,N_2785,N_274);
and U5921 (N_5921,N_1935,N_1243);
xnor U5922 (N_5922,N_942,N_1702);
nand U5923 (N_5923,N_687,N_3890);
or U5924 (N_5924,N_3797,N_1516);
and U5925 (N_5925,N_1325,N_3879);
nand U5926 (N_5926,N_786,N_3291);
or U5927 (N_5927,N_522,N_1098);
and U5928 (N_5928,N_2428,N_1202);
or U5929 (N_5929,N_2951,N_462);
xnor U5930 (N_5930,N_3972,N_879);
nor U5931 (N_5931,N_61,N_1863);
and U5932 (N_5932,N_1640,N_1965);
or U5933 (N_5933,N_2933,N_2802);
nand U5934 (N_5934,N_1570,N_2726);
xor U5935 (N_5935,N_3398,N_1168);
and U5936 (N_5936,N_1424,N_1996);
xnor U5937 (N_5937,N_439,N_3273);
and U5938 (N_5938,N_2095,N_549);
and U5939 (N_5939,N_1875,N_3743);
xnor U5940 (N_5940,N_2295,N_3311);
xnor U5941 (N_5941,N_1400,N_1595);
or U5942 (N_5942,N_2899,N_200);
nor U5943 (N_5943,N_669,N_3520);
and U5944 (N_5944,N_3982,N_2910);
nor U5945 (N_5945,N_1248,N_1745);
nand U5946 (N_5946,N_2180,N_555);
and U5947 (N_5947,N_203,N_315);
nor U5948 (N_5948,N_3684,N_3720);
or U5949 (N_5949,N_2872,N_3131);
nand U5950 (N_5950,N_542,N_3403);
nor U5951 (N_5951,N_1681,N_1103);
and U5952 (N_5952,N_485,N_724);
nor U5953 (N_5953,N_1968,N_1649);
nor U5954 (N_5954,N_2567,N_2444);
nor U5955 (N_5955,N_1087,N_827);
nand U5956 (N_5956,N_3039,N_24);
or U5957 (N_5957,N_3809,N_2935);
nor U5958 (N_5958,N_1628,N_2104);
or U5959 (N_5959,N_962,N_3770);
xnor U5960 (N_5960,N_3549,N_2004);
or U5961 (N_5961,N_3832,N_3495);
nor U5962 (N_5962,N_139,N_3927);
and U5963 (N_5963,N_1601,N_2332);
nor U5964 (N_5964,N_2106,N_3257);
or U5965 (N_5965,N_313,N_3528);
nand U5966 (N_5966,N_2764,N_3071);
or U5967 (N_5967,N_1075,N_2738);
nand U5968 (N_5968,N_2636,N_899);
nand U5969 (N_5969,N_1236,N_1603);
or U5970 (N_5970,N_2347,N_869);
or U5971 (N_5971,N_1534,N_2765);
or U5972 (N_5972,N_3717,N_3866);
or U5973 (N_5973,N_3605,N_2364);
nor U5974 (N_5974,N_1072,N_1760);
nand U5975 (N_5975,N_192,N_632);
and U5976 (N_5976,N_2219,N_3757);
nor U5977 (N_5977,N_2440,N_166);
nand U5978 (N_5978,N_3204,N_3544);
and U5979 (N_5979,N_2380,N_526);
or U5980 (N_5980,N_335,N_2317);
and U5981 (N_5981,N_1568,N_3721);
and U5982 (N_5982,N_3810,N_3295);
nor U5983 (N_5983,N_465,N_3540);
nor U5984 (N_5984,N_3491,N_3806);
or U5985 (N_5985,N_2847,N_2799);
or U5986 (N_5986,N_880,N_3043);
nor U5987 (N_5987,N_511,N_2311);
xnor U5988 (N_5988,N_1145,N_1810);
xnor U5989 (N_5989,N_2071,N_3672);
nand U5990 (N_5990,N_3659,N_3399);
nor U5991 (N_5991,N_1856,N_2985);
or U5992 (N_5992,N_2288,N_863);
and U5993 (N_5993,N_1552,N_1149);
nor U5994 (N_5994,N_2255,N_3702);
and U5995 (N_5995,N_2889,N_3101);
or U5996 (N_5996,N_2072,N_310);
or U5997 (N_5997,N_124,N_2060);
or U5998 (N_5998,N_3238,N_3974);
xnor U5999 (N_5999,N_2189,N_3527);
and U6000 (N_6000,N_1292,N_3453);
and U6001 (N_6001,N_3250,N_1231);
nor U6002 (N_6002,N_568,N_3596);
and U6003 (N_6003,N_2773,N_677);
nand U6004 (N_6004,N_31,N_3661);
nand U6005 (N_6005,N_3255,N_2715);
and U6006 (N_6006,N_2656,N_515);
nor U6007 (N_6007,N_3721,N_2928);
nand U6008 (N_6008,N_2031,N_3049);
and U6009 (N_6009,N_1534,N_164);
nor U6010 (N_6010,N_2938,N_2122);
nor U6011 (N_6011,N_3425,N_2262);
nand U6012 (N_6012,N_2604,N_578);
nor U6013 (N_6013,N_3870,N_1243);
or U6014 (N_6014,N_2912,N_144);
xnor U6015 (N_6015,N_639,N_3239);
or U6016 (N_6016,N_3826,N_435);
or U6017 (N_6017,N_1171,N_126);
nand U6018 (N_6018,N_3323,N_1602);
nand U6019 (N_6019,N_2533,N_3697);
nand U6020 (N_6020,N_1740,N_3342);
nor U6021 (N_6021,N_3369,N_3186);
and U6022 (N_6022,N_263,N_699);
and U6023 (N_6023,N_1957,N_2009);
and U6024 (N_6024,N_411,N_1463);
nand U6025 (N_6025,N_957,N_2299);
nand U6026 (N_6026,N_382,N_2784);
xnor U6027 (N_6027,N_2853,N_116);
nor U6028 (N_6028,N_1841,N_1737);
nand U6029 (N_6029,N_1941,N_202);
nand U6030 (N_6030,N_1485,N_740);
xnor U6031 (N_6031,N_3833,N_334);
or U6032 (N_6032,N_3214,N_2315);
nor U6033 (N_6033,N_3152,N_1214);
nand U6034 (N_6034,N_249,N_2915);
nor U6035 (N_6035,N_3146,N_2001);
or U6036 (N_6036,N_1784,N_2087);
xnor U6037 (N_6037,N_3728,N_3719);
nor U6038 (N_6038,N_3553,N_3325);
nor U6039 (N_6039,N_3339,N_2795);
or U6040 (N_6040,N_3747,N_3801);
and U6041 (N_6041,N_2020,N_1351);
or U6042 (N_6042,N_912,N_3100);
xnor U6043 (N_6043,N_3981,N_3249);
nor U6044 (N_6044,N_3812,N_2567);
xor U6045 (N_6045,N_3821,N_1314);
or U6046 (N_6046,N_2874,N_2086);
and U6047 (N_6047,N_3163,N_2454);
nor U6048 (N_6048,N_994,N_1614);
or U6049 (N_6049,N_3103,N_614);
nand U6050 (N_6050,N_3093,N_1854);
and U6051 (N_6051,N_2228,N_1927);
nor U6052 (N_6052,N_3478,N_3627);
xor U6053 (N_6053,N_1818,N_2211);
and U6054 (N_6054,N_3278,N_2609);
nor U6055 (N_6055,N_3964,N_706);
xnor U6056 (N_6056,N_2899,N_3508);
nand U6057 (N_6057,N_1931,N_3746);
nand U6058 (N_6058,N_2489,N_3375);
and U6059 (N_6059,N_2548,N_1565);
xor U6060 (N_6060,N_3346,N_633);
nor U6061 (N_6061,N_3354,N_1417);
and U6062 (N_6062,N_1541,N_970);
and U6063 (N_6063,N_1588,N_1218);
or U6064 (N_6064,N_1191,N_2916);
or U6065 (N_6065,N_3315,N_3489);
and U6066 (N_6066,N_1702,N_3545);
and U6067 (N_6067,N_415,N_1101);
or U6068 (N_6068,N_0,N_1779);
nand U6069 (N_6069,N_2406,N_1135);
nor U6070 (N_6070,N_1960,N_2);
nor U6071 (N_6071,N_2591,N_3280);
nor U6072 (N_6072,N_2190,N_2806);
or U6073 (N_6073,N_3853,N_3818);
or U6074 (N_6074,N_2828,N_3934);
and U6075 (N_6075,N_2212,N_1645);
or U6076 (N_6076,N_3275,N_446);
nand U6077 (N_6077,N_457,N_156);
nor U6078 (N_6078,N_3606,N_2588);
and U6079 (N_6079,N_2899,N_982);
or U6080 (N_6080,N_3485,N_7);
nand U6081 (N_6081,N_1855,N_699);
and U6082 (N_6082,N_924,N_3246);
xnor U6083 (N_6083,N_108,N_2660);
xor U6084 (N_6084,N_659,N_2399);
or U6085 (N_6085,N_2299,N_3231);
nor U6086 (N_6086,N_979,N_2983);
and U6087 (N_6087,N_856,N_227);
and U6088 (N_6088,N_681,N_2268);
nand U6089 (N_6089,N_1868,N_555);
nor U6090 (N_6090,N_1578,N_1941);
nand U6091 (N_6091,N_2111,N_3767);
or U6092 (N_6092,N_2987,N_2450);
and U6093 (N_6093,N_924,N_3656);
xor U6094 (N_6094,N_518,N_981);
or U6095 (N_6095,N_2715,N_1088);
or U6096 (N_6096,N_3814,N_1380);
nand U6097 (N_6097,N_1191,N_1875);
or U6098 (N_6098,N_248,N_664);
xnor U6099 (N_6099,N_1544,N_3265);
nor U6100 (N_6100,N_1699,N_940);
or U6101 (N_6101,N_1706,N_847);
nand U6102 (N_6102,N_1588,N_2410);
nand U6103 (N_6103,N_1054,N_1166);
and U6104 (N_6104,N_518,N_1765);
nor U6105 (N_6105,N_3478,N_3766);
or U6106 (N_6106,N_3504,N_3243);
or U6107 (N_6107,N_3244,N_986);
and U6108 (N_6108,N_3797,N_2809);
nand U6109 (N_6109,N_3092,N_2498);
xnor U6110 (N_6110,N_1863,N_3529);
or U6111 (N_6111,N_2428,N_2140);
and U6112 (N_6112,N_802,N_1667);
nor U6113 (N_6113,N_1832,N_3464);
or U6114 (N_6114,N_479,N_353);
and U6115 (N_6115,N_1960,N_3441);
and U6116 (N_6116,N_154,N_1847);
or U6117 (N_6117,N_2811,N_1252);
nand U6118 (N_6118,N_2765,N_955);
nor U6119 (N_6119,N_626,N_691);
nor U6120 (N_6120,N_191,N_974);
nand U6121 (N_6121,N_636,N_2152);
nand U6122 (N_6122,N_93,N_1286);
or U6123 (N_6123,N_2974,N_2028);
nand U6124 (N_6124,N_990,N_521);
and U6125 (N_6125,N_2552,N_2013);
nor U6126 (N_6126,N_2733,N_3945);
or U6127 (N_6127,N_1683,N_2997);
nand U6128 (N_6128,N_1264,N_3880);
nand U6129 (N_6129,N_2985,N_1238);
and U6130 (N_6130,N_258,N_2472);
or U6131 (N_6131,N_565,N_1265);
and U6132 (N_6132,N_707,N_3757);
xnor U6133 (N_6133,N_952,N_1090);
xor U6134 (N_6134,N_1738,N_3184);
or U6135 (N_6135,N_1794,N_2807);
and U6136 (N_6136,N_2557,N_3647);
xor U6137 (N_6137,N_3702,N_1012);
and U6138 (N_6138,N_3588,N_3397);
xor U6139 (N_6139,N_244,N_1205);
nor U6140 (N_6140,N_591,N_3837);
or U6141 (N_6141,N_3281,N_1076);
nand U6142 (N_6142,N_1237,N_1482);
nor U6143 (N_6143,N_1927,N_2798);
or U6144 (N_6144,N_1312,N_1712);
or U6145 (N_6145,N_2913,N_3165);
and U6146 (N_6146,N_2334,N_1556);
nand U6147 (N_6147,N_3141,N_1238);
nand U6148 (N_6148,N_821,N_301);
nand U6149 (N_6149,N_3939,N_2221);
and U6150 (N_6150,N_2144,N_155);
and U6151 (N_6151,N_3835,N_3095);
nand U6152 (N_6152,N_3155,N_1447);
nor U6153 (N_6153,N_2438,N_2940);
nor U6154 (N_6154,N_3204,N_2772);
xnor U6155 (N_6155,N_473,N_678);
nand U6156 (N_6156,N_2518,N_1351);
nand U6157 (N_6157,N_425,N_953);
nor U6158 (N_6158,N_2718,N_2100);
or U6159 (N_6159,N_2031,N_900);
nand U6160 (N_6160,N_3120,N_2107);
and U6161 (N_6161,N_2931,N_3108);
and U6162 (N_6162,N_53,N_2915);
nor U6163 (N_6163,N_344,N_3810);
nand U6164 (N_6164,N_2978,N_3031);
nor U6165 (N_6165,N_1581,N_791);
nand U6166 (N_6166,N_2204,N_736);
nor U6167 (N_6167,N_3485,N_1258);
nand U6168 (N_6168,N_2257,N_454);
and U6169 (N_6169,N_2119,N_813);
or U6170 (N_6170,N_3183,N_2738);
or U6171 (N_6171,N_1185,N_2674);
and U6172 (N_6172,N_1379,N_3618);
and U6173 (N_6173,N_1176,N_2461);
nor U6174 (N_6174,N_162,N_2203);
xor U6175 (N_6175,N_1859,N_2980);
or U6176 (N_6176,N_2546,N_3072);
nor U6177 (N_6177,N_2996,N_2355);
and U6178 (N_6178,N_3450,N_3727);
nor U6179 (N_6179,N_3466,N_3674);
nor U6180 (N_6180,N_3933,N_827);
nor U6181 (N_6181,N_3850,N_2753);
and U6182 (N_6182,N_1172,N_1767);
nand U6183 (N_6183,N_1993,N_770);
or U6184 (N_6184,N_1190,N_3160);
and U6185 (N_6185,N_2199,N_815);
or U6186 (N_6186,N_2838,N_12);
nand U6187 (N_6187,N_2601,N_805);
xnor U6188 (N_6188,N_569,N_1172);
or U6189 (N_6189,N_2849,N_1750);
nor U6190 (N_6190,N_379,N_601);
or U6191 (N_6191,N_54,N_386);
nor U6192 (N_6192,N_3507,N_644);
nor U6193 (N_6193,N_2906,N_1188);
nand U6194 (N_6194,N_1522,N_1822);
nor U6195 (N_6195,N_744,N_2244);
nor U6196 (N_6196,N_1283,N_2277);
or U6197 (N_6197,N_298,N_2055);
nand U6198 (N_6198,N_3096,N_1605);
and U6199 (N_6199,N_336,N_560);
nor U6200 (N_6200,N_804,N_476);
nand U6201 (N_6201,N_3726,N_3472);
xnor U6202 (N_6202,N_835,N_2212);
and U6203 (N_6203,N_1703,N_3659);
and U6204 (N_6204,N_2749,N_2909);
nand U6205 (N_6205,N_212,N_127);
and U6206 (N_6206,N_798,N_2642);
or U6207 (N_6207,N_2728,N_1976);
or U6208 (N_6208,N_1165,N_289);
or U6209 (N_6209,N_2576,N_3610);
xnor U6210 (N_6210,N_637,N_2992);
nand U6211 (N_6211,N_448,N_3096);
or U6212 (N_6212,N_2000,N_953);
nand U6213 (N_6213,N_2964,N_120);
and U6214 (N_6214,N_2121,N_138);
or U6215 (N_6215,N_2560,N_1907);
nor U6216 (N_6216,N_305,N_932);
and U6217 (N_6217,N_2083,N_400);
nand U6218 (N_6218,N_3739,N_2934);
nand U6219 (N_6219,N_2298,N_3646);
xnor U6220 (N_6220,N_2283,N_3982);
or U6221 (N_6221,N_893,N_943);
nor U6222 (N_6222,N_1776,N_102);
or U6223 (N_6223,N_1296,N_2091);
nand U6224 (N_6224,N_1055,N_336);
or U6225 (N_6225,N_2753,N_2260);
nand U6226 (N_6226,N_3299,N_1380);
or U6227 (N_6227,N_3694,N_1216);
xor U6228 (N_6228,N_1827,N_3089);
nand U6229 (N_6229,N_1558,N_12);
or U6230 (N_6230,N_2962,N_842);
nand U6231 (N_6231,N_2368,N_2784);
nor U6232 (N_6232,N_772,N_3186);
nor U6233 (N_6233,N_75,N_749);
nor U6234 (N_6234,N_2629,N_243);
nor U6235 (N_6235,N_3404,N_1594);
nor U6236 (N_6236,N_337,N_1508);
and U6237 (N_6237,N_2034,N_3822);
and U6238 (N_6238,N_2583,N_2484);
nor U6239 (N_6239,N_1552,N_2231);
nor U6240 (N_6240,N_1893,N_1062);
and U6241 (N_6241,N_70,N_3467);
nand U6242 (N_6242,N_2676,N_975);
nor U6243 (N_6243,N_2745,N_604);
or U6244 (N_6244,N_2391,N_2122);
nor U6245 (N_6245,N_2603,N_2171);
nor U6246 (N_6246,N_3212,N_3930);
nor U6247 (N_6247,N_3480,N_990);
nor U6248 (N_6248,N_1490,N_3881);
nor U6249 (N_6249,N_3795,N_3581);
or U6250 (N_6250,N_3296,N_1985);
or U6251 (N_6251,N_1380,N_1863);
or U6252 (N_6252,N_2186,N_785);
or U6253 (N_6253,N_2458,N_2769);
and U6254 (N_6254,N_2030,N_2814);
or U6255 (N_6255,N_1170,N_2213);
and U6256 (N_6256,N_1224,N_1248);
xnor U6257 (N_6257,N_519,N_847);
nand U6258 (N_6258,N_1387,N_1775);
and U6259 (N_6259,N_2019,N_2757);
nand U6260 (N_6260,N_58,N_1494);
and U6261 (N_6261,N_3211,N_1290);
xnor U6262 (N_6262,N_318,N_2216);
nand U6263 (N_6263,N_1729,N_2286);
nor U6264 (N_6264,N_2305,N_2929);
xor U6265 (N_6265,N_1299,N_3570);
or U6266 (N_6266,N_1718,N_2150);
nand U6267 (N_6267,N_2803,N_2779);
and U6268 (N_6268,N_739,N_1148);
or U6269 (N_6269,N_138,N_527);
or U6270 (N_6270,N_3611,N_627);
nand U6271 (N_6271,N_646,N_1272);
xnor U6272 (N_6272,N_1598,N_2352);
nor U6273 (N_6273,N_930,N_1546);
nor U6274 (N_6274,N_2390,N_1877);
nor U6275 (N_6275,N_1201,N_3520);
and U6276 (N_6276,N_498,N_2239);
nor U6277 (N_6277,N_1589,N_2856);
nand U6278 (N_6278,N_2578,N_729);
or U6279 (N_6279,N_2666,N_1520);
nor U6280 (N_6280,N_2750,N_197);
xor U6281 (N_6281,N_3515,N_854);
xnor U6282 (N_6282,N_1519,N_3596);
xor U6283 (N_6283,N_3932,N_3017);
or U6284 (N_6284,N_1962,N_1724);
nand U6285 (N_6285,N_784,N_84);
xnor U6286 (N_6286,N_1300,N_3355);
nand U6287 (N_6287,N_2818,N_3279);
or U6288 (N_6288,N_1400,N_1920);
and U6289 (N_6289,N_2488,N_218);
and U6290 (N_6290,N_394,N_1827);
nand U6291 (N_6291,N_2711,N_1373);
or U6292 (N_6292,N_1931,N_1673);
nand U6293 (N_6293,N_3509,N_3399);
or U6294 (N_6294,N_569,N_85);
nand U6295 (N_6295,N_742,N_3463);
nand U6296 (N_6296,N_1184,N_2861);
nand U6297 (N_6297,N_2232,N_1537);
xnor U6298 (N_6298,N_3572,N_920);
xnor U6299 (N_6299,N_835,N_1042);
and U6300 (N_6300,N_210,N_2488);
and U6301 (N_6301,N_3806,N_2826);
nand U6302 (N_6302,N_2096,N_487);
nand U6303 (N_6303,N_2340,N_1371);
and U6304 (N_6304,N_820,N_407);
xor U6305 (N_6305,N_2622,N_48);
or U6306 (N_6306,N_3421,N_1591);
and U6307 (N_6307,N_2093,N_2970);
or U6308 (N_6308,N_3376,N_387);
xnor U6309 (N_6309,N_1201,N_2495);
nand U6310 (N_6310,N_3172,N_2835);
or U6311 (N_6311,N_998,N_2658);
and U6312 (N_6312,N_831,N_3675);
xor U6313 (N_6313,N_1871,N_1277);
or U6314 (N_6314,N_3846,N_2691);
and U6315 (N_6315,N_392,N_1914);
and U6316 (N_6316,N_2039,N_1629);
nor U6317 (N_6317,N_3175,N_1058);
xnor U6318 (N_6318,N_2422,N_2650);
nand U6319 (N_6319,N_52,N_664);
nand U6320 (N_6320,N_1770,N_3814);
nand U6321 (N_6321,N_585,N_3917);
nand U6322 (N_6322,N_2704,N_96);
or U6323 (N_6323,N_378,N_262);
or U6324 (N_6324,N_3241,N_3728);
and U6325 (N_6325,N_852,N_600);
nor U6326 (N_6326,N_1250,N_5);
nand U6327 (N_6327,N_3390,N_1093);
and U6328 (N_6328,N_2454,N_2053);
and U6329 (N_6329,N_1198,N_2464);
and U6330 (N_6330,N_2592,N_2828);
nand U6331 (N_6331,N_1784,N_802);
and U6332 (N_6332,N_1383,N_603);
nand U6333 (N_6333,N_3029,N_1659);
or U6334 (N_6334,N_488,N_3114);
nor U6335 (N_6335,N_2065,N_3224);
or U6336 (N_6336,N_1825,N_3289);
nor U6337 (N_6337,N_3022,N_159);
and U6338 (N_6338,N_2571,N_352);
or U6339 (N_6339,N_214,N_3445);
or U6340 (N_6340,N_2826,N_2633);
nand U6341 (N_6341,N_1529,N_1438);
nand U6342 (N_6342,N_780,N_2102);
xor U6343 (N_6343,N_2595,N_3024);
and U6344 (N_6344,N_2234,N_3189);
and U6345 (N_6345,N_2988,N_92);
nor U6346 (N_6346,N_417,N_1831);
nor U6347 (N_6347,N_1861,N_3297);
nor U6348 (N_6348,N_1115,N_419);
nor U6349 (N_6349,N_79,N_2281);
nand U6350 (N_6350,N_1452,N_2451);
or U6351 (N_6351,N_3125,N_410);
nor U6352 (N_6352,N_3372,N_2095);
and U6353 (N_6353,N_256,N_2981);
and U6354 (N_6354,N_2967,N_3282);
nor U6355 (N_6355,N_3775,N_3147);
nor U6356 (N_6356,N_392,N_3228);
or U6357 (N_6357,N_825,N_1670);
nand U6358 (N_6358,N_1620,N_926);
or U6359 (N_6359,N_1516,N_2278);
and U6360 (N_6360,N_619,N_3557);
nand U6361 (N_6361,N_1015,N_1176);
xor U6362 (N_6362,N_2754,N_2787);
nand U6363 (N_6363,N_2609,N_3555);
or U6364 (N_6364,N_1959,N_3687);
xnor U6365 (N_6365,N_1873,N_505);
nor U6366 (N_6366,N_2844,N_1883);
nor U6367 (N_6367,N_392,N_3591);
nor U6368 (N_6368,N_2199,N_980);
or U6369 (N_6369,N_287,N_89);
nor U6370 (N_6370,N_3955,N_1493);
nand U6371 (N_6371,N_1851,N_1964);
or U6372 (N_6372,N_1414,N_919);
nor U6373 (N_6373,N_3447,N_3657);
nand U6374 (N_6374,N_1590,N_2006);
xnor U6375 (N_6375,N_988,N_1257);
nand U6376 (N_6376,N_2408,N_2178);
nor U6377 (N_6377,N_1063,N_2972);
or U6378 (N_6378,N_163,N_1801);
and U6379 (N_6379,N_3830,N_3014);
nand U6380 (N_6380,N_3581,N_3071);
and U6381 (N_6381,N_3305,N_1731);
or U6382 (N_6382,N_3085,N_1867);
nor U6383 (N_6383,N_576,N_538);
nor U6384 (N_6384,N_3440,N_1665);
or U6385 (N_6385,N_1291,N_3055);
or U6386 (N_6386,N_189,N_1202);
or U6387 (N_6387,N_2096,N_3917);
nand U6388 (N_6388,N_2957,N_3963);
or U6389 (N_6389,N_1477,N_190);
nor U6390 (N_6390,N_491,N_758);
nand U6391 (N_6391,N_2807,N_3013);
nand U6392 (N_6392,N_2098,N_1445);
nor U6393 (N_6393,N_1324,N_1019);
and U6394 (N_6394,N_1678,N_2005);
nor U6395 (N_6395,N_1889,N_3540);
nor U6396 (N_6396,N_801,N_634);
nand U6397 (N_6397,N_1719,N_664);
xor U6398 (N_6398,N_3520,N_714);
nand U6399 (N_6399,N_2102,N_3897);
and U6400 (N_6400,N_615,N_975);
and U6401 (N_6401,N_3319,N_2602);
xnor U6402 (N_6402,N_1384,N_1217);
nor U6403 (N_6403,N_1225,N_3045);
nor U6404 (N_6404,N_255,N_126);
or U6405 (N_6405,N_2887,N_291);
and U6406 (N_6406,N_3001,N_1805);
xor U6407 (N_6407,N_2447,N_913);
xnor U6408 (N_6408,N_1763,N_3878);
nand U6409 (N_6409,N_533,N_3824);
or U6410 (N_6410,N_3209,N_11);
xor U6411 (N_6411,N_3878,N_1163);
or U6412 (N_6412,N_1891,N_913);
and U6413 (N_6413,N_1394,N_1046);
or U6414 (N_6414,N_246,N_2734);
and U6415 (N_6415,N_689,N_251);
or U6416 (N_6416,N_2562,N_1548);
xnor U6417 (N_6417,N_2774,N_1978);
and U6418 (N_6418,N_3888,N_3974);
or U6419 (N_6419,N_2055,N_1059);
nor U6420 (N_6420,N_2893,N_2993);
nand U6421 (N_6421,N_1405,N_3496);
or U6422 (N_6422,N_2045,N_2482);
nand U6423 (N_6423,N_3039,N_1945);
and U6424 (N_6424,N_3909,N_138);
xnor U6425 (N_6425,N_3717,N_2558);
and U6426 (N_6426,N_936,N_2908);
and U6427 (N_6427,N_1264,N_2165);
and U6428 (N_6428,N_342,N_2911);
or U6429 (N_6429,N_2306,N_1938);
nand U6430 (N_6430,N_1898,N_577);
or U6431 (N_6431,N_3145,N_202);
nor U6432 (N_6432,N_525,N_181);
and U6433 (N_6433,N_321,N_1480);
or U6434 (N_6434,N_1385,N_571);
nor U6435 (N_6435,N_1196,N_2715);
nand U6436 (N_6436,N_588,N_56);
and U6437 (N_6437,N_1568,N_54);
and U6438 (N_6438,N_2671,N_574);
nor U6439 (N_6439,N_2935,N_1438);
nand U6440 (N_6440,N_2184,N_537);
nor U6441 (N_6441,N_3895,N_192);
nor U6442 (N_6442,N_3227,N_3073);
nand U6443 (N_6443,N_1984,N_618);
and U6444 (N_6444,N_1534,N_660);
and U6445 (N_6445,N_2155,N_1612);
xor U6446 (N_6446,N_1693,N_1689);
or U6447 (N_6447,N_3644,N_713);
or U6448 (N_6448,N_3936,N_348);
nand U6449 (N_6449,N_3265,N_1834);
nand U6450 (N_6450,N_3634,N_1598);
nor U6451 (N_6451,N_419,N_1423);
nor U6452 (N_6452,N_105,N_1946);
nor U6453 (N_6453,N_3465,N_747);
nand U6454 (N_6454,N_380,N_1660);
and U6455 (N_6455,N_716,N_2137);
or U6456 (N_6456,N_1235,N_1504);
xor U6457 (N_6457,N_739,N_1618);
and U6458 (N_6458,N_1785,N_28);
or U6459 (N_6459,N_3730,N_2095);
or U6460 (N_6460,N_1532,N_364);
or U6461 (N_6461,N_906,N_1006);
nor U6462 (N_6462,N_1841,N_2642);
nor U6463 (N_6463,N_217,N_3348);
nand U6464 (N_6464,N_2166,N_2746);
xnor U6465 (N_6465,N_3235,N_1278);
xnor U6466 (N_6466,N_15,N_1954);
and U6467 (N_6467,N_189,N_23);
xnor U6468 (N_6468,N_608,N_1407);
nand U6469 (N_6469,N_3715,N_2926);
nand U6470 (N_6470,N_2676,N_2224);
or U6471 (N_6471,N_2891,N_3120);
and U6472 (N_6472,N_3872,N_3654);
nand U6473 (N_6473,N_3079,N_1342);
and U6474 (N_6474,N_3469,N_546);
nand U6475 (N_6475,N_2260,N_2339);
nand U6476 (N_6476,N_584,N_2414);
nor U6477 (N_6477,N_1398,N_3414);
xor U6478 (N_6478,N_1191,N_3059);
nand U6479 (N_6479,N_2100,N_2669);
and U6480 (N_6480,N_1687,N_2949);
and U6481 (N_6481,N_1522,N_1040);
and U6482 (N_6482,N_737,N_1307);
nand U6483 (N_6483,N_3764,N_1703);
or U6484 (N_6484,N_3959,N_3064);
nand U6485 (N_6485,N_2147,N_2967);
nor U6486 (N_6486,N_1848,N_425);
and U6487 (N_6487,N_1448,N_3203);
or U6488 (N_6488,N_1619,N_626);
and U6489 (N_6489,N_498,N_1227);
nand U6490 (N_6490,N_2260,N_1144);
nor U6491 (N_6491,N_1925,N_1560);
and U6492 (N_6492,N_3164,N_3671);
nand U6493 (N_6493,N_455,N_519);
or U6494 (N_6494,N_1131,N_490);
xnor U6495 (N_6495,N_1743,N_691);
or U6496 (N_6496,N_2032,N_2992);
or U6497 (N_6497,N_1527,N_652);
and U6498 (N_6498,N_2743,N_3516);
or U6499 (N_6499,N_1158,N_3612);
nand U6500 (N_6500,N_734,N_1587);
or U6501 (N_6501,N_2408,N_2337);
xnor U6502 (N_6502,N_646,N_3728);
or U6503 (N_6503,N_3669,N_2257);
nor U6504 (N_6504,N_201,N_3018);
or U6505 (N_6505,N_1876,N_2352);
nand U6506 (N_6506,N_509,N_3587);
and U6507 (N_6507,N_3116,N_956);
xor U6508 (N_6508,N_1087,N_2654);
and U6509 (N_6509,N_2274,N_3411);
nor U6510 (N_6510,N_1182,N_755);
nor U6511 (N_6511,N_1754,N_3549);
or U6512 (N_6512,N_1380,N_2901);
nor U6513 (N_6513,N_3901,N_662);
nor U6514 (N_6514,N_804,N_1086);
nand U6515 (N_6515,N_1720,N_286);
nand U6516 (N_6516,N_2665,N_2139);
and U6517 (N_6517,N_3219,N_2474);
nand U6518 (N_6518,N_2891,N_3549);
nand U6519 (N_6519,N_1743,N_2224);
or U6520 (N_6520,N_2869,N_1206);
nand U6521 (N_6521,N_1207,N_2730);
nand U6522 (N_6522,N_695,N_2646);
nand U6523 (N_6523,N_1476,N_116);
and U6524 (N_6524,N_2853,N_2127);
and U6525 (N_6525,N_470,N_756);
nor U6526 (N_6526,N_8,N_3868);
nand U6527 (N_6527,N_1013,N_3963);
nor U6528 (N_6528,N_2808,N_952);
nor U6529 (N_6529,N_3978,N_2464);
nand U6530 (N_6530,N_2068,N_1344);
nand U6531 (N_6531,N_3506,N_1508);
nor U6532 (N_6532,N_3401,N_1896);
nor U6533 (N_6533,N_2939,N_3551);
and U6534 (N_6534,N_554,N_3181);
nor U6535 (N_6535,N_606,N_2752);
and U6536 (N_6536,N_1694,N_61);
nand U6537 (N_6537,N_2308,N_878);
nor U6538 (N_6538,N_1840,N_1557);
or U6539 (N_6539,N_1370,N_3522);
or U6540 (N_6540,N_1079,N_2971);
nor U6541 (N_6541,N_3793,N_1063);
or U6542 (N_6542,N_3839,N_3941);
nor U6543 (N_6543,N_3058,N_3191);
nand U6544 (N_6544,N_154,N_1828);
nor U6545 (N_6545,N_474,N_2005);
or U6546 (N_6546,N_2763,N_823);
and U6547 (N_6547,N_1855,N_3468);
nand U6548 (N_6548,N_2720,N_1698);
xor U6549 (N_6549,N_2114,N_512);
nor U6550 (N_6550,N_825,N_573);
nand U6551 (N_6551,N_503,N_784);
and U6552 (N_6552,N_3301,N_1980);
and U6553 (N_6553,N_724,N_3352);
and U6554 (N_6554,N_387,N_2479);
and U6555 (N_6555,N_3745,N_2553);
or U6556 (N_6556,N_1398,N_1731);
nand U6557 (N_6557,N_2833,N_2945);
or U6558 (N_6558,N_1316,N_1430);
and U6559 (N_6559,N_1894,N_934);
nor U6560 (N_6560,N_3543,N_1035);
or U6561 (N_6561,N_1084,N_2336);
nand U6562 (N_6562,N_3654,N_484);
nor U6563 (N_6563,N_3872,N_531);
nor U6564 (N_6564,N_637,N_1243);
and U6565 (N_6565,N_3083,N_914);
xor U6566 (N_6566,N_2308,N_3246);
nand U6567 (N_6567,N_1621,N_2206);
nand U6568 (N_6568,N_2587,N_304);
or U6569 (N_6569,N_3908,N_1842);
xnor U6570 (N_6570,N_740,N_2752);
nand U6571 (N_6571,N_2723,N_3234);
nand U6572 (N_6572,N_823,N_2573);
or U6573 (N_6573,N_3248,N_3982);
nor U6574 (N_6574,N_2379,N_1494);
nand U6575 (N_6575,N_1572,N_2305);
or U6576 (N_6576,N_540,N_1580);
xnor U6577 (N_6577,N_2548,N_716);
xor U6578 (N_6578,N_1059,N_2336);
nor U6579 (N_6579,N_963,N_3129);
nand U6580 (N_6580,N_3995,N_3410);
nand U6581 (N_6581,N_2736,N_911);
and U6582 (N_6582,N_2435,N_3241);
and U6583 (N_6583,N_1248,N_1929);
and U6584 (N_6584,N_3152,N_2102);
nor U6585 (N_6585,N_1649,N_2757);
and U6586 (N_6586,N_3098,N_1436);
and U6587 (N_6587,N_455,N_664);
nor U6588 (N_6588,N_2229,N_676);
or U6589 (N_6589,N_1310,N_2924);
nand U6590 (N_6590,N_1392,N_1052);
nor U6591 (N_6591,N_2737,N_586);
nand U6592 (N_6592,N_3700,N_3500);
and U6593 (N_6593,N_1524,N_1061);
and U6594 (N_6594,N_2321,N_123);
and U6595 (N_6595,N_142,N_1097);
or U6596 (N_6596,N_527,N_2643);
xnor U6597 (N_6597,N_2310,N_1295);
and U6598 (N_6598,N_2608,N_2326);
and U6599 (N_6599,N_3998,N_21);
nand U6600 (N_6600,N_1622,N_1430);
nor U6601 (N_6601,N_3875,N_2065);
and U6602 (N_6602,N_1845,N_3141);
nor U6603 (N_6603,N_428,N_168);
nor U6604 (N_6604,N_647,N_1885);
or U6605 (N_6605,N_1146,N_309);
and U6606 (N_6606,N_1306,N_1495);
xnor U6607 (N_6607,N_2988,N_3843);
or U6608 (N_6608,N_3998,N_287);
or U6609 (N_6609,N_206,N_28);
nor U6610 (N_6610,N_1501,N_1366);
or U6611 (N_6611,N_3884,N_2952);
or U6612 (N_6612,N_517,N_80);
and U6613 (N_6613,N_1992,N_2836);
and U6614 (N_6614,N_2530,N_447);
and U6615 (N_6615,N_2660,N_1620);
and U6616 (N_6616,N_338,N_236);
nor U6617 (N_6617,N_3676,N_2381);
or U6618 (N_6618,N_2671,N_1186);
nor U6619 (N_6619,N_2358,N_2589);
or U6620 (N_6620,N_1780,N_104);
or U6621 (N_6621,N_3993,N_2408);
or U6622 (N_6622,N_3006,N_3532);
xnor U6623 (N_6623,N_370,N_2142);
nor U6624 (N_6624,N_859,N_2299);
nor U6625 (N_6625,N_3944,N_2589);
and U6626 (N_6626,N_2817,N_3834);
and U6627 (N_6627,N_2616,N_3373);
nand U6628 (N_6628,N_1093,N_529);
and U6629 (N_6629,N_335,N_462);
nand U6630 (N_6630,N_1852,N_1798);
or U6631 (N_6631,N_2476,N_417);
or U6632 (N_6632,N_566,N_1594);
nand U6633 (N_6633,N_3146,N_647);
nand U6634 (N_6634,N_1925,N_1272);
nor U6635 (N_6635,N_2022,N_993);
nor U6636 (N_6636,N_1607,N_2012);
xor U6637 (N_6637,N_3214,N_2740);
nor U6638 (N_6638,N_2613,N_249);
nand U6639 (N_6639,N_630,N_627);
and U6640 (N_6640,N_3197,N_3604);
or U6641 (N_6641,N_1809,N_1397);
or U6642 (N_6642,N_2487,N_3323);
nand U6643 (N_6643,N_2685,N_1950);
or U6644 (N_6644,N_139,N_3869);
and U6645 (N_6645,N_3560,N_2574);
nand U6646 (N_6646,N_2032,N_1307);
nand U6647 (N_6647,N_2819,N_873);
nand U6648 (N_6648,N_1433,N_1638);
and U6649 (N_6649,N_1811,N_1179);
nand U6650 (N_6650,N_1394,N_712);
and U6651 (N_6651,N_3720,N_3313);
nand U6652 (N_6652,N_2613,N_1882);
xnor U6653 (N_6653,N_2662,N_2981);
nand U6654 (N_6654,N_1304,N_1174);
nand U6655 (N_6655,N_1938,N_164);
nor U6656 (N_6656,N_1515,N_3165);
and U6657 (N_6657,N_1544,N_1215);
or U6658 (N_6658,N_3713,N_311);
and U6659 (N_6659,N_778,N_2469);
and U6660 (N_6660,N_2478,N_1060);
xnor U6661 (N_6661,N_3130,N_2185);
and U6662 (N_6662,N_1805,N_604);
or U6663 (N_6663,N_2743,N_3077);
nand U6664 (N_6664,N_1903,N_3941);
or U6665 (N_6665,N_2185,N_1695);
nor U6666 (N_6666,N_1969,N_2054);
nor U6667 (N_6667,N_2197,N_447);
nand U6668 (N_6668,N_1427,N_2988);
nand U6669 (N_6669,N_2372,N_3402);
or U6670 (N_6670,N_3164,N_1824);
nand U6671 (N_6671,N_1389,N_3283);
or U6672 (N_6672,N_939,N_2127);
nand U6673 (N_6673,N_2986,N_3343);
xor U6674 (N_6674,N_664,N_976);
nand U6675 (N_6675,N_2883,N_1654);
nor U6676 (N_6676,N_3241,N_2252);
xnor U6677 (N_6677,N_577,N_1608);
or U6678 (N_6678,N_1903,N_321);
or U6679 (N_6679,N_411,N_91);
and U6680 (N_6680,N_2430,N_3076);
or U6681 (N_6681,N_828,N_3004);
nor U6682 (N_6682,N_492,N_124);
and U6683 (N_6683,N_3767,N_2744);
or U6684 (N_6684,N_610,N_1097);
nand U6685 (N_6685,N_1227,N_3564);
and U6686 (N_6686,N_3300,N_3386);
or U6687 (N_6687,N_3557,N_3740);
or U6688 (N_6688,N_2001,N_3423);
xnor U6689 (N_6689,N_1966,N_474);
nand U6690 (N_6690,N_2571,N_1839);
nand U6691 (N_6691,N_2787,N_1531);
nand U6692 (N_6692,N_1049,N_2797);
or U6693 (N_6693,N_1650,N_2760);
or U6694 (N_6694,N_2028,N_3571);
xnor U6695 (N_6695,N_2369,N_3898);
or U6696 (N_6696,N_3526,N_380);
or U6697 (N_6697,N_2493,N_2937);
xnor U6698 (N_6698,N_1420,N_1747);
nor U6699 (N_6699,N_1980,N_2175);
nand U6700 (N_6700,N_2691,N_3736);
and U6701 (N_6701,N_1366,N_2787);
xnor U6702 (N_6702,N_1045,N_2360);
xnor U6703 (N_6703,N_2457,N_1504);
xor U6704 (N_6704,N_745,N_537);
nand U6705 (N_6705,N_1077,N_2071);
nand U6706 (N_6706,N_3527,N_2964);
and U6707 (N_6707,N_302,N_1196);
or U6708 (N_6708,N_792,N_779);
and U6709 (N_6709,N_748,N_384);
or U6710 (N_6710,N_1020,N_2941);
nor U6711 (N_6711,N_1487,N_793);
xor U6712 (N_6712,N_3426,N_3757);
nand U6713 (N_6713,N_2879,N_536);
nor U6714 (N_6714,N_554,N_2816);
or U6715 (N_6715,N_2378,N_3761);
or U6716 (N_6716,N_1962,N_2669);
or U6717 (N_6717,N_1397,N_2231);
nand U6718 (N_6718,N_328,N_3891);
nand U6719 (N_6719,N_2375,N_2278);
or U6720 (N_6720,N_3767,N_2092);
xor U6721 (N_6721,N_502,N_2309);
or U6722 (N_6722,N_3599,N_575);
or U6723 (N_6723,N_111,N_1456);
and U6724 (N_6724,N_368,N_3563);
nor U6725 (N_6725,N_3214,N_108);
and U6726 (N_6726,N_24,N_2855);
or U6727 (N_6727,N_1494,N_3119);
nand U6728 (N_6728,N_842,N_3045);
or U6729 (N_6729,N_3956,N_609);
and U6730 (N_6730,N_3092,N_3528);
xnor U6731 (N_6731,N_3298,N_1127);
nand U6732 (N_6732,N_2794,N_874);
nand U6733 (N_6733,N_1740,N_3046);
or U6734 (N_6734,N_1793,N_2605);
nand U6735 (N_6735,N_2256,N_2067);
nand U6736 (N_6736,N_2258,N_1533);
nor U6737 (N_6737,N_2052,N_1302);
or U6738 (N_6738,N_1566,N_1220);
nand U6739 (N_6739,N_3631,N_840);
and U6740 (N_6740,N_1240,N_2586);
nand U6741 (N_6741,N_469,N_1262);
nor U6742 (N_6742,N_496,N_1188);
xnor U6743 (N_6743,N_2388,N_1362);
or U6744 (N_6744,N_3955,N_1792);
or U6745 (N_6745,N_3212,N_2341);
and U6746 (N_6746,N_568,N_682);
nor U6747 (N_6747,N_3987,N_64);
xnor U6748 (N_6748,N_534,N_2691);
or U6749 (N_6749,N_3052,N_3688);
nor U6750 (N_6750,N_1067,N_11);
or U6751 (N_6751,N_116,N_2226);
xor U6752 (N_6752,N_2664,N_3265);
or U6753 (N_6753,N_1692,N_3451);
or U6754 (N_6754,N_803,N_3462);
xnor U6755 (N_6755,N_242,N_704);
nand U6756 (N_6756,N_2248,N_1079);
and U6757 (N_6757,N_2765,N_943);
or U6758 (N_6758,N_1544,N_3535);
nor U6759 (N_6759,N_2779,N_3163);
and U6760 (N_6760,N_2367,N_3183);
xnor U6761 (N_6761,N_1767,N_1209);
and U6762 (N_6762,N_3075,N_974);
nand U6763 (N_6763,N_3671,N_3540);
nand U6764 (N_6764,N_3916,N_3365);
and U6765 (N_6765,N_287,N_2772);
and U6766 (N_6766,N_13,N_2365);
or U6767 (N_6767,N_1297,N_2713);
xnor U6768 (N_6768,N_3497,N_2918);
or U6769 (N_6769,N_3923,N_3446);
nand U6770 (N_6770,N_3357,N_2604);
and U6771 (N_6771,N_209,N_3832);
and U6772 (N_6772,N_3731,N_3056);
xnor U6773 (N_6773,N_1015,N_3747);
xor U6774 (N_6774,N_329,N_2977);
or U6775 (N_6775,N_3707,N_43);
or U6776 (N_6776,N_157,N_2589);
and U6777 (N_6777,N_1817,N_855);
nor U6778 (N_6778,N_1336,N_2972);
xnor U6779 (N_6779,N_3441,N_3538);
or U6780 (N_6780,N_2796,N_2214);
nand U6781 (N_6781,N_1238,N_257);
xor U6782 (N_6782,N_2632,N_3460);
xor U6783 (N_6783,N_2307,N_1151);
nor U6784 (N_6784,N_2405,N_2932);
and U6785 (N_6785,N_300,N_1886);
or U6786 (N_6786,N_2446,N_806);
nand U6787 (N_6787,N_3089,N_3880);
nor U6788 (N_6788,N_1443,N_2519);
or U6789 (N_6789,N_2604,N_824);
nor U6790 (N_6790,N_2247,N_1275);
nor U6791 (N_6791,N_2417,N_3268);
and U6792 (N_6792,N_1231,N_2139);
xor U6793 (N_6793,N_3352,N_3660);
or U6794 (N_6794,N_1423,N_2717);
and U6795 (N_6795,N_1864,N_1099);
nand U6796 (N_6796,N_3875,N_176);
and U6797 (N_6797,N_1667,N_661);
nand U6798 (N_6798,N_3620,N_2561);
xnor U6799 (N_6799,N_1676,N_584);
and U6800 (N_6800,N_3753,N_3385);
nor U6801 (N_6801,N_1255,N_881);
nor U6802 (N_6802,N_163,N_2704);
or U6803 (N_6803,N_1455,N_2483);
or U6804 (N_6804,N_2632,N_1648);
nand U6805 (N_6805,N_3683,N_3539);
xor U6806 (N_6806,N_3369,N_949);
and U6807 (N_6807,N_2654,N_3250);
nor U6808 (N_6808,N_3721,N_519);
xnor U6809 (N_6809,N_3096,N_2640);
nand U6810 (N_6810,N_985,N_47);
nand U6811 (N_6811,N_359,N_735);
nor U6812 (N_6812,N_701,N_533);
nor U6813 (N_6813,N_1410,N_2480);
nor U6814 (N_6814,N_3944,N_1315);
xor U6815 (N_6815,N_1283,N_2527);
or U6816 (N_6816,N_570,N_2427);
nand U6817 (N_6817,N_3640,N_2518);
nand U6818 (N_6818,N_1251,N_1601);
nor U6819 (N_6819,N_1334,N_1090);
and U6820 (N_6820,N_2579,N_3412);
and U6821 (N_6821,N_1408,N_540);
or U6822 (N_6822,N_412,N_3258);
or U6823 (N_6823,N_1513,N_2626);
nand U6824 (N_6824,N_350,N_880);
and U6825 (N_6825,N_3816,N_894);
or U6826 (N_6826,N_2304,N_398);
or U6827 (N_6827,N_1811,N_1227);
nor U6828 (N_6828,N_1319,N_1189);
nor U6829 (N_6829,N_2176,N_1707);
or U6830 (N_6830,N_1990,N_1654);
nand U6831 (N_6831,N_783,N_2934);
nor U6832 (N_6832,N_348,N_3226);
and U6833 (N_6833,N_1653,N_2296);
nor U6834 (N_6834,N_743,N_654);
and U6835 (N_6835,N_2660,N_24);
or U6836 (N_6836,N_3963,N_56);
xor U6837 (N_6837,N_1534,N_3260);
nand U6838 (N_6838,N_1495,N_1516);
and U6839 (N_6839,N_613,N_1185);
nor U6840 (N_6840,N_1108,N_2762);
nor U6841 (N_6841,N_2301,N_1256);
and U6842 (N_6842,N_803,N_257);
and U6843 (N_6843,N_3857,N_1667);
nor U6844 (N_6844,N_2287,N_517);
or U6845 (N_6845,N_497,N_3163);
nor U6846 (N_6846,N_448,N_2923);
nor U6847 (N_6847,N_519,N_1055);
and U6848 (N_6848,N_3332,N_111);
and U6849 (N_6849,N_1811,N_2164);
and U6850 (N_6850,N_2166,N_2203);
and U6851 (N_6851,N_140,N_3968);
nor U6852 (N_6852,N_1201,N_3262);
nor U6853 (N_6853,N_1322,N_411);
nor U6854 (N_6854,N_565,N_2338);
and U6855 (N_6855,N_3273,N_2023);
and U6856 (N_6856,N_3169,N_3610);
xnor U6857 (N_6857,N_965,N_2144);
and U6858 (N_6858,N_1452,N_3436);
or U6859 (N_6859,N_3599,N_3458);
or U6860 (N_6860,N_2315,N_3320);
or U6861 (N_6861,N_1121,N_2495);
xor U6862 (N_6862,N_409,N_2066);
nor U6863 (N_6863,N_916,N_535);
nor U6864 (N_6864,N_2868,N_2475);
and U6865 (N_6865,N_2798,N_740);
nor U6866 (N_6866,N_1304,N_994);
and U6867 (N_6867,N_3771,N_3577);
or U6868 (N_6868,N_686,N_380);
and U6869 (N_6869,N_2992,N_3053);
and U6870 (N_6870,N_2149,N_2047);
nor U6871 (N_6871,N_669,N_832);
or U6872 (N_6872,N_1254,N_3690);
and U6873 (N_6873,N_226,N_274);
or U6874 (N_6874,N_749,N_1086);
nor U6875 (N_6875,N_1795,N_3930);
and U6876 (N_6876,N_1084,N_1736);
xor U6877 (N_6877,N_497,N_272);
or U6878 (N_6878,N_3452,N_3070);
nand U6879 (N_6879,N_3710,N_1669);
and U6880 (N_6880,N_2553,N_1666);
and U6881 (N_6881,N_903,N_2298);
and U6882 (N_6882,N_3828,N_1);
nand U6883 (N_6883,N_1634,N_1845);
or U6884 (N_6884,N_2705,N_469);
nor U6885 (N_6885,N_1883,N_1972);
or U6886 (N_6886,N_3529,N_1851);
nor U6887 (N_6887,N_3749,N_1722);
and U6888 (N_6888,N_3672,N_228);
nand U6889 (N_6889,N_455,N_3929);
xnor U6890 (N_6890,N_2299,N_1181);
or U6891 (N_6891,N_1987,N_1122);
or U6892 (N_6892,N_2726,N_3597);
nand U6893 (N_6893,N_2667,N_3093);
nand U6894 (N_6894,N_3326,N_628);
or U6895 (N_6895,N_2350,N_2814);
or U6896 (N_6896,N_1415,N_829);
nand U6897 (N_6897,N_3003,N_1144);
nor U6898 (N_6898,N_2253,N_1428);
nor U6899 (N_6899,N_434,N_3610);
nor U6900 (N_6900,N_2440,N_2077);
and U6901 (N_6901,N_650,N_3120);
nor U6902 (N_6902,N_3112,N_774);
nand U6903 (N_6903,N_3319,N_205);
xor U6904 (N_6904,N_317,N_3606);
nand U6905 (N_6905,N_2322,N_485);
nand U6906 (N_6906,N_3453,N_2829);
nor U6907 (N_6907,N_2792,N_267);
nor U6908 (N_6908,N_3014,N_2333);
nor U6909 (N_6909,N_2190,N_3260);
nor U6910 (N_6910,N_769,N_3558);
or U6911 (N_6911,N_3975,N_3956);
and U6912 (N_6912,N_1511,N_3596);
or U6913 (N_6913,N_524,N_3220);
nand U6914 (N_6914,N_3984,N_3182);
and U6915 (N_6915,N_3818,N_1379);
nor U6916 (N_6916,N_3666,N_3231);
or U6917 (N_6917,N_1733,N_1398);
nand U6918 (N_6918,N_704,N_3295);
and U6919 (N_6919,N_2788,N_2885);
nand U6920 (N_6920,N_2595,N_2624);
nand U6921 (N_6921,N_983,N_3067);
nor U6922 (N_6922,N_2830,N_1170);
or U6923 (N_6923,N_649,N_1780);
nand U6924 (N_6924,N_470,N_809);
and U6925 (N_6925,N_505,N_2905);
and U6926 (N_6926,N_3097,N_2895);
and U6927 (N_6927,N_866,N_1134);
or U6928 (N_6928,N_200,N_3257);
or U6929 (N_6929,N_2403,N_3620);
nor U6930 (N_6930,N_376,N_313);
xor U6931 (N_6931,N_3906,N_1163);
or U6932 (N_6932,N_1079,N_808);
nand U6933 (N_6933,N_3391,N_3238);
and U6934 (N_6934,N_2369,N_2588);
or U6935 (N_6935,N_1453,N_3723);
nor U6936 (N_6936,N_769,N_3606);
and U6937 (N_6937,N_298,N_3614);
xnor U6938 (N_6938,N_688,N_3568);
or U6939 (N_6939,N_3408,N_2474);
or U6940 (N_6940,N_75,N_703);
and U6941 (N_6941,N_1125,N_2946);
nor U6942 (N_6942,N_2831,N_2784);
nor U6943 (N_6943,N_2802,N_2193);
and U6944 (N_6944,N_3201,N_2226);
nand U6945 (N_6945,N_1403,N_3724);
xnor U6946 (N_6946,N_1794,N_3403);
nor U6947 (N_6947,N_701,N_2415);
nand U6948 (N_6948,N_2484,N_3724);
and U6949 (N_6949,N_813,N_1967);
nor U6950 (N_6950,N_3876,N_27);
nand U6951 (N_6951,N_1790,N_3567);
or U6952 (N_6952,N_2739,N_973);
nand U6953 (N_6953,N_1139,N_3739);
nor U6954 (N_6954,N_3881,N_2914);
and U6955 (N_6955,N_490,N_3476);
or U6956 (N_6956,N_392,N_94);
nand U6957 (N_6957,N_1839,N_816);
nand U6958 (N_6958,N_2360,N_1532);
or U6959 (N_6959,N_3451,N_1847);
or U6960 (N_6960,N_38,N_1624);
nor U6961 (N_6961,N_1716,N_856);
xor U6962 (N_6962,N_627,N_2576);
and U6963 (N_6963,N_3864,N_3952);
or U6964 (N_6964,N_572,N_1229);
nor U6965 (N_6965,N_3605,N_18);
or U6966 (N_6966,N_3899,N_2020);
nand U6967 (N_6967,N_1051,N_1674);
or U6968 (N_6968,N_2116,N_461);
nand U6969 (N_6969,N_3381,N_3610);
nor U6970 (N_6970,N_2006,N_1197);
or U6971 (N_6971,N_2641,N_2988);
xnor U6972 (N_6972,N_3104,N_2273);
nor U6973 (N_6973,N_1814,N_2212);
and U6974 (N_6974,N_496,N_833);
nand U6975 (N_6975,N_2582,N_2716);
or U6976 (N_6976,N_3346,N_2311);
or U6977 (N_6977,N_184,N_2935);
nand U6978 (N_6978,N_1148,N_3565);
xnor U6979 (N_6979,N_685,N_2777);
and U6980 (N_6980,N_1270,N_780);
xnor U6981 (N_6981,N_749,N_2738);
nor U6982 (N_6982,N_3817,N_3274);
and U6983 (N_6983,N_3889,N_3575);
or U6984 (N_6984,N_3962,N_1302);
nand U6985 (N_6985,N_2419,N_1922);
nand U6986 (N_6986,N_743,N_3269);
nor U6987 (N_6987,N_2603,N_2509);
nand U6988 (N_6988,N_3656,N_473);
or U6989 (N_6989,N_1741,N_3236);
xnor U6990 (N_6990,N_1979,N_1499);
nand U6991 (N_6991,N_2372,N_3856);
nand U6992 (N_6992,N_3483,N_3065);
and U6993 (N_6993,N_334,N_1231);
nand U6994 (N_6994,N_2362,N_2211);
nor U6995 (N_6995,N_1407,N_3554);
or U6996 (N_6996,N_1496,N_1289);
xor U6997 (N_6997,N_258,N_1995);
and U6998 (N_6998,N_1599,N_3929);
xnor U6999 (N_6999,N_2456,N_184);
or U7000 (N_7000,N_47,N_967);
nand U7001 (N_7001,N_384,N_1397);
nor U7002 (N_7002,N_1538,N_2933);
or U7003 (N_7003,N_2009,N_1295);
or U7004 (N_7004,N_2693,N_1088);
and U7005 (N_7005,N_1838,N_1462);
or U7006 (N_7006,N_1751,N_2736);
and U7007 (N_7007,N_7,N_2052);
nor U7008 (N_7008,N_3387,N_2534);
and U7009 (N_7009,N_2976,N_3138);
nand U7010 (N_7010,N_285,N_2708);
nor U7011 (N_7011,N_898,N_567);
nand U7012 (N_7012,N_906,N_2670);
and U7013 (N_7013,N_2321,N_3863);
and U7014 (N_7014,N_1207,N_386);
nor U7015 (N_7015,N_3316,N_936);
nand U7016 (N_7016,N_2277,N_1734);
nand U7017 (N_7017,N_833,N_1648);
nand U7018 (N_7018,N_3022,N_1921);
xor U7019 (N_7019,N_2926,N_41);
nand U7020 (N_7020,N_144,N_3909);
xnor U7021 (N_7021,N_3318,N_3340);
nor U7022 (N_7022,N_281,N_3824);
nand U7023 (N_7023,N_1468,N_3695);
xnor U7024 (N_7024,N_1844,N_1761);
nor U7025 (N_7025,N_2808,N_2535);
nand U7026 (N_7026,N_3334,N_3094);
nor U7027 (N_7027,N_946,N_2169);
and U7028 (N_7028,N_2192,N_1837);
or U7029 (N_7029,N_2854,N_1461);
and U7030 (N_7030,N_3722,N_128);
nand U7031 (N_7031,N_1672,N_2714);
xnor U7032 (N_7032,N_2735,N_217);
nor U7033 (N_7033,N_513,N_1750);
nand U7034 (N_7034,N_3163,N_2266);
nor U7035 (N_7035,N_1088,N_1898);
nor U7036 (N_7036,N_3059,N_3379);
or U7037 (N_7037,N_2936,N_2256);
or U7038 (N_7038,N_1409,N_2899);
and U7039 (N_7039,N_2067,N_1581);
or U7040 (N_7040,N_2994,N_2310);
nor U7041 (N_7041,N_745,N_1078);
or U7042 (N_7042,N_1600,N_3846);
nor U7043 (N_7043,N_724,N_207);
or U7044 (N_7044,N_3744,N_198);
nand U7045 (N_7045,N_3671,N_469);
nand U7046 (N_7046,N_1411,N_1045);
nand U7047 (N_7047,N_693,N_869);
or U7048 (N_7048,N_835,N_2937);
nor U7049 (N_7049,N_1002,N_2934);
nand U7050 (N_7050,N_141,N_2456);
nand U7051 (N_7051,N_2769,N_1688);
and U7052 (N_7052,N_2519,N_1358);
xnor U7053 (N_7053,N_1217,N_1831);
and U7054 (N_7054,N_3536,N_809);
and U7055 (N_7055,N_2012,N_3972);
or U7056 (N_7056,N_3749,N_1280);
nor U7057 (N_7057,N_2522,N_2993);
or U7058 (N_7058,N_1315,N_2015);
nor U7059 (N_7059,N_3270,N_3292);
and U7060 (N_7060,N_486,N_1516);
xnor U7061 (N_7061,N_3237,N_71);
nand U7062 (N_7062,N_651,N_92);
and U7063 (N_7063,N_3177,N_849);
and U7064 (N_7064,N_3062,N_2799);
nand U7065 (N_7065,N_3462,N_3896);
and U7066 (N_7066,N_1851,N_2132);
xnor U7067 (N_7067,N_3619,N_420);
nand U7068 (N_7068,N_759,N_2152);
and U7069 (N_7069,N_866,N_331);
or U7070 (N_7070,N_2174,N_836);
nor U7071 (N_7071,N_3126,N_3723);
nand U7072 (N_7072,N_2945,N_161);
or U7073 (N_7073,N_3761,N_1091);
or U7074 (N_7074,N_1025,N_2139);
or U7075 (N_7075,N_1081,N_1592);
and U7076 (N_7076,N_3129,N_2450);
xnor U7077 (N_7077,N_1461,N_2163);
nand U7078 (N_7078,N_3876,N_2745);
nand U7079 (N_7079,N_516,N_2708);
and U7080 (N_7080,N_1869,N_807);
or U7081 (N_7081,N_2431,N_1771);
nand U7082 (N_7082,N_102,N_1063);
nand U7083 (N_7083,N_3995,N_1480);
xor U7084 (N_7084,N_3351,N_3653);
nand U7085 (N_7085,N_2412,N_2943);
or U7086 (N_7086,N_628,N_1154);
nand U7087 (N_7087,N_51,N_906);
or U7088 (N_7088,N_1099,N_1790);
and U7089 (N_7089,N_1342,N_38);
nor U7090 (N_7090,N_3376,N_1804);
nand U7091 (N_7091,N_972,N_2887);
or U7092 (N_7092,N_829,N_3418);
xor U7093 (N_7093,N_1982,N_33);
and U7094 (N_7094,N_2659,N_3037);
nand U7095 (N_7095,N_3851,N_573);
xnor U7096 (N_7096,N_757,N_2753);
and U7097 (N_7097,N_1128,N_3682);
nand U7098 (N_7098,N_3382,N_1871);
or U7099 (N_7099,N_461,N_2644);
and U7100 (N_7100,N_783,N_642);
or U7101 (N_7101,N_2200,N_2781);
nand U7102 (N_7102,N_441,N_1153);
or U7103 (N_7103,N_3577,N_2765);
or U7104 (N_7104,N_1348,N_2018);
nand U7105 (N_7105,N_1738,N_3120);
nand U7106 (N_7106,N_2222,N_1883);
nor U7107 (N_7107,N_3508,N_2567);
or U7108 (N_7108,N_1940,N_3963);
or U7109 (N_7109,N_3506,N_3422);
or U7110 (N_7110,N_947,N_3467);
or U7111 (N_7111,N_497,N_2923);
nand U7112 (N_7112,N_3235,N_3921);
nor U7113 (N_7113,N_579,N_2840);
nand U7114 (N_7114,N_1647,N_3665);
nor U7115 (N_7115,N_2086,N_2250);
and U7116 (N_7116,N_2085,N_229);
nor U7117 (N_7117,N_1422,N_192);
and U7118 (N_7118,N_3729,N_678);
and U7119 (N_7119,N_130,N_157);
and U7120 (N_7120,N_22,N_652);
nor U7121 (N_7121,N_3142,N_2429);
or U7122 (N_7122,N_984,N_3166);
and U7123 (N_7123,N_3517,N_2188);
xor U7124 (N_7124,N_137,N_3211);
nor U7125 (N_7125,N_673,N_3844);
nor U7126 (N_7126,N_3122,N_3257);
and U7127 (N_7127,N_3906,N_3700);
and U7128 (N_7128,N_2664,N_751);
and U7129 (N_7129,N_1387,N_1126);
and U7130 (N_7130,N_1104,N_237);
nand U7131 (N_7131,N_2862,N_3180);
nand U7132 (N_7132,N_584,N_3098);
and U7133 (N_7133,N_3544,N_121);
and U7134 (N_7134,N_1378,N_596);
nand U7135 (N_7135,N_3546,N_3398);
xnor U7136 (N_7136,N_3683,N_1123);
nand U7137 (N_7137,N_3043,N_1548);
or U7138 (N_7138,N_3383,N_1896);
and U7139 (N_7139,N_3592,N_1098);
nand U7140 (N_7140,N_3861,N_3143);
and U7141 (N_7141,N_1005,N_3894);
or U7142 (N_7142,N_1564,N_1373);
nor U7143 (N_7143,N_1452,N_2614);
nor U7144 (N_7144,N_3139,N_1522);
and U7145 (N_7145,N_3819,N_2307);
nand U7146 (N_7146,N_2963,N_2541);
xnor U7147 (N_7147,N_2415,N_2677);
nor U7148 (N_7148,N_181,N_2404);
nand U7149 (N_7149,N_3576,N_3824);
nand U7150 (N_7150,N_2289,N_3078);
nand U7151 (N_7151,N_3468,N_3754);
or U7152 (N_7152,N_921,N_2629);
nand U7153 (N_7153,N_1092,N_1591);
and U7154 (N_7154,N_2267,N_3607);
and U7155 (N_7155,N_642,N_3600);
or U7156 (N_7156,N_786,N_385);
or U7157 (N_7157,N_2820,N_2251);
xor U7158 (N_7158,N_1416,N_686);
nor U7159 (N_7159,N_440,N_1634);
xnor U7160 (N_7160,N_2058,N_3369);
or U7161 (N_7161,N_1291,N_3498);
or U7162 (N_7162,N_2751,N_20);
and U7163 (N_7163,N_2939,N_3090);
nand U7164 (N_7164,N_648,N_1096);
and U7165 (N_7165,N_850,N_1638);
nor U7166 (N_7166,N_2056,N_1540);
and U7167 (N_7167,N_1001,N_402);
nand U7168 (N_7168,N_3999,N_398);
nor U7169 (N_7169,N_647,N_2942);
nand U7170 (N_7170,N_46,N_2004);
and U7171 (N_7171,N_470,N_2463);
or U7172 (N_7172,N_2587,N_2212);
xnor U7173 (N_7173,N_2364,N_2150);
or U7174 (N_7174,N_66,N_2869);
or U7175 (N_7175,N_2589,N_1766);
and U7176 (N_7176,N_2726,N_2178);
or U7177 (N_7177,N_367,N_438);
and U7178 (N_7178,N_1067,N_4);
nand U7179 (N_7179,N_1825,N_667);
nand U7180 (N_7180,N_1564,N_2567);
and U7181 (N_7181,N_3658,N_1393);
or U7182 (N_7182,N_1051,N_2320);
or U7183 (N_7183,N_3657,N_2977);
or U7184 (N_7184,N_3430,N_754);
nand U7185 (N_7185,N_1086,N_2759);
nand U7186 (N_7186,N_1500,N_1184);
or U7187 (N_7187,N_3062,N_539);
nand U7188 (N_7188,N_2314,N_690);
nand U7189 (N_7189,N_297,N_690);
or U7190 (N_7190,N_1772,N_1866);
xor U7191 (N_7191,N_990,N_185);
nand U7192 (N_7192,N_3444,N_2556);
nand U7193 (N_7193,N_1147,N_3496);
and U7194 (N_7194,N_2302,N_3998);
xor U7195 (N_7195,N_312,N_133);
xor U7196 (N_7196,N_3075,N_2246);
and U7197 (N_7197,N_2405,N_3522);
and U7198 (N_7198,N_2085,N_1037);
or U7199 (N_7199,N_3869,N_1343);
nor U7200 (N_7200,N_554,N_2789);
and U7201 (N_7201,N_2609,N_3017);
nor U7202 (N_7202,N_809,N_3525);
and U7203 (N_7203,N_2965,N_2137);
nand U7204 (N_7204,N_2991,N_1757);
or U7205 (N_7205,N_1083,N_2439);
xor U7206 (N_7206,N_3287,N_2937);
nor U7207 (N_7207,N_1773,N_1677);
nor U7208 (N_7208,N_3003,N_1671);
or U7209 (N_7209,N_2314,N_2110);
nor U7210 (N_7210,N_2463,N_1986);
and U7211 (N_7211,N_1773,N_3553);
nor U7212 (N_7212,N_3981,N_3685);
and U7213 (N_7213,N_745,N_1606);
or U7214 (N_7214,N_2878,N_3652);
or U7215 (N_7215,N_2269,N_3487);
nor U7216 (N_7216,N_1839,N_3961);
nand U7217 (N_7217,N_2985,N_3739);
and U7218 (N_7218,N_654,N_2606);
nand U7219 (N_7219,N_3424,N_3338);
nand U7220 (N_7220,N_1704,N_98);
or U7221 (N_7221,N_2442,N_495);
nor U7222 (N_7222,N_331,N_511);
and U7223 (N_7223,N_2298,N_1617);
or U7224 (N_7224,N_1504,N_558);
and U7225 (N_7225,N_3452,N_1663);
nor U7226 (N_7226,N_973,N_1933);
and U7227 (N_7227,N_82,N_2370);
or U7228 (N_7228,N_2954,N_488);
nor U7229 (N_7229,N_1092,N_3049);
nor U7230 (N_7230,N_3642,N_1764);
or U7231 (N_7231,N_64,N_2801);
nand U7232 (N_7232,N_861,N_1971);
nor U7233 (N_7233,N_2663,N_1475);
and U7234 (N_7234,N_3708,N_2042);
nor U7235 (N_7235,N_3100,N_3074);
nand U7236 (N_7236,N_3545,N_962);
nor U7237 (N_7237,N_1630,N_607);
nand U7238 (N_7238,N_2615,N_69);
or U7239 (N_7239,N_3204,N_2577);
and U7240 (N_7240,N_2699,N_1959);
or U7241 (N_7241,N_1081,N_134);
and U7242 (N_7242,N_3441,N_3510);
or U7243 (N_7243,N_2659,N_2715);
and U7244 (N_7244,N_839,N_556);
nor U7245 (N_7245,N_788,N_1809);
and U7246 (N_7246,N_2015,N_1889);
and U7247 (N_7247,N_1453,N_3244);
and U7248 (N_7248,N_1676,N_112);
xnor U7249 (N_7249,N_3503,N_156);
or U7250 (N_7250,N_627,N_2198);
and U7251 (N_7251,N_3129,N_718);
or U7252 (N_7252,N_1013,N_934);
nand U7253 (N_7253,N_1394,N_3881);
xnor U7254 (N_7254,N_3308,N_2673);
and U7255 (N_7255,N_3195,N_1334);
or U7256 (N_7256,N_3547,N_1218);
or U7257 (N_7257,N_2060,N_1810);
or U7258 (N_7258,N_2894,N_3271);
or U7259 (N_7259,N_1664,N_1856);
nand U7260 (N_7260,N_1530,N_1788);
nor U7261 (N_7261,N_1018,N_2587);
nor U7262 (N_7262,N_742,N_3670);
nand U7263 (N_7263,N_1849,N_2444);
or U7264 (N_7264,N_1994,N_1725);
or U7265 (N_7265,N_168,N_1916);
nand U7266 (N_7266,N_808,N_3576);
and U7267 (N_7267,N_3965,N_753);
or U7268 (N_7268,N_1500,N_3893);
nor U7269 (N_7269,N_3757,N_2774);
and U7270 (N_7270,N_1757,N_2461);
or U7271 (N_7271,N_501,N_1851);
and U7272 (N_7272,N_1279,N_2298);
xnor U7273 (N_7273,N_2485,N_2753);
or U7274 (N_7274,N_3182,N_796);
or U7275 (N_7275,N_532,N_179);
nor U7276 (N_7276,N_485,N_324);
and U7277 (N_7277,N_3876,N_1811);
nor U7278 (N_7278,N_1586,N_457);
nand U7279 (N_7279,N_2366,N_2076);
or U7280 (N_7280,N_3953,N_792);
nand U7281 (N_7281,N_2439,N_3224);
and U7282 (N_7282,N_3885,N_3110);
nand U7283 (N_7283,N_2428,N_2994);
or U7284 (N_7284,N_2383,N_743);
nor U7285 (N_7285,N_2286,N_3368);
and U7286 (N_7286,N_3360,N_3143);
and U7287 (N_7287,N_217,N_3166);
xor U7288 (N_7288,N_3830,N_1600);
and U7289 (N_7289,N_3216,N_115);
nor U7290 (N_7290,N_3446,N_3509);
nor U7291 (N_7291,N_2912,N_1390);
nand U7292 (N_7292,N_2415,N_2723);
xor U7293 (N_7293,N_3416,N_3272);
or U7294 (N_7294,N_1341,N_307);
nand U7295 (N_7295,N_2774,N_3140);
and U7296 (N_7296,N_824,N_892);
nor U7297 (N_7297,N_1666,N_1859);
or U7298 (N_7298,N_408,N_1703);
xor U7299 (N_7299,N_706,N_961);
or U7300 (N_7300,N_3027,N_48);
or U7301 (N_7301,N_2814,N_2200);
nor U7302 (N_7302,N_1526,N_1378);
and U7303 (N_7303,N_3805,N_3110);
xnor U7304 (N_7304,N_3843,N_1003);
or U7305 (N_7305,N_2088,N_2392);
nand U7306 (N_7306,N_3284,N_958);
nor U7307 (N_7307,N_1554,N_544);
nor U7308 (N_7308,N_2776,N_2000);
nand U7309 (N_7309,N_1992,N_3188);
nor U7310 (N_7310,N_2433,N_1981);
nor U7311 (N_7311,N_73,N_203);
nand U7312 (N_7312,N_3012,N_210);
or U7313 (N_7313,N_2207,N_1899);
nand U7314 (N_7314,N_552,N_1346);
and U7315 (N_7315,N_512,N_653);
or U7316 (N_7316,N_748,N_476);
and U7317 (N_7317,N_3732,N_3337);
nor U7318 (N_7318,N_2688,N_2971);
nand U7319 (N_7319,N_277,N_700);
nand U7320 (N_7320,N_471,N_776);
nor U7321 (N_7321,N_2667,N_1903);
nand U7322 (N_7322,N_3927,N_2719);
xnor U7323 (N_7323,N_1,N_3332);
or U7324 (N_7324,N_464,N_395);
nor U7325 (N_7325,N_569,N_2254);
nor U7326 (N_7326,N_616,N_1043);
xor U7327 (N_7327,N_2375,N_3398);
and U7328 (N_7328,N_279,N_2799);
nand U7329 (N_7329,N_1681,N_3412);
nor U7330 (N_7330,N_911,N_2535);
nor U7331 (N_7331,N_731,N_1749);
xor U7332 (N_7332,N_2032,N_1534);
nand U7333 (N_7333,N_1245,N_1422);
nand U7334 (N_7334,N_162,N_2241);
and U7335 (N_7335,N_3379,N_3509);
or U7336 (N_7336,N_925,N_161);
xor U7337 (N_7337,N_2492,N_661);
nand U7338 (N_7338,N_3646,N_680);
and U7339 (N_7339,N_2778,N_2411);
nand U7340 (N_7340,N_3730,N_1325);
nand U7341 (N_7341,N_3496,N_3131);
or U7342 (N_7342,N_1227,N_2735);
and U7343 (N_7343,N_1188,N_1115);
nand U7344 (N_7344,N_1942,N_2054);
or U7345 (N_7345,N_427,N_3640);
nand U7346 (N_7346,N_3046,N_3494);
nand U7347 (N_7347,N_560,N_2436);
and U7348 (N_7348,N_1085,N_294);
xnor U7349 (N_7349,N_2272,N_3904);
nor U7350 (N_7350,N_3158,N_3678);
nand U7351 (N_7351,N_1144,N_560);
nor U7352 (N_7352,N_3848,N_3955);
nand U7353 (N_7353,N_1356,N_2099);
xor U7354 (N_7354,N_1134,N_401);
nand U7355 (N_7355,N_3445,N_3929);
and U7356 (N_7356,N_1582,N_3095);
and U7357 (N_7357,N_2293,N_2853);
nand U7358 (N_7358,N_1092,N_321);
nor U7359 (N_7359,N_134,N_2815);
nor U7360 (N_7360,N_785,N_546);
and U7361 (N_7361,N_1004,N_2742);
or U7362 (N_7362,N_439,N_3820);
or U7363 (N_7363,N_898,N_3884);
and U7364 (N_7364,N_3394,N_2204);
nand U7365 (N_7365,N_1318,N_1809);
or U7366 (N_7366,N_2703,N_3344);
nor U7367 (N_7367,N_297,N_1746);
nand U7368 (N_7368,N_1553,N_325);
nand U7369 (N_7369,N_432,N_1649);
nand U7370 (N_7370,N_710,N_2958);
nand U7371 (N_7371,N_3905,N_1177);
xnor U7372 (N_7372,N_170,N_3912);
and U7373 (N_7373,N_1585,N_3175);
and U7374 (N_7374,N_2402,N_531);
nor U7375 (N_7375,N_281,N_591);
nand U7376 (N_7376,N_2706,N_2329);
nand U7377 (N_7377,N_3121,N_830);
nor U7378 (N_7378,N_1929,N_2535);
and U7379 (N_7379,N_959,N_2489);
or U7380 (N_7380,N_89,N_958);
and U7381 (N_7381,N_3786,N_2978);
xor U7382 (N_7382,N_695,N_337);
and U7383 (N_7383,N_1764,N_1137);
nand U7384 (N_7384,N_2524,N_1538);
nor U7385 (N_7385,N_1114,N_1749);
nand U7386 (N_7386,N_1118,N_3005);
nand U7387 (N_7387,N_643,N_1154);
nand U7388 (N_7388,N_2697,N_181);
nand U7389 (N_7389,N_193,N_296);
nand U7390 (N_7390,N_2458,N_2035);
nor U7391 (N_7391,N_254,N_355);
and U7392 (N_7392,N_2378,N_1489);
nand U7393 (N_7393,N_2577,N_2827);
nor U7394 (N_7394,N_3393,N_3331);
nand U7395 (N_7395,N_1342,N_1520);
nand U7396 (N_7396,N_3007,N_2377);
nor U7397 (N_7397,N_3164,N_2653);
and U7398 (N_7398,N_1268,N_1910);
and U7399 (N_7399,N_2489,N_1565);
nor U7400 (N_7400,N_167,N_1149);
and U7401 (N_7401,N_3982,N_3316);
and U7402 (N_7402,N_2456,N_2794);
and U7403 (N_7403,N_180,N_428);
nand U7404 (N_7404,N_2696,N_1620);
or U7405 (N_7405,N_3408,N_2221);
nor U7406 (N_7406,N_1367,N_2429);
or U7407 (N_7407,N_1130,N_1800);
and U7408 (N_7408,N_1339,N_1922);
or U7409 (N_7409,N_1938,N_1446);
or U7410 (N_7410,N_3957,N_1660);
nand U7411 (N_7411,N_91,N_27);
xnor U7412 (N_7412,N_1025,N_1794);
xor U7413 (N_7413,N_442,N_38);
xor U7414 (N_7414,N_1641,N_271);
and U7415 (N_7415,N_3165,N_3977);
nand U7416 (N_7416,N_3245,N_507);
xor U7417 (N_7417,N_601,N_3347);
xnor U7418 (N_7418,N_1921,N_2709);
nand U7419 (N_7419,N_2144,N_143);
nand U7420 (N_7420,N_3765,N_2912);
or U7421 (N_7421,N_2928,N_3401);
nand U7422 (N_7422,N_2268,N_3800);
and U7423 (N_7423,N_148,N_2795);
and U7424 (N_7424,N_1409,N_2864);
nor U7425 (N_7425,N_2171,N_62);
nor U7426 (N_7426,N_2716,N_2769);
or U7427 (N_7427,N_2010,N_1005);
nand U7428 (N_7428,N_1815,N_3897);
or U7429 (N_7429,N_1171,N_1828);
or U7430 (N_7430,N_2727,N_1900);
or U7431 (N_7431,N_414,N_116);
nand U7432 (N_7432,N_2082,N_1213);
or U7433 (N_7433,N_2968,N_2432);
nand U7434 (N_7434,N_930,N_3158);
or U7435 (N_7435,N_1676,N_1467);
nor U7436 (N_7436,N_2947,N_1956);
xnor U7437 (N_7437,N_2979,N_3879);
or U7438 (N_7438,N_753,N_533);
or U7439 (N_7439,N_3622,N_511);
and U7440 (N_7440,N_411,N_1350);
nand U7441 (N_7441,N_386,N_2129);
and U7442 (N_7442,N_1739,N_2700);
and U7443 (N_7443,N_3018,N_872);
nand U7444 (N_7444,N_3822,N_3137);
nor U7445 (N_7445,N_2946,N_3498);
nor U7446 (N_7446,N_1314,N_680);
or U7447 (N_7447,N_1282,N_789);
nor U7448 (N_7448,N_2648,N_2424);
or U7449 (N_7449,N_917,N_2749);
or U7450 (N_7450,N_3633,N_2895);
nor U7451 (N_7451,N_566,N_2893);
or U7452 (N_7452,N_930,N_3257);
and U7453 (N_7453,N_1151,N_2857);
or U7454 (N_7454,N_1029,N_3029);
nand U7455 (N_7455,N_1111,N_1794);
nand U7456 (N_7456,N_3555,N_2537);
nor U7457 (N_7457,N_2171,N_2835);
and U7458 (N_7458,N_2983,N_48);
or U7459 (N_7459,N_1814,N_2728);
or U7460 (N_7460,N_1830,N_2660);
or U7461 (N_7461,N_2872,N_1847);
nor U7462 (N_7462,N_2023,N_1508);
nor U7463 (N_7463,N_141,N_3136);
and U7464 (N_7464,N_3790,N_3386);
nor U7465 (N_7465,N_844,N_2509);
and U7466 (N_7466,N_2752,N_2016);
or U7467 (N_7467,N_3492,N_719);
nand U7468 (N_7468,N_1367,N_3313);
nand U7469 (N_7469,N_3793,N_3293);
nand U7470 (N_7470,N_2109,N_354);
xnor U7471 (N_7471,N_1818,N_825);
nand U7472 (N_7472,N_3951,N_1908);
and U7473 (N_7473,N_3573,N_2377);
or U7474 (N_7474,N_2953,N_1302);
nor U7475 (N_7475,N_3213,N_3468);
and U7476 (N_7476,N_37,N_1535);
nor U7477 (N_7477,N_2060,N_111);
nor U7478 (N_7478,N_3967,N_1830);
or U7479 (N_7479,N_818,N_3781);
nand U7480 (N_7480,N_3549,N_290);
or U7481 (N_7481,N_2053,N_2041);
nand U7482 (N_7482,N_8,N_1617);
or U7483 (N_7483,N_3395,N_1027);
nor U7484 (N_7484,N_2363,N_567);
and U7485 (N_7485,N_122,N_2075);
nor U7486 (N_7486,N_1051,N_1958);
nand U7487 (N_7487,N_2651,N_3187);
nand U7488 (N_7488,N_210,N_47);
nor U7489 (N_7489,N_3707,N_1774);
nor U7490 (N_7490,N_3428,N_3394);
and U7491 (N_7491,N_2818,N_3137);
or U7492 (N_7492,N_438,N_741);
and U7493 (N_7493,N_2491,N_1961);
or U7494 (N_7494,N_3289,N_2505);
xnor U7495 (N_7495,N_1259,N_2416);
xor U7496 (N_7496,N_3091,N_2880);
or U7497 (N_7497,N_1597,N_3204);
nor U7498 (N_7498,N_2837,N_735);
nor U7499 (N_7499,N_1083,N_1754);
nand U7500 (N_7500,N_3123,N_1741);
nand U7501 (N_7501,N_1722,N_570);
xnor U7502 (N_7502,N_823,N_3139);
xnor U7503 (N_7503,N_3523,N_2161);
nor U7504 (N_7504,N_149,N_1985);
nand U7505 (N_7505,N_996,N_772);
nand U7506 (N_7506,N_89,N_164);
nor U7507 (N_7507,N_445,N_2354);
and U7508 (N_7508,N_1309,N_123);
and U7509 (N_7509,N_1132,N_3777);
and U7510 (N_7510,N_1928,N_3190);
nand U7511 (N_7511,N_1942,N_3289);
xnor U7512 (N_7512,N_3621,N_1081);
and U7513 (N_7513,N_379,N_1482);
xor U7514 (N_7514,N_2425,N_1576);
and U7515 (N_7515,N_2548,N_2595);
or U7516 (N_7516,N_1665,N_3284);
nand U7517 (N_7517,N_1238,N_3684);
and U7518 (N_7518,N_3299,N_2760);
xor U7519 (N_7519,N_2566,N_378);
or U7520 (N_7520,N_1116,N_2842);
or U7521 (N_7521,N_938,N_981);
and U7522 (N_7522,N_2052,N_841);
nor U7523 (N_7523,N_1664,N_1051);
nor U7524 (N_7524,N_2240,N_2628);
nor U7525 (N_7525,N_2518,N_58);
and U7526 (N_7526,N_2883,N_3174);
or U7527 (N_7527,N_743,N_3250);
or U7528 (N_7528,N_3905,N_1767);
nand U7529 (N_7529,N_1417,N_3326);
xnor U7530 (N_7530,N_73,N_1030);
and U7531 (N_7531,N_2114,N_2994);
xor U7532 (N_7532,N_24,N_1786);
nor U7533 (N_7533,N_3303,N_2953);
or U7534 (N_7534,N_570,N_1935);
or U7535 (N_7535,N_1501,N_3419);
and U7536 (N_7536,N_3101,N_1904);
nand U7537 (N_7537,N_2296,N_3330);
nor U7538 (N_7538,N_3996,N_3869);
xor U7539 (N_7539,N_311,N_2988);
or U7540 (N_7540,N_3463,N_1499);
nand U7541 (N_7541,N_3705,N_2383);
or U7542 (N_7542,N_1501,N_2871);
nand U7543 (N_7543,N_3453,N_1392);
nor U7544 (N_7544,N_2427,N_2133);
and U7545 (N_7545,N_1103,N_2337);
nor U7546 (N_7546,N_2229,N_3742);
nand U7547 (N_7547,N_3069,N_1651);
and U7548 (N_7548,N_886,N_1301);
nand U7549 (N_7549,N_2718,N_2201);
or U7550 (N_7550,N_2111,N_2228);
nand U7551 (N_7551,N_1324,N_740);
and U7552 (N_7552,N_2103,N_2379);
nor U7553 (N_7553,N_3710,N_2266);
nand U7554 (N_7554,N_3276,N_193);
xor U7555 (N_7555,N_1233,N_2155);
nor U7556 (N_7556,N_1775,N_2956);
nor U7557 (N_7557,N_1089,N_11);
xor U7558 (N_7558,N_3220,N_6);
or U7559 (N_7559,N_3994,N_3159);
and U7560 (N_7560,N_3296,N_3734);
and U7561 (N_7561,N_2293,N_2333);
and U7562 (N_7562,N_1783,N_2198);
and U7563 (N_7563,N_498,N_3221);
or U7564 (N_7564,N_1168,N_2348);
nand U7565 (N_7565,N_1343,N_2599);
nand U7566 (N_7566,N_2586,N_2775);
and U7567 (N_7567,N_3229,N_2846);
nand U7568 (N_7568,N_3513,N_3673);
nor U7569 (N_7569,N_811,N_3885);
nor U7570 (N_7570,N_3152,N_1532);
nand U7571 (N_7571,N_1384,N_2394);
nor U7572 (N_7572,N_497,N_611);
nand U7573 (N_7573,N_1396,N_2953);
nor U7574 (N_7574,N_755,N_3945);
or U7575 (N_7575,N_360,N_1747);
xnor U7576 (N_7576,N_759,N_1751);
and U7577 (N_7577,N_3339,N_2393);
and U7578 (N_7578,N_3447,N_3653);
and U7579 (N_7579,N_3684,N_3559);
or U7580 (N_7580,N_1922,N_3159);
and U7581 (N_7581,N_2923,N_2290);
nand U7582 (N_7582,N_744,N_34);
nand U7583 (N_7583,N_2987,N_3827);
and U7584 (N_7584,N_1769,N_251);
xnor U7585 (N_7585,N_789,N_706);
nand U7586 (N_7586,N_789,N_3649);
and U7587 (N_7587,N_2986,N_2994);
or U7588 (N_7588,N_869,N_1551);
and U7589 (N_7589,N_1445,N_108);
nor U7590 (N_7590,N_2556,N_3949);
or U7591 (N_7591,N_3638,N_3937);
nand U7592 (N_7592,N_1091,N_1243);
and U7593 (N_7593,N_293,N_1824);
xor U7594 (N_7594,N_3817,N_2136);
or U7595 (N_7595,N_40,N_2764);
nand U7596 (N_7596,N_1004,N_1257);
nand U7597 (N_7597,N_3560,N_2050);
nor U7598 (N_7598,N_1239,N_1484);
and U7599 (N_7599,N_2794,N_1686);
nand U7600 (N_7600,N_3396,N_761);
xor U7601 (N_7601,N_2621,N_2663);
xnor U7602 (N_7602,N_726,N_3004);
nand U7603 (N_7603,N_2756,N_1141);
and U7604 (N_7604,N_1999,N_2634);
nor U7605 (N_7605,N_1001,N_585);
and U7606 (N_7606,N_936,N_2731);
and U7607 (N_7607,N_3270,N_1975);
nor U7608 (N_7608,N_3304,N_2206);
or U7609 (N_7609,N_1704,N_2557);
and U7610 (N_7610,N_3485,N_3502);
or U7611 (N_7611,N_798,N_875);
nor U7612 (N_7612,N_813,N_1684);
nand U7613 (N_7613,N_1003,N_3926);
xnor U7614 (N_7614,N_3012,N_2796);
xor U7615 (N_7615,N_1330,N_2349);
and U7616 (N_7616,N_503,N_3847);
nand U7617 (N_7617,N_1999,N_857);
nand U7618 (N_7618,N_375,N_2909);
nand U7619 (N_7619,N_1021,N_2689);
and U7620 (N_7620,N_227,N_2355);
xor U7621 (N_7621,N_1640,N_1510);
nor U7622 (N_7622,N_949,N_3543);
or U7623 (N_7623,N_2332,N_2170);
or U7624 (N_7624,N_1805,N_92);
nand U7625 (N_7625,N_3492,N_3730);
nand U7626 (N_7626,N_1141,N_3657);
or U7627 (N_7627,N_3234,N_91);
and U7628 (N_7628,N_517,N_780);
or U7629 (N_7629,N_2735,N_1178);
nand U7630 (N_7630,N_2863,N_1334);
or U7631 (N_7631,N_2545,N_117);
and U7632 (N_7632,N_843,N_1152);
nand U7633 (N_7633,N_339,N_3324);
nor U7634 (N_7634,N_3990,N_3830);
or U7635 (N_7635,N_450,N_171);
or U7636 (N_7636,N_2889,N_2574);
and U7637 (N_7637,N_1037,N_1577);
and U7638 (N_7638,N_346,N_2890);
and U7639 (N_7639,N_81,N_3630);
or U7640 (N_7640,N_560,N_3235);
nand U7641 (N_7641,N_1560,N_3017);
or U7642 (N_7642,N_3990,N_3443);
nand U7643 (N_7643,N_2235,N_3269);
xor U7644 (N_7644,N_2468,N_3383);
nor U7645 (N_7645,N_3587,N_3271);
nand U7646 (N_7646,N_1116,N_2921);
nand U7647 (N_7647,N_3427,N_1339);
or U7648 (N_7648,N_11,N_550);
nor U7649 (N_7649,N_2045,N_1243);
and U7650 (N_7650,N_647,N_631);
or U7651 (N_7651,N_644,N_3369);
xnor U7652 (N_7652,N_2360,N_3016);
nor U7653 (N_7653,N_3039,N_1233);
nor U7654 (N_7654,N_75,N_3359);
nor U7655 (N_7655,N_1284,N_3078);
nor U7656 (N_7656,N_200,N_2939);
or U7657 (N_7657,N_2292,N_1295);
nor U7658 (N_7658,N_2726,N_79);
nor U7659 (N_7659,N_3244,N_1540);
nor U7660 (N_7660,N_3684,N_2221);
and U7661 (N_7661,N_3310,N_1287);
or U7662 (N_7662,N_3344,N_2034);
or U7663 (N_7663,N_3053,N_2930);
or U7664 (N_7664,N_2165,N_1930);
xnor U7665 (N_7665,N_661,N_2358);
and U7666 (N_7666,N_2089,N_869);
and U7667 (N_7667,N_3886,N_1056);
xor U7668 (N_7668,N_178,N_1420);
nand U7669 (N_7669,N_3166,N_3575);
and U7670 (N_7670,N_3177,N_1194);
nand U7671 (N_7671,N_2128,N_2103);
nor U7672 (N_7672,N_317,N_2063);
nand U7673 (N_7673,N_293,N_1056);
or U7674 (N_7674,N_783,N_2618);
or U7675 (N_7675,N_2543,N_574);
nor U7676 (N_7676,N_1734,N_1106);
nand U7677 (N_7677,N_1326,N_2675);
nor U7678 (N_7678,N_794,N_209);
or U7679 (N_7679,N_1285,N_61);
nand U7680 (N_7680,N_2380,N_2452);
or U7681 (N_7681,N_3939,N_524);
and U7682 (N_7682,N_3854,N_3927);
xnor U7683 (N_7683,N_3023,N_3836);
nor U7684 (N_7684,N_1905,N_1017);
nor U7685 (N_7685,N_2135,N_1098);
nand U7686 (N_7686,N_2497,N_1688);
nor U7687 (N_7687,N_1197,N_2184);
or U7688 (N_7688,N_1466,N_1144);
nor U7689 (N_7689,N_594,N_3062);
or U7690 (N_7690,N_925,N_781);
nand U7691 (N_7691,N_848,N_2486);
and U7692 (N_7692,N_2693,N_3849);
nand U7693 (N_7693,N_3008,N_2888);
nor U7694 (N_7694,N_2274,N_1690);
nor U7695 (N_7695,N_660,N_2908);
nor U7696 (N_7696,N_298,N_2227);
nor U7697 (N_7697,N_2866,N_3219);
or U7698 (N_7698,N_1590,N_1944);
nand U7699 (N_7699,N_3393,N_1624);
nand U7700 (N_7700,N_2587,N_1912);
and U7701 (N_7701,N_1857,N_3253);
xnor U7702 (N_7702,N_2818,N_2517);
nor U7703 (N_7703,N_1414,N_2017);
nand U7704 (N_7704,N_728,N_3410);
and U7705 (N_7705,N_568,N_237);
and U7706 (N_7706,N_669,N_2772);
nor U7707 (N_7707,N_1240,N_843);
nor U7708 (N_7708,N_3269,N_320);
or U7709 (N_7709,N_1253,N_245);
and U7710 (N_7710,N_3306,N_123);
nor U7711 (N_7711,N_2172,N_233);
and U7712 (N_7712,N_3631,N_2648);
and U7713 (N_7713,N_676,N_350);
nor U7714 (N_7714,N_150,N_1680);
nor U7715 (N_7715,N_2919,N_3255);
nor U7716 (N_7716,N_2114,N_319);
or U7717 (N_7717,N_2059,N_2340);
and U7718 (N_7718,N_2990,N_828);
nand U7719 (N_7719,N_3793,N_43);
or U7720 (N_7720,N_3147,N_3219);
nand U7721 (N_7721,N_15,N_1818);
or U7722 (N_7722,N_2945,N_423);
or U7723 (N_7723,N_2061,N_609);
nand U7724 (N_7724,N_3061,N_2488);
or U7725 (N_7725,N_386,N_1054);
or U7726 (N_7726,N_1113,N_1276);
xor U7727 (N_7727,N_1863,N_285);
nor U7728 (N_7728,N_3772,N_1839);
and U7729 (N_7729,N_1348,N_2818);
or U7730 (N_7730,N_1340,N_3318);
or U7731 (N_7731,N_1514,N_1778);
and U7732 (N_7732,N_1988,N_2693);
nand U7733 (N_7733,N_559,N_942);
xnor U7734 (N_7734,N_3069,N_873);
xor U7735 (N_7735,N_2756,N_2030);
or U7736 (N_7736,N_3968,N_409);
or U7737 (N_7737,N_3781,N_3214);
or U7738 (N_7738,N_1631,N_1264);
and U7739 (N_7739,N_1146,N_3601);
nand U7740 (N_7740,N_891,N_1121);
and U7741 (N_7741,N_865,N_1244);
xnor U7742 (N_7742,N_3886,N_3595);
xnor U7743 (N_7743,N_2020,N_3825);
nor U7744 (N_7744,N_2505,N_3860);
and U7745 (N_7745,N_975,N_1161);
and U7746 (N_7746,N_140,N_2019);
or U7747 (N_7747,N_114,N_2031);
nand U7748 (N_7748,N_1909,N_1607);
and U7749 (N_7749,N_2199,N_140);
or U7750 (N_7750,N_3160,N_2274);
nand U7751 (N_7751,N_3268,N_3738);
nor U7752 (N_7752,N_3795,N_91);
nor U7753 (N_7753,N_1553,N_1030);
or U7754 (N_7754,N_832,N_1576);
nor U7755 (N_7755,N_3880,N_833);
and U7756 (N_7756,N_1033,N_3874);
and U7757 (N_7757,N_38,N_3020);
and U7758 (N_7758,N_1863,N_2278);
nor U7759 (N_7759,N_3787,N_783);
nor U7760 (N_7760,N_2523,N_2699);
nor U7761 (N_7761,N_151,N_1399);
nand U7762 (N_7762,N_62,N_594);
nor U7763 (N_7763,N_3918,N_3655);
xor U7764 (N_7764,N_204,N_185);
nand U7765 (N_7765,N_3018,N_594);
and U7766 (N_7766,N_1023,N_1977);
and U7767 (N_7767,N_2027,N_1848);
nor U7768 (N_7768,N_1950,N_3381);
and U7769 (N_7769,N_674,N_3542);
nor U7770 (N_7770,N_2536,N_132);
or U7771 (N_7771,N_2726,N_1131);
or U7772 (N_7772,N_758,N_268);
or U7773 (N_7773,N_2576,N_130);
or U7774 (N_7774,N_3182,N_1199);
nand U7775 (N_7775,N_1163,N_2144);
and U7776 (N_7776,N_3896,N_3463);
and U7777 (N_7777,N_3514,N_2434);
nor U7778 (N_7778,N_1160,N_1092);
nand U7779 (N_7779,N_3532,N_461);
and U7780 (N_7780,N_409,N_2550);
nor U7781 (N_7781,N_55,N_960);
or U7782 (N_7782,N_2866,N_3768);
and U7783 (N_7783,N_629,N_1542);
nor U7784 (N_7784,N_148,N_2922);
xnor U7785 (N_7785,N_574,N_2729);
nor U7786 (N_7786,N_2577,N_431);
and U7787 (N_7787,N_1988,N_25);
and U7788 (N_7788,N_3731,N_1144);
or U7789 (N_7789,N_3995,N_2120);
or U7790 (N_7790,N_2479,N_1363);
and U7791 (N_7791,N_3681,N_1550);
nand U7792 (N_7792,N_843,N_2749);
and U7793 (N_7793,N_3255,N_2512);
nor U7794 (N_7794,N_2366,N_3808);
xnor U7795 (N_7795,N_1750,N_2049);
or U7796 (N_7796,N_3404,N_627);
nand U7797 (N_7797,N_1852,N_2541);
or U7798 (N_7798,N_3175,N_409);
nand U7799 (N_7799,N_775,N_3258);
nor U7800 (N_7800,N_3163,N_2404);
nand U7801 (N_7801,N_633,N_553);
nand U7802 (N_7802,N_877,N_1781);
or U7803 (N_7803,N_165,N_2732);
nor U7804 (N_7804,N_191,N_1002);
or U7805 (N_7805,N_1340,N_2384);
or U7806 (N_7806,N_432,N_299);
nand U7807 (N_7807,N_1008,N_2752);
and U7808 (N_7808,N_1938,N_2828);
nand U7809 (N_7809,N_3616,N_1788);
xor U7810 (N_7810,N_3200,N_1150);
nand U7811 (N_7811,N_1119,N_341);
nand U7812 (N_7812,N_2413,N_3767);
xor U7813 (N_7813,N_3456,N_3163);
or U7814 (N_7814,N_1105,N_3716);
and U7815 (N_7815,N_1544,N_2665);
and U7816 (N_7816,N_1208,N_328);
nor U7817 (N_7817,N_3963,N_3922);
nor U7818 (N_7818,N_530,N_1872);
and U7819 (N_7819,N_1388,N_2909);
or U7820 (N_7820,N_1690,N_110);
and U7821 (N_7821,N_1206,N_2173);
nand U7822 (N_7822,N_238,N_801);
nand U7823 (N_7823,N_3334,N_2519);
nand U7824 (N_7824,N_1081,N_2762);
or U7825 (N_7825,N_828,N_3431);
nand U7826 (N_7826,N_1048,N_3366);
xor U7827 (N_7827,N_1076,N_1924);
nor U7828 (N_7828,N_938,N_3512);
and U7829 (N_7829,N_459,N_2099);
or U7830 (N_7830,N_423,N_2307);
xor U7831 (N_7831,N_3388,N_3639);
or U7832 (N_7832,N_2514,N_606);
nand U7833 (N_7833,N_1904,N_132);
nand U7834 (N_7834,N_2951,N_2851);
nand U7835 (N_7835,N_3236,N_3581);
and U7836 (N_7836,N_3930,N_2286);
and U7837 (N_7837,N_689,N_1035);
and U7838 (N_7838,N_3739,N_299);
nand U7839 (N_7839,N_1984,N_3536);
or U7840 (N_7840,N_1696,N_3563);
or U7841 (N_7841,N_3025,N_657);
and U7842 (N_7842,N_2014,N_3863);
or U7843 (N_7843,N_851,N_756);
and U7844 (N_7844,N_3031,N_1939);
and U7845 (N_7845,N_3162,N_1378);
nor U7846 (N_7846,N_1486,N_249);
nor U7847 (N_7847,N_3032,N_3363);
or U7848 (N_7848,N_2797,N_1777);
nand U7849 (N_7849,N_261,N_1779);
nand U7850 (N_7850,N_799,N_3420);
or U7851 (N_7851,N_2112,N_2795);
nand U7852 (N_7852,N_3845,N_1651);
xor U7853 (N_7853,N_394,N_1157);
or U7854 (N_7854,N_2682,N_2426);
or U7855 (N_7855,N_992,N_2557);
nand U7856 (N_7856,N_1534,N_1822);
or U7857 (N_7857,N_3724,N_2430);
nand U7858 (N_7858,N_545,N_304);
nand U7859 (N_7859,N_140,N_1686);
and U7860 (N_7860,N_2,N_389);
nor U7861 (N_7861,N_2891,N_2483);
or U7862 (N_7862,N_805,N_1176);
xor U7863 (N_7863,N_3397,N_3015);
nor U7864 (N_7864,N_3612,N_1901);
and U7865 (N_7865,N_3862,N_2057);
or U7866 (N_7866,N_1427,N_2863);
and U7867 (N_7867,N_2086,N_1464);
and U7868 (N_7868,N_3631,N_1510);
and U7869 (N_7869,N_3205,N_922);
nand U7870 (N_7870,N_341,N_2465);
or U7871 (N_7871,N_367,N_3939);
or U7872 (N_7872,N_2514,N_3673);
and U7873 (N_7873,N_366,N_3150);
nand U7874 (N_7874,N_3404,N_3760);
and U7875 (N_7875,N_2714,N_1814);
or U7876 (N_7876,N_3227,N_285);
nor U7877 (N_7877,N_495,N_1129);
nor U7878 (N_7878,N_73,N_1938);
nor U7879 (N_7879,N_1116,N_1254);
nand U7880 (N_7880,N_2770,N_2835);
nor U7881 (N_7881,N_445,N_613);
or U7882 (N_7882,N_644,N_44);
or U7883 (N_7883,N_3870,N_2152);
and U7884 (N_7884,N_3538,N_2786);
and U7885 (N_7885,N_721,N_3557);
nor U7886 (N_7886,N_3761,N_3731);
and U7887 (N_7887,N_3437,N_2362);
or U7888 (N_7888,N_339,N_1706);
and U7889 (N_7889,N_1919,N_3306);
nor U7890 (N_7890,N_3178,N_1696);
nor U7891 (N_7891,N_84,N_3314);
nand U7892 (N_7892,N_179,N_2368);
or U7893 (N_7893,N_108,N_3979);
nor U7894 (N_7894,N_2599,N_1100);
nor U7895 (N_7895,N_415,N_1777);
and U7896 (N_7896,N_3929,N_832);
nor U7897 (N_7897,N_888,N_135);
nand U7898 (N_7898,N_1750,N_3376);
and U7899 (N_7899,N_1233,N_1861);
or U7900 (N_7900,N_316,N_1072);
nor U7901 (N_7901,N_2089,N_3563);
nand U7902 (N_7902,N_3811,N_732);
nand U7903 (N_7903,N_691,N_1094);
and U7904 (N_7904,N_3525,N_2463);
and U7905 (N_7905,N_3390,N_3378);
and U7906 (N_7906,N_3424,N_3032);
xor U7907 (N_7907,N_2663,N_2406);
nor U7908 (N_7908,N_1557,N_2318);
or U7909 (N_7909,N_313,N_3584);
xnor U7910 (N_7910,N_1137,N_2392);
or U7911 (N_7911,N_3961,N_90);
or U7912 (N_7912,N_2350,N_1350);
and U7913 (N_7913,N_1058,N_3186);
and U7914 (N_7914,N_1715,N_759);
or U7915 (N_7915,N_2118,N_299);
nand U7916 (N_7916,N_1372,N_2082);
xor U7917 (N_7917,N_2375,N_3267);
xnor U7918 (N_7918,N_1009,N_1762);
or U7919 (N_7919,N_2585,N_3694);
nand U7920 (N_7920,N_3694,N_1827);
nor U7921 (N_7921,N_2401,N_3057);
nor U7922 (N_7922,N_2535,N_3561);
and U7923 (N_7923,N_1999,N_146);
xnor U7924 (N_7924,N_1634,N_3773);
nand U7925 (N_7925,N_342,N_3022);
nand U7926 (N_7926,N_2347,N_1520);
nand U7927 (N_7927,N_1987,N_1346);
nor U7928 (N_7928,N_2602,N_2679);
nand U7929 (N_7929,N_3075,N_2785);
or U7930 (N_7930,N_1108,N_1022);
and U7931 (N_7931,N_1144,N_1843);
nand U7932 (N_7932,N_2684,N_3894);
nor U7933 (N_7933,N_310,N_3990);
or U7934 (N_7934,N_1586,N_1202);
xor U7935 (N_7935,N_3203,N_3338);
and U7936 (N_7936,N_1027,N_1958);
or U7937 (N_7937,N_1120,N_3769);
or U7938 (N_7938,N_3499,N_1448);
and U7939 (N_7939,N_20,N_2189);
nor U7940 (N_7940,N_3325,N_1980);
and U7941 (N_7941,N_3841,N_1496);
and U7942 (N_7942,N_3214,N_1303);
or U7943 (N_7943,N_3807,N_1232);
and U7944 (N_7944,N_2410,N_3729);
nor U7945 (N_7945,N_1820,N_131);
and U7946 (N_7946,N_1126,N_2228);
xnor U7947 (N_7947,N_1572,N_3224);
nor U7948 (N_7948,N_3345,N_2871);
and U7949 (N_7949,N_2132,N_1427);
nand U7950 (N_7950,N_3665,N_3518);
or U7951 (N_7951,N_1205,N_3616);
nand U7952 (N_7952,N_3771,N_2194);
xnor U7953 (N_7953,N_2775,N_1253);
nand U7954 (N_7954,N_898,N_2555);
and U7955 (N_7955,N_2100,N_3779);
nand U7956 (N_7956,N_2531,N_737);
xor U7957 (N_7957,N_3218,N_3880);
or U7958 (N_7958,N_136,N_3393);
or U7959 (N_7959,N_535,N_814);
and U7960 (N_7960,N_3406,N_1139);
or U7961 (N_7961,N_1272,N_2335);
nand U7962 (N_7962,N_3131,N_912);
nand U7963 (N_7963,N_2238,N_2038);
nor U7964 (N_7964,N_321,N_3600);
and U7965 (N_7965,N_53,N_2209);
and U7966 (N_7966,N_968,N_3537);
nor U7967 (N_7967,N_1506,N_3633);
nor U7968 (N_7968,N_3697,N_501);
nor U7969 (N_7969,N_1523,N_946);
or U7970 (N_7970,N_1012,N_1185);
or U7971 (N_7971,N_483,N_3306);
and U7972 (N_7972,N_969,N_1024);
and U7973 (N_7973,N_3147,N_601);
and U7974 (N_7974,N_874,N_3448);
and U7975 (N_7975,N_3320,N_3545);
nand U7976 (N_7976,N_307,N_1086);
nand U7977 (N_7977,N_2799,N_951);
nand U7978 (N_7978,N_2006,N_1596);
nand U7979 (N_7979,N_325,N_3075);
nand U7980 (N_7980,N_3111,N_389);
and U7981 (N_7981,N_2836,N_2414);
and U7982 (N_7982,N_1250,N_811);
nand U7983 (N_7983,N_1110,N_3073);
nand U7984 (N_7984,N_2770,N_1626);
nand U7985 (N_7985,N_2176,N_3141);
xnor U7986 (N_7986,N_428,N_2825);
or U7987 (N_7987,N_3154,N_2824);
nor U7988 (N_7988,N_708,N_3128);
nand U7989 (N_7989,N_1477,N_335);
and U7990 (N_7990,N_3608,N_2758);
xnor U7991 (N_7991,N_2288,N_1814);
nor U7992 (N_7992,N_351,N_3582);
or U7993 (N_7993,N_882,N_758);
or U7994 (N_7994,N_2605,N_772);
nor U7995 (N_7995,N_2097,N_1296);
and U7996 (N_7996,N_1840,N_3981);
nand U7997 (N_7997,N_2761,N_2643);
nand U7998 (N_7998,N_3344,N_188);
nor U7999 (N_7999,N_2127,N_275);
and U8000 (N_8000,N_4814,N_7410);
and U8001 (N_8001,N_7003,N_6542);
nand U8002 (N_8002,N_5227,N_6200);
nand U8003 (N_8003,N_5775,N_7538);
or U8004 (N_8004,N_4872,N_5669);
or U8005 (N_8005,N_7101,N_4026);
and U8006 (N_8006,N_7854,N_5839);
nand U8007 (N_8007,N_4428,N_6603);
nand U8008 (N_8008,N_7172,N_4082);
or U8009 (N_8009,N_5467,N_5490);
nor U8010 (N_8010,N_4306,N_4936);
or U8011 (N_8011,N_4281,N_4567);
and U8012 (N_8012,N_7114,N_7887);
nor U8013 (N_8013,N_5951,N_6206);
xor U8014 (N_8014,N_5625,N_7262);
or U8015 (N_8015,N_7122,N_7926);
nand U8016 (N_8016,N_4929,N_6855);
nand U8017 (N_8017,N_4640,N_5434);
or U8018 (N_8018,N_7374,N_5960);
nand U8019 (N_8019,N_6549,N_5177);
and U8020 (N_8020,N_7289,N_7044);
xnor U8021 (N_8021,N_4797,N_7455);
and U8022 (N_8022,N_6686,N_4406);
or U8023 (N_8023,N_6734,N_6198);
nor U8024 (N_8024,N_5794,N_6567);
xor U8025 (N_8025,N_4931,N_5009);
xnor U8026 (N_8026,N_5727,N_5256);
and U8027 (N_8027,N_5380,N_4969);
and U8028 (N_8028,N_6300,N_7297);
or U8029 (N_8029,N_6830,N_5457);
nor U8030 (N_8030,N_6562,N_6294);
nor U8031 (N_8031,N_5972,N_7023);
or U8032 (N_8032,N_7815,N_4246);
nand U8033 (N_8033,N_6307,N_5118);
nor U8034 (N_8034,N_5614,N_6420);
and U8035 (N_8035,N_5500,N_5129);
and U8036 (N_8036,N_7330,N_4351);
and U8037 (N_8037,N_5172,N_6496);
or U8038 (N_8038,N_6279,N_6651);
or U8039 (N_8039,N_4952,N_7770);
and U8040 (N_8040,N_4569,N_5059);
and U8041 (N_8041,N_7591,N_7176);
nor U8042 (N_8042,N_4553,N_6026);
nor U8043 (N_8043,N_6290,N_7655);
and U8044 (N_8044,N_5212,N_7119);
and U8045 (N_8045,N_4417,N_5957);
xnor U8046 (N_8046,N_6762,N_6646);
nand U8047 (N_8047,N_5801,N_4934);
nand U8048 (N_8048,N_7653,N_4008);
nor U8049 (N_8049,N_4856,N_6622);
nor U8050 (N_8050,N_6920,N_5431);
nor U8051 (N_8051,N_5528,N_4470);
nand U8052 (N_8052,N_7737,N_4152);
or U8053 (N_8053,N_5339,N_6856);
or U8054 (N_8054,N_7187,N_6952);
or U8055 (N_8055,N_6505,N_7869);
nor U8056 (N_8056,N_5605,N_4594);
nand U8057 (N_8057,N_6778,N_6040);
and U8058 (N_8058,N_4827,N_5593);
or U8059 (N_8059,N_7664,N_6644);
nor U8060 (N_8060,N_5132,N_5684);
nand U8061 (N_8061,N_4441,N_6400);
nand U8062 (N_8062,N_4398,N_5154);
nor U8063 (N_8063,N_4565,N_5268);
nor U8064 (N_8064,N_5848,N_5984);
and U8065 (N_8065,N_4681,N_4158);
or U8066 (N_8066,N_6370,N_5174);
xor U8067 (N_8067,N_4695,N_4545);
nand U8068 (N_8068,N_7608,N_7442);
xor U8069 (N_8069,N_7163,N_4365);
nor U8070 (N_8070,N_6469,N_4140);
and U8071 (N_8071,N_6218,N_4412);
nor U8072 (N_8072,N_4941,N_7233);
nand U8073 (N_8073,N_6533,N_7429);
and U8074 (N_8074,N_6470,N_7220);
nor U8075 (N_8075,N_6534,N_5947);
and U8076 (N_8076,N_4037,N_4064);
and U8077 (N_8077,N_6342,N_4312);
nand U8078 (N_8078,N_7822,N_5202);
nand U8079 (N_8079,N_7557,N_7102);
and U8080 (N_8080,N_6571,N_7565);
and U8081 (N_8081,N_7371,N_4943);
and U8082 (N_8082,N_5458,N_7049);
nor U8083 (N_8083,N_4182,N_4632);
nand U8084 (N_8084,N_5730,N_6994);
and U8085 (N_8085,N_5538,N_5048);
or U8086 (N_8086,N_7184,N_6833);
nor U8087 (N_8087,N_6663,N_7292);
and U8088 (N_8088,N_7633,N_7996);
nand U8089 (N_8089,N_4072,N_6798);
nand U8090 (N_8090,N_4527,N_7533);
or U8091 (N_8091,N_4546,N_7767);
nand U8092 (N_8092,N_4755,N_4834);
nand U8093 (N_8093,N_7931,N_7701);
and U8094 (N_8094,N_6321,N_4275);
nand U8095 (N_8095,N_7973,N_5636);
and U8096 (N_8096,N_5403,N_4930);
and U8097 (N_8097,N_5231,N_5163);
nand U8098 (N_8098,N_7240,N_6979);
or U8099 (N_8099,N_7331,N_7253);
or U8100 (N_8100,N_6637,N_7775);
nand U8101 (N_8101,N_6234,N_6800);
nand U8102 (N_8102,N_6283,N_7376);
nor U8103 (N_8103,N_7298,N_6878);
or U8104 (N_8104,N_6568,N_4555);
nor U8105 (N_8105,N_6377,N_4539);
nand U8106 (N_8106,N_7211,N_4901);
and U8107 (N_8107,N_5929,N_4124);
or U8108 (N_8108,N_6504,N_7452);
nand U8109 (N_8109,N_6072,N_7158);
or U8110 (N_8110,N_5854,N_4264);
nor U8111 (N_8111,N_5696,N_7895);
or U8112 (N_8112,N_5841,N_5764);
nor U8113 (N_8113,N_6412,N_4986);
nand U8114 (N_8114,N_5567,N_5607);
and U8115 (N_8115,N_6932,N_5498);
nand U8116 (N_8116,N_4487,N_7677);
and U8117 (N_8117,N_6719,N_5548);
or U8118 (N_8118,N_6532,N_6700);
xnor U8119 (N_8119,N_6907,N_7232);
nor U8120 (N_8120,N_7988,N_7636);
nand U8121 (N_8121,N_4022,N_4563);
or U8122 (N_8122,N_5735,N_7803);
nor U8123 (N_8123,N_4902,N_4877);
nor U8124 (N_8124,N_6507,N_7004);
or U8125 (N_8125,N_5452,N_4643);
nor U8126 (N_8126,N_6016,N_4100);
or U8127 (N_8127,N_5524,N_7524);
nor U8128 (N_8128,N_6195,N_6575);
xnor U8129 (N_8129,N_4376,N_6740);
and U8130 (N_8130,N_6069,N_5701);
nor U8131 (N_8131,N_4680,N_6503);
xnor U8132 (N_8132,N_5635,N_7530);
nor U8133 (N_8133,N_4481,N_5550);
or U8134 (N_8134,N_5464,N_5708);
nor U8135 (N_8135,N_7963,N_4085);
xnor U8136 (N_8136,N_5111,N_6476);
xnor U8137 (N_8137,N_5127,N_4666);
nand U8138 (N_8138,N_6695,N_5942);
nand U8139 (N_8139,N_4244,N_6940);
nor U8140 (N_8140,N_7362,N_7234);
nor U8141 (N_8141,N_4792,N_5294);
and U8142 (N_8142,N_6906,N_4075);
nand U8143 (N_8143,N_7348,N_6196);
nor U8144 (N_8144,N_6067,N_4213);
or U8145 (N_8145,N_7553,N_5358);
nor U8146 (N_8146,N_7542,N_5874);
or U8147 (N_8147,N_6024,N_4875);
nor U8148 (N_8148,N_6553,N_7175);
or U8149 (N_8149,N_6311,N_5442);
and U8150 (N_8150,N_4864,N_7453);
nand U8151 (N_8151,N_6772,N_5257);
xor U8152 (N_8152,N_4132,N_7169);
and U8153 (N_8153,N_7467,N_6053);
nor U8154 (N_8154,N_4884,N_6688);
and U8155 (N_8155,N_5752,N_7190);
nand U8156 (N_8156,N_6669,N_5046);
nand U8157 (N_8157,N_6039,N_4445);
and U8158 (N_8158,N_4767,N_4352);
and U8159 (N_8159,N_7311,N_5852);
nor U8160 (N_8160,N_7900,N_4204);
nor U8161 (N_8161,N_6965,N_4329);
and U8162 (N_8162,N_7614,N_4368);
nand U8163 (N_8163,N_4103,N_4853);
nor U8164 (N_8164,N_7412,N_6015);
and U8165 (N_8165,N_5811,N_7941);
nand U8166 (N_8166,N_5650,N_4747);
nor U8167 (N_8167,N_6025,N_7920);
nor U8168 (N_8168,N_4566,N_6705);
nand U8169 (N_8169,N_5312,N_4704);
and U8170 (N_8170,N_6163,N_5072);
or U8171 (N_8171,N_4341,N_5782);
and U8172 (N_8172,N_5050,N_6779);
nand U8173 (N_8173,N_6808,N_5749);
and U8174 (N_8174,N_7302,N_5751);
or U8175 (N_8175,N_4232,N_7250);
nor U8176 (N_8176,N_5617,N_6433);
and U8177 (N_8177,N_7112,N_5119);
and U8178 (N_8178,N_7054,N_4089);
or U8179 (N_8179,N_4160,N_5738);
and U8180 (N_8180,N_5105,N_4739);
xor U8181 (N_8181,N_4635,N_6713);
or U8182 (N_8182,N_5913,N_5864);
nand U8183 (N_8183,N_7078,N_7590);
xnor U8184 (N_8184,N_4699,N_6112);
or U8185 (N_8185,N_4027,N_4314);
xor U8186 (N_8186,N_4354,N_7487);
or U8187 (N_8187,N_6736,N_7280);
nor U8188 (N_8188,N_6879,N_5188);
and U8189 (N_8189,N_7108,N_4965);
and U8190 (N_8190,N_4679,N_5685);
nand U8191 (N_8191,N_7583,N_5598);
nand U8192 (N_8192,N_7508,N_7823);
and U8193 (N_8193,N_4601,N_7087);
or U8194 (N_8194,N_7831,N_5399);
or U8195 (N_8195,N_7623,N_6102);
xor U8196 (N_8196,N_4791,N_6814);
xor U8197 (N_8197,N_5281,N_4274);
xnor U8198 (N_8198,N_5624,N_5646);
or U8199 (N_8199,N_6452,N_7732);
and U8200 (N_8200,N_6353,N_7314);
and U8201 (N_8201,N_6293,N_4266);
nor U8202 (N_8202,N_4909,N_5580);
or U8203 (N_8203,N_4229,N_6537);
xnor U8204 (N_8204,N_7705,N_7989);
nand U8205 (N_8205,N_6891,N_5899);
or U8206 (N_8206,N_6619,N_5015);
nand U8207 (N_8207,N_5954,N_7759);
or U8208 (N_8208,N_5195,N_4967);
and U8209 (N_8209,N_6822,N_4725);
and U8210 (N_8210,N_5812,N_4393);
nor U8211 (N_8211,N_6369,N_5974);
or U8212 (N_8212,N_4392,N_6423);
or U8213 (N_8213,N_5475,N_6550);
nand U8214 (N_8214,N_5169,N_7347);
or U8215 (N_8215,N_7971,N_5832);
or U8216 (N_8216,N_7486,N_7343);
xnor U8217 (N_8217,N_4590,N_7497);
or U8218 (N_8218,N_6010,N_5769);
and U8219 (N_8219,N_7084,N_7230);
and U8220 (N_8220,N_5338,N_5734);
nand U8221 (N_8221,N_5897,N_7231);
xor U8222 (N_8222,N_5706,N_6512);
nand U8223 (N_8223,N_7121,N_5631);
or U8224 (N_8224,N_6836,N_6557);
nand U8225 (N_8225,N_7662,N_6639);
or U8226 (N_8226,N_4099,N_6632);
xor U8227 (N_8227,N_6511,N_4299);
nand U8228 (N_8228,N_5497,N_6928);
or U8229 (N_8229,N_7788,N_7974);
or U8230 (N_8230,N_6209,N_6210);
nor U8231 (N_8231,N_6176,N_7011);
nand U8232 (N_8232,N_7088,N_6388);
nand U8233 (N_8233,N_5340,N_7689);
nor U8234 (N_8234,N_7960,N_5262);
nor U8235 (N_8235,N_7561,N_6410);
or U8236 (N_8236,N_6122,N_5937);
nand U8237 (N_8237,N_7765,N_6642);
nor U8238 (N_8238,N_7801,N_4030);
nand U8239 (N_8239,N_7312,N_5980);
xnor U8240 (N_8240,N_4012,N_7946);
nor U8241 (N_8241,N_6662,N_4477);
nand U8242 (N_8242,N_5757,N_4198);
nor U8243 (N_8243,N_6472,N_7914);
nor U8244 (N_8244,N_7321,N_6819);
and U8245 (N_8245,N_5896,N_5482);
or U8246 (N_8246,N_7554,N_4781);
xor U8247 (N_8247,N_5559,N_4826);
xnor U8248 (N_8248,N_7758,N_6244);
xor U8249 (N_8249,N_6076,N_7364);
and U8250 (N_8250,N_4221,N_6109);
and U8251 (N_8251,N_7644,N_5133);
xnor U8252 (N_8252,N_7304,N_6934);
nand U8253 (N_8253,N_6881,N_6591);
and U8254 (N_8254,N_4507,N_6860);
and U8255 (N_8255,N_7413,N_7764);
nand U8256 (N_8256,N_7391,N_6461);
nor U8257 (N_8257,N_5962,N_4911);
and U8258 (N_8258,N_6893,N_4631);
nor U8259 (N_8259,N_4706,N_5224);
or U8260 (N_8260,N_5055,N_4663);
and U8261 (N_8261,N_7275,N_5967);
or U8262 (N_8262,N_4789,N_6242);
nand U8263 (N_8263,N_6479,N_7451);
and U8264 (N_8264,N_7193,N_4651);
nand U8265 (N_8265,N_6670,N_4520);
nor U8266 (N_8266,N_7249,N_6429);
nor U8267 (N_8267,N_4709,N_7006);
and U8268 (N_8268,N_7773,N_4482);
nand U8269 (N_8269,N_5779,N_6785);
or U8270 (N_8270,N_6839,N_4147);
nor U8271 (N_8271,N_7474,N_7685);
nor U8272 (N_8272,N_5400,N_7028);
and U8273 (N_8273,N_4937,N_5008);
nor U8274 (N_8274,N_6137,N_4010);
and U8275 (N_8275,N_5741,N_6153);
or U8276 (N_8276,N_7604,N_6909);
and U8277 (N_8277,N_6925,N_5337);
nor U8278 (N_8278,N_6330,N_7625);
or U8279 (N_8279,N_5756,N_7483);
or U8280 (N_8280,N_7651,N_6228);
nand U8281 (N_8281,N_6277,N_4025);
or U8282 (N_8282,N_6313,N_5043);
and U8283 (N_8283,N_4407,N_6285);
or U8284 (N_8284,N_6368,N_7837);
or U8285 (N_8285,N_5437,N_6960);
nor U8286 (N_8286,N_5014,N_5686);
nor U8287 (N_8287,N_4038,N_4782);
nor U8288 (N_8288,N_6378,N_4637);
nor U8289 (N_8289,N_6043,N_4247);
nor U8290 (N_8290,N_5608,N_5217);
nor U8291 (N_8291,N_7186,N_5153);
and U8292 (N_8292,N_7891,N_6077);
and U8293 (N_8293,N_4705,N_5724);
nor U8294 (N_8294,N_5597,N_5481);
xor U8295 (N_8295,N_5890,N_5867);
nand U8296 (N_8296,N_5547,N_6233);
or U8297 (N_8297,N_6292,N_7276);
nor U8298 (N_8298,N_6308,N_7159);
nand U8299 (N_8299,N_6064,N_5626);
and U8300 (N_8300,N_6379,N_7296);
and U8301 (N_8301,N_4815,N_7880);
and U8302 (N_8302,N_5152,N_7301);
nand U8303 (N_8303,N_6821,N_4307);
xor U8304 (N_8304,N_7050,N_6851);
or U8305 (N_8305,N_6463,N_7043);
and U8306 (N_8306,N_4169,N_4040);
or U8307 (N_8307,N_4494,N_5875);
and U8308 (N_8308,N_6185,N_7587);
nand U8309 (N_8309,N_7185,N_6494);
nor U8310 (N_8310,N_7723,N_5728);
nand U8311 (N_8311,N_6780,N_5615);
nand U8312 (N_8312,N_7797,N_6600);
and U8313 (N_8313,N_7045,N_6075);
nor U8314 (N_8314,N_4984,N_7799);
or U8315 (N_8315,N_7990,N_6214);
nand U8316 (N_8316,N_6212,N_6992);
nand U8317 (N_8317,N_5139,N_6011);
or U8318 (N_8318,N_7581,N_7541);
and U8319 (N_8319,N_6224,N_6145);
nor U8320 (N_8320,N_5765,N_4650);
nand U8321 (N_8321,N_6304,N_4642);
nor U8322 (N_8322,N_4728,N_5637);
nor U8323 (N_8323,N_5923,N_6817);
nand U8324 (N_8324,N_6708,N_7760);
xnor U8325 (N_8325,N_6968,N_7513);
or U8326 (N_8326,N_4390,N_4868);
nand U8327 (N_8327,N_6682,N_4079);
nor U8328 (N_8328,N_6601,N_5377);
or U8329 (N_8329,N_4536,N_7130);
nand U8330 (N_8330,N_7879,N_4034);
nand U8331 (N_8331,N_7389,N_6993);
or U8332 (N_8332,N_6106,N_5526);
xor U8333 (N_8333,N_6126,N_4784);
nand U8334 (N_8334,N_5304,N_5300);
and U8335 (N_8335,N_5633,N_6060);
nor U8336 (N_8336,N_7809,N_4619);
and U8337 (N_8337,N_7569,N_5440);
and U8338 (N_8338,N_6747,N_6787);
and U8339 (N_8339,N_5030,N_6358);
nand U8340 (N_8340,N_7603,N_4155);
nor U8341 (N_8341,N_7325,N_4225);
nand U8342 (N_8342,N_5351,N_7074);
xor U8343 (N_8343,N_7428,N_5991);
and U8344 (N_8344,N_5258,N_7221);
nand U8345 (N_8345,N_7745,N_4211);
and U8346 (N_8346,N_7222,N_6248);
nand U8347 (N_8347,N_5206,N_7703);
nand U8348 (N_8348,N_4774,N_7420);
nor U8349 (N_8349,N_4907,N_5423);
nand U8350 (N_8350,N_4134,N_5641);
xor U8351 (N_8351,N_6792,N_4059);
nor U8352 (N_8352,N_4763,N_7807);
or U8353 (N_8353,N_4164,N_5630);
nor U8354 (N_8354,N_6659,N_4935);
xnor U8355 (N_8355,N_7372,N_7787);
xor U8356 (N_8356,N_6487,N_6046);
and U8357 (N_8357,N_7268,N_4605);
or U8358 (N_8358,N_5681,N_7440);
nor U8359 (N_8359,N_4556,N_4421);
xnor U8360 (N_8360,N_4948,N_5697);
nand U8361 (N_8361,N_7238,N_6019);
nand U8362 (N_8362,N_5928,N_7000);
and U8363 (N_8363,N_4703,N_4617);
nor U8364 (N_8364,N_6773,N_6416);
nor U8365 (N_8365,N_6730,N_7008);
nand U8366 (N_8366,N_5619,N_7728);
or U8367 (N_8367,N_7978,N_4693);
or U8368 (N_8368,N_6633,N_7772);
or U8369 (N_8369,N_6973,N_7991);
xnor U8370 (N_8370,N_5422,N_4707);
nor U8371 (N_8371,N_4121,N_4294);
nand U8372 (N_8372,N_4777,N_6152);
and U8373 (N_8373,N_6157,N_5901);
or U8374 (N_8374,N_6021,N_6759);
xor U8375 (N_8375,N_5535,N_7719);
nand U8376 (N_8376,N_7896,N_5705);
and U8377 (N_8377,N_5505,N_4738);
nor U8378 (N_8378,N_6698,N_5193);
and U8379 (N_8379,N_5964,N_6052);
nor U8380 (N_8380,N_5448,N_7925);
nor U8381 (N_8381,N_6402,N_5621);
and U8382 (N_8382,N_5021,N_6832);
nor U8383 (N_8383,N_4687,N_5917);
nand U8384 (N_8384,N_7066,N_4544);
and U8385 (N_8385,N_7933,N_6240);
nor U8386 (N_8386,N_7295,N_4595);
nand U8387 (N_8387,N_7432,N_4073);
or U8388 (N_8388,N_5003,N_5391);
or U8389 (N_8389,N_6767,N_6204);
xor U8390 (N_8390,N_7962,N_7444);
and U8391 (N_8391,N_7443,N_4906);
and U8392 (N_8392,N_7063,N_4971);
nor U8393 (N_8393,N_5767,N_6845);
nor U8394 (N_8394,N_6810,N_4230);
or U8395 (N_8395,N_5570,N_4411);
nor U8396 (N_8396,N_6529,N_4682);
nand U8397 (N_8397,N_6750,N_4587);
xor U8398 (N_8398,N_5024,N_6205);
nor U8399 (N_8399,N_6260,N_6437);
nand U8400 (N_8400,N_4095,N_7714);
nor U8401 (N_8401,N_6193,N_4807);
nand U8402 (N_8402,N_5830,N_7954);
and U8403 (N_8403,N_7414,N_4235);
nand U8404 (N_8404,N_6811,N_4113);
or U8405 (N_8405,N_5502,N_5190);
xor U8406 (N_8406,N_7790,N_4916);
nand U8407 (N_8407,N_5722,N_7987);
nand U8408 (N_8408,N_7142,N_6162);
or U8409 (N_8409,N_4018,N_7782);
or U8410 (N_8410,N_4652,N_7201);
nor U8411 (N_8411,N_4118,N_6971);
xor U8412 (N_8412,N_6919,N_5911);
nor U8413 (N_8413,N_5125,N_7143);
nand U8414 (N_8414,N_7940,N_7713);
nor U8415 (N_8415,N_5813,N_4440);
xnor U8416 (N_8416,N_5647,N_4626);
nand U8417 (N_8417,N_6013,N_6958);
or U8418 (N_8418,N_5711,N_5350);
nand U8419 (N_8419,N_4263,N_7021);
and U8420 (N_8420,N_6607,N_7173);
or U8421 (N_8421,N_5495,N_6339);
or U8422 (N_8422,N_7965,N_6626);
nand U8423 (N_8423,N_4885,N_6357);
nor U8424 (N_8424,N_5894,N_5302);
nand U8425 (N_8425,N_4753,N_7840);
or U8426 (N_8426,N_6667,N_6638);
nand U8427 (N_8427,N_4240,N_5873);
nor U8428 (N_8428,N_6521,N_5925);
or U8429 (N_8429,N_5755,N_6314);
nor U8430 (N_8430,N_4498,N_6774);
nor U8431 (N_8431,N_5726,N_6790);
nor U8432 (N_8432,N_5750,N_5595);
nand U8433 (N_8433,N_5429,N_4394);
nor U8434 (N_8434,N_6390,N_5795);
xor U8435 (N_8435,N_7320,N_7017);
or U8436 (N_8436,N_7085,N_5223);
or U8437 (N_8437,N_6876,N_5904);
nor U8438 (N_8438,N_6381,N_7421);
and U8439 (N_8439,N_4262,N_5222);
or U8440 (N_8440,N_6628,N_5247);
nand U8441 (N_8441,N_5924,N_7205);
nor U8442 (N_8442,N_5250,N_5093);
nor U8443 (N_8443,N_5920,N_5887);
nand U8444 (N_8444,N_5889,N_4195);
nand U8445 (N_8445,N_6961,N_7069);
nand U8446 (N_8446,N_7318,N_5562);
nor U8447 (N_8447,N_5978,N_6904);
nand U8448 (N_8448,N_4522,N_5936);
xnor U8449 (N_8449,N_7329,N_6177);
or U8450 (N_8450,N_6658,N_4088);
and U8451 (N_8451,N_5472,N_4254);
and U8452 (N_8452,N_4702,N_5506);
xnor U8453 (N_8453,N_6265,N_4768);
and U8454 (N_8454,N_7096,N_6386);
and U8455 (N_8455,N_6278,N_7751);
nand U8456 (N_8456,N_5800,N_4028);
nor U8457 (N_8457,N_4379,N_5766);
and U8458 (N_8458,N_4530,N_7715);
and U8459 (N_8459,N_4883,N_5488);
or U8460 (N_8460,N_5656,N_5368);
nand U8461 (N_8461,N_5419,N_4963);
nor U8462 (N_8462,N_7917,N_6841);
and U8463 (N_8463,N_4372,N_6333);
nor U8464 (N_8464,N_5687,N_5604);
nor U8465 (N_8465,N_4296,N_4525);
and U8466 (N_8466,N_6485,N_4043);
nand U8467 (N_8467,N_5989,N_6718);
nor U8468 (N_8468,N_7607,N_6846);
or U8469 (N_8469,N_4449,N_5087);
nor U8470 (N_8470,N_7858,N_7830);
nor U8471 (N_8471,N_6871,N_5791);
and U8472 (N_8472,N_7682,N_7824);
and U8473 (N_8473,N_6144,N_6345);
nand U8474 (N_8474,N_5494,N_7447);
nand U8475 (N_8475,N_5371,N_5225);
and U8476 (N_8476,N_7881,N_7402);
and U8477 (N_8477,N_5715,N_5820);
xor U8478 (N_8478,N_5886,N_6227);
nand U8479 (N_8479,N_4190,N_7191);
and U8480 (N_8480,N_6048,N_5205);
or U8481 (N_8481,N_6825,N_7258);
nand U8482 (N_8482,N_5365,N_7843);
and U8483 (N_8483,N_6419,N_5306);
and U8484 (N_8484,N_5688,N_7073);
or U8485 (N_8485,N_5639,N_4492);
or U8486 (N_8486,N_4241,N_4286);
nor U8487 (N_8487,N_7210,N_7810);
and U8488 (N_8488,N_7194,N_5450);
and U8489 (N_8489,N_7055,N_7150);
and U8490 (N_8490,N_5314,N_4933);
and U8491 (N_8491,N_4416,N_4871);
and U8492 (N_8492,N_6953,N_4496);
and U8493 (N_8493,N_6241,N_6944);
or U8494 (N_8494,N_5141,N_4616);
nand U8495 (N_8495,N_7617,N_5233);
or U8496 (N_8496,N_5071,N_5965);
or U8497 (N_8497,N_7407,N_7161);
or U8498 (N_8498,N_4196,N_6763);
and U8499 (N_8499,N_7986,N_4451);
or U8500 (N_8500,N_4427,N_6924);
or U8501 (N_8501,N_5388,N_4759);
nand U8502 (N_8502,N_4511,N_6018);
and U8503 (N_8503,N_4997,N_7979);
and U8504 (N_8504,N_6156,N_5941);
nor U8505 (N_8505,N_7937,N_7666);
nor U8506 (N_8506,N_6595,N_7919);
and U8507 (N_8507,N_5287,N_4357);
or U8508 (N_8508,N_4456,N_6098);
xor U8509 (N_8509,N_6252,N_5968);
nor U8510 (N_8510,N_4272,N_4023);
xor U8511 (N_8511,N_4310,N_4094);
and U8512 (N_8512,N_4108,N_7835);
nand U8513 (N_8513,N_6579,N_6257);
nand U8514 (N_8514,N_6374,N_6858);
or U8515 (N_8515,N_4850,N_7450);
nor U8516 (N_8516,N_6783,N_6775);
and U8517 (N_8517,N_4953,N_5085);
and U8518 (N_8518,N_6927,N_5778);
and U8519 (N_8519,N_4570,N_6050);
and U8520 (N_8520,N_4636,N_7997);
nor U8521 (N_8521,N_6207,N_6312);
and U8522 (N_8522,N_7315,N_7378);
nor U8523 (N_8523,N_5919,N_7943);
or U8524 (N_8524,N_6362,N_7248);
or U8525 (N_8525,N_6124,N_6617);
nand U8526 (N_8526,N_4319,N_7848);
xor U8527 (N_8527,N_5863,N_4597);
or U8528 (N_8528,N_5719,N_6289);
nor U8529 (N_8529,N_7105,N_7873);
or U8530 (N_8530,N_5264,N_7503);
nand U8531 (N_8531,N_7610,N_5806);
and U8532 (N_8532,N_5215,N_5918);
or U8533 (N_8533,N_4921,N_6459);
and U8534 (N_8534,N_6753,N_6336);
and U8535 (N_8535,N_4574,N_7380);
nand U8536 (N_8536,N_4289,N_5644);
nor U8537 (N_8537,N_4946,N_4165);
or U8538 (N_8538,N_6888,N_5409);
and U8539 (N_8539,N_6148,N_6007);
or U8540 (N_8540,N_5274,N_6382);
nor U8541 (N_8541,N_6062,N_5849);
nand U8542 (N_8542,N_7392,N_7601);
and U8543 (N_8543,N_7555,N_7183);
xor U8544 (N_8544,N_7821,N_6375);
nor U8545 (N_8545,N_6477,N_7706);
nand U8546 (N_8546,N_7681,N_5040);
nor U8547 (N_8547,N_6405,N_5326);
xor U8548 (N_8548,N_6384,N_5785);
nand U8549 (N_8549,N_5704,N_4191);
nor U8550 (N_8550,N_4716,N_4991);
nor U8551 (N_8551,N_4339,N_5914);
and U8552 (N_8552,N_4894,N_4248);
nand U8553 (N_8553,N_5817,N_4389);
or U8554 (N_8554,N_5492,N_5731);
and U8555 (N_8555,N_5699,N_5138);
nor U8556 (N_8556,N_6643,N_5760);
and U8557 (N_8557,N_6418,N_7132);
xnor U8558 (N_8558,N_5483,N_5100);
xor U8559 (N_8559,N_7398,N_4343);
and U8560 (N_8560,N_4848,N_5575);
nand U8561 (N_8561,N_5844,N_5983);
nand U8562 (N_8562,N_4348,N_7437);
nor U8563 (N_8563,N_6742,N_7646);
or U8564 (N_8564,N_4446,N_6366);
and U8565 (N_8565,N_6894,N_6866);
xor U8566 (N_8566,N_7261,N_4585);
nor U8567 (N_8567,N_5108,N_5342);
nand U8568 (N_8568,N_5558,N_5855);
or U8569 (N_8569,N_7104,N_7634);
nand U8570 (N_8570,N_6587,N_7227);
or U8571 (N_8571,N_4698,N_4301);
nor U8572 (N_8572,N_4880,N_7279);
and U8573 (N_8573,N_6475,N_7040);
or U8574 (N_8574,N_7504,N_7097);
nor U8575 (N_8575,N_6840,N_6396);
nor U8576 (N_8576,N_6097,N_7079);
or U8577 (N_8577,N_7826,N_4656);
xor U8578 (N_8578,N_5572,N_6267);
nand U8579 (N_8579,N_7427,N_5948);
or U8580 (N_8580,N_4861,N_4193);
nor U8581 (N_8581,N_6031,N_6082);
nand U8582 (N_8582,N_5235,N_4168);
or U8583 (N_8583,N_7813,N_4171);
nor U8584 (N_8584,N_4057,N_7899);
and U8585 (N_8585,N_6355,N_6442);
and U8586 (N_8586,N_5045,N_6035);
nand U8587 (N_8587,N_7307,N_7585);
nor U8588 (N_8588,N_4962,N_6946);
nand U8589 (N_8589,N_5523,N_5213);
or U8590 (N_8590,N_6678,N_4292);
nand U8591 (N_8591,N_4490,N_5420);
nor U8592 (N_8592,N_6722,N_7235);
nor U8593 (N_8593,N_4485,N_7334);
and U8594 (N_8594,N_6034,N_7690);
nand U8595 (N_8595,N_7589,N_6818);
nor U8596 (N_8596,N_6738,N_4519);
xor U8597 (N_8597,N_4397,N_5555);
or U8598 (N_8598,N_5328,N_7856);
nand U8599 (N_8599,N_4086,N_5616);
and U8600 (N_8600,N_4245,N_5075);
xnor U8601 (N_8601,N_6739,N_4957);
or U8602 (N_8602,N_5311,N_5796);
and U8603 (N_8603,N_6497,N_4423);
or U8604 (N_8604,N_5892,N_7139);
or U8605 (N_8605,N_5518,N_7725);
xnor U8606 (N_8606,N_4150,N_6444);
and U8607 (N_8607,N_5052,N_7052);
nand U8608 (N_8608,N_6236,N_7667);
and U8609 (N_8609,N_4276,N_6618);
xor U8610 (N_8610,N_7597,N_5561);
nand U8611 (N_8611,N_5296,N_5496);
nand U8612 (N_8612,N_5987,N_7415);
or U8613 (N_8613,N_7403,N_4197);
or U8614 (N_8614,N_4091,N_4672);
nor U8615 (N_8615,N_6939,N_4144);
nor U8616 (N_8616,N_5185,N_7160);
or U8617 (N_8617,N_6191,N_4212);
or U8618 (N_8618,N_4015,N_4315);
nand U8619 (N_8619,N_6142,N_5916);
nor U8620 (N_8620,N_6583,N_7918);
xnor U8621 (N_8621,N_7902,N_4994);
nor U8622 (N_8622,N_7113,N_4977);
and U8623 (N_8623,N_4751,N_5946);
or U8624 (N_8624,N_4665,N_6572);
or U8625 (N_8625,N_4500,N_4316);
and U8626 (N_8626,N_4497,N_5985);
and U8627 (N_8627,N_5479,N_6984);
and U8628 (N_8628,N_6945,N_7016);
nand U8629 (N_8629,N_4216,N_5465);
and U8630 (N_8630,N_5432,N_6235);
nor U8631 (N_8631,N_5799,N_6500);
or U8632 (N_8632,N_7181,N_5444);
or U8633 (N_8633,N_4208,N_4534);
and U8634 (N_8634,N_5861,N_6699);
nand U8635 (N_8635,N_4899,N_7424);
or U8636 (N_8636,N_6393,N_7540);
xor U8637 (N_8637,N_6096,N_7224);
nand U8638 (N_8638,N_4926,N_4334);
nand U8639 (N_8639,N_7468,N_7560);
nand U8640 (N_8640,N_5988,N_6868);
nand U8641 (N_8641,N_6581,N_4471);
or U8642 (N_8642,N_7659,N_4639);
nor U8643 (N_8643,N_5891,N_5712);
nand U8644 (N_8644,N_6723,N_5123);
nor U8645 (N_8645,N_6823,N_4898);
nand U8646 (N_8646,N_5197,N_6140);
or U8647 (N_8647,N_6178,N_4420);
or U8648 (N_8648,N_5025,N_7739);
nand U8649 (N_8649,N_7922,N_6802);
and U8650 (N_8650,N_5449,N_5563);
xnor U8651 (N_8651,N_5898,N_4603);
and U8652 (N_8652,N_5390,N_6020);
nand U8653 (N_8653,N_5970,N_4543);
nand U8654 (N_8654,N_7578,N_4104);
and U8655 (N_8655,N_7956,N_6714);
nand U8656 (N_8656,N_5343,N_7370);
nand U8657 (N_8657,N_7394,N_4258);
xor U8658 (N_8658,N_5037,N_6859);
nor U8659 (N_8659,N_5167,N_4683);
or U8660 (N_8660,N_4253,N_6547);
nand U8661 (N_8661,N_6605,N_5648);
and U8662 (N_8662,N_4922,N_6558);
or U8663 (N_8663,N_7928,N_5804);
nand U8664 (N_8664,N_5658,N_7492);
nor U8665 (N_8665,N_5573,N_7596);
and U8666 (N_8666,N_4488,N_5716);
and U8667 (N_8667,N_7375,N_6488);
and U8668 (N_8668,N_7579,N_6522);
xor U8669 (N_8669,N_7393,N_4391);
nor U8670 (N_8670,N_6755,N_6789);
xnor U8671 (N_8671,N_4162,N_6058);
nand U8672 (N_8672,N_7832,N_5277);
nand U8673 (N_8673,N_7110,N_4669);
nand U8674 (N_8674,N_7323,N_4243);
or U8675 (N_8675,N_6099,N_7065);
nand U8676 (N_8676,N_6001,N_4041);
nand U8677 (N_8677,N_6287,N_5260);
nor U8678 (N_8678,N_7850,N_5622);
nand U8679 (N_8679,N_4426,N_5969);
nor U8680 (N_8680,N_4518,N_4215);
nor U8681 (N_8681,N_6766,N_4311);
nand U8682 (N_8682,N_7244,N_7128);
or U8683 (N_8683,N_4554,N_4736);
or U8684 (N_8684,N_6926,N_7022);
and U8685 (N_8685,N_4367,N_7763);
and U8686 (N_8686,N_5990,N_4432);
nand U8687 (N_8687,N_4989,N_7911);
and U8688 (N_8688,N_7382,N_5961);
nand U8689 (N_8689,N_4847,N_4336);
nand U8690 (N_8690,N_7431,N_4176);
nand U8691 (N_8691,N_5476,N_5246);
and U8692 (N_8692,N_6729,N_6431);
and U8693 (N_8693,N_6492,N_4366);
or U8694 (N_8694,N_6725,N_4608);
or U8695 (N_8695,N_4674,N_5077);
xnor U8696 (N_8696,N_5290,N_4509);
nand U8697 (N_8697,N_5551,N_7265);
nand U8698 (N_8698,N_7894,N_4893);
xnor U8699 (N_8699,N_6963,N_6413);
nor U8700 (N_8700,N_4402,N_6526);
nand U8701 (N_8701,N_6047,N_5090);
nand U8702 (N_8702,N_5284,N_6528);
or U8703 (N_8703,N_4083,N_7893);
nor U8704 (N_8704,N_6867,N_5288);
nor U8705 (N_8705,N_4837,N_4733);
or U8706 (N_8706,N_6173,N_7528);
nand U8707 (N_8707,N_7534,N_5410);
nor U8708 (N_8708,N_4776,N_7149);
or U8709 (N_8709,N_5001,N_4156);
or U8710 (N_8710,N_7007,N_7148);
xor U8711 (N_8711,N_6861,N_5515);
and U8712 (N_8712,N_7650,N_4000);
xnor U8713 (N_8713,N_5162,N_4042);
nor U8714 (N_8714,N_4535,N_6440);
and U8715 (N_8715,N_7358,N_7341);
nand U8716 (N_8716,N_6510,N_4879);
nand U8717 (N_8717,N_5305,N_7120);
nor U8718 (N_8718,N_5354,N_6991);
or U8719 (N_8719,N_5876,N_6337);
and U8720 (N_8720,N_4267,N_5265);
or U8721 (N_8721,N_5004,N_4900);
nand U8722 (N_8722,N_6079,N_6806);
or U8723 (N_8723,N_5408,N_7313);
or U8724 (N_8724,N_4982,N_5418);
nand U8725 (N_8725,N_5689,N_7789);
or U8726 (N_8726,N_6807,N_5080);
and U8727 (N_8727,N_7571,N_7921);
nor U8728 (N_8728,N_4581,N_4114);
nand U8729 (N_8729,N_4529,N_4786);
xor U8730 (N_8730,N_5543,N_5663);
xor U8731 (N_8731,N_4620,N_4764);
and U8732 (N_8732,N_5191,N_6383);
nor U8733 (N_8733,N_4288,N_6694);
nor U8734 (N_8734,N_6005,N_4434);
nand U8735 (N_8735,N_7328,N_7290);
nor U8736 (N_8736,N_7047,N_5236);
nand U8737 (N_8737,N_4501,N_7884);
and U8738 (N_8738,N_4748,N_4579);
and U8739 (N_8739,N_7668,N_7337);
or U8740 (N_8740,N_7731,N_4514);
nand U8741 (N_8741,N_4838,N_4720);
and U8742 (N_8742,N_4710,N_5675);
or U8743 (N_8743,N_5659,N_5541);
or U8744 (N_8744,N_6728,N_7551);
and U8745 (N_8745,N_6305,N_6683);
nor U8746 (N_8746,N_7849,N_7865);
and U8747 (N_8747,N_4430,N_7138);
xor U8748 (N_8748,N_4090,N_5789);
xnor U8749 (N_8749,N_5577,N_4401);
or U8750 (N_8750,N_6411,N_4200);
xor U8751 (N_8751,N_7537,N_6422);
and U8752 (N_8752,N_5023,N_7796);
and U8753 (N_8753,N_4413,N_7388);
or U8754 (N_8754,N_4468,N_7556);
or U8755 (N_8755,N_6631,N_7795);
or U8756 (N_8756,N_6447,N_4714);
nor U8757 (N_8757,N_4833,N_7466);
nand U8758 (N_8758,N_6335,N_4101);
nand U8759 (N_8759,N_6936,N_7029);
nand U8760 (N_8760,N_6404,N_4328);
nor U8761 (N_8761,N_6460,N_6466);
and U8762 (N_8762,N_4017,N_6976);
and U8763 (N_8763,N_5020,N_4116);
nor U8764 (N_8764,N_6250,N_7819);
nor U8765 (N_8765,N_6995,N_7615);
xor U8766 (N_8766,N_6654,N_4111);
and U8767 (N_8767,N_5369,N_5341);
or U8768 (N_8768,N_7934,N_6113);
nand U8769 (N_8769,N_4677,N_6263);
nand U8770 (N_8770,N_7197,N_6829);
nor U8771 (N_8771,N_7359,N_7736);
nand U8772 (N_8772,N_6194,N_5660);
or U8773 (N_8773,N_6501,N_5862);
nand U8774 (N_8774,N_7106,N_5058);
nand U8775 (N_8775,N_6552,N_4047);
nor U8776 (N_8776,N_5921,N_7284);
nand U8777 (N_8777,N_5392,N_7291);
nand U8778 (N_8778,N_5519,N_7627);
nor U8779 (N_8779,N_4664,N_5192);
nand U8780 (N_8780,N_6349,N_7336);
nand U8781 (N_8781,N_4918,N_4046);
xnor U8782 (N_8782,N_4051,N_7916);
nand U8783 (N_8783,N_7448,N_4732);
and U8784 (N_8784,N_5927,N_5124);
and U8785 (N_8785,N_4363,N_6731);
nand U8786 (N_8786,N_7209,N_6217);
and U8787 (N_8787,N_4005,N_4242);
or U8788 (N_8788,N_4237,N_5189);
nand U8789 (N_8789,N_6110,N_4335);
and U8790 (N_8790,N_5135,N_6850);
xor U8791 (N_8791,N_6439,N_5204);
xnor U8792 (N_8792,N_4742,N_7277);
nand U8793 (N_8793,N_6149,N_6029);
xor U8794 (N_8794,N_6473,N_4386);
nand U8795 (N_8795,N_4279,N_4717);
and U8796 (N_8796,N_7144,N_4476);
or U8797 (N_8797,N_7652,N_5099);
and U8798 (N_8798,N_7859,N_7781);
and U8799 (N_8799,N_6324,N_5905);
nor U8800 (N_8800,N_6158,N_6559);
or U8801 (N_8801,N_7500,N_7246);
or U8802 (N_8802,N_4817,N_4159);
nand U8803 (N_8803,N_7964,N_7287);
and U8804 (N_8804,N_5028,N_4119);
and U8805 (N_8805,N_4410,N_7923);
and U8806 (N_8806,N_6842,N_5103);
nor U8807 (N_8807,N_5594,N_7829);
and U8808 (N_8808,N_7942,N_7721);
or U8809 (N_8809,N_6499,N_7851);
or U8810 (N_8810,N_4269,N_5666);
xnor U8811 (N_8811,N_5018,N_4823);
or U8812 (N_8812,N_5881,N_5151);
nor U8813 (N_8813,N_7460,N_4188);
or U8814 (N_8814,N_4172,N_5826);
and U8815 (N_8815,N_5973,N_4192);
nor U8816 (N_8816,N_4966,N_6457);
nor U8817 (N_8817,N_5249,N_6161);
nand U8818 (N_8818,N_7727,N_7631);
or U8819 (N_8819,N_4503,N_5736);
or U8820 (N_8820,N_5166,N_5051);
or U8821 (N_8821,N_5401,N_7519);
and U8822 (N_8822,N_7214,N_6222);
and U8823 (N_8823,N_4979,N_5344);
or U8824 (N_8824,N_7241,N_4896);
nor U8825 (N_8825,N_4891,N_7502);
or U8826 (N_8826,N_4358,N_7039);
xnor U8827 (N_8827,N_6232,N_4557);
nor U8828 (N_8828,N_7605,N_5164);
and U8829 (N_8829,N_6348,N_7476);
nor U8830 (N_8830,N_5345,N_5677);
nand U8831 (N_8831,N_5883,N_5740);
xnor U8832 (N_8832,N_4323,N_7708);
xor U8833 (N_8833,N_4547,N_6332);
nor U8834 (N_8834,N_4009,N_4513);
nand U8835 (N_8835,N_6266,N_5581);
and U8836 (N_8836,N_5384,N_6545);
or U8837 (N_8837,N_7154,N_5120);
and U8838 (N_8838,N_4143,N_5469);
or U8839 (N_8839,N_4250,N_6291);
or U8840 (N_8840,N_6661,N_7441);
nand U8841 (N_8841,N_5556,N_5317);
nor U8842 (N_8842,N_5672,N_4066);
and U8843 (N_8843,N_5109,N_4115);
nand U8844 (N_8844,N_7593,N_4486);
nor U8845 (N_8845,N_7953,N_7076);
or U8846 (N_8846,N_7845,N_4179);
nand U8847 (N_8847,N_7620,N_6539);
nand U8848 (N_8848,N_7094,N_7877);
nor U8849 (N_8849,N_6280,N_6835);
nand U8850 (N_8850,N_6784,N_5933);
and U8851 (N_8851,N_5446,N_7461);
nor U8852 (N_8852,N_6625,N_4964);
or U8853 (N_8853,N_5165,N_4065);
nor U8854 (N_8854,N_7153,N_6303);
nand U8855 (N_8855,N_4475,N_6136);
xnor U8856 (N_8856,N_7091,N_4859);
nor U8857 (N_8857,N_6872,N_5857);
xor U8858 (N_8858,N_7228,N_5214);
or U8859 (N_8859,N_5805,N_6560);
nand U8860 (N_8860,N_7573,N_7031);
nor U8861 (N_8861,N_4375,N_6415);
or U8862 (N_8862,N_4054,N_6520);
nor U8863 (N_8863,N_4024,N_6516);
nor U8864 (N_8864,N_7516,N_6653);
or U8865 (N_8865,N_5297,N_6347);
and U8866 (N_8866,N_5713,N_5104);
nor U8867 (N_8867,N_5145,N_6181);
or U8868 (N_8868,N_4092,N_6288);
nand U8869 (N_8869,N_6596,N_7828);
and U8870 (N_8870,N_6154,N_4429);
and U8871 (N_8871,N_7005,N_7137);
nor U8872 (N_8872,N_4489,N_5613);
nor U8873 (N_8873,N_4615,N_6027);
or U8874 (N_8874,N_7395,N_6938);
and U8875 (N_8875,N_5816,N_6593);
and U8876 (N_8876,N_4346,N_7641);
or U8877 (N_8877,N_5334,N_6863);
nor U8878 (N_8878,N_6182,N_4126);
and U8879 (N_8879,N_6371,N_5846);
nand U8880 (N_8880,N_7217,N_5770);
nand U8881 (N_8881,N_4174,N_4839);
or U8882 (N_8882,N_4578,N_5057);
or U8883 (N_8883,N_6022,N_4750);
nand U8884 (N_8884,N_6951,N_7434);
and U8885 (N_8885,N_7836,N_4136);
and U8886 (N_8886,N_5083,N_7844);
xnor U8887 (N_8887,N_4360,N_4721);
or U8888 (N_8888,N_6115,N_7948);
or U8889 (N_8889,N_4659,N_4377);
and U8890 (N_8890,N_5335,N_5807);
xor U8891 (N_8891,N_4146,N_4913);
and U8892 (N_8892,N_4070,N_7495);
nand U8893 (N_8893,N_6151,N_7206);
nand U8894 (N_8894,N_5858,N_7564);
and U8895 (N_8895,N_7536,N_4290);
nor U8896 (N_8896,N_7648,N_5416);
nand U8897 (N_8897,N_4840,N_7529);
nand U8898 (N_8898,N_7702,N_4628);
nand U8899 (N_8899,N_6875,N_7168);
and U8900 (N_8900,N_5470,N_4453);
nand U8901 (N_8901,N_7567,N_5703);
or U8902 (N_8902,N_5252,N_6325);
or U8903 (N_8903,N_7082,N_6908);
nand U8904 (N_8904,N_4161,N_6531);
or U8905 (N_8905,N_7123,N_7482);
xor U8906 (N_8906,N_7147,N_6229);
nand U8907 (N_8907,N_4313,N_5499);
and U8908 (N_8908,N_7223,N_5831);
and U8909 (N_8909,N_4866,N_5908);
nand U8910 (N_8910,N_4189,N_5910);
or U8911 (N_8911,N_7177,N_4238);
and U8912 (N_8912,N_7980,N_7133);
and U8913 (N_8913,N_5742,N_7059);
nand U8914 (N_8914,N_4021,N_5992);
and U8915 (N_8915,N_5084,N_7155);
and U8916 (N_8916,N_7459,N_6737);
xnor U8917 (N_8917,N_6647,N_7747);
nor U8918 (N_8918,N_7225,N_5953);
nand U8919 (N_8919,N_4609,N_6484);
xnor U8920 (N_8920,N_4731,N_4455);
nor U8921 (N_8921,N_6805,N_5634);
and U8922 (N_8922,N_5243,N_6933);
or U8923 (N_8923,N_4954,N_5199);
and U8924 (N_8924,N_6623,N_7842);
and U8925 (N_8925,N_6885,N_7665);
nand U8926 (N_8926,N_7959,N_4822);
and U8927 (N_8927,N_6014,N_5116);
nor U8928 (N_8928,N_6676,N_4870);
and U8929 (N_8929,N_7030,N_7281);
nand U8930 (N_8930,N_7771,N_6671);
nor U8931 (N_8931,N_6538,N_4369);
and U8932 (N_8932,N_7932,N_7994);
or U8933 (N_8933,N_4917,N_4381);
and U8934 (N_8934,N_7905,N_7438);
nand U8935 (N_8935,N_4291,N_5569);
xnor U8936 (N_8936,N_5682,N_4863);
nor U8937 (N_8937,N_5463,N_6208);
nand U8938 (N_8938,N_5330,N_4131);
nor U8939 (N_8939,N_7686,N_6167);
nor U8940 (N_8940,N_4061,N_5940);
nand U8941 (N_8941,N_7693,N_7966);
xnor U8942 (N_8942,N_5142,N_6677);
and U8943 (N_8943,N_6754,N_7093);
and U8944 (N_8944,N_4437,N_6666);
and U8945 (N_8945,N_7373,N_4743);
nor U8946 (N_8946,N_6175,N_7995);
and U8947 (N_8947,N_5632,N_4330);
and U8948 (N_8948,N_4819,N_7272);
xor U8949 (N_8949,N_7784,N_7124);
and U8950 (N_8950,N_7092,N_5975);
nor U8951 (N_8951,N_6911,N_5649);
or U8952 (N_8952,N_6489,N_6306);
or U8953 (N_8953,N_7588,N_6286);
nor U8954 (N_8954,N_6813,N_4461);
nand U8955 (N_8955,N_6310,N_5271);
nand U8956 (N_8956,N_5674,N_7288);
and U8957 (N_8957,N_7367,N_7507);
nand U8958 (N_8958,N_4148,N_4942);
or U8959 (N_8959,N_6432,N_6350);
or U8960 (N_8960,N_4790,N_5181);
nand U8961 (N_8961,N_7867,N_7423);
nand U8962 (N_8962,N_5838,N_6536);
and U8963 (N_8963,N_4592,N_4163);
and U8964 (N_8964,N_5406,N_5710);
or U8965 (N_8965,N_6220,N_6070);
or U8966 (N_8966,N_7360,N_7129);
or U8967 (N_8967,N_7212,N_5803);
xor U8968 (N_8968,N_6996,N_4849);
nand U8969 (N_8969,N_5436,N_7236);
and U8970 (N_8970,N_4011,N_4803);
nand U8971 (N_8971,N_5031,N_4851);
nor U8972 (N_8972,N_6852,N_4972);
or U8973 (N_8973,N_6680,N_6598);
or U8974 (N_8974,N_4613,N_5827);
xor U8975 (N_8975,N_5266,N_5424);
and U8976 (N_8976,N_4096,N_7897);
or U8977 (N_8977,N_6915,N_4758);
or U8978 (N_8978,N_6687,N_6673);
and U8979 (N_8979,N_4586,N_4976);
and U8980 (N_8980,N_7695,N_7425);
and U8981 (N_8981,N_4821,N_4076);
nand U8982 (N_8982,N_7369,N_4268);
nor U8983 (N_8983,N_5915,N_5695);
and U8984 (N_8984,N_7741,N_5107);
or U8985 (N_8985,N_7594,N_4852);
or U8986 (N_8986,N_5263,N_7526);
nand U8987 (N_8987,N_7365,N_5148);
nand U8988 (N_8988,N_4689,N_6758);
and U8989 (N_8989,N_5385,N_4285);
nor U8990 (N_8990,N_6089,N_6574);
and U8991 (N_8991,N_4325,N_4130);
and U8992 (N_8992,N_4540,N_4722);
xnor U8993 (N_8993,N_6689,N_6650);
and U8994 (N_8994,N_4801,N_5501);
or U8995 (N_8995,N_7525,N_4324);
nand U8996 (N_8996,N_5038,N_6540);
or U8997 (N_8997,N_6506,N_5245);
or U8998 (N_8998,N_7699,N_7755);
and U8999 (N_8999,N_6269,N_7351);
nor U9000 (N_9000,N_7550,N_5480);
or U9001 (N_9001,N_5533,N_5733);
nand U9002 (N_9002,N_4624,N_7462);
or U9003 (N_9003,N_6107,N_4167);
or U9004 (N_9004,N_6691,N_6544);
or U9005 (N_9005,N_4779,N_5067);
nor U9006 (N_9006,N_7203,N_4857);
or U9007 (N_9007,N_4641,N_6323);
and U9008 (N_9008,N_4629,N_4460);
nor U9009 (N_9009,N_5336,N_6660);
nand U9010 (N_9010,N_6090,N_7406);
or U9011 (N_9011,N_4692,N_5062);
nand U9012 (N_9012,N_6957,N_7439);
or U9013 (N_9013,N_6594,N_7777);
or U9014 (N_9014,N_6091,N_6478);
nand U9015 (N_9015,N_4120,N_6341);
or U9016 (N_9016,N_6203,N_6273);
xnor U9017 (N_9017,N_5417,N_7387);
and U9018 (N_9018,N_7167,N_5091);
nand U9019 (N_9019,N_7913,N_4409);
nand U9020 (N_9020,N_5591,N_5771);
or U9021 (N_9021,N_6087,N_4177);
or U9022 (N_9022,N_6733,N_4062);
and U9023 (N_9023,N_5866,N_4218);
or U9024 (N_9024,N_4504,N_4772);
nand U9025 (N_9025,N_6446,N_6602);
nor U9026 (N_9026,N_5375,N_4231);
nor U9027 (N_9027,N_5934,N_7613);
nand U9028 (N_9028,N_5932,N_5007);
nand U9029 (N_9029,N_6223,N_6865);
or U9030 (N_9030,N_7612,N_6245);
nand U9031 (N_9031,N_5478,N_6120);
nand U9032 (N_9032,N_5136,N_7498);
nand U9033 (N_9033,N_5194,N_4806);
nand U9034 (N_9034,N_7239,N_5753);
and U9035 (N_9035,N_5544,N_7490);
or U9036 (N_9036,N_6387,N_6781);
and U9037 (N_9037,N_7264,N_7200);
xor U9038 (N_9038,N_5609,N_7754);
or U9039 (N_9039,N_5068,N_6801);
and U9040 (N_9040,N_5698,N_4353);
nor U9041 (N_9041,N_5179,N_6344);
nor U9042 (N_9042,N_7067,N_7509);
nor U9043 (N_9043,N_4796,N_4454);
and U9044 (N_9044,N_4373,N_4778);
nor U9045 (N_9045,N_6160,N_7547);
and U9046 (N_9046,N_7812,N_7226);
and U9047 (N_9047,N_4614,N_4561);
or U9048 (N_9048,N_4517,N_7883);
and U9049 (N_9049,N_7786,N_6331);
xnor U9050 (N_9050,N_5178,N_5683);
nand U9051 (N_9051,N_7868,N_7136);
nand U9052 (N_9052,N_4715,N_4607);
and U9053 (N_9053,N_6297,N_5066);
or U9054 (N_9054,N_7734,N_7924);
or U9055 (N_9055,N_7324,N_5856);
or U9056 (N_9056,N_5853,N_4077);
xnor U9057 (N_9057,N_7726,N_6645);
or U9058 (N_9058,N_6094,N_7174);
and U9059 (N_9059,N_5655,N_4915);
nor U9060 (N_9060,N_6709,N_7907);
nor U9061 (N_9061,N_5610,N_5286);
xnor U9062 (N_9062,N_6803,N_6436);
nor U9063 (N_9063,N_5359,N_5690);
nor U9064 (N_9064,N_6448,N_7640);
and U9065 (N_9065,N_6656,N_7552);
and U9066 (N_9066,N_6970,N_7285);
and U9067 (N_9067,N_7632,N_5017);
and U9068 (N_9068,N_6360,N_6421);
and U9069 (N_9069,N_4102,N_4462);
nand U9070 (N_9070,N_4832,N_7619);
nor U9071 (N_9071,N_4029,N_6809);
nor U9072 (N_9072,N_4770,N_4004);
nor U9073 (N_9073,N_5137,N_4573);
nand U9074 (N_9074,N_6028,N_6541);
nor U9075 (N_9075,N_7558,N_4745);
nand U9076 (N_9076,N_4019,N_6221);
nor U9077 (N_9077,N_6103,N_6696);
xnor U9078 (N_9078,N_7930,N_6380);
or U9079 (N_9079,N_5828,N_5451);
and U9080 (N_9080,N_5398,N_5299);
nand U9081 (N_9081,N_7716,N_5879);
or U9082 (N_9082,N_4050,N_4985);
and U9083 (N_9083,N_4220,N_7949);
nand U9084 (N_9084,N_4201,N_7876);
or U9085 (N_9085,N_6183,N_5629);
xor U9086 (N_9086,N_4661,N_7630);
nor U9087 (N_9087,N_5603,N_6899);
nor U9088 (N_9088,N_6427,N_4443);
nand U9089 (N_9089,N_6211,N_5692);
nand U9090 (N_9090,N_6727,N_7151);
nand U9091 (N_9091,N_6000,N_6056);
and U9092 (N_9092,N_5487,N_5516);
and U9093 (N_9093,N_5060,N_7072);
nand U9094 (N_9094,N_5036,N_5251);
xnor U9095 (N_9095,N_4436,N_7957);
nand U9096 (N_9096,N_5549,N_6848);
or U9097 (N_9097,N_5029,N_4599);
xnor U9098 (N_9098,N_6982,N_7794);
or U9099 (N_9099,N_6271,N_5276);
and U9100 (N_9100,N_5537,N_6584);
nand U9101 (N_9101,N_6892,N_4835);
nor U9102 (N_9102,N_7804,N_7635);
or U9103 (N_9103,N_6975,N_5825);
or U9104 (N_9104,N_5319,N_4433);
xor U9105 (N_9105,N_7752,N_5097);
xor U9106 (N_9106,N_6870,N_7724);
xor U9107 (N_9107,N_6057,N_5044);
or U9108 (N_9108,N_4903,N_4598);
xor U9109 (N_9109,N_6238,N_6716);
and U9110 (N_9110,N_7404,N_7464);
nor U9111 (N_9111,N_6849,N_4214);
or U9112 (N_9112,N_7456,N_4684);
or U9113 (N_9113,N_5554,N_7170);
nand U9114 (N_9114,N_6585,N_5859);
and U9115 (N_9115,N_6950,N_7435);
nand U9116 (N_9116,N_5279,N_4364);
or U9117 (N_9117,N_4927,N_5745);
nor U9118 (N_9118,N_4724,N_4016);
nor U9119 (N_9119,N_5784,N_7676);
nor U9120 (N_9120,N_5638,N_6073);
xnor U9121 (N_9121,N_5950,N_6988);
and U9122 (N_9122,N_5332,N_4355);
and U9123 (N_9123,N_5747,N_6998);
xnor U9124 (N_9124,N_5054,N_7827);
or U9125 (N_9125,N_5851,N_4795);
and U9126 (N_9126,N_5725,N_4804);
and U9127 (N_9127,N_6565,N_7712);
or U9128 (N_9128,N_6613,N_5842);
or U9129 (N_9129,N_6356,N_7354);
and U9130 (N_9130,N_4802,N_5546);
and U9131 (N_9131,N_4729,N_5836);
nand U9132 (N_9132,N_4178,N_5723);
nor U9133 (N_9133,N_6319,N_5714);
and U9134 (N_9134,N_4612,N_6967);
nand U9135 (N_9135,N_7606,N_6017);
and U9136 (N_9136,N_6215,N_6741);
or U9137 (N_9137,N_4812,N_6268);
and U9138 (N_9138,N_6367,N_5175);
nand U9139 (N_9139,N_7115,N_4564);
nor U9140 (N_9140,N_6615,N_7207);
or U9141 (N_9141,N_4007,N_5298);
xor U9142 (N_9142,N_5865,N_4327);
nor U9143 (N_9143,N_7802,N_7426);
nand U9144 (N_9144,N_7811,N_7353);
and U9145 (N_9145,N_6464,N_5397);
and U9146 (N_9146,N_6456,N_4068);
nand U9147 (N_9147,N_4448,N_5082);
and U9148 (N_9148,N_5777,N_4572);
xnor U9149 (N_9149,N_7243,N_5309);
nor U9150 (N_9150,N_4756,N_4531);
nor U9151 (N_9151,N_6338,N_7463);
nand U9152 (N_9152,N_4305,N_4625);
xor U9153 (N_9153,N_4271,N_6105);
or U9154 (N_9154,N_7164,N_6794);
and U9155 (N_9155,N_5200,N_4771);
nor U9156 (N_9156,N_6514,N_4474);
or U9157 (N_9157,N_4582,N_4107);
and U9158 (N_9158,N_7638,N_4761);
nor U9159 (N_9159,N_7499,N_4970);
and U9160 (N_9160,N_4309,N_4508);
or U9161 (N_9161,N_4800,N_5219);
nor U9162 (N_9162,N_6036,N_4154);
nor U9163 (N_9163,N_7042,N_4217);
nor U9164 (N_9164,N_4744,N_4209);
or U9165 (N_9165,N_4283,N_6481);
nor U9166 (N_9166,N_4128,N_7798);
or U9167 (N_9167,N_6059,N_7510);
and U9168 (N_9168,N_4816,N_5768);
or U9169 (N_9169,N_4713,N_5599);
and U9170 (N_9170,N_7886,N_6990);
nor U9171 (N_9171,N_7109,N_7349);
or U9172 (N_9172,N_6609,N_7750);
and U9173 (N_9173,N_6712,N_4097);
nand U9174 (N_9174,N_7019,N_4568);
nor U9175 (N_9175,N_4785,N_5661);
and U9176 (N_9176,N_5221,N_5395);
nand U9177 (N_9177,N_6641,N_5156);
nand U9178 (N_9178,N_7472,N_7575);
nand U9179 (N_9179,N_7166,N_7355);
or U9180 (N_9180,N_7189,N_6576);
nand U9181 (N_9181,N_5318,N_7117);
xor U9182 (N_9182,N_4878,N_5182);
or U9183 (N_9183,N_7386,N_7970);
nand U9184 (N_9184,N_6668,N_4780);
nor U9185 (N_9185,N_5110,N_5402);
nor U9186 (N_9186,N_7936,N_4297);
and U9187 (N_9187,N_7024,N_4112);
and U9188 (N_9188,N_6088,N_4278);
and U9189 (N_9189,N_4060,N_6599);
or U9190 (N_9190,N_4571,N_6033);
and U9191 (N_9191,N_6486,N_5588);
or U9192 (N_9192,N_7670,N_7469);
nor U9193 (N_9193,N_6104,N_4944);
nand U9194 (N_9194,N_4145,N_7156);
xor U9195 (N_9195,N_7494,N_5746);
nor U9196 (N_9196,N_4654,N_7539);
and U9197 (N_9197,N_4960,N_6877);
nand U9198 (N_9198,N_6577,N_6897);
nand U9199 (N_9199,N_4662,N_7945);
nand U9200 (N_9200,N_6042,N_5835);
and U9201 (N_9201,N_5208,N_7062);
nor U9202 (N_9202,N_7733,N_4910);
and U9203 (N_9203,N_7800,N_7696);
nand U9204 (N_9204,N_5693,N_4098);
nor U9205 (N_9205,N_4993,N_5443);
nor U9206 (N_9206,N_6247,N_5783);
or U9207 (N_9207,N_6365,N_6239);
nand U9208 (N_9208,N_7576,N_6201);
xor U9209 (N_9209,N_7532,N_7527);
and U9210 (N_9210,N_6498,N_5430);
and U9211 (N_9211,N_7618,N_6171);
or U9212 (N_9212,N_5982,N_7687);
xor U9213 (N_9213,N_6675,N_7915);
nor U9214 (N_9214,N_7910,N_6398);
nand U9215 (N_9215,N_7860,N_5414);
nor U9216 (N_9216,N_4961,N_6948);
nor U9217 (N_9217,N_6760,N_7491);
nand U9218 (N_9218,N_6826,N_7872);
and U9219 (N_9219,N_4551,N_6797);
nand U9220 (N_9220,N_4093,N_7599);
or U9221 (N_9221,N_5815,N_4479);
and U9222 (N_9222,N_6254,N_5140);
and U9223 (N_9223,N_5583,N_6701);
xor U9224 (N_9224,N_5064,N_6068);
nor U9225 (N_9225,N_7107,N_6854);
or U9226 (N_9226,N_7825,N_4844);
or U9227 (N_9227,N_5159,N_4794);
nand U9228 (N_9228,N_4149,N_5331);
or U9229 (N_9229,N_4818,N_7658);
nor U9230 (N_9230,N_5759,N_7968);
nand U9231 (N_9231,N_5653,N_7938);
nand U9232 (N_9232,N_5640,N_6189);
nor U9233 (N_9233,N_5679,N_5412);
nor U9234 (N_9234,N_4320,N_4735);
nand U9235 (N_9235,N_5943,N_6883);
nor U9236 (N_9236,N_5096,N_5995);
or U9237 (N_9237,N_4265,N_5198);
or U9238 (N_9238,N_6804,N_7909);
nand U9239 (N_9239,N_7955,N_6889);
and U9240 (N_9240,N_6438,N_6554);
and U9241 (N_9241,N_4071,N_6180);
nand U9242 (N_9242,N_6535,N_6874);
and U9243 (N_9243,N_5935,N_6329);
nor U9244 (N_9244,N_5671,N_6959);
or U9245 (N_9245,N_7152,N_5323);
nand U9246 (N_9246,N_5895,N_5620);
and U9247 (N_9247,N_5425,N_4185);
nor U9248 (N_9248,N_4505,N_7477);
nor U9249 (N_9249,N_4308,N_7259);
and U9250 (N_9250,N_4399,N_5355);
or U9251 (N_9251,N_4260,N_7306);
nand U9252 (N_9252,N_7983,N_4251);
nor U9253 (N_9253,N_4484,N_6458);
nor U9254 (N_9254,N_6721,N_6674);
and U9255 (N_9255,N_4740,N_6815);
nor U9256 (N_9256,N_5721,N_7584);
nor U9257 (N_9257,N_4558,N_5994);
xnor U9258 (N_9258,N_5694,N_4532);
and U9259 (N_9259,N_7678,N_4824);
nand U9260 (N_9260,N_4495,N_5367);
and U9261 (N_9261,N_4210,N_7611);
and U9262 (N_9262,N_7935,N_6032);
nand U9263 (N_9263,N_4206,N_6462);
and U9264 (N_9264,N_7939,N_7266);
and U9265 (N_9265,N_5680,N_6630);
xnor U9266 (N_9266,N_7833,N_6253);
nor U9267 (N_9267,N_5545,N_4001);
or U9268 (N_9268,N_4032,N_5468);
and U9269 (N_9269,N_7698,N_4186);
or U9270 (N_9270,N_5642,N_5070);
xor U9271 (N_9271,N_7600,N_6816);
and U9272 (N_9272,N_4463,N_5160);
or U9273 (N_9273,N_6174,N_5088);
nor U9274 (N_9274,N_6216,N_5427);
nor U9275 (N_9275,N_6604,N_4673);
or U9276 (N_9276,N_7400,N_6834);
and U9277 (N_9277,N_5006,N_6003);
or U9278 (N_9278,N_7270,N_4431);
nor U9279 (N_9279,N_6363,N_5042);
nor U9280 (N_9280,N_4227,N_7252);
xnor U9281 (N_9281,N_6320,N_6943);
xnor U9282 (N_9282,N_7496,N_7742);
nor U9283 (N_9283,N_5421,N_4326);
or U9284 (N_9284,N_5144,N_4862);
or U9285 (N_9285,N_4696,N_7086);
nor U9286 (N_9286,N_7729,N_4658);
nand U9287 (N_9287,N_4858,N_4385);
and U9288 (N_9288,N_4655,N_7793);
or U9289 (N_9289,N_7749,N_6768);
nand U9290 (N_9290,N_6608,N_6524);
nor U9291 (N_9291,N_5346,N_6614);
and U9292 (N_9292,N_4881,N_7661);
and U9293 (N_9293,N_6343,N_6788);
nor U9294 (N_9294,N_6474,N_7326);
xor U9295 (N_9295,N_5606,N_7972);
and U9296 (N_9296,N_5818,N_5652);
or U9297 (N_9297,N_7992,N_7204);
and U9298 (N_9298,N_4318,N_7308);
nand U9299 (N_9299,N_4383,N_6983);
xnor U9300 (N_9300,N_5394,N_5324);
nor U9301 (N_9301,N_5700,N_6326);
nor U9302 (N_9302,N_4938,N_6764);
or U9303 (N_9303,N_6495,N_7870);
nor U9304 (N_9304,N_7034,N_4350);
or U9305 (N_9305,N_7300,N_7098);
or U9306 (N_9306,N_5389,N_7060);
and U9307 (N_9307,N_4685,N_4604);
nand U9308 (N_9308,N_5665,N_6454);
nor U9309 (N_9309,N_7058,N_4226);
nor U9310 (N_9310,N_5289,N_6192);
and U9311 (N_9311,N_7511,N_6679);
nor U9312 (N_9312,N_6121,N_5938);
or U9313 (N_9313,N_7157,N_6143);
xor U9314 (N_9314,N_7269,N_5860);
and U9315 (N_9315,N_5292,N_5762);
nand U9316 (N_9316,N_4403,N_4414);
or U9317 (N_9317,N_7673,N_4949);
xnor U9318 (N_9318,N_6135,N_6776);
nor U9319 (N_9319,N_6986,N_4810);
nor U9320 (N_9320,N_5273,N_5218);
nor U9321 (N_9321,N_7783,N_5882);
and U9322 (N_9322,N_5411,N_5143);
nand U9323 (N_9323,N_6409,N_6588);
xor U9324 (N_9324,N_4593,N_5381);
or U9325 (N_9325,N_6430,N_7025);
nor U9326 (N_9326,N_7577,N_4808);
or U9327 (N_9327,N_4388,N_5833);
and U9328 (N_9328,N_5971,N_4459);
and U9329 (N_9329,N_5201,N_4987);
xnor U9330 (N_9330,N_4580,N_6649);
xnor U9331 (N_9331,N_6913,N_5005);
nor U9332 (N_9332,N_5667,N_7993);
or U9333 (N_9333,N_6693,N_4170);
nor U9334 (N_9334,N_5184,N_7283);
or U9335 (N_9335,N_6219,N_6130);
nor U9336 (N_9336,N_4760,N_4644);
xnor U9337 (N_9337,N_7213,N_6111);
nor U9338 (N_9338,N_6055,N_4347);
or U9339 (N_9339,N_5073,N_5643);
and U9340 (N_9340,N_5485,N_4257);
xor U9341 (N_9341,N_7002,N_4765);
nand U9342 (N_9342,N_5651,N_5428);
or U9343 (N_9343,N_7756,N_5248);
or U9344 (N_9344,N_5707,N_4345);
nand U9345 (N_9345,N_5743,N_5459);
and U9346 (N_9346,N_5926,N_4447);
nand U9347 (N_9347,N_7077,N_4133);
nor U9348 (N_9348,N_7001,N_5739);
or U9349 (N_9349,N_6672,N_4908);
nand U9350 (N_9350,N_5702,N_7481);
or U9351 (N_9351,N_4521,N_6551);
nand U9352 (N_9352,N_5000,N_5374);
and U9353 (N_9353,N_4591,N_4700);
or U9354 (N_9354,N_7182,N_4548);
and U9355 (N_9355,N_6295,N_7216);
and U9356 (N_9356,N_5993,N_7397);
or U9357 (N_9357,N_4559,N_7111);
xnor U9358 (N_9358,N_4438,N_6589);
nand U9359 (N_9359,N_5456,N_4138);
or U9360 (N_9360,N_5176,N_7196);
nor U9361 (N_9361,N_6786,N_5823);
and U9362 (N_9362,N_7647,N_4035);
xor U9363 (N_9363,N_6900,N_7422);
or U9364 (N_9364,N_7303,N_5902);
and U9365 (N_9365,N_7140,N_6309);
nand U9366 (N_9366,N_7436,N_4727);
xnor U9367 (N_9367,N_5553,N_6597);
nor U9368 (N_9368,N_4233,N_6898);
nor U9369 (N_9369,N_6706,N_7874);
or U9370 (N_9370,N_4252,N_4678);
xnor U9371 (N_9371,N_4184,N_7339);
and U9372 (N_9372,N_5253,N_6159);
nand U9373 (N_9373,N_5069,N_4583);
nand U9374 (N_9374,N_6184,N_5466);
xnor U9375 (N_9375,N_4647,N_6276);
nor U9376 (N_9376,N_5039,N_5089);
nor U9377 (N_9377,N_4726,N_5576);
nor U9378 (N_9378,N_5602,N_4869);
or U9379 (N_9379,N_7286,N_5522);
and U9380 (N_9380,N_7981,N_5999);
or U9381 (N_9381,N_4404,N_5763);
xor U9382 (N_9382,N_7642,N_5542);
xnor U9383 (N_9383,N_6376,N_5117);
nor U9384 (N_9384,N_4415,N_7522);
and U9385 (N_9385,N_4408,N_7546);
or U9386 (N_9386,N_6634,N_4422);
nor U9387 (N_9387,N_6450,N_5877);
xnor U9388 (N_9388,N_5761,N_5906);
nand U9389 (N_9389,N_7743,N_5361);
nand U9390 (N_9390,N_4757,N_5386);
nand U9391 (N_9391,N_7586,N_5491);
or U9392 (N_9392,N_6483,N_5508);
nor U9393 (N_9393,N_4956,N_4322);
and U9394 (N_9394,N_5691,N_5405);
or U9395 (N_9395,N_6635,N_5383);
nor U9396 (N_9396,N_7580,N_4575);
nor U9397 (N_9397,N_6270,N_5131);
or U9398 (N_9398,N_7700,N_5565);
and U9399 (N_9399,N_7340,N_6556);
and U9400 (N_9400,N_5291,N_6517);
nor U9401 (N_9401,N_7100,N_5027);
and U9402 (N_9402,N_6424,N_5372);
nor U9403 (N_9403,N_5413,N_4282);
nor U9404 (N_9404,N_5278,N_4074);
and U9405 (N_9405,N_4491,N_6008);
nor U9406 (N_9406,N_4303,N_5061);
xor U9407 (N_9407,N_6999,N_4127);
nor U9408 (N_9408,N_5564,N_6093);
nor U9409 (N_9409,N_6246,N_7626);
or U9410 (N_9410,N_5872,N_5628);
nand U9411 (N_9411,N_6710,N_4370);
nor U9412 (N_9412,N_5210,N_7127);
nor U9413 (N_9413,N_6873,N_7814);
nand U9414 (N_9414,N_4056,N_4515);
or U9415 (N_9415,N_4670,N_6230);
nand U9416 (N_9416,N_7419,N_4239);
nand U9417 (N_9417,N_7338,N_6264);
xor U9418 (N_9418,N_5981,N_6251);
and U9419 (N_9419,N_7014,N_5668);
or U9420 (N_9420,N_5161,N_6002);
and U9421 (N_9421,N_6045,N_7654);
xnor U9422 (N_9422,N_7785,N_6030);
and U9423 (N_9423,N_6141,N_7680);
and U9424 (N_9424,N_4106,N_4080);
or U9425 (N_9425,N_6555,N_7344);
and U9426 (N_9426,N_5447,N_5259);
or U9427 (N_9427,N_4300,N_5370);
and U9428 (N_9428,N_7882,N_7520);
or U9429 (N_9429,N_5869,N_7738);
nor U9430 (N_9430,N_7103,N_6408);
nand U9431 (N_9431,N_4920,N_5347);
nand U9432 (N_9432,N_7875,N_5269);
or U9433 (N_9433,N_6525,N_5772);
or U9434 (N_9434,N_4998,N_6134);
and U9435 (N_9435,N_5837,N_4973);
nand U9436 (N_9436,N_5850,N_7683);
and U9437 (N_9437,N_5230,N_7890);
nand U9438 (N_9438,N_4063,N_7255);
or U9439 (N_9439,N_5808,N_5295);
nand U9440 (N_9440,N_5618,N_7864);
or U9441 (N_9441,N_7125,N_4371);
xnor U9442 (N_9442,N_5582,N_4424);
nor U9443 (N_9443,N_7769,N_5049);
nand U9444 (N_9444,N_7889,N_7518);
nor U9445 (N_9445,N_5814,N_5320);
and U9446 (N_9446,N_7247,N_4234);
and U9447 (N_9447,N_4924,N_7639);
nand U9448 (N_9448,N_7746,N_4939);
nor U9449 (N_9449,N_6905,N_5441);
and U9450 (N_9450,N_5810,N_5507);
nor U9451 (N_9451,N_4219,N_5952);
or U9452 (N_9452,N_6471,N_4173);
and U9453 (N_9453,N_6844,N_7704);
nand U9454 (N_9454,N_5949,N_6648);
nor U9455 (N_9455,N_5063,N_7660);
or U9456 (N_9456,N_6080,N_5720);
and U9457 (N_9457,N_6955,N_6334);
nor U9458 (N_9458,N_4660,N_5329);
or U9459 (N_9459,N_4261,N_6249);
nor U9460 (N_9460,N_7446,N_7116);
nand U9461 (N_9461,N_4199,N_6401);
nand U9462 (N_9462,N_7901,N_7317);
xor U9463 (N_9463,N_5013,N_6480);
nor U9464 (N_9464,N_5353,N_7245);
and U9465 (N_9465,N_5307,N_6101);
and U9466 (N_9466,N_7776,N_7135);
nor U9467 (N_9467,N_5986,N_6302);
and U9468 (N_9468,N_4395,N_6884);
xor U9469 (N_9469,N_5909,N_4923);
nor U9470 (N_9470,N_5426,N_7242);
and U9471 (N_9471,N_5147,N_4855);
or U9472 (N_9472,N_4829,N_7032);
nor U9473 (N_9473,N_7592,N_6147);
xnor U9474 (N_9474,N_7780,N_7852);
nand U9475 (N_9475,N_7912,N_4048);
and U9476 (N_9476,N_6543,N_5781);
nor U9477 (N_9477,N_7834,N_6523);
xnor U9478 (N_9478,N_5113,N_7409);
xnor U9479 (N_9479,N_7335,N_5566);
or U9480 (N_9480,N_4842,N_4981);
xor U9481 (N_9481,N_5912,N_5155);
nand U9482 (N_9482,N_5517,N_7506);
nand U9483 (N_9483,N_6385,N_6612);
or U9484 (N_9484,N_7195,N_4142);
nand U9485 (N_9485,N_7475,N_6697);
nand U9486 (N_9486,N_7643,N_4746);
nor U9487 (N_9487,N_4450,N_6108);
nor U9488 (N_9488,N_4889,N_4552);
nand U9489 (N_9489,N_6947,N_7768);
nand U9490 (N_9490,N_5847,N_6129);
or U9491 (N_9491,N_6508,N_6083);
nor U9492 (N_9492,N_5102,N_6074);
nor U9493 (N_9493,N_5280,N_4284);
nor U9494 (N_9494,N_5939,N_4223);
nor U9495 (N_9495,N_4526,N_4418);
nor U9496 (N_9496,N_4183,N_5275);
and U9497 (N_9497,N_5378,N_7512);
or U9498 (N_9498,N_4249,N_7562);
and U9499 (N_9499,N_7958,N_4105);
nor U9500 (N_9500,N_7888,N_4820);
nor U9501 (N_9501,N_5086,N_6922);
nand U9502 (N_9502,N_6352,N_4541);
xnor U9503 (N_9503,N_5315,N_7057);
nor U9504 (N_9504,N_4904,N_7753);
nand U9505 (N_9505,N_6586,N_4153);
nand U9506 (N_9506,N_7566,N_4787);
nand U9507 (N_9507,N_5955,N_4836);
nor U9508 (N_9508,N_6169,N_6467);
nor U9509 (N_9509,N_4865,N_5034);
and U9510 (N_9510,N_4277,N_7316);
or U9511 (N_9511,N_4968,N_6606);
nor U9512 (N_9512,N_6592,N_6299);
or U9513 (N_9513,N_6226,N_5788);
and U9514 (N_9514,N_4338,N_6664);
nor U9515 (N_9515,N_5126,N_6895);
nor U9516 (N_9516,N_5026,N_6451);
and U9517 (N_9517,N_7744,N_6434);
nor U9518 (N_9518,N_6954,N_6100);
nand U9519 (N_9519,N_7256,N_5016);
xnor U9520 (N_9520,N_4387,N_6054);
nor U9521 (N_9521,N_5321,N_5645);
nor U9522 (N_9522,N_4657,N_6403);
nor U9523 (N_9523,N_7010,N_6743);
or U9524 (N_9524,N_7568,N_6770);
nand U9525 (N_9525,N_4125,N_6049);
nor U9526 (N_9526,N_7319,N_6066);
nand U9527 (N_9527,N_4959,N_4897);
and U9528 (N_9528,N_4222,N_5078);
nand U9529 (N_9529,N_4493,N_4538);
nor U9530 (N_9530,N_6041,N_7470);
xor U9531 (N_9531,N_5664,N_4478);
nor U9532 (N_9532,N_5433,N_6065);
xor U9533 (N_9533,N_5186,N_5748);
or U9534 (N_9534,N_5893,N_5531);
and U9535 (N_9535,N_6084,N_5612);
or U9536 (N_9536,N_6969,N_7035);
or U9537 (N_9537,N_4895,N_4464);
nand U9538 (N_9538,N_6749,N_7131);
or U9539 (N_9539,N_4020,N_7454);
nor U9540 (N_9540,N_7717,N_6435);
nor U9541 (N_9541,N_5180,N_4882);
nand U9542 (N_9542,N_5584,N_7041);
and U9543 (N_9543,N_4467,N_7263);
and U9544 (N_9544,N_4033,N_6509);
xor U9545 (N_9545,N_6929,N_4510);
xnor U9546 (N_9546,N_4975,N_7322);
and U9547 (N_9547,N_6127,N_5717);
or U9548 (N_9548,N_5574,N_5907);
or U9549 (N_9549,N_7099,N_5360);
or U9550 (N_9550,N_7309,N_7333);
and U9551 (N_9551,N_7033,N_7563);
nand U9552 (N_9552,N_6123,N_7327);
xor U9553 (N_9553,N_7637,N_5237);
and U9554 (N_9554,N_6150,N_6956);
or U9555 (N_9555,N_7484,N_7549);
or U9556 (N_9556,N_6519,N_6259);
nor U9557 (N_9557,N_6916,N_5255);
or U9558 (N_9558,N_4627,N_4996);
nand U9559 (N_9559,N_7056,N_5578);
nand U9560 (N_9560,N_6482,N_6392);
nor U9561 (N_9561,N_7361,N_5754);
and U9562 (N_9562,N_5484,N_4180);
nor U9563 (N_9563,N_7774,N_4502);
and U9564 (N_9564,N_7817,N_7906);
nor U9565 (N_9565,N_5888,N_7572);
or U9566 (N_9566,N_7645,N_4867);
nand U9567 (N_9567,N_7818,N_7950);
or U9568 (N_9568,N_4762,N_6681);
nand U9569 (N_9569,N_5220,N_6636);
or U9570 (N_9570,N_6769,N_5976);
nand U9571 (N_9571,N_4723,N_6843);
or U9572 (N_9572,N_5092,N_6316);
nor U9573 (N_9573,N_5183,N_4983);
nand U9574 (N_9574,N_5228,N_6824);
xnor U9575 (N_9575,N_4828,N_4588);
and U9576 (N_9576,N_5997,N_4914);
or U9577 (N_9577,N_6704,N_5527);
and U9578 (N_9578,N_6902,N_4799);
nor U9579 (N_9579,N_5316,N_7020);
nor U9580 (N_9580,N_7730,N_6490);
nor U9581 (N_9581,N_4860,N_7267);
and U9582 (N_9582,N_5366,N_7071);
and U9583 (N_9583,N_5821,N_5012);
nor U9584 (N_9584,N_5489,N_4988);
nor U9585 (N_9585,N_5387,N_7975);
and U9586 (N_9586,N_5471,N_6081);
nor U9587 (N_9587,N_5513,N_7684);
and U9588 (N_9588,N_4202,N_4945);
nand U9589 (N_9589,N_6364,N_6155);
nor U9590 (N_9590,N_5376,N_7145);
or U9591 (N_9591,N_7449,N_5238);
or U9592 (N_9592,N_6864,N_4701);
nor U9593 (N_9593,N_7544,N_6997);
xor U9594 (N_9594,N_4109,N_6426);
or U9595 (N_9595,N_6372,N_4618);
or U9596 (N_9596,N_4304,N_5592);
and U9597 (N_9597,N_4045,N_4203);
nand U9598 (N_9598,N_5196,N_6752);
nor U9599 (N_9599,N_6921,N_6629);
nor U9600 (N_9600,N_6425,N_6910);
nand U9601 (N_9601,N_7984,N_4537);
xnor U9602 (N_9602,N_7855,N_4466);
and U9603 (N_9603,N_6012,N_5670);
nor U9604 (N_9604,N_4754,N_4676);
nor U9605 (N_9605,N_6530,N_4925);
nor U9606 (N_9606,N_4084,N_6962);
nand U9607 (N_9607,N_5460,N_5333);
nand U9608 (N_9608,N_4621,N_6652);
and U9609 (N_9609,N_4549,N_6684);
or U9610 (N_9610,N_7118,N_6078);
and U9611 (N_9611,N_5396,N_7691);
nor U9612 (N_9612,N_7061,N_4166);
and U9613 (N_9613,N_4675,N_6942);
nand U9614 (N_9614,N_7806,N_4270);
nand U9615 (N_9615,N_5076,N_4932);
xor U9616 (N_9616,N_5356,N_4295);
and U9617 (N_9617,N_6301,N_5654);
nand U9618 (N_9618,N_6117,N_7735);
and U9619 (N_9619,N_4622,N_4876);
xor U9620 (N_9620,N_4058,N_6023);
nor U9621 (N_9621,N_7999,N_5600);
nand U9622 (N_9622,N_7656,N_6564);
xnor U9623 (N_9623,N_7273,N_4793);
nand U9624 (N_9624,N_6116,N_4002);
and U9625 (N_9625,N_5709,N_4317);
nor U9626 (N_9626,N_5829,N_7479);
nor U9627 (N_9627,N_6354,N_5270);
and U9628 (N_9628,N_4419,N_6131);
nor U9629 (N_9629,N_7199,N_5959);
nand U9630 (N_9630,N_7310,N_7649);
and U9631 (N_9631,N_5525,N_5963);
nor U9632 (N_9632,N_4396,N_4730);
and U9633 (N_9633,N_6624,N_7048);
or U9634 (N_9634,N_7018,N_7574);
nor U9635 (N_9635,N_6578,N_4560);
and U9636 (N_9636,N_7384,N_5171);
nand U9637 (N_9637,N_7260,N_5792);
and U9638 (N_9638,N_5357,N_7514);
or U9639 (N_9639,N_7363,N_4805);
and U9640 (N_9640,N_6987,N_7473);
and U9641 (N_9641,N_4854,N_5462);
xnor U9642 (N_9642,N_6793,N_4122);
or U9643 (N_9643,N_6791,N_5207);
and U9644 (N_9644,N_4194,N_5047);
nand U9645 (N_9645,N_6468,N_7208);
and U9646 (N_9646,N_6812,N_5729);
and U9647 (N_9647,N_6395,N_7381);
or U9648 (N_9648,N_5407,N_5445);
and U9649 (N_9649,N_7672,N_6164);
nor U9650 (N_9650,N_5776,N_7257);
nor U9651 (N_9651,N_7778,N_5254);
nor U9652 (N_9652,N_7629,N_5884);
or U9653 (N_9653,N_4458,N_5503);
nand U9654 (N_9654,N_7037,N_7791);
and U9655 (N_9655,N_5945,N_5529);
or U9656 (N_9656,N_6685,N_5002);
nand U9657 (N_9657,N_5520,N_5209);
nor U9658 (N_9658,N_7863,N_5611);
xnor U9659 (N_9659,N_5065,N_5878);
nand U9660 (N_9660,N_7053,N_7624);
nor U9661 (N_9661,N_4483,N_6935);
nor U9662 (N_9662,N_5011,N_7342);
nand U9663 (N_9663,N_7352,N_5552);
and U9664 (N_9664,N_4766,N_7679);
and U9665 (N_9665,N_4905,N_7976);
nor U9666 (N_9666,N_5282,N_6179);
nor U9667 (N_9667,N_7179,N_4912);
nor U9668 (N_9668,N_7878,N_5157);
nor U9669 (N_9669,N_7198,N_4667);
or U9670 (N_9670,N_7947,N_7171);
or U9671 (N_9671,N_4841,N_5493);
and U9672 (N_9672,N_4457,N_6799);
xnor U9673 (N_9673,N_6322,N_6004);
or U9674 (N_9674,N_6838,N_6757);
nand U9675 (N_9675,N_4919,N_5226);
nand U9676 (N_9676,N_6086,N_5128);
nand U9677 (N_9677,N_7332,N_7548);
nand U9678 (N_9678,N_6491,N_7927);
nor U9679 (N_9679,N_4333,N_7383);
nand U9680 (N_9680,N_4940,N_5510);
nor U9681 (N_9681,N_6751,N_5673);
or U9682 (N_9682,N_7985,N_5737);
and U9683 (N_9683,N_7866,N_5871);
xnor U9684 (N_9684,N_6406,N_6237);
nor U9685 (N_9685,N_6166,N_6262);
or U9686 (N_9686,N_4405,N_6744);
and U9687 (N_9687,N_7944,N_5568);
and U9688 (N_9688,N_6361,N_4634);
or U9689 (N_9689,N_6119,N_5521);
nand U9690 (N_9690,N_6063,N_4809);
xor U9691 (N_9691,N_7146,N_5382);
nor U9692 (N_9692,N_4139,N_5903);
nor U9693 (N_9693,N_5540,N_4452);
or U9694 (N_9694,N_7478,N_5149);
nand U9695 (N_9695,N_4845,N_4069);
xor U9696 (N_9696,N_5774,N_5623);
nand U9697 (N_9697,N_6937,N_6455);
xnor U9698 (N_9698,N_7820,N_5056);
nand U9699 (N_9699,N_7126,N_6453);
or U9700 (N_9700,N_6085,N_4302);
or U9701 (N_9701,N_4187,N_6831);
or U9702 (N_9702,N_5627,N_7515);
or U9703 (N_9703,N_6657,N_7904);
xor U9704 (N_9704,N_5824,N_7485);
and U9705 (N_9705,N_7582,N_5122);
nand U9706 (N_9706,N_7009,N_7488);
nor U9707 (N_9707,N_4887,N_6044);
and U9708 (N_9708,N_5310,N_6296);
and U9709 (N_9709,N_7036,N_7694);
and U9710 (N_9710,N_5798,N_7282);
and U9711 (N_9711,N_6190,N_7720);
and U9712 (N_9712,N_4031,N_5134);
nor U9713 (N_9713,N_4694,N_6690);
and U9714 (N_9714,N_5557,N_5393);
and U9715 (N_9715,N_7885,N_5130);
and U9716 (N_9716,N_7396,N_7559);
and U9717 (N_9717,N_6187,N_4141);
and U9718 (N_9718,N_5732,N_7430);
nor U9719 (N_9719,N_6315,N_5114);
and U9720 (N_9720,N_7080,N_6443);
nand U9721 (N_9721,N_4648,N_4442);
and U9722 (N_9722,N_4686,N_7871);
or U9723 (N_9723,N_7908,N_7357);
or U9724 (N_9724,N_4688,N_5170);
or U9725 (N_9725,N_6980,N_5363);
nor U9726 (N_9726,N_4129,N_5232);
nor U9727 (N_9727,N_6272,N_4049);
and U9728 (N_9728,N_5840,N_5819);
nand U9729 (N_9729,N_4359,N_6513);
nor U9730 (N_9730,N_7366,N_6414);
or U9731 (N_9731,N_6702,N_6449);
or U9732 (N_9732,N_6328,N_6139);
xor U9733 (N_9733,N_7740,N_6006);
nor U9734 (N_9734,N_7707,N_4711);
and U9735 (N_9735,N_5596,N_5079);
or U9736 (N_9736,N_5587,N_4473);
nor U9737 (N_9737,N_6502,N_6493);
or U9738 (N_9738,N_7416,N_7293);
nor U9739 (N_9739,N_5352,N_4646);
nand U9740 (N_9740,N_7857,N_7390);
and U9741 (N_9741,N_6692,N_4003);
nand U9742 (N_9742,N_4469,N_4611);
nor U9743 (N_9743,N_7408,N_4752);
and U9744 (N_9744,N_4207,N_4980);
and U9745 (N_9745,N_7251,N_6146);
xor U9746 (N_9746,N_5101,N_5797);
or U9747 (N_9747,N_7792,N_5150);
nor U9748 (N_9748,N_7385,N_5242);
nor U9749 (N_9749,N_6389,N_7215);
nor U9750 (N_9750,N_4999,N_7418);
and U9751 (N_9751,N_6327,N_4298);
xnor U9752 (N_9752,N_6985,N_6318);
nor U9753 (N_9753,N_7982,N_6977);
and U9754 (N_9754,N_6213,N_6903);
nor U9755 (N_9755,N_6197,N_4435);
nand U9756 (N_9756,N_5786,N_4378);
or U9757 (N_9757,N_7892,N_7598);
nor U9758 (N_9758,N_6515,N_6351);
xnor U9759 (N_9759,N_4205,N_7192);
and U9760 (N_9760,N_5285,N_5657);
nor U9761 (N_9761,N_6748,N_5455);
and U9762 (N_9762,N_5211,N_4596);
xor U9763 (N_9763,N_7709,N_7458);
or U9764 (N_9764,N_6715,N_5930);
nand U9765 (N_9765,N_5115,N_7089);
nor U9766 (N_9766,N_7081,N_6820);
and U9767 (N_9767,N_4813,N_4811);
nor U9768 (N_9768,N_4036,N_4236);
nor U9769 (N_9769,N_6359,N_7710);
or U9770 (N_9770,N_5272,N_5404);
and U9771 (N_9771,N_5301,N_5349);
or U9772 (N_9772,N_7162,N_5022);
nand U9773 (N_9773,N_5678,N_5486);
nor U9774 (N_9774,N_7083,N_4110);
or U9775 (N_9775,N_4151,N_4293);
or U9776 (N_9776,N_6611,N_7761);
or U9777 (N_9777,N_7711,N_6138);
nor U9778 (N_9778,N_5601,N_6225);
nor U9779 (N_9779,N_6199,N_5327);
xor U9780 (N_9780,N_5477,N_6896);
and U9781 (N_9781,N_7254,N_7015);
nand U9782 (N_9782,N_4528,N_4741);
nand U9783 (N_9783,N_5845,N_5146);
nor U9784 (N_9784,N_6989,N_5868);
nor U9785 (N_9785,N_5234,N_5203);
nor U9786 (N_9786,N_6172,N_6720);
or U9787 (N_9787,N_4668,N_4623);
nand U9788 (N_9788,N_6428,N_7399);
xor U9789 (N_9789,N_6765,N_5512);
nand U9790 (N_9790,N_5809,N_6616);
and U9791 (N_9791,N_4465,N_6640);
and U9792 (N_9792,N_4950,N_7026);
and U9793 (N_9793,N_4337,N_6274);
and U9794 (N_9794,N_4228,N_6590);
nand U9795 (N_9795,N_5944,N_4737);
nand U9796 (N_9796,N_4734,N_4444);
nor U9797 (N_9797,N_6796,N_4524);
xor U9798 (N_9798,N_6735,N_4067);
nand U9799 (N_9799,N_6391,N_5348);
and U9800 (N_9800,N_4425,N_6862);
nand U9801 (N_9801,N_5461,N_4708);
or U9802 (N_9802,N_6620,N_4014);
nand U9803 (N_9803,N_7237,N_6761);
nand U9804 (N_9804,N_5053,N_6972);
nand U9805 (N_9805,N_4995,N_6317);
nand U9806 (N_9806,N_4888,N_6745);
nor U9807 (N_9807,N_6071,N_4886);
or U9808 (N_9808,N_7271,N_5308);
nor U9809 (N_9809,N_5112,N_5585);
nor U9810 (N_9810,N_6981,N_4831);
nor U9811 (N_9811,N_7998,N_6243);
xnor U9812 (N_9812,N_5793,N_7278);
nor U9813 (N_9813,N_6707,N_5744);
nor U9814 (N_9814,N_7202,N_7847);
nor U9815 (N_9815,N_5454,N_7417);
nand U9816 (N_9816,N_7595,N_4576);
nor U9817 (N_9817,N_5362,N_5787);
or U9818 (N_9818,N_6128,N_4123);
nand U9819 (N_9819,N_4630,N_6724);
nand U9820 (N_9820,N_6795,N_6445);
and U9821 (N_9821,N_6009,N_4044);
nor U9822 (N_9822,N_4990,N_5453);
nor U9823 (N_9823,N_6923,N_6964);
nor U9824 (N_9824,N_7898,N_6837);
and U9825 (N_9825,N_6912,N_6284);
nand U9826 (N_9826,N_6373,N_4691);
nor U9827 (N_9827,N_5241,N_4769);
or U9828 (N_9828,N_5956,N_6569);
and U9829 (N_9829,N_5121,N_7134);
xnor U9830 (N_9830,N_4947,N_4356);
and U9831 (N_9831,N_4533,N_4157);
nor U9832 (N_9832,N_4775,N_4137);
or U9833 (N_9833,N_7808,N_5780);
xnor U9834 (N_9834,N_4645,N_4892);
nand U9835 (N_9835,N_7697,N_7846);
nand U9836 (N_9836,N_6397,N_5977);
or U9837 (N_9837,N_6655,N_4690);
nand U9838 (N_9838,N_7805,N_6869);
nand U9839 (N_9839,N_7531,N_6346);
and U9840 (N_9840,N_4671,N_7688);
or U9841 (N_9841,N_6732,N_7051);
and U9842 (N_9842,N_7165,N_6890);
nand U9843 (N_9843,N_5032,N_6917);
and U9844 (N_9844,N_6949,N_6465);
xnor U9845 (N_9845,N_5676,N_5041);
xor U9846 (N_9846,N_5293,N_5216);
or U9847 (N_9847,N_5098,N_7816);
nor U9848 (N_9848,N_7543,N_5590);
and U9849 (N_9849,N_4653,N_7445);
nand U9850 (N_9850,N_4718,N_5303);
and U9851 (N_9851,N_4843,N_5532);
nor U9852 (N_9852,N_7663,N_5379);
nand U9853 (N_9853,N_7722,N_5168);
and U9854 (N_9854,N_7609,N_5885);
nand U9855 (N_9855,N_6853,N_7356);
or U9856 (N_9856,N_4181,N_7766);
nor U9857 (N_9857,N_6857,N_5010);
and U9858 (N_9858,N_7489,N_4649);
or U9859 (N_9859,N_4055,N_6407);
nand U9860 (N_9860,N_4512,N_6399);
nor U9861 (N_9861,N_6231,N_7517);
nand U9862 (N_9862,N_6827,N_7762);
nor U9863 (N_9863,N_7465,N_5758);
or U9864 (N_9864,N_7345,N_6114);
nor U9865 (N_9865,N_7294,N_4928);
and U9866 (N_9866,N_5998,N_5094);
nand U9867 (N_9867,N_7839,N_7674);
nand U9868 (N_9868,N_4374,N_6886);
and U9869 (N_9869,N_5325,N_4382);
nand U9870 (N_9870,N_7501,N_5267);
and U9871 (N_9871,N_6573,N_6563);
nor U9872 (N_9872,N_4340,N_7493);
nor U9873 (N_9873,N_4499,N_5074);
or U9874 (N_9874,N_4773,N_6202);
or U9875 (N_9875,N_5966,N_4610);
and U9876 (N_9876,N_5900,N_6051);
or U9877 (N_9877,N_7046,N_4542);
and U9878 (N_9878,N_5571,N_7090);
or U9879 (N_9879,N_4331,N_5438);
nand U9880 (N_9880,N_5415,N_5880);
or U9881 (N_9881,N_7013,N_4273);
and U9882 (N_9882,N_7521,N_5435);
and U9883 (N_9883,N_6256,N_5173);
nor U9884 (N_9884,N_6918,N_4480);
nor U9885 (N_9885,N_6168,N_4380);
and U9886 (N_9886,N_6133,N_4280);
nor U9887 (N_9887,N_5019,N_5530);
nor U9888 (N_9888,N_7178,N_4577);
and U9889 (N_9889,N_6188,N_4951);
nor U9890 (N_9890,N_5095,N_4516);
nand U9891 (N_9891,N_5586,N_5261);
and U9892 (N_9892,N_6582,N_7757);
and U9893 (N_9893,N_4259,N_6887);
nand U9894 (N_9894,N_7692,N_7838);
xnor U9895 (N_9895,N_4788,N_4175);
nand U9896 (N_9896,N_5035,N_5834);
nor U9897 (N_9897,N_6037,N_7141);
and U9898 (N_9898,N_6282,N_5239);
or U9899 (N_9899,N_6417,N_7952);
or U9900 (N_9900,N_7628,N_5283);
or U9901 (N_9901,N_4978,N_6561);
or U9902 (N_9902,N_6621,N_6703);
and U9903 (N_9903,N_6726,N_4287);
nor U9904 (N_9904,N_4439,N_5822);
xnor U9905 (N_9905,N_7070,N_5802);
nand U9906 (N_9906,N_4053,N_7961);
nor U9907 (N_9907,N_6978,N_6847);
or U9908 (N_9908,N_6882,N_4830);
and U9909 (N_9909,N_6880,N_6610);
nand U9910 (N_9910,N_5662,N_5322);
nor U9911 (N_9911,N_7969,N_5539);
or U9912 (N_9912,N_5229,N_7977);
nor U9913 (N_9913,N_7377,N_5996);
or U9914 (N_9914,N_5718,N_6548);
nand U9915 (N_9915,N_4342,N_6931);
nor U9916 (N_9916,N_4550,N_6441);
and U9917 (N_9917,N_4633,N_7457);
and U9918 (N_9918,N_6914,N_6340);
xnor U9919 (N_9919,N_6165,N_6546);
or U9920 (N_9920,N_7075,N_4719);
nor U9921 (N_9921,N_6092,N_5511);
or U9922 (N_9922,N_4712,N_6580);
nor U9923 (N_9923,N_7188,N_5313);
or U9924 (N_9924,N_5106,N_4081);
nor U9925 (N_9925,N_4638,N_6901);
and U9926 (N_9926,N_7669,N_7545);
or U9927 (N_9927,N_4039,N_4384);
nand U9928 (N_9928,N_4874,N_6717);
nand U9929 (N_9929,N_6746,N_5240);
nor U9930 (N_9930,N_4846,N_4749);
and U9931 (N_9931,N_6186,N_7219);
nand U9932 (N_9932,N_4602,N_6941);
nand U9933 (N_9933,N_6930,N_4400);
nor U9934 (N_9934,N_7535,N_6095);
xnor U9935 (N_9935,N_5958,N_6627);
nand U9936 (N_9936,N_5843,N_7305);
nand U9937 (N_9937,N_7861,N_7038);
nor U9938 (N_9938,N_4006,N_4783);
nor U9939 (N_9939,N_5473,N_6261);
nand U9940 (N_9940,N_5922,N_6061);
nor U9941 (N_9941,N_7480,N_7862);
and U9942 (N_9942,N_7718,N_4873);
xor U9943 (N_9943,N_4697,N_5579);
xnor U9944 (N_9944,N_7218,N_7350);
nor U9945 (N_9945,N_7929,N_6711);
nor U9946 (N_9946,N_4135,N_7433);
xnor U9947 (N_9947,N_6118,N_5589);
nor U9948 (N_9948,N_4600,N_4825);
xnor U9949 (N_9949,N_4362,N_7405);
or U9950 (N_9950,N_7229,N_4332);
nand U9951 (N_9951,N_6974,N_6665);
nand U9952 (N_9952,N_7779,N_7853);
or U9953 (N_9953,N_7657,N_4349);
and U9954 (N_9954,N_5187,N_7602);
nand U9955 (N_9955,N_7505,N_6132);
and U9956 (N_9956,N_7523,N_4472);
or U9957 (N_9957,N_7671,N_5931);
and U9958 (N_9958,N_4523,N_4955);
or U9959 (N_9959,N_5536,N_4798);
xor U9960 (N_9960,N_5158,N_7622);
and U9961 (N_9961,N_7967,N_6771);
nand U9962 (N_9962,N_6527,N_4052);
nand U9963 (N_9963,N_7027,N_7411);
and U9964 (N_9964,N_4506,N_7471);
or U9965 (N_9965,N_4344,N_4256);
nor U9966 (N_9966,N_6275,N_7068);
or U9967 (N_9967,N_5514,N_5364);
xor U9968 (N_9968,N_6125,N_6394);
nand U9969 (N_9969,N_7570,N_5534);
and U9970 (N_9970,N_4117,N_4013);
and U9971 (N_9971,N_7621,N_6782);
or U9972 (N_9972,N_5560,N_7299);
and U9973 (N_9973,N_6828,N_6756);
and U9974 (N_9974,N_7180,N_6566);
nor U9975 (N_9975,N_5504,N_5790);
nor U9976 (N_9976,N_6258,N_7616);
and U9977 (N_9977,N_4584,N_7012);
xnor U9978 (N_9978,N_5773,N_4958);
or U9979 (N_9979,N_6777,N_7401);
nand U9980 (N_9980,N_4078,N_5870);
or U9981 (N_9981,N_5373,N_4224);
xnor U9982 (N_9982,N_4255,N_6170);
nand U9983 (N_9983,N_7379,N_7903);
nand U9984 (N_9984,N_4562,N_4992);
and U9985 (N_9985,N_7841,N_7951);
and U9986 (N_9986,N_7274,N_5244);
and U9987 (N_9987,N_5081,N_4890);
nor U9988 (N_9988,N_5033,N_6518);
nand U9989 (N_9989,N_7675,N_5439);
xnor U9990 (N_9990,N_5979,N_7064);
nor U9991 (N_9991,N_7368,N_5509);
and U9992 (N_9992,N_4361,N_6298);
nor U9993 (N_9993,N_4589,N_6570);
nand U9994 (N_9994,N_7748,N_4087);
nand U9995 (N_9995,N_4974,N_4321);
xnor U9996 (N_9996,N_5474,N_6255);
and U9997 (N_9997,N_7346,N_6966);
nor U9998 (N_9998,N_6038,N_7095);
and U9999 (N_9999,N_4606,N_6281);
or U10000 (N_10000,N_7966,N_5166);
nor U10001 (N_10001,N_7210,N_5754);
nand U10002 (N_10002,N_7882,N_4355);
nor U10003 (N_10003,N_4710,N_6196);
or U10004 (N_10004,N_4793,N_4177);
or U10005 (N_10005,N_4773,N_5462);
or U10006 (N_10006,N_6986,N_7935);
nand U10007 (N_10007,N_4073,N_6970);
nor U10008 (N_10008,N_4908,N_6865);
and U10009 (N_10009,N_4390,N_6055);
nand U10010 (N_10010,N_4845,N_7958);
or U10011 (N_10011,N_6923,N_7621);
and U10012 (N_10012,N_6175,N_6547);
or U10013 (N_10013,N_5346,N_6909);
nand U10014 (N_10014,N_6988,N_6550);
or U10015 (N_10015,N_4471,N_4969);
xnor U10016 (N_10016,N_6885,N_7902);
and U10017 (N_10017,N_4479,N_5898);
nand U10018 (N_10018,N_4187,N_5194);
nand U10019 (N_10019,N_7651,N_4570);
nor U10020 (N_10020,N_7981,N_5271);
nand U10021 (N_10021,N_4751,N_4603);
and U10022 (N_10022,N_7584,N_5882);
or U10023 (N_10023,N_7043,N_5514);
or U10024 (N_10024,N_6135,N_7158);
nor U10025 (N_10025,N_7974,N_4976);
or U10026 (N_10026,N_6191,N_5143);
nand U10027 (N_10027,N_7150,N_7169);
nor U10028 (N_10028,N_6005,N_5516);
nor U10029 (N_10029,N_5653,N_5693);
or U10030 (N_10030,N_7871,N_6455);
nor U10031 (N_10031,N_6576,N_6112);
and U10032 (N_10032,N_4260,N_7167);
xnor U10033 (N_10033,N_7984,N_5434);
and U10034 (N_10034,N_6684,N_4451);
xnor U10035 (N_10035,N_4048,N_5657);
and U10036 (N_10036,N_6082,N_4570);
xor U10037 (N_10037,N_4802,N_6619);
and U10038 (N_10038,N_7518,N_5752);
nand U10039 (N_10039,N_5618,N_5856);
nand U10040 (N_10040,N_6469,N_5618);
nand U10041 (N_10041,N_4647,N_7345);
nor U10042 (N_10042,N_5054,N_4086);
nand U10043 (N_10043,N_5079,N_5170);
nor U10044 (N_10044,N_6646,N_7106);
or U10045 (N_10045,N_6285,N_6591);
nor U10046 (N_10046,N_4122,N_4285);
nor U10047 (N_10047,N_5477,N_5522);
nor U10048 (N_10048,N_6008,N_4693);
nor U10049 (N_10049,N_6934,N_5241);
or U10050 (N_10050,N_6037,N_5544);
nor U10051 (N_10051,N_5919,N_7782);
nand U10052 (N_10052,N_4911,N_4102);
and U10053 (N_10053,N_6245,N_6879);
nand U10054 (N_10054,N_4470,N_6142);
nand U10055 (N_10055,N_7994,N_6578);
and U10056 (N_10056,N_7281,N_4967);
or U10057 (N_10057,N_4344,N_7119);
xnor U10058 (N_10058,N_6045,N_7245);
or U10059 (N_10059,N_7948,N_4654);
and U10060 (N_10060,N_4569,N_4103);
and U10061 (N_10061,N_4268,N_4194);
or U10062 (N_10062,N_5578,N_6268);
and U10063 (N_10063,N_6952,N_7960);
nand U10064 (N_10064,N_4852,N_5709);
and U10065 (N_10065,N_4285,N_5211);
nor U10066 (N_10066,N_7827,N_5356);
or U10067 (N_10067,N_4383,N_4585);
and U10068 (N_10068,N_6715,N_5048);
and U10069 (N_10069,N_5396,N_5112);
nand U10070 (N_10070,N_4699,N_7141);
nor U10071 (N_10071,N_5864,N_5854);
and U10072 (N_10072,N_7145,N_5431);
or U10073 (N_10073,N_4019,N_4041);
nor U10074 (N_10074,N_4778,N_7729);
and U10075 (N_10075,N_7068,N_6700);
and U10076 (N_10076,N_6619,N_4554);
and U10077 (N_10077,N_6918,N_6384);
and U10078 (N_10078,N_5211,N_7298);
and U10079 (N_10079,N_5417,N_6016);
and U10080 (N_10080,N_7386,N_6437);
nand U10081 (N_10081,N_7473,N_4626);
or U10082 (N_10082,N_6996,N_4755);
nand U10083 (N_10083,N_4182,N_7149);
and U10084 (N_10084,N_7240,N_4054);
and U10085 (N_10085,N_6593,N_5387);
nand U10086 (N_10086,N_6145,N_7157);
xor U10087 (N_10087,N_6924,N_5972);
or U10088 (N_10088,N_6519,N_7504);
and U10089 (N_10089,N_5416,N_7886);
nand U10090 (N_10090,N_6433,N_7017);
nor U10091 (N_10091,N_6775,N_7309);
xor U10092 (N_10092,N_6164,N_6798);
or U10093 (N_10093,N_5508,N_6198);
xnor U10094 (N_10094,N_6663,N_5176);
and U10095 (N_10095,N_7503,N_5690);
and U10096 (N_10096,N_4671,N_7012);
nand U10097 (N_10097,N_6217,N_7491);
and U10098 (N_10098,N_6060,N_6863);
or U10099 (N_10099,N_7230,N_6651);
and U10100 (N_10100,N_6598,N_5114);
nor U10101 (N_10101,N_6010,N_5924);
or U10102 (N_10102,N_5185,N_7934);
nand U10103 (N_10103,N_6249,N_5266);
nand U10104 (N_10104,N_6155,N_7375);
nand U10105 (N_10105,N_6315,N_5684);
and U10106 (N_10106,N_7013,N_4904);
nor U10107 (N_10107,N_5822,N_4464);
or U10108 (N_10108,N_5037,N_5249);
or U10109 (N_10109,N_7304,N_6084);
nor U10110 (N_10110,N_5263,N_7362);
nand U10111 (N_10111,N_5307,N_5848);
xor U10112 (N_10112,N_4530,N_7837);
and U10113 (N_10113,N_4798,N_5879);
nand U10114 (N_10114,N_4575,N_6621);
nor U10115 (N_10115,N_5148,N_4849);
and U10116 (N_10116,N_5470,N_4012);
nand U10117 (N_10117,N_4908,N_6027);
xnor U10118 (N_10118,N_6934,N_4269);
xnor U10119 (N_10119,N_5209,N_6250);
or U10120 (N_10120,N_6924,N_7869);
and U10121 (N_10121,N_6662,N_6969);
xor U10122 (N_10122,N_5572,N_6831);
nor U10123 (N_10123,N_6503,N_5798);
nor U10124 (N_10124,N_5452,N_7711);
nor U10125 (N_10125,N_6500,N_6551);
nor U10126 (N_10126,N_4412,N_7516);
and U10127 (N_10127,N_4764,N_5817);
or U10128 (N_10128,N_4740,N_6381);
and U10129 (N_10129,N_4420,N_6921);
nand U10130 (N_10130,N_6604,N_4693);
nor U10131 (N_10131,N_7082,N_5885);
or U10132 (N_10132,N_4213,N_4689);
or U10133 (N_10133,N_7076,N_7885);
and U10134 (N_10134,N_6495,N_7660);
nand U10135 (N_10135,N_7825,N_7677);
or U10136 (N_10136,N_5742,N_4403);
and U10137 (N_10137,N_6276,N_7972);
xor U10138 (N_10138,N_7741,N_5790);
and U10139 (N_10139,N_4028,N_6641);
nand U10140 (N_10140,N_6409,N_7741);
and U10141 (N_10141,N_6445,N_7875);
or U10142 (N_10142,N_5546,N_4355);
nand U10143 (N_10143,N_7424,N_5409);
nor U10144 (N_10144,N_6541,N_5005);
xor U10145 (N_10145,N_4474,N_6794);
or U10146 (N_10146,N_7457,N_6179);
and U10147 (N_10147,N_6082,N_5000);
nor U10148 (N_10148,N_4143,N_6445);
nor U10149 (N_10149,N_7782,N_4009);
nor U10150 (N_10150,N_4921,N_5333);
nor U10151 (N_10151,N_6604,N_5878);
and U10152 (N_10152,N_6425,N_7838);
or U10153 (N_10153,N_7259,N_6915);
nor U10154 (N_10154,N_5969,N_7606);
or U10155 (N_10155,N_7043,N_6573);
nand U10156 (N_10156,N_6217,N_5823);
or U10157 (N_10157,N_5046,N_5747);
and U10158 (N_10158,N_7352,N_7943);
and U10159 (N_10159,N_4479,N_4526);
nand U10160 (N_10160,N_5089,N_5563);
or U10161 (N_10161,N_7955,N_5076);
and U10162 (N_10162,N_7393,N_4712);
nand U10163 (N_10163,N_5749,N_6877);
and U10164 (N_10164,N_7829,N_7990);
and U10165 (N_10165,N_4448,N_4498);
and U10166 (N_10166,N_4894,N_4274);
nand U10167 (N_10167,N_4006,N_4122);
and U10168 (N_10168,N_6355,N_7037);
nand U10169 (N_10169,N_5236,N_7129);
and U10170 (N_10170,N_4753,N_7745);
nand U10171 (N_10171,N_7991,N_5272);
and U10172 (N_10172,N_5898,N_6257);
nor U10173 (N_10173,N_4931,N_7954);
nor U10174 (N_10174,N_5274,N_7342);
nor U10175 (N_10175,N_7123,N_7498);
or U10176 (N_10176,N_6661,N_7130);
nor U10177 (N_10177,N_6446,N_4085);
or U10178 (N_10178,N_5744,N_4653);
nor U10179 (N_10179,N_5725,N_7055);
nand U10180 (N_10180,N_7779,N_6904);
and U10181 (N_10181,N_6832,N_4968);
and U10182 (N_10182,N_6081,N_4803);
nor U10183 (N_10183,N_6686,N_5493);
nand U10184 (N_10184,N_7958,N_4328);
and U10185 (N_10185,N_7388,N_6499);
and U10186 (N_10186,N_4614,N_7714);
or U10187 (N_10187,N_7937,N_5603);
or U10188 (N_10188,N_5599,N_4990);
or U10189 (N_10189,N_5258,N_5364);
or U10190 (N_10190,N_5049,N_5168);
or U10191 (N_10191,N_7985,N_7905);
nor U10192 (N_10192,N_4216,N_4561);
nor U10193 (N_10193,N_4895,N_7531);
and U10194 (N_10194,N_4896,N_4348);
and U10195 (N_10195,N_6208,N_6762);
nand U10196 (N_10196,N_7715,N_5485);
nor U10197 (N_10197,N_7427,N_4453);
nand U10198 (N_10198,N_6903,N_7684);
nand U10199 (N_10199,N_4333,N_6638);
nor U10200 (N_10200,N_4070,N_5525);
xnor U10201 (N_10201,N_6457,N_6763);
nand U10202 (N_10202,N_5991,N_4314);
nor U10203 (N_10203,N_5751,N_5533);
nor U10204 (N_10204,N_6521,N_5783);
or U10205 (N_10205,N_6368,N_7488);
or U10206 (N_10206,N_5699,N_6396);
and U10207 (N_10207,N_6630,N_6064);
xor U10208 (N_10208,N_6420,N_5996);
nand U10209 (N_10209,N_5104,N_7759);
nand U10210 (N_10210,N_4080,N_6202);
nor U10211 (N_10211,N_6174,N_5189);
nand U10212 (N_10212,N_4335,N_7461);
nor U10213 (N_10213,N_6107,N_4214);
nor U10214 (N_10214,N_6222,N_7591);
nor U10215 (N_10215,N_6232,N_4278);
and U10216 (N_10216,N_5040,N_4481);
nand U10217 (N_10217,N_6890,N_7979);
nand U10218 (N_10218,N_7303,N_4461);
xor U10219 (N_10219,N_4635,N_6895);
nor U10220 (N_10220,N_5315,N_6145);
nor U10221 (N_10221,N_6726,N_6938);
nor U10222 (N_10222,N_7488,N_7161);
nor U10223 (N_10223,N_7318,N_5536);
or U10224 (N_10224,N_4153,N_4875);
nor U10225 (N_10225,N_4593,N_5402);
or U10226 (N_10226,N_4251,N_7085);
and U10227 (N_10227,N_5897,N_4321);
nand U10228 (N_10228,N_5177,N_5377);
nand U10229 (N_10229,N_7541,N_5172);
nor U10230 (N_10230,N_6401,N_6725);
nand U10231 (N_10231,N_7878,N_5682);
xor U10232 (N_10232,N_5074,N_6042);
or U10233 (N_10233,N_7269,N_6873);
nand U10234 (N_10234,N_6417,N_4643);
or U10235 (N_10235,N_7690,N_7129);
nor U10236 (N_10236,N_5384,N_5060);
nand U10237 (N_10237,N_5885,N_7648);
nand U10238 (N_10238,N_5575,N_4688);
nor U10239 (N_10239,N_4394,N_4049);
or U10240 (N_10240,N_6970,N_4289);
xnor U10241 (N_10241,N_7968,N_5755);
xnor U10242 (N_10242,N_4972,N_7299);
or U10243 (N_10243,N_6408,N_4941);
or U10244 (N_10244,N_4037,N_6029);
and U10245 (N_10245,N_6588,N_5269);
xor U10246 (N_10246,N_6230,N_6718);
nand U10247 (N_10247,N_4460,N_6806);
or U10248 (N_10248,N_5420,N_7563);
nor U10249 (N_10249,N_4799,N_6590);
nand U10250 (N_10250,N_6353,N_6472);
and U10251 (N_10251,N_4554,N_6545);
and U10252 (N_10252,N_4996,N_4406);
and U10253 (N_10253,N_5673,N_5024);
or U10254 (N_10254,N_6112,N_7545);
or U10255 (N_10255,N_5575,N_5375);
or U10256 (N_10256,N_4957,N_7149);
nor U10257 (N_10257,N_5403,N_4964);
and U10258 (N_10258,N_6983,N_6214);
nor U10259 (N_10259,N_4523,N_6582);
nor U10260 (N_10260,N_5816,N_4323);
xnor U10261 (N_10261,N_6648,N_6917);
nor U10262 (N_10262,N_6569,N_6233);
xnor U10263 (N_10263,N_7188,N_5256);
nor U10264 (N_10264,N_7061,N_4444);
or U10265 (N_10265,N_5965,N_6185);
or U10266 (N_10266,N_7589,N_6959);
nand U10267 (N_10267,N_4579,N_5555);
nor U10268 (N_10268,N_6962,N_7613);
and U10269 (N_10269,N_7700,N_4947);
and U10270 (N_10270,N_7013,N_5435);
or U10271 (N_10271,N_5977,N_4346);
nor U10272 (N_10272,N_5405,N_6774);
nand U10273 (N_10273,N_7061,N_5633);
nor U10274 (N_10274,N_5154,N_4392);
or U10275 (N_10275,N_5860,N_4290);
nor U10276 (N_10276,N_5335,N_6457);
xor U10277 (N_10277,N_4095,N_6546);
nor U10278 (N_10278,N_5489,N_4568);
and U10279 (N_10279,N_6939,N_5456);
nand U10280 (N_10280,N_6110,N_7615);
or U10281 (N_10281,N_5126,N_7906);
and U10282 (N_10282,N_6479,N_6923);
xor U10283 (N_10283,N_6802,N_5006);
nor U10284 (N_10284,N_7147,N_5597);
or U10285 (N_10285,N_5348,N_7563);
or U10286 (N_10286,N_6418,N_7955);
xnor U10287 (N_10287,N_6647,N_4483);
or U10288 (N_10288,N_4716,N_4298);
nand U10289 (N_10289,N_7495,N_7104);
or U10290 (N_10290,N_4939,N_7233);
or U10291 (N_10291,N_6364,N_6766);
nor U10292 (N_10292,N_4859,N_4289);
nor U10293 (N_10293,N_4740,N_6740);
nand U10294 (N_10294,N_4252,N_4158);
xnor U10295 (N_10295,N_7768,N_4852);
nand U10296 (N_10296,N_4618,N_5922);
or U10297 (N_10297,N_6314,N_4246);
or U10298 (N_10298,N_6093,N_5588);
nor U10299 (N_10299,N_6774,N_7381);
nor U10300 (N_10300,N_5290,N_7729);
and U10301 (N_10301,N_5812,N_6565);
or U10302 (N_10302,N_5097,N_4842);
nand U10303 (N_10303,N_4938,N_4653);
and U10304 (N_10304,N_6064,N_5580);
nand U10305 (N_10305,N_4144,N_4627);
nand U10306 (N_10306,N_4998,N_5290);
or U10307 (N_10307,N_5389,N_4438);
nand U10308 (N_10308,N_4576,N_5820);
and U10309 (N_10309,N_7395,N_6627);
xnor U10310 (N_10310,N_7762,N_7184);
nand U10311 (N_10311,N_6257,N_5438);
nand U10312 (N_10312,N_6935,N_5118);
nor U10313 (N_10313,N_7449,N_6963);
xnor U10314 (N_10314,N_6180,N_7739);
or U10315 (N_10315,N_7050,N_4441);
and U10316 (N_10316,N_4732,N_5855);
or U10317 (N_10317,N_7647,N_6432);
or U10318 (N_10318,N_7414,N_6296);
and U10319 (N_10319,N_5066,N_5842);
nand U10320 (N_10320,N_7586,N_7520);
nor U10321 (N_10321,N_5932,N_6527);
nand U10322 (N_10322,N_7351,N_5022);
and U10323 (N_10323,N_4109,N_6032);
and U10324 (N_10324,N_7577,N_7153);
nand U10325 (N_10325,N_7179,N_6305);
and U10326 (N_10326,N_5054,N_7959);
or U10327 (N_10327,N_7993,N_7443);
xor U10328 (N_10328,N_4358,N_5600);
or U10329 (N_10329,N_4174,N_5062);
or U10330 (N_10330,N_6389,N_4463);
and U10331 (N_10331,N_7440,N_6479);
or U10332 (N_10332,N_7081,N_6919);
or U10333 (N_10333,N_5037,N_7069);
or U10334 (N_10334,N_6418,N_6854);
nand U10335 (N_10335,N_7269,N_6976);
nand U10336 (N_10336,N_7352,N_7715);
nand U10337 (N_10337,N_6497,N_6684);
or U10338 (N_10338,N_7568,N_6696);
nor U10339 (N_10339,N_4034,N_5397);
or U10340 (N_10340,N_5002,N_6219);
nor U10341 (N_10341,N_4323,N_4050);
xor U10342 (N_10342,N_7192,N_4321);
nor U10343 (N_10343,N_6990,N_7048);
nand U10344 (N_10344,N_5636,N_7256);
nand U10345 (N_10345,N_4504,N_5920);
nand U10346 (N_10346,N_5637,N_4273);
and U10347 (N_10347,N_5507,N_4384);
nor U10348 (N_10348,N_7684,N_7357);
and U10349 (N_10349,N_5831,N_6451);
nor U10350 (N_10350,N_4706,N_6913);
nand U10351 (N_10351,N_5352,N_6853);
xor U10352 (N_10352,N_4247,N_5728);
or U10353 (N_10353,N_4799,N_4793);
xor U10354 (N_10354,N_6149,N_4390);
or U10355 (N_10355,N_4913,N_6037);
and U10356 (N_10356,N_6870,N_4676);
nor U10357 (N_10357,N_5230,N_4553);
nand U10358 (N_10358,N_7238,N_4358);
nand U10359 (N_10359,N_6681,N_7799);
and U10360 (N_10360,N_4011,N_6394);
nand U10361 (N_10361,N_6961,N_4515);
nor U10362 (N_10362,N_7429,N_4087);
nand U10363 (N_10363,N_7619,N_5327);
or U10364 (N_10364,N_7758,N_6364);
or U10365 (N_10365,N_7104,N_6197);
and U10366 (N_10366,N_5744,N_4616);
nand U10367 (N_10367,N_4079,N_5061);
nor U10368 (N_10368,N_5707,N_4260);
and U10369 (N_10369,N_7737,N_4781);
nor U10370 (N_10370,N_5974,N_5165);
nand U10371 (N_10371,N_4372,N_4881);
nor U10372 (N_10372,N_7233,N_5358);
nor U10373 (N_10373,N_4679,N_4191);
nand U10374 (N_10374,N_4223,N_5213);
or U10375 (N_10375,N_7277,N_4456);
or U10376 (N_10376,N_7105,N_4144);
or U10377 (N_10377,N_4078,N_4598);
nor U10378 (N_10378,N_4787,N_7209);
and U10379 (N_10379,N_6539,N_7095);
or U10380 (N_10380,N_6040,N_7964);
or U10381 (N_10381,N_5815,N_4624);
xnor U10382 (N_10382,N_7590,N_4157);
xnor U10383 (N_10383,N_4602,N_5500);
xnor U10384 (N_10384,N_7973,N_4046);
nor U10385 (N_10385,N_6796,N_7561);
or U10386 (N_10386,N_7930,N_7206);
or U10387 (N_10387,N_7288,N_5897);
or U10388 (N_10388,N_5041,N_4202);
xnor U10389 (N_10389,N_7500,N_5570);
nor U10390 (N_10390,N_5571,N_7363);
nor U10391 (N_10391,N_4937,N_6165);
or U10392 (N_10392,N_7486,N_5184);
nand U10393 (N_10393,N_6829,N_6634);
or U10394 (N_10394,N_7446,N_7455);
nor U10395 (N_10395,N_7181,N_7898);
nand U10396 (N_10396,N_7814,N_4206);
nor U10397 (N_10397,N_7737,N_4391);
nor U10398 (N_10398,N_6437,N_7353);
nand U10399 (N_10399,N_7248,N_5596);
and U10400 (N_10400,N_5911,N_4390);
nand U10401 (N_10401,N_4241,N_4790);
nor U10402 (N_10402,N_6389,N_5988);
nor U10403 (N_10403,N_4036,N_7756);
xnor U10404 (N_10404,N_4917,N_5192);
nor U10405 (N_10405,N_5547,N_5999);
or U10406 (N_10406,N_4439,N_6482);
nand U10407 (N_10407,N_4074,N_7606);
or U10408 (N_10408,N_7915,N_6794);
nor U10409 (N_10409,N_5101,N_6944);
or U10410 (N_10410,N_6793,N_5846);
nor U10411 (N_10411,N_4775,N_4941);
nor U10412 (N_10412,N_7055,N_5287);
or U10413 (N_10413,N_7954,N_7296);
nand U10414 (N_10414,N_5819,N_5990);
nand U10415 (N_10415,N_5044,N_6953);
nand U10416 (N_10416,N_7999,N_7038);
nor U10417 (N_10417,N_5392,N_5574);
or U10418 (N_10418,N_7867,N_6938);
or U10419 (N_10419,N_5631,N_7400);
nand U10420 (N_10420,N_4639,N_5669);
or U10421 (N_10421,N_6367,N_4539);
xor U10422 (N_10422,N_5137,N_4948);
nor U10423 (N_10423,N_4316,N_7026);
nand U10424 (N_10424,N_4640,N_4055);
nor U10425 (N_10425,N_6984,N_7673);
nand U10426 (N_10426,N_5564,N_5885);
nor U10427 (N_10427,N_4025,N_7295);
or U10428 (N_10428,N_7146,N_4781);
nand U10429 (N_10429,N_7748,N_5425);
nand U10430 (N_10430,N_4551,N_6856);
or U10431 (N_10431,N_6142,N_7736);
xor U10432 (N_10432,N_6142,N_6129);
nor U10433 (N_10433,N_5225,N_5833);
nand U10434 (N_10434,N_4257,N_6853);
and U10435 (N_10435,N_6077,N_7791);
xor U10436 (N_10436,N_5075,N_4695);
and U10437 (N_10437,N_6220,N_4122);
and U10438 (N_10438,N_6326,N_7405);
nor U10439 (N_10439,N_5255,N_5843);
and U10440 (N_10440,N_6983,N_7556);
or U10441 (N_10441,N_5745,N_5646);
or U10442 (N_10442,N_4882,N_6352);
and U10443 (N_10443,N_5279,N_4001);
nand U10444 (N_10444,N_7027,N_7786);
nand U10445 (N_10445,N_5441,N_6164);
nand U10446 (N_10446,N_5746,N_6712);
xor U10447 (N_10447,N_6839,N_6289);
nor U10448 (N_10448,N_6275,N_5817);
nand U10449 (N_10449,N_4598,N_7113);
xnor U10450 (N_10450,N_5163,N_7848);
or U10451 (N_10451,N_7288,N_4971);
or U10452 (N_10452,N_5233,N_7787);
and U10453 (N_10453,N_4090,N_5410);
nor U10454 (N_10454,N_6194,N_4882);
or U10455 (N_10455,N_5759,N_6630);
nand U10456 (N_10456,N_4314,N_7108);
nor U10457 (N_10457,N_7172,N_4685);
and U10458 (N_10458,N_7034,N_5602);
nand U10459 (N_10459,N_4166,N_7107);
nand U10460 (N_10460,N_7066,N_6128);
and U10461 (N_10461,N_6241,N_6735);
nor U10462 (N_10462,N_7112,N_5975);
nor U10463 (N_10463,N_5308,N_4915);
nor U10464 (N_10464,N_6812,N_4158);
nand U10465 (N_10465,N_6569,N_7007);
nor U10466 (N_10466,N_5941,N_7192);
nand U10467 (N_10467,N_5934,N_5004);
nor U10468 (N_10468,N_5676,N_6964);
and U10469 (N_10469,N_6571,N_7406);
or U10470 (N_10470,N_6499,N_6914);
or U10471 (N_10471,N_6695,N_4911);
and U10472 (N_10472,N_6395,N_5337);
and U10473 (N_10473,N_5268,N_6862);
xor U10474 (N_10474,N_5714,N_6704);
nor U10475 (N_10475,N_7206,N_5622);
and U10476 (N_10476,N_6545,N_5196);
nor U10477 (N_10477,N_5902,N_4965);
nand U10478 (N_10478,N_6600,N_7774);
or U10479 (N_10479,N_6040,N_6360);
or U10480 (N_10480,N_4216,N_4455);
or U10481 (N_10481,N_6033,N_5991);
nand U10482 (N_10482,N_7261,N_7259);
and U10483 (N_10483,N_7497,N_5211);
and U10484 (N_10484,N_5707,N_5060);
nand U10485 (N_10485,N_5084,N_4291);
and U10486 (N_10486,N_5871,N_7201);
or U10487 (N_10487,N_7302,N_4450);
and U10488 (N_10488,N_6555,N_5273);
or U10489 (N_10489,N_5966,N_6842);
and U10490 (N_10490,N_4389,N_4868);
nor U10491 (N_10491,N_4317,N_4051);
or U10492 (N_10492,N_6332,N_5894);
nor U10493 (N_10493,N_7492,N_7115);
nand U10494 (N_10494,N_4354,N_5057);
nor U10495 (N_10495,N_7026,N_5507);
nor U10496 (N_10496,N_5216,N_6602);
nor U10497 (N_10497,N_6635,N_5179);
and U10498 (N_10498,N_7616,N_4557);
xor U10499 (N_10499,N_6352,N_5179);
xnor U10500 (N_10500,N_6471,N_6541);
nor U10501 (N_10501,N_4694,N_5307);
or U10502 (N_10502,N_6354,N_7451);
or U10503 (N_10503,N_6777,N_6998);
nand U10504 (N_10504,N_4041,N_5974);
nand U10505 (N_10505,N_6286,N_4640);
nor U10506 (N_10506,N_7381,N_5179);
nor U10507 (N_10507,N_6961,N_7704);
nand U10508 (N_10508,N_4207,N_6486);
and U10509 (N_10509,N_5420,N_7994);
or U10510 (N_10510,N_5796,N_7615);
or U10511 (N_10511,N_4565,N_6543);
and U10512 (N_10512,N_4157,N_7356);
nor U10513 (N_10513,N_6277,N_4244);
or U10514 (N_10514,N_7356,N_6662);
and U10515 (N_10515,N_4715,N_7386);
xor U10516 (N_10516,N_5165,N_5906);
or U10517 (N_10517,N_6235,N_7786);
nand U10518 (N_10518,N_6180,N_4303);
and U10519 (N_10519,N_7597,N_7968);
and U10520 (N_10520,N_5696,N_7803);
nor U10521 (N_10521,N_4218,N_5771);
or U10522 (N_10522,N_4658,N_7640);
and U10523 (N_10523,N_7778,N_6454);
nor U10524 (N_10524,N_5664,N_7088);
nor U10525 (N_10525,N_6444,N_7346);
or U10526 (N_10526,N_5448,N_4412);
nor U10527 (N_10527,N_4410,N_4028);
xnor U10528 (N_10528,N_5075,N_7409);
nor U10529 (N_10529,N_6688,N_7151);
nor U10530 (N_10530,N_7457,N_5123);
xnor U10531 (N_10531,N_6127,N_6692);
or U10532 (N_10532,N_5411,N_6491);
nor U10533 (N_10533,N_7250,N_7294);
xor U10534 (N_10534,N_4067,N_6026);
and U10535 (N_10535,N_4507,N_6131);
nand U10536 (N_10536,N_7748,N_6990);
nand U10537 (N_10537,N_4809,N_5512);
or U10538 (N_10538,N_5247,N_4847);
xnor U10539 (N_10539,N_6799,N_5947);
or U10540 (N_10540,N_6116,N_5918);
nor U10541 (N_10541,N_7012,N_6650);
nor U10542 (N_10542,N_5467,N_5460);
or U10543 (N_10543,N_7480,N_6520);
nor U10544 (N_10544,N_7273,N_7719);
or U10545 (N_10545,N_7606,N_7281);
and U10546 (N_10546,N_4448,N_7089);
nand U10547 (N_10547,N_5859,N_6540);
or U10548 (N_10548,N_7562,N_6031);
and U10549 (N_10549,N_5532,N_5090);
nor U10550 (N_10550,N_7136,N_7409);
xnor U10551 (N_10551,N_7505,N_4703);
nand U10552 (N_10552,N_4996,N_4235);
nand U10553 (N_10553,N_5419,N_4396);
or U10554 (N_10554,N_5887,N_7799);
nor U10555 (N_10555,N_7829,N_4661);
or U10556 (N_10556,N_7585,N_6122);
nor U10557 (N_10557,N_5928,N_7018);
nor U10558 (N_10558,N_5975,N_4138);
nor U10559 (N_10559,N_6274,N_4918);
and U10560 (N_10560,N_7504,N_4109);
xnor U10561 (N_10561,N_4115,N_4866);
nand U10562 (N_10562,N_6676,N_5903);
nand U10563 (N_10563,N_5486,N_4870);
nor U10564 (N_10564,N_4822,N_5974);
nand U10565 (N_10565,N_7700,N_5977);
or U10566 (N_10566,N_4306,N_7610);
nand U10567 (N_10567,N_5990,N_7818);
or U10568 (N_10568,N_5718,N_5941);
nor U10569 (N_10569,N_6232,N_6140);
nand U10570 (N_10570,N_5804,N_4064);
and U10571 (N_10571,N_4068,N_6472);
xor U10572 (N_10572,N_7415,N_5464);
and U10573 (N_10573,N_6415,N_7595);
and U10574 (N_10574,N_6456,N_5101);
and U10575 (N_10575,N_6481,N_6715);
xnor U10576 (N_10576,N_7171,N_4841);
xor U10577 (N_10577,N_7196,N_4816);
xor U10578 (N_10578,N_7570,N_4500);
or U10579 (N_10579,N_6929,N_4362);
and U10580 (N_10580,N_4017,N_6639);
nor U10581 (N_10581,N_6104,N_6970);
and U10582 (N_10582,N_4790,N_6671);
nand U10583 (N_10583,N_5182,N_7825);
nor U10584 (N_10584,N_4608,N_7652);
nand U10585 (N_10585,N_6178,N_7375);
nor U10586 (N_10586,N_5514,N_7081);
nor U10587 (N_10587,N_7558,N_5458);
nand U10588 (N_10588,N_6446,N_6682);
xor U10589 (N_10589,N_7348,N_7865);
nand U10590 (N_10590,N_4395,N_6927);
xnor U10591 (N_10591,N_6685,N_7333);
and U10592 (N_10592,N_4685,N_5845);
and U10593 (N_10593,N_5783,N_6601);
and U10594 (N_10594,N_6854,N_7242);
and U10595 (N_10595,N_4946,N_7292);
or U10596 (N_10596,N_6732,N_4226);
nand U10597 (N_10597,N_6696,N_5215);
and U10598 (N_10598,N_7926,N_7360);
nand U10599 (N_10599,N_5167,N_4032);
xor U10600 (N_10600,N_4915,N_6518);
or U10601 (N_10601,N_7462,N_4131);
and U10602 (N_10602,N_5897,N_4902);
nand U10603 (N_10603,N_6670,N_6086);
and U10604 (N_10604,N_7306,N_6520);
nand U10605 (N_10605,N_5549,N_4378);
or U10606 (N_10606,N_7631,N_5423);
nand U10607 (N_10607,N_5570,N_4241);
nand U10608 (N_10608,N_6043,N_7906);
or U10609 (N_10609,N_6932,N_6497);
nor U10610 (N_10610,N_7902,N_7925);
nand U10611 (N_10611,N_7935,N_5107);
or U10612 (N_10612,N_6515,N_5738);
or U10613 (N_10613,N_5461,N_7420);
xnor U10614 (N_10614,N_5046,N_4798);
and U10615 (N_10615,N_7918,N_5074);
and U10616 (N_10616,N_4671,N_6123);
nor U10617 (N_10617,N_6663,N_6498);
nand U10618 (N_10618,N_6129,N_7018);
and U10619 (N_10619,N_5430,N_4683);
nor U10620 (N_10620,N_5429,N_7335);
and U10621 (N_10621,N_6314,N_7437);
nand U10622 (N_10622,N_7605,N_7613);
and U10623 (N_10623,N_5014,N_7345);
nor U10624 (N_10624,N_7456,N_4066);
nand U10625 (N_10625,N_4788,N_6372);
xor U10626 (N_10626,N_6446,N_6861);
or U10627 (N_10627,N_5050,N_4144);
and U10628 (N_10628,N_5873,N_5023);
nand U10629 (N_10629,N_5500,N_5580);
or U10630 (N_10630,N_5946,N_5844);
nor U10631 (N_10631,N_6814,N_7176);
xor U10632 (N_10632,N_6719,N_6360);
xor U10633 (N_10633,N_6960,N_5238);
and U10634 (N_10634,N_6157,N_6593);
nand U10635 (N_10635,N_4866,N_7450);
nor U10636 (N_10636,N_7695,N_6530);
and U10637 (N_10637,N_4584,N_4823);
and U10638 (N_10638,N_6644,N_7170);
and U10639 (N_10639,N_4572,N_7668);
or U10640 (N_10640,N_4810,N_5955);
nand U10641 (N_10641,N_5983,N_4036);
xor U10642 (N_10642,N_4758,N_6390);
and U10643 (N_10643,N_5082,N_4955);
and U10644 (N_10644,N_4345,N_6503);
nor U10645 (N_10645,N_4494,N_4877);
nand U10646 (N_10646,N_4943,N_5468);
xnor U10647 (N_10647,N_5787,N_6283);
xnor U10648 (N_10648,N_5485,N_4031);
or U10649 (N_10649,N_4991,N_7625);
or U10650 (N_10650,N_7043,N_7515);
nand U10651 (N_10651,N_7066,N_5724);
or U10652 (N_10652,N_7267,N_4582);
nand U10653 (N_10653,N_5648,N_5335);
nor U10654 (N_10654,N_4573,N_4058);
nand U10655 (N_10655,N_5950,N_4747);
xnor U10656 (N_10656,N_5970,N_7663);
nand U10657 (N_10657,N_6674,N_4347);
nor U10658 (N_10658,N_4144,N_5478);
or U10659 (N_10659,N_6756,N_4548);
nand U10660 (N_10660,N_4471,N_6561);
or U10661 (N_10661,N_4290,N_6693);
and U10662 (N_10662,N_5191,N_7296);
or U10663 (N_10663,N_5175,N_6254);
nand U10664 (N_10664,N_7329,N_6547);
nand U10665 (N_10665,N_4159,N_5226);
nor U10666 (N_10666,N_7192,N_6345);
nand U10667 (N_10667,N_6454,N_4689);
nand U10668 (N_10668,N_6910,N_7060);
or U10669 (N_10669,N_5595,N_4574);
nand U10670 (N_10670,N_6846,N_5052);
or U10671 (N_10671,N_4861,N_7305);
or U10672 (N_10672,N_5493,N_5806);
and U10673 (N_10673,N_4850,N_6754);
nor U10674 (N_10674,N_7905,N_7390);
nand U10675 (N_10675,N_6430,N_4323);
nand U10676 (N_10676,N_7139,N_4049);
nor U10677 (N_10677,N_5872,N_6732);
nand U10678 (N_10678,N_4351,N_6340);
and U10679 (N_10679,N_4568,N_5256);
and U10680 (N_10680,N_5306,N_5822);
or U10681 (N_10681,N_4455,N_4117);
and U10682 (N_10682,N_7897,N_6666);
or U10683 (N_10683,N_6061,N_7698);
or U10684 (N_10684,N_7291,N_7875);
xnor U10685 (N_10685,N_4623,N_5914);
nand U10686 (N_10686,N_4785,N_4549);
nor U10687 (N_10687,N_6755,N_4560);
and U10688 (N_10688,N_5655,N_7304);
or U10689 (N_10689,N_5720,N_7974);
or U10690 (N_10690,N_5286,N_4670);
nor U10691 (N_10691,N_7682,N_5999);
xor U10692 (N_10692,N_6932,N_6282);
nand U10693 (N_10693,N_5675,N_6699);
nor U10694 (N_10694,N_6136,N_7120);
nand U10695 (N_10695,N_5107,N_4783);
and U10696 (N_10696,N_4858,N_4716);
nand U10697 (N_10697,N_7943,N_7550);
or U10698 (N_10698,N_7687,N_7686);
xor U10699 (N_10699,N_7088,N_7274);
and U10700 (N_10700,N_7127,N_5859);
nor U10701 (N_10701,N_7240,N_7048);
or U10702 (N_10702,N_6183,N_5040);
nand U10703 (N_10703,N_7632,N_6478);
nand U10704 (N_10704,N_4291,N_7008);
or U10705 (N_10705,N_6462,N_7375);
xnor U10706 (N_10706,N_5753,N_7382);
nor U10707 (N_10707,N_4493,N_5480);
and U10708 (N_10708,N_4787,N_5262);
nand U10709 (N_10709,N_6692,N_4416);
and U10710 (N_10710,N_6104,N_7929);
and U10711 (N_10711,N_4003,N_4890);
nor U10712 (N_10712,N_4813,N_6781);
nor U10713 (N_10713,N_4504,N_7082);
nand U10714 (N_10714,N_4784,N_7991);
or U10715 (N_10715,N_4958,N_6647);
nand U10716 (N_10716,N_5583,N_7672);
nor U10717 (N_10717,N_4990,N_5797);
xor U10718 (N_10718,N_6805,N_4739);
and U10719 (N_10719,N_5141,N_5235);
xnor U10720 (N_10720,N_5639,N_7802);
or U10721 (N_10721,N_5411,N_5682);
nor U10722 (N_10722,N_7799,N_4709);
or U10723 (N_10723,N_5860,N_5368);
nand U10724 (N_10724,N_6293,N_6414);
nand U10725 (N_10725,N_5167,N_7573);
or U10726 (N_10726,N_7174,N_6508);
nor U10727 (N_10727,N_5179,N_6996);
nor U10728 (N_10728,N_4540,N_4307);
nand U10729 (N_10729,N_5625,N_5323);
and U10730 (N_10730,N_6748,N_6359);
and U10731 (N_10731,N_6356,N_6754);
nand U10732 (N_10732,N_7218,N_5529);
or U10733 (N_10733,N_5190,N_6162);
nor U10734 (N_10734,N_4861,N_5452);
nand U10735 (N_10735,N_7488,N_5867);
nor U10736 (N_10736,N_7515,N_6463);
or U10737 (N_10737,N_5188,N_4333);
nor U10738 (N_10738,N_5359,N_5826);
nor U10739 (N_10739,N_4045,N_7797);
nor U10740 (N_10740,N_4771,N_5213);
and U10741 (N_10741,N_6765,N_7820);
or U10742 (N_10742,N_4087,N_5444);
and U10743 (N_10743,N_7688,N_6279);
nor U10744 (N_10744,N_6245,N_7384);
xor U10745 (N_10745,N_7487,N_5218);
and U10746 (N_10746,N_6786,N_6834);
nand U10747 (N_10747,N_7948,N_5328);
or U10748 (N_10748,N_7983,N_5806);
nor U10749 (N_10749,N_6181,N_4029);
and U10750 (N_10750,N_6605,N_6950);
nand U10751 (N_10751,N_7440,N_5951);
or U10752 (N_10752,N_6640,N_5074);
nand U10753 (N_10753,N_4978,N_6288);
nand U10754 (N_10754,N_5418,N_6938);
and U10755 (N_10755,N_7156,N_4799);
and U10756 (N_10756,N_5738,N_4741);
and U10757 (N_10757,N_4650,N_4767);
nand U10758 (N_10758,N_4522,N_7654);
nor U10759 (N_10759,N_4095,N_7437);
and U10760 (N_10760,N_4752,N_5385);
nand U10761 (N_10761,N_7586,N_4903);
nor U10762 (N_10762,N_5204,N_5632);
nand U10763 (N_10763,N_4186,N_5154);
and U10764 (N_10764,N_6449,N_6861);
or U10765 (N_10765,N_4705,N_4457);
nor U10766 (N_10766,N_6593,N_5203);
nor U10767 (N_10767,N_7377,N_5972);
or U10768 (N_10768,N_5114,N_5051);
nand U10769 (N_10769,N_6864,N_7765);
xor U10770 (N_10770,N_7877,N_5069);
nor U10771 (N_10771,N_4154,N_5364);
nand U10772 (N_10772,N_7580,N_5796);
or U10773 (N_10773,N_7794,N_5930);
nor U10774 (N_10774,N_4796,N_4649);
xor U10775 (N_10775,N_6451,N_4153);
or U10776 (N_10776,N_4538,N_7105);
nor U10777 (N_10777,N_4000,N_6375);
xnor U10778 (N_10778,N_5550,N_7625);
nor U10779 (N_10779,N_5336,N_6075);
or U10780 (N_10780,N_5204,N_4439);
nor U10781 (N_10781,N_5425,N_5128);
and U10782 (N_10782,N_4260,N_4057);
nand U10783 (N_10783,N_6714,N_5550);
and U10784 (N_10784,N_7797,N_6335);
nand U10785 (N_10785,N_6295,N_5720);
nand U10786 (N_10786,N_7420,N_7157);
or U10787 (N_10787,N_5240,N_4677);
nand U10788 (N_10788,N_4572,N_6108);
nand U10789 (N_10789,N_4068,N_7358);
or U10790 (N_10790,N_7416,N_5866);
or U10791 (N_10791,N_7555,N_7114);
and U10792 (N_10792,N_5300,N_7428);
nand U10793 (N_10793,N_7462,N_6978);
or U10794 (N_10794,N_6049,N_4659);
nor U10795 (N_10795,N_5075,N_7335);
nor U10796 (N_10796,N_5895,N_7233);
nand U10797 (N_10797,N_7521,N_7436);
nand U10798 (N_10798,N_5269,N_7278);
nor U10799 (N_10799,N_6803,N_6807);
xnor U10800 (N_10800,N_7504,N_5663);
and U10801 (N_10801,N_7590,N_6061);
nand U10802 (N_10802,N_4253,N_4709);
xor U10803 (N_10803,N_7726,N_5377);
or U10804 (N_10804,N_5915,N_5238);
or U10805 (N_10805,N_6321,N_5749);
and U10806 (N_10806,N_7908,N_4340);
and U10807 (N_10807,N_4643,N_4779);
and U10808 (N_10808,N_5703,N_4199);
and U10809 (N_10809,N_4487,N_6361);
nor U10810 (N_10810,N_4587,N_5095);
nor U10811 (N_10811,N_4840,N_6372);
or U10812 (N_10812,N_7005,N_6815);
nand U10813 (N_10813,N_6490,N_6840);
nor U10814 (N_10814,N_7106,N_7978);
or U10815 (N_10815,N_6942,N_4645);
and U10816 (N_10816,N_7597,N_7937);
or U10817 (N_10817,N_5427,N_5368);
and U10818 (N_10818,N_6406,N_5189);
nor U10819 (N_10819,N_7671,N_4905);
xor U10820 (N_10820,N_4136,N_4798);
nand U10821 (N_10821,N_4756,N_5842);
or U10822 (N_10822,N_5764,N_7284);
and U10823 (N_10823,N_5312,N_7462);
nor U10824 (N_10824,N_4718,N_6941);
nand U10825 (N_10825,N_5281,N_5666);
nand U10826 (N_10826,N_7430,N_4718);
nand U10827 (N_10827,N_6612,N_7226);
nand U10828 (N_10828,N_4025,N_6781);
nand U10829 (N_10829,N_7308,N_6554);
nor U10830 (N_10830,N_7804,N_6565);
nor U10831 (N_10831,N_5327,N_4011);
nor U10832 (N_10832,N_7691,N_6893);
or U10833 (N_10833,N_4257,N_4114);
or U10834 (N_10834,N_4003,N_7990);
and U10835 (N_10835,N_6658,N_5513);
nand U10836 (N_10836,N_5475,N_4073);
nand U10837 (N_10837,N_7517,N_7529);
xnor U10838 (N_10838,N_5091,N_7330);
nand U10839 (N_10839,N_7877,N_7676);
or U10840 (N_10840,N_6774,N_6768);
xor U10841 (N_10841,N_5112,N_4237);
nand U10842 (N_10842,N_4712,N_7957);
nor U10843 (N_10843,N_4207,N_7633);
or U10844 (N_10844,N_7377,N_7646);
nand U10845 (N_10845,N_7497,N_6312);
or U10846 (N_10846,N_7802,N_5181);
nor U10847 (N_10847,N_6140,N_7406);
nor U10848 (N_10848,N_5072,N_7229);
nor U10849 (N_10849,N_5855,N_5882);
xor U10850 (N_10850,N_5749,N_4349);
nand U10851 (N_10851,N_4506,N_6577);
or U10852 (N_10852,N_7569,N_4029);
or U10853 (N_10853,N_6531,N_4808);
nor U10854 (N_10854,N_4927,N_4474);
nor U10855 (N_10855,N_4236,N_4478);
nor U10856 (N_10856,N_5259,N_6010);
nor U10857 (N_10857,N_4834,N_5660);
nor U10858 (N_10858,N_7807,N_5967);
and U10859 (N_10859,N_7523,N_4737);
nand U10860 (N_10860,N_7198,N_5776);
nand U10861 (N_10861,N_4173,N_5755);
or U10862 (N_10862,N_5601,N_5115);
or U10863 (N_10863,N_5508,N_7653);
nand U10864 (N_10864,N_6807,N_4598);
and U10865 (N_10865,N_5141,N_5937);
nor U10866 (N_10866,N_7117,N_7795);
and U10867 (N_10867,N_5668,N_5107);
nand U10868 (N_10868,N_6157,N_4575);
and U10869 (N_10869,N_4034,N_7660);
nor U10870 (N_10870,N_5511,N_7593);
nor U10871 (N_10871,N_7537,N_4161);
nor U10872 (N_10872,N_6947,N_5740);
or U10873 (N_10873,N_6712,N_6979);
nand U10874 (N_10874,N_6400,N_6158);
and U10875 (N_10875,N_6682,N_6723);
nand U10876 (N_10876,N_7118,N_7712);
and U10877 (N_10877,N_5079,N_5893);
nand U10878 (N_10878,N_7047,N_4062);
nor U10879 (N_10879,N_7623,N_4106);
nand U10880 (N_10880,N_4215,N_7659);
and U10881 (N_10881,N_5288,N_6372);
nand U10882 (N_10882,N_4643,N_6728);
or U10883 (N_10883,N_4234,N_4139);
and U10884 (N_10884,N_4076,N_6186);
xnor U10885 (N_10885,N_5056,N_7107);
xnor U10886 (N_10886,N_6097,N_4874);
and U10887 (N_10887,N_7254,N_4813);
nand U10888 (N_10888,N_6187,N_5363);
nor U10889 (N_10889,N_7185,N_4441);
and U10890 (N_10890,N_6208,N_7826);
or U10891 (N_10891,N_7714,N_6162);
nand U10892 (N_10892,N_7361,N_4077);
and U10893 (N_10893,N_6484,N_4019);
nor U10894 (N_10894,N_4382,N_5790);
and U10895 (N_10895,N_6534,N_7441);
or U10896 (N_10896,N_6967,N_5575);
and U10897 (N_10897,N_4045,N_7720);
and U10898 (N_10898,N_7435,N_5313);
xor U10899 (N_10899,N_4310,N_6715);
or U10900 (N_10900,N_6187,N_6623);
and U10901 (N_10901,N_7007,N_7174);
and U10902 (N_10902,N_7168,N_4096);
nand U10903 (N_10903,N_6617,N_5293);
nand U10904 (N_10904,N_6908,N_4035);
nand U10905 (N_10905,N_7175,N_7677);
nor U10906 (N_10906,N_6107,N_7475);
or U10907 (N_10907,N_5428,N_5086);
nor U10908 (N_10908,N_4783,N_7639);
nand U10909 (N_10909,N_4212,N_6221);
and U10910 (N_10910,N_4227,N_5549);
nor U10911 (N_10911,N_6642,N_5141);
and U10912 (N_10912,N_4866,N_5946);
or U10913 (N_10913,N_7644,N_5619);
or U10914 (N_10914,N_6543,N_6488);
nor U10915 (N_10915,N_5697,N_6179);
nor U10916 (N_10916,N_7034,N_5577);
and U10917 (N_10917,N_5145,N_7969);
or U10918 (N_10918,N_5294,N_5044);
and U10919 (N_10919,N_7197,N_5677);
nor U10920 (N_10920,N_6511,N_6840);
and U10921 (N_10921,N_6963,N_6823);
nand U10922 (N_10922,N_6551,N_5981);
nor U10923 (N_10923,N_5482,N_6014);
and U10924 (N_10924,N_4461,N_5047);
or U10925 (N_10925,N_4988,N_6537);
nor U10926 (N_10926,N_7854,N_4199);
and U10927 (N_10927,N_4104,N_4678);
and U10928 (N_10928,N_4371,N_5700);
or U10929 (N_10929,N_4349,N_7988);
and U10930 (N_10930,N_6847,N_4520);
nand U10931 (N_10931,N_6554,N_5584);
nor U10932 (N_10932,N_5232,N_7246);
and U10933 (N_10933,N_6164,N_6785);
and U10934 (N_10934,N_7642,N_6782);
or U10935 (N_10935,N_4489,N_7782);
xor U10936 (N_10936,N_7346,N_7349);
nand U10937 (N_10937,N_4645,N_7353);
nand U10938 (N_10938,N_7290,N_6768);
nand U10939 (N_10939,N_7367,N_4951);
nand U10940 (N_10940,N_6118,N_6819);
or U10941 (N_10941,N_7941,N_5289);
xnor U10942 (N_10942,N_5657,N_5790);
and U10943 (N_10943,N_5225,N_5517);
and U10944 (N_10944,N_7154,N_4246);
or U10945 (N_10945,N_5576,N_4464);
or U10946 (N_10946,N_7425,N_7150);
nor U10947 (N_10947,N_5713,N_4813);
xnor U10948 (N_10948,N_7693,N_7064);
nor U10949 (N_10949,N_5030,N_6809);
nor U10950 (N_10950,N_4655,N_5084);
nand U10951 (N_10951,N_6726,N_7407);
nand U10952 (N_10952,N_7232,N_6736);
or U10953 (N_10953,N_4325,N_5221);
or U10954 (N_10954,N_6049,N_5004);
or U10955 (N_10955,N_6703,N_6584);
nand U10956 (N_10956,N_4777,N_5750);
or U10957 (N_10957,N_5295,N_5140);
and U10958 (N_10958,N_7882,N_5992);
and U10959 (N_10959,N_5299,N_5137);
and U10960 (N_10960,N_7679,N_5585);
nand U10961 (N_10961,N_5986,N_6688);
or U10962 (N_10962,N_7290,N_4718);
xnor U10963 (N_10963,N_4425,N_7715);
or U10964 (N_10964,N_5189,N_7209);
and U10965 (N_10965,N_5469,N_4379);
and U10966 (N_10966,N_5813,N_5973);
nand U10967 (N_10967,N_4213,N_7682);
and U10968 (N_10968,N_4656,N_4293);
xnor U10969 (N_10969,N_7614,N_7616);
and U10970 (N_10970,N_6749,N_4160);
or U10971 (N_10971,N_5399,N_6023);
nand U10972 (N_10972,N_5297,N_4661);
nor U10973 (N_10973,N_5124,N_5623);
and U10974 (N_10974,N_5271,N_5375);
or U10975 (N_10975,N_7519,N_4446);
and U10976 (N_10976,N_7663,N_5070);
nand U10977 (N_10977,N_7147,N_7644);
xor U10978 (N_10978,N_7884,N_4248);
and U10979 (N_10979,N_5034,N_4640);
nor U10980 (N_10980,N_4145,N_6188);
or U10981 (N_10981,N_4454,N_7793);
or U10982 (N_10982,N_7809,N_5594);
nor U10983 (N_10983,N_6114,N_5666);
nor U10984 (N_10984,N_4161,N_7128);
nand U10985 (N_10985,N_6913,N_5720);
nor U10986 (N_10986,N_5348,N_5613);
nor U10987 (N_10987,N_4429,N_6829);
nor U10988 (N_10988,N_4265,N_5128);
nor U10989 (N_10989,N_7885,N_4644);
nand U10990 (N_10990,N_4361,N_7816);
nor U10991 (N_10991,N_4303,N_6108);
and U10992 (N_10992,N_7381,N_6802);
and U10993 (N_10993,N_5029,N_6768);
and U10994 (N_10994,N_4289,N_4624);
or U10995 (N_10995,N_6607,N_6533);
and U10996 (N_10996,N_6240,N_7604);
nand U10997 (N_10997,N_6093,N_6881);
nor U10998 (N_10998,N_7299,N_5851);
nand U10999 (N_10999,N_5605,N_5539);
and U11000 (N_11000,N_7429,N_6202);
xnor U11001 (N_11001,N_4613,N_4002);
xor U11002 (N_11002,N_6701,N_5849);
or U11003 (N_11003,N_7030,N_4392);
nor U11004 (N_11004,N_7093,N_5353);
or U11005 (N_11005,N_4489,N_7038);
nor U11006 (N_11006,N_5844,N_6746);
nand U11007 (N_11007,N_5995,N_4873);
nor U11008 (N_11008,N_6436,N_5127);
and U11009 (N_11009,N_4627,N_7182);
nor U11010 (N_11010,N_4321,N_7831);
nor U11011 (N_11011,N_4436,N_6762);
nor U11012 (N_11012,N_4510,N_5211);
nand U11013 (N_11013,N_6543,N_7026);
nand U11014 (N_11014,N_6879,N_5283);
or U11015 (N_11015,N_4868,N_7558);
nand U11016 (N_11016,N_5954,N_5720);
and U11017 (N_11017,N_7671,N_5405);
nand U11018 (N_11018,N_6027,N_6911);
or U11019 (N_11019,N_5207,N_6396);
xnor U11020 (N_11020,N_4233,N_4734);
nand U11021 (N_11021,N_5624,N_7607);
nand U11022 (N_11022,N_5708,N_7446);
xor U11023 (N_11023,N_4245,N_4737);
or U11024 (N_11024,N_5387,N_4012);
or U11025 (N_11025,N_7038,N_4465);
and U11026 (N_11026,N_4645,N_6546);
nor U11027 (N_11027,N_5228,N_5892);
nor U11028 (N_11028,N_4114,N_7468);
and U11029 (N_11029,N_4749,N_7853);
and U11030 (N_11030,N_4081,N_4946);
xor U11031 (N_11031,N_4371,N_6145);
nand U11032 (N_11032,N_7501,N_7282);
and U11033 (N_11033,N_4645,N_5591);
and U11034 (N_11034,N_5643,N_4763);
and U11035 (N_11035,N_5689,N_7105);
nand U11036 (N_11036,N_6307,N_5306);
or U11037 (N_11037,N_4176,N_7886);
nor U11038 (N_11038,N_5883,N_4514);
or U11039 (N_11039,N_7444,N_4517);
nor U11040 (N_11040,N_5579,N_5825);
nand U11041 (N_11041,N_5077,N_4920);
and U11042 (N_11042,N_6247,N_6329);
and U11043 (N_11043,N_5725,N_5211);
xor U11044 (N_11044,N_5094,N_7570);
nor U11045 (N_11045,N_5567,N_6479);
and U11046 (N_11046,N_4579,N_7975);
nand U11047 (N_11047,N_6717,N_5269);
nor U11048 (N_11048,N_6156,N_5854);
or U11049 (N_11049,N_6172,N_5725);
nand U11050 (N_11050,N_6817,N_7173);
or U11051 (N_11051,N_5299,N_4066);
and U11052 (N_11052,N_7452,N_4345);
nor U11053 (N_11053,N_4300,N_5320);
nand U11054 (N_11054,N_4030,N_5559);
and U11055 (N_11055,N_4928,N_4131);
nand U11056 (N_11056,N_7055,N_5597);
nor U11057 (N_11057,N_5208,N_4672);
and U11058 (N_11058,N_4145,N_7872);
nand U11059 (N_11059,N_4274,N_6775);
or U11060 (N_11060,N_7630,N_4240);
nand U11061 (N_11061,N_7501,N_4792);
nor U11062 (N_11062,N_7618,N_4166);
xnor U11063 (N_11063,N_7842,N_7989);
and U11064 (N_11064,N_4518,N_4218);
and U11065 (N_11065,N_4374,N_5414);
and U11066 (N_11066,N_6403,N_4242);
or U11067 (N_11067,N_6132,N_5093);
and U11068 (N_11068,N_7416,N_7342);
and U11069 (N_11069,N_4784,N_5038);
nor U11070 (N_11070,N_5977,N_4810);
nor U11071 (N_11071,N_7565,N_6375);
nand U11072 (N_11072,N_4572,N_5572);
or U11073 (N_11073,N_5416,N_6679);
or U11074 (N_11074,N_6099,N_6200);
or U11075 (N_11075,N_4519,N_7417);
and U11076 (N_11076,N_5246,N_5533);
xnor U11077 (N_11077,N_7606,N_5845);
xnor U11078 (N_11078,N_4986,N_6134);
xor U11079 (N_11079,N_5352,N_7080);
xnor U11080 (N_11080,N_7167,N_5493);
or U11081 (N_11081,N_4452,N_4309);
and U11082 (N_11082,N_5808,N_7328);
and U11083 (N_11083,N_7592,N_5535);
nor U11084 (N_11084,N_4998,N_4666);
nand U11085 (N_11085,N_7192,N_4573);
or U11086 (N_11086,N_5349,N_7527);
nand U11087 (N_11087,N_6117,N_7850);
xnor U11088 (N_11088,N_4912,N_4176);
nor U11089 (N_11089,N_7302,N_4504);
nand U11090 (N_11090,N_7476,N_7117);
and U11091 (N_11091,N_6398,N_6688);
and U11092 (N_11092,N_7737,N_6744);
and U11093 (N_11093,N_5578,N_4199);
and U11094 (N_11094,N_5789,N_5329);
nor U11095 (N_11095,N_5177,N_4948);
and U11096 (N_11096,N_4784,N_7193);
or U11097 (N_11097,N_7854,N_4635);
and U11098 (N_11098,N_4581,N_5895);
nand U11099 (N_11099,N_6791,N_6414);
nor U11100 (N_11100,N_6115,N_5613);
and U11101 (N_11101,N_7053,N_6025);
or U11102 (N_11102,N_7818,N_5700);
nor U11103 (N_11103,N_4355,N_4037);
or U11104 (N_11104,N_4024,N_4747);
xor U11105 (N_11105,N_5502,N_4743);
xnor U11106 (N_11106,N_7404,N_5041);
nand U11107 (N_11107,N_6653,N_5546);
or U11108 (N_11108,N_6874,N_5747);
xor U11109 (N_11109,N_4706,N_7248);
and U11110 (N_11110,N_7653,N_7386);
nand U11111 (N_11111,N_7785,N_7809);
nor U11112 (N_11112,N_7555,N_5494);
or U11113 (N_11113,N_6875,N_6610);
or U11114 (N_11114,N_4240,N_7271);
or U11115 (N_11115,N_4679,N_5544);
or U11116 (N_11116,N_7553,N_6619);
or U11117 (N_11117,N_4322,N_7497);
and U11118 (N_11118,N_5606,N_4190);
and U11119 (N_11119,N_5730,N_6736);
nor U11120 (N_11120,N_6116,N_5975);
or U11121 (N_11121,N_4853,N_6660);
or U11122 (N_11122,N_7800,N_6668);
and U11123 (N_11123,N_6044,N_7197);
nand U11124 (N_11124,N_7319,N_7155);
nand U11125 (N_11125,N_7218,N_4635);
nor U11126 (N_11126,N_5522,N_4131);
nor U11127 (N_11127,N_7318,N_4748);
and U11128 (N_11128,N_7865,N_6377);
xor U11129 (N_11129,N_4496,N_7606);
xnor U11130 (N_11130,N_5282,N_5324);
or U11131 (N_11131,N_7947,N_5077);
xor U11132 (N_11132,N_5505,N_4117);
or U11133 (N_11133,N_7978,N_6170);
xnor U11134 (N_11134,N_5960,N_5032);
xnor U11135 (N_11135,N_6244,N_7316);
xor U11136 (N_11136,N_5918,N_5786);
nor U11137 (N_11137,N_6422,N_5343);
nor U11138 (N_11138,N_5444,N_4854);
nor U11139 (N_11139,N_5125,N_7329);
nand U11140 (N_11140,N_5887,N_5478);
or U11141 (N_11141,N_5715,N_7114);
or U11142 (N_11142,N_4256,N_4692);
or U11143 (N_11143,N_6016,N_7709);
nor U11144 (N_11144,N_7349,N_5923);
nor U11145 (N_11145,N_6527,N_4846);
nand U11146 (N_11146,N_5656,N_6010);
or U11147 (N_11147,N_7323,N_4743);
nor U11148 (N_11148,N_6433,N_6184);
nor U11149 (N_11149,N_5493,N_4253);
and U11150 (N_11150,N_6518,N_6187);
nor U11151 (N_11151,N_4196,N_7164);
or U11152 (N_11152,N_6527,N_7941);
xor U11153 (N_11153,N_6086,N_7666);
and U11154 (N_11154,N_4007,N_5130);
xnor U11155 (N_11155,N_4989,N_4301);
and U11156 (N_11156,N_4329,N_5715);
nand U11157 (N_11157,N_7608,N_4384);
xor U11158 (N_11158,N_5991,N_5261);
or U11159 (N_11159,N_5005,N_5239);
nor U11160 (N_11160,N_5158,N_4013);
or U11161 (N_11161,N_4441,N_7551);
and U11162 (N_11162,N_4931,N_5369);
nor U11163 (N_11163,N_5677,N_7558);
nor U11164 (N_11164,N_4139,N_6223);
and U11165 (N_11165,N_7266,N_4689);
and U11166 (N_11166,N_6959,N_4588);
nor U11167 (N_11167,N_4999,N_7975);
nand U11168 (N_11168,N_5585,N_7535);
or U11169 (N_11169,N_4007,N_6942);
nor U11170 (N_11170,N_5338,N_4871);
nand U11171 (N_11171,N_4363,N_5386);
nor U11172 (N_11172,N_7867,N_4478);
and U11173 (N_11173,N_6220,N_5900);
or U11174 (N_11174,N_4173,N_4724);
nor U11175 (N_11175,N_4394,N_6209);
and U11176 (N_11176,N_4274,N_4736);
and U11177 (N_11177,N_7354,N_7003);
nand U11178 (N_11178,N_5608,N_7141);
or U11179 (N_11179,N_7126,N_4957);
or U11180 (N_11180,N_4320,N_6631);
nand U11181 (N_11181,N_4216,N_7111);
nor U11182 (N_11182,N_4370,N_5187);
nor U11183 (N_11183,N_5997,N_4560);
nand U11184 (N_11184,N_7173,N_5397);
nor U11185 (N_11185,N_7761,N_7308);
and U11186 (N_11186,N_6602,N_5823);
and U11187 (N_11187,N_7152,N_7935);
nor U11188 (N_11188,N_6476,N_5027);
nand U11189 (N_11189,N_6999,N_6811);
nand U11190 (N_11190,N_7122,N_5406);
and U11191 (N_11191,N_5191,N_7981);
nand U11192 (N_11192,N_4818,N_5126);
nand U11193 (N_11193,N_5897,N_4975);
nand U11194 (N_11194,N_4572,N_5613);
nand U11195 (N_11195,N_7305,N_6669);
and U11196 (N_11196,N_4689,N_4477);
nor U11197 (N_11197,N_6391,N_4287);
xnor U11198 (N_11198,N_6365,N_6048);
nand U11199 (N_11199,N_5621,N_6592);
xnor U11200 (N_11200,N_5936,N_7445);
or U11201 (N_11201,N_5719,N_4445);
xor U11202 (N_11202,N_6544,N_6860);
or U11203 (N_11203,N_6716,N_6321);
nand U11204 (N_11204,N_6506,N_7965);
nand U11205 (N_11205,N_4417,N_7055);
or U11206 (N_11206,N_5970,N_4979);
xor U11207 (N_11207,N_5206,N_4450);
and U11208 (N_11208,N_4464,N_4727);
nand U11209 (N_11209,N_7020,N_7904);
or U11210 (N_11210,N_4974,N_4581);
and U11211 (N_11211,N_7087,N_6345);
nand U11212 (N_11212,N_4432,N_7245);
and U11213 (N_11213,N_7849,N_7290);
and U11214 (N_11214,N_5163,N_4920);
nand U11215 (N_11215,N_7273,N_7912);
nand U11216 (N_11216,N_5492,N_6901);
xor U11217 (N_11217,N_4062,N_7430);
and U11218 (N_11218,N_6074,N_6457);
or U11219 (N_11219,N_6269,N_7601);
nor U11220 (N_11220,N_6979,N_5309);
or U11221 (N_11221,N_6901,N_6543);
or U11222 (N_11222,N_5080,N_5990);
or U11223 (N_11223,N_6488,N_4369);
or U11224 (N_11224,N_6556,N_6870);
or U11225 (N_11225,N_7634,N_5092);
and U11226 (N_11226,N_7520,N_7223);
xnor U11227 (N_11227,N_5862,N_5758);
nor U11228 (N_11228,N_4686,N_6521);
or U11229 (N_11229,N_4849,N_6976);
xor U11230 (N_11230,N_4540,N_5205);
nand U11231 (N_11231,N_4829,N_7889);
and U11232 (N_11232,N_5962,N_6304);
or U11233 (N_11233,N_7878,N_7605);
or U11234 (N_11234,N_4085,N_5983);
nand U11235 (N_11235,N_5383,N_5565);
nor U11236 (N_11236,N_5978,N_7174);
or U11237 (N_11237,N_6288,N_6854);
and U11238 (N_11238,N_7939,N_4504);
or U11239 (N_11239,N_7961,N_6363);
nand U11240 (N_11240,N_6234,N_5006);
xor U11241 (N_11241,N_4204,N_7757);
or U11242 (N_11242,N_5574,N_7703);
xor U11243 (N_11243,N_4170,N_4311);
and U11244 (N_11244,N_6514,N_5159);
and U11245 (N_11245,N_6701,N_7044);
and U11246 (N_11246,N_7885,N_7603);
nor U11247 (N_11247,N_6052,N_4689);
or U11248 (N_11248,N_4882,N_4973);
nand U11249 (N_11249,N_6215,N_6796);
nand U11250 (N_11250,N_4634,N_6707);
or U11251 (N_11251,N_6693,N_6011);
nor U11252 (N_11252,N_4443,N_7855);
nor U11253 (N_11253,N_7584,N_4721);
or U11254 (N_11254,N_4817,N_6341);
or U11255 (N_11255,N_7739,N_7265);
nor U11256 (N_11256,N_7044,N_5772);
xor U11257 (N_11257,N_7918,N_7219);
xor U11258 (N_11258,N_6127,N_6445);
and U11259 (N_11259,N_6128,N_6468);
and U11260 (N_11260,N_7028,N_7553);
or U11261 (N_11261,N_7741,N_5349);
or U11262 (N_11262,N_5275,N_5272);
nand U11263 (N_11263,N_4942,N_6318);
or U11264 (N_11264,N_6712,N_6498);
and U11265 (N_11265,N_4617,N_6695);
and U11266 (N_11266,N_5424,N_5825);
and U11267 (N_11267,N_4121,N_7745);
and U11268 (N_11268,N_6896,N_6240);
xor U11269 (N_11269,N_4259,N_7084);
nor U11270 (N_11270,N_4792,N_7003);
xor U11271 (N_11271,N_5924,N_6209);
nor U11272 (N_11272,N_5660,N_6130);
and U11273 (N_11273,N_5248,N_6483);
nor U11274 (N_11274,N_6733,N_6921);
and U11275 (N_11275,N_4445,N_4244);
or U11276 (N_11276,N_5460,N_7633);
nor U11277 (N_11277,N_4909,N_5785);
and U11278 (N_11278,N_4983,N_6392);
and U11279 (N_11279,N_7977,N_4473);
nor U11280 (N_11280,N_6499,N_7205);
or U11281 (N_11281,N_4681,N_6992);
nand U11282 (N_11282,N_5928,N_7068);
and U11283 (N_11283,N_7781,N_5371);
nand U11284 (N_11284,N_5438,N_4630);
nor U11285 (N_11285,N_4164,N_5756);
and U11286 (N_11286,N_6266,N_6852);
and U11287 (N_11287,N_4251,N_6961);
and U11288 (N_11288,N_4639,N_6664);
nand U11289 (N_11289,N_4151,N_4046);
nand U11290 (N_11290,N_6401,N_7859);
or U11291 (N_11291,N_4433,N_7299);
xor U11292 (N_11292,N_4262,N_5618);
nor U11293 (N_11293,N_6250,N_4038);
or U11294 (N_11294,N_6151,N_5550);
and U11295 (N_11295,N_5991,N_6866);
xor U11296 (N_11296,N_7008,N_4692);
nand U11297 (N_11297,N_5409,N_6281);
or U11298 (N_11298,N_7323,N_7470);
nand U11299 (N_11299,N_6999,N_5573);
and U11300 (N_11300,N_4453,N_6011);
or U11301 (N_11301,N_4754,N_6707);
or U11302 (N_11302,N_5788,N_7190);
and U11303 (N_11303,N_5588,N_6921);
nor U11304 (N_11304,N_4152,N_6765);
nand U11305 (N_11305,N_4754,N_6841);
and U11306 (N_11306,N_4233,N_7956);
nand U11307 (N_11307,N_7131,N_4378);
or U11308 (N_11308,N_6000,N_6291);
xor U11309 (N_11309,N_6239,N_6892);
and U11310 (N_11310,N_6178,N_4215);
and U11311 (N_11311,N_6265,N_6431);
nor U11312 (N_11312,N_7533,N_6325);
nor U11313 (N_11313,N_5299,N_5637);
and U11314 (N_11314,N_4366,N_7478);
xor U11315 (N_11315,N_7793,N_5705);
nor U11316 (N_11316,N_5426,N_4024);
nor U11317 (N_11317,N_5355,N_5771);
nand U11318 (N_11318,N_5126,N_7077);
or U11319 (N_11319,N_7717,N_4926);
or U11320 (N_11320,N_7120,N_5739);
or U11321 (N_11321,N_4150,N_4488);
or U11322 (N_11322,N_6523,N_7388);
or U11323 (N_11323,N_4446,N_6633);
or U11324 (N_11324,N_5081,N_7043);
and U11325 (N_11325,N_5331,N_5956);
and U11326 (N_11326,N_6100,N_4864);
nand U11327 (N_11327,N_4088,N_4918);
nor U11328 (N_11328,N_7541,N_6557);
nor U11329 (N_11329,N_7937,N_7399);
xnor U11330 (N_11330,N_5686,N_4257);
xor U11331 (N_11331,N_6534,N_4539);
nor U11332 (N_11332,N_7750,N_7662);
nand U11333 (N_11333,N_5484,N_5030);
or U11334 (N_11334,N_5571,N_7175);
nor U11335 (N_11335,N_7308,N_5563);
nand U11336 (N_11336,N_4916,N_4655);
nor U11337 (N_11337,N_5977,N_4982);
or U11338 (N_11338,N_6623,N_4199);
and U11339 (N_11339,N_7703,N_7015);
and U11340 (N_11340,N_7201,N_6344);
or U11341 (N_11341,N_4288,N_5680);
and U11342 (N_11342,N_6627,N_7702);
and U11343 (N_11343,N_7047,N_7423);
or U11344 (N_11344,N_6288,N_4305);
nor U11345 (N_11345,N_5483,N_7936);
nor U11346 (N_11346,N_7957,N_4496);
nand U11347 (N_11347,N_5798,N_7885);
and U11348 (N_11348,N_7273,N_5706);
xor U11349 (N_11349,N_4077,N_6548);
or U11350 (N_11350,N_5535,N_7288);
or U11351 (N_11351,N_4095,N_5340);
nand U11352 (N_11352,N_7148,N_7542);
xor U11353 (N_11353,N_4483,N_7268);
nor U11354 (N_11354,N_5476,N_4067);
nor U11355 (N_11355,N_5576,N_6857);
nand U11356 (N_11356,N_4008,N_6850);
xor U11357 (N_11357,N_6621,N_6263);
nand U11358 (N_11358,N_4095,N_6356);
nand U11359 (N_11359,N_6320,N_5719);
nand U11360 (N_11360,N_6570,N_7560);
nand U11361 (N_11361,N_4602,N_5496);
and U11362 (N_11362,N_6583,N_6984);
xor U11363 (N_11363,N_6766,N_7408);
xnor U11364 (N_11364,N_5757,N_6958);
and U11365 (N_11365,N_5951,N_4332);
nand U11366 (N_11366,N_6515,N_5437);
or U11367 (N_11367,N_4202,N_4275);
or U11368 (N_11368,N_5217,N_7327);
or U11369 (N_11369,N_5733,N_5100);
nand U11370 (N_11370,N_7283,N_5026);
nor U11371 (N_11371,N_4236,N_7438);
nor U11372 (N_11372,N_4350,N_7607);
and U11373 (N_11373,N_4441,N_6110);
and U11374 (N_11374,N_4669,N_7751);
or U11375 (N_11375,N_5339,N_7093);
and U11376 (N_11376,N_6369,N_6053);
nand U11377 (N_11377,N_5456,N_4019);
nor U11378 (N_11378,N_4909,N_5334);
nand U11379 (N_11379,N_4338,N_5675);
nor U11380 (N_11380,N_5570,N_4418);
and U11381 (N_11381,N_7290,N_4726);
and U11382 (N_11382,N_5204,N_4672);
or U11383 (N_11383,N_4240,N_4252);
or U11384 (N_11384,N_4347,N_7138);
and U11385 (N_11385,N_7630,N_7437);
or U11386 (N_11386,N_4655,N_4687);
and U11387 (N_11387,N_5357,N_7269);
nor U11388 (N_11388,N_4684,N_7421);
or U11389 (N_11389,N_5861,N_6110);
nor U11390 (N_11390,N_4288,N_4853);
nor U11391 (N_11391,N_7557,N_5714);
xor U11392 (N_11392,N_7288,N_5873);
xor U11393 (N_11393,N_7278,N_5179);
and U11394 (N_11394,N_7866,N_7935);
nor U11395 (N_11395,N_7833,N_5046);
nor U11396 (N_11396,N_4144,N_6878);
and U11397 (N_11397,N_4672,N_4769);
nand U11398 (N_11398,N_6050,N_5813);
and U11399 (N_11399,N_4656,N_7508);
or U11400 (N_11400,N_6991,N_6874);
xor U11401 (N_11401,N_7958,N_7002);
xor U11402 (N_11402,N_4543,N_7956);
nand U11403 (N_11403,N_6299,N_7757);
and U11404 (N_11404,N_6142,N_6501);
nor U11405 (N_11405,N_4634,N_4735);
nand U11406 (N_11406,N_4566,N_7458);
nand U11407 (N_11407,N_5029,N_5333);
nand U11408 (N_11408,N_7117,N_5966);
or U11409 (N_11409,N_5154,N_6922);
nor U11410 (N_11410,N_6141,N_7629);
and U11411 (N_11411,N_5458,N_5787);
or U11412 (N_11412,N_7055,N_7785);
nor U11413 (N_11413,N_5523,N_6210);
nor U11414 (N_11414,N_5445,N_4163);
and U11415 (N_11415,N_5775,N_6036);
and U11416 (N_11416,N_6427,N_5583);
or U11417 (N_11417,N_4002,N_4934);
nand U11418 (N_11418,N_4161,N_7148);
and U11419 (N_11419,N_5659,N_6273);
or U11420 (N_11420,N_4143,N_7942);
nor U11421 (N_11421,N_5194,N_7370);
or U11422 (N_11422,N_7940,N_5160);
nand U11423 (N_11423,N_5719,N_7511);
or U11424 (N_11424,N_4612,N_5698);
xor U11425 (N_11425,N_7196,N_7104);
and U11426 (N_11426,N_5232,N_7855);
nor U11427 (N_11427,N_5277,N_5482);
or U11428 (N_11428,N_7472,N_7150);
and U11429 (N_11429,N_4686,N_7148);
xor U11430 (N_11430,N_4332,N_7044);
nand U11431 (N_11431,N_7181,N_4165);
or U11432 (N_11432,N_7962,N_6522);
or U11433 (N_11433,N_6731,N_6344);
and U11434 (N_11434,N_7474,N_7289);
or U11435 (N_11435,N_4299,N_5568);
nor U11436 (N_11436,N_4901,N_7013);
xnor U11437 (N_11437,N_7352,N_7119);
nor U11438 (N_11438,N_6096,N_6013);
and U11439 (N_11439,N_5439,N_4690);
xor U11440 (N_11440,N_4455,N_5990);
or U11441 (N_11441,N_6425,N_4828);
nor U11442 (N_11442,N_6609,N_4655);
nand U11443 (N_11443,N_7244,N_7562);
xnor U11444 (N_11444,N_6450,N_6270);
or U11445 (N_11445,N_4074,N_4635);
nand U11446 (N_11446,N_5255,N_5045);
or U11447 (N_11447,N_7272,N_7278);
nand U11448 (N_11448,N_6870,N_6294);
and U11449 (N_11449,N_6229,N_6302);
or U11450 (N_11450,N_6364,N_5733);
and U11451 (N_11451,N_7347,N_5895);
and U11452 (N_11452,N_6940,N_4405);
xnor U11453 (N_11453,N_5762,N_7267);
and U11454 (N_11454,N_4084,N_5642);
nand U11455 (N_11455,N_5256,N_5225);
and U11456 (N_11456,N_4149,N_4888);
and U11457 (N_11457,N_7141,N_5069);
or U11458 (N_11458,N_5894,N_7464);
or U11459 (N_11459,N_6241,N_5931);
nand U11460 (N_11460,N_5492,N_6133);
or U11461 (N_11461,N_7217,N_6094);
nand U11462 (N_11462,N_4076,N_4083);
xnor U11463 (N_11463,N_5776,N_6787);
xnor U11464 (N_11464,N_5463,N_7449);
nor U11465 (N_11465,N_7227,N_6095);
nand U11466 (N_11466,N_4567,N_6407);
and U11467 (N_11467,N_6311,N_7984);
nand U11468 (N_11468,N_6604,N_7557);
nand U11469 (N_11469,N_6567,N_6833);
and U11470 (N_11470,N_4413,N_5682);
nor U11471 (N_11471,N_4752,N_4774);
and U11472 (N_11472,N_7887,N_4038);
xor U11473 (N_11473,N_4494,N_4684);
and U11474 (N_11474,N_6540,N_6501);
xnor U11475 (N_11475,N_6409,N_5257);
nand U11476 (N_11476,N_7223,N_7134);
nand U11477 (N_11477,N_4147,N_7401);
nor U11478 (N_11478,N_4723,N_6429);
nand U11479 (N_11479,N_6794,N_5619);
or U11480 (N_11480,N_5310,N_7194);
nor U11481 (N_11481,N_7208,N_6062);
nand U11482 (N_11482,N_6218,N_4167);
nor U11483 (N_11483,N_7569,N_5865);
nor U11484 (N_11484,N_7746,N_6497);
nand U11485 (N_11485,N_5928,N_7311);
or U11486 (N_11486,N_6464,N_5434);
or U11487 (N_11487,N_4194,N_5597);
nand U11488 (N_11488,N_6491,N_7329);
and U11489 (N_11489,N_6248,N_7914);
nor U11490 (N_11490,N_7854,N_7317);
or U11491 (N_11491,N_6573,N_5870);
nor U11492 (N_11492,N_5965,N_6504);
and U11493 (N_11493,N_6373,N_4998);
and U11494 (N_11494,N_5932,N_6654);
or U11495 (N_11495,N_5284,N_7126);
or U11496 (N_11496,N_7459,N_7174);
nand U11497 (N_11497,N_4494,N_5230);
xor U11498 (N_11498,N_5931,N_5299);
nand U11499 (N_11499,N_6307,N_6338);
and U11500 (N_11500,N_4584,N_5454);
nand U11501 (N_11501,N_4538,N_5992);
and U11502 (N_11502,N_4216,N_6431);
xnor U11503 (N_11503,N_4655,N_4902);
or U11504 (N_11504,N_4149,N_4672);
or U11505 (N_11505,N_4311,N_5898);
or U11506 (N_11506,N_5824,N_6272);
nor U11507 (N_11507,N_6444,N_7055);
nand U11508 (N_11508,N_4639,N_6139);
nand U11509 (N_11509,N_7593,N_4492);
nor U11510 (N_11510,N_5295,N_7834);
or U11511 (N_11511,N_7204,N_5395);
nor U11512 (N_11512,N_5410,N_7758);
and U11513 (N_11513,N_6258,N_5356);
or U11514 (N_11514,N_7946,N_6097);
nand U11515 (N_11515,N_5787,N_6643);
nor U11516 (N_11516,N_7780,N_6336);
nand U11517 (N_11517,N_6083,N_5418);
and U11518 (N_11518,N_4456,N_5771);
nand U11519 (N_11519,N_7148,N_7665);
and U11520 (N_11520,N_6717,N_5289);
nor U11521 (N_11521,N_6334,N_5108);
nor U11522 (N_11522,N_7540,N_5239);
xnor U11523 (N_11523,N_6941,N_6387);
or U11524 (N_11524,N_5833,N_6850);
or U11525 (N_11525,N_6181,N_7465);
and U11526 (N_11526,N_7861,N_6129);
or U11527 (N_11527,N_7451,N_4220);
and U11528 (N_11528,N_7072,N_7503);
nor U11529 (N_11529,N_4397,N_5388);
nand U11530 (N_11530,N_5816,N_4266);
and U11531 (N_11531,N_7865,N_6279);
nor U11532 (N_11532,N_6339,N_6524);
nor U11533 (N_11533,N_6980,N_6302);
or U11534 (N_11534,N_4152,N_7826);
nand U11535 (N_11535,N_6036,N_4664);
nand U11536 (N_11536,N_6164,N_5568);
nor U11537 (N_11537,N_6545,N_5332);
xor U11538 (N_11538,N_6180,N_5853);
nand U11539 (N_11539,N_7328,N_7954);
nor U11540 (N_11540,N_5865,N_5614);
and U11541 (N_11541,N_6976,N_7142);
or U11542 (N_11542,N_7600,N_6576);
or U11543 (N_11543,N_5837,N_5455);
or U11544 (N_11544,N_7026,N_5060);
nor U11545 (N_11545,N_4068,N_6954);
nor U11546 (N_11546,N_7962,N_5526);
xnor U11547 (N_11547,N_4947,N_7898);
nand U11548 (N_11548,N_7027,N_5858);
xor U11549 (N_11549,N_7667,N_5518);
and U11550 (N_11550,N_6309,N_5670);
nand U11551 (N_11551,N_6653,N_6529);
and U11552 (N_11552,N_6054,N_5879);
nand U11553 (N_11553,N_5586,N_4851);
nand U11554 (N_11554,N_4032,N_4533);
or U11555 (N_11555,N_6638,N_4816);
and U11556 (N_11556,N_5813,N_5752);
or U11557 (N_11557,N_4736,N_5937);
or U11558 (N_11558,N_4532,N_6803);
nand U11559 (N_11559,N_4791,N_7173);
or U11560 (N_11560,N_5860,N_4796);
nor U11561 (N_11561,N_4126,N_7084);
or U11562 (N_11562,N_6518,N_5122);
or U11563 (N_11563,N_5877,N_7690);
or U11564 (N_11564,N_5085,N_6550);
nor U11565 (N_11565,N_4202,N_4440);
and U11566 (N_11566,N_5102,N_4107);
and U11567 (N_11567,N_7877,N_4247);
and U11568 (N_11568,N_5107,N_4977);
and U11569 (N_11569,N_7975,N_4944);
nand U11570 (N_11570,N_7455,N_7142);
or U11571 (N_11571,N_4659,N_6652);
or U11572 (N_11572,N_6760,N_5496);
or U11573 (N_11573,N_4943,N_4567);
and U11574 (N_11574,N_5073,N_4249);
nand U11575 (N_11575,N_5671,N_7333);
nand U11576 (N_11576,N_4957,N_5243);
xor U11577 (N_11577,N_5282,N_5847);
and U11578 (N_11578,N_4938,N_4988);
and U11579 (N_11579,N_7617,N_7598);
nand U11580 (N_11580,N_7623,N_6167);
nand U11581 (N_11581,N_4608,N_7649);
nand U11582 (N_11582,N_5846,N_5841);
xor U11583 (N_11583,N_7055,N_6847);
xor U11584 (N_11584,N_5296,N_6661);
nor U11585 (N_11585,N_4381,N_4926);
nand U11586 (N_11586,N_5474,N_5096);
or U11587 (N_11587,N_6925,N_7572);
and U11588 (N_11588,N_6212,N_7139);
nand U11589 (N_11589,N_7155,N_4191);
nand U11590 (N_11590,N_6079,N_7233);
nor U11591 (N_11591,N_7304,N_7845);
and U11592 (N_11592,N_7595,N_7231);
nand U11593 (N_11593,N_5087,N_5692);
and U11594 (N_11594,N_7000,N_5095);
and U11595 (N_11595,N_7848,N_5612);
and U11596 (N_11596,N_5446,N_6649);
nor U11597 (N_11597,N_5370,N_5595);
nand U11598 (N_11598,N_6578,N_7408);
and U11599 (N_11599,N_6892,N_5821);
xor U11600 (N_11600,N_5661,N_7951);
xor U11601 (N_11601,N_5070,N_7623);
nor U11602 (N_11602,N_5057,N_5025);
or U11603 (N_11603,N_6781,N_5462);
or U11604 (N_11604,N_5248,N_6375);
nor U11605 (N_11605,N_7643,N_5874);
and U11606 (N_11606,N_5253,N_6494);
or U11607 (N_11607,N_7896,N_5377);
and U11608 (N_11608,N_6120,N_6593);
nand U11609 (N_11609,N_4441,N_7611);
and U11610 (N_11610,N_4748,N_5635);
or U11611 (N_11611,N_5605,N_5951);
nand U11612 (N_11612,N_7338,N_7123);
nor U11613 (N_11613,N_6389,N_5612);
and U11614 (N_11614,N_4157,N_4913);
nand U11615 (N_11615,N_5185,N_4746);
and U11616 (N_11616,N_6046,N_7062);
or U11617 (N_11617,N_6699,N_4559);
and U11618 (N_11618,N_6777,N_4803);
and U11619 (N_11619,N_4416,N_6334);
or U11620 (N_11620,N_7086,N_4270);
or U11621 (N_11621,N_4061,N_5391);
nand U11622 (N_11622,N_7005,N_7924);
xor U11623 (N_11623,N_6893,N_7610);
nor U11624 (N_11624,N_7018,N_4439);
and U11625 (N_11625,N_5465,N_6436);
nand U11626 (N_11626,N_4801,N_4096);
and U11627 (N_11627,N_7572,N_4216);
and U11628 (N_11628,N_7585,N_6665);
and U11629 (N_11629,N_7360,N_4238);
and U11630 (N_11630,N_6039,N_7312);
nand U11631 (N_11631,N_6010,N_4993);
or U11632 (N_11632,N_7374,N_4173);
xor U11633 (N_11633,N_4397,N_5952);
or U11634 (N_11634,N_4407,N_7299);
nor U11635 (N_11635,N_4522,N_6371);
xor U11636 (N_11636,N_6895,N_4147);
or U11637 (N_11637,N_5276,N_6911);
nor U11638 (N_11638,N_5747,N_5898);
or U11639 (N_11639,N_4092,N_7679);
nor U11640 (N_11640,N_7493,N_4074);
or U11641 (N_11641,N_6916,N_6404);
or U11642 (N_11642,N_5707,N_6241);
nor U11643 (N_11643,N_6153,N_6570);
nor U11644 (N_11644,N_4422,N_4819);
or U11645 (N_11645,N_7325,N_6291);
and U11646 (N_11646,N_7469,N_7914);
and U11647 (N_11647,N_5028,N_7000);
nand U11648 (N_11648,N_7633,N_7145);
or U11649 (N_11649,N_5502,N_7157);
and U11650 (N_11650,N_4204,N_4861);
and U11651 (N_11651,N_6871,N_5244);
xor U11652 (N_11652,N_7529,N_7700);
and U11653 (N_11653,N_7337,N_6009);
and U11654 (N_11654,N_7247,N_6515);
nor U11655 (N_11655,N_6682,N_7580);
and U11656 (N_11656,N_4785,N_4774);
nor U11657 (N_11657,N_4332,N_4779);
xor U11658 (N_11658,N_5922,N_5343);
nor U11659 (N_11659,N_7375,N_7968);
and U11660 (N_11660,N_5736,N_4273);
nor U11661 (N_11661,N_4409,N_7434);
nand U11662 (N_11662,N_6677,N_7956);
or U11663 (N_11663,N_5883,N_4455);
or U11664 (N_11664,N_6737,N_7128);
nor U11665 (N_11665,N_6516,N_6975);
nand U11666 (N_11666,N_7366,N_7691);
nor U11667 (N_11667,N_7679,N_5374);
nor U11668 (N_11668,N_4897,N_7550);
xnor U11669 (N_11669,N_4828,N_4145);
or U11670 (N_11670,N_7284,N_6926);
nor U11671 (N_11671,N_5442,N_5945);
and U11672 (N_11672,N_4060,N_4092);
xnor U11673 (N_11673,N_4371,N_5287);
and U11674 (N_11674,N_5291,N_4402);
and U11675 (N_11675,N_4330,N_6378);
nand U11676 (N_11676,N_5331,N_4456);
and U11677 (N_11677,N_7142,N_6942);
nand U11678 (N_11678,N_4221,N_4905);
nor U11679 (N_11679,N_5642,N_5520);
nand U11680 (N_11680,N_7864,N_4763);
nor U11681 (N_11681,N_5391,N_4613);
nand U11682 (N_11682,N_6602,N_7270);
xnor U11683 (N_11683,N_4582,N_6861);
or U11684 (N_11684,N_6141,N_5109);
nor U11685 (N_11685,N_5528,N_4683);
nand U11686 (N_11686,N_4905,N_7304);
nand U11687 (N_11687,N_7211,N_6189);
and U11688 (N_11688,N_5241,N_6089);
nand U11689 (N_11689,N_6542,N_4493);
nand U11690 (N_11690,N_4216,N_4085);
or U11691 (N_11691,N_6733,N_5049);
or U11692 (N_11692,N_5895,N_7961);
and U11693 (N_11693,N_6981,N_5086);
and U11694 (N_11694,N_7654,N_7658);
nand U11695 (N_11695,N_7523,N_7515);
and U11696 (N_11696,N_5852,N_6876);
or U11697 (N_11697,N_4426,N_5832);
and U11698 (N_11698,N_4198,N_7327);
and U11699 (N_11699,N_4681,N_6010);
nand U11700 (N_11700,N_5611,N_7944);
and U11701 (N_11701,N_7583,N_4130);
nor U11702 (N_11702,N_4383,N_4463);
nor U11703 (N_11703,N_5038,N_6596);
nor U11704 (N_11704,N_5215,N_6250);
nand U11705 (N_11705,N_6816,N_7308);
nor U11706 (N_11706,N_5457,N_6917);
or U11707 (N_11707,N_4213,N_4535);
nor U11708 (N_11708,N_4171,N_4991);
xnor U11709 (N_11709,N_7794,N_7122);
or U11710 (N_11710,N_5739,N_5997);
nor U11711 (N_11711,N_4068,N_6299);
nor U11712 (N_11712,N_5579,N_6727);
or U11713 (N_11713,N_5601,N_6044);
xnor U11714 (N_11714,N_6988,N_6479);
nand U11715 (N_11715,N_5898,N_4957);
nand U11716 (N_11716,N_5876,N_4597);
nor U11717 (N_11717,N_6686,N_4516);
and U11718 (N_11718,N_4585,N_6323);
nand U11719 (N_11719,N_7269,N_6213);
nor U11720 (N_11720,N_6099,N_4035);
or U11721 (N_11721,N_7765,N_6662);
nand U11722 (N_11722,N_5535,N_7339);
nor U11723 (N_11723,N_5925,N_5734);
and U11724 (N_11724,N_4940,N_7689);
nor U11725 (N_11725,N_5693,N_5436);
nand U11726 (N_11726,N_4859,N_6055);
and U11727 (N_11727,N_4833,N_5566);
nor U11728 (N_11728,N_7792,N_4803);
or U11729 (N_11729,N_5625,N_5055);
nor U11730 (N_11730,N_5226,N_6514);
nor U11731 (N_11731,N_6295,N_4976);
nand U11732 (N_11732,N_4504,N_6501);
nand U11733 (N_11733,N_7632,N_4472);
nand U11734 (N_11734,N_4045,N_4095);
and U11735 (N_11735,N_7023,N_6185);
nor U11736 (N_11736,N_5198,N_7444);
or U11737 (N_11737,N_5875,N_6096);
nor U11738 (N_11738,N_6904,N_4412);
nand U11739 (N_11739,N_5845,N_5104);
nand U11740 (N_11740,N_4338,N_4676);
nand U11741 (N_11741,N_6584,N_6818);
nand U11742 (N_11742,N_5731,N_6010);
and U11743 (N_11743,N_7312,N_6870);
or U11744 (N_11744,N_4550,N_7392);
nor U11745 (N_11745,N_6754,N_5161);
nor U11746 (N_11746,N_6228,N_6367);
nand U11747 (N_11747,N_5402,N_7524);
nor U11748 (N_11748,N_6002,N_5102);
xor U11749 (N_11749,N_6573,N_7174);
nor U11750 (N_11750,N_7437,N_5141);
nor U11751 (N_11751,N_6026,N_4189);
or U11752 (N_11752,N_4113,N_7831);
xor U11753 (N_11753,N_4959,N_7903);
nand U11754 (N_11754,N_7120,N_7184);
nor U11755 (N_11755,N_4764,N_5129);
nand U11756 (N_11756,N_7564,N_5403);
nor U11757 (N_11757,N_4319,N_6734);
xor U11758 (N_11758,N_6598,N_7184);
and U11759 (N_11759,N_5484,N_4769);
and U11760 (N_11760,N_7357,N_5888);
nand U11761 (N_11761,N_6156,N_5936);
nand U11762 (N_11762,N_7729,N_7826);
or U11763 (N_11763,N_7420,N_4306);
xor U11764 (N_11764,N_6072,N_4020);
nor U11765 (N_11765,N_7642,N_6727);
or U11766 (N_11766,N_7682,N_6304);
nand U11767 (N_11767,N_4654,N_5969);
or U11768 (N_11768,N_5826,N_5294);
nor U11769 (N_11769,N_7367,N_7388);
nand U11770 (N_11770,N_5540,N_7704);
and U11771 (N_11771,N_7769,N_5182);
and U11772 (N_11772,N_6708,N_4172);
and U11773 (N_11773,N_6555,N_5333);
and U11774 (N_11774,N_6967,N_5652);
and U11775 (N_11775,N_4987,N_4256);
nor U11776 (N_11776,N_5495,N_5280);
and U11777 (N_11777,N_7788,N_7381);
xor U11778 (N_11778,N_6167,N_4586);
or U11779 (N_11779,N_7714,N_4500);
nor U11780 (N_11780,N_7006,N_4701);
and U11781 (N_11781,N_7029,N_4125);
or U11782 (N_11782,N_7334,N_7600);
and U11783 (N_11783,N_4648,N_6070);
or U11784 (N_11784,N_7526,N_5758);
and U11785 (N_11785,N_6385,N_6832);
and U11786 (N_11786,N_4911,N_6002);
and U11787 (N_11787,N_7090,N_6987);
and U11788 (N_11788,N_6401,N_5626);
nor U11789 (N_11789,N_4120,N_4486);
or U11790 (N_11790,N_6743,N_5925);
nor U11791 (N_11791,N_7735,N_6213);
or U11792 (N_11792,N_5047,N_7684);
or U11793 (N_11793,N_6745,N_4109);
and U11794 (N_11794,N_5298,N_7746);
nand U11795 (N_11795,N_6416,N_7085);
nand U11796 (N_11796,N_5302,N_4778);
nor U11797 (N_11797,N_4186,N_7967);
or U11798 (N_11798,N_7316,N_6462);
and U11799 (N_11799,N_7576,N_5173);
nand U11800 (N_11800,N_6821,N_5780);
xnor U11801 (N_11801,N_4563,N_6738);
nand U11802 (N_11802,N_4792,N_4482);
nand U11803 (N_11803,N_6435,N_4821);
nor U11804 (N_11804,N_6217,N_4136);
and U11805 (N_11805,N_5161,N_4126);
nor U11806 (N_11806,N_7428,N_6473);
and U11807 (N_11807,N_5651,N_7318);
xor U11808 (N_11808,N_5389,N_4298);
or U11809 (N_11809,N_4233,N_6371);
nand U11810 (N_11810,N_6665,N_7991);
or U11811 (N_11811,N_6942,N_4035);
or U11812 (N_11812,N_5936,N_5061);
or U11813 (N_11813,N_5793,N_7588);
nor U11814 (N_11814,N_6045,N_4946);
or U11815 (N_11815,N_5225,N_6152);
or U11816 (N_11816,N_4028,N_7037);
and U11817 (N_11817,N_5649,N_7131);
xnor U11818 (N_11818,N_6559,N_7965);
and U11819 (N_11819,N_4916,N_7971);
and U11820 (N_11820,N_7325,N_5871);
nor U11821 (N_11821,N_5208,N_4645);
or U11822 (N_11822,N_5884,N_6066);
nor U11823 (N_11823,N_6271,N_6121);
or U11824 (N_11824,N_7650,N_7059);
nor U11825 (N_11825,N_4311,N_5300);
xor U11826 (N_11826,N_6659,N_4295);
and U11827 (N_11827,N_5491,N_6400);
nor U11828 (N_11828,N_4067,N_6193);
nand U11829 (N_11829,N_7449,N_5192);
and U11830 (N_11830,N_6614,N_5817);
and U11831 (N_11831,N_4160,N_4090);
or U11832 (N_11832,N_5178,N_4164);
and U11833 (N_11833,N_4654,N_6778);
nor U11834 (N_11834,N_5842,N_6207);
nor U11835 (N_11835,N_4292,N_6223);
and U11836 (N_11836,N_5968,N_6283);
or U11837 (N_11837,N_6055,N_7050);
nand U11838 (N_11838,N_6893,N_6219);
or U11839 (N_11839,N_4057,N_7069);
and U11840 (N_11840,N_4283,N_6532);
or U11841 (N_11841,N_4431,N_6849);
or U11842 (N_11842,N_5474,N_6074);
or U11843 (N_11843,N_4937,N_5255);
or U11844 (N_11844,N_7679,N_6947);
nand U11845 (N_11845,N_5720,N_7253);
or U11846 (N_11846,N_5484,N_7149);
nor U11847 (N_11847,N_7014,N_5111);
or U11848 (N_11848,N_4800,N_7464);
nand U11849 (N_11849,N_6909,N_4101);
or U11850 (N_11850,N_4219,N_5593);
nor U11851 (N_11851,N_7435,N_7035);
nor U11852 (N_11852,N_5937,N_6314);
nand U11853 (N_11853,N_4118,N_4654);
nand U11854 (N_11854,N_7053,N_7595);
or U11855 (N_11855,N_7061,N_7887);
or U11856 (N_11856,N_7851,N_6844);
nor U11857 (N_11857,N_6056,N_4976);
and U11858 (N_11858,N_4091,N_7377);
or U11859 (N_11859,N_5401,N_4593);
nor U11860 (N_11860,N_7975,N_4016);
and U11861 (N_11861,N_6117,N_6478);
or U11862 (N_11862,N_4782,N_5560);
nand U11863 (N_11863,N_5034,N_5443);
or U11864 (N_11864,N_4551,N_4209);
nand U11865 (N_11865,N_6896,N_7826);
and U11866 (N_11866,N_5867,N_7663);
or U11867 (N_11867,N_7121,N_7105);
nor U11868 (N_11868,N_7146,N_7389);
or U11869 (N_11869,N_7346,N_5874);
nand U11870 (N_11870,N_6071,N_7522);
or U11871 (N_11871,N_4707,N_6723);
nor U11872 (N_11872,N_6690,N_4415);
xor U11873 (N_11873,N_4623,N_7334);
nand U11874 (N_11874,N_7479,N_6311);
or U11875 (N_11875,N_7991,N_6296);
xnor U11876 (N_11876,N_4858,N_4305);
nor U11877 (N_11877,N_6087,N_7084);
and U11878 (N_11878,N_7973,N_6583);
xnor U11879 (N_11879,N_4940,N_6589);
or U11880 (N_11880,N_6706,N_6090);
nand U11881 (N_11881,N_6180,N_5371);
xor U11882 (N_11882,N_6910,N_6124);
and U11883 (N_11883,N_4515,N_6850);
nand U11884 (N_11884,N_4682,N_4371);
nor U11885 (N_11885,N_7698,N_6082);
nor U11886 (N_11886,N_5787,N_6472);
or U11887 (N_11887,N_6154,N_7474);
nand U11888 (N_11888,N_6649,N_7850);
nor U11889 (N_11889,N_7072,N_4197);
xnor U11890 (N_11890,N_4114,N_5863);
xnor U11891 (N_11891,N_7865,N_7945);
or U11892 (N_11892,N_5309,N_6062);
nand U11893 (N_11893,N_7710,N_5761);
nor U11894 (N_11894,N_6556,N_4989);
xor U11895 (N_11895,N_4873,N_6017);
and U11896 (N_11896,N_6582,N_7409);
and U11897 (N_11897,N_4911,N_4557);
xor U11898 (N_11898,N_6200,N_6392);
nor U11899 (N_11899,N_4107,N_7305);
nor U11900 (N_11900,N_7142,N_7974);
and U11901 (N_11901,N_5086,N_5071);
or U11902 (N_11902,N_6691,N_4229);
nor U11903 (N_11903,N_6117,N_5560);
nand U11904 (N_11904,N_4039,N_7839);
nor U11905 (N_11905,N_4250,N_7826);
and U11906 (N_11906,N_7409,N_7969);
nand U11907 (N_11907,N_4161,N_7797);
or U11908 (N_11908,N_6387,N_4896);
nor U11909 (N_11909,N_6742,N_5497);
nor U11910 (N_11910,N_7949,N_5993);
nand U11911 (N_11911,N_7794,N_5422);
or U11912 (N_11912,N_7559,N_7172);
nand U11913 (N_11913,N_4823,N_4276);
and U11914 (N_11914,N_5943,N_7984);
and U11915 (N_11915,N_7734,N_6218);
and U11916 (N_11916,N_4865,N_7516);
nor U11917 (N_11917,N_6134,N_4395);
and U11918 (N_11918,N_6939,N_6513);
and U11919 (N_11919,N_5561,N_4904);
xnor U11920 (N_11920,N_5054,N_7939);
nor U11921 (N_11921,N_7340,N_4727);
nor U11922 (N_11922,N_5623,N_7837);
nor U11923 (N_11923,N_4416,N_5644);
nand U11924 (N_11924,N_5943,N_6841);
nor U11925 (N_11925,N_7587,N_7780);
and U11926 (N_11926,N_4926,N_7334);
nor U11927 (N_11927,N_7292,N_6638);
nor U11928 (N_11928,N_6192,N_6850);
nor U11929 (N_11929,N_4384,N_7937);
or U11930 (N_11930,N_6737,N_7869);
and U11931 (N_11931,N_5699,N_6287);
nor U11932 (N_11932,N_4223,N_6765);
nand U11933 (N_11933,N_5095,N_7887);
or U11934 (N_11934,N_6851,N_5619);
nand U11935 (N_11935,N_5263,N_5433);
and U11936 (N_11936,N_6746,N_6611);
and U11937 (N_11937,N_5155,N_4667);
nand U11938 (N_11938,N_5611,N_6935);
and U11939 (N_11939,N_6122,N_7220);
and U11940 (N_11940,N_6696,N_5316);
nand U11941 (N_11941,N_7221,N_6750);
and U11942 (N_11942,N_6646,N_5301);
or U11943 (N_11943,N_4003,N_5765);
or U11944 (N_11944,N_7742,N_4317);
nor U11945 (N_11945,N_4579,N_6677);
nor U11946 (N_11946,N_5094,N_7704);
nand U11947 (N_11947,N_5660,N_4778);
nand U11948 (N_11948,N_4981,N_6492);
and U11949 (N_11949,N_4481,N_7708);
and U11950 (N_11950,N_6566,N_5872);
and U11951 (N_11951,N_7093,N_4051);
nor U11952 (N_11952,N_7807,N_6908);
and U11953 (N_11953,N_4921,N_6201);
or U11954 (N_11954,N_5699,N_5981);
nand U11955 (N_11955,N_7379,N_5909);
or U11956 (N_11956,N_7356,N_7093);
and U11957 (N_11957,N_7910,N_6928);
or U11958 (N_11958,N_6643,N_6785);
nand U11959 (N_11959,N_4105,N_7356);
xnor U11960 (N_11960,N_7291,N_4700);
or U11961 (N_11961,N_4549,N_5909);
nand U11962 (N_11962,N_7192,N_6286);
nor U11963 (N_11963,N_4434,N_7471);
or U11964 (N_11964,N_5683,N_4868);
xor U11965 (N_11965,N_6667,N_6145);
nor U11966 (N_11966,N_4941,N_4434);
xor U11967 (N_11967,N_6378,N_4350);
or U11968 (N_11968,N_7344,N_5122);
and U11969 (N_11969,N_6298,N_5166);
xnor U11970 (N_11970,N_4223,N_4683);
or U11971 (N_11971,N_7106,N_5926);
nand U11972 (N_11972,N_7826,N_4206);
nor U11973 (N_11973,N_5973,N_5681);
and U11974 (N_11974,N_7192,N_7721);
and U11975 (N_11975,N_6894,N_5405);
or U11976 (N_11976,N_5151,N_7899);
and U11977 (N_11977,N_7826,N_5822);
nand U11978 (N_11978,N_4269,N_7000);
nand U11979 (N_11979,N_6134,N_5898);
xnor U11980 (N_11980,N_4986,N_5067);
and U11981 (N_11981,N_6254,N_6291);
or U11982 (N_11982,N_7957,N_5547);
or U11983 (N_11983,N_5865,N_6105);
nor U11984 (N_11984,N_6149,N_6374);
nand U11985 (N_11985,N_7607,N_7980);
nand U11986 (N_11986,N_5324,N_6258);
or U11987 (N_11987,N_5985,N_4737);
xnor U11988 (N_11988,N_5286,N_7822);
or U11989 (N_11989,N_5853,N_5814);
or U11990 (N_11990,N_5165,N_4596);
nand U11991 (N_11991,N_7068,N_5116);
xor U11992 (N_11992,N_4785,N_7921);
or U11993 (N_11993,N_6309,N_4954);
nor U11994 (N_11994,N_7458,N_7628);
or U11995 (N_11995,N_5788,N_5461);
or U11996 (N_11996,N_7368,N_7271);
and U11997 (N_11997,N_6455,N_5903);
nand U11998 (N_11998,N_5470,N_4602);
nor U11999 (N_11999,N_6338,N_6075);
nor U12000 (N_12000,N_8813,N_11871);
or U12001 (N_12001,N_8597,N_8009);
nand U12002 (N_12002,N_11701,N_9619);
nand U12003 (N_12003,N_10910,N_11323);
or U12004 (N_12004,N_9540,N_10147);
xnor U12005 (N_12005,N_11511,N_9927);
xnor U12006 (N_12006,N_9232,N_10134);
and U12007 (N_12007,N_8335,N_11410);
or U12008 (N_12008,N_11003,N_9018);
and U12009 (N_12009,N_9177,N_10677);
nor U12010 (N_12010,N_8300,N_8368);
or U12011 (N_12011,N_10660,N_8843);
xnor U12012 (N_12012,N_9035,N_8964);
or U12013 (N_12013,N_9276,N_11508);
xnor U12014 (N_12014,N_8556,N_10383);
xnor U12015 (N_12015,N_10672,N_8747);
nand U12016 (N_12016,N_9911,N_11050);
or U12017 (N_12017,N_10690,N_11202);
or U12018 (N_12018,N_8148,N_8541);
nand U12019 (N_12019,N_11691,N_10011);
or U12020 (N_12020,N_11320,N_8583);
and U12021 (N_12021,N_8827,N_10356);
and U12022 (N_12022,N_9153,N_9077);
and U12023 (N_12023,N_11772,N_9214);
and U12024 (N_12024,N_11617,N_8432);
or U12025 (N_12025,N_8135,N_10069);
and U12026 (N_12026,N_11499,N_10237);
nand U12027 (N_12027,N_11404,N_9994);
nor U12028 (N_12028,N_11147,N_11067);
nand U12029 (N_12029,N_10859,N_8077);
or U12030 (N_12030,N_10131,N_8088);
xnor U12031 (N_12031,N_11221,N_9109);
or U12032 (N_12032,N_9612,N_11056);
nand U12033 (N_12033,N_9262,N_10145);
nor U12034 (N_12034,N_11406,N_10937);
nand U12035 (N_12035,N_11207,N_11969);
or U12036 (N_12036,N_8938,N_9854);
and U12037 (N_12037,N_10430,N_9590);
nand U12038 (N_12038,N_8347,N_9773);
or U12039 (N_12039,N_8861,N_11110);
and U12040 (N_12040,N_10819,N_9939);
nor U12041 (N_12041,N_11914,N_8988);
nor U12042 (N_12042,N_11861,N_8808);
and U12043 (N_12043,N_11562,N_11084);
or U12044 (N_12044,N_10346,N_8134);
nand U12045 (N_12045,N_10454,N_9302);
nor U12046 (N_12046,N_8119,N_9755);
or U12047 (N_12047,N_8174,N_8914);
and U12048 (N_12048,N_8224,N_9506);
and U12049 (N_12049,N_8099,N_9861);
nand U12050 (N_12050,N_11875,N_11703);
and U12051 (N_12051,N_8168,N_9986);
nor U12052 (N_12052,N_8971,N_11642);
xor U12053 (N_12053,N_9389,N_8092);
and U12054 (N_12054,N_10641,N_10728);
xor U12055 (N_12055,N_11866,N_10727);
nand U12056 (N_12056,N_8950,N_9547);
xnor U12057 (N_12057,N_9410,N_11347);
or U12058 (N_12058,N_8535,N_10038);
xor U12059 (N_12059,N_8820,N_9334);
or U12060 (N_12060,N_9467,N_8001);
or U12061 (N_12061,N_11242,N_10911);
or U12062 (N_12062,N_8703,N_8452);
or U12063 (N_12063,N_8522,N_9909);
or U12064 (N_12064,N_9455,N_9408);
nor U12065 (N_12065,N_10741,N_8891);
and U12066 (N_12066,N_9373,N_10206);
and U12067 (N_12067,N_8336,N_8725);
nand U12068 (N_12068,N_11695,N_9576);
or U12069 (N_12069,N_9426,N_11466);
xor U12070 (N_12070,N_11124,N_10758);
nand U12071 (N_12071,N_8763,N_10839);
or U12072 (N_12072,N_10675,N_9258);
xnor U12073 (N_12073,N_11724,N_9943);
nand U12074 (N_12074,N_8577,N_11343);
nand U12075 (N_12075,N_11089,N_10879);
nand U12076 (N_12076,N_9793,N_10415);
nand U12077 (N_12077,N_10354,N_8275);
xor U12078 (N_12078,N_10045,N_11986);
or U12079 (N_12079,N_11713,N_10973);
and U12080 (N_12080,N_10496,N_10938);
nand U12081 (N_12081,N_11967,N_8289);
and U12082 (N_12082,N_11057,N_11693);
or U12083 (N_12083,N_10136,N_9891);
and U12084 (N_12084,N_8338,N_8481);
xnor U12085 (N_12085,N_8952,N_8345);
or U12086 (N_12086,N_8052,N_8666);
xor U12087 (N_12087,N_8061,N_9197);
or U12088 (N_12088,N_8467,N_10593);
xnor U12089 (N_12089,N_11767,N_8068);
xnor U12090 (N_12090,N_8093,N_9688);
nand U12091 (N_12091,N_10546,N_11328);
or U12092 (N_12092,N_11162,N_9341);
nor U12093 (N_12093,N_11414,N_9299);
or U12094 (N_12094,N_9108,N_10046);
nor U12095 (N_12095,N_10708,N_10407);
nor U12096 (N_12096,N_8206,N_8863);
xnor U12097 (N_12097,N_10271,N_11224);
and U12098 (N_12098,N_11658,N_11243);
or U12099 (N_12099,N_10850,N_9818);
and U12100 (N_12100,N_8558,N_11337);
or U12101 (N_12101,N_9697,N_8881);
and U12102 (N_12102,N_8854,N_10693);
nor U12103 (N_12103,N_9963,N_10132);
nor U12104 (N_12104,N_9951,N_10670);
nand U12105 (N_12105,N_10023,N_9736);
nand U12106 (N_12106,N_10860,N_9451);
nand U12107 (N_12107,N_9990,N_9100);
and U12108 (N_12108,N_9388,N_11058);
or U12109 (N_12109,N_10054,N_11201);
nand U12110 (N_12110,N_9575,N_8448);
nor U12111 (N_12111,N_11816,N_8635);
nand U12112 (N_12112,N_9694,N_10994);
xor U12113 (N_12113,N_11315,N_9032);
or U12114 (N_12114,N_9156,N_11311);
and U12115 (N_12115,N_10807,N_8401);
nand U12116 (N_12116,N_9545,N_10156);
xor U12117 (N_12117,N_8816,N_8757);
and U12118 (N_12118,N_8250,N_9304);
or U12119 (N_12119,N_10041,N_11012);
nor U12120 (N_12120,N_8931,N_10781);
nor U12121 (N_12121,N_11291,N_9558);
or U12122 (N_12122,N_9744,N_11572);
and U12123 (N_12123,N_9811,N_11900);
nor U12124 (N_12124,N_9283,N_11533);
nand U12125 (N_12125,N_8160,N_9526);
nor U12126 (N_12126,N_10296,N_8679);
or U12127 (N_12127,N_11000,N_11262);
nand U12128 (N_12128,N_10886,N_8949);
and U12129 (N_12129,N_10352,N_11752);
nor U12130 (N_12130,N_10272,N_9541);
nor U12131 (N_12131,N_10836,N_10684);
nand U12132 (N_12132,N_9358,N_11220);
nor U12133 (N_12133,N_10800,N_10328);
or U12134 (N_12134,N_11237,N_9192);
or U12135 (N_12135,N_11033,N_10682);
nand U12136 (N_12136,N_10788,N_11746);
nor U12137 (N_12137,N_9556,N_8766);
nand U12138 (N_12138,N_8210,N_8291);
or U12139 (N_12139,N_11500,N_8887);
and U12140 (N_12140,N_9960,N_10516);
xnor U12141 (N_12141,N_8053,N_10082);
nor U12142 (N_12142,N_9791,N_10390);
xor U12143 (N_12143,N_8181,N_8711);
or U12144 (N_12144,N_11122,N_11775);
nand U12145 (N_12145,N_8268,N_11281);
and U12146 (N_12146,N_8500,N_8909);
or U12147 (N_12147,N_10412,N_9667);
nand U12148 (N_12148,N_9290,N_11269);
nand U12149 (N_12149,N_11796,N_10561);
and U12150 (N_12150,N_11626,N_10729);
nor U12151 (N_12151,N_10774,N_9549);
and U12152 (N_12152,N_11132,N_10611);
and U12153 (N_12153,N_11388,N_11360);
or U12154 (N_12154,N_8604,N_9086);
or U12155 (N_12155,N_10101,N_11023);
or U12156 (N_12156,N_10289,N_10386);
nand U12157 (N_12157,N_11459,N_9132);
xnor U12158 (N_12158,N_9537,N_8959);
nor U12159 (N_12159,N_8376,N_11167);
xor U12160 (N_12160,N_10278,N_9899);
and U12161 (N_12161,N_9785,N_10901);
and U12162 (N_12162,N_9011,N_9001);
and U12163 (N_12163,N_11120,N_9727);
xor U12164 (N_12164,N_11799,N_9259);
nor U12165 (N_12165,N_11706,N_10640);
or U12166 (N_12166,N_11219,N_11541);
and U12167 (N_12167,N_10077,N_10548);
xnor U12168 (N_12168,N_11098,N_11893);
nor U12169 (N_12169,N_11725,N_8407);
and U12170 (N_12170,N_10923,N_8672);
nor U12171 (N_12171,N_9554,N_8613);
and U12172 (N_12172,N_9106,N_9980);
or U12173 (N_12173,N_8779,N_11905);
and U12174 (N_12174,N_8408,N_11214);
and U12175 (N_12175,N_8348,N_8239);
and U12176 (N_12176,N_10264,N_11608);
and U12177 (N_12177,N_10713,N_9870);
xnor U12178 (N_12178,N_9300,N_8150);
nor U12179 (N_12179,N_10441,N_9336);
and U12180 (N_12180,N_10019,N_10018);
and U12181 (N_12181,N_11524,N_11685);
nand U12182 (N_12182,N_8457,N_11088);
or U12183 (N_12183,N_8502,N_8791);
nand U12184 (N_12184,N_9265,N_8020);
or U12185 (N_12185,N_10298,N_10429);
nand U12186 (N_12186,N_9551,N_9956);
and U12187 (N_12187,N_9977,N_10432);
nand U12188 (N_12188,N_8418,N_9401);
nor U12189 (N_12189,N_8127,N_9116);
or U12190 (N_12190,N_10811,N_8625);
and U12191 (N_12191,N_10266,N_11616);
nand U12192 (N_12192,N_9913,N_10766);
nor U12193 (N_12193,N_8006,N_8724);
nor U12194 (N_12194,N_8618,N_9435);
nor U12195 (N_12195,N_9841,N_10616);
and U12196 (N_12196,N_11631,N_11478);
nor U12197 (N_12197,N_8341,N_8086);
nand U12198 (N_12198,N_9127,N_10532);
and U12199 (N_12199,N_9031,N_10455);
and U12200 (N_12200,N_11377,N_11559);
nor U12201 (N_12201,N_11356,N_10381);
or U12202 (N_12202,N_8393,N_8149);
or U12203 (N_12203,N_8510,N_10529);
nand U12204 (N_12204,N_9488,N_10104);
or U12205 (N_12205,N_11303,N_9428);
and U12206 (N_12206,N_9607,N_8975);
and U12207 (N_12207,N_8745,N_8799);
nor U12208 (N_12208,N_9042,N_10985);
nor U12209 (N_12209,N_8389,N_8734);
nor U12210 (N_12210,N_10358,N_9118);
and U12211 (N_12211,N_8449,N_10128);
or U12212 (N_12212,N_8155,N_8851);
and U12213 (N_12213,N_10436,N_10148);
and U12214 (N_12214,N_8531,N_8069);
or U12215 (N_12215,N_11896,N_11462);
and U12216 (N_12216,N_8632,N_8411);
xor U12217 (N_12217,N_9840,N_11427);
and U12218 (N_12218,N_10783,N_9338);
or U12219 (N_12219,N_9738,N_9495);
nor U12220 (N_12220,N_10825,N_11546);
nand U12221 (N_12221,N_8424,N_11665);
and U12222 (N_12222,N_10085,N_8298);
and U12223 (N_12223,N_9940,N_10342);
nor U12224 (N_12224,N_9346,N_9926);
or U12225 (N_12225,N_8044,N_9037);
or U12226 (N_12226,N_9313,N_8888);
nand U12227 (N_12227,N_10559,N_10989);
and U12228 (N_12228,N_8285,N_8790);
xor U12229 (N_12229,N_9459,N_9616);
nand U12230 (N_12230,N_10004,N_11881);
or U12231 (N_12231,N_10756,N_11763);
and U12232 (N_12232,N_9016,N_9089);
or U12233 (N_12233,N_10120,N_9181);
and U12234 (N_12234,N_11826,N_8494);
nand U12235 (N_12235,N_10040,N_8018);
or U12236 (N_12236,N_9280,N_11346);
or U12237 (N_12237,N_8417,N_8762);
nand U12238 (N_12238,N_8292,N_8100);
and U12239 (N_12239,N_10957,N_11699);
nand U12240 (N_12240,N_8744,N_10830);
nand U12241 (N_12241,N_11362,N_11198);
xnor U12242 (N_12242,N_9725,N_9687);
and U12243 (N_12243,N_9344,N_9124);
or U12244 (N_12244,N_11635,N_8640);
and U12245 (N_12245,N_10541,N_11102);
nor U12246 (N_12246,N_10870,N_9119);
and U12247 (N_12247,N_8079,N_10715);
or U12248 (N_12248,N_9593,N_8933);
nand U12249 (N_12249,N_9111,N_9163);
xor U12250 (N_12250,N_9524,N_9708);
or U12251 (N_12251,N_11750,N_8855);
or U12252 (N_12252,N_11068,N_8874);
nor U12253 (N_12253,N_10487,N_8824);
nor U12254 (N_12254,N_11059,N_10469);
nor U12255 (N_12255,N_8805,N_9752);
or U12256 (N_12256,N_9808,N_8430);
xor U12257 (N_12257,N_8939,N_9824);
or U12258 (N_12258,N_10008,N_8850);
nor U12259 (N_12259,N_9843,N_8777);
xor U12260 (N_12260,N_9157,N_9166);
nor U12261 (N_12261,N_11731,N_11456);
xnor U12262 (N_12262,N_8165,N_9501);
or U12263 (N_12263,N_10891,N_9850);
nor U12264 (N_12264,N_8450,N_11127);
xor U12265 (N_12265,N_10627,N_9099);
nor U12266 (N_12266,N_8587,N_9005);
and U12267 (N_12267,N_10501,N_11189);
or U12268 (N_12268,N_9178,N_11501);
and U12269 (N_12269,N_11906,N_11946);
and U12270 (N_12270,N_9930,N_9269);
and U12271 (N_12271,N_8839,N_10287);
nor U12272 (N_12272,N_10301,N_8471);
nand U12273 (N_12273,N_11191,N_9047);
and U12274 (N_12274,N_10417,N_11686);
and U12275 (N_12275,N_8492,N_10483);
or U12276 (N_12276,N_9151,N_8444);
xor U12277 (N_12277,N_9226,N_8845);
nor U12278 (N_12278,N_11381,N_9933);
xor U12279 (N_12279,N_11705,N_11854);
and U12280 (N_12280,N_11828,N_11421);
nor U12281 (N_12281,N_8066,N_11727);
nor U12282 (N_12282,N_11983,N_10709);
and U12283 (N_12283,N_11436,N_10404);
and U12284 (N_12284,N_10798,N_11199);
nand U12285 (N_12285,N_9757,N_8037);
and U12286 (N_12286,N_8897,N_9603);
nor U12287 (N_12287,N_11718,N_9182);
and U12288 (N_12288,N_9239,N_11489);
and U12289 (N_12289,N_11047,N_10138);
or U12290 (N_12290,N_10314,N_11390);
and U12291 (N_12291,N_9393,N_8704);
and U12292 (N_12292,N_10574,N_9268);
nand U12293 (N_12293,N_9491,N_8657);
xor U12294 (N_12294,N_11288,N_8366);
and U12295 (N_12295,N_9746,N_10599);
or U12296 (N_12296,N_8241,N_11391);
and U12297 (N_12297,N_8176,N_11113);
and U12298 (N_12298,N_11105,N_9286);
and U12299 (N_12299,N_10714,N_9470);
nor U12300 (N_12300,N_10090,N_8563);
nor U12301 (N_12301,N_8797,N_11254);
nand U12302 (N_12302,N_10519,N_10312);
nand U12303 (N_12303,N_8919,N_11299);
xnor U12304 (N_12304,N_11240,N_11045);
xor U12305 (N_12305,N_9219,N_8167);
or U12306 (N_12306,N_11134,N_9764);
or U12307 (N_12307,N_10880,N_8385);
and U12308 (N_12308,N_8955,N_10423);
or U12309 (N_12309,N_9997,N_10244);
nor U12310 (N_12310,N_10367,N_10854);
nand U12311 (N_12311,N_9270,N_11136);
or U12312 (N_12312,N_11259,N_9985);
nand U12313 (N_12313,N_11819,N_10315);
or U12314 (N_12314,N_10198,N_11095);
and U12315 (N_12315,N_11223,N_8673);
and U12316 (N_12316,N_11643,N_8078);
xor U12317 (N_12317,N_9272,N_10621);
nor U12318 (N_12318,N_8621,N_11869);
xor U12319 (N_12319,N_10213,N_8178);
and U12320 (N_12320,N_9029,N_11402);
or U12321 (N_12321,N_9665,N_10292);
nand U12322 (N_12322,N_9320,N_9503);
nand U12323 (N_12323,N_10340,N_11283);
nor U12324 (N_12324,N_8683,N_11368);
nand U12325 (N_12325,N_8474,N_10100);
nor U12326 (N_12326,N_11352,N_9924);
nand U12327 (N_12327,N_9199,N_11780);
nand U12328 (N_12328,N_11788,N_8876);
and U12329 (N_12329,N_8163,N_8445);
and U12330 (N_12330,N_10634,N_11521);
and U12331 (N_12331,N_10248,N_9555);
nor U12332 (N_12332,N_9550,N_9816);
or U12333 (N_12333,N_11115,N_9150);
nor U12334 (N_12334,N_8670,N_11185);
and U12335 (N_12335,N_10558,N_10176);
nor U12336 (N_12336,N_8076,N_10130);
or U12337 (N_12337,N_9789,N_8332);
nand U12338 (N_12338,N_8764,N_8866);
nand U12339 (N_12339,N_11968,N_10170);
and U12340 (N_12340,N_8459,N_10928);
nand U12341 (N_12341,N_9456,N_8030);
and U12342 (N_12342,N_10782,N_9525);
and U12343 (N_12343,N_11837,N_10965);
nand U12344 (N_12344,N_9059,N_8840);
nand U12345 (N_12345,N_10916,N_11304);
nor U12346 (N_12346,N_9264,N_11895);
nand U12347 (N_12347,N_9314,N_9460);
or U12348 (N_12348,N_9916,N_11632);
and U12349 (N_12349,N_9027,N_9235);
nor U12350 (N_12350,N_11492,N_9093);
xnor U12351 (N_12351,N_9819,N_8025);
or U12352 (N_12352,N_8442,N_10052);
and U12353 (N_12353,N_11082,N_10117);
and U12354 (N_12354,N_10304,N_10614);
nor U12355 (N_12355,N_9374,N_10012);
and U12356 (N_12356,N_10983,N_9063);
and U12357 (N_12357,N_9677,N_9121);
or U12358 (N_12358,N_8247,N_11812);
nand U12359 (N_12359,N_10349,N_10696);
or U12360 (N_12360,N_10321,N_8246);
nor U12361 (N_12361,N_9632,N_8647);
or U12362 (N_12362,N_9068,N_9759);
and U12363 (N_12363,N_10745,N_11026);
nor U12364 (N_12364,N_9002,N_11104);
and U12365 (N_12365,N_8046,N_10030);
and U12366 (N_12366,N_11548,N_9586);
nand U12367 (N_12367,N_9630,N_11971);
nor U12368 (N_12368,N_10944,N_10632);
xnor U12369 (N_12369,N_11553,N_10853);
and U12370 (N_12370,N_8911,N_9141);
or U12371 (N_12371,N_10053,N_11878);
nor U12372 (N_12372,N_8981,N_11678);
nor U12373 (N_12373,N_10482,N_10344);
nand U12374 (N_12374,N_10801,N_8743);
or U12375 (N_12375,N_8537,N_10168);
nand U12376 (N_12376,N_10918,N_10635);
nand U12377 (N_12377,N_8141,N_10262);
or U12378 (N_12378,N_9648,N_8190);
nand U12379 (N_12379,N_9303,N_10309);
and U12380 (N_12380,N_11251,N_9686);
and U12381 (N_12381,N_9365,N_11129);
xor U12382 (N_12382,N_8473,N_11962);
or U12383 (N_12383,N_10179,N_8781);
nor U12384 (N_12384,N_8352,N_11322);
or U12385 (N_12385,N_8831,N_8898);
and U12386 (N_12386,N_8982,N_10195);
nor U12387 (N_12387,N_10688,N_8458);
nor U12388 (N_12388,N_8833,N_9340);
and U12389 (N_12389,N_10981,N_10215);
or U12390 (N_12390,N_11934,N_10236);
or U12391 (N_12391,N_8288,N_10705);
nor U12392 (N_12392,N_10153,N_11929);
nand U12393 (N_12393,N_10007,N_9613);
nand U12394 (N_12394,N_8259,N_11439);
nor U12395 (N_12395,N_10355,N_11446);
or U12396 (N_12396,N_10975,N_10096);
nand U12397 (N_12397,N_10687,N_10259);
nand U12398 (N_12398,N_11180,N_8050);
nor U12399 (N_12399,N_9003,N_10765);
nor U12400 (N_12400,N_8547,N_10458);
nand U12401 (N_12401,N_11190,N_8049);
xor U12402 (N_12402,N_11771,N_10031);
nand U12403 (N_12403,N_11013,N_9568);
or U12404 (N_12404,N_8598,N_10322);
nor U12405 (N_12405,N_11923,N_9790);
or U12406 (N_12406,N_10929,N_8399);
or U12407 (N_12407,N_10409,N_8652);
and U12408 (N_12408,N_10803,N_9233);
or U12409 (N_12409,N_10284,N_9581);
nand U12410 (N_12410,N_9777,N_9802);
and U12411 (N_12411,N_11942,N_8186);
xor U12412 (N_12412,N_11966,N_10171);
and U12413 (N_12413,N_8642,N_9247);
nor U12414 (N_12414,N_9498,N_8143);
nand U12415 (N_12415,N_10695,N_10067);
or U12416 (N_12416,N_10711,N_8260);
nand U12417 (N_12417,N_9889,N_9598);
or U12418 (N_12418,N_8624,N_9477);
xor U12419 (N_12419,N_10764,N_9323);
and U12420 (N_12420,N_9698,N_9375);
nor U12421 (N_12421,N_8789,N_9782);
and U12422 (N_12422,N_8434,N_8630);
or U12423 (N_12423,N_8235,N_10968);
or U12424 (N_12424,N_9045,N_11843);
nand U12425 (N_12425,N_10645,N_8042);
and U12426 (N_12426,N_9567,N_9775);
and U12427 (N_12427,N_9306,N_11076);
nor U12428 (N_12428,N_8649,N_9317);
xor U12429 (N_12429,N_10657,N_8834);
and U12430 (N_12430,N_8665,N_11822);
nor U12431 (N_12431,N_11970,N_11505);
and U12432 (N_12432,N_10662,N_11809);
nand U12433 (N_12433,N_11825,N_11275);
or U12434 (N_12434,N_8782,N_8969);
or U12435 (N_12435,N_9982,N_11075);
nor U12436 (N_12436,N_8356,N_8189);
and U12437 (N_12437,N_8973,N_9359);
and U12438 (N_12438,N_8655,N_10654);
and U12439 (N_12439,N_8865,N_11776);
xnor U12440 (N_12440,N_11048,N_10752);
nand U12441 (N_12441,N_8152,N_9385);
nor U12442 (N_12442,N_9050,N_8126);
nand U12443 (N_12443,N_11282,N_8586);
nor U12444 (N_12444,N_11135,N_10946);
nand U12445 (N_12445,N_11956,N_11800);
nand U12446 (N_12446,N_10163,N_11785);
nand U12447 (N_12447,N_11870,N_10047);
or U12448 (N_12448,N_10375,N_11580);
xnor U12449 (N_12449,N_10235,N_11358);
and U12450 (N_12450,N_11657,N_9240);
nand U12451 (N_12451,N_9021,N_10393);
nand U12452 (N_12452,N_11890,N_10299);
nand U12453 (N_12453,N_8187,N_10922);
nand U12454 (N_12454,N_9523,N_11022);
nor U12455 (N_12455,N_10828,N_11086);
nor U12456 (N_12456,N_11714,N_8440);
and U12457 (N_12457,N_8608,N_11417);
nand U12458 (N_12458,N_11755,N_8570);
and U12459 (N_12459,N_9921,N_9025);
nor U12460 (N_12460,N_9577,N_9273);
and U12461 (N_12461,N_9362,N_10350);
and U12462 (N_12462,N_10306,N_9674);
xnor U12463 (N_12463,N_8357,N_8261);
nor U12464 (N_12464,N_10202,N_10904);
nor U12465 (N_12465,N_11692,N_10651);
or U12466 (N_12466,N_11290,N_9511);
or U12467 (N_12467,N_10392,N_8661);
nand U12468 (N_12468,N_8395,N_10478);
and U12469 (N_12469,N_10095,N_8084);
xnor U12470 (N_12470,N_8306,N_10775);
nor U12471 (N_12471,N_10827,N_8231);
or U12472 (N_12472,N_11241,N_11248);
or U12473 (N_12473,N_9784,N_11049);
or U12474 (N_12474,N_10335,N_11051);
and U12475 (N_12475,N_9172,N_11376);
and U12476 (N_12476,N_8836,N_10185);
and U12477 (N_12477,N_11715,N_10232);
nor U12478 (N_12478,N_8266,N_9309);
and U12479 (N_12479,N_10964,N_9461);
nor U12480 (N_12480,N_8859,N_8374);
nor U12481 (N_12481,N_8381,N_10174);
nor U12482 (N_12482,N_9446,N_9879);
nor U12483 (N_12483,N_10468,N_9017);
and U12484 (N_12484,N_11882,N_9753);
or U12485 (N_12485,N_11979,N_8849);
and U12486 (N_12486,N_10691,N_8947);
nand U12487 (N_12487,N_10846,N_11868);
nand U12488 (N_12488,N_10217,N_9787);
and U12489 (N_12489,N_9342,N_9571);
nand U12490 (N_12490,N_9778,N_11130);
and U12491 (N_12491,N_10024,N_8132);
nor U12492 (N_12492,N_11677,N_9378);
nand U12493 (N_12493,N_8142,N_11513);
xor U12494 (N_12494,N_10999,N_8024);
nand U12495 (N_12495,N_10698,N_11422);
or U12496 (N_12496,N_8659,N_10377);
xnor U12497 (N_12497,N_8740,N_11667);
xnor U12498 (N_12498,N_9020,N_8530);
or U12499 (N_12499,N_10777,N_10379);
nand U12500 (N_12500,N_10545,N_9391);
and U12501 (N_12501,N_10181,N_9227);
nand U12502 (N_12502,N_11060,N_10866);
or U12503 (N_12503,N_10977,N_9134);
nand U12504 (N_12504,N_9740,N_10589);
nor U12505 (N_12505,N_9962,N_8671);
nor U12506 (N_12506,N_11891,N_11842);
nor U12507 (N_12507,N_10255,N_10463);
or U12508 (N_12508,N_9250,N_11070);
nand U12509 (N_12509,N_9497,N_11836);
and U12510 (N_12510,N_11668,N_9041);
or U12511 (N_12511,N_10167,N_10721);
and U12512 (N_12512,N_9583,N_11814);
and U12513 (N_12513,N_9440,N_11054);
or U12514 (N_12514,N_9033,N_9403);
xor U12515 (N_12515,N_8172,N_9833);
or U12516 (N_12516,N_10336,N_8410);
nor U12517 (N_12517,N_9120,N_9996);
or U12518 (N_12518,N_10732,N_10700);
and U12519 (N_12519,N_10094,N_10816);
or U12520 (N_12520,N_9076,N_11133);
xnor U12521 (N_12521,N_11008,N_11471);
and U12522 (N_12522,N_8344,N_8662);
nor U12523 (N_12523,N_10277,N_9957);
xnor U12524 (N_12524,N_9734,N_9476);
nand U12525 (N_12525,N_11121,N_9636);
or U12526 (N_12526,N_11194,N_10933);
nand U12527 (N_12527,N_10180,N_10348);
or U12528 (N_12528,N_9248,N_8340);
and U12529 (N_12529,N_11948,N_11073);
and U12530 (N_12530,N_11634,N_8462);
or U12531 (N_12531,N_9768,N_9453);
xnor U12532 (N_12532,N_10233,N_9448);
nand U12533 (N_12533,N_10789,N_10097);
and U12534 (N_12534,N_9409,N_8311);
xor U12535 (N_12535,N_8198,N_11899);
nand U12536 (N_12536,N_9504,N_10753);
and U12537 (N_12537,N_11472,N_9329);
nand U12538 (N_12538,N_8159,N_8516);
nor U12539 (N_12539,N_9009,N_10617);
or U12540 (N_12540,N_9781,N_8317);
nor U12541 (N_12541,N_11255,N_10622);
and U12542 (N_12542,N_8480,N_11044);
nor U12543 (N_12543,N_8035,N_8606);
or U12544 (N_12544,N_9902,N_11403);
xor U12545 (N_12545,N_9903,N_10435);
nor U12546 (N_12546,N_8039,N_11558);
nand U12547 (N_12547,N_8622,N_9263);
nor U12548 (N_12548,N_10659,N_9974);
or U12549 (N_12549,N_11025,N_10308);
xor U12550 (N_12550,N_11071,N_11739);
nor U12551 (N_12551,N_10992,N_9737);
xor U12552 (N_12552,N_11921,N_9465);
nand U12553 (N_12553,N_9788,N_11372);
nor U12554 (N_12554,N_8294,N_8379);
nand U12555 (N_12555,N_10840,N_10895);
xnor U12556 (N_12556,N_11576,N_11864);
nand U12557 (N_12557,N_8677,N_11614);
or U12558 (N_12558,N_8986,N_9103);
nor U12559 (N_12559,N_11306,N_11627);
nand U12560 (N_12560,N_8612,N_9369);
or U12561 (N_12561,N_11247,N_11512);
or U12562 (N_12562,N_8080,N_11902);
nor U12563 (N_12563,N_10784,N_8526);
or U12564 (N_12564,N_11126,N_9402);
nor U12565 (N_12565,N_10327,N_9601);
nor U12566 (N_12566,N_11438,N_9395);
nor U12567 (N_12567,N_10251,N_9335);
nand U12568 (N_12568,N_8644,N_9611);
or U12569 (N_12569,N_8775,N_8323);
and U12570 (N_12570,N_9896,N_8438);
xor U12571 (N_12571,N_8989,N_8394);
or U12572 (N_12572,N_11159,N_11774);
nor U12573 (N_12573,N_9308,N_9260);
nand U12574 (N_12574,N_11590,N_8974);
or U12575 (N_12575,N_11383,N_10834);
nor U12576 (N_12576,N_9014,N_10523);
nand U12577 (N_12577,N_9552,N_10122);
nand U12578 (N_12578,N_11445,N_9542);
or U12579 (N_12579,N_10884,N_10118);
nand U12580 (N_12580,N_8905,N_9416);
nor U12581 (N_12581,N_11607,N_8269);
nor U12582 (N_12582,N_10338,N_9642);
nor U12583 (N_12583,N_11609,N_9976);
xnor U12584 (N_12584,N_9762,N_10326);
nand U12585 (N_12585,N_8048,N_8509);
nand U12586 (N_12586,N_8114,N_10526);
or U12587 (N_12587,N_11732,N_9710);
nor U12588 (N_12588,N_11172,N_10456);
and U12589 (N_12589,N_10442,N_11435);
nor U12590 (N_12590,N_11645,N_9969);
nand U12591 (N_12591,N_10162,N_9056);
or U12592 (N_12592,N_11448,N_10329);
and U12593 (N_12593,N_11443,N_9890);
or U12594 (N_12594,N_9715,N_10974);
nor U12595 (N_12595,N_8490,N_8566);
or U12596 (N_12596,N_10759,N_10397);
nor U12597 (N_12597,N_10737,N_10520);
or U12598 (N_12598,N_11203,N_11066);
and U12599 (N_12599,N_10290,N_8871);
nor U12600 (N_12600,N_9893,N_11256);
nand U12601 (N_12601,N_10360,N_9249);
nor U12602 (N_12602,N_11334,N_11065);
or U12603 (N_12603,N_8603,N_8497);
nand U12604 (N_12604,N_9625,N_11257);
or U12605 (N_12605,N_9652,N_9995);
nand U12606 (N_12606,N_8397,N_9815);
nor U12607 (N_12607,N_8592,N_8170);
and U12608 (N_12608,N_11557,N_9364);
xnor U12609 (N_12609,N_11985,N_11234);
and U12610 (N_12610,N_8890,N_8954);
or U12611 (N_12611,N_9324,N_9168);
and U12612 (N_12612,N_10658,N_11035);
nor U12613 (N_12613,N_9729,N_10595);
and U12614 (N_12614,N_10742,N_10250);
or U12615 (N_12615,N_11420,N_10856);
or U12616 (N_12616,N_10316,N_10005);
or U12617 (N_12617,N_9681,N_9221);
and U12618 (N_12618,N_9049,N_11218);
nand U12619 (N_12619,N_11494,N_10920);
or U12620 (N_12620,N_11589,N_9973);
nand U12621 (N_12621,N_8788,N_8343);
nor U12622 (N_12622,N_8334,N_11037);
or U12623 (N_12623,N_10802,N_11940);
nand U12624 (N_12624,N_11502,N_11759);
nor U12625 (N_12625,N_11014,N_10425);
and U12626 (N_12626,N_9596,N_11318);
nand U12627 (N_12627,N_8108,N_8427);
and U12628 (N_12628,N_10630,N_8984);
or U12629 (N_12629,N_10845,N_9657);
or U12630 (N_12630,N_8551,N_8869);
or U12631 (N_12631,N_8404,N_9267);
or U12632 (N_12632,N_8912,N_10852);
or U12633 (N_12633,N_10580,N_11361);
or U12634 (N_12634,N_8154,N_10439);
nand U12635 (N_12635,N_10748,N_11423);
nand U12636 (N_12636,N_9855,N_9914);
and U12637 (N_12637,N_10517,N_9829);
and U12638 (N_12638,N_10538,N_10459);
xor U12639 (N_12639,N_9572,N_11313);
xor U12640 (N_12640,N_10971,N_11584);
and U12641 (N_12641,N_11545,N_10150);
nor U12642 (N_12642,N_8978,N_10105);
xor U12643 (N_12643,N_8870,N_9548);
and U12644 (N_12644,N_11998,N_10592);
nor U12645 (N_12645,N_10035,N_8626);
xnor U12646 (N_12646,N_8333,N_8525);
xor U12647 (N_12647,N_10135,N_11651);
xnor U12648 (N_12648,N_10586,N_11989);
and U12649 (N_12649,N_9090,N_11260);
and U12650 (N_12650,N_10530,N_10499);
nor U12651 (N_12651,N_10744,N_8431);
nand U12652 (N_12652,N_11855,N_8240);
nand U12653 (N_12653,N_10931,N_11293);
nand U12654 (N_12654,N_8877,N_8922);
nor U12655 (N_12655,N_11716,N_9941);
nor U12656 (N_12656,N_8498,N_8382);
or U12657 (N_12657,N_11904,N_8997);
or U12658 (N_12658,N_8388,N_11151);
and U12659 (N_12659,N_11173,N_10607);
nor U12660 (N_12660,N_11758,N_10534);
nor U12661 (N_12661,N_10927,N_10686);
nand U12662 (N_12662,N_9952,N_9154);
or U12663 (N_12663,N_11458,N_8596);
xnor U12664 (N_12664,N_10028,N_9000);
nor U12665 (N_12665,N_8879,N_8852);
nor U12666 (N_12666,N_10305,N_10193);
xor U12667 (N_12667,N_9457,N_9865);
nor U12668 (N_12668,N_10331,N_11338);
nor U12669 (N_12669,N_8064,N_8243);
or U12670 (N_12670,N_8628,N_8862);
nand U12671 (N_12671,N_11165,N_10258);
xnor U12672 (N_12672,N_9096,N_11487);
xor U12673 (N_12673,N_11138,N_10668);
nor U12674 (N_12674,N_11215,N_10453);
or U12675 (N_12675,N_8214,N_11270);
nor U12676 (N_12676,N_9285,N_10648);
or U12677 (N_12677,N_10406,N_8892);
and U12678 (N_12678,N_10139,N_10378);
and U12679 (N_12679,N_9938,N_9915);
or U12680 (N_12680,N_11528,N_10133);
and U12681 (N_12681,N_9312,N_8282);
nand U12682 (N_12682,N_11092,N_10547);
or U12683 (N_12683,N_11465,N_9679);
or U12684 (N_12684,N_11479,N_11833);
or U12685 (N_12685,N_10824,N_8676);
nor U12686 (N_12686,N_11717,N_11093);
and U12687 (N_12687,N_11392,N_8830);
nand U12688 (N_12688,N_10751,N_8043);
and U12689 (N_12689,N_10666,N_8138);
xor U12690 (N_12690,N_9083,N_8325);
nor U12691 (N_12691,N_11876,N_8016);
nor U12692 (N_12692,N_9966,N_8370);
nand U12693 (N_12693,N_11885,N_8880);
or U12694 (N_12694,N_9888,N_9852);
nor U12695 (N_12695,N_9222,N_9418);
and U12696 (N_12696,N_9361,N_8742);
nand U12697 (N_12697,N_10142,N_9209);
nor U12698 (N_12698,N_10112,N_10629);
or U12699 (N_12699,N_10725,N_8972);
and U12700 (N_12700,N_8695,N_11108);
nand U12701 (N_12701,N_11624,N_8557);
or U12702 (N_12702,N_10584,N_11641);
or U12703 (N_12703,N_9205,N_8355);
nand U12704 (N_12704,N_11728,N_9700);
and U12705 (N_12705,N_10609,N_9449);
or U12706 (N_12706,N_10678,N_11139);
nor U12707 (N_12707,N_9165,N_8706);
xor U12708 (N_12708,N_8991,N_11688);
nor U12709 (N_12709,N_9936,N_10942);
or U12710 (N_12710,N_10152,N_11179);
xnor U12711 (N_12711,N_9809,N_11698);
xor U12712 (N_12712,N_8476,N_8310);
nand U12713 (N_12713,N_10875,N_10917);
nand U12714 (N_12714,N_10722,N_8297);
nor U12715 (N_12715,N_9637,N_10527);
nor U12716 (N_12716,N_11996,N_9856);
nand U12717 (N_12717,N_10792,N_10477);
nand U12718 (N_12718,N_8101,N_8123);
or U12719 (N_12719,N_10932,N_11887);
and U12720 (N_12720,N_11228,N_8184);
xnor U12721 (N_12721,N_11027,N_9386);
and U12722 (N_12722,N_10461,N_10187);
xor U12723 (N_12723,N_9720,N_8362);
nand U12724 (N_12724,N_9770,N_8047);
and U12725 (N_12725,N_9191,N_11660);
nor U12726 (N_12726,N_10685,N_8609);
xnor U12727 (N_12727,N_8219,N_10243);
or U12728 (N_12728,N_10050,N_9360);
or U12729 (N_12729,N_8511,N_11784);
nor U12730 (N_12730,N_10497,N_10669);
nor U12731 (N_12731,N_11208,N_9383);
and U12732 (N_12732,N_8696,N_10650);
nand U12733 (N_12733,N_9942,N_11123);
and U12734 (N_12734,N_10779,N_8529);
nand U12735 (N_12735,N_11253,N_10405);
and U12736 (N_12736,N_11783,N_8400);
nor U12737 (N_12737,N_11389,N_10647);
xnor U12738 (N_12738,N_11230,N_11949);
nor U12739 (N_12739,N_9521,N_8857);
and U12740 (N_12740,N_9595,N_10806);
or U12741 (N_12741,N_11170,N_11197);
nand U12742 (N_12742,N_10169,N_11231);
xnor U12743 (N_12743,N_8501,N_8464);
or U12744 (N_12744,N_10491,N_11813);
and U12745 (N_12745,N_11090,N_11454);
or U12746 (N_12746,N_10771,N_10991);
nor U12747 (N_12747,N_11939,N_11803);
nor U12748 (N_12748,N_10536,N_8716);
or U12749 (N_12749,N_11031,N_11474);
or U12750 (N_12750,N_9745,N_8505);
nand U12751 (N_12751,N_8667,N_9142);
nand U12752 (N_12752,N_10882,N_10786);
and U12753 (N_12753,N_10474,N_9534);
or U12754 (N_12754,N_11623,N_11103);
nor U12755 (N_12755,N_8995,N_8726);
or U12756 (N_12756,N_10029,N_8908);
and U12757 (N_12757,N_8928,N_11879);
nor U12758 (N_12758,N_9807,N_10494);
nand U12759 (N_12759,N_10893,N_9073);
nor U12760 (N_12760,N_11865,N_11625);
nor U12761 (N_12761,N_10470,N_10661);
and U12762 (N_12762,N_11192,N_8783);
nand U12763 (N_12763,N_10370,N_8060);
nand U12764 (N_12764,N_10785,N_11567);
nand U12765 (N_12765,N_8276,N_9038);
nand U12766 (N_12766,N_8689,N_8723);
and U12767 (N_12767,N_9203,N_9800);
nand U12768 (N_12768,N_10502,N_11081);
nand U12769 (N_12769,N_8528,N_8545);
nand U12770 (N_12770,N_8493,N_10569);
or U12771 (N_12771,N_8878,N_11476);
xnor U12772 (N_12772,N_10485,N_9765);
nor U12773 (N_12773,N_9631,N_8283);
or U12774 (N_12774,N_10770,N_9424);
nor U12775 (N_12775,N_11773,N_9430);
and U12776 (N_12776,N_11824,N_10063);
nor U12777 (N_12777,N_10699,N_10663);
or U12778 (N_12778,N_10080,N_9015);
or U12779 (N_12779,N_9301,N_9661);
or U12780 (N_12780,N_9198,N_10763);
nand U12781 (N_12781,N_11764,N_8456);
and U12782 (N_12782,N_8383,N_10374);
nor U12783 (N_12783,N_9133,N_10419);
nand U12784 (N_12784,N_10347,N_11493);
nor U12785 (N_12785,N_11907,N_9712);
and U12786 (N_12786,N_10544,N_8710);
nand U12787 (N_12787,N_10391,N_9822);
or U12788 (N_12788,N_10146,N_10898);
xnor U12789 (N_12789,N_9158,N_8523);
or U12790 (N_12790,N_9112,N_8934);
nor U12791 (N_12791,N_11520,N_11867);
nor U12792 (N_12792,N_9771,N_8158);
nor U12793 (N_12793,N_9823,N_10165);
and U12794 (N_12794,N_8962,N_11074);
nor U12795 (N_12795,N_8091,N_8166);
and U12796 (N_12796,N_9585,N_11164);
or U12797 (N_12797,N_9482,N_10333);
or U12798 (N_12798,N_9094,N_9419);
or U12799 (N_12799,N_8280,N_9748);
nor U12800 (N_12800,N_9519,N_9858);
nor U12801 (N_12801,N_8453,N_9356);
nor U12802 (N_12802,N_8403,N_10637);
nor U12803 (N_12803,N_8203,N_10197);
or U12804 (N_12804,N_10978,N_9212);
and U12805 (N_12805,N_10857,N_9866);
or U12806 (N_12806,N_11982,N_11880);
and U12807 (N_12807,N_8392,N_10718);
and U12808 (N_12808,N_9174,N_8882);
nand U12809 (N_12809,N_9717,N_9143);
nand U12810 (N_12810,N_9786,N_11452);
and U12811 (N_12811,N_10762,N_10015);
or U12812 (N_12812,N_8157,N_10638);
nand U12813 (N_12813,N_10510,N_10597);
and U12814 (N_12814,N_9876,N_11782);
or U12815 (N_12815,N_10452,N_11272);
nand U12816 (N_12816,N_8844,N_8965);
nand U12817 (N_12817,N_11936,N_8886);
nor U12818 (N_12818,N_10664,N_10295);
nand U12819 (N_12819,N_11114,N_9468);
nor U12820 (N_12820,N_9517,N_9450);
and U12821 (N_12821,N_9293,N_10207);
nor U12822 (N_12822,N_11595,N_8371);
and U12823 (N_12823,N_10102,N_11371);
and U12824 (N_12824,N_8835,N_11153);
and U12825 (N_12825,N_10208,N_8082);
nand U12826 (N_12826,N_8248,N_11655);
nand U12827 (N_12827,N_11652,N_8234);
nor U12828 (N_12828,N_11612,N_10088);
nand U12829 (N_12829,N_10205,N_10141);
nor U12830 (N_12830,N_8121,N_11514);
nand U12831 (N_12831,N_11053,N_9798);
nand U12832 (N_12832,N_8414,N_11808);
or U12833 (N_12833,N_11640,N_8718);
and U12834 (N_12834,N_9774,N_11155);
and U12835 (N_12835,N_10943,N_8654);
nand U12836 (N_12836,N_10039,N_9414);
and U12837 (N_12837,N_9139,N_11945);
or U12838 (N_12838,N_9489,N_11602);
and U12839 (N_12839,N_11375,N_10194);
nand U12840 (N_12840,N_10563,N_11309);
nand U12841 (N_12841,N_9443,N_11146);
and U12842 (N_12842,N_10062,N_8737);
nor U12843 (N_12843,N_11778,N_11469);
and U12844 (N_12844,N_11831,N_11168);
xor U12845 (N_12845,N_11245,N_11265);
nand U12846 (N_12846,N_11296,N_10915);
nand U12847 (N_12847,N_9756,N_10364);
and U12848 (N_12848,N_9051,N_8924);
or U12849 (N_12849,N_10707,N_8921);
xor U12850 (N_12850,N_8314,N_11615);
or U12851 (N_12851,N_11964,N_8012);
nand U12852 (N_12852,N_10283,N_10633);
and U12853 (N_12853,N_9490,N_10076);
xor U12854 (N_12854,N_9307,N_10772);
nand U12855 (N_12855,N_11284,N_8197);
nand U12856 (N_12856,N_11488,N_11077);
or U12857 (N_12857,N_11839,N_11149);
or U12858 (N_12858,N_10767,N_8353);
nor U12859 (N_12859,N_10231,N_9690);
and U12860 (N_12860,N_11292,N_11527);
nor U12861 (N_12861,N_9868,N_8639);
and U12862 (N_12862,N_11294,N_9458);
xor U12863 (N_12863,N_10382,N_8331);
nand U12864 (N_12864,N_8633,N_8842);
nand U12865 (N_12865,N_10066,N_10221);
or U12866 (N_12866,N_11182,N_10403);
xor U12867 (N_12867,N_9863,N_8063);
nand U12868 (N_12868,N_10549,N_10954);
or U12869 (N_12869,N_8120,N_10768);
and U12870 (N_12870,N_8075,N_10268);
and U12871 (N_12871,N_11004,N_9337);
nor U12872 (N_12872,N_8182,N_8322);
nor U12873 (N_12873,N_11367,N_11143);
or U12874 (N_12874,N_9623,N_10060);
and U12875 (N_12875,N_11163,N_8697);
nor U12876 (N_12876,N_10164,N_9546);
nand U12877 (N_12877,N_8051,N_8342);
or U12878 (N_12878,N_9513,N_9886);
nand U12879 (N_12879,N_9217,N_10224);
nor U12880 (N_12880,N_8699,N_8139);
and U12881 (N_12881,N_10110,N_8810);
nand U12882 (N_12882,N_10457,N_8646);
nand U12883 (N_12883,N_9835,N_9557);
nand U12884 (N_12884,N_9706,N_10318);
nand U12885 (N_12885,N_9989,N_11850);
nor U12886 (N_12886,N_10006,N_8552);
nor U12887 (N_12887,N_11735,N_11212);
nand U12888 (N_12888,N_10021,N_11483);
nand U12889 (N_12889,N_8801,N_10903);
and U12890 (N_12890,N_9321,N_10411);
nor U12891 (N_12891,N_10506,N_9684);
or U12892 (N_12892,N_8985,N_10706);
and U12893 (N_12893,N_8913,N_11926);
or U12894 (N_12894,N_11737,N_11877);
and U12895 (N_12895,N_9431,N_9164);
or U12896 (N_12896,N_8771,N_10444);
xor U12897 (N_12897,N_10440,N_8795);
or U12898 (N_12898,N_11633,N_10734);
xnor U12899 (N_12899,N_11910,N_10246);
and U12900 (N_12900,N_9008,N_9656);
xor U12901 (N_12901,N_9243,N_8899);
or U12902 (N_12902,N_10897,N_9487);
and U12903 (N_12903,N_9368,N_11517);
nor U12904 (N_12904,N_10161,N_9367);
and U12905 (N_12905,N_9208,N_11571);
or U12906 (N_12906,N_10003,N_9231);
nor U12907 (N_12907,N_11005,N_8720);
or U12908 (N_12908,N_9935,N_9380);
xnor U12909 (N_12909,N_9183,N_8146);
and U12910 (N_12910,N_11894,N_9533);
nand U12911 (N_12911,N_9574,N_10395);
and U12912 (N_12912,N_9210,N_11709);
or U12913 (N_12913,N_8688,N_9887);
nor U12914 (N_12914,N_10849,N_11412);
and U12915 (N_12915,N_8098,N_9683);
nand U12916 (N_12916,N_9322,N_8817);
nand U12917 (N_12917,N_9695,N_8847);
xor U12918 (N_12918,N_11229,N_10014);
nor U12919 (N_12919,N_9054,N_10871);
and U12920 (N_12920,N_8837,N_11853);
and U12921 (N_12921,N_10022,N_11930);
nor U12922 (N_12922,N_8961,N_11018);
and U12923 (N_12923,N_8918,N_9672);
nand U12924 (N_12924,N_9588,N_11111);
nor U12925 (N_12925,N_11028,N_10906);
nand U12926 (N_12926,N_8281,N_9949);
nand U12927 (N_12927,N_10293,N_8568);
nor U12928 (N_12928,N_10106,N_10821);
nor U12929 (N_12929,N_10279,N_10902);
xor U12930 (N_12930,N_8893,N_8620);
and U12931 (N_12931,N_8301,N_9609);
and U12932 (N_12932,N_8749,N_8273);
nor U12933 (N_12933,N_8022,N_11917);
nor U12934 (N_12934,N_8290,N_11554);
or U12935 (N_12935,N_11336,N_9872);
nand U12936 (N_12936,N_8324,N_10323);
or U12937 (N_12937,N_10987,N_9834);
and U12938 (N_12938,N_9743,N_8315);
or U12939 (N_12939,N_8391,N_11760);
xor U12940 (N_12940,N_9711,N_8129);
and U12941 (N_12941,N_8935,N_11972);
nand U12942 (N_12942,N_11395,N_8787);
and U12943 (N_12943,N_10934,N_11574);
or U12944 (N_12944,N_8998,N_8602);
xor U12945 (N_12945,N_10955,N_11563);
and U12946 (N_12946,N_9271,N_11310);
xnor U12947 (N_12947,N_8034,N_9714);
nor U12948 (N_12948,N_11366,N_9130);
nand U12949 (N_12949,N_8549,N_11083);
xor U12950 (N_12950,N_11560,N_11659);
or U12951 (N_12951,N_9343,N_10525);
nor U12952 (N_12952,N_9254,N_10649);
and U12953 (N_12953,N_10874,N_10438);
and U12954 (N_12954,N_9713,N_9847);
nand U12955 (N_12955,N_11484,N_10143);
nand U12956 (N_12956,N_8096,N_9937);
nor U12957 (N_12957,N_9085,N_11561);
xnor U12958 (N_12958,N_11064,N_11384);
nor U12959 (N_12959,N_8369,N_8406);
nand U12960 (N_12960,N_8687,N_11960);
and U12961 (N_12961,N_11017,N_11411);
and U12962 (N_12962,N_8443,N_10984);
nor U12963 (N_12963,N_10158,N_9563);
and U12964 (N_12964,N_8513,N_8446);
xor U12965 (N_12965,N_10498,N_9971);
and U12966 (N_12966,N_11961,N_9202);
nand U12967 (N_12967,N_10324,N_9900);
xnor U12968 (N_12968,N_10941,N_11938);
xnor U12969 (N_12969,N_11726,N_9415);
nand U12970 (N_12970,N_9175,N_10034);
nand U12971 (N_12971,N_8809,N_8534);
nand U12972 (N_12972,N_9189,N_8033);
and U12973 (N_12973,N_11957,N_8103);
or U12974 (N_12974,N_8930,N_9669);
nor U12975 (N_12975,N_10869,N_10508);
xor U12976 (N_12976,N_11431,N_11719);
and U12977 (N_12977,N_9155,N_8519);
nand U12978 (N_12978,N_8337,N_11152);
and U12979 (N_12979,N_9528,N_10565);
or U12980 (N_12980,N_9662,N_10325);
nand U12981 (N_12981,N_9400,N_8572);
nor U12982 (N_12982,N_9685,N_10481);
nor U12983 (N_12983,N_8730,N_8107);
and U12984 (N_12984,N_11470,N_10473);
and U12985 (N_12985,N_9053,N_11437);
nand U12986 (N_12986,N_10925,N_8106);
or U12987 (N_12987,N_10320,N_8804);
and U12988 (N_12988,N_10808,N_10449);
nand U12989 (N_12989,N_9606,N_10947);
xnor U12990 (N_12990,N_10512,N_11680);
xor U12991 (N_12991,N_8253,N_11396);
nand U12992 (N_12992,N_11588,N_10177);
and U12993 (N_12993,N_9381,N_10079);
nor U12994 (N_12994,N_10600,N_9107);
or U12995 (N_12995,N_9584,N_10228);
or U12996 (N_12996,N_11174,N_10855);
or U12997 (N_12997,N_10433,N_9007);
or U12998 (N_12998,N_8599,N_8786);
or U12999 (N_12999,N_8770,N_11738);
xnor U13000 (N_13000,N_9998,N_11582);
and U13001 (N_13001,N_10504,N_11394);
nor U13002 (N_13002,N_9411,N_9279);
nor U13003 (N_13003,N_8684,N_11080);
nor U13004 (N_13004,N_11526,N_10909);
and U13005 (N_13005,N_11540,N_10842);
and U13006 (N_13006,N_8177,N_9610);
and U13007 (N_13007,N_10002,N_8700);
and U13008 (N_13008,N_8477,N_10413);
and U13009 (N_13009,N_9959,N_10178);
nand U13010 (N_13010,N_8233,N_10307);
nand U13011 (N_13011,N_11308,N_11628);
or U13012 (N_13012,N_9954,N_8994);
nor U13013 (N_13013,N_10140,N_9266);
or U13014 (N_13014,N_8562,N_8867);
nand U13015 (N_13015,N_10493,N_10930);
nor U13016 (N_13016,N_9159,N_9627);
nor U13017 (N_13017,N_11285,N_8496);
xor U13018 (N_13018,N_11510,N_10204);
nand U13019 (N_13019,N_10188,N_11118);
or U13020 (N_13020,N_9553,N_8286);
nand U13021 (N_13021,N_9261,N_8483);
nor U13022 (N_13022,N_8951,N_10061);
nand U13023 (N_13023,N_11638,N_10881);
nand U13024 (N_13024,N_11787,N_11770);
nor U13025 (N_13025,N_10936,N_9839);
and U13026 (N_13026,N_8611,N_10797);
and U13027 (N_13027,N_10982,N_8738);
and U13028 (N_13028,N_11844,N_9067);
or U13029 (N_13029,N_10056,N_9961);
or U13030 (N_13030,N_11592,N_11119);
or U13031 (N_13031,N_8402,N_8461);
nand U13032 (N_13032,N_11205,N_10796);
or U13033 (N_13033,N_8517,N_10495);
nand U13034 (N_13034,N_11112,N_8681);
nor U13035 (N_13035,N_10332,N_11425);
and U13036 (N_13036,N_9968,N_10631);
or U13037 (N_13037,N_8463,N_9527);
xnor U13038 (N_13038,N_9722,N_10747);
nand U13039 (N_13039,N_11145,N_10750);
and U13040 (N_13040,N_9923,N_10211);
nor U13041 (N_13041,N_9149,N_11756);
or U13042 (N_13042,N_8386,N_11817);
or U13043 (N_13043,N_10201,N_11419);
and U13044 (N_13044,N_9597,N_11838);
nor U13045 (N_13045,N_9485,N_10400);
and U13046 (N_13046,N_11873,N_10240);
nand U13047 (N_13047,N_11674,N_9794);
and U13048 (N_13048,N_11274,N_8279);
nor U13049 (N_13049,N_8904,N_8377);
or U13050 (N_13050,N_9152,N_10953);
and U13051 (N_13051,N_10551,N_10673);
nand U13052 (N_13052,N_9206,N_11244);
or U13053 (N_13053,N_9433,N_11029);
or U13054 (N_13054,N_11621,N_8637);
nor U13055 (N_13055,N_11357,N_9475);
nor U13056 (N_13056,N_8823,N_9592);
or U13057 (N_13057,N_10070,N_9842);
nor U13058 (N_13058,N_11043,N_8115);
or U13059 (N_13059,N_8263,N_10261);
nand U13060 (N_13060,N_10812,N_9148);
or U13061 (N_13061,N_9814,N_10108);
nor U13062 (N_13062,N_11106,N_9817);
and U13063 (N_13063,N_11830,N_9934);
nor U13064 (N_13064,N_8105,N_8754);
or U13065 (N_13065,N_11820,N_11794);
nand U13066 (N_13066,N_9351,N_10365);
xor U13067 (N_13067,N_11821,N_10843);
nor U13068 (N_13068,N_8217,N_11974);
xor U13069 (N_13069,N_9026,N_10921);
and U13070 (N_13070,N_10078,N_9022);
and U13071 (N_13071,N_11925,N_9413);
nand U13072 (N_13072,N_10626,N_11097);
nand U13073 (N_13073,N_11712,N_8731);
nor U13074 (N_13074,N_11525,N_8883);
and U13075 (N_13075,N_10043,N_10137);
and U13076 (N_13076,N_11578,N_11317);
nor U13077 (N_13077,N_9147,N_9146);
or U13078 (N_13078,N_8527,N_10418);
and U13079 (N_13079,N_10899,N_9749);
or U13080 (N_13080,N_8800,N_10239);
nor U13081 (N_13081,N_9844,N_9721);
and U13082 (N_13082,N_10778,N_9048);
and U13083 (N_13083,N_10552,N_9398);
xnor U13084 (N_13084,N_9806,N_10864);
or U13085 (N_13085,N_8305,N_11733);
xnor U13086 (N_13086,N_11829,N_11549);
or U13087 (N_13087,N_8868,N_11261);
nor U13088 (N_13088,N_8482,N_11177);
or U13089 (N_13089,N_11131,N_11761);
and U13090 (N_13090,N_8860,N_11909);
and U13091 (N_13091,N_11332,N_8435);
nand U13092 (N_13092,N_10209,N_8752);
and U13093 (N_13093,N_8811,N_8225);
and U13094 (N_13094,N_11397,N_10260);
nor U13095 (N_13095,N_11300,N_10588);
nand U13096 (N_13096,N_11141,N_9566);
and U13097 (N_13097,N_11342,N_10467);
and U13098 (N_13098,N_10480,N_10972);
nand U13099 (N_13099,N_11286,N_10443);
nand U13100 (N_13100,N_8722,N_8569);
or U13101 (N_13101,N_11919,N_9473);
or U13102 (N_13102,N_9105,N_9578);
nand U13103 (N_13103,N_9813,N_10212);
xnor U13104 (N_13104,N_9072,N_10253);
or U13105 (N_13105,N_10183,N_8321);
or U13106 (N_13106,N_9091,N_8023);
nor U13107 (N_13107,N_10585,N_10273);
or U13108 (N_13108,N_9692,N_11455);
nor U13109 (N_13109,N_9126,N_10203);
nor U13110 (N_13110,N_10275,N_8238);
nor U13111 (N_13111,N_11434,N_11975);
xnor U13112 (N_13112,N_9084,N_9644);
xor U13113 (N_13113,N_8721,N_8508);
nor U13114 (N_13114,N_10590,N_11032);
nand U13115 (N_13115,N_9967,N_8265);
or U13116 (N_13116,N_11648,N_10234);
nand U13117 (N_13117,N_10848,N_9075);
nor U13118 (N_13118,N_8573,N_8466);
xor U13119 (N_13119,N_8719,N_9626);
and U13120 (N_13120,N_11644,N_9062);
nand U13121 (N_13121,N_8112,N_8729);
and U13122 (N_13122,N_9123,N_9950);
nor U13123 (N_13123,N_9639,N_10956);
nor U13124 (N_13124,N_8873,N_11137);
or U13125 (N_13125,N_10341,N_10603);
nand U13126 (N_13126,N_9161,N_9620);
or U13127 (N_13127,N_11804,N_11441);
nand U13128 (N_13128,N_9953,N_8590);
and U13129 (N_13129,N_9931,N_8983);
xor U13130 (N_13130,N_8256,N_9405);
nand U13131 (N_13131,N_11933,N_11072);
nand U13132 (N_13132,N_8007,N_9673);
and U13133 (N_13133,N_10542,N_11931);
nor U13134 (N_13134,N_8668,N_8504);
nor U13135 (N_13135,N_9666,N_10252);
nor U13136 (N_13136,N_11006,N_10887);
and U13137 (N_13137,N_11675,N_10111);
or U13138 (N_13138,N_9718,N_9040);
and U13139 (N_13139,N_10437,N_11704);
or U13140 (N_13140,N_8254,N_11551);
and U13141 (N_13141,N_8616,N_8208);
nor U13142 (N_13142,N_9196,N_8207);
nor U13143 (N_13143,N_8707,N_11382);
or U13144 (N_13144,N_9958,N_10701);
or U13145 (N_13145,N_10103,N_9353);
nand U13146 (N_13146,N_9831,N_10026);
nand U13147 (N_13147,N_8161,N_11477);
nor U13148 (N_13148,N_8479,N_9311);
or U13149 (N_13149,N_9760,N_8221);
nor U13150 (N_13150,N_8543,N_11952);
nor U13151 (N_13151,N_9538,N_10081);
xor U13152 (N_13152,N_8083,N_9377);
or U13153 (N_13153,N_8992,N_9836);
nand U13154 (N_13154,N_11408,N_9675);
or U13155 (N_13155,N_8439,N_9643);
or U13156 (N_13156,N_11858,N_9704);
nand U13157 (N_13157,N_10646,N_11213);
nand U13158 (N_13158,N_10625,N_8581);
nand U13159 (N_13159,N_10059,N_10716);
and U13160 (N_13160,N_11464,N_10037);
or U13161 (N_13161,N_9531,N_11475);
nand U13162 (N_13162,N_10072,N_11670);
and U13163 (N_13163,N_8307,N_10151);
nand U13164 (N_13164,N_11144,N_11807);
nor U13165 (N_13165,N_8085,N_8137);
and U13166 (N_13166,N_10394,N_9867);
nor U13167 (N_13167,N_9135,N_8433);
and U13168 (N_13168,N_11847,N_11507);
nor U13169 (N_13169,N_9825,N_8045);
nand U13170 (N_13170,N_9905,N_9862);
nand U13171 (N_13171,N_10065,N_9061);
xnor U13172 (N_13172,N_11314,N_9618);
nor U13173 (N_13173,N_11480,N_10286);
nand U13174 (N_13174,N_9082,N_8561);
or U13175 (N_13175,N_8957,N_8212);
nand U13176 (N_13176,N_10620,N_11798);
nor U13177 (N_13177,N_8937,N_10739);
and U13178 (N_13178,N_9726,N_9237);
and U13179 (N_13179,N_11007,N_8320);
xnor U13180 (N_13180,N_11233,N_11630);
and U13181 (N_13181,N_10683,N_11175);
nand U13182 (N_13182,N_11708,N_10229);
and U13183 (N_13183,N_11606,N_9442);
nor U13184 (N_13184,N_11331,N_9255);
xor U13185 (N_13185,N_9179,N_9654);
nor U13186 (N_13186,N_9928,N_11684);
nand U13187 (N_13187,N_10368,N_9701);
nor U13188 (N_13188,N_9328,N_8507);
nor U13189 (N_13189,N_9167,N_9897);
nor U13190 (N_13190,N_9515,N_9246);
nand U13191 (N_13191,N_9799,N_10247);
nor U13192 (N_13192,N_9331,N_9615);
and U13193 (N_13193,N_9315,N_8475);
or U13194 (N_13194,N_9560,N_8634);
or U13195 (N_13195,N_9190,N_8588);
nand U13196 (N_13196,N_10805,N_9922);
nor U13197 (N_13197,N_11852,N_10710);
nand U13198 (N_13198,N_8227,N_10330);
or U13199 (N_13199,N_8784,N_10555);
nor U13200 (N_13200,N_9832,N_10970);
and U13201 (N_13201,N_9013,N_10363);
or U13202 (N_13202,N_10199,N_11555);
xnor U13203 (N_13203,N_9608,N_9535);
nor U13204 (N_13204,N_8216,N_8318);
or U13205 (N_13205,N_9795,N_10126);
nor U13206 (N_13206,N_10791,N_8802);
and U13207 (N_13207,N_9479,N_8367);
and U13208 (N_13208,N_11186,N_10402);
nor U13209 (N_13209,N_9676,N_11950);
and U13210 (N_13210,N_9236,N_9892);
or U13211 (N_13211,N_10704,N_10979);
and U13212 (N_13212,N_8117,N_11569);
or U13213 (N_13213,N_11196,N_9562);
nand U13214 (N_13214,N_10939,N_10189);
and U13215 (N_13215,N_11109,N_9763);
and U13216 (N_13216,N_10521,N_9906);
xor U13217 (N_13217,N_8610,N_11663);
nor U13218 (N_13218,N_10804,N_10450);
or U13219 (N_13219,N_8521,N_10424);
or U13220 (N_13220,N_8691,N_8073);
nor U13221 (N_13221,N_9895,N_9204);
and U13222 (N_13222,N_11235,N_10479);
or U13223 (N_13223,N_9006,N_11903);
nor U13224 (N_13224,N_8576,N_10274);
nor U13225 (N_13225,N_10562,N_11271);
or U13226 (N_13226,N_11405,N_10385);
or U13227 (N_13227,N_11091,N_8015);
and U13228 (N_13228,N_9871,N_11544);
xor U13229 (N_13229,N_9228,N_11673);
nor U13230 (N_13230,N_8872,N_10522);
nor U13231 (N_13231,N_10254,N_11195);
nor U13232 (N_13232,N_9176,N_10794);
or U13233 (N_13233,N_10263,N_8313);
nor U13234 (N_13234,N_10294,N_8943);
or U13235 (N_13235,N_9463,N_9486);
and U13236 (N_13236,N_11085,N_8070);
and U13237 (N_13237,N_8204,N_11039);
and U13238 (N_13238,N_10540,N_8821);
xnor U13239 (N_13239,N_8365,N_10594);
or U13240 (N_13240,N_8520,N_10462);
nor U13241 (N_13241,N_8000,N_8312);
and U13242 (N_13242,N_11042,N_10610);
xor U13243 (N_13243,N_11295,N_9732);
nand U13244 (N_13244,N_9432,N_9838);
xor U13245 (N_13245,N_8413,N_8584);
and U13246 (N_13246,N_11661,N_10219);
xnor U13247 (N_13247,N_11429,N_8690);
nand U13248 (N_13248,N_9754,N_9144);
or U13249 (N_13249,N_9074,N_8278);
xor U13250 (N_13250,N_10572,N_9137);
xor U13251 (N_13251,N_11997,N_8650);
or U13252 (N_13252,N_8124,N_9439);
or U13253 (N_13253,N_10032,N_9981);
or U13254 (N_13254,N_9471,N_10598);
and U13255 (N_13255,N_9318,N_11365);
and U13256 (N_13256,N_11959,N_9821);
or U13257 (N_13257,N_11834,N_10717);
or U13258 (N_13258,N_8062,N_11587);
and U13259 (N_13259,N_10524,N_11312);
nor U13260 (N_13260,N_11984,N_10908);
and U13261 (N_13261,N_10894,N_11566);
and U13262 (N_13262,N_9864,N_10962);
or U13263 (N_13263,N_10535,N_8999);
nor U13264 (N_13264,N_10357,N_11874);
and U13265 (N_13265,N_8244,N_8532);
nand U13266 (N_13266,N_8623,N_8564);
nor U13267 (N_13267,N_11063,N_11009);
and U13268 (N_13268,N_9780,N_11806);
or U13269 (N_13269,N_9352,N_10723);
nor U13270 (N_13270,N_8485,N_8153);
and U13271 (N_13271,N_8200,N_8363);
and U13272 (N_13272,N_10218,N_8309);
or U13273 (N_13273,N_8832,N_11898);
nand U13274 (N_13274,N_11266,N_10431);
and U13275 (N_13275,N_8663,N_10858);
nor U13276 (N_13276,N_8993,N_10642);
and U13277 (N_13277,N_10186,N_9184);
nor U13278 (N_13278,N_8571,N_9769);
nand U13279 (N_13279,N_11786,N_10583);
or U13280 (N_13280,N_8636,N_11236);
nor U13281 (N_13281,N_9420,N_8040);
or U13282 (N_13282,N_8454,N_9220);
or U13283 (N_13283,N_10576,N_11278);
nand U13284 (N_13284,N_11506,N_11987);
nand U13285 (N_13285,N_11498,N_10676);
nor U13286 (N_13286,N_8316,N_11187);
nor U13287 (N_13287,N_9422,N_9539);
nor U13288 (N_13288,N_11924,N_9188);
nand U13289 (N_13289,N_9447,N_10838);
nand U13290 (N_13290,N_11603,N_9384);
and U13291 (N_13291,N_10949,N_8104);
nor U13292 (N_13292,N_8798,N_10384);
and U13293 (N_13293,N_11426,N_8339);
and U13294 (N_13294,N_10225,N_8425);
nor U13295 (N_13295,N_11062,N_10896);
or U13296 (N_13296,N_9739,N_8232);
nand U13297 (N_13297,N_9058,N_8173);
or U13298 (N_13298,N_11001,N_11653);
nor U13299 (N_13299,N_10892,N_11676);
or U13300 (N_13300,N_10192,N_10388);
xor U13301 (N_13301,N_11398,N_9078);
nand U13302 (N_13302,N_9929,N_11268);
nor U13303 (N_13303,N_9345,N_8199);
and U13304 (N_13304,N_10780,N_10160);
nor U13305 (N_13305,N_10738,N_9908);
nand U13306 (N_13306,N_10570,N_8472);
nand U13307 (N_13307,N_8140,N_8057);
or U13308 (N_13308,N_10511,N_11542);
nor U13309 (N_13309,N_8929,N_11401);
nand U13310 (N_13310,N_9522,N_8271);
nand U13311 (N_13311,N_11757,N_10303);
or U13312 (N_13312,N_8429,N_10822);
nand U13313 (N_13313,N_9122,N_10109);
nand U13314 (N_13314,N_11539,N_11222);
nand U13315 (N_13315,N_10556,N_11901);
xnor U13316 (N_13316,N_9529,N_9741);
nand U13317 (N_13317,N_8358,N_9065);
or U13318 (N_13318,N_8948,N_9880);
xor U13319 (N_13319,N_9901,N_11543);
or U13320 (N_13320,N_8548,N_11671);
and U13321 (N_13321,N_10890,N_8255);
nand U13322 (N_13322,N_11486,N_11697);
or U13323 (N_13323,N_11485,N_9417);
and U13324 (N_13324,N_8218,N_9984);
and U13325 (N_13325,N_8648,N_10608);
nand U13326 (N_13326,N_8815,N_10993);
nor U13327 (N_13327,N_8026,N_10173);
xnor U13328 (N_13328,N_8072,N_8567);
or U13329 (N_13329,N_9628,N_8664);
nor U13330 (N_13330,N_9730,N_11380);
and U13331 (N_13331,N_8296,N_10269);
nor U13332 (N_13332,N_11734,N_11078);
and U13333 (N_13333,N_10952,N_9605);
and U13334 (N_13334,N_9678,N_8109);
and U13335 (N_13335,N_8008,N_9594);
xor U13336 (N_13336,N_10098,N_9723);
or U13337 (N_13337,N_11101,N_11249);
nand U13338 (N_13338,N_9493,N_10914);
nand U13339 (N_13339,N_11450,N_10414);
and U13340 (N_13340,N_8390,N_9325);
or U13341 (N_13341,N_11019,N_11765);
nor U13342 (N_13342,N_8956,N_8751);
and U13343 (N_13343,N_8491,N_10027);
nand U13344 (N_13344,N_9185,N_9707);
and U13345 (N_13345,N_10907,N_8130);
and U13346 (N_13346,N_8478,N_11226);
nand U13347 (N_13347,N_9932,N_11781);
nor U13348 (N_13348,N_11886,N_8776);
nand U13349 (N_13349,N_10730,N_10310);
and U13350 (N_13350,N_11769,N_11264);
and U13351 (N_13351,N_10754,N_11791);
nor U13352 (N_13352,N_11184,N_10068);
nor U13353 (N_13353,N_11154,N_9622);
and U13354 (N_13354,N_9514,N_11790);
xor U13355 (N_13355,N_9079,N_10073);
and U13356 (N_13356,N_11888,N_8220);
or U13357 (N_13357,N_10434,N_11801);
xor U13358 (N_13358,N_10016,N_11840);
or U13359 (N_13359,N_8329,N_8032);
nor U13360 (N_13360,N_10571,N_8515);
and U13361 (N_13361,N_10810,N_9747);
nor U13362 (N_13362,N_11639,N_8660);
nand U13363 (N_13363,N_8151,N_9894);
nor U13364 (N_13364,N_8853,N_9399);
xor U13365 (N_13365,N_11305,N_10835);
or U13366 (N_13366,N_11355,N_10505);
nand U13367 (N_13367,N_8826,N_8503);
and U13368 (N_13368,N_10242,N_9948);
nand U13369 (N_13369,N_10553,N_9028);
nor U13370 (N_13370,N_10317,N_10665);
xor U13371 (N_13371,N_10484,N_8694);
and U13372 (N_13372,N_11148,N_11370);
nor U13373 (N_13373,N_8188,N_9394);
or U13374 (N_13374,N_11345,N_8436);
nor U13375 (N_13375,N_8580,N_9693);
or U13376 (N_13376,N_8071,N_9194);
nand U13377 (N_13377,N_9518,N_8065);
xor U13378 (N_13378,N_9230,N_10851);
xor U13379 (N_13379,N_10865,N_8169);
and U13380 (N_13380,N_10000,N_10528);
nand U13381 (N_13381,N_9653,N_9993);
or U13382 (N_13382,N_11690,N_10919);
and U13383 (N_13383,N_10557,N_9733);
nor U13384 (N_13384,N_10868,N_9761);
nand U13385 (N_13385,N_9646,N_11302);
nor U13386 (N_13386,N_10878,N_9474);
or U13387 (N_13387,N_11687,N_9671);
or U13388 (N_13388,N_9327,N_9110);
or U13389 (N_13389,N_11504,N_8470);
nor U13390 (N_13390,N_11629,N_10885);
and U13391 (N_13391,N_8979,N_11916);
nand U13392 (N_13392,N_9339,N_10124);
nand U13393 (N_13393,N_8594,N_11463);
or U13394 (N_13394,N_10129,N_11335);
xor U13395 (N_13395,N_11239,N_10125);
nand U13396 (N_13396,N_9972,N_8560);
nand U13397 (N_13397,N_10420,N_10166);
nand U13398 (N_13398,N_9530,N_11460);
nor U13399 (N_13399,N_10847,N_8923);
or U13400 (N_13400,N_11932,N_11547);
nand U13401 (N_13401,N_10114,N_10863);
or U13402 (N_13402,N_10820,N_10960);
nand U13403 (N_13403,N_11156,N_9851);
nor U13404 (N_13404,N_8506,N_10900);
and U13405 (N_13405,N_9195,N_9655);
and U13406 (N_13406,N_10238,N_10655);
and U13407 (N_13407,N_8601,N_8761);
and U13408 (N_13408,N_8765,N_10113);
nand U13409 (N_13409,N_8295,N_9348);
nor U13410 (N_13410,N_10998,N_10624);
or U13411 (N_13411,N_11351,N_11204);
nand U13412 (N_13412,N_10966,N_9846);
or U13413 (N_13413,N_9898,N_8778);
nor U13414 (N_13414,N_9289,N_8125);
and U13415 (N_13415,N_9087,N_9983);
or U13416 (N_13416,N_10604,N_11669);
or U13417 (N_13417,N_9186,N_10288);
nand U13418 (N_13418,N_11321,N_10339);
xor U13419 (N_13419,N_9429,N_9910);
or U13420 (N_13420,N_11349,N_8327);
nor U13421 (N_13421,N_10245,N_8733);
nor U13422 (N_13422,N_8884,N_10831);
nand U13423 (N_13423,N_10817,N_10285);
nand U13424 (N_13424,N_8944,N_10093);
nor U13425 (N_13425,N_10184,N_9946);
and U13426 (N_13426,N_8116,N_11378);
nor U13427 (N_13427,N_8354,N_8095);
and U13428 (N_13428,N_11415,N_11449);
and U13429 (N_13429,N_10601,N_11802);
or U13430 (N_13430,N_9095,N_10844);
nand U13431 (N_13431,N_10048,N_8674);
nand U13432 (N_13432,N_9162,N_9801);
nand U13433 (N_13433,N_10230,N_10787);
and U13434 (N_13434,N_11330,N_10518);
or U13435 (N_13435,N_10997,N_9492);
nor U13436 (N_13436,N_8812,N_11792);
or U13437 (N_13437,N_8251,N_9092);
nand U13438 (N_13438,N_10539,N_11430);
or U13439 (N_13439,N_8759,N_8420);
and U13440 (N_13440,N_10566,N_8715);
and U13441 (N_13441,N_11647,N_11884);
xor U13442 (N_13442,N_10940,N_9427);
or U13443 (N_13443,N_11577,N_9030);
and U13444 (N_13444,N_8736,N_11748);
and U13445 (N_13445,N_11702,N_8910);
nand U13446 (N_13446,N_9407,N_9292);
or U13447 (N_13447,N_9406,N_11777);
nand U13448 (N_13448,N_10913,N_11556);
and U13449 (N_13449,N_11387,N_8524);
and U13450 (N_13450,N_11125,N_10564);
and U13451 (N_13451,N_11447,N_11683);
and U13452 (N_13452,N_11922,N_10190);
or U13453 (N_13453,N_11353,N_10216);
nor U13454 (N_13454,N_11995,N_9310);
or U13455 (N_13455,N_9036,N_10877);
and U13456 (N_13456,N_11666,N_11863);
nor U13457 (N_13457,N_11301,N_11795);
nand U13458 (N_13458,N_11515,N_10372);
or U13459 (N_13459,N_10049,N_8056);
or U13460 (N_13460,N_11169,N_10841);
nand U13461 (N_13461,N_9857,N_10702);
and U13462 (N_13462,N_9758,N_10740);
and U13463 (N_13463,N_8669,N_11568);
or U13464 (N_13464,N_9947,N_10280);
nand U13465 (N_13465,N_9988,N_8814);
nand U13466 (N_13466,N_9055,N_11797);
nand U13467 (N_13467,N_9296,N_11519);
nor U13468 (N_13468,N_9070,N_11565);
or U13469 (N_13469,N_11210,N_8713);
nor U13470 (N_13470,N_9437,N_11183);
nor U13471 (N_13471,N_8409,N_11810);
or U13472 (N_13472,N_9703,N_9193);
nand U13473 (N_13473,N_8739,N_11069);
nand U13474 (N_13474,N_9869,N_8074);
nor U13475 (N_13475,N_10214,N_10963);
nor U13476 (N_13476,N_9918,N_9629);
and U13477 (N_13477,N_10667,N_11664);
and U13478 (N_13478,N_11473,N_8735);
nor U13479 (N_13479,N_11988,N_10422);
and U13480 (N_13480,N_10119,N_9875);
nor U13481 (N_13481,N_8372,N_10996);
or U13482 (N_13482,N_11823,N_9039);
or U13483 (N_13483,N_10492,N_11841);
or U13484 (N_13484,N_11158,N_9582);
nand U13485 (N_13485,N_11662,N_10175);
and U13486 (N_13486,N_10064,N_9288);
or U13487 (N_13487,N_11846,N_9885);
nor U13488 (N_13488,N_9349,N_10464);
nor U13489 (N_13489,N_9589,N_9696);
and U13490 (N_13490,N_11481,N_11650);
or U13491 (N_13491,N_10500,N_11298);
or U13492 (N_13492,N_10793,N_8027);
nand U13493 (N_13493,N_11672,N_11981);
xnor U13494 (N_13494,N_11211,N_11711);
nor U13495 (N_13495,N_11227,N_11400);
or U13496 (N_13496,N_10256,N_10951);
and U13497 (N_13497,N_11965,N_11457);
and U13498 (N_13498,N_11178,N_8196);
and U13499 (N_13499,N_8293,N_8267);
nand U13500 (N_13500,N_10476,N_9796);
or U13501 (N_13501,N_11604,N_9735);
nor U13502 (N_13502,N_10618,N_10769);
nand U13503 (N_13503,N_8709,N_8544);
and U13504 (N_13504,N_8785,N_11747);
or U13505 (N_13505,N_8539,N_10513);
nand U13506 (N_13506,N_11532,N_10613);
nor U13507 (N_13507,N_11263,N_10596);
and U13508 (N_13508,N_11928,N_9297);
and U13509 (N_13509,N_8945,N_11087);
or U13510 (N_13510,N_11021,N_10489);
nor U13511 (N_13511,N_9999,N_9830);
or U13512 (N_13512,N_10876,N_11344);
and U13513 (N_13513,N_11193,N_11600);
nor U13514 (N_13514,N_9668,N_11754);
nand U13515 (N_13515,N_8113,N_8692);
and U13516 (N_13516,N_11217,N_8760);
and U13517 (N_13517,N_10421,N_11171);
and U13518 (N_13518,N_10554,N_10883);
nand U13519 (N_13519,N_9505,N_11325);
or U13520 (N_13520,N_10182,N_10337);
and U13521 (N_13521,N_8773,N_11100);
or U13522 (N_13522,N_8055,N_10416);
xnor U13523 (N_13523,N_9201,N_11618);
and U13524 (N_13524,N_8917,N_8727);
or U13525 (N_13525,N_11341,N_9561);
or U13526 (N_13526,N_9392,N_10652);
nor U13527 (N_13527,N_10042,N_8488);
and U13528 (N_13528,N_10733,N_10656);
nor U13529 (N_13529,N_11913,N_11522);
nor U13530 (N_13530,N_10815,N_8223);
xor U13531 (N_13531,N_11991,N_11529);
xor U13532 (N_13532,N_9827,N_10089);
and U13533 (N_13533,N_8807,N_10369);
or U13534 (N_13534,N_10653,N_9635);
or U13535 (N_13535,N_8538,N_11117);
nand U13536 (N_13536,N_9512,N_11297);
nor U13537 (N_13537,N_8631,N_11851);
and U13538 (N_13538,N_8468,N_9354);
nor U13539 (N_13539,N_11079,N_8236);
and U13540 (N_13540,N_10428,N_10009);
and U13541 (N_13541,N_8202,N_11944);
nor U13542 (N_13542,N_10619,N_8423);
nand U13543 (N_13543,N_11010,N_8089);
or U13544 (N_13544,N_8645,N_9462);
nand U13545 (N_13545,N_8900,N_9805);
nand U13546 (N_13546,N_10912,N_11613);
nand U13547 (N_13547,N_9117,N_9225);
nand U13548 (N_13548,N_11041,N_9670);
xor U13549 (N_13549,N_10623,N_8249);
nor U13550 (N_13550,N_8732,N_8803);
and U13551 (N_13551,N_10578,N_8416);
and U13552 (N_13552,N_11046,N_11943);
or U13553 (N_13553,N_11428,N_10776);
or U13554 (N_13554,N_11364,N_9559);
nor U13555 (N_13555,N_8617,N_8946);
and U13556 (N_13556,N_9319,N_9820);
and U13557 (N_13557,N_10313,N_10267);
nor U13558 (N_13558,N_8578,N_9257);
nand U13559 (N_13559,N_10509,N_10127);
nor U13560 (N_13560,N_11099,N_8237);
nand U13561 (N_13561,N_9284,N_9445);
nor U13562 (N_13562,N_10823,N_8768);
and U13563 (N_13563,N_11176,N_8518);
nand U13564 (N_13564,N_9638,N_11339);
xor U13565 (N_13565,N_11845,N_11994);
nand U13566 (N_13566,N_9565,N_8252);
or U13567 (N_13567,N_11181,N_8901);
or U13568 (N_13568,N_10643,N_9387);
and U13569 (N_13569,N_9355,N_11935);
nand U13570 (N_13570,N_10980,N_9664);
nor U13571 (N_13571,N_11537,N_10674);
and U13572 (N_13572,N_8222,N_10680);
or U13573 (N_13573,N_11779,N_11700);
or U13574 (N_13574,N_9587,N_11319);
and U13575 (N_13575,N_10829,N_11920);
or U13576 (N_13576,N_10465,N_9366);
nor U13577 (N_13577,N_8600,N_8110);
nor U13578 (N_13578,N_10371,N_10282);
nor U13579 (N_13579,N_9234,N_9241);
or U13580 (N_13580,N_8185,N_8550);
or U13581 (N_13581,N_8122,N_8118);
and U13582 (N_13582,N_8175,N_9251);
or U13583 (N_13583,N_10813,N_8553);
xnor U13584 (N_13584,N_9370,N_11096);
and U13585 (N_13585,N_8230,N_9371);
or U13586 (N_13586,N_8514,N_8131);
nor U13587 (N_13587,N_8996,N_9812);
nand U13588 (N_13588,N_9783,N_8419);
nand U13589 (N_13589,N_8780,N_8907);
or U13590 (N_13590,N_11973,N_9689);
or U13591 (N_13591,N_10475,N_8194);
nor U13592 (N_13592,N_10533,N_10591);
nor U13593 (N_13593,N_8895,N_10020);
xor U13594 (N_13594,N_11958,N_11289);
nor U13595 (N_13595,N_11941,N_9483);
and U13596 (N_13596,N_9256,N_9978);
nor U13597 (N_13597,N_9052,N_9965);
and U13598 (N_13598,N_10573,N_8903);
nor U13599 (N_13599,N_9173,N_11002);
or U13600 (N_13600,N_10743,N_8213);
nor U13601 (N_13601,N_11953,N_10837);
or U13602 (N_13602,N_9472,N_9060);
and U13603 (N_13603,N_8004,N_8274);
xnor U13604 (N_13604,N_11040,N_9452);
or U13605 (N_13605,N_8349,N_10343);
and U13606 (N_13606,N_11805,N_8287);
nor U13607 (N_13607,N_9397,N_11762);
nor U13608 (N_13608,N_8828,N_11744);
nor U13609 (N_13609,N_8029,N_10579);
nand U13610 (N_13610,N_11250,N_10345);
nor U13611 (N_13611,N_8209,N_9294);
nand U13612 (N_13612,N_10010,N_8746);
nor U13613 (N_13613,N_11915,N_8455);
and U13614 (N_13614,N_10986,N_9295);
nor U13615 (N_13615,N_10121,N_9536);
or U13616 (N_13616,N_10531,N_9633);
nand U13617 (N_13617,N_10905,N_10396);
or U13618 (N_13618,N_9944,N_11579);
or U13619 (N_13619,N_11575,N_10703);
nor U13620 (N_13620,N_9242,N_8976);
nand U13621 (N_13621,N_9853,N_10319);
and U13622 (N_13622,N_10719,N_10084);
nor U13623 (N_13623,N_9454,N_8960);
nor U13624 (N_13624,N_11326,N_8147);
xnor U13625 (N_13625,N_8698,N_8925);
nor U13626 (N_13626,N_9716,N_8284);
nor U13627 (N_13627,N_8257,N_11536);
nand U13628 (N_13628,N_8013,N_10757);
xnor U13629 (N_13629,N_8554,N_11373);
nand U13630 (N_13630,N_10694,N_9882);
or U13631 (N_13631,N_10083,N_9516);
nor U13632 (N_13632,N_8205,N_11789);
and U13633 (N_13633,N_8841,N_10200);
nor U13634 (N_13634,N_11622,N_8591);
and U13635 (N_13635,N_9602,N_9647);
nor U13636 (N_13636,N_9101,N_9104);
nor U13637 (N_13637,N_11369,N_11407);
or U13638 (N_13638,N_8171,N_8546);
or U13639 (N_13639,N_11516,N_10380);
nand U13640 (N_13640,N_9160,N_8864);
and U13641 (N_13641,N_10086,N_11937);
xor U13642 (N_13642,N_8941,N_8258);
and U13643 (N_13643,N_9544,N_9171);
and U13644 (N_13644,N_11413,N_8302);
and U13645 (N_13645,N_8932,N_8211);
or U13646 (N_13646,N_9044,N_9510);
and U13647 (N_13647,N_10159,N_11503);
and U13648 (N_13648,N_11591,N_11534);
nor U13649 (N_13649,N_11509,N_11374);
or U13650 (N_13650,N_10115,N_10862);
nor U13651 (N_13651,N_9573,N_9218);
xnor U13652 (N_13652,N_10191,N_10222);
or U13653 (N_13653,N_11818,N_9187);
nor U13654 (N_13654,N_11518,N_10560);
nand U13655 (N_13655,N_10809,N_10373);
or U13656 (N_13656,N_8705,N_11722);
or U13657 (N_13657,N_9709,N_11720);
nor U13658 (N_13658,N_8036,N_11619);
nand U13659 (N_13659,N_8128,N_8010);
nand U13660 (N_13660,N_11276,N_10755);
nor U13661 (N_13661,N_9849,N_10427);
nor U13662 (N_13662,N_10144,N_10051);
or U13663 (N_13663,N_8856,N_8818);
and U13664 (N_13664,N_9742,N_9634);
nor U13665 (N_13665,N_10092,N_8619);
or U13666 (N_13666,N_9350,N_10515);
xnor U13667 (N_13667,N_8953,N_9848);
or U13668 (N_13668,N_9509,N_8717);
nand U13669 (N_13669,N_8958,N_11161);
or U13670 (N_13670,N_10017,N_8987);
xor U13671 (N_13671,N_11573,N_9229);
nor U13672 (N_13672,N_9125,N_8885);
nor U13673 (N_13673,N_10990,N_11359);
nor U13674 (N_13674,N_9478,N_11889);
nor U13675 (N_13675,N_8303,N_9012);
and U13676 (N_13676,N_8003,N_8542);
nand U13677 (N_13677,N_9658,N_9494);
nor U13678 (N_13678,N_11954,N_8201);
nand U13679 (N_13679,N_11743,N_9200);
or U13680 (N_13680,N_11570,N_9779);
nor U13681 (N_13681,N_9992,N_11768);
nand U13682 (N_13682,N_10399,N_11955);
and U13683 (N_13683,N_8041,N_11585);
nor U13684 (N_13684,N_9614,N_10013);
nor U13685 (N_13685,N_9097,N_11340);
xor U13686 (N_13686,N_10543,N_9480);
and U13687 (N_13687,N_9347,N_10055);
and U13688 (N_13688,N_11034,N_8422);
and U13689 (N_13689,N_9088,N_9964);
nand U13690 (N_13690,N_10446,N_11656);
or U13691 (N_13691,N_11892,N_8575);
nor U13692 (N_13692,N_9955,N_10359);
or U13693 (N_13693,N_8005,N_8970);
and U13694 (N_13694,N_11897,N_9859);
nor U13695 (N_13695,N_11689,N_9728);
xnor U13696 (N_13696,N_11277,N_11859);
nor U13697 (N_13697,N_8846,N_10451);
nand U13698 (N_13698,N_8769,N_10025);
and U13699 (N_13699,N_10926,N_10731);
or U13700 (N_13700,N_11977,N_11766);
or U13701 (N_13701,N_11024,N_9382);
or U13702 (N_13702,N_8593,N_11857);
or U13703 (N_13703,N_8702,N_11128);
and U13704 (N_13704,N_11710,N_10291);
or U13705 (N_13705,N_8605,N_9138);
or U13706 (N_13706,N_8896,N_11999);
or U13707 (N_13707,N_10426,N_9064);
or U13708 (N_13708,N_9874,N_10749);
and U13709 (N_13709,N_11350,N_9333);
and U13710 (N_13710,N_11416,N_8902);
or U13711 (N_13711,N_10976,N_9224);
nor U13712 (N_13712,N_8906,N_9873);
or U13713 (N_13713,N_10639,N_11535);
and U13714 (N_13714,N_8714,N_11052);
nor U13715 (N_13715,N_11327,N_9238);
nand U13716 (N_13716,N_10257,N_8772);
and U13717 (N_13717,N_8806,N_9287);
xnor U13718 (N_13718,N_9372,N_8741);
and U13719 (N_13719,N_10924,N_9797);
nor U13720 (N_13720,N_11599,N_9169);
nand U13721 (N_13721,N_9599,N_11721);
and U13722 (N_13722,N_11538,N_9917);
nand U13723 (N_13723,N_8875,N_11225);
or U13724 (N_13724,N_10123,N_9543);
or U13725 (N_13725,N_9080,N_8916);
or U13726 (N_13726,N_11379,N_11160);
or U13727 (N_13727,N_8136,N_8081);
nor U13728 (N_13728,N_10724,N_9081);
or U13729 (N_13729,N_10366,N_9680);
or U13730 (N_13730,N_8629,N_8451);
and U13731 (N_13731,N_11036,N_8936);
and U13732 (N_13732,N_10961,N_10950);
nor U13733 (N_13733,N_11273,N_11015);
nand U13734 (N_13734,N_10602,N_8680);
nor U13735 (N_13735,N_9223,N_9244);
and U13736 (N_13736,N_10362,N_9569);
nor U13737 (N_13737,N_10149,N_9751);
nand U13738 (N_13738,N_8094,N_11811);
nand U13739 (N_13739,N_8595,N_9621);
and U13740 (N_13740,N_11216,N_8038);
xnor U13741 (N_13741,N_9170,N_8058);
nor U13742 (N_13742,N_8328,N_11433);
nand U13743 (N_13743,N_9213,N_8179);
xnor U13744 (N_13744,N_10720,N_9912);
or U13745 (N_13745,N_8412,N_10935);
or U13746 (N_13746,N_10577,N_10581);
nor U13747 (N_13747,N_8685,N_9772);
nand U13748 (N_13748,N_11550,N_8927);
or U13749 (N_13749,N_9500,N_8346);
and U13750 (N_13750,N_10210,N_10172);
or U13751 (N_13751,N_11442,N_9291);
and U13752 (N_13752,N_10071,N_11238);
and U13753 (N_13753,N_8102,N_10612);
nand U13754 (N_13754,N_8087,N_10302);
nor U13755 (N_13755,N_9275,N_10334);
and U13756 (N_13756,N_9245,N_10033);
and U13757 (N_13757,N_10736,N_8054);
and U13758 (N_13758,N_11107,N_11908);
nor U13759 (N_13759,N_9145,N_11793);
and U13760 (N_13760,N_10297,N_11736);
nor U13761 (N_13761,N_11140,N_11287);
nor U13762 (N_13762,N_9481,N_10503);
and U13763 (N_13763,N_9659,N_9591);
xor U13764 (N_13764,N_9298,N_10567);
and U13765 (N_13765,N_10460,N_11011);
or U13766 (N_13766,N_9180,N_8653);
and U13767 (N_13767,N_11016,N_11348);
nand U13768 (N_13768,N_8858,N_9660);
or U13769 (N_13769,N_8755,N_11586);
nand U13770 (N_13770,N_8270,N_9129);
and U13771 (N_13771,N_9140,N_10832);
xor U13772 (N_13772,N_10587,N_10265);
nor U13773 (N_13773,N_8215,N_9215);
and U13774 (N_13774,N_10948,N_9023);
or U13775 (N_13775,N_10995,N_8426);
and U13776 (N_13776,N_10644,N_11206);
nand U13777 (N_13777,N_11020,N_9115);
or U13778 (N_13778,N_9277,N_9860);
and U13779 (N_13779,N_9884,N_10099);
nand U13780 (N_13780,N_9019,N_11531);
and U13781 (N_13781,N_8693,N_10220);
and U13782 (N_13782,N_8486,N_8487);
and U13783 (N_13783,N_11610,N_11611);
or U13784 (N_13784,N_9600,N_8966);
or U13785 (N_13785,N_9332,N_8990);
or U13786 (N_13786,N_11729,N_9496);
nand U13787 (N_13787,N_11594,N_9098);
nor U13788 (N_13788,N_11927,N_11530);
nor U13789 (N_13789,N_10311,N_10376);
and U13790 (N_13790,N_11620,N_10760);
nand U13791 (N_13791,N_8164,N_11753);
nor U13792 (N_13792,N_8589,N_8643);
nand U13793 (N_13793,N_9883,N_8019);
nor U13794 (N_13794,N_8822,N_10057);
and U13795 (N_13795,N_8627,N_10471);
nor U13796 (N_13796,N_8133,N_8750);
nor U13797 (N_13797,N_9436,N_8396);
and U13798 (N_13798,N_8229,N_8838);
nand U13799 (N_13799,N_9421,N_11848);
or U13800 (N_13800,N_9316,N_9507);
and U13801 (N_13801,N_10689,N_11598);
and U13802 (N_13802,N_9881,N_11461);
and U13803 (N_13803,N_8299,N_10550);
xor U13804 (N_13804,N_10606,N_9363);
nor U13805 (N_13805,N_11963,N_8262);
nor U13806 (N_13806,N_10833,N_8889);
nand U13807 (N_13807,N_8145,N_11827);
nor U13808 (N_13808,N_8792,N_9376);
or U13809 (N_13809,N_10605,N_9379);
xnor U13810 (N_13810,N_9499,N_9904);
xor U13811 (N_13811,N_9434,N_9131);
nor U13812 (N_13812,N_9113,N_9425);
nand U13813 (N_13813,N_8495,N_11947);
nand U13814 (N_13814,N_10091,N_9828);
and U13815 (N_13815,N_10074,N_10889);
and U13816 (N_13816,N_9803,N_9580);
or U13817 (N_13817,N_9570,N_9699);
nor U13818 (N_13818,N_11581,N_10398);
and U13819 (N_13819,N_8242,N_8193);
nor U13820 (N_13820,N_8428,N_10773);
nand U13821 (N_13821,N_10488,N_9441);
and U13822 (N_13822,N_10387,N_11467);
nand U13823 (N_13823,N_11883,N_10746);
and U13824 (N_13824,N_9624,N_9532);
xnor U13825 (N_13825,N_8375,N_10568);
nand U13826 (N_13826,N_10967,N_8380);
or U13827 (N_13827,N_11993,N_8272);
and U13828 (N_13828,N_10389,N_10790);
nand U13829 (N_13829,N_11636,N_8675);
nand U13830 (N_13830,N_9640,N_10628);
xnor U13831 (N_13831,N_8712,N_8378);
or U13832 (N_13832,N_9776,N_9508);
nand U13833 (N_13833,N_9804,N_9767);
and U13834 (N_13834,N_11696,N_8794);
nand U13835 (N_13835,N_11749,N_8441);
xor U13836 (N_13836,N_8264,N_9412);
xor U13837 (N_13837,N_9837,N_8796);
and U13838 (N_13838,N_11393,N_8195);
nor U13839 (N_13839,N_8748,N_10116);
xor U13840 (N_13840,N_10969,N_9423);
and U13841 (N_13841,N_9945,N_8579);
nand U13842 (N_13842,N_8014,N_9252);
and U13843 (N_13843,N_11849,N_9650);
nor U13844 (N_13844,N_9136,N_10514);
nand U13845 (N_13845,N_8686,N_9719);
nand U13846 (N_13846,N_11605,N_9750);
nand U13847 (N_13847,N_9404,N_10945);
or U13848 (N_13848,N_8067,N_8651);
and U13849 (N_13849,N_9114,N_8387);
or U13850 (N_13850,N_9305,N_9326);
and U13851 (N_13851,N_9641,N_9979);
xor U13852 (N_13852,N_8245,N_8536);
and U13853 (N_13853,N_11637,N_8753);
and U13854 (N_13854,N_8977,N_9649);
nand U13855 (N_13855,N_9617,N_8405);
or U13856 (N_13856,N_10697,N_9330);
nor U13857 (N_13857,N_8512,N_10575);
nor U13858 (N_13858,N_8228,N_9651);
and U13859 (N_13859,N_10223,N_11815);
xor U13860 (N_13860,N_11232,N_11654);
or U13861 (N_13861,N_9216,N_9604);
and U13862 (N_13862,N_11482,N_8825);
and U13863 (N_13863,N_11723,N_8829);
or U13864 (N_13864,N_11157,N_11258);
nor U13865 (N_13865,N_8304,N_11307);
and U13866 (N_13866,N_11496,N_11912);
xnor U13867 (N_13867,N_11316,N_10735);
and U13868 (N_13868,N_11188,N_11497);
xor U13869 (N_13869,N_11564,N_9502);
nor U13870 (N_13870,N_11742,N_8351);
or U13871 (N_13871,N_11399,N_9878);
nor U13872 (N_13872,N_8191,N_8967);
and U13873 (N_13873,N_8565,N_10087);
nand U13874 (N_13874,N_11038,N_11745);
nand U13875 (N_13875,N_11490,N_8447);
and U13876 (N_13876,N_10490,N_10988);
or U13877 (N_13877,N_11386,N_9253);
xnor U13878 (N_13878,N_9691,N_8926);
and U13879 (N_13879,N_9682,N_10276);
or U13880 (N_13880,N_10799,N_10818);
nor U13881 (N_13881,N_11679,N_10445);
nand U13882 (N_13882,N_9991,N_8469);
nand U13883 (N_13883,N_8614,N_11267);
or U13884 (N_13884,N_10227,N_11860);
nor U13885 (N_13885,N_11418,N_10353);
nand U13886 (N_13886,N_11166,N_8011);
and U13887 (N_13887,N_11150,N_11583);
or U13888 (N_13888,N_8398,N_11730);
or U13889 (N_13889,N_11911,N_10226);
or U13890 (N_13890,N_8361,N_9907);
nor U13891 (N_13891,N_11856,N_10681);
and U13892 (N_13892,N_9357,N_8894);
or U13893 (N_13893,N_9024,N_10692);
nor U13894 (N_13894,N_10472,N_9705);
and U13895 (N_13895,N_10872,N_8656);
or U13896 (N_13896,N_11363,N_11055);
nand U13897 (N_13897,N_8489,N_9046);
and U13898 (N_13898,N_11740,N_11832);
or U13899 (N_13899,N_11990,N_10615);
and U13900 (N_13900,N_8638,N_8028);
or U13901 (N_13901,N_8415,N_8942);
nand U13902 (N_13902,N_10671,N_10075);
nand U13903 (N_13903,N_9396,N_8156);
and U13904 (N_13904,N_10814,N_11409);
nand U13905 (N_13905,N_9645,N_9211);
xor U13906 (N_13906,N_11444,N_10958);
nor U13907 (N_13907,N_11468,N_8180);
and U13908 (N_13908,N_9920,N_9102);
nor U13909 (N_13909,N_11597,N_11246);
or U13910 (N_13910,N_8373,N_9207);
nor U13911 (N_13911,N_8499,N_11682);
and U13912 (N_13912,N_8920,N_8226);
nand U13913 (N_13913,N_8540,N_10361);
and U13914 (N_13914,N_10155,N_10447);
nand U13915 (N_13915,N_8756,N_9469);
nor U13916 (N_13916,N_10507,N_11324);
nand U13917 (N_13917,N_11872,N_11552);
or U13918 (N_13918,N_9877,N_11333);
xnor U13919 (N_13919,N_10401,N_9987);
xnor U13920 (N_13920,N_11593,N_8017);
nor U13921 (N_13921,N_8585,N_10351);
or U13922 (N_13922,N_8421,N_10410);
nor U13923 (N_13923,N_8465,N_11200);
and U13924 (N_13924,N_9043,N_8484);
nand U13925 (N_13925,N_10448,N_8326);
and U13926 (N_13926,N_9484,N_9810);
xnor U13927 (N_13927,N_11432,N_9057);
nor U13928 (N_13928,N_10679,N_10196);
and U13929 (N_13929,N_8774,N_11142);
xor U13930 (N_13930,N_10636,N_10154);
nor U13931 (N_13931,N_8059,N_10249);
or U13932 (N_13932,N_8460,N_9970);
nand U13933 (N_13933,N_9663,N_10466);
nand U13934 (N_13934,N_11681,N_9274);
and U13935 (N_13935,N_10241,N_11992);
and U13936 (N_13936,N_8555,N_8980);
or U13937 (N_13937,N_9004,N_9444);
nand U13938 (N_13938,N_9034,N_10537);
nor U13939 (N_13939,N_10058,N_9281);
or U13940 (N_13940,N_8364,N_8559);
nor U13941 (N_13941,N_11385,N_8682);
nand U13942 (N_13942,N_8308,N_10726);
and U13943 (N_13943,N_10300,N_8359);
xnor U13944 (N_13944,N_11976,N_11951);
and U13945 (N_13945,N_9466,N_9731);
nand U13946 (N_13946,N_8574,N_9464);
or U13947 (N_13947,N_10873,N_8678);
nor U13948 (N_13948,N_9845,N_11741);
and U13949 (N_13949,N_9564,N_8183);
and U13950 (N_13950,N_8090,N_8192);
and U13951 (N_13951,N_10044,N_10795);
and U13952 (N_13952,N_11649,N_9520);
and U13953 (N_13953,N_11601,N_11094);
nand U13954 (N_13954,N_8533,N_8615);
nor U13955 (N_13955,N_9071,N_8031);
nand U13956 (N_13956,N_9390,N_10888);
nand U13957 (N_13957,N_8915,N_11329);
nor U13958 (N_13958,N_11495,N_8758);
xor U13959 (N_13959,N_9069,N_10157);
nor U13960 (N_13960,N_10270,N_11280);
and U13961 (N_13961,N_8111,N_9282);
and U13962 (N_13962,N_10486,N_11424);
nor U13963 (N_13963,N_8319,N_11451);
nor U13964 (N_13964,N_10001,N_8162);
and U13965 (N_13965,N_8384,N_8144);
nor U13966 (N_13966,N_9925,N_8767);
nand U13967 (N_13967,N_11523,N_11646);
and U13968 (N_13968,N_10712,N_8848);
nand U13969 (N_13969,N_11980,N_11354);
nor U13970 (N_13970,N_8658,N_11978);
and U13971 (N_13971,N_10281,N_9792);
or U13972 (N_13972,N_11116,N_10861);
or U13973 (N_13973,N_10867,N_11453);
xnor U13974 (N_13974,N_8963,N_11440);
and U13975 (N_13975,N_11209,N_11751);
or U13976 (N_13976,N_9128,N_11491);
and U13977 (N_13977,N_9826,N_10761);
or U13978 (N_13978,N_9010,N_8582);
nor U13979 (N_13979,N_8728,N_11918);
nor U13980 (N_13980,N_8968,N_9975);
and U13981 (N_13981,N_8940,N_8097);
xor U13982 (N_13982,N_8708,N_10826);
nor U13983 (N_13983,N_8330,N_9278);
and U13984 (N_13984,N_8819,N_11862);
nand U13985 (N_13985,N_11252,N_9702);
and U13986 (N_13986,N_10036,N_8002);
nor U13987 (N_13987,N_11707,N_9919);
and U13988 (N_13988,N_11835,N_8793);
nor U13989 (N_13989,N_11030,N_8701);
or U13990 (N_13990,N_11596,N_8350);
and U13991 (N_13991,N_9579,N_8021);
nand U13992 (N_13992,N_8607,N_8277);
nor U13993 (N_13993,N_11694,N_10959);
nor U13994 (N_13994,N_10408,N_9066);
and U13995 (N_13995,N_10107,N_10582);
nand U13996 (N_13996,N_8641,N_11061);
and U13997 (N_13997,N_8437,N_9766);
nand U13998 (N_13998,N_11279,N_8360);
and U13999 (N_13999,N_9724,N_9438);
nand U14000 (N_14000,N_10628,N_11843);
nor U14001 (N_14001,N_9941,N_11298);
and U14002 (N_14002,N_8867,N_9073);
nor U14003 (N_14003,N_9452,N_8863);
nor U14004 (N_14004,N_8061,N_10044);
xor U14005 (N_14005,N_8327,N_11599);
xnor U14006 (N_14006,N_11054,N_8240);
and U14007 (N_14007,N_9762,N_11717);
xnor U14008 (N_14008,N_11975,N_10852);
and U14009 (N_14009,N_9920,N_10558);
and U14010 (N_14010,N_9095,N_9819);
or U14011 (N_14011,N_8462,N_9477);
and U14012 (N_14012,N_10653,N_9058);
nor U14013 (N_14013,N_10018,N_11696);
or U14014 (N_14014,N_9305,N_10696);
xnor U14015 (N_14015,N_8290,N_9481);
or U14016 (N_14016,N_10778,N_11315);
nor U14017 (N_14017,N_11993,N_9816);
nor U14018 (N_14018,N_8120,N_9350);
nand U14019 (N_14019,N_11924,N_9851);
or U14020 (N_14020,N_9136,N_9983);
and U14021 (N_14021,N_8908,N_8498);
nand U14022 (N_14022,N_8049,N_10550);
nand U14023 (N_14023,N_11167,N_10036);
nand U14024 (N_14024,N_8963,N_9124);
or U14025 (N_14025,N_11620,N_10678);
nand U14026 (N_14026,N_11934,N_9834);
and U14027 (N_14027,N_10616,N_8531);
xnor U14028 (N_14028,N_10927,N_10624);
nor U14029 (N_14029,N_9689,N_8220);
nor U14030 (N_14030,N_9697,N_11313);
or U14031 (N_14031,N_8889,N_8826);
or U14032 (N_14032,N_8301,N_11149);
and U14033 (N_14033,N_11942,N_10561);
nand U14034 (N_14034,N_9821,N_9036);
nand U14035 (N_14035,N_11015,N_11602);
or U14036 (N_14036,N_8174,N_8813);
or U14037 (N_14037,N_9815,N_8299);
and U14038 (N_14038,N_10549,N_11242);
nor U14039 (N_14039,N_8663,N_8096);
and U14040 (N_14040,N_8462,N_11389);
and U14041 (N_14041,N_10429,N_8487);
nor U14042 (N_14042,N_8254,N_8123);
nand U14043 (N_14043,N_10059,N_11155);
nand U14044 (N_14044,N_11775,N_11723);
and U14045 (N_14045,N_11518,N_9254);
xor U14046 (N_14046,N_8020,N_9720);
nor U14047 (N_14047,N_10367,N_11553);
or U14048 (N_14048,N_10515,N_11594);
nor U14049 (N_14049,N_10842,N_9952);
nand U14050 (N_14050,N_8855,N_11044);
or U14051 (N_14051,N_8167,N_9085);
nand U14052 (N_14052,N_9382,N_9161);
and U14053 (N_14053,N_11929,N_10559);
and U14054 (N_14054,N_10508,N_10857);
nand U14055 (N_14055,N_9735,N_9780);
nor U14056 (N_14056,N_11492,N_8629);
xor U14057 (N_14057,N_8094,N_9764);
or U14058 (N_14058,N_8845,N_11929);
and U14059 (N_14059,N_11360,N_9343);
nor U14060 (N_14060,N_8509,N_8743);
nand U14061 (N_14061,N_8923,N_10278);
or U14062 (N_14062,N_10816,N_8141);
and U14063 (N_14063,N_11856,N_11150);
nor U14064 (N_14064,N_9597,N_10894);
and U14065 (N_14065,N_10717,N_8467);
nor U14066 (N_14066,N_8064,N_11007);
and U14067 (N_14067,N_11655,N_9633);
nor U14068 (N_14068,N_10195,N_8892);
nor U14069 (N_14069,N_8045,N_8017);
nand U14070 (N_14070,N_9908,N_11865);
nor U14071 (N_14071,N_9573,N_9422);
nand U14072 (N_14072,N_8514,N_9075);
nand U14073 (N_14073,N_10422,N_8035);
xnor U14074 (N_14074,N_10160,N_9898);
xnor U14075 (N_14075,N_11845,N_11650);
nand U14076 (N_14076,N_9501,N_11949);
xor U14077 (N_14077,N_11647,N_11977);
and U14078 (N_14078,N_11749,N_9590);
or U14079 (N_14079,N_9013,N_11539);
nand U14080 (N_14080,N_9645,N_10181);
nor U14081 (N_14081,N_8386,N_8281);
and U14082 (N_14082,N_8881,N_10456);
nor U14083 (N_14083,N_10365,N_8722);
nand U14084 (N_14084,N_10113,N_8740);
xor U14085 (N_14085,N_8710,N_10503);
or U14086 (N_14086,N_11510,N_10419);
nand U14087 (N_14087,N_9536,N_9561);
or U14088 (N_14088,N_10524,N_8936);
and U14089 (N_14089,N_9048,N_9542);
xnor U14090 (N_14090,N_10443,N_10278);
and U14091 (N_14091,N_10316,N_11895);
and U14092 (N_14092,N_8197,N_10935);
or U14093 (N_14093,N_10327,N_10844);
nor U14094 (N_14094,N_11959,N_8666);
or U14095 (N_14095,N_9819,N_11503);
xnor U14096 (N_14096,N_11312,N_9372);
and U14097 (N_14097,N_11681,N_11265);
or U14098 (N_14098,N_11090,N_10273);
or U14099 (N_14099,N_9870,N_11390);
nor U14100 (N_14100,N_11082,N_9174);
nand U14101 (N_14101,N_9674,N_10538);
nand U14102 (N_14102,N_10729,N_8388);
nor U14103 (N_14103,N_9187,N_11229);
nand U14104 (N_14104,N_10412,N_8817);
nand U14105 (N_14105,N_10235,N_9993);
or U14106 (N_14106,N_11631,N_11296);
nor U14107 (N_14107,N_9110,N_8101);
xor U14108 (N_14108,N_8943,N_8917);
nor U14109 (N_14109,N_9869,N_11436);
and U14110 (N_14110,N_8676,N_9710);
and U14111 (N_14111,N_8102,N_8427);
and U14112 (N_14112,N_11576,N_9844);
nand U14113 (N_14113,N_8157,N_9337);
nor U14114 (N_14114,N_11962,N_9572);
and U14115 (N_14115,N_11877,N_10682);
or U14116 (N_14116,N_10951,N_9709);
nor U14117 (N_14117,N_8672,N_8616);
or U14118 (N_14118,N_10636,N_8319);
nor U14119 (N_14119,N_11930,N_9967);
and U14120 (N_14120,N_10103,N_9154);
or U14121 (N_14121,N_11291,N_11608);
and U14122 (N_14122,N_11325,N_10236);
nor U14123 (N_14123,N_10800,N_11086);
and U14124 (N_14124,N_10386,N_8933);
nand U14125 (N_14125,N_9310,N_8892);
xor U14126 (N_14126,N_10544,N_11174);
xor U14127 (N_14127,N_11071,N_8478);
nand U14128 (N_14128,N_11833,N_8354);
xnor U14129 (N_14129,N_10688,N_11106);
nand U14130 (N_14130,N_9850,N_9220);
or U14131 (N_14131,N_9155,N_9024);
nand U14132 (N_14132,N_9341,N_10212);
xor U14133 (N_14133,N_9944,N_11734);
nand U14134 (N_14134,N_8744,N_11884);
and U14135 (N_14135,N_11974,N_8105);
xor U14136 (N_14136,N_10971,N_10739);
nor U14137 (N_14137,N_11440,N_9522);
and U14138 (N_14138,N_9765,N_8364);
nor U14139 (N_14139,N_11733,N_10771);
or U14140 (N_14140,N_11732,N_9681);
nor U14141 (N_14141,N_8497,N_9608);
and U14142 (N_14142,N_11711,N_10055);
or U14143 (N_14143,N_10725,N_10739);
xnor U14144 (N_14144,N_8289,N_9532);
and U14145 (N_14145,N_8456,N_10232);
nor U14146 (N_14146,N_11163,N_11814);
nand U14147 (N_14147,N_10546,N_9467);
and U14148 (N_14148,N_8274,N_10814);
or U14149 (N_14149,N_10696,N_10474);
and U14150 (N_14150,N_9802,N_11421);
nor U14151 (N_14151,N_10308,N_9218);
or U14152 (N_14152,N_8206,N_10925);
and U14153 (N_14153,N_10026,N_11143);
nor U14154 (N_14154,N_9189,N_8072);
nor U14155 (N_14155,N_11072,N_10580);
xor U14156 (N_14156,N_11668,N_9808);
xnor U14157 (N_14157,N_9163,N_10855);
nand U14158 (N_14158,N_8417,N_9694);
or U14159 (N_14159,N_9454,N_10639);
nor U14160 (N_14160,N_10225,N_10617);
nand U14161 (N_14161,N_10380,N_10757);
and U14162 (N_14162,N_8987,N_10260);
or U14163 (N_14163,N_8544,N_11425);
nand U14164 (N_14164,N_9967,N_10367);
and U14165 (N_14165,N_11173,N_10166);
and U14166 (N_14166,N_8371,N_8828);
and U14167 (N_14167,N_9376,N_9388);
or U14168 (N_14168,N_11193,N_11815);
nand U14169 (N_14169,N_8520,N_10721);
xnor U14170 (N_14170,N_9585,N_10632);
or U14171 (N_14171,N_9557,N_10976);
xnor U14172 (N_14172,N_10108,N_8535);
and U14173 (N_14173,N_8410,N_11931);
nor U14174 (N_14174,N_8030,N_8667);
nor U14175 (N_14175,N_11529,N_11705);
and U14176 (N_14176,N_10276,N_11162);
or U14177 (N_14177,N_8888,N_11750);
nor U14178 (N_14178,N_10442,N_8560);
xnor U14179 (N_14179,N_11098,N_10928);
or U14180 (N_14180,N_8414,N_10112);
nor U14181 (N_14181,N_10370,N_11965);
nand U14182 (N_14182,N_10544,N_11687);
xor U14183 (N_14183,N_8483,N_11436);
and U14184 (N_14184,N_8305,N_11663);
or U14185 (N_14185,N_8501,N_10407);
and U14186 (N_14186,N_11187,N_9621);
nand U14187 (N_14187,N_8698,N_11543);
nor U14188 (N_14188,N_8575,N_11718);
xor U14189 (N_14189,N_10397,N_10893);
nor U14190 (N_14190,N_10309,N_8764);
xor U14191 (N_14191,N_11129,N_8627);
or U14192 (N_14192,N_8121,N_8733);
nor U14193 (N_14193,N_9076,N_10174);
xor U14194 (N_14194,N_10468,N_9487);
or U14195 (N_14195,N_8981,N_11580);
nand U14196 (N_14196,N_10404,N_8584);
or U14197 (N_14197,N_9013,N_8362);
and U14198 (N_14198,N_11303,N_9379);
or U14199 (N_14199,N_11606,N_11762);
and U14200 (N_14200,N_10772,N_10908);
nand U14201 (N_14201,N_11367,N_10564);
nor U14202 (N_14202,N_8488,N_9661);
and U14203 (N_14203,N_10035,N_11566);
and U14204 (N_14204,N_8088,N_10731);
or U14205 (N_14205,N_8303,N_9544);
and U14206 (N_14206,N_11882,N_11221);
nand U14207 (N_14207,N_8033,N_9999);
or U14208 (N_14208,N_9519,N_11089);
or U14209 (N_14209,N_10259,N_11273);
and U14210 (N_14210,N_8392,N_11055);
xor U14211 (N_14211,N_9586,N_11427);
or U14212 (N_14212,N_11485,N_11227);
and U14213 (N_14213,N_11826,N_9892);
nand U14214 (N_14214,N_11809,N_8071);
nand U14215 (N_14215,N_11957,N_9016);
nor U14216 (N_14216,N_8912,N_11941);
or U14217 (N_14217,N_10827,N_11242);
nand U14218 (N_14218,N_8481,N_10702);
or U14219 (N_14219,N_10230,N_8188);
or U14220 (N_14220,N_8166,N_10832);
and U14221 (N_14221,N_11128,N_11646);
and U14222 (N_14222,N_9368,N_10423);
nand U14223 (N_14223,N_8720,N_9964);
xnor U14224 (N_14224,N_9490,N_8508);
and U14225 (N_14225,N_9490,N_10582);
or U14226 (N_14226,N_10434,N_11120);
nor U14227 (N_14227,N_10782,N_11699);
or U14228 (N_14228,N_11526,N_8127);
and U14229 (N_14229,N_8856,N_8144);
nor U14230 (N_14230,N_11244,N_8291);
nor U14231 (N_14231,N_9339,N_9949);
and U14232 (N_14232,N_8151,N_9550);
and U14233 (N_14233,N_9238,N_10178);
or U14234 (N_14234,N_9385,N_10596);
or U14235 (N_14235,N_11892,N_10268);
and U14236 (N_14236,N_10921,N_11913);
nor U14237 (N_14237,N_10443,N_8197);
nand U14238 (N_14238,N_11607,N_10757);
xnor U14239 (N_14239,N_9264,N_10077);
xnor U14240 (N_14240,N_8551,N_8845);
or U14241 (N_14241,N_11972,N_9570);
xor U14242 (N_14242,N_11752,N_11380);
or U14243 (N_14243,N_8186,N_8050);
nor U14244 (N_14244,N_10484,N_11515);
or U14245 (N_14245,N_11060,N_10581);
nor U14246 (N_14246,N_10905,N_8979);
nor U14247 (N_14247,N_8515,N_11224);
or U14248 (N_14248,N_10281,N_9217);
nor U14249 (N_14249,N_9309,N_8976);
nor U14250 (N_14250,N_9252,N_8117);
or U14251 (N_14251,N_8892,N_8768);
and U14252 (N_14252,N_8433,N_11698);
and U14253 (N_14253,N_10768,N_11145);
nor U14254 (N_14254,N_9481,N_9228);
or U14255 (N_14255,N_10975,N_9904);
or U14256 (N_14256,N_8066,N_8334);
or U14257 (N_14257,N_10898,N_11489);
or U14258 (N_14258,N_8645,N_10421);
nor U14259 (N_14259,N_9493,N_9413);
or U14260 (N_14260,N_9951,N_11415);
and U14261 (N_14261,N_10301,N_11009);
or U14262 (N_14262,N_8977,N_8239);
nand U14263 (N_14263,N_9118,N_10100);
or U14264 (N_14264,N_9027,N_10029);
and U14265 (N_14265,N_9427,N_10957);
and U14266 (N_14266,N_8382,N_11948);
and U14267 (N_14267,N_9515,N_11867);
xnor U14268 (N_14268,N_9401,N_8459);
or U14269 (N_14269,N_8291,N_9089);
nand U14270 (N_14270,N_8165,N_11773);
nand U14271 (N_14271,N_10534,N_9672);
nand U14272 (N_14272,N_10830,N_10659);
nand U14273 (N_14273,N_8541,N_9671);
nand U14274 (N_14274,N_10112,N_11934);
nor U14275 (N_14275,N_10150,N_10405);
and U14276 (N_14276,N_11738,N_10227);
and U14277 (N_14277,N_9390,N_10483);
xnor U14278 (N_14278,N_11256,N_10454);
or U14279 (N_14279,N_10545,N_9101);
or U14280 (N_14280,N_9568,N_8513);
nor U14281 (N_14281,N_8923,N_8903);
nor U14282 (N_14282,N_11600,N_10368);
nand U14283 (N_14283,N_10050,N_9925);
nor U14284 (N_14284,N_8366,N_8160);
nor U14285 (N_14285,N_8126,N_8923);
nand U14286 (N_14286,N_11971,N_11924);
xnor U14287 (N_14287,N_11969,N_8291);
and U14288 (N_14288,N_10799,N_8926);
or U14289 (N_14289,N_8890,N_8196);
or U14290 (N_14290,N_10137,N_11871);
and U14291 (N_14291,N_11517,N_8220);
nand U14292 (N_14292,N_11043,N_10176);
and U14293 (N_14293,N_9030,N_8702);
nand U14294 (N_14294,N_10060,N_8472);
nand U14295 (N_14295,N_8711,N_9711);
xnor U14296 (N_14296,N_10222,N_9149);
nand U14297 (N_14297,N_10624,N_10937);
or U14298 (N_14298,N_9471,N_8405);
nand U14299 (N_14299,N_8837,N_11696);
nor U14300 (N_14300,N_11210,N_9844);
or U14301 (N_14301,N_9875,N_9992);
nand U14302 (N_14302,N_9301,N_10919);
nand U14303 (N_14303,N_11007,N_11215);
xnor U14304 (N_14304,N_9925,N_10069);
and U14305 (N_14305,N_9876,N_10949);
or U14306 (N_14306,N_9091,N_11831);
nor U14307 (N_14307,N_11210,N_8514);
and U14308 (N_14308,N_9594,N_8484);
nor U14309 (N_14309,N_11826,N_9908);
nand U14310 (N_14310,N_8842,N_11748);
or U14311 (N_14311,N_11024,N_9927);
or U14312 (N_14312,N_9739,N_10357);
and U14313 (N_14313,N_11917,N_8414);
and U14314 (N_14314,N_11403,N_9907);
nor U14315 (N_14315,N_10520,N_8406);
and U14316 (N_14316,N_11801,N_11044);
or U14317 (N_14317,N_11007,N_8143);
and U14318 (N_14318,N_10779,N_11611);
xor U14319 (N_14319,N_8165,N_8612);
nor U14320 (N_14320,N_8481,N_11803);
nor U14321 (N_14321,N_11246,N_10793);
or U14322 (N_14322,N_11758,N_10423);
or U14323 (N_14323,N_11262,N_8415);
xnor U14324 (N_14324,N_9226,N_11801);
and U14325 (N_14325,N_9861,N_10619);
or U14326 (N_14326,N_9789,N_9529);
or U14327 (N_14327,N_8876,N_10529);
and U14328 (N_14328,N_9914,N_8907);
or U14329 (N_14329,N_9714,N_10483);
or U14330 (N_14330,N_8757,N_9901);
xor U14331 (N_14331,N_11198,N_8783);
xnor U14332 (N_14332,N_8615,N_9752);
and U14333 (N_14333,N_9422,N_10577);
nor U14334 (N_14334,N_9815,N_11450);
nor U14335 (N_14335,N_10851,N_9734);
nand U14336 (N_14336,N_10930,N_9451);
and U14337 (N_14337,N_8943,N_10747);
or U14338 (N_14338,N_10156,N_11165);
nand U14339 (N_14339,N_11097,N_9210);
and U14340 (N_14340,N_11238,N_8605);
xor U14341 (N_14341,N_11947,N_10353);
nand U14342 (N_14342,N_8182,N_11359);
and U14343 (N_14343,N_9927,N_10006);
nor U14344 (N_14344,N_9323,N_8291);
or U14345 (N_14345,N_9735,N_10304);
and U14346 (N_14346,N_9345,N_10868);
and U14347 (N_14347,N_9718,N_8374);
nand U14348 (N_14348,N_8408,N_10882);
nor U14349 (N_14349,N_10726,N_11887);
nand U14350 (N_14350,N_8754,N_11570);
nand U14351 (N_14351,N_10049,N_11722);
nand U14352 (N_14352,N_10263,N_10795);
and U14353 (N_14353,N_10110,N_11577);
nor U14354 (N_14354,N_9301,N_8485);
xor U14355 (N_14355,N_9780,N_10494);
and U14356 (N_14356,N_9756,N_8204);
and U14357 (N_14357,N_11403,N_11321);
nor U14358 (N_14358,N_10768,N_11794);
nand U14359 (N_14359,N_10894,N_10660);
or U14360 (N_14360,N_10892,N_11991);
xor U14361 (N_14361,N_8034,N_8375);
and U14362 (N_14362,N_11532,N_9599);
or U14363 (N_14363,N_11915,N_11743);
nand U14364 (N_14364,N_10090,N_10368);
nor U14365 (N_14365,N_8229,N_9693);
and U14366 (N_14366,N_10038,N_11702);
xor U14367 (N_14367,N_11703,N_8610);
nor U14368 (N_14368,N_10964,N_11535);
nand U14369 (N_14369,N_11512,N_11496);
nand U14370 (N_14370,N_8408,N_10629);
nor U14371 (N_14371,N_10248,N_8257);
nor U14372 (N_14372,N_11097,N_11830);
nor U14373 (N_14373,N_10491,N_11430);
nand U14374 (N_14374,N_8045,N_10770);
and U14375 (N_14375,N_10959,N_11182);
xor U14376 (N_14376,N_8625,N_9350);
nand U14377 (N_14377,N_11237,N_8345);
nor U14378 (N_14378,N_11033,N_11844);
and U14379 (N_14379,N_10592,N_10144);
nand U14380 (N_14380,N_9014,N_9462);
nand U14381 (N_14381,N_10115,N_10970);
or U14382 (N_14382,N_11752,N_11496);
and U14383 (N_14383,N_10627,N_11329);
xor U14384 (N_14384,N_11956,N_8465);
or U14385 (N_14385,N_8933,N_11238);
nand U14386 (N_14386,N_9368,N_11646);
nor U14387 (N_14387,N_11211,N_8468);
nor U14388 (N_14388,N_11859,N_9423);
xor U14389 (N_14389,N_8511,N_10498);
and U14390 (N_14390,N_10500,N_9162);
nand U14391 (N_14391,N_8884,N_9071);
and U14392 (N_14392,N_9714,N_8500);
nand U14393 (N_14393,N_11355,N_8601);
nor U14394 (N_14394,N_8165,N_9138);
and U14395 (N_14395,N_11819,N_11770);
or U14396 (N_14396,N_11420,N_11514);
and U14397 (N_14397,N_8052,N_8279);
and U14398 (N_14398,N_8664,N_8509);
nor U14399 (N_14399,N_10339,N_10184);
nor U14400 (N_14400,N_11677,N_11556);
nand U14401 (N_14401,N_10874,N_11175);
or U14402 (N_14402,N_11365,N_9821);
and U14403 (N_14403,N_10353,N_10995);
xnor U14404 (N_14404,N_9178,N_11754);
nor U14405 (N_14405,N_8608,N_8044);
nand U14406 (N_14406,N_10955,N_10152);
and U14407 (N_14407,N_8205,N_10587);
nor U14408 (N_14408,N_10193,N_9479);
and U14409 (N_14409,N_8432,N_11458);
and U14410 (N_14410,N_9831,N_8634);
xnor U14411 (N_14411,N_9249,N_10516);
nor U14412 (N_14412,N_10336,N_11341);
and U14413 (N_14413,N_10069,N_10717);
and U14414 (N_14414,N_11552,N_9210);
nor U14415 (N_14415,N_9408,N_11860);
and U14416 (N_14416,N_10377,N_10389);
nor U14417 (N_14417,N_8392,N_8079);
nor U14418 (N_14418,N_10310,N_11165);
nand U14419 (N_14419,N_8027,N_11880);
nand U14420 (N_14420,N_9661,N_10257);
nor U14421 (N_14421,N_11134,N_8608);
and U14422 (N_14422,N_11060,N_9866);
nor U14423 (N_14423,N_11585,N_10152);
and U14424 (N_14424,N_11740,N_10419);
or U14425 (N_14425,N_9409,N_10029);
or U14426 (N_14426,N_10188,N_11585);
nor U14427 (N_14427,N_11345,N_8773);
or U14428 (N_14428,N_10723,N_10619);
or U14429 (N_14429,N_11542,N_9222);
or U14430 (N_14430,N_9336,N_11848);
or U14431 (N_14431,N_8127,N_10142);
or U14432 (N_14432,N_10185,N_8114);
and U14433 (N_14433,N_9632,N_10306);
or U14434 (N_14434,N_11870,N_10470);
xor U14435 (N_14435,N_11616,N_10159);
or U14436 (N_14436,N_11394,N_9159);
xor U14437 (N_14437,N_9631,N_8402);
and U14438 (N_14438,N_9390,N_10365);
or U14439 (N_14439,N_10348,N_11801);
xor U14440 (N_14440,N_11844,N_11864);
nor U14441 (N_14441,N_11721,N_11865);
nor U14442 (N_14442,N_9706,N_9958);
and U14443 (N_14443,N_11729,N_11855);
and U14444 (N_14444,N_9397,N_8878);
or U14445 (N_14445,N_9154,N_9136);
nand U14446 (N_14446,N_10219,N_8793);
xor U14447 (N_14447,N_9013,N_8008);
nor U14448 (N_14448,N_10908,N_11067);
nor U14449 (N_14449,N_11385,N_8231);
nand U14450 (N_14450,N_10591,N_11435);
or U14451 (N_14451,N_11244,N_8500);
or U14452 (N_14452,N_10835,N_8850);
nor U14453 (N_14453,N_8465,N_11174);
nor U14454 (N_14454,N_10138,N_10334);
nand U14455 (N_14455,N_8104,N_8265);
and U14456 (N_14456,N_11856,N_10047);
or U14457 (N_14457,N_9361,N_11310);
and U14458 (N_14458,N_8635,N_9272);
or U14459 (N_14459,N_8240,N_8829);
nor U14460 (N_14460,N_9560,N_9910);
nor U14461 (N_14461,N_8491,N_10138);
and U14462 (N_14462,N_8207,N_9121);
and U14463 (N_14463,N_10251,N_10522);
nor U14464 (N_14464,N_9981,N_10508);
nor U14465 (N_14465,N_10651,N_11591);
and U14466 (N_14466,N_8186,N_8061);
nand U14467 (N_14467,N_8334,N_8771);
nand U14468 (N_14468,N_10708,N_10631);
xnor U14469 (N_14469,N_8499,N_10409);
nor U14470 (N_14470,N_9920,N_8666);
and U14471 (N_14471,N_11813,N_9571);
nand U14472 (N_14472,N_9840,N_8947);
and U14473 (N_14473,N_8080,N_10456);
xnor U14474 (N_14474,N_11928,N_11965);
or U14475 (N_14475,N_10179,N_8735);
or U14476 (N_14476,N_8315,N_11528);
and U14477 (N_14477,N_9675,N_11578);
nor U14478 (N_14478,N_8386,N_11344);
xor U14479 (N_14479,N_8676,N_8845);
or U14480 (N_14480,N_10520,N_10588);
xor U14481 (N_14481,N_8332,N_11721);
and U14482 (N_14482,N_9040,N_10916);
nor U14483 (N_14483,N_11410,N_8096);
nor U14484 (N_14484,N_9845,N_8753);
nand U14485 (N_14485,N_10078,N_11746);
xnor U14486 (N_14486,N_8385,N_11800);
or U14487 (N_14487,N_10996,N_10613);
and U14488 (N_14488,N_8496,N_10066);
nor U14489 (N_14489,N_10246,N_11317);
or U14490 (N_14490,N_10195,N_10268);
xnor U14491 (N_14491,N_8227,N_8179);
or U14492 (N_14492,N_8699,N_9689);
or U14493 (N_14493,N_8984,N_11165);
nand U14494 (N_14494,N_11297,N_11541);
or U14495 (N_14495,N_9814,N_8785);
and U14496 (N_14496,N_9729,N_9022);
and U14497 (N_14497,N_8574,N_11785);
and U14498 (N_14498,N_8722,N_9442);
nor U14499 (N_14499,N_11309,N_9380);
or U14500 (N_14500,N_9603,N_10951);
and U14501 (N_14501,N_8156,N_8546);
or U14502 (N_14502,N_9790,N_9007);
nor U14503 (N_14503,N_9822,N_11801);
or U14504 (N_14504,N_8118,N_10911);
nor U14505 (N_14505,N_8331,N_8298);
xor U14506 (N_14506,N_11803,N_9351);
and U14507 (N_14507,N_11965,N_9313);
and U14508 (N_14508,N_9673,N_11489);
and U14509 (N_14509,N_9182,N_9473);
or U14510 (N_14510,N_10807,N_9064);
nand U14511 (N_14511,N_10704,N_8232);
nor U14512 (N_14512,N_11706,N_8381);
nor U14513 (N_14513,N_10633,N_9476);
and U14514 (N_14514,N_8359,N_10815);
nand U14515 (N_14515,N_11514,N_8677);
nor U14516 (N_14516,N_9329,N_9129);
or U14517 (N_14517,N_8581,N_8815);
nor U14518 (N_14518,N_10901,N_8705);
and U14519 (N_14519,N_9480,N_8096);
or U14520 (N_14520,N_9801,N_8521);
and U14521 (N_14521,N_11937,N_10245);
nand U14522 (N_14522,N_9654,N_9615);
or U14523 (N_14523,N_10550,N_10374);
nor U14524 (N_14524,N_9123,N_8505);
nor U14525 (N_14525,N_11048,N_11331);
and U14526 (N_14526,N_9870,N_9250);
and U14527 (N_14527,N_10672,N_9903);
or U14528 (N_14528,N_9967,N_8396);
and U14529 (N_14529,N_10163,N_8142);
or U14530 (N_14530,N_9376,N_10517);
nor U14531 (N_14531,N_11901,N_11128);
and U14532 (N_14532,N_8455,N_9470);
and U14533 (N_14533,N_9321,N_11021);
or U14534 (N_14534,N_8160,N_8589);
nor U14535 (N_14535,N_8245,N_9479);
xnor U14536 (N_14536,N_9139,N_8449);
nand U14537 (N_14537,N_8115,N_11155);
and U14538 (N_14538,N_10179,N_10903);
or U14539 (N_14539,N_8358,N_10220);
nor U14540 (N_14540,N_9564,N_9473);
nor U14541 (N_14541,N_11582,N_8882);
or U14542 (N_14542,N_10731,N_8598);
nor U14543 (N_14543,N_10483,N_9314);
nand U14544 (N_14544,N_8249,N_8290);
or U14545 (N_14545,N_10793,N_8323);
and U14546 (N_14546,N_11517,N_10187);
and U14547 (N_14547,N_8304,N_8539);
xnor U14548 (N_14548,N_8028,N_10655);
nor U14549 (N_14549,N_8123,N_10407);
nor U14550 (N_14550,N_11452,N_9172);
and U14551 (N_14551,N_10550,N_9763);
or U14552 (N_14552,N_9638,N_9498);
or U14553 (N_14553,N_10719,N_8394);
nand U14554 (N_14554,N_11773,N_10737);
nor U14555 (N_14555,N_9735,N_10389);
or U14556 (N_14556,N_8003,N_9241);
xnor U14557 (N_14557,N_10070,N_8374);
nor U14558 (N_14558,N_10300,N_10539);
nand U14559 (N_14559,N_8945,N_9822);
and U14560 (N_14560,N_10786,N_9169);
or U14561 (N_14561,N_10032,N_8616);
and U14562 (N_14562,N_8036,N_11037);
and U14563 (N_14563,N_8958,N_8217);
nand U14564 (N_14564,N_8314,N_9699);
nand U14565 (N_14565,N_8319,N_11218);
and U14566 (N_14566,N_10748,N_8934);
or U14567 (N_14567,N_8365,N_9203);
nand U14568 (N_14568,N_9588,N_10968);
nand U14569 (N_14569,N_11408,N_8626);
or U14570 (N_14570,N_10043,N_10928);
or U14571 (N_14571,N_8610,N_8192);
xnor U14572 (N_14572,N_10124,N_9377);
nor U14573 (N_14573,N_9099,N_9164);
nand U14574 (N_14574,N_8846,N_9674);
and U14575 (N_14575,N_10598,N_10778);
nand U14576 (N_14576,N_8148,N_10430);
xnor U14577 (N_14577,N_8412,N_10127);
and U14578 (N_14578,N_9639,N_11627);
nor U14579 (N_14579,N_8901,N_9830);
or U14580 (N_14580,N_10064,N_8139);
or U14581 (N_14581,N_9090,N_11248);
nor U14582 (N_14582,N_11733,N_9134);
and U14583 (N_14583,N_10326,N_10221);
and U14584 (N_14584,N_8923,N_8781);
nor U14585 (N_14585,N_8603,N_11525);
or U14586 (N_14586,N_10541,N_8361);
nor U14587 (N_14587,N_11423,N_9560);
nand U14588 (N_14588,N_9885,N_8918);
or U14589 (N_14589,N_11020,N_10565);
nor U14590 (N_14590,N_10968,N_11290);
and U14591 (N_14591,N_10251,N_10000);
nor U14592 (N_14592,N_11602,N_10649);
nand U14593 (N_14593,N_11754,N_10412);
or U14594 (N_14594,N_10428,N_8453);
nand U14595 (N_14595,N_8768,N_11086);
or U14596 (N_14596,N_11462,N_10320);
nor U14597 (N_14597,N_10935,N_9912);
and U14598 (N_14598,N_10305,N_8043);
and U14599 (N_14599,N_9072,N_11878);
nor U14600 (N_14600,N_11937,N_11678);
nor U14601 (N_14601,N_11404,N_8514);
nor U14602 (N_14602,N_10197,N_10209);
nor U14603 (N_14603,N_10795,N_8706);
xnor U14604 (N_14604,N_9959,N_10420);
xor U14605 (N_14605,N_10048,N_10861);
xnor U14606 (N_14606,N_9959,N_9445);
xor U14607 (N_14607,N_8733,N_10073);
nor U14608 (N_14608,N_11715,N_9928);
xnor U14609 (N_14609,N_9092,N_9925);
or U14610 (N_14610,N_8823,N_8354);
nor U14611 (N_14611,N_8655,N_8000);
and U14612 (N_14612,N_8528,N_9443);
nand U14613 (N_14613,N_8489,N_10300);
nor U14614 (N_14614,N_9106,N_11738);
and U14615 (N_14615,N_10911,N_8135);
nand U14616 (N_14616,N_9826,N_9100);
and U14617 (N_14617,N_8304,N_8061);
nor U14618 (N_14618,N_8013,N_11536);
or U14619 (N_14619,N_8847,N_8020);
nor U14620 (N_14620,N_8140,N_8228);
or U14621 (N_14621,N_9664,N_8871);
nor U14622 (N_14622,N_9585,N_10996);
nor U14623 (N_14623,N_11944,N_10373);
and U14624 (N_14624,N_11235,N_10613);
nor U14625 (N_14625,N_9545,N_9396);
or U14626 (N_14626,N_9876,N_9259);
xnor U14627 (N_14627,N_8089,N_10281);
and U14628 (N_14628,N_8874,N_11479);
nor U14629 (N_14629,N_9181,N_9548);
and U14630 (N_14630,N_8081,N_11842);
nor U14631 (N_14631,N_10584,N_8576);
nand U14632 (N_14632,N_11078,N_11990);
and U14633 (N_14633,N_9224,N_9620);
nor U14634 (N_14634,N_8942,N_10097);
and U14635 (N_14635,N_8368,N_10248);
nor U14636 (N_14636,N_10485,N_9902);
and U14637 (N_14637,N_9574,N_10043);
nor U14638 (N_14638,N_11138,N_8754);
and U14639 (N_14639,N_8928,N_8573);
nand U14640 (N_14640,N_8651,N_9764);
xnor U14641 (N_14641,N_11705,N_10819);
and U14642 (N_14642,N_8162,N_10642);
nor U14643 (N_14643,N_8393,N_10242);
and U14644 (N_14644,N_10166,N_10533);
or U14645 (N_14645,N_8507,N_8096);
nand U14646 (N_14646,N_8062,N_8738);
or U14647 (N_14647,N_11788,N_11554);
or U14648 (N_14648,N_10678,N_11637);
nand U14649 (N_14649,N_10007,N_9037);
or U14650 (N_14650,N_10758,N_9004);
nor U14651 (N_14651,N_10976,N_10638);
nor U14652 (N_14652,N_10581,N_11986);
nor U14653 (N_14653,N_9790,N_10445);
or U14654 (N_14654,N_9314,N_11010);
or U14655 (N_14655,N_8225,N_8035);
or U14656 (N_14656,N_11171,N_10220);
or U14657 (N_14657,N_8741,N_9769);
and U14658 (N_14658,N_10657,N_10897);
nor U14659 (N_14659,N_10994,N_8848);
nor U14660 (N_14660,N_10303,N_8357);
nand U14661 (N_14661,N_11857,N_8683);
nand U14662 (N_14662,N_8605,N_9837);
nor U14663 (N_14663,N_9259,N_11069);
nand U14664 (N_14664,N_9034,N_11471);
nand U14665 (N_14665,N_9141,N_11159);
nor U14666 (N_14666,N_9568,N_8365);
and U14667 (N_14667,N_10555,N_11471);
nor U14668 (N_14668,N_8022,N_8051);
nor U14669 (N_14669,N_8403,N_10459);
or U14670 (N_14670,N_10563,N_11234);
or U14671 (N_14671,N_9192,N_8779);
xor U14672 (N_14672,N_9155,N_8429);
nand U14673 (N_14673,N_11553,N_10861);
and U14674 (N_14674,N_8177,N_8647);
nor U14675 (N_14675,N_9024,N_9422);
nand U14676 (N_14676,N_10275,N_9007);
nor U14677 (N_14677,N_10328,N_9821);
nor U14678 (N_14678,N_9990,N_11852);
and U14679 (N_14679,N_9364,N_8134);
nand U14680 (N_14680,N_10610,N_11990);
nand U14681 (N_14681,N_8298,N_9431);
nor U14682 (N_14682,N_9800,N_11613);
nor U14683 (N_14683,N_11842,N_8713);
nand U14684 (N_14684,N_10539,N_8566);
nor U14685 (N_14685,N_11564,N_11489);
xor U14686 (N_14686,N_9711,N_8014);
xnor U14687 (N_14687,N_9306,N_11661);
or U14688 (N_14688,N_11326,N_9025);
and U14689 (N_14689,N_10168,N_8615);
nand U14690 (N_14690,N_10534,N_10720);
or U14691 (N_14691,N_8391,N_10512);
and U14692 (N_14692,N_10797,N_10165);
nor U14693 (N_14693,N_8019,N_8001);
nand U14694 (N_14694,N_9520,N_8009);
nand U14695 (N_14695,N_8519,N_9302);
nand U14696 (N_14696,N_8605,N_8292);
or U14697 (N_14697,N_11222,N_8777);
nor U14698 (N_14698,N_9047,N_8281);
or U14699 (N_14699,N_8130,N_8719);
or U14700 (N_14700,N_8333,N_11056);
nor U14701 (N_14701,N_9847,N_8996);
or U14702 (N_14702,N_8135,N_9903);
xnor U14703 (N_14703,N_10826,N_9201);
nand U14704 (N_14704,N_9852,N_11508);
and U14705 (N_14705,N_10172,N_8034);
or U14706 (N_14706,N_8927,N_9165);
and U14707 (N_14707,N_10642,N_11113);
nand U14708 (N_14708,N_9656,N_11572);
and U14709 (N_14709,N_10083,N_10304);
and U14710 (N_14710,N_11495,N_11716);
and U14711 (N_14711,N_11873,N_10582);
or U14712 (N_14712,N_10036,N_11117);
nand U14713 (N_14713,N_10563,N_10304);
nand U14714 (N_14714,N_11593,N_8456);
xor U14715 (N_14715,N_11194,N_10030);
nand U14716 (N_14716,N_8695,N_10244);
or U14717 (N_14717,N_11557,N_11489);
nand U14718 (N_14718,N_10993,N_9286);
or U14719 (N_14719,N_8049,N_11170);
nand U14720 (N_14720,N_10613,N_11682);
nand U14721 (N_14721,N_10355,N_11966);
nand U14722 (N_14722,N_9419,N_9266);
nor U14723 (N_14723,N_11682,N_8174);
and U14724 (N_14724,N_8681,N_10796);
nor U14725 (N_14725,N_9716,N_10277);
and U14726 (N_14726,N_8787,N_10021);
nand U14727 (N_14727,N_10758,N_9145);
nand U14728 (N_14728,N_11666,N_8255);
or U14729 (N_14729,N_9749,N_11460);
and U14730 (N_14730,N_9046,N_9156);
nand U14731 (N_14731,N_11852,N_8293);
nand U14732 (N_14732,N_11225,N_8002);
and U14733 (N_14733,N_8828,N_9245);
and U14734 (N_14734,N_8737,N_9805);
xnor U14735 (N_14735,N_8782,N_8183);
or U14736 (N_14736,N_11392,N_9785);
or U14737 (N_14737,N_8238,N_9408);
xnor U14738 (N_14738,N_10138,N_10061);
nor U14739 (N_14739,N_9863,N_8437);
nand U14740 (N_14740,N_8129,N_9469);
or U14741 (N_14741,N_11686,N_10028);
nand U14742 (N_14742,N_11916,N_10197);
xor U14743 (N_14743,N_8315,N_9402);
nand U14744 (N_14744,N_10502,N_8667);
nand U14745 (N_14745,N_8040,N_9453);
nor U14746 (N_14746,N_10655,N_8136);
or U14747 (N_14747,N_11774,N_9744);
or U14748 (N_14748,N_11715,N_8006);
nor U14749 (N_14749,N_10237,N_9664);
nor U14750 (N_14750,N_11501,N_9643);
or U14751 (N_14751,N_8339,N_8609);
or U14752 (N_14752,N_11228,N_11312);
nand U14753 (N_14753,N_10200,N_8685);
and U14754 (N_14754,N_10690,N_11159);
nand U14755 (N_14755,N_10610,N_11901);
and U14756 (N_14756,N_10297,N_8980);
nand U14757 (N_14757,N_9789,N_8290);
nor U14758 (N_14758,N_8071,N_10424);
and U14759 (N_14759,N_10647,N_11510);
nor U14760 (N_14760,N_8778,N_9492);
and U14761 (N_14761,N_9302,N_8878);
and U14762 (N_14762,N_11368,N_10842);
and U14763 (N_14763,N_9861,N_11331);
xor U14764 (N_14764,N_11279,N_9668);
or U14765 (N_14765,N_11961,N_11692);
nand U14766 (N_14766,N_10248,N_9715);
or U14767 (N_14767,N_11456,N_10675);
or U14768 (N_14768,N_8988,N_11991);
and U14769 (N_14769,N_11743,N_9616);
or U14770 (N_14770,N_10778,N_8845);
nand U14771 (N_14771,N_9012,N_9586);
or U14772 (N_14772,N_8966,N_8359);
nor U14773 (N_14773,N_9451,N_10700);
or U14774 (N_14774,N_8652,N_10434);
nor U14775 (N_14775,N_10031,N_11513);
nor U14776 (N_14776,N_11389,N_11212);
xnor U14777 (N_14777,N_8228,N_11241);
nand U14778 (N_14778,N_11253,N_8719);
xnor U14779 (N_14779,N_8645,N_11223);
and U14780 (N_14780,N_10168,N_9143);
xor U14781 (N_14781,N_11994,N_9783);
nor U14782 (N_14782,N_11623,N_11795);
nand U14783 (N_14783,N_8223,N_11067);
nand U14784 (N_14784,N_8334,N_9585);
nand U14785 (N_14785,N_8300,N_8363);
nor U14786 (N_14786,N_11503,N_10637);
and U14787 (N_14787,N_11661,N_9945);
or U14788 (N_14788,N_8493,N_9228);
xor U14789 (N_14789,N_11450,N_11279);
and U14790 (N_14790,N_10943,N_8838);
nand U14791 (N_14791,N_11646,N_8936);
nor U14792 (N_14792,N_9106,N_11542);
and U14793 (N_14793,N_11110,N_8194);
or U14794 (N_14794,N_10596,N_8319);
or U14795 (N_14795,N_11229,N_9782);
and U14796 (N_14796,N_8914,N_10377);
and U14797 (N_14797,N_10086,N_10679);
nand U14798 (N_14798,N_11098,N_11032);
or U14799 (N_14799,N_8962,N_8507);
and U14800 (N_14800,N_8616,N_8430);
or U14801 (N_14801,N_8128,N_9110);
nor U14802 (N_14802,N_10914,N_9534);
or U14803 (N_14803,N_10054,N_10311);
nor U14804 (N_14804,N_8368,N_11853);
and U14805 (N_14805,N_10666,N_11467);
xor U14806 (N_14806,N_11257,N_9951);
nand U14807 (N_14807,N_10115,N_9602);
or U14808 (N_14808,N_9062,N_8121);
and U14809 (N_14809,N_11417,N_11551);
nand U14810 (N_14810,N_9327,N_8228);
xor U14811 (N_14811,N_9483,N_11030);
and U14812 (N_14812,N_8947,N_10560);
nor U14813 (N_14813,N_11458,N_11465);
nand U14814 (N_14814,N_10947,N_8160);
nand U14815 (N_14815,N_10972,N_8140);
or U14816 (N_14816,N_9632,N_10505);
or U14817 (N_14817,N_9471,N_8869);
or U14818 (N_14818,N_11322,N_9488);
nand U14819 (N_14819,N_11446,N_11403);
nand U14820 (N_14820,N_8889,N_8231);
or U14821 (N_14821,N_10779,N_10954);
or U14822 (N_14822,N_11404,N_9919);
and U14823 (N_14823,N_9631,N_8311);
nand U14824 (N_14824,N_10237,N_9414);
nand U14825 (N_14825,N_10197,N_9007);
xnor U14826 (N_14826,N_9568,N_8444);
xnor U14827 (N_14827,N_11086,N_9698);
and U14828 (N_14828,N_8248,N_8524);
or U14829 (N_14829,N_9507,N_9629);
xor U14830 (N_14830,N_9561,N_10536);
nand U14831 (N_14831,N_10291,N_9447);
and U14832 (N_14832,N_9856,N_11986);
and U14833 (N_14833,N_11451,N_8012);
or U14834 (N_14834,N_10842,N_9396);
xnor U14835 (N_14835,N_10499,N_10390);
and U14836 (N_14836,N_8615,N_9017);
nand U14837 (N_14837,N_10846,N_11360);
or U14838 (N_14838,N_8446,N_10006);
nand U14839 (N_14839,N_11710,N_9753);
nand U14840 (N_14840,N_10646,N_11451);
xor U14841 (N_14841,N_8393,N_10385);
and U14842 (N_14842,N_8687,N_8293);
nor U14843 (N_14843,N_11911,N_11320);
or U14844 (N_14844,N_10602,N_8686);
and U14845 (N_14845,N_11025,N_9187);
nand U14846 (N_14846,N_8834,N_10472);
xor U14847 (N_14847,N_10113,N_9805);
nor U14848 (N_14848,N_9061,N_9226);
or U14849 (N_14849,N_11539,N_10216);
nand U14850 (N_14850,N_9661,N_11564);
nand U14851 (N_14851,N_8266,N_11679);
nor U14852 (N_14852,N_9712,N_8023);
xor U14853 (N_14853,N_10416,N_9988);
nand U14854 (N_14854,N_8280,N_9122);
or U14855 (N_14855,N_9017,N_9743);
nor U14856 (N_14856,N_10179,N_9276);
nor U14857 (N_14857,N_10686,N_8636);
and U14858 (N_14858,N_11951,N_10379);
nor U14859 (N_14859,N_9718,N_10461);
or U14860 (N_14860,N_8846,N_11685);
xnor U14861 (N_14861,N_10440,N_8898);
and U14862 (N_14862,N_11649,N_11226);
nor U14863 (N_14863,N_8925,N_9882);
and U14864 (N_14864,N_9549,N_8228);
nor U14865 (N_14865,N_10613,N_9060);
and U14866 (N_14866,N_10654,N_8793);
nand U14867 (N_14867,N_10717,N_10994);
nor U14868 (N_14868,N_11839,N_10917);
or U14869 (N_14869,N_11451,N_10949);
or U14870 (N_14870,N_11142,N_11151);
nand U14871 (N_14871,N_9478,N_11462);
nand U14872 (N_14872,N_8875,N_11329);
or U14873 (N_14873,N_9803,N_8377);
nor U14874 (N_14874,N_8150,N_11373);
and U14875 (N_14875,N_10113,N_8454);
or U14876 (N_14876,N_11368,N_8340);
nand U14877 (N_14877,N_9996,N_8467);
nand U14878 (N_14878,N_10391,N_8625);
or U14879 (N_14879,N_8858,N_10431);
and U14880 (N_14880,N_10384,N_8783);
or U14881 (N_14881,N_9515,N_8910);
xnor U14882 (N_14882,N_10950,N_8679);
or U14883 (N_14883,N_11317,N_11448);
nand U14884 (N_14884,N_8135,N_10675);
nor U14885 (N_14885,N_9185,N_9968);
nand U14886 (N_14886,N_10218,N_9337);
and U14887 (N_14887,N_8432,N_11681);
nand U14888 (N_14888,N_8283,N_9978);
or U14889 (N_14889,N_10211,N_10108);
and U14890 (N_14890,N_9833,N_8685);
xor U14891 (N_14891,N_11041,N_9884);
and U14892 (N_14892,N_8172,N_11303);
or U14893 (N_14893,N_11991,N_11648);
and U14894 (N_14894,N_9211,N_9034);
and U14895 (N_14895,N_10003,N_8130);
or U14896 (N_14896,N_9765,N_10481);
or U14897 (N_14897,N_10803,N_11459);
nor U14898 (N_14898,N_9683,N_10258);
nand U14899 (N_14899,N_8697,N_10874);
or U14900 (N_14900,N_11669,N_9005);
nor U14901 (N_14901,N_8667,N_11776);
nor U14902 (N_14902,N_9703,N_10979);
and U14903 (N_14903,N_10374,N_8494);
nor U14904 (N_14904,N_8842,N_8738);
nand U14905 (N_14905,N_10058,N_8331);
nor U14906 (N_14906,N_9282,N_10641);
and U14907 (N_14907,N_8157,N_11261);
nand U14908 (N_14908,N_10887,N_9788);
xnor U14909 (N_14909,N_11307,N_9734);
and U14910 (N_14910,N_10397,N_8298);
nand U14911 (N_14911,N_11282,N_11084);
nand U14912 (N_14912,N_9119,N_10206);
or U14913 (N_14913,N_9374,N_8140);
nor U14914 (N_14914,N_11545,N_9684);
or U14915 (N_14915,N_11567,N_8664);
nand U14916 (N_14916,N_10711,N_8154);
and U14917 (N_14917,N_9715,N_11939);
or U14918 (N_14918,N_8695,N_11529);
nor U14919 (N_14919,N_9216,N_10123);
nor U14920 (N_14920,N_8115,N_11209);
or U14921 (N_14921,N_10783,N_8453);
and U14922 (N_14922,N_9308,N_8746);
nor U14923 (N_14923,N_8339,N_9735);
nor U14924 (N_14924,N_11371,N_9806);
nand U14925 (N_14925,N_8258,N_9607);
nor U14926 (N_14926,N_11912,N_9616);
or U14927 (N_14927,N_11143,N_8468);
and U14928 (N_14928,N_11902,N_8538);
nand U14929 (N_14929,N_11012,N_8044);
xor U14930 (N_14930,N_10658,N_8412);
nand U14931 (N_14931,N_9278,N_10632);
and U14932 (N_14932,N_10958,N_8840);
and U14933 (N_14933,N_10927,N_9842);
nor U14934 (N_14934,N_9871,N_11204);
xnor U14935 (N_14935,N_10125,N_10009);
nand U14936 (N_14936,N_8504,N_10970);
nand U14937 (N_14937,N_8677,N_11496);
nand U14938 (N_14938,N_8386,N_11551);
xor U14939 (N_14939,N_8072,N_11405);
xor U14940 (N_14940,N_10178,N_11070);
nand U14941 (N_14941,N_8447,N_8563);
nand U14942 (N_14942,N_11440,N_9670);
or U14943 (N_14943,N_8076,N_10023);
nand U14944 (N_14944,N_9454,N_8567);
nand U14945 (N_14945,N_9992,N_9989);
or U14946 (N_14946,N_9489,N_10697);
nand U14947 (N_14947,N_11686,N_10258);
nand U14948 (N_14948,N_11370,N_8811);
nor U14949 (N_14949,N_10968,N_11224);
and U14950 (N_14950,N_8833,N_11727);
and U14951 (N_14951,N_8047,N_11779);
nand U14952 (N_14952,N_11425,N_8302);
and U14953 (N_14953,N_9682,N_9563);
and U14954 (N_14954,N_10447,N_11251);
or U14955 (N_14955,N_8871,N_9037);
nand U14956 (N_14956,N_11846,N_10605);
nand U14957 (N_14957,N_9756,N_8951);
or U14958 (N_14958,N_10589,N_10647);
or U14959 (N_14959,N_8826,N_9088);
nor U14960 (N_14960,N_10510,N_8437);
nor U14961 (N_14961,N_11958,N_9448);
xnor U14962 (N_14962,N_10607,N_9825);
nor U14963 (N_14963,N_10101,N_8527);
nor U14964 (N_14964,N_10250,N_11175);
nand U14965 (N_14965,N_8386,N_11217);
and U14966 (N_14966,N_8884,N_9017);
nor U14967 (N_14967,N_8858,N_9748);
nand U14968 (N_14968,N_10091,N_11341);
and U14969 (N_14969,N_8170,N_10882);
xnor U14970 (N_14970,N_9852,N_9374);
xnor U14971 (N_14971,N_10284,N_10215);
and U14972 (N_14972,N_9362,N_8117);
and U14973 (N_14973,N_9324,N_10400);
or U14974 (N_14974,N_10974,N_9084);
or U14975 (N_14975,N_9994,N_9264);
and U14976 (N_14976,N_8879,N_8021);
xnor U14977 (N_14977,N_10741,N_11971);
xnor U14978 (N_14978,N_10314,N_8555);
nor U14979 (N_14979,N_9603,N_9482);
nand U14980 (N_14980,N_8857,N_11290);
nand U14981 (N_14981,N_8893,N_9222);
and U14982 (N_14982,N_10266,N_9261);
or U14983 (N_14983,N_8353,N_9160);
nor U14984 (N_14984,N_10489,N_8060);
nor U14985 (N_14985,N_10694,N_9635);
nor U14986 (N_14986,N_9673,N_10256);
or U14987 (N_14987,N_10895,N_10510);
nand U14988 (N_14988,N_8634,N_11022);
and U14989 (N_14989,N_9715,N_10386);
nor U14990 (N_14990,N_8792,N_9162);
and U14991 (N_14991,N_10622,N_11746);
nand U14992 (N_14992,N_10029,N_11139);
or U14993 (N_14993,N_10922,N_11943);
or U14994 (N_14994,N_11159,N_10117);
nor U14995 (N_14995,N_11345,N_11753);
nand U14996 (N_14996,N_9798,N_11728);
xor U14997 (N_14997,N_8089,N_11956);
nor U14998 (N_14998,N_9254,N_10091);
nand U14999 (N_14999,N_8383,N_9769);
or U15000 (N_15000,N_8842,N_9103);
nand U15001 (N_15001,N_11098,N_9930);
and U15002 (N_15002,N_8214,N_8885);
or U15003 (N_15003,N_9959,N_9836);
nor U15004 (N_15004,N_9027,N_8830);
nand U15005 (N_15005,N_10886,N_9731);
nand U15006 (N_15006,N_11385,N_10073);
nor U15007 (N_15007,N_10731,N_10148);
nor U15008 (N_15008,N_9698,N_8087);
nor U15009 (N_15009,N_8686,N_9387);
or U15010 (N_15010,N_11718,N_8897);
nor U15011 (N_15011,N_9922,N_10932);
nor U15012 (N_15012,N_8169,N_8076);
or U15013 (N_15013,N_8395,N_9440);
xor U15014 (N_15014,N_9850,N_8713);
or U15015 (N_15015,N_9850,N_11412);
and U15016 (N_15016,N_8427,N_10253);
nand U15017 (N_15017,N_8507,N_8219);
nor U15018 (N_15018,N_11461,N_10473);
xnor U15019 (N_15019,N_10858,N_8480);
xnor U15020 (N_15020,N_8691,N_9053);
and U15021 (N_15021,N_9060,N_11810);
nor U15022 (N_15022,N_8728,N_8209);
nand U15023 (N_15023,N_9405,N_11909);
nor U15024 (N_15024,N_11872,N_11250);
xnor U15025 (N_15025,N_10311,N_8242);
nand U15026 (N_15026,N_11643,N_10972);
xor U15027 (N_15027,N_8379,N_9492);
nand U15028 (N_15028,N_11227,N_8336);
nor U15029 (N_15029,N_8368,N_9407);
and U15030 (N_15030,N_11533,N_10109);
nor U15031 (N_15031,N_11425,N_11487);
nand U15032 (N_15032,N_11717,N_10896);
nand U15033 (N_15033,N_10290,N_8002);
nor U15034 (N_15034,N_11620,N_11811);
and U15035 (N_15035,N_9136,N_9191);
and U15036 (N_15036,N_8301,N_9785);
nand U15037 (N_15037,N_8088,N_10682);
and U15038 (N_15038,N_8654,N_9374);
nand U15039 (N_15039,N_9264,N_10336);
nor U15040 (N_15040,N_10944,N_9984);
or U15041 (N_15041,N_9326,N_8680);
nor U15042 (N_15042,N_10298,N_9498);
nand U15043 (N_15043,N_9899,N_11242);
or U15044 (N_15044,N_10707,N_9035);
or U15045 (N_15045,N_10561,N_9707);
nand U15046 (N_15046,N_9978,N_11933);
and U15047 (N_15047,N_8503,N_10956);
and U15048 (N_15048,N_11875,N_9240);
and U15049 (N_15049,N_10288,N_9041);
and U15050 (N_15050,N_11309,N_8548);
nand U15051 (N_15051,N_10550,N_11393);
nor U15052 (N_15052,N_9371,N_11564);
or U15053 (N_15053,N_11984,N_9114);
nor U15054 (N_15054,N_10913,N_10370);
or U15055 (N_15055,N_10769,N_8408);
nand U15056 (N_15056,N_8458,N_8419);
and U15057 (N_15057,N_8508,N_9412);
and U15058 (N_15058,N_8263,N_11121);
and U15059 (N_15059,N_10104,N_10849);
or U15060 (N_15060,N_8215,N_10717);
nand U15061 (N_15061,N_8057,N_11695);
nor U15062 (N_15062,N_9814,N_9173);
and U15063 (N_15063,N_11172,N_9505);
or U15064 (N_15064,N_11197,N_8204);
nor U15065 (N_15065,N_8934,N_8761);
or U15066 (N_15066,N_8999,N_8496);
and U15067 (N_15067,N_11525,N_10069);
nor U15068 (N_15068,N_9082,N_8125);
or U15069 (N_15069,N_11297,N_11670);
and U15070 (N_15070,N_8167,N_9447);
or U15071 (N_15071,N_9605,N_8516);
or U15072 (N_15072,N_10801,N_11049);
nor U15073 (N_15073,N_10572,N_11067);
and U15074 (N_15074,N_10324,N_10784);
or U15075 (N_15075,N_9742,N_8696);
nor U15076 (N_15076,N_9836,N_11371);
nor U15077 (N_15077,N_8793,N_9913);
or U15078 (N_15078,N_9239,N_8238);
nand U15079 (N_15079,N_10154,N_10802);
nor U15080 (N_15080,N_9033,N_9626);
nor U15081 (N_15081,N_10672,N_10522);
or U15082 (N_15082,N_8228,N_9068);
nor U15083 (N_15083,N_8657,N_9928);
or U15084 (N_15084,N_8255,N_8060);
nand U15085 (N_15085,N_9733,N_9739);
xor U15086 (N_15086,N_8314,N_10801);
nor U15087 (N_15087,N_11649,N_11704);
or U15088 (N_15088,N_10980,N_9230);
or U15089 (N_15089,N_10271,N_10900);
and U15090 (N_15090,N_10199,N_11073);
nand U15091 (N_15091,N_8695,N_9819);
xor U15092 (N_15092,N_9089,N_9897);
nor U15093 (N_15093,N_11712,N_9110);
nor U15094 (N_15094,N_9275,N_10437);
and U15095 (N_15095,N_8977,N_10948);
and U15096 (N_15096,N_9397,N_9919);
or U15097 (N_15097,N_8952,N_11500);
or U15098 (N_15098,N_10619,N_11476);
or U15099 (N_15099,N_8260,N_11906);
and U15100 (N_15100,N_9630,N_11528);
nand U15101 (N_15101,N_10456,N_8160);
nor U15102 (N_15102,N_9591,N_10322);
or U15103 (N_15103,N_11778,N_11246);
and U15104 (N_15104,N_8788,N_9589);
and U15105 (N_15105,N_11308,N_9790);
and U15106 (N_15106,N_10693,N_11769);
and U15107 (N_15107,N_9950,N_9587);
or U15108 (N_15108,N_10370,N_9307);
nor U15109 (N_15109,N_8944,N_9808);
or U15110 (N_15110,N_8696,N_11609);
nand U15111 (N_15111,N_9881,N_9439);
and U15112 (N_15112,N_10264,N_9955);
nor U15113 (N_15113,N_11457,N_10857);
and U15114 (N_15114,N_11932,N_9473);
nand U15115 (N_15115,N_11446,N_8706);
xnor U15116 (N_15116,N_8101,N_10043);
nand U15117 (N_15117,N_10442,N_10156);
nand U15118 (N_15118,N_9773,N_10151);
and U15119 (N_15119,N_10767,N_11112);
nor U15120 (N_15120,N_9182,N_9693);
and U15121 (N_15121,N_11236,N_9907);
nand U15122 (N_15122,N_10711,N_8115);
or U15123 (N_15123,N_11786,N_10540);
or U15124 (N_15124,N_11833,N_10273);
nand U15125 (N_15125,N_11770,N_11470);
and U15126 (N_15126,N_9303,N_8576);
or U15127 (N_15127,N_8295,N_8201);
or U15128 (N_15128,N_8173,N_11726);
or U15129 (N_15129,N_11693,N_11376);
or U15130 (N_15130,N_8757,N_9856);
nand U15131 (N_15131,N_10294,N_8572);
or U15132 (N_15132,N_10615,N_10250);
or U15133 (N_15133,N_10697,N_8024);
nor U15134 (N_15134,N_9052,N_8656);
or U15135 (N_15135,N_10922,N_10415);
or U15136 (N_15136,N_9198,N_9884);
or U15137 (N_15137,N_9818,N_10193);
nand U15138 (N_15138,N_10161,N_9117);
and U15139 (N_15139,N_11039,N_9321);
or U15140 (N_15140,N_10233,N_11822);
nor U15141 (N_15141,N_9484,N_8596);
or U15142 (N_15142,N_8164,N_9951);
and U15143 (N_15143,N_9749,N_10664);
nand U15144 (N_15144,N_11326,N_10290);
and U15145 (N_15145,N_8394,N_8669);
nor U15146 (N_15146,N_9517,N_8856);
and U15147 (N_15147,N_8100,N_11811);
and U15148 (N_15148,N_8959,N_10510);
nor U15149 (N_15149,N_9106,N_9876);
or U15150 (N_15150,N_9105,N_8118);
xor U15151 (N_15151,N_9907,N_11010);
or U15152 (N_15152,N_8863,N_8723);
nand U15153 (N_15153,N_9384,N_11683);
or U15154 (N_15154,N_9598,N_8858);
nand U15155 (N_15155,N_10005,N_8972);
nor U15156 (N_15156,N_11920,N_10015);
and U15157 (N_15157,N_10520,N_8422);
nor U15158 (N_15158,N_10718,N_9677);
xor U15159 (N_15159,N_10098,N_8582);
or U15160 (N_15160,N_9043,N_10167);
nand U15161 (N_15161,N_9942,N_9115);
nand U15162 (N_15162,N_9053,N_8455);
and U15163 (N_15163,N_11227,N_10124);
nand U15164 (N_15164,N_11635,N_10051);
and U15165 (N_15165,N_10194,N_11357);
or U15166 (N_15166,N_11782,N_11082);
and U15167 (N_15167,N_11380,N_8254);
and U15168 (N_15168,N_9735,N_8509);
xor U15169 (N_15169,N_10372,N_8910);
xor U15170 (N_15170,N_9031,N_11083);
or U15171 (N_15171,N_11306,N_10213);
nor U15172 (N_15172,N_11067,N_10292);
nor U15173 (N_15173,N_8315,N_9756);
nand U15174 (N_15174,N_8412,N_11111);
xor U15175 (N_15175,N_11610,N_11462);
xnor U15176 (N_15176,N_8220,N_11196);
and U15177 (N_15177,N_9984,N_11094);
nor U15178 (N_15178,N_10806,N_10039);
nor U15179 (N_15179,N_10725,N_9001);
or U15180 (N_15180,N_10330,N_9947);
or U15181 (N_15181,N_11771,N_9359);
nand U15182 (N_15182,N_10480,N_11785);
or U15183 (N_15183,N_9923,N_10236);
nand U15184 (N_15184,N_8690,N_10748);
nand U15185 (N_15185,N_9061,N_9662);
nor U15186 (N_15186,N_11023,N_9416);
nand U15187 (N_15187,N_10096,N_8388);
or U15188 (N_15188,N_9842,N_9754);
and U15189 (N_15189,N_11468,N_11128);
and U15190 (N_15190,N_10793,N_9059);
and U15191 (N_15191,N_9403,N_9156);
and U15192 (N_15192,N_10920,N_11942);
nand U15193 (N_15193,N_11763,N_10600);
and U15194 (N_15194,N_10441,N_8293);
nor U15195 (N_15195,N_8130,N_9702);
and U15196 (N_15196,N_8768,N_8582);
nand U15197 (N_15197,N_9133,N_8742);
nor U15198 (N_15198,N_11457,N_10451);
nor U15199 (N_15199,N_11375,N_8676);
nor U15200 (N_15200,N_8207,N_10253);
xnor U15201 (N_15201,N_9315,N_10331);
nor U15202 (N_15202,N_8045,N_9351);
and U15203 (N_15203,N_10342,N_9336);
or U15204 (N_15204,N_11081,N_8191);
or U15205 (N_15205,N_8725,N_8900);
nor U15206 (N_15206,N_9421,N_9363);
or U15207 (N_15207,N_11646,N_10853);
and U15208 (N_15208,N_9172,N_10720);
or U15209 (N_15209,N_10903,N_9728);
xnor U15210 (N_15210,N_11631,N_10625);
and U15211 (N_15211,N_10367,N_8358);
nor U15212 (N_15212,N_9848,N_11337);
nand U15213 (N_15213,N_9957,N_9771);
or U15214 (N_15214,N_10547,N_9513);
nand U15215 (N_15215,N_8961,N_9913);
and U15216 (N_15216,N_8788,N_11387);
or U15217 (N_15217,N_9597,N_8739);
xor U15218 (N_15218,N_8618,N_8269);
and U15219 (N_15219,N_11768,N_8925);
or U15220 (N_15220,N_8163,N_8509);
nor U15221 (N_15221,N_11845,N_9339);
xor U15222 (N_15222,N_11076,N_8636);
or U15223 (N_15223,N_11180,N_9642);
nor U15224 (N_15224,N_10506,N_11631);
or U15225 (N_15225,N_9244,N_11611);
nor U15226 (N_15226,N_9451,N_11819);
nor U15227 (N_15227,N_8251,N_8806);
and U15228 (N_15228,N_9967,N_9171);
or U15229 (N_15229,N_8240,N_11310);
and U15230 (N_15230,N_9877,N_11497);
and U15231 (N_15231,N_8608,N_11979);
nor U15232 (N_15232,N_11946,N_11631);
nor U15233 (N_15233,N_10785,N_9128);
xor U15234 (N_15234,N_11291,N_10517);
and U15235 (N_15235,N_11518,N_11215);
xor U15236 (N_15236,N_9509,N_10176);
nand U15237 (N_15237,N_9838,N_9028);
or U15238 (N_15238,N_11700,N_10078);
nand U15239 (N_15239,N_11411,N_9090);
nor U15240 (N_15240,N_8594,N_8072);
or U15241 (N_15241,N_8575,N_9337);
or U15242 (N_15242,N_10080,N_11067);
nand U15243 (N_15243,N_10181,N_9382);
xnor U15244 (N_15244,N_8997,N_10411);
and U15245 (N_15245,N_8684,N_8445);
and U15246 (N_15246,N_9391,N_10339);
xnor U15247 (N_15247,N_11548,N_10892);
and U15248 (N_15248,N_11971,N_9171);
nand U15249 (N_15249,N_8931,N_11407);
or U15250 (N_15250,N_10384,N_9651);
nor U15251 (N_15251,N_8940,N_9807);
xor U15252 (N_15252,N_11353,N_8983);
nand U15253 (N_15253,N_9246,N_9996);
and U15254 (N_15254,N_10164,N_8632);
or U15255 (N_15255,N_9527,N_11455);
or U15256 (N_15256,N_10126,N_10164);
and U15257 (N_15257,N_10919,N_9283);
or U15258 (N_15258,N_9807,N_11663);
xor U15259 (N_15259,N_11950,N_9364);
nand U15260 (N_15260,N_10944,N_9273);
xnor U15261 (N_15261,N_11915,N_11299);
and U15262 (N_15262,N_11319,N_8562);
and U15263 (N_15263,N_10823,N_10568);
nor U15264 (N_15264,N_8141,N_10309);
nand U15265 (N_15265,N_9170,N_10967);
and U15266 (N_15266,N_10279,N_10606);
or U15267 (N_15267,N_11565,N_9472);
or U15268 (N_15268,N_11359,N_11019);
or U15269 (N_15269,N_8398,N_8288);
nor U15270 (N_15270,N_8303,N_11291);
or U15271 (N_15271,N_9962,N_9114);
or U15272 (N_15272,N_10974,N_11560);
and U15273 (N_15273,N_10694,N_11833);
and U15274 (N_15274,N_8957,N_10409);
nor U15275 (N_15275,N_11794,N_9665);
or U15276 (N_15276,N_8955,N_10387);
nand U15277 (N_15277,N_9916,N_11935);
nand U15278 (N_15278,N_8390,N_9805);
nand U15279 (N_15279,N_11372,N_11059);
nand U15280 (N_15280,N_9281,N_8694);
and U15281 (N_15281,N_11980,N_11750);
nand U15282 (N_15282,N_11643,N_8291);
and U15283 (N_15283,N_8779,N_8978);
nor U15284 (N_15284,N_11077,N_10213);
nor U15285 (N_15285,N_8222,N_9995);
or U15286 (N_15286,N_9228,N_10965);
or U15287 (N_15287,N_9401,N_9216);
or U15288 (N_15288,N_9087,N_8917);
nand U15289 (N_15289,N_8748,N_11519);
or U15290 (N_15290,N_11401,N_11352);
xor U15291 (N_15291,N_10895,N_8912);
nand U15292 (N_15292,N_11175,N_9308);
and U15293 (N_15293,N_9451,N_9797);
or U15294 (N_15294,N_11453,N_11336);
xor U15295 (N_15295,N_8412,N_8122);
or U15296 (N_15296,N_9028,N_11999);
nand U15297 (N_15297,N_9628,N_8690);
or U15298 (N_15298,N_10150,N_11474);
nand U15299 (N_15299,N_8590,N_10733);
or U15300 (N_15300,N_9633,N_8008);
nor U15301 (N_15301,N_10191,N_9285);
nand U15302 (N_15302,N_8159,N_8327);
xnor U15303 (N_15303,N_9031,N_9920);
nand U15304 (N_15304,N_10331,N_10487);
xnor U15305 (N_15305,N_9785,N_11530);
and U15306 (N_15306,N_9079,N_9146);
or U15307 (N_15307,N_8718,N_11716);
xnor U15308 (N_15308,N_10937,N_8311);
and U15309 (N_15309,N_10301,N_11224);
nor U15310 (N_15310,N_9876,N_10654);
nor U15311 (N_15311,N_8935,N_8097);
and U15312 (N_15312,N_11602,N_10862);
or U15313 (N_15313,N_8083,N_10011);
or U15314 (N_15314,N_10995,N_8806);
nand U15315 (N_15315,N_8969,N_8575);
nor U15316 (N_15316,N_9205,N_10560);
nor U15317 (N_15317,N_11116,N_9209);
nor U15318 (N_15318,N_9977,N_10906);
and U15319 (N_15319,N_9087,N_10864);
nor U15320 (N_15320,N_8434,N_11917);
or U15321 (N_15321,N_10779,N_11380);
nor U15322 (N_15322,N_10760,N_8372);
and U15323 (N_15323,N_11774,N_11138);
nand U15324 (N_15324,N_8157,N_9367);
and U15325 (N_15325,N_10536,N_8385);
or U15326 (N_15326,N_11533,N_11563);
nand U15327 (N_15327,N_9856,N_10043);
xor U15328 (N_15328,N_9413,N_9597);
nand U15329 (N_15329,N_9249,N_8678);
nor U15330 (N_15330,N_8526,N_10995);
nand U15331 (N_15331,N_11860,N_8807);
nand U15332 (N_15332,N_9437,N_11240);
nand U15333 (N_15333,N_10277,N_11744);
or U15334 (N_15334,N_10281,N_8396);
and U15335 (N_15335,N_9106,N_10868);
nand U15336 (N_15336,N_11043,N_10943);
or U15337 (N_15337,N_9636,N_8465);
nor U15338 (N_15338,N_8305,N_8463);
or U15339 (N_15339,N_9210,N_10179);
nand U15340 (N_15340,N_9283,N_11229);
nor U15341 (N_15341,N_11398,N_8456);
or U15342 (N_15342,N_11288,N_11804);
or U15343 (N_15343,N_10715,N_8293);
nor U15344 (N_15344,N_10304,N_8503);
nor U15345 (N_15345,N_11511,N_10910);
nor U15346 (N_15346,N_8984,N_11570);
xnor U15347 (N_15347,N_11549,N_11281);
nand U15348 (N_15348,N_8444,N_9538);
nor U15349 (N_15349,N_8589,N_9582);
or U15350 (N_15350,N_10530,N_10939);
nor U15351 (N_15351,N_11435,N_11656);
or U15352 (N_15352,N_9995,N_9743);
nand U15353 (N_15353,N_11386,N_9450);
xor U15354 (N_15354,N_9805,N_9487);
nand U15355 (N_15355,N_9816,N_9251);
nor U15356 (N_15356,N_8412,N_9297);
and U15357 (N_15357,N_11098,N_8312);
nand U15358 (N_15358,N_8410,N_10140);
or U15359 (N_15359,N_8803,N_9233);
and U15360 (N_15360,N_10139,N_11845);
or U15361 (N_15361,N_11754,N_11353);
nor U15362 (N_15362,N_9124,N_11152);
nand U15363 (N_15363,N_9986,N_10110);
nand U15364 (N_15364,N_8757,N_11311);
nand U15365 (N_15365,N_8483,N_8213);
nor U15366 (N_15366,N_10367,N_9797);
nand U15367 (N_15367,N_10206,N_10282);
nand U15368 (N_15368,N_10841,N_11290);
nand U15369 (N_15369,N_8230,N_9400);
nor U15370 (N_15370,N_11618,N_11215);
or U15371 (N_15371,N_9403,N_10648);
and U15372 (N_15372,N_11435,N_10915);
and U15373 (N_15373,N_11640,N_11565);
and U15374 (N_15374,N_11209,N_9048);
nor U15375 (N_15375,N_11278,N_11436);
and U15376 (N_15376,N_8368,N_10238);
and U15377 (N_15377,N_11987,N_8108);
nand U15378 (N_15378,N_10301,N_10934);
xnor U15379 (N_15379,N_9660,N_9059);
and U15380 (N_15380,N_8052,N_10155);
and U15381 (N_15381,N_9419,N_11730);
or U15382 (N_15382,N_8673,N_11582);
nor U15383 (N_15383,N_11754,N_11674);
or U15384 (N_15384,N_9095,N_11866);
nand U15385 (N_15385,N_11631,N_8740);
nand U15386 (N_15386,N_8349,N_8929);
nor U15387 (N_15387,N_8543,N_8929);
nand U15388 (N_15388,N_8729,N_10541);
nor U15389 (N_15389,N_9007,N_10038);
nor U15390 (N_15390,N_11567,N_8412);
nand U15391 (N_15391,N_10914,N_9219);
xor U15392 (N_15392,N_11505,N_9694);
nand U15393 (N_15393,N_11645,N_8663);
nand U15394 (N_15394,N_9518,N_10320);
and U15395 (N_15395,N_9325,N_8307);
nor U15396 (N_15396,N_9404,N_10443);
nor U15397 (N_15397,N_8279,N_9924);
nand U15398 (N_15398,N_11261,N_9938);
and U15399 (N_15399,N_9749,N_9822);
nand U15400 (N_15400,N_10696,N_8924);
and U15401 (N_15401,N_10000,N_10061);
nor U15402 (N_15402,N_10996,N_10976);
and U15403 (N_15403,N_10379,N_11566);
nand U15404 (N_15404,N_9619,N_11741);
or U15405 (N_15405,N_8023,N_11094);
or U15406 (N_15406,N_8676,N_9802);
and U15407 (N_15407,N_11033,N_8699);
or U15408 (N_15408,N_10234,N_9300);
nor U15409 (N_15409,N_11333,N_11502);
or U15410 (N_15410,N_8001,N_10682);
nor U15411 (N_15411,N_10281,N_11923);
and U15412 (N_15412,N_10105,N_8516);
or U15413 (N_15413,N_8434,N_8726);
nand U15414 (N_15414,N_9553,N_10209);
and U15415 (N_15415,N_8779,N_8955);
or U15416 (N_15416,N_10437,N_8807);
nand U15417 (N_15417,N_9305,N_11955);
or U15418 (N_15418,N_8888,N_8151);
nand U15419 (N_15419,N_9989,N_10649);
and U15420 (N_15420,N_8556,N_10767);
nand U15421 (N_15421,N_11928,N_9519);
and U15422 (N_15422,N_9882,N_8222);
nand U15423 (N_15423,N_9473,N_11528);
or U15424 (N_15424,N_11168,N_8343);
or U15425 (N_15425,N_11292,N_8575);
and U15426 (N_15426,N_9157,N_9271);
nor U15427 (N_15427,N_8998,N_8326);
nand U15428 (N_15428,N_11028,N_10681);
nand U15429 (N_15429,N_8802,N_11842);
nor U15430 (N_15430,N_10160,N_11619);
nor U15431 (N_15431,N_10526,N_9967);
nand U15432 (N_15432,N_11671,N_9946);
nor U15433 (N_15433,N_10943,N_9906);
nand U15434 (N_15434,N_10780,N_8889);
and U15435 (N_15435,N_10168,N_10540);
and U15436 (N_15436,N_10706,N_8237);
nand U15437 (N_15437,N_11359,N_8516);
or U15438 (N_15438,N_8033,N_10797);
nand U15439 (N_15439,N_8478,N_8907);
and U15440 (N_15440,N_10626,N_11824);
xnor U15441 (N_15441,N_11357,N_8905);
and U15442 (N_15442,N_8182,N_10378);
nand U15443 (N_15443,N_10297,N_10393);
or U15444 (N_15444,N_8337,N_9355);
nand U15445 (N_15445,N_11454,N_10013);
and U15446 (N_15446,N_9099,N_11648);
or U15447 (N_15447,N_11030,N_11531);
or U15448 (N_15448,N_11757,N_9601);
nor U15449 (N_15449,N_10058,N_10999);
nor U15450 (N_15450,N_9790,N_8571);
nor U15451 (N_15451,N_11923,N_8878);
nor U15452 (N_15452,N_10253,N_10609);
xor U15453 (N_15453,N_8921,N_8904);
nor U15454 (N_15454,N_10947,N_10321);
nor U15455 (N_15455,N_11095,N_9300);
nor U15456 (N_15456,N_9583,N_10089);
xor U15457 (N_15457,N_9917,N_8542);
and U15458 (N_15458,N_9109,N_11958);
nand U15459 (N_15459,N_9403,N_11803);
nor U15460 (N_15460,N_10084,N_8878);
and U15461 (N_15461,N_9554,N_10546);
or U15462 (N_15462,N_10567,N_11440);
nand U15463 (N_15463,N_8327,N_11145);
or U15464 (N_15464,N_8281,N_10785);
nor U15465 (N_15465,N_9747,N_8694);
nor U15466 (N_15466,N_10154,N_9870);
nor U15467 (N_15467,N_9227,N_9369);
nor U15468 (N_15468,N_8449,N_11119);
and U15469 (N_15469,N_8187,N_8129);
and U15470 (N_15470,N_8764,N_9102);
nor U15471 (N_15471,N_10283,N_8912);
xor U15472 (N_15472,N_9156,N_10814);
and U15473 (N_15473,N_11385,N_8527);
or U15474 (N_15474,N_9102,N_11562);
nand U15475 (N_15475,N_10898,N_11246);
or U15476 (N_15476,N_8910,N_11687);
nand U15477 (N_15477,N_9725,N_9219);
nand U15478 (N_15478,N_8955,N_11438);
or U15479 (N_15479,N_10969,N_10283);
and U15480 (N_15480,N_10091,N_9667);
and U15481 (N_15481,N_8534,N_11152);
xor U15482 (N_15482,N_8646,N_11767);
nor U15483 (N_15483,N_9008,N_11400);
nand U15484 (N_15484,N_11433,N_9283);
or U15485 (N_15485,N_10696,N_9491);
nor U15486 (N_15486,N_8400,N_8953);
nand U15487 (N_15487,N_11799,N_11341);
or U15488 (N_15488,N_10355,N_11106);
nand U15489 (N_15489,N_8848,N_9040);
and U15490 (N_15490,N_10842,N_10221);
nor U15491 (N_15491,N_9951,N_8006);
nor U15492 (N_15492,N_10919,N_11491);
and U15493 (N_15493,N_8080,N_9687);
or U15494 (N_15494,N_11311,N_11455);
or U15495 (N_15495,N_10941,N_11417);
and U15496 (N_15496,N_11393,N_10692);
or U15497 (N_15497,N_11144,N_8201);
xnor U15498 (N_15498,N_10561,N_9248);
or U15499 (N_15499,N_9187,N_9626);
nand U15500 (N_15500,N_10205,N_11296);
and U15501 (N_15501,N_8497,N_8813);
nand U15502 (N_15502,N_9077,N_10692);
and U15503 (N_15503,N_8272,N_10130);
nand U15504 (N_15504,N_8984,N_8271);
nor U15505 (N_15505,N_8405,N_10319);
xnor U15506 (N_15506,N_10624,N_8815);
xnor U15507 (N_15507,N_10186,N_10656);
or U15508 (N_15508,N_9324,N_9338);
nor U15509 (N_15509,N_11580,N_8158);
nand U15510 (N_15510,N_11177,N_10582);
nand U15511 (N_15511,N_9668,N_11642);
and U15512 (N_15512,N_8514,N_8200);
and U15513 (N_15513,N_10834,N_11079);
or U15514 (N_15514,N_10620,N_10642);
or U15515 (N_15515,N_11330,N_9835);
or U15516 (N_15516,N_10842,N_8465);
nand U15517 (N_15517,N_8445,N_10315);
nor U15518 (N_15518,N_10856,N_10987);
or U15519 (N_15519,N_11815,N_11204);
and U15520 (N_15520,N_11476,N_8043);
and U15521 (N_15521,N_10760,N_9886);
nand U15522 (N_15522,N_9583,N_11948);
and U15523 (N_15523,N_8976,N_11089);
nor U15524 (N_15524,N_10042,N_8625);
nor U15525 (N_15525,N_8544,N_11663);
and U15526 (N_15526,N_9098,N_11704);
or U15527 (N_15527,N_10932,N_9639);
and U15528 (N_15528,N_9429,N_9007);
or U15529 (N_15529,N_11162,N_9957);
and U15530 (N_15530,N_8181,N_8954);
or U15531 (N_15531,N_9472,N_10321);
nand U15532 (N_15532,N_11981,N_10475);
or U15533 (N_15533,N_10458,N_10265);
or U15534 (N_15534,N_11253,N_10942);
nand U15535 (N_15535,N_11075,N_11533);
nand U15536 (N_15536,N_11228,N_9458);
nand U15537 (N_15537,N_9961,N_9601);
nor U15538 (N_15538,N_8241,N_9361);
nand U15539 (N_15539,N_11412,N_10628);
or U15540 (N_15540,N_11649,N_9741);
or U15541 (N_15541,N_8344,N_10398);
and U15542 (N_15542,N_10846,N_9330);
or U15543 (N_15543,N_10624,N_9055);
nor U15544 (N_15544,N_11077,N_11474);
xnor U15545 (N_15545,N_10858,N_8372);
or U15546 (N_15546,N_8821,N_11426);
and U15547 (N_15547,N_8607,N_9745);
or U15548 (N_15548,N_11420,N_8876);
and U15549 (N_15549,N_8199,N_10237);
and U15550 (N_15550,N_8972,N_9832);
nand U15551 (N_15551,N_11979,N_8844);
or U15552 (N_15552,N_8427,N_10602);
nor U15553 (N_15553,N_10893,N_11301);
and U15554 (N_15554,N_11397,N_11846);
or U15555 (N_15555,N_8173,N_8821);
or U15556 (N_15556,N_9599,N_9778);
or U15557 (N_15557,N_11554,N_11735);
nand U15558 (N_15558,N_10293,N_10408);
and U15559 (N_15559,N_11948,N_8117);
xor U15560 (N_15560,N_10342,N_11955);
nor U15561 (N_15561,N_11904,N_11315);
xor U15562 (N_15562,N_8441,N_10050);
and U15563 (N_15563,N_9209,N_11233);
and U15564 (N_15564,N_8517,N_11373);
or U15565 (N_15565,N_10994,N_8749);
or U15566 (N_15566,N_8270,N_9325);
or U15567 (N_15567,N_11716,N_8708);
or U15568 (N_15568,N_10896,N_8902);
nor U15569 (N_15569,N_8250,N_8660);
and U15570 (N_15570,N_11754,N_11042);
nand U15571 (N_15571,N_10518,N_10963);
nand U15572 (N_15572,N_11275,N_8995);
or U15573 (N_15573,N_9678,N_8675);
xor U15574 (N_15574,N_11454,N_10914);
nor U15575 (N_15575,N_9023,N_11304);
and U15576 (N_15576,N_11877,N_11335);
nand U15577 (N_15577,N_10874,N_11648);
or U15578 (N_15578,N_9018,N_10252);
or U15579 (N_15579,N_10154,N_9493);
and U15580 (N_15580,N_10226,N_11915);
nand U15581 (N_15581,N_8598,N_8551);
nor U15582 (N_15582,N_8532,N_8483);
nor U15583 (N_15583,N_8232,N_8284);
nand U15584 (N_15584,N_8480,N_11815);
and U15585 (N_15585,N_11067,N_8215);
or U15586 (N_15586,N_10485,N_8521);
and U15587 (N_15587,N_9687,N_8254);
and U15588 (N_15588,N_11904,N_11894);
or U15589 (N_15589,N_9458,N_10061);
and U15590 (N_15590,N_11327,N_8806);
and U15591 (N_15591,N_11114,N_9895);
and U15592 (N_15592,N_9309,N_11696);
xor U15593 (N_15593,N_8371,N_9234);
xor U15594 (N_15594,N_10807,N_9906);
nand U15595 (N_15595,N_8060,N_11754);
and U15596 (N_15596,N_8265,N_10260);
and U15597 (N_15597,N_8390,N_9415);
xor U15598 (N_15598,N_8575,N_11990);
nor U15599 (N_15599,N_8212,N_9186);
or U15600 (N_15600,N_9698,N_10531);
or U15601 (N_15601,N_11029,N_8103);
nor U15602 (N_15602,N_10587,N_8584);
or U15603 (N_15603,N_11249,N_11316);
nor U15604 (N_15604,N_10816,N_10889);
and U15605 (N_15605,N_10700,N_8565);
and U15606 (N_15606,N_11770,N_10781);
or U15607 (N_15607,N_8401,N_10152);
nor U15608 (N_15608,N_11702,N_9255);
and U15609 (N_15609,N_10043,N_9186);
and U15610 (N_15610,N_10054,N_10019);
and U15611 (N_15611,N_11395,N_10954);
or U15612 (N_15612,N_11329,N_9106);
nand U15613 (N_15613,N_8519,N_10230);
nor U15614 (N_15614,N_11116,N_9194);
and U15615 (N_15615,N_9984,N_9047);
and U15616 (N_15616,N_11400,N_8157);
nor U15617 (N_15617,N_9598,N_9521);
nor U15618 (N_15618,N_10382,N_8784);
nand U15619 (N_15619,N_10585,N_10583);
nand U15620 (N_15620,N_8327,N_8071);
xnor U15621 (N_15621,N_10049,N_9604);
nor U15622 (N_15622,N_9220,N_8889);
xor U15623 (N_15623,N_8746,N_11003);
or U15624 (N_15624,N_11233,N_8941);
nor U15625 (N_15625,N_8316,N_9424);
nand U15626 (N_15626,N_9717,N_9939);
nand U15627 (N_15627,N_8492,N_10945);
nand U15628 (N_15628,N_10070,N_9609);
nor U15629 (N_15629,N_11837,N_10012);
nand U15630 (N_15630,N_10096,N_8945);
and U15631 (N_15631,N_11178,N_8506);
or U15632 (N_15632,N_10765,N_10899);
nand U15633 (N_15633,N_9771,N_10831);
nor U15634 (N_15634,N_9482,N_11730);
nand U15635 (N_15635,N_9594,N_11047);
nor U15636 (N_15636,N_8649,N_8449);
nand U15637 (N_15637,N_8439,N_8934);
xor U15638 (N_15638,N_11186,N_11624);
nand U15639 (N_15639,N_9693,N_11765);
and U15640 (N_15640,N_11798,N_10274);
nand U15641 (N_15641,N_8452,N_10833);
nand U15642 (N_15642,N_9432,N_9441);
xnor U15643 (N_15643,N_10246,N_9290);
and U15644 (N_15644,N_10383,N_9466);
or U15645 (N_15645,N_10192,N_11946);
and U15646 (N_15646,N_11738,N_9220);
and U15647 (N_15647,N_11888,N_10489);
or U15648 (N_15648,N_11557,N_11552);
and U15649 (N_15649,N_11312,N_9158);
and U15650 (N_15650,N_11525,N_9426);
and U15651 (N_15651,N_11327,N_8857);
or U15652 (N_15652,N_11946,N_8107);
nand U15653 (N_15653,N_11918,N_11379);
nor U15654 (N_15654,N_11713,N_9388);
nor U15655 (N_15655,N_11542,N_10361);
nor U15656 (N_15656,N_11676,N_11489);
and U15657 (N_15657,N_8668,N_10968);
and U15658 (N_15658,N_10003,N_8508);
and U15659 (N_15659,N_10985,N_8613);
nor U15660 (N_15660,N_10109,N_9775);
and U15661 (N_15661,N_10296,N_8957);
and U15662 (N_15662,N_10910,N_8541);
nor U15663 (N_15663,N_9016,N_9519);
nand U15664 (N_15664,N_10168,N_8934);
and U15665 (N_15665,N_9074,N_11276);
and U15666 (N_15666,N_11696,N_9979);
xnor U15667 (N_15667,N_9163,N_9520);
xor U15668 (N_15668,N_11258,N_8460);
xnor U15669 (N_15669,N_8382,N_10284);
xnor U15670 (N_15670,N_8008,N_11447);
nor U15671 (N_15671,N_9186,N_11178);
or U15672 (N_15672,N_9396,N_9673);
nand U15673 (N_15673,N_8136,N_11678);
and U15674 (N_15674,N_11296,N_9755);
and U15675 (N_15675,N_11210,N_8465);
xor U15676 (N_15676,N_9778,N_10815);
or U15677 (N_15677,N_9770,N_10438);
xnor U15678 (N_15678,N_10128,N_11598);
or U15679 (N_15679,N_10781,N_9973);
and U15680 (N_15680,N_11820,N_8265);
nand U15681 (N_15681,N_11720,N_10004);
or U15682 (N_15682,N_10236,N_9192);
nand U15683 (N_15683,N_11761,N_11968);
nand U15684 (N_15684,N_8949,N_8151);
or U15685 (N_15685,N_9019,N_11647);
and U15686 (N_15686,N_11574,N_9072);
xor U15687 (N_15687,N_11230,N_9078);
nand U15688 (N_15688,N_9671,N_9751);
or U15689 (N_15689,N_10662,N_8999);
nand U15690 (N_15690,N_9569,N_8282);
nand U15691 (N_15691,N_8906,N_10098);
nand U15692 (N_15692,N_9166,N_9760);
nand U15693 (N_15693,N_9423,N_10054);
xor U15694 (N_15694,N_11541,N_10247);
or U15695 (N_15695,N_10914,N_10947);
nor U15696 (N_15696,N_9437,N_8692);
and U15697 (N_15697,N_10136,N_11975);
xnor U15698 (N_15698,N_11417,N_8039);
or U15699 (N_15699,N_8469,N_9972);
and U15700 (N_15700,N_9097,N_11768);
and U15701 (N_15701,N_10658,N_8508);
nand U15702 (N_15702,N_9374,N_10933);
and U15703 (N_15703,N_9497,N_8476);
xnor U15704 (N_15704,N_10878,N_8277);
nand U15705 (N_15705,N_9527,N_10427);
or U15706 (N_15706,N_9065,N_9187);
nand U15707 (N_15707,N_9199,N_10759);
nor U15708 (N_15708,N_11393,N_11197);
nand U15709 (N_15709,N_8660,N_11749);
and U15710 (N_15710,N_11548,N_8603);
nand U15711 (N_15711,N_10205,N_9391);
and U15712 (N_15712,N_8030,N_10021);
nor U15713 (N_15713,N_9607,N_10759);
nand U15714 (N_15714,N_9454,N_10582);
nor U15715 (N_15715,N_10556,N_10633);
and U15716 (N_15716,N_11372,N_9419);
nor U15717 (N_15717,N_8246,N_10899);
or U15718 (N_15718,N_11442,N_11939);
nor U15719 (N_15719,N_9030,N_10701);
nand U15720 (N_15720,N_9689,N_9984);
and U15721 (N_15721,N_10136,N_11043);
nor U15722 (N_15722,N_8090,N_10615);
or U15723 (N_15723,N_8588,N_10577);
or U15724 (N_15724,N_8118,N_10331);
nor U15725 (N_15725,N_9023,N_11033);
or U15726 (N_15726,N_11456,N_9773);
nor U15727 (N_15727,N_8001,N_10380);
nor U15728 (N_15728,N_9804,N_11997);
and U15729 (N_15729,N_8821,N_8804);
and U15730 (N_15730,N_10742,N_10624);
xor U15731 (N_15731,N_8543,N_9694);
nand U15732 (N_15732,N_10529,N_10324);
nor U15733 (N_15733,N_10710,N_11365);
or U15734 (N_15734,N_8466,N_8781);
nor U15735 (N_15735,N_9988,N_11590);
nand U15736 (N_15736,N_11827,N_9842);
nand U15737 (N_15737,N_11689,N_8889);
or U15738 (N_15738,N_10892,N_8689);
nor U15739 (N_15739,N_11536,N_10325);
or U15740 (N_15740,N_9933,N_11920);
nand U15741 (N_15741,N_9043,N_11665);
or U15742 (N_15742,N_9415,N_11043);
or U15743 (N_15743,N_10593,N_10441);
nor U15744 (N_15744,N_10147,N_10648);
nand U15745 (N_15745,N_10833,N_8538);
and U15746 (N_15746,N_8963,N_9648);
nand U15747 (N_15747,N_8718,N_9893);
or U15748 (N_15748,N_8761,N_8714);
and U15749 (N_15749,N_9641,N_10029);
nand U15750 (N_15750,N_10153,N_10874);
or U15751 (N_15751,N_8103,N_8077);
or U15752 (N_15752,N_8686,N_11605);
or U15753 (N_15753,N_9293,N_11447);
xnor U15754 (N_15754,N_9266,N_11241);
or U15755 (N_15755,N_9511,N_9649);
and U15756 (N_15756,N_8571,N_8524);
nand U15757 (N_15757,N_10814,N_11839);
xnor U15758 (N_15758,N_10583,N_8623);
or U15759 (N_15759,N_11807,N_8233);
or U15760 (N_15760,N_11490,N_10103);
nor U15761 (N_15761,N_8657,N_9678);
nor U15762 (N_15762,N_8879,N_8792);
nand U15763 (N_15763,N_11570,N_11993);
and U15764 (N_15764,N_9771,N_9264);
nand U15765 (N_15765,N_10457,N_9934);
nor U15766 (N_15766,N_10085,N_9180);
nand U15767 (N_15767,N_10329,N_9599);
and U15768 (N_15768,N_10072,N_10911);
or U15769 (N_15769,N_9790,N_10451);
or U15770 (N_15770,N_8351,N_8244);
xor U15771 (N_15771,N_9989,N_10701);
nor U15772 (N_15772,N_9508,N_8611);
nor U15773 (N_15773,N_8744,N_9899);
nand U15774 (N_15774,N_10461,N_8246);
or U15775 (N_15775,N_8496,N_9226);
or U15776 (N_15776,N_10490,N_8431);
and U15777 (N_15777,N_8441,N_9132);
nor U15778 (N_15778,N_11837,N_11938);
and U15779 (N_15779,N_8734,N_8581);
nand U15780 (N_15780,N_8267,N_11219);
nand U15781 (N_15781,N_11942,N_9765);
nor U15782 (N_15782,N_11155,N_9801);
and U15783 (N_15783,N_10005,N_10194);
and U15784 (N_15784,N_8059,N_9270);
or U15785 (N_15785,N_8578,N_8625);
nor U15786 (N_15786,N_8137,N_11937);
or U15787 (N_15787,N_10794,N_9921);
nand U15788 (N_15788,N_11324,N_8534);
and U15789 (N_15789,N_9727,N_9377);
nor U15790 (N_15790,N_11208,N_8748);
nand U15791 (N_15791,N_9168,N_8061);
xor U15792 (N_15792,N_11036,N_10887);
xnor U15793 (N_15793,N_10454,N_11318);
xnor U15794 (N_15794,N_9125,N_11962);
nand U15795 (N_15795,N_8189,N_11296);
nand U15796 (N_15796,N_9834,N_9332);
or U15797 (N_15797,N_8516,N_8754);
or U15798 (N_15798,N_8442,N_11644);
nand U15799 (N_15799,N_8834,N_8586);
or U15800 (N_15800,N_10957,N_9959);
and U15801 (N_15801,N_8185,N_8499);
nor U15802 (N_15802,N_8259,N_8791);
and U15803 (N_15803,N_10533,N_8346);
nor U15804 (N_15804,N_10903,N_10187);
and U15805 (N_15805,N_9490,N_9942);
or U15806 (N_15806,N_10654,N_8966);
and U15807 (N_15807,N_11421,N_11808);
or U15808 (N_15808,N_8735,N_11757);
nand U15809 (N_15809,N_10170,N_11025);
and U15810 (N_15810,N_9237,N_11552);
nand U15811 (N_15811,N_8330,N_8936);
nand U15812 (N_15812,N_9931,N_9405);
and U15813 (N_15813,N_10465,N_9480);
nor U15814 (N_15814,N_10512,N_10272);
nor U15815 (N_15815,N_11934,N_11275);
nor U15816 (N_15816,N_9547,N_9431);
nor U15817 (N_15817,N_10920,N_9270);
nand U15818 (N_15818,N_8079,N_9592);
xnor U15819 (N_15819,N_10538,N_8105);
and U15820 (N_15820,N_11035,N_8595);
and U15821 (N_15821,N_9174,N_8662);
or U15822 (N_15822,N_11250,N_10415);
or U15823 (N_15823,N_11106,N_9340);
or U15824 (N_15824,N_8759,N_8929);
and U15825 (N_15825,N_9966,N_10822);
nor U15826 (N_15826,N_11775,N_8508);
nor U15827 (N_15827,N_9332,N_10300);
nand U15828 (N_15828,N_9482,N_11373);
or U15829 (N_15829,N_9091,N_11133);
nand U15830 (N_15830,N_9755,N_11791);
xor U15831 (N_15831,N_8425,N_8799);
nor U15832 (N_15832,N_8225,N_11605);
nand U15833 (N_15833,N_8316,N_10931);
or U15834 (N_15834,N_11371,N_10478);
and U15835 (N_15835,N_9310,N_10174);
and U15836 (N_15836,N_11968,N_10364);
nand U15837 (N_15837,N_10175,N_11543);
nor U15838 (N_15838,N_8083,N_10824);
and U15839 (N_15839,N_10831,N_10741);
xor U15840 (N_15840,N_8331,N_10644);
and U15841 (N_15841,N_9958,N_9133);
and U15842 (N_15842,N_9838,N_11246);
nand U15843 (N_15843,N_8372,N_11609);
nor U15844 (N_15844,N_9108,N_8243);
or U15845 (N_15845,N_9812,N_10365);
and U15846 (N_15846,N_10961,N_10190);
nor U15847 (N_15847,N_9006,N_8873);
or U15848 (N_15848,N_8298,N_8323);
nand U15849 (N_15849,N_11059,N_10143);
nand U15850 (N_15850,N_8142,N_8059);
or U15851 (N_15851,N_8725,N_9038);
nand U15852 (N_15852,N_10354,N_9057);
nor U15853 (N_15853,N_9230,N_11751);
or U15854 (N_15854,N_8628,N_11783);
nand U15855 (N_15855,N_8187,N_9669);
or U15856 (N_15856,N_9482,N_11438);
and U15857 (N_15857,N_9255,N_8411);
nand U15858 (N_15858,N_10462,N_10851);
and U15859 (N_15859,N_9016,N_9393);
nor U15860 (N_15860,N_10766,N_11327);
nand U15861 (N_15861,N_11158,N_9485);
and U15862 (N_15862,N_8026,N_9474);
and U15863 (N_15863,N_9568,N_10904);
nor U15864 (N_15864,N_9925,N_9023);
and U15865 (N_15865,N_9553,N_8946);
or U15866 (N_15866,N_10313,N_8203);
and U15867 (N_15867,N_9322,N_10854);
nand U15868 (N_15868,N_11874,N_8753);
nor U15869 (N_15869,N_10529,N_11378);
nor U15870 (N_15870,N_8190,N_8877);
xnor U15871 (N_15871,N_8636,N_8717);
or U15872 (N_15872,N_9737,N_8672);
nor U15873 (N_15873,N_11351,N_8591);
xor U15874 (N_15874,N_10788,N_11271);
nor U15875 (N_15875,N_10935,N_8553);
nand U15876 (N_15876,N_10513,N_10939);
nor U15877 (N_15877,N_9409,N_9437);
nor U15878 (N_15878,N_11443,N_9433);
and U15879 (N_15879,N_11270,N_8894);
nand U15880 (N_15880,N_11056,N_9741);
or U15881 (N_15881,N_8229,N_8502);
and U15882 (N_15882,N_9727,N_11384);
nor U15883 (N_15883,N_9768,N_10776);
or U15884 (N_15884,N_8167,N_8087);
xnor U15885 (N_15885,N_9192,N_11272);
nand U15886 (N_15886,N_9841,N_10051);
nand U15887 (N_15887,N_8875,N_8095);
or U15888 (N_15888,N_11768,N_8814);
or U15889 (N_15889,N_10263,N_10021);
or U15890 (N_15890,N_9693,N_11391);
nor U15891 (N_15891,N_10377,N_10886);
xnor U15892 (N_15892,N_8873,N_11736);
or U15893 (N_15893,N_10848,N_11433);
and U15894 (N_15894,N_9748,N_9866);
nand U15895 (N_15895,N_10611,N_10537);
nand U15896 (N_15896,N_8487,N_11295);
nor U15897 (N_15897,N_9989,N_10656);
and U15898 (N_15898,N_8184,N_10163);
or U15899 (N_15899,N_8623,N_8593);
or U15900 (N_15900,N_8758,N_11435);
or U15901 (N_15901,N_8359,N_8446);
nand U15902 (N_15902,N_11676,N_11040);
or U15903 (N_15903,N_8456,N_9507);
nor U15904 (N_15904,N_10919,N_11437);
nor U15905 (N_15905,N_9346,N_9855);
or U15906 (N_15906,N_10346,N_8228);
nor U15907 (N_15907,N_9165,N_8523);
nand U15908 (N_15908,N_10885,N_8290);
and U15909 (N_15909,N_9571,N_10228);
xor U15910 (N_15910,N_11215,N_9725);
and U15911 (N_15911,N_9794,N_8338);
nand U15912 (N_15912,N_9454,N_11737);
nor U15913 (N_15913,N_11987,N_11913);
nor U15914 (N_15914,N_10954,N_9060);
nand U15915 (N_15915,N_8807,N_11413);
or U15916 (N_15916,N_9492,N_9675);
or U15917 (N_15917,N_8766,N_8112);
nor U15918 (N_15918,N_10778,N_8189);
or U15919 (N_15919,N_11467,N_10760);
and U15920 (N_15920,N_9844,N_8693);
nor U15921 (N_15921,N_10759,N_9965);
nand U15922 (N_15922,N_8447,N_9741);
nand U15923 (N_15923,N_10169,N_8891);
or U15924 (N_15924,N_8538,N_9204);
and U15925 (N_15925,N_11686,N_11899);
xor U15926 (N_15926,N_11716,N_8228);
or U15927 (N_15927,N_11053,N_8112);
nor U15928 (N_15928,N_10918,N_11587);
or U15929 (N_15929,N_10501,N_10283);
nor U15930 (N_15930,N_9400,N_9567);
or U15931 (N_15931,N_9136,N_9028);
and U15932 (N_15932,N_10829,N_9637);
nand U15933 (N_15933,N_11197,N_10431);
nor U15934 (N_15934,N_11343,N_8965);
nor U15935 (N_15935,N_9830,N_9284);
or U15936 (N_15936,N_9950,N_11443);
and U15937 (N_15937,N_9199,N_11847);
xnor U15938 (N_15938,N_11097,N_11273);
nand U15939 (N_15939,N_10484,N_10389);
xor U15940 (N_15940,N_11768,N_8739);
and U15941 (N_15941,N_9369,N_10310);
and U15942 (N_15942,N_11822,N_9454);
nand U15943 (N_15943,N_8227,N_9395);
xor U15944 (N_15944,N_11457,N_10661);
and U15945 (N_15945,N_10001,N_8063);
and U15946 (N_15946,N_10844,N_8388);
or U15947 (N_15947,N_11964,N_10489);
xnor U15948 (N_15948,N_9740,N_9952);
or U15949 (N_15949,N_8716,N_9125);
nor U15950 (N_15950,N_11739,N_9481);
and U15951 (N_15951,N_10000,N_8524);
or U15952 (N_15952,N_9932,N_8831);
and U15953 (N_15953,N_10831,N_8467);
nand U15954 (N_15954,N_10622,N_10700);
nor U15955 (N_15955,N_9645,N_10227);
nor U15956 (N_15956,N_8119,N_8399);
nand U15957 (N_15957,N_11344,N_10821);
and U15958 (N_15958,N_9594,N_8694);
and U15959 (N_15959,N_10810,N_8335);
nor U15960 (N_15960,N_11462,N_11145);
nor U15961 (N_15961,N_9176,N_8507);
nor U15962 (N_15962,N_10474,N_8255);
and U15963 (N_15963,N_10660,N_10407);
and U15964 (N_15964,N_10084,N_9837);
nand U15965 (N_15965,N_8058,N_9050);
or U15966 (N_15966,N_11983,N_9854);
and U15967 (N_15967,N_11461,N_10571);
or U15968 (N_15968,N_8461,N_8978);
nor U15969 (N_15969,N_9566,N_11873);
nand U15970 (N_15970,N_10667,N_11532);
or U15971 (N_15971,N_10513,N_8035);
xnor U15972 (N_15972,N_8200,N_9091);
nor U15973 (N_15973,N_8044,N_9875);
nand U15974 (N_15974,N_10905,N_11671);
or U15975 (N_15975,N_8989,N_11215);
nor U15976 (N_15976,N_8074,N_9723);
and U15977 (N_15977,N_8975,N_9895);
nand U15978 (N_15978,N_9727,N_8504);
and U15979 (N_15979,N_11088,N_9803);
nor U15980 (N_15980,N_10352,N_11581);
nand U15981 (N_15981,N_10750,N_11784);
nor U15982 (N_15982,N_8587,N_11447);
or U15983 (N_15983,N_10577,N_8905);
or U15984 (N_15984,N_9373,N_8342);
or U15985 (N_15985,N_8917,N_11371);
nand U15986 (N_15986,N_11244,N_8131);
nor U15987 (N_15987,N_9646,N_9752);
nand U15988 (N_15988,N_11139,N_8790);
xnor U15989 (N_15989,N_11364,N_10291);
nand U15990 (N_15990,N_11178,N_8652);
nor U15991 (N_15991,N_11716,N_10542);
nand U15992 (N_15992,N_8799,N_10155);
nand U15993 (N_15993,N_8391,N_8469);
and U15994 (N_15994,N_10858,N_9115);
nand U15995 (N_15995,N_10636,N_10614);
or U15996 (N_15996,N_11161,N_8046);
and U15997 (N_15997,N_10091,N_8476);
or U15998 (N_15998,N_9436,N_8233);
nor U15999 (N_15999,N_11706,N_10189);
or U16000 (N_16000,N_15576,N_12472);
nor U16001 (N_16001,N_14405,N_12285);
nand U16002 (N_16002,N_12769,N_13991);
nand U16003 (N_16003,N_13579,N_13434);
xnor U16004 (N_16004,N_12501,N_15135);
and U16005 (N_16005,N_12827,N_13056);
nor U16006 (N_16006,N_14417,N_12594);
or U16007 (N_16007,N_13531,N_14304);
or U16008 (N_16008,N_14049,N_12502);
xor U16009 (N_16009,N_15674,N_13730);
or U16010 (N_16010,N_15333,N_13700);
and U16011 (N_16011,N_12199,N_14727);
nor U16012 (N_16012,N_15728,N_14174);
nand U16013 (N_16013,N_14345,N_13822);
and U16014 (N_16014,N_14792,N_12499);
xnor U16015 (N_16015,N_15398,N_15341);
nand U16016 (N_16016,N_12049,N_12336);
nor U16017 (N_16017,N_15336,N_14778);
or U16018 (N_16018,N_15298,N_12666);
or U16019 (N_16019,N_13975,N_12609);
xnor U16020 (N_16020,N_15979,N_15820);
and U16021 (N_16021,N_14670,N_13852);
or U16022 (N_16022,N_14609,N_14218);
and U16023 (N_16023,N_14807,N_14175);
and U16024 (N_16024,N_12069,N_12102);
nor U16025 (N_16025,N_14229,N_13359);
nor U16026 (N_16026,N_15683,N_15774);
or U16027 (N_16027,N_14921,N_13503);
and U16028 (N_16028,N_15896,N_12346);
or U16029 (N_16029,N_12053,N_15313);
or U16030 (N_16030,N_15953,N_13820);
or U16031 (N_16031,N_12129,N_14150);
xnor U16032 (N_16032,N_13270,N_13356);
nand U16033 (N_16033,N_14989,N_15575);
nand U16034 (N_16034,N_15003,N_15569);
or U16035 (N_16035,N_14893,N_12086);
nor U16036 (N_16036,N_14286,N_12838);
nor U16037 (N_16037,N_15046,N_15191);
xor U16038 (N_16038,N_15409,N_15723);
and U16039 (N_16039,N_13707,N_12717);
or U16040 (N_16040,N_14167,N_15706);
or U16041 (N_16041,N_15022,N_12245);
or U16042 (N_16042,N_12247,N_15417);
and U16043 (N_16043,N_12214,N_12698);
nor U16044 (N_16044,N_15442,N_13732);
or U16045 (N_16045,N_14940,N_14669);
nor U16046 (N_16046,N_13363,N_12396);
and U16047 (N_16047,N_14904,N_14388);
xnor U16048 (N_16048,N_15180,N_14080);
nor U16049 (N_16049,N_13818,N_14235);
xor U16050 (N_16050,N_14672,N_12019);
nand U16051 (N_16051,N_15759,N_13386);
or U16052 (N_16052,N_12018,N_13457);
and U16053 (N_16053,N_14973,N_14566);
nand U16054 (N_16054,N_13888,N_12063);
nor U16055 (N_16055,N_14008,N_13927);
or U16056 (N_16056,N_15045,N_15512);
nand U16057 (N_16057,N_13519,N_13087);
nand U16058 (N_16058,N_15929,N_15270);
nand U16059 (N_16059,N_13211,N_15996);
and U16060 (N_16060,N_14818,N_15105);
and U16061 (N_16061,N_15932,N_15631);
or U16062 (N_16062,N_14086,N_14574);
and U16063 (N_16063,N_12401,N_12050);
nand U16064 (N_16064,N_13950,N_14976);
and U16065 (N_16065,N_12082,N_13045);
or U16066 (N_16066,N_14564,N_15315);
nor U16067 (N_16067,N_12466,N_15424);
and U16068 (N_16068,N_12606,N_12337);
nand U16069 (N_16069,N_14529,N_13153);
xor U16070 (N_16070,N_15717,N_15472);
nor U16071 (N_16071,N_12378,N_14758);
and U16072 (N_16072,N_13227,N_13310);
or U16073 (N_16073,N_14024,N_12475);
nor U16074 (N_16074,N_14913,N_13920);
and U16075 (N_16075,N_12601,N_12469);
or U16076 (N_16076,N_12960,N_12851);
or U16077 (N_16077,N_12052,N_15700);
and U16078 (N_16078,N_14541,N_15858);
nor U16079 (N_16079,N_15921,N_13872);
and U16080 (N_16080,N_12309,N_14039);
or U16081 (N_16081,N_12222,N_14467);
and U16082 (N_16082,N_15773,N_15986);
xnor U16083 (N_16083,N_12560,N_14013);
nor U16084 (N_16084,N_14485,N_12414);
nor U16085 (N_16085,N_13664,N_15878);
nand U16086 (N_16086,N_14108,N_13005);
nand U16087 (N_16087,N_13725,N_15915);
and U16088 (N_16088,N_12744,N_15547);
xor U16089 (N_16089,N_13701,N_15006);
nand U16090 (N_16090,N_12459,N_15361);
nand U16091 (N_16091,N_12572,N_14078);
or U16092 (N_16092,N_14740,N_14223);
or U16093 (N_16093,N_12300,N_14867);
or U16094 (N_16094,N_13615,N_15276);
nor U16095 (N_16095,N_15543,N_15194);
and U16096 (N_16096,N_13084,N_14850);
xor U16097 (N_16097,N_14801,N_12238);
nor U16098 (N_16098,N_15934,N_12142);
xor U16099 (N_16099,N_15756,N_15474);
or U16100 (N_16100,N_13362,N_13151);
xnor U16101 (N_16101,N_13248,N_14996);
or U16102 (N_16102,N_12479,N_12356);
and U16103 (N_16103,N_13892,N_12143);
or U16104 (N_16104,N_15714,N_14949);
and U16105 (N_16105,N_12507,N_13574);
or U16106 (N_16106,N_14776,N_12638);
nor U16107 (N_16107,N_12713,N_15889);
nor U16108 (N_16108,N_14780,N_12435);
nor U16109 (N_16109,N_13952,N_14253);
or U16110 (N_16110,N_14052,N_14279);
or U16111 (N_16111,N_15779,N_15578);
or U16112 (N_16112,N_13719,N_12650);
xor U16113 (N_16113,N_13633,N_12637);
and U16114 (N_16114,N_12779,N_14927);
nor U16115 (N_16115,N_12492,N_15603);
or U16116 (N_16116,N_12514,N_15427);
or U16117 (N_16117,N_15084,N_12589);
and U16118 (N_16118,N_14946,N_14377);
and U16119 (N_16119,N_15102,N_13619);
or U16120 (N_16120,N_13302,N_13047);
and U16121 (N_16121,N_15615,N_12946);
xor U16122 (N_16122,N_12966,N_14370);
or U16123 (N_16123,N_13516,N_15583);
nand U16124 (N_16124,N_12442,N_12703);
nor U16125 (N_16125,N_14611,N_13346);
and U16126 (N_16126,N_13609,N_12944);
nor U16127 (N_16127,N_13777,N_13969);
and U16128 (N_16128,N_15869,N_14181);
or U16129 (N_16129,N_13058,N_13557);
nand U16130 (N_16130,N_12994,N_15726);
nor U16131 (N_16131,N_14518,N_12563);
nand U16132 (N_16132,N_14910,N_14042);
and U16133 (N_16133,N_15043,N_14667);
and U16134 (N_16134,N_12370,N_13951);
nand U16135 (N_16135,N_12029,N_15136);
nand U16136 (N_16136,N_13641,N_13051);
nor U16137 (N_16137,N_13342,N_15055);
xor U16138 (N_16138,N_15223,N_12316);
nand U16139 (N_16139,N_12242,N_12424);
nor U16140 (N_16140,N_14966,N_14885);
nand U16141 (N_16141,N_12977,N_15415);
nor U16142 (N_16142,N_14096,N_14010);
nand U16143 (N_16143,N_12799,N_12896);
nor U16144 (N_16144,N_13405,N_15019);
nand U16145 (N_16145,N_14040,N_12901);
nand U16146 (N_16146,N_15852,N_15179);
nand U16147 (N_16147,N_15231,N_12125);
or U16148 (N_16148,N_15499,N_13150);
and U16149 (N_16149,N_12193,N_12882);
nand U16150 (N_16150,N_15923,N_13745);
nor U16151 (N_16151,N_12458,N_15351);
nand U16152 (N_16152,N_12537,N_12067);
nor U16153 (N_16153,N_15160,N_13974);
or U16154 (N_16154,N_12229,N_14714);
or U16155 (N_16155,N_13761,N_15633);
xnor U16156 (N_16156,N_14214,N_15991);
or U16157 (N_16157,N_13008,N_15324);
xor U16158 (N_16158,N_13219,N_13322);
and U16159 (N_16159,N_12167,N_15225);
nor U16160 (N_16160,N_13953,N_14819);
and U16161 (N_16161,N_15173,N_12165);
nor U16162 (N_16162,N_14043,N_14307);
xnor U16163 (N_16163,N_15579,N_15804);
and U16164 (N_16164,N_12282,N_12998);
nand U16165 (N_16165,N_12813,N_13274);
and U16166 (N_16166,N_13088,N_12073);
or U16167 (N_16167,N_12766,N_13569);
and U16168 (N_16168,N_13788,N_15665);
or U16169 (N_16169,N_14948,N_14607);
xnor U16170 (N_16170,N_13597,N_15263);
xnor U16171 (N_16171,N_15154,N_13348);
nor U16172 (N_16172,N_15377,N_15766);
and U16173 (N_16173,N_14400,N_12568);
or U16174 (N_16174,N_14455,N_13325);
xor U16175 (N_16175,N_15822,N_14551);
or U16176 (N_16176,N_12433,N_14955);
nor U16177 (N_16177,N_12444,N_15807);
nand U16178 (N_16178,N_12982,N_13981);
nand U16179 (N_16179,N_12451,N_12513);
and U16180 (N_16180,N_12824,N_12719);
or U16181 (N_16181,N_14606,N_13210);
and U16182 (N_16182,N_12675,N_13759);
nor U16183 (N_16183,N_14757,N_14349);
nand U16184 (N_16184,N_14652,N_14384);
nand U16185 (N_16185,N_15604,N_12663);
and U16186 (N_16186,N_13517,N_12658);
or U16187 (N_16187,N_12000,N_12907);
nor U16188 (N_16188,N_15172,N_15972);
or U16189 (N_16189,N_14216,N_12128);
nand U16190 (N_16190,N_13285,N_13738);
and U16191 (N_16191,N_13768,N_14489);
and U16192 (N_16192,N_12906,N_14779);
or U16193 (N_16193,N_14933,N_15992);
or U16194 (N_16194,N_15634,N_14688);
and U16195 (N_16195,N_14673,N_15314);
or U16196 (N_16196,N_13033,N_12106);
xnor U16197 (N_16197,N_12196,N_14200);
xor U16198 (N_16198,N_15275,N_12494);
and U16199 (N_16199,N_14392,N_15190);
nand U16200 (N_16200,N_15110,N_15124);
or U16201 (N_16201,N_14368,N_14480);
nand U16202 (N_16202,N_14726,N_14593);
nor U16203 (N_16203,N_13241,N_15023);
and U16204 (N_16204,N_12613,N_14020);
nand U16205 (N_16205,N_13100,N_12967);
and U16206 (N_16206,N_14563,N_14891);
nor U16207 (N_16207,N_12175,N_15966);
and U16208 (N_16208,N_14502,N_14659);
and U16209 (N_16209,N_14746,N_13709);
nor U16210 (N_16210,N_13422,N_13407);
and U16211 (N_16211,N_13445,N_13965);
or U16212 (N_16212,N_14531,N_15647);
or U16213 (N_16213,N_15357,N_12884);
and U16214 (N_16214,N_15788,N_14944);
nor U16215 (N_16215,N_12376,N_15515);
nor U16216 (N_16216,N_15943,N_15380);
nor U16217 (N_16217,N_14750,N_14894);
and U16218 (N_16218,N_13804,N_13774);
or U16219 (N_16219,N_13547,N_15158);
nand U16220 (N_16220,N_13435,N_12312);
nand U16221 (N_16221,N_12344,N_12553);
and U16222 (N_16222,N_14087,N_15808);
xor U16223 (N_16223,N_12060,N_15217);
or U16224 (N_16224,N_15591,N_12530);
nor U16225 (N_16225,N_13402,N_15643);
xor U16226 (N_16226,N_14613,N_15289);
and U16227 (N_16227,N_12023,N_12954);
nand U16228 (N_16228,N_14333,N_13424);
nand U16229 (N_16229,N_14775,N_13308);
nand U16230 (N_16230,N_13311,N_13881);
nand U16231 (N_16231,N_13935,N_14097);
or U16232 (N_16232,N_12878,N_15493);
and U16233 (N_16233,N_13145,N_12375);
and U16234 (N_16234,N_13318,N_12622);
xnor U16235 (N_16235,N_13024,N_12176);
nor U16236 (N_16236,N_13332,N_14215);
or U16237 (N_16237,N_13490,N_13198);
nor U16238 (N_16238,N_14019,N_12207);
or U16239 (N_16239,N_12938,N_12042);
or U16240 (N_16240,N_12693,N_12620);
or U16241 (N_16241,N_14460,N_12263);
or U16242 (N_16242,N_15260,N_15396);
nor U16243 (N_16243,N_14748,N_12992);
or U16244 (N_16244,N_13875,N_15708);
or U16245 (N_16245,N_14856,N_15977);
and U16246 (N_16246,N_15024,N_14284);
nand U16247 (N_16247,N_14412,N_12130);
nor U16248 (N_16248,N_15900,N_15983);
or U16249 (N_16249,N_15737,N_12173);
or U16250 (N_16250,N_15407,N_13081);
or U16251 (N_16251,N_13521,N_15834);
nand U16252 (N_16252,N_12662,N_13723);
nand U16253 (N_16253,N_12251,N_14029);
nand U16254 (N_16254,N_13762,N_14387);
nor U16255 (N_16255,N_14883,N_14092);
or U16256 (N_16256,N_15588,N_14555);
xor U16257 (N_16257,N_12921,N_12699);
and U16258 (N_16258,N_14539,N_12372);
and U16259 (N_16259,N_15711,N_14126);
and U16260 (N_16260,N_12495,N_14676);
nand U16261 (N_16261,N_14114,N_15234);
nand U16262 (N_16262,N_13161,N_14419);
nor U16263 (N_16263,N_14472,N_13312);
nand U16264 (N_16264,N_15486,N_12075);
xor U16265 (N_16265,N_13658,N_13763);
nand U16266 (N_16266,N_12640,N_14596);
nor U16267 (N_16267,N_13358,N_13224);
nor U16268 (N_16268,N_15686,N_15743);
or U16269 (N_16269,N_15893,N_15233);
nand U16270 (N_16270,N_14974,N_13940);
or U16271 (N_16271,N_12116,N_13937);
xnor U16272 (N_16272,N_15961,N_15300);
nand U16273 (N_16273,N_14064,N_12743);
nand U16274 (N_16274,N_15599,N_13623);
nand U16275 (N_16275,N_15664,N_14381);
or U16276 (N_16276,N_12014,N_15497);
nor U16277 (N_16277,N_12162,N_12305);
nand U16278 (N_16278,N_15137,N_13685);
and U16279 (N_16279,N_12110,N_13070);
or U16280 (N_16280,N_12150,N_13233);
or U16281 (N_16281,N_13671,N_14000);
or U16282 (N_16282,N_13131,N_12817);
nand U16283 (N_16283,N_13186,N_15806);
nand U16284 (N_16284,N_13423,N_12091);
nor U16285 (N_16285,N_12085,N_13933);
xnor U16286 (N_16286,N_13269,N_15076);
or U16287 (N_16287,N_14487,N_13827);
and U16288 (N_16288,N_14737,N_15195);
nor U16289 (N_16289,N_14859,N_13982);
or U16290 (N_16290,N_13526,N_14295);
xor U16291 (N_16291,N_13113,N_14265);
and U16292 (N_16292,N_12135,N_15397);
nor U16293 (N_16293,N_15495,N_14890);
or U16294 (N_16294,N_12296,N_12178);
nor U16295 (N_16295,N_12152,N_14720);
and U16296 (N_16296,N_14407,N_14644);
and U16297 (N_16297,N_15177,N_12707);
xnor U16298 (N_16298,N_14511,N_13589);
and U16299 (N_16299,N_14700,N_12618);
nor U16300 (N_16300,N_14364,N_13463);
nor U16301 (N_16301,N_15060,N_14122);
and U16302 (N_16302,N_13060,N_13976);
nor U16303 (N_16303,N_13440,N_12677);
nor U16304 (N_16304,N_15635,N_15293);
and U16305 (N_16305,N_13347,N_15485);
nor U16306 (N_16306,N_14597,N_14712);
nor U16307 (N_16307,N_12752,N_15079);
and U16308 (N_16308,N_14236,N_12984);
or U16309 (N_16309,N_15391,N_15481);
or U16310 (N_16310,N_14881,N_13205);
or U16311 (N_16311,N_15386,N_13866);
and U16312 (N_16312,N_15720,N_14725);
nor U16313 (N_16313,N_14862,N_13978);
nor U16314 (N_16314,N_15856,N_14066);
and U16315 (N_16315,N_15555,N_12093);
or U16316 (N_16316,N_13271,N_12664);
nand U16317 (N_16317,N_13438,N_15245);
nand U16318 (N_16318,N_14865,N_14423);
or U16319 (N_16319,N_15450,N_15026);
nor U16320 (N_16320,N_15439,N_15688);
nor U16321 (N_16321,N_15404,N_15107);
nand U16322 (N_16322,N_12980,N_15265);
and U16323 (N_16323,N_13986,N_12936);
xor U16324 (N_16324,N_13054,N_14129);
or U16325 (N_16325,N_14468,N_15403);
and U16326 (N_16326,N_15238,N_14697);
xnor U16327 (N_16327,N_15216,N_14264);
or U16328 (N_16328,N_12169,N_12270);
nand U16329 (N_16329,N_12930,N_14664);
xnor U16330 (N_16330,N_13742,N_13166);
or U16331 (N_16331,N_15811,N_14627);
or U16332 (N_16332,N_14083,N_14575);
nand U16333 (N_16333,N_13061,N_15307);
nand U16334 (N_16334,N_12676,N_14646);
nor U16335 (N_16335,N_12841,N_14567);
nor U16336 (N_16336,N_13048,N_14988);
and U16337 (N_16337,N_14889,N_15385);
or U16338 (N_16338,N_13596,N_15328);
nand U16339 (N_16339,N_12345,N_12225);
or U16340 (N_16340,N_13637,N_13169);
nor U16341 (N_16341,N_13068,N_12145);
nor U16342 (N_16342,N_13416,N_15652);
nand U16343 (N_16343,N_12504,N_14391);
nand U16344 (N_16344,N_15566,N_12006);
xnor U16345 (N_16345,N_15843,N_15951);
nor U16346 (N_16346,N_13506,N_14523);
nand U16347 (N_16347,N_13839,N_12800);
nand U16348 (N_16348,N_12335,N_13335);
or U16349 (N_16349,N_15058,N_15798);
xor U16350 (N_16350,N_14866,N_13580);
and U16351 (N_16351,N_12999,N_14009);
nor U16352 (N_16352,N_14911,N_14586);
and U16353 (N_16353,N_12136,N_13731);
or U16354 (N_16354,N_15264,N_13512);
and U16355 (N_16355,N_13858,N_12518);
or U16356 (N_16356,N_15950,N_15701);
nor U16357 (N_16357,N_13317,N_13213);
nor U16358 (N_16358,N_13002,N_15317);
and U16359 (N_16359,N_15475,N_14619);
and U16360 (N_16360,N_14399,N_13484);
nor U16361 (N_16361,N_12593,N_14736);
or U16362 (N_16362,N_14558,N_13706);
or U16363 (N_16363,N_15152,N_13472);
nand U16364 (N_16364,N_15483,N_12619);
xnor U16365 (N_16365,N_12600,N_15099);
nand U16366 (N_16366,N_13543,N_15468);
and U16367 (N_16367,N_14482,N_14496);
nor U16368 (N_16368,N_12022,N_15732);
nor U16369 (N_16369,N_15917,N_15757);
and U16370 (N_16370,N_14657,N_13104);
nor U16371 (N_16371,N_14420,N_15623);
nand U16372 (N_16372,N_15242,N_12058);
xor U16373 (N_16373,N_14002,N_15203);
nor U16374 (N_16374,N_12416,N_14478);
nor U16375 (N_16375,N_14047,N_13411);
or U16376 (N_16376,N_12089,N_12555);
and U16377 (N_16377,N_12816,N_12291);
nand U16378 (N_16378,N_14084,N_13660);
nand U16379 (N_16379,N_14195,N_13697);
or U16380 (N_16380,N_13261,N_12721);
nand U16381 (N_16381,N_13963,N_13518);
or U16382 (N_16382,N_12531,N_15340);
and U16383 (N_16383,N_15198,N_13214);
or U16384 (N_16384,N_14051,N_13598);
nand U16385 (N_16385,N_14585,N_13663);
and U16386 (N_16386,N_12587,N_13582);
or U16387 (N_16387,N_14683,N_12301);
nand U16388 (N_16388,N_12055,N_13275);
nor U16389 (N_16389,N_13586,N_12661);
or U16390 (N_16390,N_15009,N_15622);
nor U16391 (N_16391,N_14484,N_15800);
nor U16392 (N_16392,N_12048,N_14924);
and U16393 (N_16393,N_14240,N_12852);
and U16394 (N_16394,N_14794,N_14569);
and U16395 (N_16395,N_15283,N_12184);
nand U16396 (N_16396,N_14838,N_14624);
nand U16397 (N_16397,N_13590,N_13456);
nand U16398 (N_16398,N_12182,N_13090);
or U16399 (N_16399,N_15814,N_15850);
nor U16400 (N_16400,N_14958,N_15736);
or U16401 (N_16401,N_12480,N_14825);
or U16402 (N_16402,N_14771,N_12750);
or U16403 (N_16403,N_13865,N_13454);
nand U16404 (N_16404,N_14612,N_13736);
nor U16405 (N_16405,N_14959,N_13606);
nand U16406 (N_16406,N_13230,N_14262);
or U16407 (N_16407,N_13505,N_13139);
nand U16408 (N_16408,N_12860,N_15860);
nand U16409 (N_16409,N_12298,N_15832);
nand U16410 (N_16410,N_14581,N_14063);
nand U16411 (N_16411,N_12651,N_13035);
nor U16412 (N_16412,N_13134,N_14906);
and U16413 (N_16413,N_13541,N_13357);
or U16414 (N_16414,N_13766,N_14273);
and U16415 (N_16415,N_13328,N_15657);
and U16416 (N_16416,N_14061,N_13137);
and U16417 (N_16417,N_12784,N_14728);
and U16418 (N_16418,N_13595,N_12987);
or U16419 (N_16419,N_15227,N_12447);
nor U16420 (N_16420,N_15362,N_13018);
nor U16421 (N_16421,N_15716,N_14239);
or U16422 (N_16422,N_14654,N_12158);
nand U16423 (N_16423,N_15861,N_13259);
and U16424 (N_16424,N_15488,N_13813);
and U16425 (N_16425,N_12007,N_13999);
nand U16426 (N_16426,N_14155,N_12484);
and U16427 (N_16427,N_15430,N_15738);
and U16428 (N_16428,N_12672,N_12163);
nor U16429 (N_16429,N_14414,N_12087);
nor U16430 (N_16430,N_14538,N_13130);
nand U16431 (N_16431,N_14133,N_14639);
nand U16432 (N_16432,N_13123,N_14565);
xor U16433 (N_16433,N_15709,N_13471);
or U16434 (N_16434,N_13752,N_15597);
and U16435 (N_16435,N_13349,N_12945);
nor U16436 (N_16436,N_14591,N_13148);
or U16437 (N_16437,N_15540,N_15329);
or U16438 (N_16438,N_13204,N_15589);
or U16439 (N_16439,N_13117,N_15687);
nand U16440 (N_16440,N_15596,N_12066);
nand U16441 (N_16441,N_15908,N_13909);
nand U16442 (N_16442,N_15343,N_14444);
nor U16443 (N_16443,N_15914,N_14269);
nand U16444 (N_16444,N_12154,N_13334);
nand U16445 (N_16445,N_15819,N_15465);
nand U16446 (N_16446,N_12684,N_15114);
xor U16447 (N_16447,N_14693,N_14431);
and U16448 (N_16448,N_13288,N_15368);
or U16449 (N_16449,N_12823,N_12126);
nand U16450 (N_16450,N_14733,N_12617);
nand U16451 (N_16451,N_14961,N_14608);
and U16452 (N_16452,N_14684,N_13942);
xnor U16453 (N_16453,N_15432,N_15150);
nor U16454 (N_16454,N_14202,N_14159);
and U16455 (N_16455,N_15031,N_15406);
and U16456 (N_16456,N_15985,N_14230);
nor U16457 (N_16457,N_12171,N_14124);
nand U16458 (N_16458,N_14787,N_14335);
or U16459 (N_16459,N_15502,N_12198);
nand U16460 (N_16460,N_14760,N_14777);
nor U16461 (N_16461,N_14062,N_13040);
or U16462 (N_16462,N_12139,N_15719);
nor U16463 (N_16463,N_14969,N_14984);
nand U16464 (N_16464,N_12105,N_12262);
and U16465 (N_16465,N_13877,N_15952);
nand U16466 (N_16466,N_14248,N_13878);
nand U16467 (N_16467,N_14360,N_12715);
and U16468 (N_16468,N_14982,N_13258);
or U16469 (N_16469,N_15744,N_13876);
xnor U16470 (N_16470,N_12566,N_12909);
or U16471 (N_16471,N_15678,N_15496);
or U16472 (N_16472,N_13437,N_15292);
xor U16473 (N_16473,N_15739,N_12935);
and U16474 (N_16474,N_12762,N_14620);
nor U16475 (N_16475,N_12728,N_13724);
nor U16476 (N_16476,N_12529,N_13716);
or U16477 (N_16477,N_12791,N_12685);
nor U16478 (N_16478,N_12054,N_14105);
xor U16479 (N_16479,N_13483,N_14418);
nor U16480 (N_16480,N_12765,N_12850);
nor U16481 (N_16481,N_15519,N_14774);
or U16482 (N_16482,N_15119,N_13996);
nor U16483 (N_16483,N_14542,N_14638);
nand U16484 (N_16484,N_15140,N_15214);
and U16485 (N_16485,N_15715,N_14300);
nand U16486 (N_16486,N_12760,N_14032);
nor U16487 (N_16487,N_13159,N_15106);
or U16488 (N_16488,N_14337,N_12079);
or U16489 (N_16489,N_13795,N_12233);
nor U16490 (N_16490,N_13020,N_12787);
nor U16491 (N_16491,N_12815,N_12814);
or U16492 (N_16492,N_14600,N_14823);
and U16493 (N_16493,N_12928,N_13196);
and U16494 (N_16494,N_12038,N_15890);
nand U16495 (N_16495,N_12315,N_13523);
nand U16496 (N_16496,N_12072,N_15973);
and U16497 (N_16497,N_12916,N_13031);
nand U16498 (N_16498,N_15164,N_12395);
nand U16499 (N_16499,N_14767,N_14630);
nor U16500 (N_16500,N_12697,N_14686);
and U16501 (N_16501,N_12485,N_13636);
nor U16502 (N_16502,N_13247,N_14182);
nor U16503 (N_16503,N_12598,N_15197);
nand U16504 (N_16504,N_12491,N_12151);
nor U16505 (N_16505,N_14427,N_14193);
nor U16506 (N_16506,N_15218,N_14705);
nand U16507 (N_16507,N_14028,N_12348);
xnor U16508 (N_16508,N_13617,N_14187);
or U16509 (N_16509,N_13502,N_15587);
nand U16510 (N_16510,N_13620,N_13215);
or U16511 (N_16511,N_13497,N_14835);
xor U16512 (N_16512,N_15322,N_14396);
and U16513 (N_16513,N_15848,N_13917);
and U16514 (N_16514,N_12460,N_12763);
and U16515 (N_16515,N_12796,N_14292);
and U16516 (N_16516,N_12463,N_12716);
nor U16517 (N_16517,N_15379,N_12218);
nor U16518 (N_16518,N_15091,N_14219);
nor U16519 (N_16519,N_13232,N_15538);
nand U16520 (N_16520,N_14470,N_14544);
nor U16521 (N_16521,N_15021,N_13811);
nor U16522 (N_16522,N_12856,N_12887);
and U16523 (N_16523,N_15503,N_15937);
nand U16524 (N_16524,N_14785,N_15121);
and U16525 (N_16525,N_14462,N_13065);
and U16526 (N_16526,N_13262,N_12867);
or U16527 (N_16527,N_12738,N_13593);
or U16528 (N_16528,N_13380,N_13944);
and U16529 (N_16529,N_12359,N_14527);
nand U16530 (N_16530,N_12639,N_13115);
xor U16531 (N_16531,N_12869,N_12596);
nor U16532 (N_16532,N_15211,N_12798);
xnor U16533 (N_16533,N_14473,N_12180);
or U16534 (N_16534,N_12673,N_15416);
nor U16535 (N_16535,N_13540,N_12532);
or U16536 (N_16536,N_15199,N_15767);
and U16537 (N_16537,N_14125,N_13879);
nor U16538 (N_16538,N_13231,N_13767);
and U16539 (N_16539,N_12794,N_14254);
nand U16540 (N_16540,N_14056,N_14509);
nand U16541 (N_16541,N_14185,N_13789);
or U16542 (N_16542,N_15826,N_15629);
nand U16543 (N_16543,N_15375,N_12610);
or U16544 (N_16544,N_13737,N_14553);
and U16545 (N_16545,N_13552,N_12217);
xnor U16546 (N_16546,N_12340,N_14724);
nand U16547 (N_16547,N_14492,N_13964);
nor U16548 (N_16548,N_14385,N_15096);
nand U16549 (N_16549,N_13443,N_12669);
nand U16550 (N_16550,N_14011,N_15243);
and U16551 (N_16551,N_13988,N_14072);
nand U16552 (N_16552,N_15374,N_13116);
and U16553 (N_16553,N_12240,N_13093);
nor U16554 (N_16554,N_13371,N_12837);
nand U16555 (N_16555,N_14098,N_12174);
nand U16556 (N_16556,N_15250,N_15466);
xnor U16557 (N_16557,N_12523,N_15193);
nand U16558 (N_16558,N_13441,N_14900);
nand U16559 (N_16559,N_15567,N_12381);
nand U16560 (N_16560,N_13947,N_13336);
nand U16561 (N_16561,N_12259,N_12428);
and U16562 (N_16562,N_13674,N_13149);
nand U16563 (N_16563,N_14449,N_12777);
or U16564 (N_16564,N_14351,N_14633);
nor U16565 (N_16565,N_13429,N_13538);
and U16566 (N_16566,N_13199,N_12213);
nor U16567 (N_16567,N_13741,N_12119);
and U16568 (N_16568,N_14177,N_13297);
nor U16569 (N_16569,N_14658,N_15443);
nor U16570 (N_16570,N_13010,N_13279);
and U16571 (N_16571,N_15241,N_12995);
and U16572 (N_16572,N_12864,N_14208);
nand U16573 (N_16573,N_13249,N_14037);
xnor U16574 (N_16574,N_12024,N_12283);
xor U16575 (N_16575,N_12803,N_15610);
and U16576 (N_16576,N_13042,N_12210);
and U16577 (N_16577,N_12855,N_14004);
nor U16578 (N_16578,N_13832,N_14112);
or U16579 (N_16579,N_13218,N_15421);
nor U16580 (N_16580,N_14871,N_15143);
xor U16581 (N_16581,N_15365,N_13603);
nor U16582 (N_16582,N_15461,N_15785);
or U16583 (N_16583,N_14799,N_14812);
nor U16584 (N_16584,N_14549,N_12755);
and U16585 (N_16585,N_14465,N_14160);
and U16586 (N_16586,N_12527,N_12915);
nor U16587 (N_16587,N_14451,N_15747);
and U16588 (N_16588,N_13473,N_14962);
and U16589 (N_16589,N_13077,N_14698);
xnor U16590 (N_16590,N_13803,N_12741);
nor U16591 (N_16591,N_13874,N_12043);
or U16592 (N_16592,N_15907,N_12940);
or U16593 (N_16593,N_14005,N_15489);
nor U16594 (N_16594,N_13368,N_12266);
nand U16595 (N_16595,N_14831,N_13583);
nor U16596 (N_16596,N_13182,N_12605);
or U16597 (N_16597,N_15065,N_12123);
nand U16598 (N_16598,N_13726,N_12274);
nand U16599 (N_16599,N_13188,N_14144);
nand U16600 (N_16600,N_14901,N_13770);
nand U16601 (N_16601,N_14934,N_15240);
and U16602 (N_16602,N_14796,N_15239);
nand U16603 (N_16603,N_15413,N_12403);
nor U16604 (N_16604,N_12013,N_12700);
nand U16605 (N_16605,N_15220,N_14164);
nand U16606 (N_16606,N_13539,N_12608);
or U16607 (N_16607,N_13102,N_12387);
and U16608 (N_16608,N_14715,N_13556);
or U16609 (N_16609,N_13053,N_12399);
and U16610 (N_16610,N_15772,N_12026);
nor U16611 (N_16611,N_12581,N_14583);
xnor U16612 (N_16612,N_13025,N_14355);
nor U16613 (N_16613,N_14907,N_13785);
or U16614 (N_16614,N_12657,N_13945);
nor U16615 (N_16615,N_14204,N_14655);
and U16616 (N_16616,N_13256,N_15894);
nand U16617 (N_16617,N_14251,N_15684);
nor U16618 (N_16618,N_13345,N_12419);
and U16619 (N_16619,N_15011,N_15444);
nor U16620 (N_16620,N_15038,N_12725);
nand U16621 (N_16621,N_13432,N_15845);
nor U16622 (N_16622,N_15866,N_15188);
or U16623 (N_16623,N_13147,N_15844);
and U16624 (N_16624,N_15614,N_14640);
nand U16625 (N_16625,N_14532,N_15369);
and U16626 (N_16626,N_14788,N_14389);
xnor U16627 (N_16627,N_14571,N_14975);
xor U16628 (N_16628,N_14457,N_13192);
xnor U16629 (N_16629,N_15000,N_12505);
and U16630 (N_16630,N_13189,N_15696);
xor U16631 (N_16631,N_12642,N_12612);
and U16632 (N_16632,N_15904,N_12411);
nand U16633 (N_16633,N_14915,N_12584);
xnor U16634 (N_16634,N_15414,N_12234);
or U16635 (N_16635,N_14828,N_15482);
nand U16636 (N_16636,N_15734,N_12561);
nand U16637 (N_16637,N_14888,N_12759);
nor U16638 (N_16638,N_14995,N_13775);
or U16639 (N_16639,N_15897,N_12100);
nor U16640 (N_16640,N_15261,N_14846);
or U16641 (N_16641,N_13234,N_14860);
or U16642 (N_16642,N_12432,N_12510);
nor U16643 (N_16643,N_14817,N_13943);
nand U16644 (N_16644,N_13848,N_15068);
nor U16645 (N_16645,N_12363,N_15760);
nand U16646 (N_16646,N_12037,N_15436);
or U16647 (N_16647,N_13870,N_15557);
nor U16648 (N_16648,N_15580,N_14461);
or U16649 (N_16649,N_15144,N_15942);
nor U16650 (N_16650,N_12865,N_13733);
nor U16651 (N_16651,N_14067,N_15693);
xor U16652 (N_16652,N_12201,N_15722);
nor U16653 (N_16653,N_12334,N_13050);
nor U16654 (N_16654,N_13379,N_12807);
and U16655 (N_16655,N_14853,N_15507);
xnor U16656 (N_16656,N_14815,N_14790);
and U16657 (N_16657,N_15252,N_15093);
nand U16658 (N_16658,N_14168,N_15842);
nand U16659 (N_16659,N_14170,N_15247);
nand U16660 (N_16660,N_13455,N_12107);
and U16661 (N_16661,N_15857,N_14699);
and U16662 (N_16662,N_14302,N_15458);
nand U16663 (N_16663,N_14272,N_14301);
and U16664 (N_16664,N_12261,N_12467);
or U16665 (N_16665,N_14212,N_13520);
nand U16666 (N_16666,N_13885,N_12338);
nor U16667 (N_16667,N_13853,N_14756);
nor U16668 (N_16668,N_13849,N_13178);
nand U16669 (N_16669,N_14617,N_12875);
xnor U16670 (N_16670,N_13754,N_12267);
nor U16671 (N_16671,N_12295,N_14550);
nor U16672 (N_16672,N_12981,N_14491);
nand U16673 (N_16673,N_13389,N_14142);
or U16674 (N_16674,N_12390,N_15690);
nor U16675 (N_16675,N_13904,N_12034);
or U16676 (N_16676,N_13837,N_14991);
nand U16677 (N_16677,N_15139,N_13897);
nand U16678 (N_16678,N_14833,N_13929);
nor U16679 (N_16679,N_13801,N_14971);
xor U16680 (N_16680,N_12062,N_14861);
or U16681 (N_16681,N_12811,N_12758);
or U16682 (N_16682,N_12051,N_12454);
xnor U16683 (N_16683,N_14556,N_14401);
nand U16684 (N_16684,N_13340,N_12567);
nand U16685 (N_16685,N_13649,N_13283);
nand U16686 (N_16686,N_13889,N_13015);
xnor U16687 (N_16687,N_15667,N_15879);
or U16688 (N_16688,N_12192,N_14937);
nor U16689 (N_16689,N_12496,N_12456);
nand U16690 (N_16690,N_14576,N_12326);
xnor U16691 (N_16691,N_15087,N_12586);
or U16692 (N_16692,N_14786,N_15565);
nor U16693 (N_16693,N_14605,N_13983);
nor U16694 (N_16694,N_15697,N_15441);
and U16695 (N_16695,N_14763,N_14822);
nand U16696 (N_16696,N_12871,N_12493);
nand U16697 (N_16697,N_13686,N_12287);
and U16698 (N_16698,N_14708,N_12094);
xor U16699 (N_16699,N_14386,N_15200);
or U16700 (N_16700,N_12969,N_12439);
nor U16701 (N_16701,N_14501,N_15425);
and U16702 (N_16702,N_14843,N_12101);
or U16703 (N_16703,N_14089,N_15978);
and U16704 (N_16704,N_12515,N_13462);
and U16705 (N_16705,N_12170,N_13417);
nor U16706 (N_16706,N_12032,N_14326);
or U16707 (N_16707,N_14653,N_15312);
and U16708 (N_16708,N_15204,N_12078);
nand U16709 (N_16709,N_15163,N_14075);
nand U16710 (N_16710,N_12912,N_13998);
and U16711 (N_16711,N_13220,N_13442);
or U16712 (N_16712,N_12888,N_14956);
xnor U16713 (N_16713,N_12547,N_14325);
nor U16714 (N_16714,N_12932,N_15922);
or U16715 (N_16715,N_14434,N_15269);
nand U16716 (N_16716,N_14402,N_14148);
nand U16717 (N_16717,N_12288,N_14849);
xnor U16718 (N_16718,N_12616,N_15660);
nor U16719 (N_16719,N_15492,N_14314);
and U16720 (N_16720,N_14506,N_15162);
or U16721 (N_16721,N_13669,N_15630);
or U16722 (N_16722,N_12179,N_15794);
nor U16723 (N_16723,N_15699,N_12249);
and U16724 (N_16724,N_13680,N_15980);
or U16725 (N_16725,N_13522,N_15434);
nand U16726 (N_16726,N_12629,N_12453);
and U16727 (N_16727,N_13152,N_15888);
and U16728 (N_16728,N_14674,N_15749);
or U16729 (N_16729,N_13304,N_13038);
xnor U16730 (N_16730,N_13451,N_12534);
and U16731 (N_16731,N_15902,N_15067);
nand U16732 (N_16732,N_14366,N_13562);
nand U16733 (N_16733,N_15183,N_13654);
or U16734 (N_16734,N_14497,N_14732);
nand U16735 (N_16735,N_15146,N_15178);
nand U16736 (N_16736,N_14811,N_12397);
nor U16737 (N_16737,N_14093,N_13403);
nand U16738 (N_16738,N_14217,N_13922);
nand U16739 (N_16739,N_15207,N_12825);
and U16740 (N_16740,N_12955,N_15624);
or U16741 (N_16741,N_13532,N_15764);
or U16742 (N_16742,N_12748,N_14250);
nand U16743 (N_16743,N_12056,N_13600);
nand U16744 (N_16744,N_12273,N_13242);
nand U16745 (N_16745,N_14963,N_13968);
nand U16746 (N_16746,N_12761,N_15334);
nand U16747 (N_16747,N_14027,N_14258);
and U16748 (N_16748,N_12470,N_14731);
and U16749 (N_16749,N_15827,N_14433);
or U16750 (N_16750,N_15816,N_12859);
nand U16751 (N_16751,N_15556,N_13846);
nand U16752 (N_16752,N_12324,N_15304);
xor U16753 (N_16753,N_12446,N_13385);
and U16754 (N_16754,N_15906,N_12783);
or U16755 (N_16755,N_13175,N_13027);
or U16756 (N_16756,N_15835,N_13162);
and U16757 (N_16757,N_15456,N_12556);
xor U16758 (N_16758,N_13781,N_12636);
or U16759 (N_16759,N_15305,N_13281);
nand U16760 (N_16760,N_14440,N_13133);
or U16761 (N_16761,N_14045,N_12092);
xnor U16762 (N_16762,N_15617,N_12889);
nand U16763 (N_16763,N_14115,N_15872);
nor U16764 (N_16764,N_12509,N_15303);
nor U16765 (N_16765,N_12625,N_13703);
and U16766 (N_16766,N_14415,N_13108);
xor U16767 (N_16767,N_13936,N_14450);
and U16768 (N_16768,N_12172,N_12362);
and U16769 (N_16769,N_14839,N_13343);
and U16770 (N_16770,N_15671,N_13729);
nor U16771 (N_16771,N_12828,N_14094);
or U16772 (N_16772,N_13821,N_14662);
and U16773 (N_16773,N_12917,N_12353);
nand U16774 (N_16774,N_14044,N_12329);
nor U16775 (N_16775,N_14874,N_12571);
or U16776 (N_16776,N_13467,N_15859);
nand U16777 (N_16777,N_14334,N_14987);
and U16778 (N_16778,N_12028,N_14663);
or U16779 (N_16779,N_13604,N_15875);
nor U16780 (N_16780,N_15731,N_15539);
nor U16781 (N_16781,N_12468,N_15372);
nor U16782 (N_16782,N_15125,N_14394);
nand U16783 (N_16783,N_15874,N_14347);
or U16784 (N_16784,N_13525,N_15054);
or U16785 (N_16785,N_15222,N_14764);
or U16786 (N_16786,N_12756,N_13533);
nor U16787 (N_16787,N_15337,N_14886);
nor U16788 (N_16788,N_13787,N_15967);
xor U16789 (N_16789,N_12227,N_12792);
and U16790 (N_16790,N_14425,N_15073);
nor U16791 (N_16791,N_15851,N_15524);
or U16792 (N_16792,N_13459,N_15355);
and U16793 (N_16793,N_15257,N_12208);
or U16794 (N_16794,N_13221,N_13399);
and U16795 (N_16795,N_15015,N_12255);
or U16796 (N_16796,N_14079,N_14338);
or U16797 (N_16797,N_13255,N_13694);
or U16798 (N_16798,N_14410,N_14055);
or U16799 (N_16799,N_13656,N_14559);
or U16800 (N_16800,N_13643,N_14299);
nand U16801 (N_16801,N_15039,N_15763);
nand U16802 (N_16802,N_15658,N_15670);
or U16803 (N_16803,N_14997,N_13509);
nor U16804 (N_16804,N_14783,N_15750);
or U16805 (N_16805,N_15048,N_13049);
nor U16806 (N_16806,N_12157,N_13911);
or U16807 (N_16807,N_12557,N_13174);
or U16808 (N_16808,N_12415,N_14521);
nand U16809 (N_16809,N_13683,N_14577);
nor U16810 (N_16810,N_12010,N_14820);
and U16811 (N_16811,N_12720,N_12420);
nor U16812 (N_16812,N_13806,N_14119);
and U16813 (N_16813,N_12754,N_14206);
nand U16814 (N_16814,N_12314,N_14131);
or U16815 (N_16815,N_12706,N_15871);
nand U16816 (N_16816,N_12108,N_13425);
nand U16817 (N_16817,N_12235,N_13681);
nand U16818 (N_16818,N_14376,N_14829);
nand U16819 (N_16819,N_14046,N_13382);
and U16820 (N_16820,N_15882,N_15438);
and U16821 (N_16821,N_14713,N_15830);
and U16822 (N_16822,N_15209,N_12194);
and U16823 (N_16823,N_15014,N_14939);
or U16824 (N_16824,N_15010,N_14117);
nand U16825 (N_16825,N_15095,N_12244);
nand U16826 (N_16826,N_15212,N_13946);
xnor U16827 (N_16827,N_15751,N_14162);
or U16828 (N_16828,N_12785,N_14595);
nand U16829 (N_16829,N_15956,N_14499);
xnor U16830 (N_16830,N_12205,N_15778);
nand U16831 (N_16831,N_14348,N_14471);
nand U16832 (N_16832,N_14721,N_12307);
nand U16833 (N_16833,N_15447,N_12628);
or U16834 (N_16834,N_15457,N_12243);
xor U16835 (N_16835,N_13023,N_12965);
and U16836 (N_16836,N_13043,N_13817);
nor U16837 (N_16837,N_15650,N_13272);
and U16838 (N_16838,N_13714,N_13823);
nor U16839 (N_16839,N_15668,N_15755);
and U16840 (N_16840,N_13962,N_13309);
and U16841 (N_16841,N_12789,N_13784);
or U16842 (N_16842,N_15295,N_15358);
nor U16843 (N_16843,N_15862,N_14318);
nor U16844 (N_16844,N_13501,N_12734);
nor U16845 (N_16845,N_14165,N_14429);
and U16846 (N_16846,N_12241,N_13327);
nand U16847 (N_16847,N_12718,N_13844);
or U16848 (N_16848,N_14139,N_12774);
nor U16849 (N_16849,N_15128,N_14287);
xor U16850 (N_16850,N_12310,N_13124);
and U16851 (N_16851,N_13941,N_14130);
nand U16852 (N_16852,N_15987,N_14935);
or U16853 (N_16853,N_13101,N_13780);
nor U16854 (N_16854,N_13277,N_15044);
or U16855 (N_16855,N_13118,N_15625);
nor U16856 (N_16856,N_12690,N_14312);
or U16857 (N_16857,N_13480,N_15100);
or U16858 (N_16858,N_13355,N_13461);
nor U16859 (N_16859,N_13374,N_14718);
xor U16860 (N_16860,N_15402,N_13800);
and U16861 (N_16861,N_15968,N_14015);
xor U16862 (N_16862,N_12747,N_12772);
nor U16863 (N_16863,N_13544,N_14908);
nand U16864 (N_16864,N_12570,N_15616);
and U16865 (N_16865,N_12035,N_13086);
and U16866 (N_16866,N_13326,N_14977);
or U16867 (N_16867,N_12412,N_12948);
nor U16868 (N_16868,N_12972,N_15226);
or U16869 (N_16869,N_12371,N_13548);
nor U16870 (N_16870,N_13551,N_13535);
nand U16871 (N_16871,N_14257,N_13850);
and U16872 (N_16872,N_15659,N_15388);
nor U16873 (N_16873,N_13657,N_14437);
nand U16874 (N_16874,N_12839,N_15661);
or U16875 (N_16875,N_15564,N_14844);
or U16876 (N_16876,N_12452,N_13067);
nand U16877 (N_16877,N_14928,N_13628);
nand U16878 (N_16878,N_12449,N_15762);
or U16879 (N_16879,N_12894,N_12924);
nor U16880 (N_16880,N_12751,N_15272);
nor U16881 (N_16881,N_15870,N_12365);
or U16882 (N_16882,N_14350,N_13482);
and U16883 (N_16883,N_12327,N_14526);
nand U16884 (N_16884,N_14957,N_12036);
nand U16885 (N_16885,N_14610,N_15306);
nand U16886 (N_16886,N_14876,N_12297);
xor U16887 (N_16887,N_15873,N_14719);
nor U16888 (N_16888,N_14628,N_12521);
or U16889 (N_16889,N_12979,N_12095);
or U16890 (N_16890,N_12558,N_15998);
or U16891 (N_16891,N_14268,N_13805);
and U16892 (N_16892,N_14845,N_12588);
xor U16893 (N_16893,N_14036,N_15679);
nor U16894 (N_16894,N_12786,N_15013);
nand U16895 (N_16895,N_15363,N_14903);
or U16896 (N_16896,N_15847,N_15215);
nor U16897 (N_16897,N_12425,N_14224);
nor U16898 (N_16898,N_15501,N_13354);
xor U16899 (N_16899,N_13601,N_14916);
or U16900 (N_16900,N_13105,N_14321);
nand U16901 (N_16901,N_12764,N_15171);
and U16902 (N_16902,N_14281,N_14001);
nand U16903 (N_16903,N_13171,N_14466);
nor U16904 (N_16904,N_13553,N_15536);
or U16905 (N_16905,N_15518,N_14766);
nand U16906 (N_16906,N_12726,N_13244);
nor U16907 (N_16907,N_12525,N_15941);
nor U16908 (N_16908,N_12868,N_14276);
xor U16909 (N_16909,N_14280,N_13698);
and U16910 (N_16910,N_13388,N_14864);
and U16911 (N_16911,N_15092,N_15418);
and U16912 (N_16912,N_13479,N_15611);
or U16913 (N_16913,N_15149,N_13602);
and U16914 (N_16914,N_12166,N_13786);
or U16915 (N_16915,N_15741,N_15718);
nor U16916 (N_16916,N_15562,N_14759);
or U16917 (N_16917,N_12576,N_14329);
nand U16918 (N_16918,N_12191,N_13995);
nand U16919 (N_16919,N_14873,N_12614);
and U16920 (N_16920,N_14369,N_15071);
nand U16921 (N_16921,N_14941,N_15948);
nor U16922 (N_16922,N_12668,N_12988);
nand U16923 (N_16923,N_14323,N_14649);
nor U16924 (N_16924,N_13282,N_13675);
or U16925 (N_16925,N_13939,N_13465);
nand U16926 (N_16926,N_15568,N_14762);
nand U16927 (N_16927,N_12302,N_12843);
nor U16928 (N_16928,N_12264,N_12899);
and U16929 (N_16929,N_15053,N_12870);
or U16930 (N_16930,N_15410,N_13647);
or U16931 (N_16931,N_15419,N_13702);
nor U16932 (N_16932,N_15408,N_15669);
xnor U16933 (N_16933,N_15098,N_12797);
nand U16934 (N_16934,N_12692,N_13111);
or U16935 (N_16935,N_15428,N_12925);
nor U16936 (N_16936,N_15422,N_12384);
nor U16937 (N_16937,N_12729,N_14026);
xnor U16938 (N_16938,N_14424,N_13573);
or U16939 (N_16939,N_12648,N_12404);
or U16940 (N_16940,N_13421,N_15885);
and U16941 (N_16941,N_12339,N_12232);
nand U16942 (N_16942,N_12161,N_12188);
nand U16943 (N_16943,N_12423,N_12578);
nand U16944 (N_16944,N_12025,N_15927);
and U16945 (N_16945,N_15691,N_12290);
and U16946 (N_16946,N_14246,N_14702);
or U16947 (N_16947,N_14735,N_14464);
or U16948 (N_16948,N_15648,N_15533);
xor U16949 (N_16949,N_15449,N_14517);
or U16950 (N_16950,N_12632,N_12074);
nor U16951 (N_16951,N_12795,N_14189);
nor U16952 (N_16952,N_12308,N_15730);
nand U16953 (N_16953,N_13142,N_14868);
and U16954 (N_16954,N_13799,N_12835);
and U16955 (N_16955,N_13705,N_13436);
nor U16956 (N_16956,N_12656,N_15288);
nand U16957 (N_16957,N_14426,N_14554);
nand U16958 (N_16958,N_13254,N_13401);
or U16959 (N_16959,N_14824,N_12708);
nor U16960 (N_16960,N_15228,N_15517);
nor U16961 (N_16961,N_14711,N_12746);
nor U16962 (N_16962,N_13592,N_15213);
and U16963 (N_16963,N_13253,N_14495);
nor U16964 (N_16964,N_12076,N_12059);
or U16965 (N_16965,N_14568,N_12711);
and U16966 (N_16966,N_14572,N_14680);
xnor U16967 (N_16967,N_14875,N_13838);
or U16968 (N_16968,N_15018,N_12922);
and U16969 (N_16969,N_12471,N_14570);
nor U16970 (N_16970,N_12739,N_15075);
xnor U16971 (N_16971,N_13676,N_15296);
nor U16972 (N_16972,N_12908,N_15030);
nand U16973 (N_16973,N_12109,N_12840);
nand U16974 (N_16974,N_13728,N_12462);
nor U16975 (N_16975,N_15266,N_13468);
xor U16976 (N_16976,N_12782,N_15854);
nand U16977 (N_16977,N_15733,N_15251);
or U16978 (N_16978,N_15235,N_14920);
and U16979 (N_16979,N_15563,N_15354);
and U16980 (N_16980,N_13708,N_14994);
nand U16981 (N_16981,N_14156,N_12549);
nor U16982 (N_16982,N_14514,N_13469);
or U16983 (N_16983,N_15256,N_13052);
nor U16984 (N_16984,N_12688,N_15913);
and U16985 (N_16985,N_13704,N_12248);
nand U16986 (N_16986,N_13488,N_14416);
and U16987 (N_16987,N_13496,N_12806);
nand U16988 (N_16988,N_15924,N_13138);
and U16989 (N_16989,N_15219,N_12354);
nand U16990 (N_16990,N_14228,N_13212);
nor U16991 (N_16991,N_13760,N_13771);
nor U16992 (N_16992,N_15455,N_12592);
nor U16993 (N_16993,N_12902,N_12607);
and U16994 (N_16994,N_13078,N_13032);
nor U16995 (N_16995,N_15846,N_12776);
nand U16996 (N_16996,N_15877,N_12961);
nor U16997 (N_16997,N_15127,N_15281);
nor U16998 (N_16998,N_13985,N_13915);
and U16999 (N_16999,N_14267,N_13956);
xor U17000 (N_17000,N_13973,N_14393);
nand U17001 (N_17001,N_12065,N_12402);
nor U17002 (N_17002,N_13246,N_14120);
or U17003 (N_17003,N_14102,N_14535);
nor U17004 (N_17004,N_12985,N_12942);
nand U17005 (N_17005,N_15551,N_15132);
or U17006 (N_17006,N_12886,N_12061);
or U17007 (N_17007,N_13464,N_14194);
nand U17008 (N_17008,N_13769,N_12350);
nor U17009 (N_17009,N_14540,N_13791);
nor U17010 (N_17010,N_15974,N_13928);
or U17011 (N_17011,N_13252,N_12138);
nand U17012 (N_17012,N_14584,N_13143);
nor U17013 (N_17013,N_13650,N_13507);
xnor U17014 (N_17014,N_15350,N_12124);
and U17015 (N_17015,N_14729,N_14111);
xor U17016 (N_17016,N_14226,N_14327);
nor U17017 (N_17017,N_14932,N_13537);
or U17018 (N_17018,N_12421,N_12862);
nor U17019 (N_17019,N_15761,N_15817);
and U17020 (N_17020,N_12088,N_14069);
or U17021 (N_17021,N_13453,N_13477);
and U17022 (N_17022,N_14259,N_14858);
nor U17023 (N_17023,N_13500,N_12986);
nor U17024 (N_17024,N_14081,N_14953);
nand U17025 (N_17025,N_12320,N_15176);
nand U17026 (N_17026,N_12332,N_13127);
or U17027 (N_17027,N_15954,N_15028);
nor U17028 (N_17028,N_15765,N_15309);
nand U17029 (N_17029,N_15645,N_13645);
and U17030 (N_17030,N_12275,N_13755);
or U17031 (N_17031,N_14180,N_12630);
nand U17032 (N_17032,N_12096,N_12903);
or U17033 (N_17033,N_13487,N_15549);
nor U17034 (N_17034,N_13173,N_13753);
nand U17035 (N_17035,N_13383,N_12964);
nor U17036 (N_17036,N_15849,N_12393);
and U17037 (N_17037,N_13625,N_14773);
nand U17038 (N_17038,N_14695,N_13037);
nand U17039 (N_17039,N_13826,N_14985);
and U17040 (N_17040,N_15206,N_13854);
nand U17041 (N_17041,N_15585,N_12276);
nor U17042 (N_17042,N_12313,N_12910);
and U17043 (N_17043,N_14528,N_15109);
and U17044 (N_17044,N_14007,N_12559);
nand U17045 (N_17045,N_15142,N_14618);
nor U17046 (N_17046,N_15721,N_12064);
or U17047 (N_17047,N_12246,N_12422);
or U17048 (N_17048,N_14313,N_14054);
or U17049 (N_17049,N_15208,N_15531);
and U17050 (N_17050,N_14179,N_15145);
nor U17051 (N_17051,N_14380,N_15327);
and U17052 (N_17052,N_15982,N_13106);
and U17053 (N_17053,N_15008,N_12574);
nor U17054 (N_17054,N_14877,N_13691);
nor U17055 (N_17055,N_12386,N_14879);
nand U17056 (N_17056,N_14050,N_13659);
nor U17057 (N_17057,N_12097,N_15799);
or U17058 (N_17058,N_15277,N_15994);
or U17059 (N_17059,N_15704,N_12858);
nand U17060 (N_17060,N_15931,N_13916);
or U17061 (N_17061,N_14041,N_13750);
or U17062 (N_17062,N_15572,N_14809);
or U17063 (N_17063,N_15600,N_14031);
and U17064 (N_17064,N_14741,N_14238);
or U17065 (N_17065,N_14260,N_15463);
nand U17066 (N_17066,N_13372,N_13082);
or U17067 (N_17067,N_12603,N_14367);
or U17068 (N_17068,N_12045,N_12357);
nor U17069 (N_17069,N_12508,N_15134);
nand U17070 (N_17070,N_14816,N_12546);
and U17071 (N_17071,N_12317,N_14362);
nor U17072 (N_17072,N_14145,N_14500);
nand U17073 (N_17073,N_13170,N_13626);
nor U17074 (N_17074,N_14947,N_15713);
or U17075 (N_17075,N_12407,N_14942);
or U17076 (N_17076,N_15801,N_13829);
nor U17077 (N_17077,N_15294,N_15069);
and U17078 (N_17078,N_12239,N_13565);
xnor U17079 (N_17079,N_12562,N_12216);
and U17080 (N_17080,N_13614,N_15740);
and U17081 (N_17081,N_13426,N_14798);
nand U17082 (N_17082,N_12183,N_14814);
and U17083 (N_17083,N_15812,N_14522);
nand U17084 (N_17084,N_15965,N_12260);
and U17085 (N_17085,N_13329,N_12230);
and U17086 (N_17086,N_13972,N_13337);
and U17087 (N_17087,N_12790,N_13938);
nor U17088 (N_17088,N_14344,N_12141);
nand U17089 (N_17089,N_15389,N_13333);
or U17090 (N_17090,N_15899,N_15237);
or U17091 (N_17091,N_15249,N_13012);
nor U17092 (N_17092,N_12299,N_12206);
nor U17093 (N_17093,N_15594,N_13250);
or U17094 (N_17094,N_14587,N_14623);
and U17095 (N_17095,N_15542,N_15962);
nand U17096 (N_17096,N_15685,N_14631);
and U17097 (N_17097,N_12528,N_15007);
and U17098 (N_17098,N_15609,N_15122);
nand U17099 (N_17099,N_15147,N_12185);
and U17100 (N_17100,N_14510,N_14579);
and U17101 (N_17101,N_12660,N_15282);
and U17102 (N_17102,N_12512,N_13530);
or U17103 (N_17103,N_12159,N_12654);
xor U17104 (N_17104,N_15618,N_13474);
xor U17105 (N_17105,N_12279,N_12963);
and U17106 (N_17106,N_14936,N_12341);
and U17107 (N_17107,N_13833,N_13009);
nor U17108 (N_17108,N_13901,N_14203);
and U17109 (N_17109,N_13273,N_13743);
nor U17110 (N_17110,N_13840,N_14025);
and U17111 (N_17111,N_14772,N_15323);
nand U17112 (N_17112,N_15352,N_13687);
xor U17113 (N_17113,N_15577,N_13560);
and U17114 (N_17114,N_14547,N_12004);
and U17115 (N_17115,N_12579,N_14227);
nor U17116 (N_17116,N_13631,N_13289);
or U17117 (N_17117,N_15311,N_14634);
xnor U17118 (N_17118,N_13581,N_13545);
or U17119 (N_17119,N_14243,N_15695);
nand U17120 (N_17120,N_12595,N_14560);
nand U17121 (N_17121,N_15232,N_13263);
nand U17122 (N_17122,N_13129,N_14469);
nor U17123 (N_17123,N_14516,N_15905);
or U17124 (N_17124,N_12258,N_15823);
nand U17125 (N_17125,N_13819,N_15346);
nand U17126 (N_17126,N_13576,N_14677);
nor U17127 (N_17127,N_15971,N_14197);
and U17128 (N_17128,N_13367,N_12793);
nor U17129 (N_17129,N_13842,N_15392);
nor U17130 (N_17130,N_14747,N_12373);
nor U17131 (N_17131,N_14053,N_12970);
nand U17132 (N_17132,N_12111,N_14622);
and U17133 (N_17133,N_13793,N_14926);
nand U17134 (N_17134,N_12426,N_13661);
and U17135 (N_17135,N_12121,N_12958);
nor U17136 (N_17136,N_13611,N_13696);
or U17137 (N_17137,N_15705,N_15196);
nor U17138 (N_17138,N_13360,N_13001);
nand U17139 (N_17139,N_13984,N_12920);
nor U17140 (N_17140,N_15279,N_13217);
nor U17141 (N_17141,N_15815,N_12997);
nor U17142 (N_17142,N_14751,N_15984);
nand U17143 (N_17143,N_13857,N_15742);
or U17144 (N_17144,N_15940,N_14625);
xor U17145 (N_17145,N_15694,N_13096);
and U17146 (N_17146,N_15520,N_14332);
or U17147 (N_17147,N_13667,N_14317);
xor U17148 (N_17148,N_14453,N_15129);
or U17149 (N_17149,N_13172,N_13855);
nor U17150 (N_17150,N_13203,N_15156);
and U17151 (N_17151,N_15490,N_12646);
nor U17152 (N_17152,N_13264,N_12682);
nand U17153 (N_17153,N_13395,N_15636);
nor U17154 (N_17154,N_13914,N_13154);
nand U17155 (N_17155,N_15508,N_13959);
nor U17156 (N_17156,N_12554,N_14813);
or U17157 (N_17157,N_14810,N_15793);
nand U17158 (N_17158,N_15813,N_12550);
nand U17159 (N_17159,N_13163,N_12645);
and U17160 (N_17160,N_15605,N_15286);
xnor U17161 (N_17161,N_15892,N_15527);
or U17162 (N_17162,N_12015,N_12388);
and U17163 (N_17163,N_13377,N_14599);
or U17164 (N_17164,N_15025,N_15901);
nand U17165 (N_17165,N_13415,N_13073);
and U17166 (N_17166,N_15348,N_13670);
nand U17167 (N_17167,N_15595,N_14205);
and U17168 (N_17168,N_14656,N_14452);
nand U17169 (N_17169,N_13955,N_13924);
and U17170 (N_17170,N_14244,N_13918);
xnor U17171 (N_17171,N_13635,N_12873);
nand U17172 (N_17172,N_14895,N_14311);
xor U17173 (N_17173,N_15254,N_14641);
nor U17174 (N_17174,N_14803,N_14328);
and U17175 (N_17175,N_14972,N_15607);
or U17176 (N_17176,N_13764,N_13536);
or U17177 (N_17177,N_12890,N_13080);
nor U17178 (N_17178,N_13085,N_15675);
or U17179 (N_17179,N_12104,N_15271);
and U17180 (N_17180,N_13064,N_12391);
or U17181 (N_17181,N_13245,N_12413);
nand U17182 (N_17182,N_15113,N_14293);
or U17183 (N_17183,N_15072,N_12934);
and U17184 (N_17184,N_13039,N_15867);
nor U17185 (N_17185,N_15326,N_12524);
nand U17186 (N_17186,N_12927,N_15185);
and U17187 (N_17187,N_12583,N_15258);
xor U17188 (N_17188,N_12187,N_14166);
xor U17189 (N_17189,N_14834,N_12377);
nand U17190 (N_17190,N_13028,N_12257);
and U17191 (N_17191,N_13413,N_15344);
or U17192 (N_17192,N_12949,N_13306);
or U17193 (N_17193,N_13994,N_13235);
nand U17194 (N_17194,N_14282,N_14395);
nand U17195 (N_17195,N_13678,N_14330);
xnor U17196 (N_17196,N_13381,N_13923);
and U17197 (N_17197,N_12853,N_14557);
nand U17198 (N_17198,N_12519,N_14968);
or U17199 (N_17199,N_15035,N_13990);
or U17200 (N_17200,N_12146,N_13307);
nand U17201 (N_17201,N_15462,N_12221);
xnor U17202 (N_17202,N_14739,N_13608);
nor U17203 (N_17203,N_15453,N_15725);
xnor U17204 (N_17204,N_12127,N_13017);
nor U17205 (N_17205,N_13672,N_14507);
nor U17206 (N_17206,N_14459,N_12781);
nor U17207 (N_17207,N_12542,N_12272);
nor U17208 (N_17208,N_15586,N_14255);
and U17209 (N_17209,N_15366,N_13191);
nor U17210 (N_17210,N_15057,N_15186);
nor U17211 (N_17211,N_12749,N_12971);
and U17212 (N_17212,N_12005,N_14382);
or U17213 (N_17213,N_14637,N_15865);
or U17214 (N_17214,N_12464,N_13948);
or U17215 (N_17215,N_13567,N_13392);
nor U17216 (N_17216,N_14169,N_12822);
xor U17217 (N_17217,N_12808,N_13873);
xnor U17218 (N_17218,N_13128,N_12294);
and U17219 (N_17219,N_15229,N_12535);
or U17220 (N_17220,N_15712,N_15074);
or U17221 (N_17221,N_13651,N_12913);
nand U17222 (N_17222,N_15787,N_14690);
and U17223 (N_17223,N_14356,N_15839);
nor U17224 (N_17224,N_14960,N_15753);
nand U17225 (N_17225,N_12117,N_14979);
nor U17226 (N_17226,N_15534,N_12691);
or U17227 (N_17227,N_12880,N_14100);
or U17228 (N_17228,N_15824,N_12897);
and U17229 (N_17229,N_12836,N_12580);
xnor U17230 (N_17230,N_12250,N_15426);
nand U17231 (N_17231,N_13624,N_15005);
nand U17232 (N_17232,N_14038,N_15581);
or U17233 (N_17233,N_14483,N_15598);
nor U17234 (N_17234,N_14882,N_12394);
and U17235 (N_17235,N_14795,N_14978);
or U17236 (N_17236,N_12565,N_14912);
or U17237 (N_17237,N_13278,N_13208);
xor U17238 (N_17238,N_13157,N_13420);
nand U17239 (N_17239,N_13066,N_15570);
nor U17240 (N_17240,N_13610,N_12770);
nor U17241 (N_17241,N_14443,N_14059);
nand U17242 (N_17242,N_14077,N_12231);
and U17243 (N_17243,N_12030,N_13913);
nor U17244 (N_17244,N_14661,N_15103);
nor U17245 (N_17245,N_14065,N_13782);
or U17246 (N_17246,N_12833,N_15381);
xnor U17247 (N_17247,N_14363,N_15521);
nand U17248 (N_17248,N_13588,N_14872);
or U17249 (N_17249,N_15770,N_15553);
or U17250 (N_17250,N_14476,N_14319);
xor U17251 (N_17251,N_12604,N_15606);
or U17252 (N_17252,N_15912,N_13396);
or U17253 (N_17253,N_14188,N_14887);
xor U17254 (N_17254,N_14033,N_14207);
and U17255 (N_17255,N_15797,N_15990);
or U17256 (N_17256,N_15086,N_14651);
nand U17257 (N_17257,N_14088,N_15574);
nand U17258 (N_17258,N_14588,N_13016);
nor U17259 (N_17259,N_12417,N_12953);
and U17260 (N_17260,N_13412,N_13893);
nand U17261 (N_17261,N_12653,N_15863);
and U17262 (N_17262,N_13206,N_14022);
nor U17263 (N_17263,N_13907,N_12627);
xor U17264 (N_17264,N_14562,N_13778);
nand U17265 (N_17265,N_13912,N_12538);
or U17266 (N_17266,N_14857,N_15729);
nor U17267 (N_17267,N_15523,N_13301);
nor U17268 (N_17268,N_13140,N_13094);
nor U17269 (N_17269,N_13075,N_12219);
and U17270 (N_17270,N_13063,N_14095);
and U17271 (N_17271,N_13692,N_14383);
nand U17272 (N_17272,N_13834,N_12369);
or U17273 (N_17273,N_12876,N_14463);
and U17274 (N_17274,N_12533,N_13400);
nor U17275 (N_17275,N_12448,N_14456);
and U17276 (N_17276,N_14172,N_14745);
xnor U17277 (N_17277,N_12778,N_14706);
nand U17278 (N_17278,N_14441,N_14504);
and U17279 (N_17279,N_15612,N_15321);
or U17280 (N_17280,N_13749,N_13450);
nand U17281 (N_17281,N_13638,N_13575);
xnor U17282 (N_17282,N_12914,N_14841);
and U17283 (N_17283,N_13041,N_13114);
nand U17284 (N_17284,N_12775,N_13779);
nand U17285 (N_17285,N_12325,N_12503);
nand U17286 (N_17286,N_15637,N_12905);
or U17287 (N_17287,N_14546,N_15201);
and U17288 (N_17288,N_13110,N_13091);
or U17289 (N_17289,N_14445,N_12001);
xnor U17290 (N_17290,N_15510,N_14770);
or U17291 (N_17291,N_14621,N_12220);
nand U17292 (N_17292,N_15151,N_13585);
and U17293 (N_17293,N_13428,N_14135);
nor U17294 (N_17294,N_13478,N_12039);
or U17295 (N_17295,N_12854,N_15378);
nand U17296 (N_17296,N_14503,N_14744);
nor U17297 (N_17297,N_13721,N_15947);
nand U17298 (N_17298,N_14354,N_13418);
nand U17299 (N_17299,N_13966,N_15818);
xnor U17300 (N_17300,N_12011,N_14515);
and U17301 (N_17301,N_14636,N_12857);
xor U17302 (N_17302,N_12788,N_15316);
nand U17303 (N_17303,N_15666,N_14992);
and U17304 (N_17304,N_13572,N_15945);
xor U17305 (N_17305,N_13689,N_15267);
nand U17306 (N_17306,N_13298,N_13119);
and U17307 (N_17307,N_12409,N_14769);
nor U17308 (N_17308,N_12181,N_12740);
or U17309 (N_17309,N_13748,N_13120);
and U17310 (N_17310,N_12957,N_13587);
and U17311 (N_17311,N_14371,N_12536);
xnor U17312 (N_17312,N_15029,N_13776);
or U17313 (N_17313,N_15561,N_12951);
nor U17314 (N_17314,N_13452,N_13265);
nor U17315 (N_17315,N_13880,N_12893);
nor U17316 (N_17316,N_15064,N_14964);
or U17317 (N_17317,N_13491,N_12368);
xor U17318 (N_17318,N_15771,N_12434);
xor U17319 (N_17319,N_13794,N_13896);
and U17320 (N_17320,N_12943,N_15790);
and U17321 (N_17321,N_12821,N_14919);
nand U17322 (N_17322,N_13808,N_13653);
xnor U17323 (N_17323,N_13856,N_12084);
nand U17324 (N_17324,N_12695,N_15592);
nand U17325 (N_17325,N_12112,N_15926);
nor U17326 (N_17326,N_13200,N_14552);
nor U17327 (N_17327,N_12236,N_15117);
and U17328 (N_17328,N_15632,N_12631);
nand U17329 (N_17329,N_12497,N_15584);
or U17330 (N_17330,N_14413,N_13499);
nor U17331 (N_17331,N_14589,N_12709);
nand U17332 (N_17332,N_15809,N_15431);
and U17333 (N_17333,N_14365,N_13970);
nor U17334 (N_17334,N_13616,N_12486);
or U17335 (N_17335,N_13549,N_13629);
or U17336 (N_17336,N_14140,N_13534);
nor U17337 (N_17337,N_13393,N_14709);
nor U17338 (N_17338,N_15702,N_13494);
nor U17339 (N_17339,N_14397,N_12098);
or U17340 (N_17340,N_14006,N_13934);
nor U17341 (N_17341,N_15939,N_15390);
nor U17342 (N_17342,N_15168,N_15925);
nor U17343 (N_17343,N_13375,N_12431);
or U17344 (N_17344,N_13195,N_12866);
xor U17345 (N_17345,N_14409,N_12189);
or U17346 (N_17346,N_14848,N_15210);
nor U17347 (N_17347,N_15085,N_13932);
or U17348 (N_17348,N_14014,N_14106);
nor U17349 (N_17349,N_12644,N_15437);
xor U17350 (N_17350,N_15320,N_14800);
and U17351 (N_17351,N_12842,N_13099);
or U17352 (N_17352,N_14012,N_12517);
nor U17353 (N_17353,N_13931,N_15593);
nand U17354 (N_17354,N_15202,N_13699);
or U17355 (N_17355,N_13980,N_15828);
and U17356 (N_17356,N_12990,N_14298);
nand U17357 (N_17357,N_15707,N_15016);
and U17358 (N_17358,N_12577,N_12343);
nor U17359 (N_17359,N_15278,N_12483);
nor U17360 (N_17360,N_15646,N_14582);
and U17361 (N_17361,N_14561,N_15063);
and U17362 (N_17362,N_14603,N_13527);
or U17363 (N_17363,N_12849,N_13074);
nand U17364 (N_17364,N_15032,N_15627);
or U17365 (N_17365,N_13295,N_13225);
and U17366 (N_17366,N_13409,N_15308);
nor U17367 (N_17367,N_12848,N_12976);
xor U17368 (N_17368,N_14232,N_13644);
nand U17369 (N_17369,N_13164,N_13097);
and U17370 (N_17370,N_12237,N_12724);
nand U17371 (N_17371,N_14289,N_14003);
nor U17372 (N_17372,N_14998,N_14950);
nand U17373 (N_17373,N_14832,N_12681);
and U17374 (N_17374,N_12278,N_14525);
nor U17375 (N_17375,N_13599,N_13902);
nor U17376 (N_17376,N_14121,N_14840);
or U17377 (N_17377,N_12364,N_12696);
and U17378 (N_17378,N_14696,N_12303);
or U17379 (N_17379,N_12702,N_14073);
and U17380 (N_17380,N_15752,N_13353);
nor U17381 (N_17381,N_13201,N_15727);
nand U17382 (N_17382,N_15066,N_12745);
or U17383 (N_17383,N_15620,N_15284);
nor U17384 (N_17384,N_12352,N_12277);
or U17385 (N_17385,N_15960,N_14261);
or U17386 (N_17386,N_12812,N_13361);
nand U17387 (N_17387,N_12488,N_15864);
xnor U17388 (N_17388,N_13294,N_13824);
nor U17389 (N_17389,N_13618,N_12455);
nand U17390 (N_17390,N_13316,N_15059);
nor U17391 (N_17391,N_15440,N_12200);
or U17392 (N_17392,N_14681,N_13887);
and U17393 (N_17393,N_15936,N_12212);
nor U17394 (N_17394,N_14378,N_13863);
nor U17395 (N_17395,N_12506,N_15516);
nor U17396 (N_17396,N_12929,N_13338);
or U17397 (N_17397,N_12268,N_13268);
and U17398 (N_17398,N_15051,N_15682);
nor U17399 (N_17399,N_15473,N_14048);
nand U17400 (N_17400,N_12705,N_15012);
and U17401 (N_17401,N_14592,N_12831);
or U17402 (N_17402,N_13003,N_15400);
or U17403 (N_17403,N_15446,N_15020);
nor U17404 (N_17404,N_13734,N_13757);
and U17405 (N_17405,N_14076,N_15192);
and U17406 (N_17406,N_12624,N_15464);
and U17407 (N_17407,N_12863,N_13427);
or U17408 (N_17408,N_14430,N_12498);
and U17409 (N_17409,N_14548,N_15644);
nor U17410 (N_17410,N_14458,N_15886);
or U17411 (N_17411,N_14945,N_15356);
nand U17412 (N_17412,N_15782,N_15810);
nor U17413 (N_17413,N_13930,N_12590);
xnor U17414 (N_17414,N_15353,N_15078);
nand U17415 (N_17415,N_15181,N_12623);
and U17416 (N_17416,N_13000,N_13792);
or U17417 (N_17417,N_13034,N_15522);
nand U17418 (N_17418,N_12443,N_12164);
nand U17419 (N_17419,N_15995,N_12223);
or U17420 (N_17420,N_13315,N_12900);
nand U17421 (N_17421,N_13197,N_14198);
and U17422 (N_17422,N_13783,N_14981);
or U17423 (N_17423,N_12768,N_12427);
xor U17424 (N_17424,N_13486,N_13408);
nor U17425 (N_17425,N_13890,N_13292);
nand U17426 (N_17426,N_15108,N_12802);
nor U17427 (N_17427,N_14128,N_12068);
or U17428 (N_17428,N_14060,N_12292);
nor U17429 (N_17429,N_12392,N_13810);
or U17430 (N_17430,N_15050,N_14324);
nor U17431 (N_17431,N_14863,N_12330);
nand U17432 (N_17432,N_14017,N_15399);
nor U17433 (N_17433,N_12385,N_14021);
and U17434 (N_17434,N_12665,N_15184);
or U17435 (N_17435,N_12349,N_12647);
or U17436 (N_17436,N_14734,N_15347);
xor U17437 (N_17437,N_14707,N_13373);
and U17438 (N_17438,N_14704,N_13485);
or U17439 (N_17439,N_12008,N_15958);
nand U17440 (N_17440,N_12923,N_15274);
and U17441 (N_17441,N_14601,N_14446);
or U17442 (N_17442,N_13960,N_12877);
and U17443 (N_17443,N_13323,N_13109);
nand U17444 (N_17444,N_15786,N_15230);
or U17445 (N_17445,N_12430,N_13891);
or U17446 (N_17446,N_12652,N_15783);
nor U17447 (N_17447,N_14545,N_15469);
nand U17448 (N_17448,N_12952,N_14643);
and U17449 (N_17449,N_13954,N_15959);
or U17450 (N_17450,N_14710,N_15608);
or U17451 (N_17451,N_15070,N_13571);
nor U17452 (N_17452,N_13239,N_14925);
nor U17453 (N_17453,N_14660,N_15769);
or U17454 (N_17454,N_15042,N_15676);
nand U17455 (N_17455,N_13510,N_12975);
and U17456 (N_17456,N_14023,N_14716);
nand U17457 (N_17457,N_15981,N_12319);
and U17458 (N_17458,N_13514,N_12830);
nor U17459 (N_17459,N_15115,N_14357);
or U17460 (N_17460,N_13584,N_15345);
and U17461 (N_17461,N_14914,N_12366);
or U17462 (N_17462,N_13662,N_15081);
or U17463 (N_17463,N_12680,N_13883);
nand U17464 (N_17464,N_15429,N_14738);
xor U17465 (N_17465,N_13352,N_14967);
or U17466 (N_17466,N_15649,N_12989);
nand U17467 (N_17467,N_13809,N_14030);
nand U17468 (N_17468,N_14428,N_14058);
nor U17469 (N_17469,N_12641,N_15881);
nor U17470 (N_17470,N_12360,N_13648);
nand U17471 (N_17471,N_15454,N_14153);
nand U17472 (N_17472,N_15130,N_13493);
nor U17473 (N_17473,N_13122,N_15796);
nand U17474 (N_17474,N_14110,N_13103);
nor U17475 (N_17475,N_13958,N_12003);
or U17476 (N_17476,N_14665,N_15833);
or U17477 (N_17477,N_13430,N_14322);
and U17478 (N_17478,N_12898,N_13807);
xnor U17479 (N_17479,N_15559,N_12153);
xor U17480 (N_17480,N_14804,N_15034);
or U17481 (N_17481,N_13007,N_14404);
or U17482 (N_17482,N_15677,N_12203);
nor U17483 (N_17483,N_15529,N_15001);
nand U17484 (N_17484,N_14970,N_12482);
or U17485 (N_17485,N_13384,N_13319);
or U17486 (N_17486,N_14602,N_13886);
nand U17487 (N_17487,N_12626,N_13181);
or U17488 (N_17488,N_12683,N_12311);
or U17489 (N_17489,N_15698,N_15302);
or U17490 (N_17490,N_15975,N_13177);
nor U17491 (N_17491,N_12347,N_14277);
nor U17492 (N_17492,N_14104,N_13030);
or U17493 (N_17493,N_13076,N_13860);
and U17494 (N_17494,N_15002,N_13489);
nand U17495 (N_17495,N_12895,N_14493);
nor U17496 (N_17496,N_13160,N_14898);
nand U17497 (N_17497,N_15036,N_15359);
nand U17498 (N_17498,N_15653,N_15525);
and U17499 (N_17499,N_13508,N_13299);
nand U17500 (N_17500,N_12597,N_15898);
nand U17501 (N_17501,N_13622,N_15118);
nor U17502 (N_17502,N_12410,N_12256);
or U17503 (N_17503,N_14827,N_14635);
nor U17504 (N_17504,N_13369,N_13207);
and U17505 (N_17505,N_15500,N_15911);
nor U17506 (N_17506,N_12655,N_13222);
nor U17507 (N_17507,N_14536,N_15993);
nor U17508 (N_17508,N_14252,N_14722);
nor U17509 (N_17509,N_12704,N_12367);
and U17510 (N_17510,N_15236,N_13165);
nor U17511 (N_17511,N_15777,N_12228);
nand U17512 (N_17512,N_13550,N_13071);
or U17513 (N_17513,N_15672,N_15545);
nand U17514 (N_17514,N_12265,N_13238);
nor U17515 (N_17515,N_12722,N_12819);
nand U17516 (N_17516,N_15056,N_12575);
nand U17517 (N_17517,N_13906,N_13351);
and U17518 (N_17518,N_12541,N_14435);
nand U17519 (N_17519,N_13243,N_13688);
or U17520 (N_17520,N_13798,N_15537);
and U17521 (N_17521,N_15423,N_12634);
nand U17522 (N_17522,N_13062,N_13089);
nand U17523 (N_17523,N_12885,N_12027);
nand U17524 (N_17524,N_15930,N_12081);
and U17525 (N_17525,N_14157,N_13796);
nand U17526 (N_17526,N_13815,N_12476);
nor U17527 (N_17527,N_15433,N_14632);
xor U17528 (N_17528,N_13564,N_14340);
or U17529 (N_17529,N_14993,N_13004);
nand U17530 (N_17530,N_12473,N_12818);
and U17531 (N_17531,N_14134,N_14221);
or U17532 (N_17532,N_12844,N_14190);
nor U17533 (N_17533,N_12993,N_13019);
nor U17534 (N_17534,N_13542,N_13476);
nor U17535 (N_17535,N_14508,N_14220);
xor U17536 (N_17536,N_12380,N_13957);
nor U17537 (N_17537,N_14929,N_15090);
and U17538 (N_17538,N_14448,N_12947);
nor U17539 (N_17539,N_14723,N_15169);
and U17540 (N_17540,N_12160,N_12318);
and U17541 (N_17541,N_15840,N_14271);
nor U17542 (N_17542,N_14118,N_13135);
nand U17543 (N_17543,N_15935,N_15395);
nand U17544 (N_17544,N_14176,N_14909);
or U17545 (N_17545,N_14647,N_13321);
nor U17546 (N_17546,N_14701,N_13167);
xnor U17547 (N_17547,N_14146,N_14103);
nand U17548 (N_17548,N_14411,N_14374);
nor U17549 (N_17549,N_12041,N_15692);
or U17550 (N_17550,N_14136,N_14598);
nand U17551 (N_17551,N_14245,N_13727);
xnor U17552 (N_17552,N_13397,N_15689);
nor U17553 (N_17553,N_14331,N_15651);
and U17554 (N_17554,N_12211,N_15376);
or U17555 (N_17555,N_12002,N_12040);
and U17556 (N_17556,N_15101,N_15435);
nand U17557 (N_17557,N_15748,N_14897);
nand U17558 (N_17558,N_13180,N_14353);
nor U17559 (N_17559,N_14127,N_14791);
and U17560 (N_17560,N_14479,N_13176);
and U17561 (N_17561,N_14352,N_12323);
nor U17562 (N_17562,N_15626,N_12254);
or U17563 (N_17563,N_15784,N_15938);
nand U17564 (N_17564,N_15448,N_13391);
and U17565 (N_17565,N_15335,N_14359);
and U17566 (N_17566,N_13216,N_12701);
nand U17567 (N_17567,N_14474,N_15373);
nand U17568 (N_17568,N_12017,N_15639);
or U17569 (N_17569,N_15768,N_13652);
nand U17570 (N_17570,N_14802,N_15552);
or U17571 (N_17571,N_14346,N_13621);
and U17572 (N_17572,N_12602,N_15964);
xnor U17573 (N_17573,N_12436,N_13344);
nand U17574 (N_17574,N_14143,N_13921);
or U17575 (N_17575,N_13014,N_15781);
nor U17576 (N_17576,N_12926,N_14703);
or U17577 (N_17577,N_15452,N_15970);
xnor U17578 (N_17578,N_13446,N_13925);
nand U17579 (N_17579,N_14439,N_15558);
or U17580 (N_17580,N_13046,N_15451);
or U17581 (N_17581,N_12156,N_12286);
nand U17582 (N_17582,N_13410,N_15401);
or U17583 (N_17583,N_12398,N_12361);
nand U17584 (N_17584,N_12809,N_12983);
or U17585 (N_17585,N_13083,N_12400);
and U17586 (N_17586,N_13578,N_12195);
and U17587 (N_17587,N_13251,N_15273);
and U17588 (N_17588,N_12694,N_14486);
nand U17589 (N_17589,N_15775,N_14178);
xor U17590 (N_17590,N_13899,N_13125);
nand U17591 (N_17591,N_13903,N_12114);
or U17592 (N_17592,N_12342,N_12132);
or U17593 (N_17593,N_13773,N_14930);
xor U17594 (N_17594,N_13098,N_13739);
or U17595 (N_17595,N_12810,N_15656);
nand U17596 (N_17596,N_15126,N_15655);
nand U17597 (N_17597,N_14242,N_15836);
and U17598 (N_17598,N_14917,N_12939);
and U17599 (N_17599,N_12742,N_13112);
nor U17600 (N_17600,N_13444,N_15838);
or U17601 (N_17601,N_14070,N_15887);
and U17602 (N_17602,N_13495,N_14573);
xnor U17603 (N_17603,N_14403,N_13155);
xnor U17604 (N_17604,N_12118,N_14285);
nor U17605 (N_17605,N_15514,N_15153);
or U17606 (N_17606,N_12148,N_14847);
and U17607 (N_17607,N_13561,N_12956);
nand U17608 (N_17608,N_12687,N_15370);
nand U17609 (N_17609,N_15919,N_15802);
nand U17610 (N_17610,N_15654,N_13715);
nor U17611 (N_17611,N_13460,N_15047);
xnor U17612 (N_17612,N_12351,N_12635);
nand U17613 (N_17613,N_15663,N_14163);
and U17614 (N_17614,N_14438,N_14196);
nor U17615 (N_17615,N_12978,N_12773);
xnor U17616 (N_17616,N_15175,N_15205);
xor U17617 (N_17617,N_12904,N_13668);
and U17618 (N_17618,N_15933,N_13513);
nor U17619 (N_17619,N_13961,N_15868);
xor U17620 (N_17620,N_15628,N_13677);
and U17621 (N_17621,N_13894,N_12012);
or U17622 (N_17622,N_15120,N_14361);
and U17623 (N_17623,N_12911,N_12686);
xor U17624 (N_17624,N_15041,N_12140);
nand U17625 (N_17625,N_12333,N_12883);
nor U17626 (N_17626,N_13712,N_14520);
and U17627 (N_17627,N_12621,N_12551);
or U17628 (N_17628,N_12991,N_15837);
and U17629 (N_17629,N_13226,N_12599);
nor U17630 (N_17630,N_14211,N_15590);
and U17631 (N_17631,N_12544,N_15989);
nand U17632 (N_17632,N_13366,N_13260);
nor U17633 (N_17633,N_13646,N_13859);
nor U17634 (N_17634,N_13711,N_13695);
and U17635 (N_17635,N_12382,N_15310);
xnor U17636 (N_17636,N_12861,N_14870);
and U17637 (N_17637,N_12962,N_14275);
nor U17638 (N_17638,N_12408,N_14943);
nand U17639 (N_17639,N_12071,N_13751);
nand U17640 (N_17640,N_13679,N_15976);
nand U17641 (N_17641,N_14421,N_14090);
or U17642 (N_17642,N_13339,N_12122);
and U17643 (N_17643,N_12804,N_15513);
and U17644 (N_17644,N_14650,N_14149);
nor U17645 (N_17645,N_12280,N_13293);
and U17646 (N_17646,N_14590,N_14278);
and U17647 (N_17647,N_13642,N_15460);
nand U17648 (N_17648,N_13286,N_14113);
xnor U17649 (N_17649,N_15855,N_13665);
or U17650 (N_17650,N_12569,N_12516);
nand U17651 (N_17651,N_12545,N_12383);
and U17652 (N_17652,N_13718,N_15601);
nand U17653 (N_17653,N_15342,N_15083);
nand U17654 (N_17654,N_13267,N_13710);
or U17655 (N_17655,N_14158,N_13168);
and U17656 (N_17656,N_13376,N_13320);
or U17657 (N_17657,N_14494,N_13570);
nand U17658 (N_17658,N_15299,N_13772);
nand U17659 (N_17659,N_13324,N_12009);
nand U17660 (N_17660,N_12689,N_13814);
or U17661 (N_17661,N_12548,N_13977);
or U17662 (N_17662,N_14490,N_12306);
or U17663 (N_17663,N_13209,N_15112);
or U17664 (N_17664,N_14922,N_13266);
and U17665 (N_17665,N_13079,N_15821);
or U17666 (N_17666,N_12450,N_15918);
and U17667 (N_17667,N_14454,N_12736);
nor U17668 (N_17668,N_15484,N_13021);
nor U17669 (N_17669,N_13864,N_15477);
or U17670 (N_17670,N_15548,N_14537);
or U17671 (N_17671,N_14234,N_12611);
and U17672 (N_17672,N_15033,N_13577);
or U17673 (N_17673,N_14225,N_13095);
or U17674 (N_17674,N_14616,N_14797);
nor U17675 (N_17675,N_13284,N_12155);
xor U17676 (N_17676,N_15049,N_12591);
and U17677 (N_17677,N_14691,N_14668);
xor U17678 (N_17678,N_12845,N_13414);
xor U17679 (N_17679,N_14016,N_15642);
nand U17680 (N_17680,N_13044,N_12678);
and U17681 (N_17681,N_15290,N_13202);
or U17682 (N_17682,N_14199,N_12020);
nand U17683 (N_17683,N_12441,N_15526);
nand U17684 (N_17684,N_15349,N_12543);
xor U17685 (N_17685,N_13406,N_15382);
nand U17686 (N_17686,N_14892,N_15619);
and U17687 (N_17687,N_14339,N_14294);
nand U17688 (N_17688,N_13882,N_13900);
or U17689 (N_17689,N_14902,N_13554);
nor U17690 (N_17690,N_13158,N_13919);
and U17691 (N_17691,N_14679,N_14151);
nand U17692 (N_17692,N_12712,N_14161);
nand U17693 (N_17693,N_14256,N_12730);
nor U17694 (N_17694,N_14475,N_12177);
or U17695 (N_17695,N_13092,N_15554);
and U17696 (N_17696,N_15138,N_14085);
or U17697 (N_17697,N_13365,N_12131);
xnor U17698 (N_17698,N_13555,N_15420);
xnor U17699 (N_17699,N_13156,N_13190);
nand U17700 (N_17700,N_14291,N_12021);
xor U17701 (N_17701,N_15221,N_14071);
nand U17702 (N_17702,N_12643,N_14247);
or U17703 (N_17703,N_12832,N_15116);
nand U17704 (N_17704,N_13861,N_13528);
nand U17705 (N_17705,N_14210,N_14851);
nand U17706 (N_17706,N_14512,N_13713);
and U17707 (N_17707,N_12115,N_13447);
and U17708 (N_17708,N_14233,N_14694);
or U17709 (N_17709,N_15703,N_12190);
nor U17710 (N_17710,N_14854,N_14821);
xnor U17711 (N_17711,N_13228,N_13022);
or U17712 (N_17712,N_13908,N_13612);
and U17713 (N_17713,N_14481,N_15895);
or U17714 (N_17714,N_14109,N_14761);
nand U17715 (N_17715,N_15505,N_14035);
nand U17716 (N_17716,N_13006,N_12033);
and U17717 (N_17717,N_14116,N_14952);
or U17718 (N_17718,N_13558,N_14191);
xor U17719 (N_17719,N_12289,N_14099);
or U17720 (N_17720,N_13036,N_15157);
nand U17721 (N_17721,N_13449,N_15550);
nand U17722 (N_17722,N_14855,N_13816);
nand U17723 (N_17723,N_12090,N_15319);
or U17724 (N_17724,N_12679,N_15371);
and U17725 (N_17725,N_12044,N_12202);
nor U17726 (N_17726,N_12737,N_12046);
nor U17727 (N_17727,N_14498,N_15909);
nor U17728 (N_17728,N_15097,N_13287);
or U17729 (N_17729,N_13790,N_14954);
nand U17730 (N_17730,N_15541,N_15903);
and U17731 (N_17731,N_13634,N_13845);
and U17732 (N_17732,N_12520,N_15471);
or U17733 (N_17733,N_15511,N_13314);
nor U17734 (N_17734,N_12649,N_12224);
or U17735 (N_17735,N_15535,N_14884);
and U17736 (N_17736,N_14692,N_15478);
nor U17737 (N_17737,N_14717,N_13350);
nor U17738 (N_17738,N_13690,N_14543);
and U17739 (N_17739,N_13187,N_14682);
and U17740 (N_17740,N_12474,N_14237);
xnor U17741 (N_17741,N_13280,N_12834);
and U17742 (N_17742,N_12522,N_15111);
nor U17743 (N_17743,N_15331,N_12573);
nand U17744 (N_17744,N_12481,N_13841);
and U17745 (N_17745,N_15259,N_12891);
and U17746 (N_17746,N_15004,N_12973);
nand U17747 (N_17747,N_15776,N_14918);
nand U17748 (N_17748,N_13236,N_13722);
and U17749 (N_17749,N_15825,N_14675);
or U17750 (N_17750,N_14806,N_12355);
nand U17751 (N_17751,N_13851,N_14513);
nand U17752 (N_17752,N_15880,N_14931);
nor U17753 (N_17753,N_15803,N_13830);
and U17754 (N_17754,N_14358,N_13867);
nand U17755 (N_17755,N_12826,N_15470);
nand U17756 (N_17756,N_14091,N_13237);
nor U17757 (N_17757,N_14316,N_13898);
nor U17758 (N_17758,N_12322,N_14980);
and U17759 (N_17759,N_14315,N_14171);
or U17760 (N_17760,N_15040,N_12099);
or U17761 (N_17761,N_14249,N_15189);
nor U17762 (N_17762,N_15253,N_14530);
xor U17763 (N_17763,N_12149,N_12321);
nor U17764 (N_17764,N_14184,N_15393);
or U17765 (N_17765,N_13868,N_13747);
and U17766 (N_17766,N_14152,N_13825);
and U17767 (N_17767,N_13276,N_12457);
xnor U17768 (N_17768,N_14341,N_14689);
nor U17769 (N_17769,N_14306,N_12429);
and U17770 (N_17770,N_14878,N_15077);
or U17771 (N_17771,N_13640,N_14132);
nor U17772 (N_17772,N_14154,N_12767);
nand U17773 (N_17773,N_15944,N_15360);
nor U17774 (N_17774,N_15248,N_15573);
or U17775 (N_17775,N_15224,N_12874);
nand U17776 (N_17776,N_14408,N_15673);
nor U17777 (N_17777,N_15141,N_13949);
nor U17778 (N_17778,N_13057,N_15387);
and U17779 (N_17779,N_12919,N_14034);
nor U17780 (N_17780,N_15148,N_15166);
nor U17781 (N_17781,N_12133,N_15724);
and U17782 (N_17782,N_14782,N_15509);
nor U17783 (N_17783,N_14578,N_14789);
and U17784 (N_17784,N_13448,N_12253);
and U17785 (N_17785,N_15480,N_15853);
and U17786 (N_17786,N_15089,N_13144);
or U17787 (N_17787,N_15080,N_15988);
or U17788 (N_17788,N_14905,N_13223);
xor U17789 (N_17789,N_14678,N_12144);
nor U17790 (N_17790,N_14297,N_15662);
or U17791 (N_17791,N_13758,N_15088);
nand U17792 (N_17792,N_14752,N_13591);
and U17793 (N_17793,N_15287,N_13179);
or U17794 (N_17794,N_12103,N_13666);
nor U17795 (N_17795,N_14068,N_13481);
nand U17796 (N_17796,N_12080,N_15182);
or U17797 (N_17797,N_14379,N_12585);
or U17798 (N_17798,N_13240,N_14398);
and U17799 (N_17799,N_12304,N_13141);
and U17800 (N_17800,N_15957,N_15339);
or U17801 (N_17801,N_13511,N_15494);
nand U17802 (N_17802,N_15133,N_15621);
and U17803 (N_17803,N_12879,N_12293);
xnor U17804 (N_17804,N_12872,N_13605);
and U17805 (N_17805,N_15332,N_12974);
or U17806 (N_17806,N_13566,N_13979);
xnor U17807 (N_17807,N_12281,N_14406);
nand U17808 (N_17808,N_15459,N_14263);
nand U17809 (N_17809,N_14320,N_13884);
and U17810 (N_17810,N_14614,N_15244);
nor U17811 (N_17811,N_12757,N_13433);
nor U17812 (N_17812,N_13059,N_15530);
nor U17813 (N_17813,N_15613,N_15131);
or U17814 (N_17814,N_13802,N_15017);
and U17815 (N_17815,N_15571,N_12465);
nand U17816 (N_17816,N_14990,N_14123);
or U17817 (N_17817,N_12070,N_15268);
nor U17818 (N_17818,N_13398,N_14137);
or U17819 (N_17819,N_13735,N_12077);
xor U17820 (N_17820,N_15165,N_15949);
nor U17821 (N_17821,N_15255,N_13987);
and U17822 (N_17822,N_12445,N_12120);
or U17823 (N_17823,N_12331,N_12552);
or U17824 (N_17824,N_13756,N_15841);
xor U17825 (N_17825,N_15602,N_15528);
or U17826 (N_17826,N_15476,N_13183);
xnor U17827 (N_17827,N_14648,N_13475);
nand U17828 (N_17828,N_13504,N_12406);
and U17829 (N_17829,N_12405,N_12358);
nand U17830 (N_17830,N_15641,N_14754);
nor U17831 (N_17831,N_15997,N_15506);
xnor U17832 (N_17832,N_13132,N_14375);
xnor U17833 (N_17833,N_15037,N_14138);
nand U17834 (N_17834,N_12582,N_13387);
nand U17835 (N_17835,N_12477,N_14594);
and U17836 (N_17836,N_13895,N_12996);
or U17837 (N_17837,N_15504,N_14082);
or U17838 (N_17838,N_13673,N_13185);
xor U17839 (N_17839,N_15383,N_12829);
or U17840 (N_17840,N_13812,N_13026);
and U17841 (N_17841,N_13717,N_15280);
nor U17842 (N_17842,N_14615,N_13419);
nor U17843 (N_17843,N_12933,N_12633);
xnor U17844 (N_17844,N_13682,N_12269);
or U17845 (N_17845,N_12540,N_13404);
or U17846 (N_17846,N_13121,N_12134);
xnor U17847 (N_17847,N_12379,N_12328);
nand U17848 (N_17848,N_14183,N_13568);
and U17849 (N_17849,N_13394,N_14671);
nand U17850 (N_17850,N_12941,N_14604);
nor U17851 (N_17851,N_15920,N_14749);
and U17852 (N_17852,N_13632,N_13072);
or U17853 (N_17853,N_13330,N_12271);
xor U17854 (N_17854,N_12659,N_13146);
nor U17855 (N_17855,N_15123,N_14533);
or U17856 (N_17856,N_13997,N_15394);
nor U17857 (N_17857,N_12168,N_15325);
nand U17858 (N_17858,N_12931,N_15640);
nor U17859 (N_17859,N_12083,N_13905);
or U17860 (N_17860,N_12057,N_12733);
nor U17861 (N_17861,N_13720,N_14372);
nor U17862 (N_17862,N_15167,N_15412);
or U17863 (N_17863,N_13370,N_14442);
or U17864 (N_17864,N_15297,N_14186);
or U17865 (N_17865,N_15884,N_14983);
nand U17866 (N_17866,N_15384,N_13828);
nor U17867 (N_17867,N_15969,N_12031);
or U17868 (N_17868,N_14173,N_13013);
or U17869 (N_17869,N_14270,N_13613);
xor U17870 (N_17870,N_15364,N_13194);
xnor U17871 (N_17871,N_15170,N_12731);
nand U17872 (N_17872,N_12197,N_15159);
nor U17873 (N_17873,N_12735,N_13524);
nand U17874 (N_17874,N_14666,N_15467);
xnor U17875 (N_17875,N_15582,N_13341);
nor U17876 (N_17876,N_12950,N_15916);
or U17877 (N_17877,N_12846,N_13257);
nor U17878 (N_17878,N_14645,N_14896);
and U17879 (N_17879,N_15876,N_15789);
nand U17880 (N_17880,N_14629,N_15487);
and U17881 (N_17881,N_12723,N_15498);
and U17882 (N_17882,N_15891,N_13693);
xor U17883 (N_17883,N_13910,N_15061);
or U17884 (N_17884,N_13529,N_14830);
or U17885 (N_17885,N_12137,N_12418);
xor U17886 (N_17886,N_14923,N_14765);
or U17887 (N_17887,N_14274,N_13847);
nor U17888 (N_17888,N_12892,N_15318);
or U17889 (N_17889,N_12881,N_13871);
or U17890 (N_17890,N_12487,N_14101);
nand U17891 (N_17891,N_12780,N_13331);
nand U17892 (N_17892,N_12727,N_14390);
or U17893 (N_17893,N_15027,N_14580);
xor U17894 (N_17894,N_14826,N_12389);
or U17895 (N_17895,N_13466,N_15638);
or U17896 (N_17896,N_13229,N_14753);
nand U17897 (N_17897,N_15411,N_13926);
and U17898 (N_17898,N_12438,N_13291);
and U17899 (N_17899,N_14519,N_12016);
nor U17900 (N_17900,N_14308,N_12710);
or U17901 (N_17901,N_13303,N_15710);
nor U17902 (N_17902,N_15187,N_15174);
nand U17903 (N_17903,N_13627,N_12186);
and U17904 (N_17904,N_15999,N_14305);
and U17905 (N_17905,N_13594,N_15946);
nand U17906 (N_17906,N_14743,N_13989);
or U17907 (N_17907,N_14899,N_12968);
nand U17908 (N_17908,N_12204,N_14626);
nand U17909 (N_17909,N_15246,N_12937);
nand U17910 (N_17910,N_12440,N_15928);
nand U17911 (N_17911,N_13869,N_14057);
xor U17912 (N_17912,N_14213,N_12215);
or U17913 (N_17913,N_13992,N_13364);
and U17914 (N_17914,N_12564,N_12674);
and U17915 (N_17915,N_14074,N_13559);
nor U17916 (N_17916,N_14869,N_15883);
and U17917 (N_17917,N_13193,N_15746);
xnor U17918 (N_17918,N_13971,N_14432);
nand U17919 (N_17919,N_12801,N_13296);
and U17920 (N_17920,N_12959,N_15792);
nor U17921 (N_17921,N_15681,N_12047);
or U17922 (N_17922,N_14488,N_12847);
or U17923 (N_17923,N_14784,N_12113);
nand U17924 (N_17924,N_12226,N_12667);
nand U17925 (N_17925,N_15291,N_13563);
nor U17926 (N_17926,N_14477,N_12500);
and U17927 (N_17927,N_13011,N_15338);
or U17928 (N_17928,N_14793,N_14781);
xnor U17929 (N_17929,N_12511,N_14373);
nor U17930 (N_17930,N_13607,N_12526);
and U17931 (N_17931,N_15285,N_12771);
xor U17932 (N_17932,N_14303,N_13069);
nor U17933 (N_17933,N_15831,N_14938);
nor U17934 (N_17934,N_14201,N_14742);
and U17935 (N_17935,N_14837,N_12209);
or U17936 (N_17936,N_15795,N_13546);
and U17937 (N_17937,N_13184,N_13740);
nor U17938 (N_17938,N_14642,N_13300);
nand U17939 (N_17939,N_14018,N_14290);
nor U17940 (N_17940,N_15546,N_15544);
nor U17941 (N_17941,N_15745,N_14965);
nor U17942 (N_17942,N_14107,N_12671);
nor U17943 (N_17943,N_12615,N_13431);
nand U17944 (N_17944,N_13290,N_14343);
nand U17945 (N_17945,N_13765,N_15560);
nand U17946 (N_17946,N_12539,N_15955);
nor U17947 (N_17947,N_13639,N_14524);
or U17948 (N_17948,N_12753,N_13993);
and U17949 (N_17949,N_13305,N_14842);
nand U17950 (N_17950,N_15829,N_14685);
or U17951 (N_17951,N_14342,N_13126);
and U17952 (N_17952,N_14755,N_13835);
nor U17953 (N_17953,N_14309,N_13498);
and U17954 (N_17954,N_13458,N_13029);
or U17955 (N_17955,N_14951,N_14436);
and U17956 (N_17956,N_12714,N_15094);
nand U17957 (N_17957,N_13313,N_14209);
nand U17958 (N_17958,N_14336,N_15680);
or U17959 (N_17959,N_12489,N_14880);
nand U17960 (N_17960,N_13744,N_15155);
and U17961 (N_17961,N_13797,N_14141);
nor U17962 (N_17962,N_12437,N_15104);
nand U17963 (N_17963,N_15262,N_13107);
nand U17964 (N_17964,N_13470,N_13136);
and U17965 (N_17965,N_15791,N_14986);
or U17966 (N_17966,N_14288,N_14836);
and U17967 (N_17967,N_13378,N_15735);
and U17968 (N_17968,N_12918,N_14805);
and U17969 (N_17969,N_14310,N_14147);
or U17970 (N_17970,N_15330,N_13967);
and U17971 (N_17971,N_13492,N_15758);
or U17972 (N_17972,N_15805,N_13655);
or U17973 (N_17973,N_13836,N_14808);
nand U17974 (N_17974,N_12670,N_14231);
or U17975 (N_17975,N_15405,N_15532);
and U17976 (N_17976,N_12490,N_14283);
and U17977 (N_17977,N_14730,N_15445);
or U17978 (N_17978,N_15082,N_12147);
nor U17979 (N_17979,N_13055,N_12805);
nor U17980 (N_17980,N_15062,N_14852);
or U17981 (N_17981,N_14447,N_14422);
and U17982 (N_17982,N_12732,N_15301);
nor U17983 (N_17983,N_13843,N_14768);
and U17984 (N_17984,N_15754,N_12478);
and U17985 (N_17985,N_13390,N_14241);
nor U17986 (N_17986,N_14505,N_14687);
nand U17987 (N_17987,N_13630,N_14266);
nor U17988 (N_17988,N_13746,N_12820);
nor U17989 (N_17989,N_14192,N_13515);
nor U17990 (N_17990,N_15910,N_14999);
or U17991 (N_17991,N_15161,N_12252);
nand U17992 (N_17992,N_12284,N_13684);
nand U17993 (N_17993,N_15963,N_14222);
nand U17994 (N_17994,N_15367,N_13439);
xor U17995 (N_17995,N_12461,N_14534);
xnor U17996 (N_17996,N_13831,N_15052);
nor U17997 (N_17997,N_12374,N_15491);
nor U17998 (N_17998,N_15780,N_13862);
and U17999 (N_17999,N_14296,N_15479);
nand U18000 (N_18000,N_12224,N_14702);
nor U18001 (N_18001,N_15357,N_13264);
xnor U18002 (N_18002,N_12910,N_14043);
nand U18003 (N_18003,N_13379,N_13996);
nor U18004 (N_18004,N_12483,N_12914);
nor U18005 (N_18005,N_13181,N_15614);
and U18006 (N_18006,N_12734,N_14041);
nand U18007 (N_18007,N_14696,N_15566);
nor U18008 (N_18008,N_14497,N_14184);
nand U18009 (N_18009,N_13941,N_15478);
nand U18010 (N_18010,N_13340,N_12001);
and U18011 (N_18011,N_13655,N_12104);
nand U18012 (N_18012,N_13326,N_14825);
nand U18013 (N_18013,N_15087,N_15522);
and U18014 (N_18014,N_14273,N_13008);
xnor U18015 (N_18015,N_12129,N_13231);
nand U18016 (N_18016,N_12447,N_12720);
nor U18017 (N_18017,N_15824,N_13933);
or U18018 (N_18018,N_14143,N_14186);
nand U18019 (N_18019,N_15706,N_12248);
nand U18020 (N_18020,N_15007,N_13981);
nand U18021 (N_18021,N_13096,N_14238);
xor U18022 (N_18022,N_13323,N_15618);
nor U18023 (N_18023,N_15178,N_12650);
or U18024 (N_18024,N_15687,N_15554);
nand U18025 (N_18025,N_14171,N_14927);
nand U18026 (N_18026,N_14301,N_14489);
and U18027 (N_18027,N_13806,N_12107);
nor U18028 (N_18028,N_15623,N_14482);
and U18029 (N_18029,N_15784,N_14744);
nor U18030 (N_18030,N_13952,N_15035);
nand U18031 (N_18031,N_14276,N_15679);
or U18032 (N_18032,N_12884,N_14442);
and U18033 (N_18033,N_15842,N_13281);
or U18034 (N_18034,N_14178,N_14242);
nor U18035 (N_18035,N_13946,N_14134);
and U18036 (N_18036,N_14041,N_13564);
xnor U18037 (N_18037,N_14468,N_15806);
nor U18038 (N_18038,N_15572,N_12918);
and U18039 (N_18039,N_14030,N_14322);
and U18040 (N_18040,N_15245,N_14933);
nor U18041 (N_18041,N_12276,N_15857);
nand U18042 (N_18042,N_13926,N_12908);
nand U18043 (N_18043,N_14991,N_13396);
nor U18044 (N_18044,N_15367,N_15140);
nor U18045 (N_18045,N_12056,N_14644);
and U18046 (N_18046,N_12475,N_12939);
or U18047 (N_18047,N_13651,N_14046);
or U18048 (N_18048,N_14660,N_14385);
and U18049 (N_18049,N_13232,N_12901);
xnor U18050 (N_18050,N_15292,N_12735);
or U18051 (N_18051,N_14817,N_15993);
xor U18052 (N_18052,N_14554,N_12979);
nand U18053 (N_18053,N_15987,N_15308);
and U18054 (N_18054,N_12437,N_13562);
nand U18055 (N_18055,N_14295,N_12000);
xnor U18056 (N_18056,N_14916,N_13368);
nor U18057 (N_18057,N_15379,N_15018);
and U18058 (N_18058,N_15498,N_12060);
nor U18059 (N_18059,N_12511,N_15827);
nand U18060 (N_18060,N_12964,N_13209);
and U18061 (N_18061,N_14198,N_13447);
and U18062 (N_18062,N_15849,N_12999);
and U18063 (N_18063,N_12646,N_13112);
nor U18064 (N_18064,N_12050,N_15115);
or U18065 (N_18065,N_12212,N_15105);
nand U18066 (N_18066,N_14403,N_14969);
and U18067 (N_18067,N_13345,N_13151);
nand U18068 (N_18068,N_15466,N_13264);
xor U18069 (N_18069,N_12610,N_15808);
nor U18070 (N_18070,N_12036,N_12948);
xnor U18071 (N_18071,N_13371,N_14193);
xor U18072 (N_18072,N_13409,N_13864);
nand U18073 (N_18073,N_13144,N_12542);
nand U18074 (N_18074,N_14874,N_13081);
and U18075 (N_18075,N_12871,N_12430);
or U18076 (N_18076,N_12116,N_14474);
or U18077 (N_18077,N_15685,N_12065);
and U18078 (N_18078,N_15616,N_13174);
or U18079 (N_18079,N_15361,N_15786);
nor U18080 (N_18080,N_14967,N_13142);
nand U18081 (N_18081,N_13817,N_13599);
or U18082 (N_18082,N_12086,N_14499);
and U18083 (N_18083,N_13784,N_14028);
nand U18084 (N_18084,N_13768,N_15600);
nor U18085 (N_18085,N_12040,N_14328);
nor U18086 (N_18086,N_13296,N_14299);
or U18087 (N_18087,N_13232,N_12898);
nand U18088 (N_18088,N_12632,N_15444);
and U18089 (N_18089,N_12628,N_12298);
xor U18090 (N_18090,N_14944,N_13390);
nand U18091 (N_18091,N_15531,N_13469);
xor U18092 (N_18092,N_14706,N_13562);
and U18093 (N_18093,N_15212,N_12921);
and U18094 (N_18094,N_13141,N_14696);
xor U18095 (N_18095,N_12367,N_14699);
nor U18096 (N_18096,N_13172,N_15212);
and U18097 (N_18097,N_13159,N_15497);
xnor U18098 (N_18098,N_15723,N_12179);
nor U18099 (N_18099,N_12620,N_13515);
nor U18100 (N_18100,N_14654,N_15671);
xnor U18101 (N_18101,N_14584,N_13584);
or U18102 (N_18102,N_12806,N_12013);
and U18103 (N_18103,N_13990,N_12258);
or U18104 (N_18104,N_15080,N_13001);
nor U18105 (N_18105,N_13324,N_13185);
or U18106 (N_18106,N_15560,N_13915);
nor U18107 (N_18107,N_13448,N_14372);
and U18108 (N_18108,N_13009,N_14732);
nand U18109 (N_18109,N_12718,N_15217);
xnor U18110 (N_18110,N_14217,N_14120);
and U18111 (N_18111,N_13386,N_12884);
or U18112 (N_18112,N_15072,N_15820);
or U18113 (N_18113,N_12678,N_14451);
or U18114 (N_18114,N_13908,N_15914);
nor U18115 (N_18115,N_14384,N_14803);
xnor U18116 (N_18116,N_14530,N_13568);
or U18117 (N_18117,N_13025,N_14182);
nor U18118 (N_18118,N_15045,N_14638);
or U18119 (N_18119,N_12089,N_13525);
nand U18120 (N_18120,N_15340,N_15216);
and U18121 (N_18121,N_14115,N_13581);
nor U18122 (N_18122,N_12428,N_14775);
nand U18123 (N_18123,N_15379,N_14477);
nand U18124 (N_18124,N_15670,N_12579);
and U18125 (N_18125,N_15998,N_13348);
or U18126 (N_18126,N_13246,N_12521);
or U18127 (N_18127,N_15263,N_15563);
and U18128 (N_18128,N_13299,N_14670);
and U18129 (N_18129,N_14951,N_15982);
nor U18130 (N_18130,N_13280,N_14810);
nand U18131 (N_18131,N_13351,N_12071);
xnor U18132 (N_18132,N_14615,N_13653);
or U18133 (N_18133,N_13893,N_13239);
nor U18134 (N_18134,N_15220,N_14036);
nor U18135 (N_18135,N_13746,N_13904);
or U18136 (N_18136,N_15564,N_12608);
nor U18137 (N_18137,N_12963,N_13334);
xnor U18138 (N_18138,N_12355,N_14522);
nand U18139 (N_18139,N_13865,N_15301);
nand U18140 (N_18140,N_12942,N_12152);
and U18141 (N_18141,N_13072,N_15759);
or U18142 (N_18142,N_12102,N_14150);
xnor U18143 (N_18143,N_15060,N_15175);
nor U18144 (N_18144,N_12184,N_15826);
nand U18145 (N_18145,N_15458,N_14410);
and U18146 (N_18146,N_12653,N_13888);
or U18147 (N_18147,N_15343,N_14972);
or U18148 (N_18148,N_15683,N_12153);
and U18149 (N_18149,N_15445,N_15915);
or U18150 (N_18150,N_12383,N_12217);
and U18151 (N_18151,N_12554,N_15910);
nand U18152 (N_18152,N_12637,N_15000);
nor U18153 (N_18153,N_13448,N_12679);
nand U18154 (N_18154,N_15323,N_14849);
xnor U18155 (N_18155,N_12191,N_14961);
or U18156 (N_18156,N_15168,N_13051);
and U18157 (N_18157,N_14728,N_14065);
nand U18158 (N_18158,N_13045,N_14579);
nor U18159 (N_18159,N_15369,N_15822);
or U18160 (N_18160,N_12496,N_14520);
and U18161 (N_18161,N_15478,N_15766);
or U18162 (N_18162,N_12644,N_13250);
nor U18163 (N_18163,N_14691,N_13272);
xnor U18164 (N_18164,N_13859,N_15016);
nor U18165 (N_18165,N_15224,N_14017);
nand U18166 (N_18166,N_15254,N_14605);
and U18167 (N_18167,N_14735,N_13579);
or U18168 (N_18168,N_15607,N_12262);
nor U18169 (N_18169,N_13021,N_12962);
or U18170 (N_18170,N_15226,N_12091);
nor U18171 (N_18171,N_12994,N_13540);
nand U18172 (N_18172,N_14825,N_14310);
and U18173 (N_18173,N_12322,N_13520);
and U18174 (N_18174,N_15102,N_14590);
or U18175 (N_18175,N_14138,N_14364);
or U18176 (N_18176,N_12921,N_13803);
or U18177 (N_18177,N_15112,N_14176);
or U18178 (N_18178,N_13889,N_13916);
and U18179 (N_18179,N_14214,N_14270);
xor U18180 (N_18180,N_13141,N_12516);
or U18181 (N_18181,N_12258,N_14720);
nand U18182 (N_18182,N_15132,N_12153);
nand U18183 (N_18183,N_13489,N_13414);
nor U18184 (N_18184,N_12376,N_15195);
and U18185 (N_18185,N_12240,N_14661);
nand U18186 (N_18186,N_13134,N_14857);
and U18187 (N_18187,N_13880,N_14273);
or U18188 (N_18188,N_13984,N_14697);
and U18189 (N_18189,N_14715,N_13112);
nand U18190 (N_18190,N_15534,N_12938);
nand U18191 (N_18191,N_14043,N_13747);
nand U18192 (N_18192,N_15864,N_12201);
and U18193 (N_18193,N_12739,N_15498);
nor U18194 (N_18194,N_12052,N_13575);
or U18195 (N_18195,N_15106,N_13736);
and U18196 (N_18196,N_15812,N_12515);
and U18197 (N_18197,N_13076,N_15872);
and U18198 (N_18198,N_15638,N_14828);
nand U18199 (N_18199,N_12073,N_13748);
nand U18200 (N_18200,N_14264,N_12250);
or U18201 (N_18201,N_15477,N_12141);
nand U18202 (N_18202,N_12265,N_15600);
and U18203 (N_18203,N_12590,N_13253);
nor U18204 (N_18204,N_15434,N_13964);
or U18205 (N_18205,N_13824,N_15220);
or U18206 (N_18206,N_14424,N_13093);
or U18207 (N_18207,N_13450,N_14817);
nand U18208 (N_18208,N_15068,N_15142);
or U18209 (N_18209,N_15741,N_14035);
and U18210 (N_18210,N_13597,N_15624);
nor U18211 (N_18211,N_15037,N_12721);
nor U18212 (N_18212,N_12221,N_14946);
or U18213 (N_18213,N_13087,N_14820);
nand U18214 (N_18214,N_13566,N_14142);
and U18215 (N_18215,N_12135,N_12158);
nor U18216 (N_18216,N_15859,N_12818);
nor U18217 (N_18217,N_14973,N_12137);
nand U18218 (N_18218,N_13479,N_12846);
nand U18219 (N_18219,N_14326,N_12411);
or U18220 (N_18220,N_12777,N_12566);
and U18221 (N_18221,N_15444,N_12968);
or U18222 (N_18222,N_15324,N_15246);
or U18223 (N_18223,N_12455,N_15383);
or U18224 (N_18224,N_14869,N_12150);
nand U18225 (N_18225,N_14287,N_12337);
nor U18226 (N_18226,N_12981,N_15860);
xor U18227 (N_18227,N_14521,N_12864);
and U18228 (N_18228,N_14112,N_15903);
nand U18229 (N_18229,N_15687,N_13312);
or U18230 (N_18230,N_12698,N_13960);
nor U18231 (N_18231,N_12118,N_15163);
xor U18232 (N_18232,N_13576,N_13869);
and U18233 (N_18233,N_14626,N_14961);
nor U18234 (N_18234,N_13571,N_14613);
nand U18235 (N_18235,N_15570,N_13765);
and U18236 (N_18236,N_15962,N_15171);
or U18237 (N_18237,N_14486,N_12657);
nor U18238 (N_18238,N_13271,N_14504);
or U18239 (N_18239,N_15990,N_12324);
nor U18240 (N_18240,N_15600,N_12437);
nand U18241 (N_18241,N_15152,N_14333);
and U18242 (N_18242,N_15982,N_15747);
xor U18243 (N_18243,N_12685,N_13288);
nor U18244 (N_18244,N_15500,N_12984);
or U18245 (N_18245,N_13291,N_14815);
nor U18246 (N_18246,N_12192,N_13551);
xnor U18247 (N_18247,N_15153,N_15037);
nor U18248 (N_18248,N_12464,N_13371);
nand U18249 (N_18249,N_13780,N_15583);
nand U18250 (N_18250,N_14857,N_13845);
nand U18251 (N_18251,N_14318,N_14625);
nor U18252 (N_18252,N_12577,N_15429);
and U18253 (N_18253,N_13126,N_12972);
xor U18254 (N_18254,N_12901,N_12832);
nor U18255 (N_18255,N_12494,N_13457);
nand U18256 (N_18256,N_12016,N_12565);
or U18257 (N_18257,N_15501,N_13912);
or U18258 (N_18258,N_12519,N_14761);
or U18259 (N_18259,N_15394,N_15900);
or U18260 (N_18260,N_12028,N_15177);
nand U18261 (N_18261,N_13018,N_14622);
and U18262 (N_18262,N_14366,N_12621);
and U18263 (N_18263,N_15285,N_14665);
or U18264 (N_18264,N_15338,N_14658);
or U18265 (N_18265,N_13653,N_13248);
nand U18266 (N_18266,N_14110,N_12211);
or U18267 (N_18267,N_12022,N_13271);
or U18268 (N_18268,N_14147,N_12739);
or U18269 (N_18269,N_14609,N_14923);
and U18270 (N_18270,N_13949,N_14677);
xor U18271 (N_18271,N_12264,N_12193);
and U18272 (N_18272,N_15999,N_15841);
or U18273 (N_18273,N_14812,N_14263);
and U18274 (N_18274,N_14940,N_14408);
and U18275 (N_18275,N_13604,N_13968);
or U18276 (N_18276,N_15250,N_12552);
nor U18277 (N_18277,N_15641,N_15989);
nand U18278 (N_18278,N_13960,N_12295);
and U18279 (N_18279,N_12302,N_13907);
xnor U18280 (N_18280,N_15954,N_13694);
and U18281 (N_18281,N_15478,N_12897);
xnor U18282 (N_18282,N_13364,N_13045);
nand U18283 (N_18283,N_12686,N_14318);
xor U18284 (N_18284,N_14962,N_12283);
xor U18285 (N_18285,N_12788,N_13011);
and U18286 (N_18286,N_13153,N_12776);
or U18287 (N_18287,N_15667,N_15297);
and U18288 (N_18288,N_12237,N_12424);
or U18289 (N_18289,N_13457,N_15088);
or U18290 (N_18290,N_12563,N_15002);
and U18291 (N_18291,N_15648,N_14174);
nand U18292 (N_18292,N_15096,N_13396);
nand U18293 (N_18293,N_12635,N_15985);
nor U18294 (N_18294,N_12388,N_13373);
xor U18295 (N_18295,N_12612,N_12827);
nand U18296 (N_18296,N_14696,N_12674);
and U18297 (N_18297,N_12341,N_15752);
and U18298 (N_18298,N_15731,N_15855);
nand U18299 (N_18299,N_15658,N_15077);
nor U18300 (N_18300,N_12778,N_14702);
xor U18301 (N_18301,N_15923,N_15507);
and U18302 (N_18302,N_13052,N_12808);
or U18303 (N_18303,N_14921,N_14485);
nor U18304 (N_18304,N_12316,N_13059);
or U18305 (N_18305,N_12566,N_12549);
nor U18306 (N_18306,N_12349,N_14015);
nor U18307 (N_18307,N_13168,N_13051);
xnor U18308 (N_18308,N_13705,N_15289);
nor U18309 (N_18309,N_14583,N_13786);
nand U18310 (N_18310,N_14442,N_15835);
or U18311 (N_18311,N_14882,N_12788);
or U18312 (N_18312,N_13878,N_14801);
nand U18313 (N_18313,N_13683,N_15667);
and U18314 (N_18314,N_12560,N_15257);
and U18315 (N_18315,N_12024,N_12069);
nand U18316 (N_18316,N_12462,N_15470);
nand U18317 (N_18317,N_14152,N_15605);
xnor U18318 (N_18318,N_14570,N_15412);
and U18319 (N_18319,N_12899,N_14263);
nand U18320 (N_18320,N_15682,N_13773);
nor U18321 (N_18321,N_12843,N_12606);
and U18322 (N_18322,N_15567,N_15354);
nor U18323 (N_18323,N_14170,N_15078);
and U18324 (N_18324,N_15807,N_15752);
nand U18325 (N_18325,N_15871,N_14782);
nor U18326 (N_18326,N_12378,N_13190);
or U18327 (N_18327,N_14015,N_13380);
nand U18328 (N_18328,N_14141,N_14018);
xnor U18329 (N_18329,N_15233,N_14338);
nand U18330 (N_18330,N_14968,N_15578);
nand U18331 (N_18331,N_13493,N_13993);
nand U18332 (N_18332,N_15672,N_14117);
nor U18333 (N_18333,N_12315,N_13049);
xor U18334 (N_18334,N_15125,N_15284);
and U18335 (N_18335,N_13591,N_15593);
and U18336 (N_18336,N_14820,N_12180);
nand U18337 (N_18337,N_15301,N_14219);
or U18338 (N_18338,N_15183,N_12083);
or U18339 (N_18339,N_13154,N_15899);
nand U18340 (N_18340,N_13716,N_15325);
nor U18341 (N_18341,N_14980,N_14348);
or U18342 (N_18342,N_12451,N_13074);
or U18343 (N_18343,N_14523,N_14005);
xor U18344 (N_18344,N_12029,N_15709);
or U18345 (N_18345,N_14123,N_12613);
and U18346 (N_18346,N_13234,N_13284);
nor U18347 (N_18347,N_12553,N_14950);
nor U18348 (N_18348,N_13989,N_13415);
nand U18349 (N_18349,N_12532,N_15571);
and U18350 (N_18350,N_14986,N_12067);
nor U18351 (N_18351,N_12610,N_14921);
nand U18352 (N_18352,N_15449,N_14223);
xor U18353 (N_18353,N_13457,N_13866);
nand U18354 (N_18354,N_13956,N_15573);
nand U18355 (N_18355,N_14699,N_13670);
nor U18356 (N_18356,N_12359,N_15752);
nor U18357 (N_18357,N_14199,N_15424);
or U18358 (N_18358,N_13010,N_15726);
nand U18359 (N_18359,N_13254,N_14332);
nor U18360 (N_18360,N_15352,N_15178);
nor U18361 (N_18361,N_15695,N_15944);
nor U18362 (N_18362,N_13588,N_14948);
or U18363 (N_18363,N_13777,N_13229);
and U18364 (N_18364,N_15072,N_14746);
or U18365 (N_18365,N_14120,N_12603);
and U18366 (N_18366,N_14236,N_13619);
xor U18367 (N_18367,N_12469,N_14271);
nand U18368 (N_18368,N_15888,N_12910);
or U18369 (N_18369,N_15746,N_15611);
and U18370 (N_18370,N_12276,N_12843);
and U18371 (N_18371,N_13397,N_13965);
or U18372 (N_18372,N_13597,N_15836);
or U18373 (N_18373,N_14075,N_15322);
nor U18374 (N_18374,N_13383,N_13595);
xor U18375 (N_18375,N_15374,N_14151);
and U18376 (N_18376,N_13722,N_12601);
or U18377 (N_18377,N_14029,N_12506);
nand U18378 (N_18378,N_13553,N_12699);
nor U18379 (N_18379,N_15238,N_14563);
and U18380 (N_18380,N_15366,N_12847);
nor U18381 (N_18381,N_14475,N_12475);
or U18382 (N_18382,N_12748,N_12227);
or U18383 (N_18383,N_15740,N_12118);
nand U18384 (N_18384,N_13738,N_14790);
nor U18385 (N_18385,N_14016,N_15174);
and U18386 (N_18386,N_12683,N_12396);
or U18387 (N_18387,N_13390,N_14197);
and U18388 (N_18388,N_13450,N_14673);
and U18389 (N_18389,N_14142,N_15599);
or U18390 (N_18390,N_15801,N_12806);
or U18391 (N_18391,N_14876,N_15116);
nand U18392 (N_18392,N_12391,N_14700);
nor U18393 (N_18393,N_13333,N_13941);
nand U18394 (N_18394,N_13903,N_12411);
or U18395 (N_18395,N_12982,N_14048);
and U18396 (N_18396,N_15308,N_15604);
and U18397 (N_18397,N_12409,N_12052);
and U18398 (N_18398,N_15275,N_13494);
nand U18399 (N_18399,N_15884,N_13221);
nor U18400 (N_18400,N_13772,N_13393);
or U18401 (N_18401,N_12253,N_15670);
and U18402 (N_18402,N_15688,N_14541);
nand U18403 (N_18403,N_15655,N_13885);
xnor U18404 (N_18404,N_12278,N_12895);
nand U18405 (N_18405,N_15151,N_15070);
and U18406 (N_18406,N_14442,N_14561);
or U18407 (N_18407,N_14746,N_15754);
xor U18408 (N_18408,N_15741,N_14211);
or U18409 (N_18409,N_15918,N_12856);
or U18410 (N_18410,N_14746,N_12524);
and U18411 (N_18411,N_12372,N_13708);
nand U18412 (N_18412,N_14597,N_14679);
nor U18413 (N_18413,N_12190,N_14585);
nand U18414 (N_18414,N_12196,N_13336);
and U18415 (N_18415,N_15595,N_12398);
and U18416 (N_18416,N_13630,N_12974);
xnor U18417 (N_18417,N_12669,N_15227);
nand U18418 (N_18418,N_12424,N_13961);
and U18419 (N_18419,N_13690,N_12982);
nand U18420 (N_18420,N_14951,N_14430);
nand U18421 (N_18421,N_13607,N_15983);
xor U18422 (N_18422,N_13090,N_15835);
or U18423 (N_18423,N_13685,N_15527);
nor U18424 (N_18424,N_12440,N_13579);
and U18425 (N_18425,N_12900,N_15577);
nor U18426 (N_18426,N_14189,N_15758);
nor U18427 (N_18427,N_15244,N_15349);
or U18428 (N_18428,N_15269,N_13136);
nor U18429 (N_18429,N_13409,N_12637);
xnor U18430 (N_18430,N_12554,N_15315);
or U18431 (N_18431,N_15728,N_13919);
and U18432 (N_18432,N_13627,N_13507);
nor U18433 (N_18433,N_15739,N_13525);
nand U18434 (N_18434,N_13127,N_13672);
and U18435 (N_18435,N_12344,N_15562);
nand U18436 (N_18436,N_15559,N_15315);
and U18437 (N_18437,N_12760,N_12854);
xnor U18438 (N_18438,N_13469,N_14223);
nand U18439 (N_18439,N_14972,N_15205);
nor U18440 (N_18440,N_12149,N_15394);
xor U18441 (N_18441,N_15337,N_12684);
nand U18442 (N_18442,N_14154,N_15767);
and U18443 (N_18443,N_13086,N_15585);
and U18444 (N_18444,N_14612,N_15420);
and U18445 (N_18445,N_15151,N_14048);
nand U18446 (N_18446,N_13894,N_13889);
nor U18447 (N_18447,N_12606,N_14035);
nor U18448 (N_18448,N_15958,N_13307);
nor U18449 (N_18449,N_14868,N_14985);
or U18450 (N_18450,N_13840,N_14020);
nor U18451 (N_18451,N_12996,N_13836);
or U18452 (N_18452,N_14100,N_15042);
nor U18453 (N_18453,N_14912,N_14313);
and U18454 (N_18454,N_12828,N_14751);
or U18455 (N_18455,N_14092,N_12058);
and U18456 (N_18456,N_14763,N_14198);
nand U18457 (N_18457,N_14862,N_12459);
nor U18458 (N_18458,N_13536,N_12838);
xor U18459 (N_18459,N_12197,N_14626);
or U18460 (N_18460,N_13290,N_12062);
nand U18461 (N_18461,N_15098,N_14893);
or U18462 (N_18462,N_15700,N_14970);
and U18463 (N_18463,N_14377,N_14785);
xor U18464 (N_18464,N_12031,N_12995);
or U18465 (N_18465,N_14279,N_13156);
nand U18466 (N_18466,N_15545,N_15090);
xnor U18467 (N_18467,N_12101,N_13690);
or U18468 (N_18468,N_15321,N_15393);
and U18469 (N_18469,N_13007,N_15791);
nand U18470 (N_18470,N_13303,N_12053);
and U18471 (N_18471,N_13133,N_14013);
and U18472 (N_18472,N_14495,N_15960);
and U18473 (N_18473,N_13344,N_14802);
nand U18474 (N_18474,N_15006,N_13436);
and U18475 (N_18475,N_15836,N_14173);
xnor U18476 (N_18476,N_15605,N_12802);
and U18477 (N_18477,N_13980,N_14116);
nand U18478 (N_18478,N_12779,N_14447);
nor U18479 (N_18479,N_12307,N_15809);
nor U18480 (N_18480,N_15071,N_14546);
or U18481 (N_18481,N_12830,N_12578);
nor U18482 (N_18482,N_12912,N_14336);
or U18483 (N_18483,N_15427,N_13055);
nor U18484 (N_18484,N_15938,N_15678);
and U18485 (N_18485,N_12405,N_12383);
nor U18486 (N_18486,N_15792,N_15442);
or U18487 (N_18487,N_15863,N_13954);
nor U18488 (N_18488,N_14873,N_14877);
or U18489 (N_18489,N_12547,N_14544);
nand U18490 (N_18490,N_12725,N_15478);
and U18491 (N_18491,N_14346,N_13709);
xor U18492 (N_18492,N_15611,N_15780);
nor U18493 (N_18493,N_14554,N_13189);
xor U18494 (N_18494,N_12046,N_13346);
and U18495 (N_18495,N_12974,N_15052);
nor U18496 (N_18496,N_12928,N_13138);
and U18497 (N_18497,N_14130,N_12922);
and U18498 (N_18498,N_12773,N_14349);
nor U18499 (N_18499,N_14118,N_15245);
xor U18500 (N_18500,N_14116,N_12046);
or U18501 (N_18501,N_12500,N_12192);
or U18502 (N_18502,N_15957,N_14181);
or U18503 (N_18503,N_14749,N_14743);
xor U18504 (N_18504,N_14255,N_14551);
xor U18505 (N_18505,N_15884,N_14192);
or U18506 (N_18506,N_13717,N_13338);
or U18507 (N_18507,N_14731,N_12340);
nor U18508 (N_18508,N_13027,N_15316);
and U18509 (N_18509,N_12115,N_13086);
nand U18510 (N_18510,N_13477,N_13163);
nand U18511 (N_18511,N_14567,N_13822);
xnor U18512 (N_18512,N_15532,N_14962);
nor U18513 (N_18513,N_14574,N_12511);
nor U18514 (N_18514,N_14543,N_14558);
and U18515 (N_18515,N_14034,N_15263);
nor U18516 (N_18516,N_12437,N_14330);
or U18517 (N_18517,N_14343,N_14358);
or U18518 (N_18518,N_15777,N_14490);
nand U18519 (N_18519,N_12280,N_13285);
and U18520 (N_18520,N_12832,N_14147);
or U18521 (N_18521,N_15274,N_12837);
nand U18522 (N_18522,N_15991,N_15564);
nor U18523 (N_18523,N_12077,N_13592);
or U18524 (N_18524,N_13543,N_12875);
nand U18525 (N_18525,N_12870,N_12315);
or U18526 (N_18526,N_14260,N_12898);
nor U18527 (N_18527,N_12294,N_12613);
nor U18528 (N_18528,N_12973,N_14828);
xnor U18529 (N_18529,N_15894,N_13593);
xor U18530 (N_18530,N_13290,N_14369);
nor U18531 (N_18531,N_12213,N_14813);
nor U18532 (N_18532,N_12250,N_13452);
or U18533 (N_18533,N_13387,N_12404);
or U18534 (N_18534,N_12518,N_12491);
nor U18535 (N_18535,N_15742,N_13800);
nand U18536 (N_18536,N_13802,N_15696);
or U18537 (N_18537,N_13252,N_13559);
nor U18538 (N_18538,N_15466,N_14438);
or U18539 (N_18539,N_12190,N_12626);
xor U18540 (N_18540,N_14993,N_15367);
and U18541 (N_18541,N_13162,N_13695);
xnor U18542 (N_18542,N_15711,N_14303);
or U18543 (N_18543,N_14543,N_14764);
and U18544 (N_18544,N_15263,N_15189);
nor U18545 (N_18545,N_12311,N_12371);
nor U18546 (N_18546,N_14739,N_14138);
and U18547 (N_18547,N_15286,N_12502);
and U18548 (N_18548,N_14026,N_13037);
nand U18549 (N_18549,N_12454,N_14064);
nor U18550 (N_18550,N_12694,N_13780);
and U18551 (N_18551,N_13946,N_13925);
nand U18552 (N_18552,N_12954,N_15683);
nand U18553 (N_18553,N_14934,N_15324);
nor U18554 (N_18554,N_14832,N_13482);
nor U18555 (N_18555,N_14852,N_14045);
and U18556 (N_18556,N_12215,N_15454);
nor U18557 (N_18557,N_15359,N_13441);
or U18558 (N_18558,N_12109,N_15894);
nor U18559 (N_18559,N_14246,N_14807);
nor U18560 (N_18560,N_12800,N_14774);
or U18561 (N_18561,N_14477,N_15081);
and U18562 (N_18562,N_13557,N_15215);
or U18563 (N_18563,N_15148,N_14845);
xnor U18564 (N_18564,N_12742,N_13274);
or U18565 (N_18565,N_15219,N_14684);
and U18566 (N_18566,N_12485,N_14102);
or U18567 (N_18567,N_14905,N_14390);
nor U18568 (N_18568,N_12909,N_14439);
nor U18569 (N_18569,N_15476,N_13940);
and U18570 (N_18570,N_12322,N_15211);
or U18571 (N_18571,N_14417,N_14728);
nor U18572 (N_18572,N_12270,N_12506);
nand U18573 (N_18573,N_14107,N_13949);
and U18574 (N_18574,N_15117,N_14020);
nor U18575 (N_18575,N_15754,N_12793);
nand U18576 (N_18576,N_14333,N_13392);
nor U18577 (N_18577,N_12496,N_14600);
and U18578 (N_18578,N_15717,N_12889);
nand U18579 (N_18579,N_14870,N_15487);
or U18580 (N_18580,N_12288,N_12591);
nand U18581 (N_18581,N_15530,N_14737);
nand U18582 (N_18582,N_14996,N_14529);
and U18583 (N_18583,N_12454,N_15549);
or U18584 (N_18584,N_12662,N_13098);
and U18585 (N_18585,N_12777,N_14238);
or U18586 (N_18586,N_15392,N_13545);
nor U18587 (N_18587,N_12861,N_15731);
nor U18588 (N_18588,N_15229,N_12480);
nor U18589 (N_18589,N_14633,N_13666);
xnor U18590 (N_18590,N_14140,N_12101);
and U18591 (N_18591,N_14896,N_12864);
and U18592 (N_18592,N_13089,N_13052);
nor U18593 (N_18593,N_15782,N_14630);
nor U18594 (N_18594,N_12741,N_12872);
and U18595 (N_18595,N_12313,N_15140);
and U18596 (N_18596,N_14000,N_12449);
and U18597 (N_18597,N_15456,N_12632);
nand U18598 (N_18598,N_12674,N_13757);
or U18599 (N_18599,N_13116,N_15092);
or U18600 (N_18600,N_13278,N_13440);
nor U18601 (N_18601,N_15531,N_15282);
xnor U18602 (N_18602,N_12290,N_14542);
nand U18603 (N_18603,N_12083,N_14222);
nor U18604 (N_18604,N_15500,N_15185);
nor U18605 (N_18605,N_15348,N_12267);
xor U18606 (N_18606,N_12288,N_12961);
nor U18607 (N_18607,N_12031,N_13328);
nand U18608 (N_18608,N_12871,N_15366);
nand U18609 (N_18609,N_12275,N_13004);
nor U18610 (N_18610,N_12915,N_15353);
or U18611 (N_18611,N_14345,N_12220);
and U18612 (N_18612,N_15738,N_14464);
nand U18613 (N_18613,N_15081,N_14907);
or U18614 (N_18614,N_13992,N_14998);
nor U18615 (N_18615,N_12337,N_14490);
and U18616 (N_18616,N_12510,N_14593);
nand U18617 (N_18617,N_14305,N_14396);
and U18618 (N_18618,N_14200,N_13619);
and U18619 (N_18619,N_15464,N_13016);
nor U18620 (N_18620,N_13273,N_14016);
xor U18621 (N_18621,N_14431,N_14238);
xnor U18622 (N_18622,N_15033,N_12681);
nand U18623 (N_18623,N_14410,N_15037);
and U18624 (N_18624,N_13278,N_13280);
nand U18625 (N_18625,N_15707,N_13552);
nor U18626 (N_18626,N_14268,N_12652);
and U18627 (N_18627,N_12044,N_14474);
and U18628 (N_18628,N_14952,N_14618);
nor U18629 (N_18629,N_13846,N_13801);
or U18630 (N_18630,N_14025,N_15188);
nor U18631 (N_18631,N_14746,N_13737);
nand U18632 (N_18632,N_13371,N_13057);
nand U18633 (N_18633,N_15656,N_13193);
and U18634 (N_18634,N_13041,N_13795);
nor U18635 (N_18635,N_15684,N_12998);
nor U18636 (N_18636,N_15272,N_15768);
nor U18637 (N_18637,N_14864,N_15376);
and U18638 (N_18638,N_12768,N_13108);
nand U18639 (N_18639,N_15784,N_12008);
and U18640 (N_18640,N_13378,N_14930);
and U18641 (N_18641,N_13832,N_12095);
and U18642 (N_18642,N_12277,N_14343);
nor U18643 (N_18643,N_12765,N_15423);
and U18644 (N_18644,N_15785,N_13429);
nor U18645 (N_18645,N_13553,N_14691);
xor U18646 (N_18646,N_13127,N_13026);
or U18647 (N_18647,N_14498,N_14567);
nor U18648 (N_18648,N_12202,N_14387);
nor U18649 (N_18649,N_13110,N_15360);
and U18650 (N_18650,N_13320,N_14479);
nand U18651 (N_18651,N_12918,N_14457);
nor U18652 (N_18652,N_14692,N_13874);
nor U18653 (N_18653,N_12146,N_14931);
or U18654 (N_18654,N_15903,N_14741);
and U18655 (N_18655,N_12176,N_12806);
nand U18656 (N_18656,N_12101,N_12745);
and U18657 (N_18657,N_13091,N_15958);
or U18658 (N_18658,N_14941,N_14437);
xnor U18659 (N_18659,N_14158,N_12567);
nor U18660 (N_18660,N_13794,N_15405);
or U18661 (N_18661,N_15108,N_14672);
nor U18662 (N_18662,N_13806,N_13556);
nand U18663 (N_18663,N_15638,N_12118);
nor U18664 (N_18664,N_12282,N_15936);
or U18665 (N_18665,N_13498,N_15967);
or U18666 (N_18666,N_13699,N_13483);
and U18667 (N_18667,N_15924,N_15444);
and U18668 (N_18668,N_14476,N_14472);
and U18669 (N_18669,N_12578,N_12122);
nor U18670 (N_18670,N_15008,N_13665);
nor U18671 (N_18671,N_13286,N_15202);
nor U18672 (N_18672,N_14244,N_14230);
and U18673 (N_18673,N_15213,N_15369);
xnor U18674 (N_18674,N_14972,N_12464);
or U18675 (N_18675,N_12484,N_14970);
and U18676 (N_18676,N_15488,N_13017);
xnor U18677 (N_18677,N_14171,N_14510);
nand U18678 (N_18678,N_12030,N_15736);
nand U18679 (N_18679,N_15729,N_15030);
and U18680 (N_18680,N_12938,N_14578);
nand U18681 (N_18681,N_12223,N_13113);
xor U18682 (N_18682,N_14699,N_14865);
nor U18683 (N_18683,N_12377,N_13929);
or U18684 (N_18684,N_12416,N_15337);
nor U18685 (N_18685,N_15867,N_14208);
nand U18686 (N_18686,N_14412,N_13486);
or U18687 (N_18687,N_14063,N_14697);
or U18688 (N_18688,N_14892,N_13025);
nor U18689 (N_18689,N_15849,N_14197);
nand U18690 (N_18690,N_15969,N_14384);
xnor U18691 (N_18691,N_13792,N_13264);
nand U18692 (N_18692,N_14478,N_15534);
and U18693 (N_18693,N_14679,N_15112);
nor U18694 (N_18694,N_12153,N_13805);
or U18695 (N_18695,N_12502,N_15572);
or U18696 (N_18696,N_12878,N_14216);
or U18697 (N_18697,N_12413,N_13466);
nor U18698 (N_18698,N_13550,N_12175);
nor U18699 (N_18699,N_13374,N_12427);
nand U18700 (N_18700,N_15391,N_14004);
and U18701 (N_18701,N_15125,N_14545);
nor U18702 (N_18702,N_12882,N_15115);
or U18703 (N_18703,N_15892,N_12494);
or U18704 (N_18704,N_15230,N_13080);
nand U18705 (N_18705,N_12637,N_15300);
or U18706 (N_18706,N_15534,N_13912);
nand U18707 (N_18707,N_14980,N_15796);
nand U18708 (N_18708,N_15500,N_14411);
nor U18709 (N_18709,N_13161,N_13295);
nand U18710 (N_18710,N_12478,N_12744);
nor U18711 (N_18711,N_15729,N_14123);
or U18712 (N_18712,N_14518,N_12810);
nor U18713 (N_18713,N_14999,N_14884);
nor U18714 (N_18714,N_13017,N_12284);
nor U18715 (N_18715,N_13376,N_12248);
nor U18716 (N_18716,N_14301,N_13335);
or U18717 (N_18717,N_14238,N_15145);
and U18718 (N_18718,N_15787,N_13939);
nand U18719 (N_18719,N_13906,N_15553);
and U18720 (N_18720,N_12661,N_14742);
nor U18721 (N_18721,N_13470,N_12498);
and U18722 (N_18722,N_12772,N_12283);
nor U18723 (N_18723,N_12868,N_13372);
and U18724 (N_18724,N_13797,N_14597);
nor U18725 (N_18725,N_12080,N_13306);
and U18726 (N_18726,N_12643,N_14139);
nor U18727 (N_18727,N_14992,N_12083);
nor U18728 (N_18728,N_14021,N_12732);
and U18729 (N_18729,N_14347,N_13617);
and U18730 (N_18730,N_12911,N_15467);
and U18731 (N_18731,N_12379,N_12573);
and U18732 (N_18732,N_14065,N_12221);
and U18733 (N_18733,N_15599,N_14751);
and U18734 (N_18734,N_13682,N_14238);
or U18735 (N_18735,N_12611,N_14085);
and U18736 (N_18736,N_14942,N_13252);
nor U18737 (N_18737,N_12387,N_15127);
or U18738 (N_18738,N_13524,N_14494);
nand U18739 (N_18739,N_15650,N_13500);
and U18740 (N_18740,N_12849,N_13654);
or U18741 (N_18741,N_15230,N_15750);
and U18742 (N_18742,N_13008,N_13730);
nor U18743 (N_18743,N_14605,N_15366);
nand U18744 (N_18744,N_12492,N_15671);
xor U18745 (N_18745,N_14869,N_12528);
xor U18746 (N_18746,N_12965,N_15707);
or U18747 (N_18747,N_13466,N_14678);
nor U18748 (N_18748,N_13633,N_14537);
and U18749 (N_18749,N_13535,N_15395);
xor U18750 (N_18750,N_14551,N_12036);
nand U18751 (N_18751,N_12287,N_15358);
and U18752 (N_18752,N_13816,N_12905);
nand U18753 (N_18753,N_12401,N_13058);
nand U18754 (N_18754,N_13267,N_15586);
xor U18755 (N_18755,N_14615,N_12336);
nand U18756 (N_18756,N_12255,N_14601);
nor U18757 (N_18757,N_12190,N_15494);
or U18758 (N_18758,N_12022,N_13124);
and U18759 (N_18759,N_15241,N_15294);
or U18760 (N_18760,N_12013,N_15675);
nand U18761 (N_18761,N_15781,N_14154);
and U18762 (N_18762,N_13569,N_14146);
or U18763 (N_18763,N_12636,N_12109);
or U18764 (N_18764,N_15173,N_12479);
and U18765 (N_18765,N_13230,N_15494);
and U18766 (N_18766,N_15776,N_15421);
or U18767 (N_18767,N_13661,N_13038);
nor U18768 (N_18768,N_14301,N_13648);
or U18769 (N_18769,N_14961,N_15835);
xor U18770 (N_18770,N_15796,N_14344);
nand U18771 (N_18771,N_15061,N_13052);
or U18772 (N_18772,N_15628,N_12236);
nor U18773 (N_18773,N_14465,N_12886);
xor U18774 (N_18774,N_13257,N_14812);
and U18775 (N_18775,N_15211,N_15078);
xnor U18776 (N_18776,N_14167,N_14864);
nand U18777 (N_18777,N_14091,N_12491);
nor U18778 (N_18778,N_14811,N_12684);
nand U18779 (N_18779,N_14517,N_15780);
nand U18780 (N_18780,N_15880,N_12410);
nand U18781 (N_18781,N_14412,N_14670);
nand U18782 (N_18782,N_12237,N_14272);
or U18783 (N_18783,N_13906,N_13729);
nor U18784 (N_18784,N_12393,N_13090);
nand U18785 (N_18785,N_12636,N_13489);
nor U18786 (N_18786,N_14149,N_14425);
nor U18787 (N_18787,N_14975,N_14854);
or U18788 (N_18788,N_14627,N_15449);
nor U18789 (N_18789,N_12853,N_15353);
xor U18790 (N_18790,N_14897,N_15663);
or U18791 (N_18791,N_12202,N_14980);
nor U18792 (N_18792,N_14661,N_13042);
and U18793 (N_18793,N_15869,N_12538);
nand U18794 (N_18794,N_15915,N_13747);
and U18795 (N_18795,N_15378,N_14906);
or U18796 (N_18796,N_12546,N_13738);
xor U18797 (N_18797,N_14411,N_12973);
nand U18798 (N_18798,N_12363,N_15624);
nor U18799 (N_18799,N_12613,N_15303);
nor U18800 (N_18800,N_14847,N_14853);
and U18801 (N_18801,N_15046,N_12161);
nor U18802 (N_18802,N_14190,N_14562);
or U18803 (N_18803,N_14444,N_13223);
and U18804 (N_18804,N_12786,N_14770);
nor U18805 (N_18805,N_14326,N_15864);
nor U18806 (N_18806,N_12601,N_15521);
and U18807 (N_18807,N_12532,N_15607);
nor U18808 (N_18808,N_13898,N_15060);
nand U18809 (N_18809,N_12145,N_13066);
xor U18810 (N_18810,N_12066,N_14530);
nand U18811 (N_18811,N_12588,N_14605);
nor U18812 (N_18812,N_14967,N_14438);
or U18813 (N_18813,N_14890,N_14447);
xor U18814 (N_18814,N_13453,N_13930);
or U18815 (N_18815,N_12211,N_15698);
and U18816 (N_18816,N_13989,N_12735);
nand U18817 (N_18817,N_14661,N_15130);
nand U18818 (N_18818,N_14474,N_15075);
nor U18819 (N_18819,N_15138,N_13418);
nor U18820 (N_18820,N_14713,N_14423);
and U18821 (N_18821,N_14753,N_14047);
nor U18822 (N_18822,N_13202,N_13693);
xnor U18823 (N_18823,N_13025,N_15470);
nor U18824 (N_18824,N_13935,N_13448);
xnor U18825 (N_18825,N_15862,N_14632);
or U18826 (N_18826,N_15466,N_12683);
or U18827 (N_18827,N_15216,N_14544);
nand U18828 (N_18828,N_15455,N_14725);
nand U18829 (N_18829,N_12538,N_14591);
nor U18830 (N_18830,N_15544,N_13395);
nand U18831 (N_18831,N_15591,N_13198);
xor U18832 (N_18832,N_12573,N_15429);
nor U18833 (N_18833,N_13577,N_15251);
or U18834 (N_18834,N_15586,N_13234);
nor U18835 (N_18835,N_13024,N_12195);
and U18836 (N_18836,N_13108,N_12060);
nor U18837 (N_18837,N_14813,N_15653);
nor U18838 (N_18838,N_13787,N_13488);
or U18839 (N_18839,N_12816,N_15918);
nand U18840 (N_18840,N_13492,N_15826);
xor U18841 (N_18841,N_12500,N_15444);
nand U18842 (N_18842,N_15399,N_14042);
and U18843 (N_18843,N_14641,N_13677);
nor U18844 (N_18844,N_14616,N_14534);
nand U18845 (N_18845,N_12529,N_14562);
or U18846 (N_18846,N_12650,N_13487);
xor U18847 (N_18847,N_15516,N_15008);
nand U18848 (N_18848,N_15194,N_14731);
and U18849 (N_18849,N_12502,N_13620);
or U18850 (N_18850,N_15630,N_12688);
and U18851 (N_18851,N_14040,N_15896);
nor U18852 (N_18852,N_13213,N_13667);
or U18853 (N_18853,N_13735,N_13338);
or U18854 (N_18854,N_15631,N_14313);
nor U18855 (N_18855,N_14375,N_14974);
nand U18856 (N_18856,N_12877,N_13676);
nor U18857 (N_18857,N_15141,N_13873);
or U18858 (N_18858,N_15574,N_15713);
or U18859 (N_18859,N_12005,N_14697);
and U18860 (N_18860,N_13924,N_13537);
nand U18861 (N_18861,N_14696,N_14426);
xnor U18862 (N_18862,N_14559,N_12349);
nand U18863 (N_18863,N_14556,N_15389);
and U18864 (N_18864,N_12899,N_15694);
nand U18865 (N_18865,N_15809,N_13972);
or U18866 (N_18866,N_12763,N_15404);
nor U18867 (N_18867,N_12618,N_15638);
nor U18868 (N_18868,N_13108,N_13111);
nor U18869 (N_18869,N_14390,N_12530);
or U18870 (N_18870,N_12055,N_15128);
nand U18871 (N_18871,N_15766,N_15485);
and U18872 (N_18872,N_15348,N_14677);
and U18873 (N_18873,N_15253,N_14634);
nor U18874 (N_18874,N_15485,N_13669);
xnor U18875 (N_18875,N_14857,N_12062);
or U18876 (N_18876,N_13645,N_14275);
and U18877 (N_18877,N_15005,N_13409);
nand U18878 (N_18878,N_13556,N_15332);
or U18879 (N_18879,N_13951,N_13887);
and U18880 (N_18880,N_15321,N_13541);
nand U18881 (N_18881,N_14049,N_15346);
or U18882 (N_18882,N_14478,N_12703);
and U18883 (N_18883,N_12394,N_12090);
nand U18884 (N_18884,N_15691,N_15052);
or U18885 (N_18885,N_15981,N_14626);
or U18886 (N_18886,N_13267,N_14226);
nand U18887 (N_18887,N_13408,N_15097);
nor U18888 (N_18888,N_13042,N_14337);
or U18889 (N_18889,N_14552,N_12625);
or U18890 (N_18890,N_12245,N_12313);
and U18891 (N_18891,N_13358,N_13726);
nand U18892 (N_18892,N_15334,N_15347);
and U18893 (N_18893,N_12218,N_14955);
nor U18894 (N_18894,N_14687,N_12141);
nor U18895 (N_18895,N_14506,N_13616);
xnor U18896 (N_18896,N_14592,N_14808);
nor U18897 (N_18897,N_15729,N_13373);
nor U18898 (N_18898,N_12628,N_15667);
or U18899 (N_18899,N_13833,N_13291);
and U18900 (N_18900,N_14692,N_12207);
nor U18901 (N_18901,N_15109,N_12387);
xnor U18902 (N_18902,N_15783,N_15861);
and U18903 (N_18903,N_12489,N_15765);
nand U18904 (N_18904,N_14427,N_12740);
nor U18905 (N_18905,N_15453,N_13835);
or U18906 (N_18906,N_15232,N_14969);
or U18907 (N_18907,N_12824,N_13500);
nand U18908 (N_18908,N_12303,N_12926);
xnor U18909 (N_18909,N_12155,N_15312);
or U18910 (N_18910,N_15780,N_14793);
and U18911 (N_18911,N_14503,N_14657);
nor U18912 (N_18912,N_15568,N_15175);
nor U18913 (N_18913,N_15027,N_13508);
nand U18914 (N_18914,N_14476,N_13365);
or U18915 (N_18915,N_14142,N_13063);
or U18916 (N_18916,N_12891,N_13971);
xor U18917 (N_18917,N_12214,N_12280);
nand U18918 (N_18918,N_13207,N_12096);
nand U18919 (N_18919,N_12847,N_14111);
nor U18920 (N_18920,N_14068,N_13651);
or U18921 (N_18921,N_13995,N_13918);
and U18922 (N_18922,N_15402,N_14360);
or U18923 (N_18923,N_15040,N_15599);
nand U18924 (N_18924,N_15059,N_14070);
nand U18925 (N_18925,N_12277,N_12091);
or U18926 (N_18926,N_14455,N_12113);
and U18927 (N_18927,N_15394,N_13127);
nor U18928 (N_18928,N_15699,N_15850);
xnor U18929 (N_18929,N_13442,N_15560);
and U18930 (N_18930,N_13951,N_14635);
or U18931 (N_18931,N_13548,N_15954);
nand U18932 (N_18932,N_12391,N_15931);
nor U18933 (N_18933,N_14953,N_15838);
and U18934 (N_18934,N_13885,N_14517);
and U18935 (N_18935,N_14135,N_15683);
nand U18936 (N_18936,N_14366,N_12528);
nand U18937 (N_18937,N_12366,N_13565);
nand U18938 (N_18938,N_14797,N_12392);
nand U18939 (N_18939,N_12186,N_15226);
nor U18940 (N_18940,N_12042,N_14096);
nor U18941 (N_18941,N_12950,N_14579);
xnor U18942 (N_18942,N_15464,N_14012);
or U18943 (N_18943,N_15852,N_12244);
and U18944 (N_18944,N_13408,N_15443);
nor U18945 (N_18945,N_15899,N_12870);
nand U18946 (N_18946,N_15900,N_12324);
nor U18947 (N_18947,N_12524,N_12866);
or U18948 (N_18948,N_14520,N_13702);
or U18949 (N_18949,N_12820,N_15771);
nand U18950 (N_18950,N_15776,N_14355);
or U18951 (N_18951,N_13735,N_14462);
and U18952 (N_18952,N_15180,N_15508);
and U18953 (N_18953,N_15786,N_13507);
or U18954 (N_18954,N_13256,N_12085);
or U18955 (N_18955,N_12787,N_14554);
nor U18956 (N_18956,N_13192,N_12057);
nor U18957 (N_18957,N_12532,N_14319);
or U18958 (N_18958,N_12116,N_15015);
nor U18959 (N_18959,N_15629,N_14617);
or U18960 (N_18960,N_14011,N_13844);
or U18961 (N_18961,N_15726,N_15220);
xnor U18962 (N_18962,N_12276,N_14509);
nand U18963 (N_18963,N_15098,N_13509);
nor U18964 (N_18964,N_13250,N_13576);
nand U18965 (N_18965,N_12683,N_12576);
and U18966 (N_18966,N_12881,N_14433);
and U18967 (N_18967,N_15125,N_15422);
nand U18968 (N_18968,N_14686,N_15519);
and U18969 (N_18969,N_13156,N_12512);
xnor U18970 (N_18970,N_12207,N_12073);
nor U18971 (N_18971,N_12839,N_13076);
nand U18972 (N_18972,N_13682,N_15672);
nor U18973 (N_18973,N_14866,N_14661);
xnor U18974 (N_18974,N_12591,N_15193);
or U18975 (N_18975,N_12277,N_13534);
nor U18976 (N_18976,N_14417,N_15843);
nand U18977 (N_18977,N_13084,N_15790);
or U18978 (N_18978,N_15191,N_15352);
nand U18979 (N_18979,N_12787,N_15912);
or U18980 (N_18980,N_13850,N_12038);
nand U18981 (N_18981,N_13904,N_15931);
and U18982 (N_18982,N_13015,N_12865);
nand U18983 (N_18983,N_15774,N_12415);
xnor U18984 (N_18984,N_15551,N_14056);
or U18985 (N_18985,N_13571,N_12501);
and U18986 (N_18986,N_13571,N_14961);
nand U18987 (N_18987,N_14211,N_14441);
and U18988 (N_18988,N_12438,N_12296);
and U18989 (N_18989,N_13891,N_12897);
nand U18990 (N_18990,N_12725,N_14631);
and U18991 (N_18991,N_13522,N_13883);
or U18992 (N_18992,N_14624,N_15790);
or U18993 (N_18993,N_15784,N_15172);
nand U18994 (N_18994,N_12843,N_14646);
or U18995 (N_18995,N_12443,N_13687);
xor U18996 (N_18996,N_12778,N_12642);
or U18997 (N_18997,N_14920,N_15073);
nor U18998 (N_18998,N_12795,N_14797);
or U18999 (N_18999,N_13730,N_14598);
nand U19000 (N_19000,N_14275,N_15407);
and U19001 (N_19001,N_15333,N_13289);
and U19002 (N_19002,N_15067,N_13273);
xnor U19003 (N_19003,N_13908,N_12712);
and U19004 (N_19004,N_12629,N_13046);
nor U19005 (N_19005,N_14484,N_14946);
nor U19006 (N_19006,N_15016,N_15435);
nand U19007 (N_19007,N_15915,N_13797);
nand U19008 (N_19008,N_12534,N_15000);
or U19009 (N_19009,N_15671,N_14102);
or U19010 (N_19010,N_13556,N_13548);
nor U19011 (N_19011,N_12684,N_14117);
nor U19012 (N_19012,N_15972,N_12079);
nand U19013 (N_19013,N_12360,N_13172);
or U19014 (N_19014,N_14823,N_12606);
nor U19015 (N_19015,N_13477,N_13385);
or U19016 (N_19016,N_14611,N_13158);
nor U19017 (N_19017,N_13823,N_12032);
nor U19018 (N_19018,N_13661,N_14353);
xnor U19019 (N_19019,N_13147,N_12201);
or U19020 (N_19020,N_13004,N_14862);
nand U19021 (N_19021,N_14481,N_15652);
nor U19022 (N_19022,N_12226,N_14044);
nor U19023 (N_19023,N_14743,N_14847);
nand U19024 (N_19024,N_14003,N_13006);
or U19025 (N_19025,N_14168,N_15325);
or U19026 (N_19026,N_15706,N_13725);
nor U19027 (N_19027,N_15221,N_15860);
nand U19028 (N_19028,N_13640,N_15976);
or U19029 (N_19029,N_13206,N_13285);
or U19030 (N_19030,N_14380,N_15818);
or U19031 (N_19031,N_14791,N_12595);
nand U19032 (N_19032,N_14058,N_13188);
nor U19033 (N_19033,N_14639,N_13326);
nor U19034 (N_19034,N_13036,N_15890);
nand U19035 (N_19035,N_14457,N_12926);
and U19036 (N_19036,N_14252,N_13881);
nand U19037 (N_19037,N_14605,N_13231);
and U19038 (N_19038,N_15936,N_13640);
xor U19039 (N_19039,N_15350,N_13969);
nor U19040 (N_19040,N_12355,N_14090);
and U19041 (N_19041,N_12000,N_14063);
and U19042 (N_19042,N_15622,N_12566);
nor U19043 (N_19043,N_14299,N_13054);
and U19044 (N_19044,N_12704,N_15512);
nand U19045 (N_19045,N_13215,N_14801);
nor U19046 (N_19046,N_12725,N_15281);
xnor U19047 (N_19047,N_12555,N_13944);
nor U19048 (N_19048,N_12288,N_14706);
xnor U19049 (N_19049,N_14318,N_15117);
and U19050 (N_19050,N_12216,N_13452);
or U19051 (N_19051,N_13374,N_12603);
or U19052 (N_19052,N_12576,N_12454);
nor U19053 (N_19053,N_12696,N_12207);
nand U19054 (N_19054,N_13109,N_15953);
nor U19055 (N_19055,N_13170,N_14433);
or U19056 (N_19056,N_12657,N_14805);
xnor U19057 (N_19057,N_13226,N_14967);
nor U19058 (N_19058,N_12137,N_14859);
nor U19059 (N_19059,N_12405,N_12801);
or U19060 (N_19060,N_14508,N_14511);
or U19061 (N_19061,N_13913,N_14994);
xor U19062 (N_19062,N_14424,N_15185);
nor U19063 (N_19063,N_12357,N_13263);
or U19064 (N_19064,N_14282,N_15407);
or U19065 (N_19065,N_15584,N_14352);
nand U19066 (N_19066,N_14602,N_12287);
xor U19067 (N_19067,N_14766,N_12537);
xnor U19068 (N_19068,N_13328,N_14840);
and U19069 (N_19069,N_15728,N_14686);
nor U19070 (N_19070,N_12053,N_12168);
and U19071 (N_19071,N_15827,N_14511);
and U19072 (N_19072,N_12026,N_12424);
or U19073 (N_19073,N_12164,N_13209);
nand U19074 (N_19074,N_14098,N_12325);
and U19075 (N_19075,N_13958,N_12433);
nand U19076 (N_19076,N_14579,N_13446);
and U19077 (N_19077,N_14436,N_13607);
nor U19078 (N_19078,N_13600,N_14245);
and U19079 (N_19079,N_13256,N_15737);
nand U19080 (N_19080,N_15592,N_12861);
or U19081 (N_19081,N_12735,N_14608);
nand U19082 (N_19082,N_12604,N_14407);
and U19083 (N_19083,N_15417,N_13503);
nand U19084 (N_19084,N_12368,N_13503);
nand U19085 (N_19085,N_12258,N_14983);
and U19086 (N_19086,N_14750,N_12447);
nor U19087 (N_19087,N_13852,N_13544);
nand U19088 (N_19088,N_14560,N_12983);
and U19089 (N_19089,N_14784,N_12114);
or U19090 (N_19090,N_14361,N_13940);
nand U19091 (N_19091,N_14330,N_13101);
nand U19092 (N_19092,N_12958,N_13388);
nand U19093 (N_19093,N_14336,N_13727);
and U19094 (N_19094,N_15877,N_12018);
or U19095 (N_19095,N_13820,N_12226);
nor U19096 (N_19096,N_14480,N_13100);
nand U19097 (N_19097,N_13002,N_15049);
nor U19098 (N_19098,N_13382,N_12291);
and U19099 (N_19099,N_12500,N_13959);
and U19100 (N_19100,N_14587,N_15198);
nor U19101 (N_19101,N_15826,N_14893);
nand U19102 (N_19102,N_13236,N_12519);
or U19103 (N_19103,N_15684,N_13495);
and U19104 (N_19104,N_12845,N_13751);
or U19105 (N_19105,N_12514,N_13688);
xnor U19106 (N_19106,N_12146,N_13823);
nand U19107 (N_19107,N_15134,N_14080);
and U19108 (N_19108,N_12098,N_12642);
nor U19109 (N_19109,N_12973,N_15401);
or U19110 (N_19110,N_12306,N_14084);
nor U19111 (N_19111,N_14862,N_15461);
or U19112 (N_19112,N_15129,N_15242);
or U19113 (N_19113,N_12323,N_14494);
nor U19114 (N_19114,N_13189,N_12674);
or U19115 (N_19115,N_12950,N_15361);
nor U19116 (N_19116,N_14465,N_14463);
nor U19117 (N_19117,N_13309,N_14942);
nand U19118 (N_19118,N_12771,N_15253);
or U19119 (N_19119,N_13312,N_14751);
nor U19120 (N_19120,N_14253,N_12474);
nor U19121 (N_19121,N_15814,N_15848);
xnor U19122 (N_19122,N_12857,N_13516);
and U19123 (N_19123,N_12546,N_13560);
nand U19124 (N_19124,N_12530,N_14997);
and U19125 (N_19125,N_15098,N_15288);
nand U19126 (N_19126,N_13454,N_13311);
or U19127 (N_19127,N_13468,N_12054);
or U19128 (N_19128,N_14897,N_13587);
nor U19129 (N_19129,N_14871,N_12588);
and U19130 (N_19130,N_13386,N_15796);
and U19131 (N_19131,N_14731,N_15705);
nor U19132 (N_19132,N_15984,N_12701);
or U19133 (N_19133,N_15734,N_15336);
or U19134 (N_19134,N_12033,N_13080);
and U19135 (N_19135,N_14156,N_12504);
or U19136 (N_19136,N_13155,N_13615);
nand U19137 (N_19137,N_14871,N_13226);
or U19138 (N_19138,N_15471,N_15918);
nand U19139 (N_19139,N_12433,N_12427);
xor U19140 (N_19140,N_15575,N_14118);
xnor U19141 (N_19141,N_13821,N_14318);
nor U19142 (N_19142,N_15188,N_13871);
and U19143 (N_19143,N_13042,N_12424);
nand U19144 (N_19144,N_14868,N_13848);
or U19145 (N_19145,N_13063,N_15301);
nor U19146 (N_19146,N_14530,N_15626);
nand U19147 (N_19147,N_13022,N_13124);
nand U19148 (N_19148,N_15534,N_12340);
xor U19149 (N_19149,N_15137,N_14792);
xnor U19150 (N_19150,N_13732,N_12860);
and U19151 (N_19151,N_12462,N_14647);
nor U19152 (N_19152,N_15701,N_15789);
and U19153 (N_19153,N_13880,N_14668);
nor U19154 (N_19154,N_12035,N_14670);
xnor U19155 (N_19155,N_15223,N_13292);
xnor U19156 (N_19156,N_15666,N_14501);
nand U19157 (N_19157,N_14419,N_12904);
nand U19158 (N_19158,N_14371,N_12983);
nor U19159 (N_19159,N_12847,N_15910);
nor U19160 (N_19160,N_15879,N_15505);
or U19161 (N_19161,N_14314,N_14647);
nand U19162 (N_19162,N_14071,N_15328);
nor U19163 (N_19163,N_15221,N_15758);
and U19164 (N_19164,N_15970,N_15249);
nand U19165 (N_19165,N_15398,N_15737);
nor U19166 (N_19166,N_13480,N_14082);
or U19167 (N_19167,N_14895,N_15798);
and U19168 (N_19168,N_12701,N_12680);
and U19169 (N_19169,N_12452,N_13890);
xor U19170 (N_19170,N_15826,N_15094);
or U19171 (N_19171,N_12572,N_14721);
or U19172 (N_19172,N_12830,N_15731);
or U19173 (N_19173,N_12675,N_13253);
and U19174 (N_19174,N_15714,N_12435);
nor U19175 (N_19175,N_12874,N_14073);
and U19176 (N_19176,N_12600,N_14366);
or U19177 (N_19177,N_13190,N_15235);
or U19178 (N_19178,N_14138,N_14312);
nand U19179 (N_19179,N_13157,N_13401);
or U19180 (N_19180,N_15072,N_15796);
or U19181 (N_19181,N_13127,N_15665);
nor U19182 (N_19182,N_15069,N_15598);
and U19183 (N_19183,N_12428,N_15033);
nand U19184 (N_19184,N_15805,N_12711);
nor U19185 (N_19185,N_13082,N_13091);
nor U19186 (N_19186,N_12954,N_13849);
or U19187 (N_19187,N_14172,N_13032);
nor U19188 (N_19188,N_15992,N_14417);
nor U19189 (N_19189,N_14921,N_14832);
nor U19190 (N_19190,N_14792,N_14766);
nor U19191 (N_19191,N_15440,N_14942);
nor U19192 (N_19192,N_15185,N_15324);
and U19193 (N_19193,N_14802,N_14973);
and U19194 (N_19194,N_15601,N_15884);
or U19195 (N_19195,N_15987,N_13614);
or U19196 (N_19196,N_15273,N_12153);
nor U19197 (N_19197,N_14510,N_13823);
nor U19198 (N_19198,N_14617,N_15704);
nor U19199 (N_19199,N_12696,N_14006);
nor U19200 (N_19200,N_13308,N_13482);
nor U19201 (N_19201,N_15276,N_12594);
or U19202 (N_19202,N_15235,N_15569);
xnor U19203 (N_19203,N_12878,N_15667);
nand U19204 (N_19204,N_12528,N_13834);
or U19205 (N_19205,N_12691,N_14796);
or U19206 (N_19206,N_12936,N_13746);
and U19207 (N_19207,N_13318,N_12921);
and U19208 (N_19208,N_15907,N_14615);
nand U19209 (N_19209,N_12817,N_15730);
nor U19210 (N_19210,N_13980,N_12486);
or U19211 (N_19211,N_15218,N_13738);
nor U19212 (N_19212,N_12320,N_15128);
or U19213 (N_19213,N_13213,N_12276);
nor U19214 (N_19214,N_13359,N_15037);
and U19215 (N_19215,N_15775,N_12282);
or U19216 (N_19216,N_13247,N_14394);
nor U19217 (N_19217,N_13885,N_13584);
nand U19218 (N_19218,N_13812,N_14935);
or U19219 (N_19219,N_12141,N_14564);
nor U19220 (N_19220,N_13935,N_12102);
or U19221 (N_19221,N_15030,N_15761);
or U19222 (N_19222,N_13021,N_15365);
or U19223 (N_19223,N_15460,N_12585);
nor U19224 (N_19224,N_14333,N_14789);
or U19225 (N_19225,N_12901,N_12238);
nor U19226 (N_19226,N_12311,N_14862);
and U19227 (N_19227,N_12633,N_15572);
or U19228 (N_19228,N_13027,N_15290);
or U19229 (N_19229,N_14111,N_13188);
and U19230 (N_19230,N_15503,N_15842);
xor U19231 (N_19231,N_14055,N_14909);
or U19232 (N_19232,N_14692,N_13942);
nand U19233 (N_19233,N_15466,N_15761);
nor U19234 (N_19234,N_15608,N_13297);
nand U19235 (N_19235,N_15851,N_14498);
nand U19236 (N_19236,N_15628,N_15917);
or U19237 (N_19237,N_14744,N_12158);
or U19238 (N_19238,N_15202,N_15383);
nor U19239 (N_19239,N_15376,N_14156);
and U19240 (N_19240,N_15948,N_12795);
and U19241 (N_19241,N_13906,N_14564);
and U19242 (N_19242,N_15277,N_13687);
and U19243 (N_19243,N_14259,N_13109);
and U19244 (N_19244,N_13136,N_13192);
or U19245 (N_19245,N_12704,N_12412);
and U19246 (N_19246,N_13022,N_15618);
or U19247 (N_19247,N_12624,N_12952);
nand U19248 (N_19248,N_12085,N_13487);
nand U19249 (N_19249,N_15439,N_12901);
or U19250 (N_19250,N_15887,N_14841);
or U19251 (N_19251,N_14005,N_15998);
or U19252 (N_19252,N_15858,N_14576);
or U19253 (N_19253,N_12938,N_15170);
and U19254 (N_19254,N_15772,N_14351);
nor U19255 (N_19255,N_14118,N_12588);
and U19256 (N_19256,N_12084,N_12242);
nor U19257 (N_19257,N_14109,N_15506);
nor U19258 (N_19258,N_13625,N_14055);
and U19259 (N_19259,N_13383,N_13088);
xor U19260 (N_19260,N_15593,N_15366);
nand U19261 (N_19261,N_12386,N_12115);
and U19262 (N_19262,N_14933,N_14399);
or U19263 (N_19263,N_14064,N_15166);
xnor U19264 (N_19264,N_12647,N_14180);
nor U19265 (N_19265,N_14638,N_13616);
xnor U19266 (N_19266,N_12962,N_13725);
and U19267 (N_19267,N_13768,N_15785);
or U19268 (N_19268,N_12296,N_12269);
nor U19269 (N_19269,N_15675,N_13473);
or U19270 (N_19270,N_14079,N_13598);
and U19271 (N_19271,N_15293,N_12257);
nand U19272 (N_19272,N_14501,N_14197);
nor U19273 (N_19273,N_13460,N_13080);
or U19274 (N_19274,N_15645,N_13294);
or U19275 (N_19275,N_13179,N_13261);
and U19276 (N_19276,N_13420,N_12279);
nor U19277 (N_19277,N_13103,N_14626);
and U19278 (N_19278,N_13640,N_13406);
and U19279 (N_19279,N_13309,N_15767);
or U19280 (N_19280,N_15019,N_12734);
xnor U19281 (N_19281,N_15395,N_13626);
or U19282 (N_19282,N_13842,N_13649);
and U19283 (N_19283,N_15535,N_13169);
and U19284 (N_19284,N_15197,N_12905);
or U19285 (N_19285,N_14109,N_15377);
xnor U19286 (N_19286,N_13282,N_12972);
and U19287 (N_19287,N_14455,N_15418);
nand U19288 (N_19288,N_13388,N_15176);
nor U19289 (N_19289,N_14238,N_14031);
nand U19290 (N_19290,N_13772,N_12300);
and U19291 (N_19291,N_14622,N_14337);
xor U19292 (N_19292,N_13416,N_15162);
nor U19293 (N_19293,N_12421,N_15064);
nand U19294 (N_19294,N_14623,N_12588);
and U19295 (N_19295,N_12249,N_13519);
nand U19296 (N_19296,N_14476,N_14357);
and U19297 (N_19297,N_14079,N_12454);
nor U19298 (N_19298,N_14814,N_12570);
or U19299 (N_19299,N_15391,N_15356);
nand U19300 (N_19300,N_12986,N_15621);
and U19301 (N_19301,N_15060,N_12002);
or U19302 (N_19302,N_13199,N_15068);
and U19303 (N_19303,N_15156,N_13386);
or U19304 (N_19304,N_13607,N_13815);
or U19305 (N_19305,N_13578,N_13392);
or U19306 (N_19306,N_12790,N_13129);
and U19307 (N_19307,N_14514,N_12696);
nor U19308 (N_19308,N_13572,N_14849);
nand U19309 (N_19309,N_15094,N_14900);
and U19310 (N_19310,N_15988,N_15326);
or U19311 (N_19311,N_15117,N_14026);
and U19312 (N_19312,N_14638,N_14716);
or U19313 (N_19313,N_12371,N_14867);
and U19314 (N_19314,N_15659,N_12267);
or U19315 (N_19315,N_12922,N_14968);
or U19316 (N_19316,N_15780,N_12251);
nand U19317 (N_19317,N_15706,N_13445);
or U19318 (N_19318,N_15761,N_13351);
and U19319 (N_19319,N_15509,N_15216);
nor U19320 (N_19320,N_14497,N_15465);
nor U19321 (N_19321,N_12484,N_15346);
nor U19322 (N_19322,N_12729,N_15621);
xnor U19323 (N_19323,N_14511,N_15797);
and U19324 (N_19324,N_13160,N_14348);
nor U19325 (N_19325,N_14717,N_13782);
nor U19326 (N_19326,N_13783,N_12322);
nand U19327 (N_19327,N_13361,N_15321);
nor U19328 (N_19328,N_15614,N_12379);
or U19329 (N_19329,N_13777,N_12459);
or U19330 (N_19330,N_12941,N_12256);
or U19331 (N_19331,N_13109,N_15841);
and U19332 (N_19332,N_14369,N_14639);
or U19333 (N_19333,N_14295,N_14925);
nand U19334 (N_19334,N_14300,N_13126);
or U19335 (N_19335,N_15455,N_13173);
nand U19336 (N_19336,N_12467,N_13851);
nand U19337 (N_19337,N_12410,N_12580);
or U19338 (N_19338,N_13338,N_15626);
or U19339 (N_19339,N_14564,N_14370);
nor U19340 (N_19340,N_14202,N_14535);
or U19341 (N_19341,N_14003,N_15767);
xor U19342 (N_19342,N_12006,N_13780);
nor U19343 (N_19343,N_15659,N_14604);
nand U19344 (N_19344,N_14202,N_13801);
nor U19345 (N_19345,N_12736,N_15141);
or U19346 (N_19346,N_15409,N_14590);
or U19347 (N_19347,N_14974,N_15676);
nor U19348 (N_19348,N_14966,N_15530);
nand U19349 (N_19349,N_12761,N_13763);
or U19350 (N_19350,N_15247,N_14848);
or U19351 (N_19351,N_13074,N_14448);
nand U19352 (N_19352,N_15522,N_14294);
nor U19353 (N_19353,N_13097,N_12544);
xor U19354 (N_19354,N_12750,N_14588);
and U19355 (N_19355,N_15690,N_12068);
and U19356 (N_19356,N_13260,N_15989);
nand U19357 (N_19357,N_12762,N_15518);
xnor U19358 (N_19358,N_12250,N_12791);
nor U19359 (N_19359,N_13353,N_12191);
or U19360 (N_19360,N_12106,N_13562);
nor U19361 (N_19361,N_15616,N_13066);
nor U19362 (N_19362,N_13308,N_12733);
nand U19363 (N_19363,N_13884,N_15543);
nor U19364 (N_19364,N_13515,N_15251);
and U19365 (N_19365,N_14584,N_15835);
nand U19366 (N_19366,N_12808,N_14576);
xnor U19367 (N_19367,N_13704,N_13817);
nand U19368 (N_19368,N_13455,N_15235);
or U19369 (N_19369,N_15520,N_14582);
nand U19370 (N_19370,N_13061,N_13956);
nand U19371 (N_19371,N_12165,N_14250);
and U19372 (N_19372,N_14776,N_12201);
nand U19373 (N_19373,N_14036,N_13740);
or U19374 (N_19374,N_13035,N_13743);
nor U19375 (N_19375,N_12775,N_12573);
and U19376 (N_19376,N_13414,N_12864);
xor U19377 (N_19377,N_13866,N_15688);
or U19378 (N_19378,N_13295,N_12513);
nor U19379 (N_19379,N_12279,N_14331);
nor U19380 (N_19380,N_13114,N_12654);
nor U19381 (N_19381,N_15969,N_12278);
nand U19382 (N_19382,N_12348,N_13362);
nor U19383 (N_19383,N_12724,N_12291);
and U19384 (N_19384,N_15376,N_14343);
nand U19385 (N_19385,N_14353,N_12343);
nor U19386 (N_19386,N_14166,N_14265);
xor U19387 (N_19387,N_14616,N_13837);
xor U19388 (N_19388,N_13020,N_14224);
and U19389 (N_19389,N_15399,N_15717);
or U19390 (N_19390,N_13765,N_13463);
and U19391 (N_19391,N_14549,N_15848);
nand U19392 (N_19392,N_12411,N_15274);
and U19393 (N_19393,N_14218,N_15741);
and U19394 (N_19394,N_12768,N_14625);
nor U19395 (N_19395,N_13201,N_13752);
nor U19396 (N_19396,N_12743,N_12313);
and U19397 (N_19397,N_15303,N_13292);
or U19398 (N_19398,N_13267,N_13109);
or U19399 (N_19399,N_13104,N_12649);
or U19400 (N_19400,N_12278,N_14281);
and U19401 (N_19401,N_13262,N_14856);
or U19402 (N_19402,N_14015,N_14164);
nor U19403 (N_19403,N_13957,N_15505);
nand U19404 (N_19404,N_14518,N_14679);
and U19405 (N_19405,N_14240,N_12343);
xnor U19406 (N_19406,N_12633,N_14317);
or U19407 (N_19407,N_14673,N_15332);
and U19408 (N_19408,N_14979,N_15838);
nand U19409 (N_19409,N_14785,N_14438);
xor U19410 (N_19410,N_12714,N_14729);
or U19411 (N_19411,N_13052,N_14009);
nor U19412 (N_19412,N_15900,N_12266);
nand U19413 (N_19413,N_15125,N_13070);
nor U19414 (N_19414,N_14194,N_12031);
and U19415 (N_19415,N_13283,N_15785);
nor U19416 (N_19416,N_13583,N_15738);
and U19417 (N_19417,N_14865,N_13202);
and U19418 (N_19418,N_15145,N_14370);
nand U19419 (N_19419,N_12574,N_15493);
and U19420 (N_19420,N_14188,N_13436);
and U19421 (N_19421,N_15600,N_14254);
and U19422 (N_19422,N_14906,N_12184);
nand U19423 (N_19423,N_15146,N_13136);
xnor U19424 (N_19424,N_15277,N_12871);
or U19425 (N_19425,N_12520,N_14339);
or U19426 (N_19426,N_12340,N_15428);
and U19427 (N_19427,N_12649,N_14991);
and U19428 (N_19428,N_13637,N_13691);
nor U19429 (N_19429,N_14836,N_13973);
nand U19430 (N_19430,N_15513,N_12358);
nor U19431 (N_19431,N_13408,N_15001);
or U19432 (N_19432,N_13076,N_15025);
nor U19433 (N_19433,N_13574,N_12307);
and U19434 (N_19434,N_13206,N_12954);
or U19435 (N_19435,N_13649,N_14839);
nor U19436 (N_19436,N_13249,N_13020);
or U19437 (N_19437,N_13277,N_14949);
and U19438 (N_19438,N_13721,N_12297);
nor U19439 (N_19439,N_12814,N_13320);
or U19440 (N_19440,N_13693,N_12102);
or U19441 (N_19441,N_12982,N_12000);
nor U19442 (N_19442,N_15720,N_12361);
or U19443 (N_19443,N_13706,N_12217);
and U19444 (N_19444,N_14766,N_14866);
nor U19445 (N_19445,N_12583,N_12486);
or U19446 (N_19446,N_13290,N_14602);
and U19447 (N_19447,N_13405,N_13765);
or U19448 (N_19448,N_15923,N_13831);
or U19449 (N_19449,N_13052,N_15556);
and U19450 (N_19450,N_12524,N_14147);
and U19451 (N_19451,N_12919,N_12742);
nor U19452 (N_19452,N_14765,N_14312);
nand U19453 (N_19453,N_14568,N_13218);
or U19454 (N_19454,N_14859,N_15137);
or U19455 (N_19455,N_14832,N_15584);
nand U19456 (N_19456,N_14356,N_14763);
nor U19457 (N_19457,N_15095,N_15500);
or U19458 (N_19458,N_14245,N_12022);
nand U19459 (N_19459,N_12041,N_12113);
nor U19460 (N_19460,N_14825,N_12661);
nand U19461 (N_19461,N_13183,N_12360);
and U19462 (N_19462,N_14557,N_12059);
and U19463 (N_19463,N_12894,N_13381);
nor U19464 (N_19464,N_13143,N_13182);
or U19465 (N_19465,N_14418,N_13329);
xnor U19466 (N_19466,N_15403,N_15725);
nand U19467 (N_19467,N_14486,N_12903);
nand U19468 (N_19468,N_13564,N_12281);
or U19469 (N_19469,N_12932,N_12865);
xnor U19470 (N_19470,N_13678,N_15352);
and U19471 (N_19471,N_15041,N_12728);
nor U19472 (N_19472,N_14718,N_13460);
and U19473 (N_19473,N_13947,N_12892);
nor U19474 (N_19474,N_12082,N_15057);
nand U19475 (N_19475,N_15032,N_15980);
nand U19476 (N_19476,N_14527,N_15569);
nor U19477 (N_19477,N_13315,N_12084);
and U19478 (N_19478,N_13407,N_13610);
or U19479 (N_19479,N_12402,N_14642);
or U19480 (N_19480,N_15176,N_14776);
nor U19481 (N_19481,N_12236,N_15334);
nand U19482 (N_19482,N_12075,N_14968);
nand U19483 (N_19483,N_13246,N_15497);
xnor U19484 (N_19484,N_15845,N_12498);
or U19485 (N_19485,N_14797,N_15080);
nand U19486 (N_19486,N_14795,N_13743);
nor U19487 (N_19487,N_14387,N_12027);
xnor U19488 (N_19488,N_13078,N_15370);
nand U19489 (N_19489,N_13384,N_15835);
nand U19490 (N_19490,N_15665,N_14387);
xnor U19491 (N_19491,N_14744,N_13911);
or U19492 (N_19492,N_12325,N_12830);
and U19493 (N_19493,N_13263,N_12800);
and U19494 (N_19494,N_13709,N_14066);
nor U19495 (N_19495,N_15730,N_13597);
and U19496 (N_19496,N_15945,N_15202);
or U19497 (N_19497,N_13534,N_12764);
nand U19498 (N_19498,N_13024,N_13365);
nor U19499 (N_19499,N_12374,N_14989);
nand U19500 (N_19500,N_14116,N_13791);
nor U19501 (N_19501,N_14667,N_15894);
or U19502 (N_19502,N_13494,N_13350);
and U19503 (N_19503,N_15992,N_12941);
nor U19504 (N_19504,N_13818,N_12835);
nor U19505 (N_19505,N_12794,N_14213);
xnor U19506 (N_19506,N_14544,N_14504);
and U19507 (N_19507,N_12082,N_14921);
nor U19508 (N_19508,N_13939,N_14801);
nor U19509 (N_19509,N_12744,N_14995);
or U19510 (N_19510,N_14702,N_15608);
nor U19511 (N_19511,N_12890,N_14539);
nor U19512 (N_19512,N_12096,N_13133);
and U19513 (N_19513,N_15994,N_13005);
nand U19514 (N_19514,N_14274,N_13085);
and U19515 (N_19515,N_15208,N_13325);
and U19516 (N_19516,N_15961,N_12820);
and U19517 (N_19517,N_15495,N_15037);
nor U19518 (N_19518,N_15046,N_12667);
and U19519 (N_19519,N_12970,N_12583);
nand U19520 (N_19520,N_14476,N_13185);
and U19521 (N_19521,N_15155,N_15680);
xor U19522 (N_19522,N_14575,N_13997);
or U19523 (N_19523,N_14045,N_13121);
or U19524 (N_19524,N_13941,N_14869);
nor U19525 (N_19525,N_12851,N_13186);
nand U19526 (N_19526,N_14812,N_13298);
nand U19527 (N_19527,N_15556,N_12122);
nor U19528 (N_19528,N_15032,N_15367);
or U19529 (N_19529,N_13920,N_13503);
nand U19530 (N_19530,N_13927,N_14761);
and U19531 (N_19531,N_12090,N_15330);
nand U19532 (N_19532,N_15204,N_12895);
or U19533 (N_19533,N_15099,N_15395);
nand U19534 (N_19534,N_12768,N_12857);
xnor U19535 (N_19535,N_14830,N_14764);
and U19536 (N_19536,N_14128,N_15729);
or U19537 (N_19537,N_12585,N_12139);
nand U19538 (N_19538,N_13162,N_13074);
nand U19539 (N_19539,N_14416,N_12307);
nand U19540 (N_19540,N_13721,N_12925);
nand U19541 (N_19541,N_15341,N_12816);
nor U19542 (N_19542,N_15221,N_13870);
nand U19543 (N_19543,N_12058,N_13518);
and U19544 (N_19544,N_14854,N_13802);
nand U19545 (N_19545,N_15426,N_15301);
or U19546 (N_19546,N_15291,N_12985);
nor U19547 (N_19547,N_12736,N_14029);
nand U19548 (N_19548,N_15340,N_13108);
or U19549 (N_19549,N_15040,N_14241);
nand U19550 (N_19550,N_12299,N_14959);
nor U19551 (N_19551,N_13274,N_12060);
and U19552 (N_19552,N_15721,N_13478);
nor U19553 (N_19553,N_14410,N_14478);
or U19554 (N_19554,N_12322,N_15894);
nand U19555 (N_19555,N_13165,N_14715);
or U19556 (N_19556,N_15151,N_15243);
nand U19557 (N_19557,N_14672,N_13689);
or U19558 (N_19558,N_15417,N_12692);
or U19559 (N_19559,N_13970,N_12223);
nor U19560 (N_19560,N_14482,N_14560);
or U19561 (N_19561,N_15001,N_13249);
and U19562 (N_19562,N_15401,N_13399);
and U19563 (N_19563,N_14607,N_14474);
or U19564 (N_19564,N_13300,N_15774);
and U19565 (N_19565,N_12765,N_14602);
and U19566 (N_19566,N_13543,N_12600);
xnor U19567 (N_19567,N_15214,N_13741);
nor U19568 (N_19568,N_13435,N_12063);
nand U19569 (N_19569,N_14838,N_14532);
and U19570 (N_19570,N_15124,N_13645);
xnor U19571 (N_19571,N_12155,N_12688);
and U19572 (N_19572,N_13967,N_15790);
xnor U19573 (N_19573,N_13869,N_13486);
nor U19574 (N_19574,N_15547,N_13284);
nand U19575 (N_19575,N_15124,N_15335);
nor U19576 (N_19576,N_14910,N_15397);
nor U19577 (N_19577,N_15058,N_14978);
nand U19578 (N_19578,N_14463,N_14877);
nand U19579 (N_19579,N_12263,N_14432);
nand U19580 (N_19580,N_13245,N_14531);
nor U19581 (N_19581,N_15709,N_14891);
nor U19582 (N_19582,N_14452,N_14075);
nand U19583 (N_19583,N_14782,N_14990);
nand U19584 (N_19584,N_14068,N_14963);
nor U19585 (N_19585,N_14687,N_12800);
or U19586 (N_19586,N_14696,N_12081);
nor U19587 (N_19587,N_14719,N_14413);
and U19588 (N_19588,N_13601,N_12309);
or U19589 (N_19589,N_12637,N_14501);
nand U19590 (N_19590,N_13034,N_15770);
and U19591 (N_19591,N_14064,N_15780);
or U19592 (N_19592,N_15803,N_13808);
nor U19593 (N_19593,N_13970,N_14585);
and U19594 (N_19594,N_12248,N_15678);
nand U19595 (N_19595,N_13679,N_12560);
and U19596 (N_19596,N_14804,N_13701);
nand U19597 (N_19597,N_15446,N_12970);
or U19598 (N_19598,N_13599,N_14176);
or U19599 (N_19599,N_15134,N_13114);
xnor U19600 (N_19600,N_12162,N_15981);
nand U19601 (N_19601,N_15121,N_12533);
or U19602 (N_19602,N_15719,N_12504);
and U19603 (N_19603,N_13236,N_14179);
nand U19604 (N_19604,N_13818,N_14437);
xor U19605 (N_19605,N_15246,N_15513);
or U19606 (N_19606,N_15382,N_13148);
nand U19607 (N_19607,N_14515,N_15257);
or U19608 (N_19608,N_14604,N_15030);
or U19609 (N_19609,N_12994,N_13189);
nor U19610 (N_19610,N_15824,N_13110);
and U19611 (N_19611,N_15835,N_13251);
or U19612 (N_19612,N_14894,N_12313);
nand U19613 (N_19613,N_12892,N_13650);
or U19614 (N_19614,N_13642,N_14934);
nor U19615 (N_19615,N_12174,N_13103);
or U19616 (N_19616,N_15975,N_15380);
and U19617 (N_19617,N_12690,N_14685);
nand U19618 (N_19618,N_12770,N_13722);
and U19619 (N_19619,N_13956,N_12998);
or U19620 (N_19620,N_15030,N_13071);
or U19621 (N_19621,N_13654,N_13678);
and U19622 (N_19622,N_12056,N_12377);
nor U19623 (N_19623,N_14299,N_15133);
and U19624 (N_19624,N_15265,N_12711);
or U19625 (N_19625,N_15446,N_14535);
nand U19626 (N_19626,N_14079,N_15152);
nand U19627 (N_19627,N_12482,N_12303);
or U19628 (N_19628,N_12183,N_13364);
nand U19629 (N_19629,N_15193,N_12295);
xor U19630 (N_19630,N_15263,N_12853);
nor U19631 (N_19631,N_12142,N_14408);
and U19632 (N_19632,N_14320,N_13233);
or U19633 (N_19633,N_12475,N_13681);
nand U19634 (N_19634,N_12497,N_15416);
nand U19635 (N_19635,N_15617,N_14595);
nor U19636 (N_19636,N_15851,N_15316);
nand U19637 (N_19637,N_14461,N_12016);
and U19638 (N_19638,N_14997,N_13627);
and U19639 (N_19639,N_12810,N_14740);
and U19640 (N_19640,N_12571,N_12819);
or U19641 (N_19641,N_13135,N_12770);
nand U19642 (N_19642,N_15207,N_13660);
nand U19643 (N_19643,N_15430,N_13811);
nor U19644 (N_19644,N_14299,N_15575);
or U19645 (N_19645,N_14058,N_15250);
nand U19646 (N_19646,N_15610,N_13708);
nor U19647 (N_19647,N_13859,N_14635);
nand U19648 (N_19648,N_12111,N_12016);
or U19649 (N_19649,N_13125,N_13153);
or U19650 (N_19650,N_15548,N_14925);
nor U19651 (N_19651,N_13224,N_13359);
and U19652 (N_19652,N_14973,N_12622);
nor U19653 (N_19653,N_14792,N_13236);
or U19654 (N_19654,N_15772,N_15153);
nor U19655 (N_19655,N_15512,N_15883);
and U19656 (N_19656,N_15487,N_15563);
nand U19657 (N_19657,N_12989,N_14034);
or U19658 (N_19658,N_12665,N_12307);
or U19659 (N_19659,N_12068,N_12066);
xnor U19660 (N_19660,N_14475,N_14467);
and U19661 (N_19661,N_14754,N_14809);
or U19662 (N_19662,N_15012,N_14611);
or U19663 (N_19663,N_15917,N_13609);
nor U19664 (N_19664,N_15831,N_13014);
and U19665 (N_19665,N_12457,N_13494);
or U19666 (N_19666,N_14528,N_12794);
and U19667 (N_19667,N_14826,N_13237);
nand U19668 (N_19668,N_13776,N_12136);
and U19669 (N_19669,N_15985,N_14527);
nand U19670 (N_19670,N_14461,N_15053);
nand U19671 (N_19671,N_15310,N_13157);
and U19672 (N_19672,N_14369,N_14082);
or U19673 (N_19673,N_13471,N_14664);
and U19674 (N_19674,N_13027,N_13810);
and U19675 (N_19675,N_13160,N_14120);
nand U19676 (N_19676,N_14080,N_12414);
nand U19677 (N_19677,N_15366,N_12015);
xnor U19678 (N_19678,N_15686,N_14100);
nand U19679 (N_19679,N_15263,N_12525);
nor U19680 (N_19680,N_13987,N_12368);
xor U19681 (N_19681,N_14199,N_15924);
nand U19682 (N_19682,N_15059,N_14603);
xnor U19683 (N_19683,N_14609,N_12270);
or U19684 (N_19684,N_13387,N_13630);
nor U19685 (N_19685,N_15044,N_15606);
and U19686 (N_19686,N_12781,N_12379);
nor U19687 (N_19687,N_15584,N_13456);
or U19688 (N_19688,N_14250,N_14185);
nand U19689 (N_19689,N_13714,N_15633);
nor U19690 (N_19690,N_14970,N_13357);
and U19691 (N_19691,N_13857,N_15823);
and U19692 (N_19692,N_15678,N_14925);
and U19693 (N_19693,N_15033,N_15614);
nor U19694 (N_19694,N_13869,N_15350);
and U19695 (N_19695,N_14594,N_14239);
and U19696 (N_19696,N_13657,N_15486);
xor U19697 (N_19697,N_13776,N_12283);
nor U19698 (N_19698,N_13224,N_12637);
and U19699 (N_19699,N_12100,N_12700);
nor U19700 (N_19700,N_14069,N_15197);
nor U19701 (N_19701,N_14098,N_13391);
and U19702 (N_19702,N_14557,N_15444);
and U19703 (N_19703,N_14747,N_14583);
nor U19704 (N_19704,N_14235,N_13048);
nand U19705 (N_19705,N_14756,N_15654);
or U19706 (N_19706,N_13310,N_13927);
or U19707 (N_19707,N_13061,N_15617);
or U19708 (N_19708,N_13946,N_13176);
nand U19709 (N_19709,N_13486,N_15274);
xor U19710 (N_19710,N_14127,N_15522);
nand U19711 (N_19711,N_13926,N_14858);
nor U19712 (N_19712,N_13545,N_13793);
nor U19713 (N_19713,N_13686,N_13386);
nor U19714 (N_19714,N_15172,N_14333);
nand U19715 (N_19715,N_14444,N_12970);
nor U19716 (N_19716,N_12862,N_14711);
nand U19717 (N_19717,N_15026,N_12145);
and U19718 (N_19718,N_14132,N_13134);
nand U19719 (N_19719,N_14073,N_14368);
nor U19720 (N_19720,N_15668,N_12942);
nor U19721 (N_19721,N_12315,N_14565);
or U19722 (N_19722,N_13743,N_12652);
nand U19723 (N_19723,N_15050,N_15816);
or U19724 (N_19724,N_12525,N_12866);
and U19725 (N_19725,N_13158,N_12238);
nand U19726 (N_19726,N_14565,N_12555);
nor U19727 (N_19727,N_12105,N_15697);
xnor U19728 (N_19728,N_12369,N_12722);
nand U19729 (N_19729,N_13865,N_12972);
xnor U19730 (N_19730,N_15806,N_14971);
or U19731 (N_19731,N_13879,N_12037);
and U19732 (N_19732,N_14210,N_14263);
and U19733 (N_19733,N_12680,N_12599);
nand U19734 (N_19734,N_14120,N_14126);
xnor U19735 (N_19735,N_15215,N_14850);
or U19736 (N_19736,N_15561,N_14283);
or U19737 (N_19737,N_12576,N_12356);
nand U19738 (N_19738,N_14786,N_13898);
nor U19739 (N_19739,N_14606,N_13028);
nor U19740 (N_19740,N_13021,N_13665);
and U19741 (N_19741,N_12776,N_15118);
and U19742 (N_19742,N_12327,N_14498);
nor U19743 (N_19743,N_15576,N_14035);
nor U19744 (N_19744,N_14776,N_15884);
nand U19745 (N_19745,N_12026,N_15523);
or U19746 (N_19746,N_14484,N_15867);
nand U19747 (N_19747,N_15775,N_14696);
nor U19748 (N_19748,N_13195,N_14201);
or U19749 (N_19749,N_14438,N_14949);
nor U19750 (N_19750,N_14748,N_12350);
and U19751 (N_19751,N_12976,N_15599);
and U19752 (N_19752,N_13618,N_12711);
or U19753 (N_19753,N_15757,N_15674);
xor U19754 (N_19754,N_13737,N_13939);
nor U19755 (N_19755,N_13724,N_14278);
nand U19756 (N_19756,N_15324,N_14412);
or U19757 (N_19757,N_13312,N_13320);
nor U19758 (N_19758,N_12246,N_13396);
and U19759 (N_19759,N_14641,N_13380);
nor U19760 (N_19760,N_15509,N_13193);
nor U19761 (N_19761,N_12168,N_15650);
or U19762 (N_19762,N_12478,N_12025);
xor U19763 (N_19763,N_13912,N_14299);
xor U19764 (N_19764,N_15082,N_13823);
and U19765 (N_19765,N_12021,N_13687);
nor U19766 (N_19766,N_13109,N_14638);
nand U19767 (N_19767,N_12545,N_12562);
nand U19768 (N_19768,N_15761,N_13729);
nand U19769 (N_19769,N_12814,N_13824);
and U19770 (N_19770,N_14893,N_12134);
or U19771 (N_19771,N_15806,N_14855);
and U19772 (N_19772,N_15701,N_15486);
nand U19773 (N_19773,N_15813,N_12293);
and U19774 (N_19774,N_12918,N_15705);
and U19775 (N_19775,N_12291,N_15675);
xnor U19776 (N_19776,N_15248,N_15256);
xnor U19777 (N_19777,N_15144,N_14581);
and U19778 (N_19778,N_14264,N_12487);
nor U19779 (N_19779,N_14682,N_12338);
and U19780 (N_19780,N_15224,N_15797);
and U19781 (N_19781,N_15294,N_15382);
nor U19782 (N_19782,N_13555,N_12913);
or U19783 (N_19783,N_13217,N_15816);
xnor U19784 (N_19784,N_14917,N_13824);
nor U19785 (N_19785,N_15637,N_15162);
or U19786 (N_19786,N_13978,N_12488);
nor U19787 (N_19787,N_13578,N_15263);
or U19788 (N_19788,N_15496,N_15932);
or U19789 (N_19789,N_12833,N_12838);
or U19790 (N_19790,N_14640,N_15267);
and U19791 (N_19791,N_14056,N_15107);
nor U19792 (N_19792,N_15261,N_13290);
or U19793 (N_19793,N_15647,N_15049);
xor U19794 (N_19794,N_12128,N_12715);
nor U19795 (N_19795,N_15521,N_13974);
or U19796 (N_19796,N_13811,N_13907);
nor U19797 (N_19797,N_12870,N_14675);
and U19798 (N_19798,N_15773,N_12693);
xor U19799 (N_19799,N_15004,N_15400);
nor U19800 (N_19800,N_15870,N_15270);
nor U19801 (N_19801,N_15244,N_15763);
and U19802 (N_19802,N_14257,N_13986);
nand U19803 (N_19803,N_13615,N_14556);
and U19804 (N_19804,N_14695,N_13995);
nor U19805 (N_19805,N_15401,N_15244);
or U19806 (N_19806,N_12846,N_12134);
nand U19807 (N_19807,N_12292,N_14213);
nand U19808 (N_19808,N_14783,N_13289);
and U19809 (N_19809,N_13460,N_12251);
nor U19810 (N_19810,N_14339,N_13938);
and U19811 (N_19811,N_12474,N_12877);
and U19812 (N_19812,N_15275,N_15085);
and U19813 (N_19813,N_15971,N_12428);
nand U19814 (N_19814,N_12162,N_14749);
and U19815 (N_19815,N_13006,N_13914);
or U19816 (N_19816,N_12955,N_12061);
or U19817 (N_19817,N_15204,N_13608);
or U19818 (N_19818,N_12613,N_15298);
nand U19819 (N_19819,N_13014,N_14844);
or U19820 (N_19820,N_14400,N_14903);
xnor U19821 (N_19821,N_14455,N_14019);
or U19822 (N_19822,N_14452,N_13569);
nor U19823 (N_19823,N_14419,N_14311);
nand U19824 (N_19824,N_12030,N_15847);
nor U19825 (N_19825,N_12359,N_13598);
nand U19826 (N_19826,N_14948,N_14282);
nor U19827 (N_19827,N_13789,N_12853);
or U19828 (N_19828,N_15140,N_15090);
and U19829 (N_19829,N_14993,N_13723);
nand U19830 (N_19830,N_15822,N_12697);
and U19831 (N_19831,N_12511,N_13754);
xnor U19832 (N_19832,N_14218,N_12224);
nor U19833 (N_19833,N_14635,N_14084);
xor U19834 (N_19834,N_15640,N_13937);
xnor U19835 (N_19835,N_13712,N_15897);
nor U19836 (N_19836,N_12958,N_14445);
nor U19837 (N_19837,N_15125,N_12235);
and U19838 (N_19838,N_13034,N_12233);
nand U19839 (N_19839,N_14952,N_15905);
and U19840 (N_19840,N_15993,N_15878);
or U19841 (N_19841,N_14014,N_15728);
and U19842 (N_19842,N_14561,N_15297);
nor U19843 (N_19843,N_13565,N_14561);
nand U19844 (N_19844,N_12554,N_12162);
nand U19845 (N_19845,N_13325,N_12444);
and U19846 (N_19846,N_13425,N_12002);
and U19847 (N_19847,N_15711,N_13100);
nor U19848 (N_19848,N_13979,N_13246);
or U19849 (N_19849,N_15803,N_13382);
and U19850 (N_19850,N_14081,N_15136);
xnor U19851 (N_19851,N_12703,N_15448);
xnor U19852 (N_19852,N_14783,N_15087);
nand U19853 (N_19853,N_15477,N_12091);
or U19854 (N_19854,N_12666,N_15513);
nor U19855 (N_19855,N_13810,N_12462);
nand U19856 (N_19856,N_12155,N_14803);
nor U19857 (N_19857,N_13659,N_15657);
and U19858 (N_19858,N_12725,N_15067);
nand U19859 (N_19859,N_13822,N_13358);
nor U19860 (N_19860,N_12037,N_14792);
nor U19861 (N_19861,N_12566,N_15932);
or U19862 (N_19862,N_12077,N_15167);
or U19863 (N_19863,N_13357,N_13198);
and U19864 (N_19864,N_12260,N_12520);
or U19865 (N_19865,N_13473,N_14629);
nand U19866 (N_19866,N_14305,N_14302);
or U19867 (N_19867,N_13190,N_14938);
nor U19868 (N_19868,N_12100,N_14853);
nor U19869 (N_19869,N_12647,N_14752);
and U19870 (N_19870,N_14529,N_13501);
nor U19871 (N_19871,N_15909,N_12461);
nor U19872 (N_19872,N_14317,N_12780);
nand U19873 (N_19873,N_13885,N_15133);
or U19874 (N_19874,N_13417,N_14330);
or U19875 (N_19875,N_12717,N_13141);
nand U19876 (N_19876,N_13135,N_15591);
and U19877 (N_19877,N_14176,N_14746);
nand U19878 (N_19878,N_14431,N_13804);
and U19879 (N_19879,N_14026,N_12379);
nand U19880 (N_19880,N_15113,N_12311);
nor U19881 (N_19881,N_12991,N_14830);
or U19882 (N_19882,N_15564,N_15741);
or U19883 (N_19883,N_15564,N_15520);
and U19884 (N_19884,N_15101,N_14063);
or U19885 (N_19885,N_14385,N_14989);
or U19886 (N_19886,N_15946,N_12455);
or U19887 (N_19887,N_13860,N_15783);
nand U19888 (N_19888,N_12284,N_14396);
xnor U19889 (N_19889,N_12967,N_15469);
nand U19890 (N_19890,N_15368,N_14277);
and U19891 (N_19891,N_12768,N_13453);
xor U19892 (N_19892,N_15334,N_14958);
or U19893 (N_19893,N_14268,N_12695);
nor U19894 (N_19894,N_12476,N_12640);
nor U19895 (N_19895,N_13420,N_12800);
and U19896 (N_19896,N_13068,N_12466);
nor U19897 (N_19897,N_14893,N_15341);
or U19898 (N_19898,N_14659,N_13713);
nand U19899 (N_19899,N_12925,N_15327);
and U19900 (N_19900,N_12411,N_12673);
nand U19901 (N_19901,N_12915,N_13006);
nor U19902 (N_19902,N_14256,N_15273);
xnor U19903 (N_19903,N_12555,N_14073);
or U19904 (N_19904,N_15951,N_12447);
or U19905 (N_19905,N_15239,N_13702);
xor U19906 (N_19906,N_14551,N_13040);
xor U19907 (N_19907,N_13980,N_15794);
nand U19908 (N_19908,N_13172,N_14986);
or U19909 (N_19909,N_14809,N_14381);
nor U19910 (N_19910,N_12524,N_13271);
xor U19911 (N_19911,N_13737,N_12030);
nand U19912 (N_19912,N_14423,N_15470);
nand U19913 (N_19913,N_15106,N_14268);
or U19914 (N_19914,N_14618,N_14862);
and U19915 (N_19915,N_13944,N_14658);
nand U19916 (N_19916,N_14769,N_12352);
or U19917 (N_19917,N_12556,N_13300);
or U19918 (N_19918,N_14317,N_14699);
and U19919 (N_19919,N_12922,N_14259);
and U19920 (N_19920,N_14172,N_15473);
and U19921 (N_19921,N_12140,N_14604);
and U19922 (N_19922,N_12084,N_12326);
and U19923 (N_19923,N_15560,N_13913);
or U19924 (N_19924,N_12445,N_14127);
or U19925 (N_19925,N_12747,N_14635);
xnor U19926 (N_19926,N_13389,N_14503);
nor U19927 (N_19927,N_15267,N_13800);
nor U19928 (N_19928,N_12547,N_13581);
nand U19929 (N_19929,N_13084,N_15721);
nand U19930 (N_19930,N_13846,N_14765);
nor U19931 (N_19931,N_14730,N_13689);
xor U19932 (N_19932,N_14577,N_15114);
xnor U19933 (N_19933,N_13948,N_15351);
or U19934 (N_19934,N_14439,N_13990);
or U19935 (N_19935,N_12189,N_12150);
and U19936 (N_19936,N_13255,N_12606);
nand U19937 (N_19937,N_15469,N_14141);
nand U19938 (N_19938,N_14449,N_13866);
nor U19939 (N_19939,N_12104,N_12991);
and U19940 (N_19940,N_13326,N_15062);
nor U19941 (N_19941,N_15287,N_14601);
xor U19942 (N_19942,N_14692,N_15228);
and U19943 (N_19943,N_14377,N_12356);
or U19944 (N_19944,N_13412,N_14678);
and U19945 (N_19945,N_15195,N_14237);
or U19946 (N_19946,N_15893,N_15709);
and U19947 (N_19947,N_15242,N_15299);
nand U19948 (N_19948,N_15603,N_12190);
nor U19949 (N_19949,N_12284,N_15786);
xnor U19950 (N_19950,N_13181,N_13508);
or U19951 (N_19951,N_14392,N_12280);
nor U19952 (N_19952,N_14724,N_13718);
or U19953 (N_19953,N_14399,N_12456);
or U19954 (N_19954,N_12143,N_15844);
nor U19955 (N_19955,N_12168,N_12217);
nand U19956 (N_19956,N_13918,N_12482);
nand U19957 (N_19957,N_12636,N_15749);
nand U19958 (N_19958,N_13327,N_15522);
and U19959 (N_19959,N_15417,N_15158);
and U19960 (N_19960,N_12132,N_12629);
nand U19961 (N_19961,N_13587,N_14499);
nor U19962 (N_19962,N_14011,N_13340);
nor U19963 (N_19963,N_14270,N_15594);
or U19964 (N_19964,N_15769,N_15824);
or U19965 (N_19965,N_14084,N_12631);
and U19966 (N_19966,N_15548,N_15708);
and U19967 (N_19967,N_15880,N_13775);
nor U19968 (N_19968,N_12015,N_14590);
xnor U19969 (N_19969,N_15690,N_12827);
nand U19970 (N_19970,N_15576,N_15419);
and U19971 (N_19971,N_13106,N_12566);
or U19972 (N_19972,N_15595,N_12810);
nand U19973 (N_19973,N_12602,N_14915);
nor U19974 (N_19974,N_13247,N_12255);
nor U19975 (N_19975,N_14175,N_12725);
nor U19976 (N_19976,N_14398,N_13666);
or U19977 (N_19977,N_13179,N_13565);
and U19978 (N_19978,N_12786,N_15280);
xor U19979 (N_19979,N_13218,N_12104);
xnor U19980 (N_19980,N_14296,N_13082);
nor U19981 (N_19981,N_13620,N_14221);
nand U19982 (N_19982,N_13610,N_14503);
nand U19983 (N_19983,N_13681,N_12923);
nand U19984 (N_19984,N_13567,N_15055);
and U19985 (N_19985,N_13689,N_15630);
nor U19986 (N_19986,N_14136,N_15152);
nor U19987 (N_19987,N_14735,N_14572);
nand U19988 (N_19988,N_15586,N_14227);
or U19989 (N_19989,N_15218,N_14655);
nand U19990 (N_19990,N_13132,N_15998);
nor U19991 (N_19991,N_15726,N_13701);
nor U19992 (N_19992,N_13824,N_15972);
nor U19993 (N_19993,N_14584,N_12864);
or U19994 (N_19994,N_13314,N_12624);
nor U19995 (N_19995,N_12433,N_12445);
and U19996 (N_19996,N_14788,N_13897);
nor U19997 (N_19997,N_14674,N_14580);
nand U19998 (N_19998,N_13315,N_15808);
or U19999 (N_19999,N_15330,N_14407);
or UO_0 (O_0,N_16927,N_19802);
nor UO_1 (O_1,N_18544,N_19635);
and UO_2 (O_2,N_19069,N_18638);
nand UO_3 (O_3,N_16339,N_17625);
nand UO_4 (O_4,N_19173,N_18237);
and UO_5 (O_5,N_18923,N_16215);
nor UO_6 (O_6,N_17218,N_17225);
xnor UO_7 (O_7,N_16144,N_17581);
or UO_8 (O_8,N_16479,N_16801);
or UO_9 (O_9,N_16537,N_18150);
or UO_10 (O_10,N_16253,N_17338);
nand UO_11 (O_11,N_19454,N_16994);
nand UO_12 (O_12,N_19497,N_17854);
nand UO_13 (O_13,N_16976,N_19111);
or UO_14 (O_14,N_16422,N_16500);
and UO_15 (O_15,N_19983,N_17888);
nand UO_16 (O_16,N_18689,N_19153);
nand UO_17 (O_17,N_17297,N_16607);
or UO_18 (O_18,N_17857,N_16900);
or UO_19 (O_19,N_17066,N_16409);
and UO_20 (O_20,N_19797,N_16876);
or UO_21 (O_21,N_18363,N_18169);
nand UO_22 (O_22,N_18655,N_19106);
or UO_23 (O_23,N_16275,N_16972);
and UO_24 (O_24,N_17903,N_18490);
nand UO_25 (O_25,N_19676,N_19927);
or UO_26 (O_26,N_19700,N_16267);
xor UO_27 (O_27,N_17173,N_19114);
nor UO_28 (O_28,N_16341,N_16269);
xor UO_29 (O_29,N_18778,N_19589);
nand UO_30 (O_30,N_19396,N_19368);
or UO_31 (O_31,N_19036,N_16757);
xnor UO_32 (O_32,N_19437,N_16733);
and UO_33 (O_33,N_18652,N_18178);
and UO_34 (O_34,N_19044,N_16162);
xor UO_35 (O_35,N_19350,N_18665);
or UO_36 (O_36,N_18011,N_18849);
nor UO_37 (O_37,N_17547,N_17586);
or UO_38 (O_38,N_19076,N_16213);
nor UO_39 (O_39,N_16728,N_18523);
nand UO_40 (O_40,N_18780,N_19161);
nand UO_41 (O_41,N_18010,N_17263);
nor UO_42 (O_42,N_18838,N_19181);
xor UO_43 (O_43,N_17315,N_17734);
xor UO_44 (O_44,N_19914,N_18208);
nor UO_45 (O_45,N_18503,N_16735);
nand UO_46 (O_46,N_19549,N_18513);
or UO_47 (O_47,N_18160,N_18984);
nor UO_48 (O_48,N_17606,N_17317);
nand UO_49 (O_49,N_16989,N_17559);
xor UO_50 (O_50,N_17591,N_17298);
and UO_51 (O_51,N_16217,N_19159);
xnor UO_52 (O_52,N_19449,N_17920);
or UO_53 (O_53,N_18775,N_17406);
or UO_54 (O_54,N_16055,N_17032);
nor UO_55 (O_55,N_18432,N_16608);
nand UO_56 (O_56,N_18392,N_19451);
xor UO_57 (O_57,N_18221,N_19593);
nor UO_58 (O_58,N_19464,N_17147);
nand UO_59 (O_59,N_18761,N_17222);
xnor UO_60 (O_60,N_16390,N_19766);
nand UO_61 (O_61,N_17480,N_16738);
or UO_62 (O_62,N_16291,N_18265);
nor UO_63 (O_63,N_16377,N_16872);
nor UO_64 (O_64,N_18582,N_19493);
nand UO_65 (O_65,N_16957,N_17042);
nor UO_66 (O_66,N_17486,N_16060);
nand UO_67 (O_67,N_17993,N_17733);
nor UO_68 (O_68,N_17724,N_16788);
nor UO_69 (O_69,N_18342,N_19892);
nand UO_70 (O_70,N_16312,N_18380);
and UO_71 (O_71,N_17487,N_17189);
nand UO_72 (O_72,N_18765,N_19308);
nor UO_73 (O_73,N_19572,N_16464);
nor UO_74 (O_74,N_18646,N_19525);
or UO_75 (O_75,N_18969,N_17580);
and UO_76 (O_76,N_17550,N_16015);
and UO_77 (O_77,N_19431,N_16914);
or UO_78 (O_78,N_19697,N_17195);
nand UO_79 (O_79,N_16476,N_18797);
or UO_80 (O_80,N_19100,N_19316);
or UO_81 (O_81,N_17514,N_18678);
nor UO_82 (O_82,N_16486,N_19801);
nor UO_83 (O_83,N_16621,N_17398);
nand UO_84 (O_84,N_19864,N_18602);
and UO_85 (O_85,N_19299,N_18867);
nor UO_86 (O_86,N_17275,N_17707);
nor UO_87 (O_87,N_19188,N_18756);
nand UO_88 (O_88,N_16897,N_19861);
nor UO_89 (O_89,N_17078,N_18478);
nor UO_90 (O_90,N_16261,N_18177);
nand UO_91 (O_91,N_16962,N_18938);
nand UO_92 (O_92,N_17118,N_17468);
nand UO_93 (O_93,N_16798,N_19664);
nor UO_94 (O_94,N_19381,N_18092);
nor UO_95 (O_95,N_18215,N_19942);
xor UO_96 (O_96,N_16321,N_19195);
xor UO_97 (O_97,N_17153,N_19594);
nor UO_98 (O_98,N_17385,N_16161);
nand UO_99 (O_99,N_17822,N_18660);
and UO_100 (O_100,N_19614,N_19947);
nand UO_101 (O_101,N_19756,N_19535);
nor UO_102 (O_102,N_18805,N_17171);
or UO_103 (O_103,N_18324,N_19580);
nand UO_104 (O_104,N_19783,N_19731);
and UO_105 (O_105,N_19187,N_16128);
nand UO_106 (O_106,N_17249,N_16909);
or UO_107 (O_107,N_17785,N_16841);
nor UO_108 (O_108,N_17867,N_17889);
nor UO_109 (O_109,N_18101,N_18136);
and UO_110 (O_110,N_16455,N_17834);
or UO_111 (O_111,N_17403,N_17124);
nor UO_112 (O_112,N_19209,N_16330);
or UO_113 (O_113,N_18421,N_18212);
nor UO_114 (O_114,N_17271,N_18257);
nand UO_115 (O_115,N_17200,N_19498);
or UO_116 (O_116,N_19415,N_16838);
xnor UO_117 (O_117,N_17278,N_19787);
xor UO_118 (O_118,N_16651,N_18075);
xor UO_119 (O_119,N_19315,N_17191);
and UO_120 (O_120,N_19799,N_16539);
nand UO_121 (O_121,N_16629,N_16765);
nor UO_122 (O_122,N_17425,N_18123);
nor UO_123 (O_123,N_18524,N_19835);
or UO_124 (O_124,N_16222,N_19006);
nand UO_125 (O_125,N_18773,N_19110);
nand UO_126 (O_126,N_16137,N_18796);
nor UO_127 (O_127,N_19786,N_16238);
or UO_128 (O_128,N_18271,N_16953);
nand UO_129 (O_129,N_19280,N_17073);
xor UO_130 (O_130,N_19823,N_16378);
and UO_131 (O_131,N_16038,N_16940);
and UO_132 (O_132,N_19653,N_18337);
nor UO_133 (O_133,N_17201,N_16535);
or UO_134 (O_134,N_16787,N_16856);
nor UO_135 (O_135,N_17915,N_19333);
nand UO_136 (O_136,N_18681,N_18076);
and UO_137 (O_137,N_18433,N_19916);
or UO_138 (O_138,N_16984,N_16100);
nor UO_139 (O_139,N_16742,N_16916);
or UO_140 (O_140,N_16827,N_16285);
and UO_141 (O_141,N_16487,N_17035);
nand UO_142 (O_142,N_16103,N_18167);
nor UO_143 (O_143,N_18930,N_17618);
nor UO_144 (O_144,N_17143,N_17146);
nor UO_145 (O_145,N_19618,N_18273);
or UO_146 (O_146,N_19105,N_18145);
nand UO_147 (O_147,N_19936,N_18514);
nand UO_148 (O_148,N_18522,N_18133);
nand UO_149 (O_149,N_18924,N_19900);
or UO_150 (O_150,N_18767,N_18632);
and UO_151 (O_151,N_16620,N_18459);
xor UO_152 (O_152,N_16094,N_19112);
or UO_153 (O_153,N_18072,N_17764);
and UO_154 (O_154,N_18233,N_17387);
and UO_155 (O_155,N_19721,N_19046);
and UO_156 (O_156,N_16702,N_17163);
or UO_157 (O_157,N_16048,N_16926);
nor UO_158 (O_158,N_17941,N_19042);
and UO_159 (O_159,N_19517,N_16525);
nand UO_160 (O_160,N_16745,N_17177);
and UO_161 (O_161,N_17790,N_16337);
nand UO_162 (O_162,N_16711,N_19893);
xor UO_163 (O_163,N_19930,N_17028);
nand UO_164 (O_164,N_17861,N_18134);
xor UO_165 (O_165,N_19544,N_18279);
nor UO_166 (O_166,N_18998,N_16781);
nor UO_167 (O_167,N_17156,N_18376);
or UO_168 (O_168,N_17906,N_17870);
or UO_169 (O_169,N_19443,N_16043);
and UO_170 (O_170,N_19859,N_17865);
nand UO_171 (O_171,N_18567,N_17248);
or UO_172 (O_172,N_19142,N_18083);
or UO_173 (O_173,N_17560,N_17700);
nand UO_174 (O_174,N_19473,N_17182);
or UO_175 (O_175,N_16397,N_18809);
or UO_176 (O_176,N_16573,N_17197);
and UO_177 (O_177,N_17869,N_16230);
and UO_178 (O_178,N_16670,N_17240);
or UO_179 (O_179,N_19248,N_17001);
and UO_180 (O_180,N_19379,N_16344);
or UO_181 (O_181,N_19180,N_18776);
or UO_182 (O_182,N_19027,N_16502);
or UO_183 (O_183,N_16513,N_16085);
or UO_184 (O_184,N_16718,N_19842);
xor UO_185 (O_185,N_18369,N_16859);
xnor UO_186 (O_186,N_17310,N_18926);
nor UO_187 (O_187,N_16430,N_17755);
and UO_188 (O_188,N_18149,N_16287);
nand UO_189 (O_189,N_17646,N_18774);
and UO_190 (O_190,N_18953,N_18240);
nand UO_191 (O_191,N_18539,N_17098);
nor UO_192 (O_192,N_17166,N_17352);
nor UO_193 (O_193,N_19353,N_17185);
and UO_194 (O_194,N_19639,N_16700);
and UO_195 (O_195,N_18563,N_19685);
and UO_196 (O_196,N_16325,N_17285);
xnor UO_197 (O_197,N_18649,N_18738);
and UO_198 (O_198,N_19662,N_19107);
nand UO_199 (O_199,N_19122,N_19926);
or UO_200 (O_200,N_19845,N_18473);
xnor UO_201 (O_201,N_19829,N_17070);
and UO_202 (O_202,N_19463,N_19837);
nand UO_203 (O_203,N_17244,N_19509);
or UO_204 (O_204,N_19072,N_18398);
and UO_205 (O_205,N_18744,N_19274);
and UO_206 (O_206,N_16208,N_19256);
and UO_207 (O_207,N_17928,N_17303);
nor UO_208 (O_208,N_17706,N_18635);
nor UO_209 (O_209,N_18364,N_16165);
and UO_210 (O_210,N_17718,N_16991);
xor UO_211 (O_211,N_17830,N_16488);
and UO_212 (O_212,N_19411,N_19850);
nand UO_213 (O_213,N_17904,N_19601);
xor UO_214 (O_214,N_19230,N_18664);
nor UO_215 (O_215,N_17509,N_17927);
or UO_216 (O_216,N_16109,N_18970);
xnor UO_217 (O_217,N_16681,N_16760);
nor UO_218 (O_218,N_16066,N_16080);
or UO_219 (O_219,N_16126,N_16402);
nand UO_220 (O_220,N_16532,N_17626);
nor UO_221 (O_221,N_18294,N_19022);
nand UO_222 (O_222,N_19945,N_19887);
and UO_223 (O_223,N_17630,N_17256);
or UO_224 (O_224,N_18734,N_18086);
nor UO_225 (O_225,N_18572,N_18746);
nor UO_226 (O_226,N_16522,N_16861);
nor UO_227 (O_227,N_17100,N_17607);
and UO_228 (O_228,N_18877,N_17172);
nor UO_229 (O_229,N_18583,N_16857);
nand UO_230 (O_230,N_18856,N_18094);
or UO_231 (O_231,N_16361,N_19420);
or UO_232 (O_232,N_19149,N_16617);
and UO_233 (O_233,N_19476,N_18210);
or UO_234 (O_234,N_18782,N_17539);
nand UO_235 (O_235,N_17094,N_18601);
or UO_236 (O_236,N_19569,N_16610);
xnor UO_237 (O_237,N_19247,N_18585);
or UO_238 (O_238,N_18165,N_19693);
nand UO_239 (O_239,N_17392,N_17134);
or UO_240 (O_240,N_16188,N_18549);
nor UO_241 (O_241,N_16258,N_19706);
or UO_242 (O_242,N_18708,N_17307);
or UO_243 (O_243,N_16709,N_19583);
nor UO_244 (O_244,N_16364,N_18203);
nand UO_245 (O_245,N_18573,N_17939);
nor UO_246 (O_246,N_16392,N_17199);
and UO_247 (O_247,N_19421,N_16968);
nand UO_248 (O_248,N_18770,N_18079);
or UO_249 (O_249,N_19559,N_16353);
or UO_250 (O_250,N_17350,N_17916);
nor UO_251 (O_251,N_18834,N_17531);
nand UO_252 (O_252,N_17577,N_17322);
and UO_253 (O_253,N_19692,N_17292);
nand UO_254 (O_254,N_18625,N_19956);
nor UO_255 (O_255,N_19527,N_16919);
nand UO_256 (O_256,N_18329,N_18644);
nand UO_257 (O_257,N_17252,N_19494);
xor UO_258 (O_258,N_17578,N_19041);
nand UO_259 (O_259,N_18587,N_16021);
or UO_260 (O_260,N_17803,N_16963);
and UO_261 (O_261,N_17731,N_19375);
or UO_262 (O_262,N_17568,N_17912);
or UO_263 (O_263,N_18758,N_16234);
or UO_264 (O_264,N_19546,N_18736);
nand UO_265 (O_265,N_17662,N_18084);
nor UO_266 (O_266,N_16075,N_17858);
nand UO_267 (O_267,N_18052,N_17407);
or UO_268 (O_268,N_18619,N_17769);
or UO_269 (O_269,N_16945,N_18491);
or UO_270 (O_270,N_18304,N_19975);
and UO_271 (O_271,N_18438,N_19907);
nor UO_272 (O_272,N_16682,N_17132);
or UO_273 (O_273,N_17207,N_19393);
nor UO_274 (O_274,N_18124,N_18568);
and UO_275 (O_275,N_18760,N_18351);
nand UO_276 (O_276,N_17289,N_17048);
or UO_277 (O_277,N_18263,N_19383);
xnor UO_278 (O_278,N_18295,N_17893);
nand UO_279 (O_279,N_17072,N_16491);
and UO_280 (O_280,N_18201,N_18229);
nor UO_281 (O_281,N_17800,N_17148);
and UO_282 (O_282,N_16047,N_16351);
nor UO_283 (O_283,N_17461,N_17507);
or UO_284 (O_284,N_17695,N_18395);
xnor UO_285 (O_285,N_18799,N_19796);
nand UO_286 (O_286,N_17367,N_19874);
nand UO_287 (O_287,N_16264,N_18489);
nor UO_288 (O_288,N_19918,N_19322);
xor UO_289 (O_289,N_19143,N_16317);
or UO_290 (O_290,N_17672,N_17670);
or UO_291 (O_291,N_17023,N_17235);
or UO_292 (O_292,N_19960,N_16866);
nand UO_293 (O_293,N_16619,N_16133);
or UO_294 (O_294,N_19735,N_17313);
and UO_295 (O_295,N_18220,N_16041);
nor UO_296 (O_296,N_17737,N_17573);
nor UO_297 (O_297,N_17515,N_18691);
nand UO_298 (O_298,N_19698,N_18002);
and UO_299 (O_299,N_16555,N_18197);
and UO_300 (O_300,N_19656,N_18902);
nand UO_301 (O_301,N_18496,N_18061);
nor UO_302 (O_302,N_18735,N_18190);
nand UO_303 (O_303,N_19913,N_18358);
nor UO_304 (O_304,N_17575,N_17549);
nor UO_305 (O_305,N_19867,N_17837);
nor UO_306 (O_306,N_18727,N_17886);
nand UO_307 (O_307,N_17015,N_16673);
and UO_308 (O_308,N_17880,N_18748);
nand UO_309 (O_309,N_19284,N_18250);
nor UO_310 (O_310,N_19467,N_16400);
nor UO_311 (O_311,N_16444,N_17829);
nor UO_312 (O_312,N_19189,N_19007);
nand UO_313 (O_313,N_19880,N_19577);
or UO_314 (O_314,N_19031,N_16674);
nor UO_315 (O_315,N_18670,N_17752);
and UO_316 (O_316,N_16497,N_18538);
nor UO_317 (O_317,N_17205,N_16921);
or UO_318 (O_318,N_16858,N_18087);
nor UO_319 (O_319,N_18246,N_16379);
or UO_320 (O_320,N_16791,N_16245);
xnor UO_321 (O_321,N_19456,N_16393);
or UO_322 (O_322,N_19165,N_16756);
nand UO_323 (O_323,N_18298,N_16563);
or UO_324 (O_324,N_19726,N_18707);
xor UO_325 (O_325,N_17610,N_17597);
nand UO_326 (O_326,N_16106,N_19070);
nand UO_327 (O_327,N_17418,N_16218);
and UO_328 (O_328,N_18786,N_19896);
or UO_329 (O_329,N_17125,N_17566);
and UO_330 (O_330,N_19255,N_16045);
nor UO_331 (O_331,N_16837,N_19462);
nand UO_332 (O_332,N_18403,N_17410);
or UO_333 (O_333,N_16216,N_17596);
and UO_334 (O_334,N_17684,N_18267);
nor UO_335 (O_335,N_18128,N_17457);
and UO_336 (O_336,N_16068,N_19533);
or UO_337 (O_337,N_18534,N_18604);
or UO_338 (O_338,N_16835,N_18719);
nand UO_339 (O_339,N_16202,N_17828);
or UO_340 (O_340,N_18559,N_17046);
nor UO_341 (O_341,N_16928,N_19037);
xor UO_342 (O_342,N_17698,N_17295);
and UO_343 (O_343,N_18091,N_16741);
or UO_344 (O_344,N_18182,N_17603);
nand UO_345 (O_345,N_19419,N_17756);
or UO_346 (O_346,N_19005,N_17429);
nor UO_347 (O_347,N_16567,N_16243);
nand UO_348 (O_348,N_16039,N_19374);
nand UO_349 (O_349,N_16214,N_17004);
xnor UO_350 (O_350,N_17192,N_19434);
nor UO_351 (O_351,N_16751,N_18600);
nand UO_352 (O_352,N_16394,N_18181);
nor UO_353 (O_353,N_19258,N_17114);
and UO_354 (O_354,N_18898,N_16889);
and UO_355 (O_355,N_17679,N_16210);
xor UO_356 (O_356,N_17704,N_16528);
and UO_357 (O_357,N_19313,N_18439);
and UO_358 (O_358,N_17516,N_16707);
and UO_359 (O_359,N_17950,N_18289);
nand UO_360 (O_360,N_16286,N_17103);
nand UO_361 (O_361,N_18561,N_17930);
nand UO_362 (O_362,N_16730,N_19788);
nand UO_363 (O_363,N_17759,N_19403);
nor UO_364 (O_364,N_19581,N_16524);
nand UO_365 (O_365,N_18135,N_19665);
or UO_366 (O_366,N_18402,N_17699);
nor UO_367 (O_367,N_19970,N_19879);
and UO_368 (O_368,N_16772,N_17556);
xor UO_369 (O_369,N_18677,N_19045);
and UO_370 (O_370,N_19470,N_17652);
xor UO_371 (O_371,N_16187,N_16521);
or UO_372 (O_372,N_19441,N_17284);
nor UO_373 (O_373,N_17017,N_18219);
and UO_374 (O_374,N_17989,N_17126);
or UO_375 (O_375,N_16884,N_19125);
xnor UO_376 (O_376,N_16970,N_16863);
xor UO_377 (O_377,N_18308,N_19634);
nand UO_378 (O_378,N_16587,N_19598);
or UO_379 (O_379,N_16583,N_18952);
nand UO_380 (O_380,N_19741,N_18495);
or UO_381 (O_381,N_19172,N_18252);
xnor UO_382 (O_382,N_18798,N_16936);
xor UO_383 (O_383,N_16604,N_17663);
nand UO_384 (O_384,N_18527,N_16153);
or UO_385 (O_385,N_18116,N_18310);
nand UO_386 (O_386,N_18792,N_16731);
nand UO_387 (O_387,N_16118,N_16578);
nand UO_388 (O_388,N_18469,N_19862);
or UO_389 (O_389,N_17446,N_17839);
or UO_390 (O_390,N_18096,N_17938);
nor UO_391 (O_391,N_18204,N_16495);
and UO_392 (O_392,N_17376,N_17499);
nand UO_393 (O_393,N_18547,N_18187);
nor UO_394 (O_394,N_17542,N_18880);
nor UO_395 (O_395,N_18418,N_18319);
or UO_396 (O_396,N_19144,N_16618);
nor UO_397 (O_397,N_19827,N_19919);
nor UO_398 (O_398,N_19097,N_16997);
nand UO_399 (O_399,N_19809,N_17453);
nor UO_400 (O_400,N_19283,N_16265);
nand UO_401 (O_401,N_18893,N_19009);
nor UO_402 (O_402,N_17361,N_17783);
xnor UO_403 (O_403,N_16037,N_19026);
nand UO_404 (O_404,N_17423,N_18785);
nor UO_405 (O_405,N_19273,N_18725);
nor UO_406 (O_406,N_19344,N_18891);
nand UO_407 (O_407,N_16182,N_16070);
and UO_408 (O_408,N_18662,N_16538);
and UO_409 (O_409,N_16964,N_17943);
xor UO_410 (O_410,N_19643,N_17341);
or UO_411 (O_411,N_18099,N_18982);
nand UO_412 (O_412,N_17365,N_18009);
or UO_413 (O_413,N_18750,N_17878);
or UO_414 (O_414,N_17805,N_18841);
nor UO_415 (O_415,N_19596,N_16763);
nor UO_416 (O_416,N_18234,N_17633);
nor UO_417 (O_417,N_16652,N_18093);
and UO_418 (O_418,N_18617,N_19860);
and UO_419 (O_419,N_17465,N_17657);
or UO_420 (O_420,N_19061,N_18528);
and UO_421 (O_421,N_17064,N_16151);
and UO_422 (O_422,N_17772,N_19645);
or UO_423 (O_423,N_19060,N_18261);
xor UO_424 (O_424,N_17037,N_18599);
nor UO_425 (O_425,N_18777,N_19674);
and UO_426 (O_426,N_16633,N_17428);
nand UO_427 (O_427,N_16333,N_16295);
nor UO_428 (O_428,N_16168,N_19051);
or UO_429 (O_429,N_17122,N_19220);
xor UO_430 (O_430,N_16823,N_19412);
nor UO_431 (O_431,N_19478,N_17144);
or UO_432 (O_432,N_19136,N_16115);
nand UO_433 (O_433,N_16120,N_17600);
and UO_434 (O_434,N_19152,N_18757);
xnor UO_435 (O_435,N_18512,N_19890);
and UO_436 (O_436,N_17331,N_17239);
or UO_437 (O_437,N_19318,N_19361);
nand UO_438 (O_438,N_17007,N_16104);
or UO_439 (O_439,N_19789,N_19855);
nand UO_440 (O_440,N_16340,N_16107);
nor UO_441 (O_441,N_16967,N_16813);
or UO_442 (O_442,N_16616,N_19959);
nand UO_443 (O_443,N_16313,N_19993);
or UO_444 (O_444,N_19366,N_18480);
and UO_445 (O_445,N_19120,N_17820);
nor UO_446 (O_446,N_16249,N_16675);
and UO_447 (O_447,N_17230,N_16913);
and UO_448 (O_448,N_18932,N_16877);
nor UO_449 (O_449,N_17948,N_19182);
or UO_450 (O_450,N_17680,N_16565);
or UO_451 (O_451,N_19428,N_17613);
or UO_452 (O_452,N_18465,N_18876);
or UO_453 (O_453,N_19196,N_19048);
nand UO_454 (O_454,N_19782,N_17588);
xnor UO_455 (O_455,N_18163,N_16319);
and UO_456 (O_456,N_17965,N_17877);
nor UO_457 (O_457,N_19904,N_18255);
or UO_458 (O_458,N_19241,N_19438);
and UO_459 (O_459,N_17827,N_18929);
nor UO_460 (O_460,N_19513,N_17748);
nor UO_461 (O_461,N_18022,N_16247);
xor UO_462 (O_462,N_17665,N_19894);
or UO_463 (O_463,N_17779,N_18471);
nor UO_464 (O_464,N_19099,N_16358);
or UO_465 (O_465,N_17027,N_19372);
nand UO_466 (O_466,N_19417,N_17008);
or UO_467 (O_467,N_18593,N_16640);
nand UO_468 (O_468,N_16074,N_17570);
and UO_469 (O_469,N_16803,N_18715);
and UO_470 (O_470,N_18726,N_17330);
nand UO_471 (O_471,N_18989,N_16359);
xnor UO_472 (O_472,N_16059,N_17299);
and UO_473 (O_473,N_16995,N_16322);
nor UO_474 (O_474,N_19516,N_19429);
nor UO_475 (O_475,N_16958,N_19177);
xor UO_476 (O_476,N_18223,N_19277);
nor UO_477 (O_477,N_17841,N_19092);
or UO_478 (O_478,N_17051,N_16193);
nand UO_479 (O_479,N_18436,N_18540);
nor UO_480 (O_480,N_16316,N_19263);
and UO_481 (O_481,N_19600,N_18657);
nand UO_482 (O_482,N_19290,N_16676);
nor UO_483 (O_483,N_19649,N_19734);
nor UO_484 (O_484,N_18122,N_17236);
nor UO_485 (O_485,N_19029,N_17843);
and UO_486 (O_486,N_16227,N_18499);
nand UO_487 (O_487,N_18518,N_16931);
and UO_488 (O_488,N_19039,N_18978);
nor UO_489 (O_489,N_19605,N_17746);
nand UO_490 (O_490,N_17543,N_19327);
nand UO_491 (O_491,N_16084,N_16804);
nor UO_492 (O_492,N_19033,N_18535);
and UO_493 (O_493,N_18029,N_16292);
nor UO_494 (O_494,N_18966,N_16105);
nand UO_495 (O_495,N_18947,N_16374);
and UO_496 (O_496,N_16680,N_18847);
xor UO_497 (O_497,N_18425,N_18068);
or UO_498 (O_498,N_19468,N_19184);
nor UO_499 (O_499,N_18317,N_19973);
nor UO_500 (O_500,N_19948,N_18207);
or UO_501 (O_501,N_18276,N_19080);
xor UO_502 (O_502,N_18218,N_16978);
or UO_503 (O_503,N_16974,N_17998);
nor UO_504 (O_504,N_16200,N_18916);
or UO_505 (O_505,N_17211,N_19518);
or UO_506 (O_506,N_16833,N_16669);
or UO_507 (O_507,N_19268,N_18082);
nand UO_508 (O_508,N_19621,N_16642);
or UO_509 (O_509,N_17395,N_19560);
and UO_510 (O_510,N_18505,N_19901);
nor UO_511 (O_511,N_16417,N_18227);
nor UO_512 (O_512,N_19307,N_18357);
or UO_513 (O_513,N_18245,N_17823);
or UO_514 (O_514,N_19836,N_16766);
nor UO_515 (O_515,N_17243,N_17005);
nand UO_516 (O_516,N_17815,N_18270);
nor UO_517 (O_517,N_16752,N_16644);
nor UO_518 (O_518,N_17842,N_19608);
xnor UO_519 (O_519,N_17674,N_17811);
or UO_520 (O_520,N_17554,N_16095);
or UO_521 (O_521,N_17902,N_18615);
or UO_522 (O_522,N_18764,N_17855);
nand UO_523 (O_523,N_16905,N_17876);
and UO_524 (O_524,N_17572,N_18275);
nand UO_525 (O_525,N_19906,N_16613);
and UO_526 (O_526,N_16309,N_18486);
or UO_527 (O_527,N_17713,N_18334);
nand UO_528 (O_528,N_17648,N_19853);
nor UO_529 (O_529,N_17587,N_16879);
nor UO_530 (O_530,N_19469,N_18914);
and UO_531 (O_531,N_17666,N_17788);
nor UO_532 (O_532,N_18339,N_18118);
nand UO_533 (O_533,N_16557,N_17951);
and UO_534 (O_534,N_17728,N_18413);
nand UO_535 (O_535,N_16429,N_16271);
nand UO_536 (O_536,N_16469,N_19712);
and UO_537 (O_537,N_17874,N_18808);
nor UO_538 (O_538,N_16704,N_16591);
and UO_539 (O_539,N_16551,N_19348);
or UO_540 (O_540,N_19086,N_19296);
nand UO_541 (O_541,N_17983,N_16049);
nor UO_542 (O_542,N_19312,N_17975);
nand UO_543 (O_543,N_19320,N_17901);
nor UO_544 (O_544,N_18069,N_17949);
and UO_545 (O_545,N_17266,N_16320);
or UO_546 (O_546,N_16482,N_16442);
nand UO_547 (O_547,N_17832,N_19213);
nand UO_548 (O_548,N_16014,N_19895);
or UO_549 (O_549,N_17866,N_16472);
or UO_550 (O_550,N_17936,N_18696);
or UO_551 (O_551,N_16774,N_18866);
and UO_552 (O_552,N_19261,N_16242);
nor UO_553 (O_553,N_18226,N_18054);
or UO_554 (O_554,N_18132,N_17849);
nor UO_555 (O_555,N_18047,N_19126);
nand UO_556 (O_556,N_16975,N_16492);
or UO_557 (O_557,N_18171,N_18830);
nand UO_558 (O_558,N_17782,N_18080);
nand UO_559 (O_559,N_17723,N_17540);
nor UO_560 (O_560,N_17641,N_17845);
nand UO_561 (O_561,N_17671,N_18147);
nand UO_562 (O_562,N_19309,N_18694);
nor UO_563 (O_563,N_17444,N_19378);
nor UO_564 (O_564,N_16058,N_16383);
xor UO_565 (O_565,N_17627,N_19212);
or UO_566 (O_566,N_17334,N_16270);
nor UO_567 (O_567,N_19576,N_17614);
or UO_568 (O_568,N_18318,N_17133);
nand UO_569 (O_569,N_17168,N_16362);
nor UO_570 (O_570,N_18366,N_17537);
nor UO_571 (O_571,N_18249,N_19311);
nor UO_572 (O_572,N_16724,N_16179);
or UO_573 (O_573,N_17179,N_19233);
or UO_574 (O_574,N_16689,N_18872);
nand UO_575 (O_575,N_19422,N_19713);
or UO_576 (O_576,N_16634,N_16920);
nand UO_577 (O_577,N_17555,N_17489);
xnor UO_578 (O_578,N_18004,N_17853);
or UO_579 (O_579,N_18125,N_17598);
and UO_580 (O_580,N_17055,N_16520);
or UO_581 (O_581,N_16943,N_16854);
nor UO_582 (O_582,N_19838,N_18931);
nand UO_583 (O_583,N_18592,N_16420);
nor UO_584 (O_584,N_19358,N_18328);
nor UO_585 (O_585,N_17819,N_18065);
xor UO_586 (O_586,N_19298,N_18236);
nor UO_587 (O_587,N_17360,N_19185);
nand UO_588 (O_588,N_16307,N_18879);
nor UO_589 (O_589,N_19201,N_18697);
nand UO_590 (O_590,N_18071,N_17569);
and UO_591 (O_591,N_16770,N_17054);
nand UO_592 (O_592,N_18892,N_18375);
or UO_593 (O_593,N_16101,N_18404);
nand UO_594 (O_594,N_18521,N_18558);
nor UO_595 (O_595,N_18679,N_16529);
and UO_596 (O_596,N_16283,N_16893);
nand UO_597 (O_597,N_17529,N_18511);
or UO_598 (O_598,N_17106,N_17019);
or UO_599 (O_599,N_17014,N_18759);
nor UO_600 (O_600,N_18813,N_19760);
and UO_601 (O_601,N_17957,N_16667);
or UO_602 (O_602,N_18791,N_16786);
nand UO_603 (O_603,N_16138,N_18494);
or UO_604 (O_604,N_17527,N_18312);
or UO_605 (O_605,N_17332,N_19672);
nand UO_606 (O_606,N_19382,N_16175);
xnor UO_607 (O_607,N_19515,N_18837);
nor UO_608 (O_608,N_18700,N_17386);
and UO_609 (O_609,N_17860,N_19285);
nand UO_610 (O_610,N_16518,N_18386);
and UO_611 (O_611,N_16743,N_18596);
or UO_612 (O_612,N_17897,N_18348);
or UO_613 (O_613,N_19831,N_18482);
or UO_614 (O_614,N_16544,N_17617);
nand UO_615 (O_615,N_17921,N_19000);
nand UO_616 (O_616,N_19254,N_18170);
and UO_617 (O_617,N_17661,N_17375);
or UO_618 (O_618,N_19733,N_17622);
xnor UO_619 (O_619,N_18565,N_16448);
nor UO_620 (O_620,N_18968,N_19194);
or UO_621 (O_621,N_18579,N_17582);
or UO_622 (O_622,N_19132,N_16747);
or UO_623 (O_623,N_18095,N_18863);
nor UO_624 (O_624,N_19334,N_18620);
nand UO_625 (O_625,N_18705,N_17440);
or UO_626 (O_626,N_19976,N_16032);
or UO_627 (O_627,N_16881,N_17150);
xor UO_628 (O_628,N_17676,N_17914);
and UO_629 (O_629,N_16471,N_16462);
nor UO_630 (O_630,N_19567,N_18933);
nor UO_631 (O_631,N_19673,N_18821);
nor UO_632 (O_632,N_17808,N_19408);
or UO_633 (O_633,N_19661,N_17296);
nand UO_634 (O_634,N_19304,N_18416);
nand UO_635 (O_635,N_16812,N_17393);
and UO_636 (O_636,N_16596,N_19650);
or UO_637 (O_637,N_18393,N_16435);
and UO_638 (O_638,N_16338,N_17442);
nand UO_639 (O_639,N_16553,N_17775);
or UO_640 (O_640,N_19763,N_17340);
or UO_641 (O_641,N_18526,N_16922);
or UO_642 (O_642,N_19291,N_18603);
nor UO_643 (O_643,N_17594,N_18571);
nand UO_644 (O_644,N_18554,N_19595);
nand UO_645 (O_645,N_17161,N_16830);
or UO_646 (O_646,N_19465,N_16713);
and UO_647 (O_647,N_19587,N_19084);
nand UO_648 (O_648,N_19708,N_19197);
and UO_649 (O_649,N_18016,N_19511);
nor UO_650 (O_650,N_16860,N_17167);
or UO_651 (O_651,N_18476,N_19982);
nand UO_652 (O_652,N_16932,N_16018);
and UO_653 (O_653,N_18908,N_17655);
xor UO_654 (O_654,N_18846,N_17040);
nor UO_655 (O_655,N_18857,N_19878);
or UO_656 (O_656,N_16348,N_17291);
or UO_657 (O_657,N_19950,N_19905);
or UO_658 (O_658,N_18698,N_19236);
or UO_659 (O_659,N_18037,N_16369);
nor UO_660 (O_660,N_17565,N_18917);
and UO_661 (O_661,N_17021,N_17438);
nand UO_662 (O_662,N_19556,N_19295);
nor UO_663 (O_663,N_16198,N_18186);
nor UO_664 (O_664,N_16543,N_17116);
or UO_665 (O_665,N_19380,N_18400);
nand UO_666 (O_666,N_17532,N_16719);
or UO_667 (O_667,N_17306,N_17612);
nor UO_668 (O_668,N_16092,N_17896);
nor UO_669 (O_669,N_19071,N_18860);
or UO_670 (O_670,N_16599,N_17036);
or UO_671 (O_671,N_17926,N_16020);
or UO_672 (O_672,N_19816,N_19971);
nand UO_673 (O_673,N_19539,N_18607);
nor UO_674 (O_674,N_19828,N_18869);
or UO_675 (O_675,N_16000,N_16452);
or UO_676 (O_676,N_18305,N_19014);
and UO_677 (O_677,N_18258,N_19364);
nor UO_678 (O_678,N_16425,N_19389);
or UO_679 (O_679,N_19998,N_16614);
nand UO_680 (O_680,N_16332,N_16887);
and UO_681 (O_681,N_18426,N_18802);
and UO_682 (O_682,N_19682,N_18377);
or UO_683 (O_683,N_17319,N_16282);
or UO_684 (O_684,N_17813,N_18654);
nand UO_685 (O_685,N_16758,N_17213);
nor UO_686 (O_686,N_18272,N_17378);
nor UO_687 (O_687,N_18997,N_16904);
and UO_688 (O_688,N_19418,N_18306);
or UO_689 (O_689,N_18980,N_16844);
and UO_690 (O_690,N_18394,N_16457);
nor UO_691 (O_691,N_17210,N_17441);
xor UO_692 (O_692,N_17136,N_18290);
nand UO_693 (O_693,N_17183,N_16099);
and UO_694 (O_694,N_17604,N_18987);
or UO_695 (O_695,N_19753,N_18622);
nand UO_696 (O_696,N_17247,N_16167);
and UO_697 (O_697,N_19885,N_16122);
xor UO_698 (O_698,N_19994,N_16470);
nand UO_699 (O_699,N_18687,N_16971);
nor UO_700 (O_700,N_16134,N_18936);
nand UO_701 (O_701,N_17259,N_16371);
xor UO_702 (O_702,N_16329,N_19453);
nand UO_703 (O_703,N_17002,N_17944);
and UO_704 (O_704,N_18843,N_19575);
nor UO_705 (O_705,N_16664,N_17504);
xnor UO_706 (O_706,N_16396,N_17826);
nand UO_707 (O_707,N_17417,N_19617);
or UO_708 (O_708,N_16278,N_17033);
nor UO_709 (O_709,N_19660,N_18161);
and UO_710 (O_710,N_19772,N_16851);
or UO_711 (O_711,N_17485,N_18205);
nor UO_712 (O_712,N_18352,N_17345);
or UO_713 (O_713,N_19395,N_19922);
and UO_714 (O_714,N_17682,N_16558);
or UO_715 (O_715,N_17634,N_16658);
and UO_716 (O_716,N_19972,N_16413);
nor UO_717 (O_717,N_16220,N_18993);
nand UO_718 (O_718,N_17714,N_16566);
and UO_719 (O_719,N_16155,N_19267);
nand UO_720 (O_720,N_16917,N_16706);
nand UO_721 (O_721,N_17882,N_16121);
and UO_722 (O_722,N_17954,N_17856);
xnor UO_723 (O_723,N_17447,N_17162);
and UO_724 (O_724,N_19769,N_18051);
and UO_725 (O_725,N_19004,N_17273);
nand UO_726 (O_726,N_16447,N_17763);
and UO_727 (O_727,N_18214,N_16892);
or UO_728 (O_728,N_16009,N_17864);
and UO_729 (O_729,N_18935,N_17804);
xor UO_730 (O_730,N_17389,N_19388);
xnor UO_731 (O_731,N_16896,N_17545);
nor UO_732 (O_732,N_19329,N_17462);
nand UO_733 (O_733,N_19440,N_19123);
or UO_734 (O_734,N_16815,N_18343);
and UO_735 (O_735,N_18533,N_19915);
or UO_736 (O_736,N_17501,N_17430);
and UO_737 (O_737,N_16342,N_18153);
xnor UO_738 (O_738,N_17640,N_19392);
xnor UO_739 (O_739,N_16089,N_19636);
and UO_740 (O_740,N_17859,N_17774);
or UO_741 (O_741,N_19848,N_16147);
and UO_742 (O_742,N_16843,N_16346);
xor UO_743 (O_743,N_16903,N_19147);
or UO_744 (O_744,N_19953,N_19938);
or UO_745 (O_745,N_17203,N_17105);
nand UO_746 (O_746,N_18692,N_19481);
nand UO_747 (O_747,N_16454,N_16349);
and UO_748 (O_748,N_17404,N_19657);
nand UO_749 (O_749,N_18024,N_17789);
nand UO_750 (O_750,N_16712,N_18286);
nor UO_751 (O_751,N_18320,N_17262);
nor UO_752 (O_752,N_16114,N_18260);
nor UO_753 (O_753,N_16156,N_16477);
and UO_754 (O_754,N_16164,N_16979);
or UO_755 (O_755,N_19191,N_16441);
xor UO_756 (O_756,N_16955,N_16343);
nor UO_757 (O_757,N_19371,N_19238);
or UO_758 (O_758,N_18466,N_16570);
xnor UO_759 (O_759,N_18189,N_17097);
and UO_760 (O_760,N_17492,N_18299);
nor UO_761 (O_761,N_18280,N_19871);
nand UO_762 (O_762,N_18349,N_16499);
or UO_763 (O_763,N_18672,N_19514);
nand UO_764 (O_764,N_19563,N_18451);
nand UO_765 (O_765,N_18444,N_18828);
or UO_766 (O_766,N_16357,N_18862);
nor UO_767 (O_767,N_16415,N_16228);
nand UO_768 (O_768,N_19755,N_18259);
nand UO_769 (O_769,N_17084,N_17422);
nand UO_770 (O_770,N_19016,N_16716);
or UO_771 (O_771,N_19920,N_17863);
or UO_772 (O_772,N_16368,N_17705);
or UO_773 (O_773,N_17371,N_19707);
nor UO_774 (O_774,N_19025,N_18942);
nor UO_775 (O_775,N_19503,N_18129);
and UO_776 (O_776,N_16862,N_17420);
or UO_777 (O_777,N_16481,N_16305);
nand UO_778 (O_778,N_19219,N_18974);
and UO_779 (O_779,N_17847,N_16985);
nor UO_780 (O_780,N_18141,N_16880);
or UO_781 (O_781,N_18504,N_18943);
and UO_782 (O_782,N_19336,N_16690);
or UO_783 (O_783,N_18463,N_17708);
or UO_784 (O_784,N_16852,N_17802);
or UO_785 (O_785,N_18415,N_19955);
or UO_786 (O_786,N_17443,N_17357);
or UO_787 (O_787,N_17890,N_19049);
nand UO_788 (O_788,N_16078,N_16431);
and UO_789 (O_789,N_16426,N_19359);
nand UO_790 (O_790,N_18159,N_16818);
or UO_791 (O_791,N_17223,N_18239);
nor UO_792 (O_792,N_17437,N_19113);
nand UO_793 (O_793,N_17621,N_18142);
and UO_794 (O_794,N_16401,N_17316);
or UO_795 (O_795,N_17274,N_16173);
nor UO_796 (O_796,N_18810,N_19625);
nand UO_797 (O_797,N_18484,N_19690);
or UO_798 (O_798,N_17494,N_16749);
nor UO_799 (O_799,N_19774,N_18812);
nand UO_800 (O_800,N_18327,N_17962);
nand UO_801 (O_801,N_17946,N_17382);
and UO_802 (O_802,N_16526,N_19175);
and UO_803 (O_803,N_17762,N_19602);
and UO_804 (O_804,N_16192,N_17956);
and UO_805 (O_805,N_18313,N_19777);
nand UO_806 (O_806,N_16777,N_18457);
xnor UO_807 (O_807,N_17076,N_19654);
and UO_808 (O_808,N_16507,N_18884);
and UO_809 (O_809,N_17309,N_17260);
or UO_810 (O_810,N_17968,N_17401);
xnor UO_811 (O_811,N_17477,N_16710);
and UO_812 (O_812,N_16110,N_18743);
or UO_813 (O_813,N_19669,N_16022);
nand UO_814 (O_814,N_19824,N_17396);
xnor UO_815 (O_815,N_18994,N_19186);
and UO_816 (O_816,N_17071,N_19081);
nor UO_817 (O_817,N_19215,N_17377);
or UO_818 (O_818,N_18723,N_17905);
nand UO_819 (O_819,N_18021,N_19536);
or UO_820 (O_820,N_16508,N_19804);
or UO_821 (O_821,N_19540,N_19554);
nor UO_822 (O_822,N_18623,N_19257);
nand UO_823 (O_823,N_16373,N_17329);
nand UO_824 (O_824,N_19506,N_18067);
or UO_825 (O_825,N_17484,N_18253);
and UO_826 (O_826,N_19121,N_19640);
and UO_827 (O_827,N_18577,N_17045);
nand UO_828 (O_828,N_17445,N_18217);
or UO_829 (O_829,N_19530,N_16871);
and UO_830 (O_830,N_16067,N_19356);
or UO_831 (O_831,N_17736,N_16910);
nor UO_832 (O_832,N_19074,N_17776);
and UO_833 (O_833,N_17451,N_18784);
nand UO_834 (O_834,N_16598,N_16744);
nand UO_835 (O_835,N_16071,N_19803);
and UO_836 (O_836,N_16514,N_16952);
nor UO_837 (O_837,N_19779,N_19812);
nor UO_838 (O_838,N_18381,N_18379);
or UO_839 (O_839,N_18296,N_18373);
or UO_840 (O_840,N_19821,N_16873);
nor UO_841 (O_841,N_19999,N_17681);
xnor UO_842 (O_842,N_16512,N_18235);
nor UO_843 (O_843,N_16139,N_16160);
or UO_844 (O_844,N_17777,N_18613);
nor UO_845 (O_845,N_17277,N_16256);
nand UO_846 (O_846,N_19725,N_18428);
and UO_847 (O_847,N_18703,N_16272);
and UO_848 (O_848,N_17127,N_18992);
nand UO_849 (O_849,N_17952,N_17216);
nor UO_850 (O_850,N_18078,N_18854);
or UO_851 (O_851,N_17088,N_16334);
nand UO_852 (O_852,N_16294,N_18097);
xor UO_853 (O_853,N_18768,N_17624);
and UO_854 (O_854,N_17615,N_17228);
and UO_855 (O_855,N_16891,N_17978);
nand UO_856 (O_856,N_16419,N_16898);
nor UO_857 (O_857,N_19303,N_16181);
or UO_858 (O_858,N_18669,N_16593);
and UO_859 (O_859,N_17751,N_17020);
nand UO_860 (O_860,N_17658,N_19840);
nor UO_861 (O_861,N_17693,N_17999);
nand UO_862 (O_862,N_19227,N_17656);
and UO_863 (O_863,N_19523,N_19432);
and UO_864 (O_864,N_18695,N_18148);
nand UO_865 (O_865,N_19032,N_19163);
nor UO_866 (O_866,N_16982,N_17563);
and UO_867 (O_867,N_16714,N_19474);
or UO_868 (O_868,N_18302,N_17498);
or UO_869 (O_869,N_18031,N_17653);
xor UO_870 (O_870,N_17502,N_16946);
nand UO_871 (O_871,N_17589,N_18581);
nor UO_872 (O_872,N_19775,N_19626);
and UO_873 (O_873,N_19190,N_18832);
xor UO_874 (O_874,N_18365,N_19573);
nand UO_875 (O_875,N_17348,N_19902);
or UO_876 (O_876,N_18015,N_19765);
nand UO_877 (O_877,N_17523,N_19495);
nand UO_878 (O_878,N_16509,N_19974);
nand UO_879 (O_879,N_18005,N_17709);
or UO_880 (O_880,N_17741,N_16993);
or UO_881 (O_881,N_18111,N_18209);
and UO_882 (O_882,N_17198,N_16950);
nor UO_883 (O_883,N_16510,N_17250);
and UO_884 (O_884,N_18384,N_16405);
nand UO_885 (O_885,N_18594,N_18606);
nand UO_886 (O_886,N_16350,N_16912);
or UO_887 (O_887,N_18545,N_16406);
or UO_888 (O_888,N_16250,N_19486);
nand UO_889 (O_889,N_19718,N_16458);
or UO_890 (O_890,N_16407,N_16308);
xnor UO_891 (O_891,N_19732,N_18944);
and UO_892 (O_892,N_17970,N_17269);
nor UO_893 (O_893,N_17513,N_16627);
nor UO_894 (O_894,N_18070,N_17955);
nand UO_895 (O_895,N_16637,N_16890);
and UO_896 (O_896,N_16708,N_19479);
and UO_897 (O_897,N_18729,N_19819);
nand UO_898 (O_898,N_19425,N_18089);
or UO_899 (O_899,N_16533,N_17987);
nor UO_900 (O_900,N_19226,N_18835);
or UO_901 (O_901,N_17190,N_18332);
and UO_902 (O_902,N_19160,N_16523);
and UO_903 (O_903,N_17364,N_16806);
or UO_904 (O_904,N_17031,N_18291);
nor UO_905 (O_905,N_19271,N_17351);
nand UO_906 (O_906,N_18506,N_16622);
and UO_907 (O_907,N_16473,N_17405);
and UO_908 (O_908,N_17984,N_19929);
xnor UO_909 (O_909,N_16800,N_19030);
nand UO_910 (O_910,N_19992,N_16864);
nand UO_911 (O_911,N_19442,N_17801);
nand UO_912 (O_912,N_19040,N_19492);
xor UO_913 (O_913,N_16934,N_16692);
nor UO_914 (O_914,N_17892,N_18887);
nor UO_915 (O_915,N_19193,N_19253);
nand UO_916 (O_916,N_19736,N_16792);
nor UO_917 (O_917,N_17346,N_16540);
and UO_918 (O_918,N_19164,N_17608);
or UO_919 (O_919,N_17188,N_17852);
and UO_920 (O_920,N_19210,N_19670);
or UO_921 (O_921,N_19884,N_16194);
nand UO_922 (O_922,N_18307,N_16846);
nor UO_923 (O_923,N_19211,N_19475);
nor UO_924 (O_924,N_16336,N_19727);
xnor UO_925 (O_925,N_17909,N_18447);
nor UO_926 (O_926,N_17760,N_16484);
or UO_927 (O_927,N_17686,N_16840);
or UO_928 (O_928,N_16780,N_17013);
nand UO_929 (O_929,N_16767,N_19541);
xnor UO_930 (O_930,N_18803,N_19711);
or UO_931 (O_931,N_17321,N_18651);
nor UO_932 (O_932,N_16446,N_19472);
xor UO_933 (O_933,N_17931,N_17796);
nor UO_934 (O_934,N_19528,N_18042);
and UO_935 (O_935,N_16306,N_16129);
nand UO_936 (O_936,N_16550,N_19963);
and UO_937 (O_937,N_17564,N_17794);
nor UO_938 (O_938,N_18454,N_18557);
nand UO_939 (O_939,N_19485,N_18910);
nand UO_940 (O_940,N_18073,N_16467);
nand UO_941 (O_941,N_16050,N_16775);
and UO_942 (O_942,N_19749,N_17895);
or UO_943 (O_943,N_16693,N_17062);
nor UO_944 (O_944,N_18199,N_17493);
and UO_945 (O_945,N_19606,N_18461);
nor UO_946 (O_946,N_16146,N_16279);
and UO_947 (O_947,N_18714,N_16648);
nand UO_948 (O_948,N_19232,N_17110);
nor UO_949 (O_949,N_16177,N_17716);
and UO_950 (O_950,N_17180,N_16990);
or UO_951 (O_951,N_16569,N_18839);
and UO_952 (O_952,N_18045,N_19205);
nand UO_953 (O_953,N_16874,N_18595);
nand UO_954 (O_954,N_17687,N_16375);
xor UO_955 (O_955,N_18508,N_18060);
nor UO_956 (O_956,N_19666,N_16042);
nor UO_957 (O_957,N_17257,N_17356);
and UO_958 (O_958,N_18643,N_19908);
or UO_959 (O_959,N_19109,N_17997);
and UO_960 (O_960,N_16252,N_18848);
xor UO_961 (O_961,N_17336,N_18243);
and UO_962 (O_962,N_18520,N_17347);
or UO_963 (O_963,N_18983,N_19306);
xnor UO_964 (O_964,N_18157,N_18590);
and UO_965 (O_965,N_16645,N_17044);
and UO_966 (O_966,N_16205,N_18164);
nand UO_967 (O_967,N_16759,N_17318);
xnor UO_968 (O_968,N_19776,N_17043);
or UO_969 (O_969,N_18264,N_17053);
or UO_970 (O_970,N_17720,N_16082);
nand UO_971 (O_971,N_18269,N_16113);
or UO_972 (O_972,N_18420,N_19139);
and UO_973 (O_973,N_19206,N_17717);
and UO_974 (O_974,N_17506,N_18875);
and UO_975 (O_975,N_16376,N_19034);
or UO_976 (O_976,N_18772,N_18222);
nor UO_977 (O_977,N_18035,N_16817);
nand UO_978 (O_978,N_19409,N_16363);
nand UO_979 (O_979,N_17380,N_18941);
or UO_980 (O_980,N_19198,N_16035);
and UO_981 (O_981,N_18675,N_17868);
nor UO_982 (O_982,N_17632,N_16643);
nand UO_983 (O_983,N_16750,N_19857);
and UO_984 (O_984,N_19889,N_18367);
nor UO_985 (O_985,N_16490,N_18293);
nand UO_986 (O_986,N_19647,N_16190);
nor UO_987 (O_987,N_19243,N_19578);
and UO_988 (O_988,N_19001,N_19954);
and UO_989 (O_989,N_17452,N_16822);
nor UO_990 (O_990,N_19758,N_17985);
nand UO_991 (O_991,N_17469,N_19746);
nor UO_992 (O_992,N_19287,N_18321);
xor UO_993 (O_993,N_18845,N_18228);
and UO_994 (O_994,N_18552,N_17456);
or UO_995 (O_995,N_17848,N_18894);
nand UO_996 (O_996,N_19909,N_17039);
or UO_997 (O_997,N_17991,N_16414);
nor UO_998 (O_998,N_18127,N_19370);
nor UO_999 (O_999,N_17784,N_18030);
nand UO_1000 (O_1000,N_18206,N_18281);
or UO_1001 (O_1001,N_17358,N_18483);
nand UO_1002 (O_1002,N_18138,N_18699);
and UO_1003 (O_1003,N_16848,N_19297);
or UO_1004 (O_1004,N_18437,N_18008);
nand UO_1005 (O_1005,N_17835,N_18474);
xnor UO_1006 (O_1006,N_16671,N_16260);
xor UO_1007 (O_1007,N_18556,N_17538);
nand UO_1008 (O_1008,N_17953,N_16226);
and UO_1009 (O_1009,N_18990,N_16211);
nor UO_1010 (O_1010,N_16184,N_18690);
or UO_1011 (O_1011,N_16577,N_16869);
and UO_1012 (O_1012,N_19079,N_16753);
nor UO_1013 (O_1013,N_16240,N_18783);
or UO_1014 (O_1014,N_17454,N_18516);
and UO_1015 (O_1015,N_16427,N_17458);
or UO_1016 (O_1016,N_19265,N_18733);
and UO_1017 (O_1017,N_17061,N_19286);
and UO_1018 (O_1018,N_16918,N_16157);
nand UO_1019 (O_1019,N_18440,N_19314);
and UO_1020 (O_1020,N_18749,N_19912);
nand UO_1021 (O_1021,N_16545,N_19877);
nor UO_1022 (O_1022,N_18977,N_16755);
and UO_1023 (O_1023,N_16628,N_16412);
xor UO_1024 (O_1024,N_16290,N_18262);
nand UO_1025 (O_1025,N_16456,N_18642);
nand UO_1026 (O_1026,N_18361,N_18175);
or UO_1027 (O_1027,N_19924,N_17012);
xnor UO_1028 (O_1028,N_17280,N_17673);
and UO_1029 (O_1029,N_16268,N_16820);
nor UO_1030 (O_1030,N_17511,N_19851);
or UO_1031 (O_1031,N_18794,N_18949);
nand UO_1032 (O_1032,N_17320,N_18685);
nor UO_1033 (O_1033,N_19130,N_17433);
nor UO_1034 (O_1034,N_19288,N_17958);
or UO_1035 (O_1035,N_19678,N_17719);
and UO_1036 (O_1036,N_16746,N_19990);
or UO_1037 (O_1037,N_17268,N_16395);
xnor UO_1038 (O_1038,N_18541,N_19592);
nor UO_1039 (O_1039,N_19115,N_17328);
and UO_1040 (O_1040,N_17754,N_17379);
or UO_1041 (O_1041,N_17994,N_19278);
and UO_1042 (O_1042,N_19204,N_17181);
or UO_1043 (O_1043,N_19326,N_16855);
and UO_1044 (O_1044,N_18507,N_16051);
nor UO_1045 (O_1045,N_18475,N_19002);
nand UO_1046 (O_1046,N_17068,N_19101);
and UO_1047 (O_1047,N_19133,N_16301);
and UO_1048 (O_1048,N_19856,N_19338);
and UO_1049 (O_1049,N_16355,N_16259);
or UO_1050 (O_1050,N_19134,N_17973);
and UO_1051 (O_1051,N_18618,N_16300);
nor UO_1052 (O_1052,N_19349,N_16723);
and UO_1053 (O_1053,N_16923,N_19489);
or UO_1054 (O_1054,N_17164,N_18954);
nor UO_1055 (O_1055,N_19652,N_16836);
nand UO_1056 (O_1056,N_19762,N_19362);
and UO_1057 (O_1057,N_19761,N_16548);
or UO_1058 (O_1058,N_19124,N_18144);
or UO_1059 (O_1059,N_17918,N_16001);
xor UO_1060 (O_1060,N_16816,N_19543);
nor UO_1061 (O_1061,N_17986,N_16748);
nor UO_1062 (O_1062,N_18333,N_19671);
or UO_1063 (O_1063,N_19882,N_19701);
and UO_1064 (O_1064,N_18597,N_17818);
xor UO_1065 (O_1065,N_19519,N_16232);
nand UO_1066 (O_1066,N_16849,N_19010);
or UO_1067 (O_1067,N_18419,N_16036);
nor UO_1068 (O_1068,N_17374,N_16438);
and UO_1069 (O_1069,N_18755,N_16609);
nor UO_1070 (O_1070,N_18282,N_17231);
nor UO_1071 (O_1071,N_18452,N_16799);
nand UO_1072 (O_1072,N_16531,N_16040);
nor UO_1073 (O_1073,N_19694,N_19747);
nor UO_1074 (O_1074,N_18981,N_19754);
nand UO_1075 (O_1075,N_18322,N_17727);
and UO_1076 (O_1076,N_18450,N_18922);
and UO_1077 (O_1077,N_18003,N_17178);
or UO_1078 (O_1078,N_18771,N_16453);
nand UO_1079 (O_1079,N_19616,N_18676);
and UO_1080 (O_1080,N_18731,N_18886);
and UO_1081 (O_1081,N_19301,N_19817);
or UO_1082 (O_1082,N_17739,N_19452);
nor UO_1083 (O_1083,N_17932,N_19064);
or UO_1084 (O_1084,N_16907,N_18338);
nand UO_1085 (O_1085,N_18017,N_18530);
and UO_1086 (O_1086,N_19138,N_16195);
or UO_1087 (O_1087,N_16273,N_16605);
nor UO_1088 (O_1088,N_16498,N_19704);
nand UO_1089 (O_1089,N_18912,N_16882);
nand UO_1090 (O_1090,N_17034,N_18179);
nand UO_1091 (O_1091,N_19719,N_17817);
nand UO_1092 (O_1092,N_16298,N_17237);
nand UO_1093 (O_1093,N_17186,N_16326);
nand UO_1094 (O_1094,N_16574,N_17388);
or UO_1095 (O_1095,N_18336,N_16280);
xnor UO_1096 (O_1096,N_16180,N_18680);
and UO_1097 (O_1097,N_16635,N_18789);
and UO_1098 (O_1098,N_18074,N_17304);
or UO_1099 (O_1099,N_16511,N_18090);
or UO_1100 (O_1100,N_19968,N_18827);
nand UO_1101 (O_1101,N_17668,N_16465);
nand UO_1102 (O_1102,N_18973,N_17561);
nand UO_1103 (O_1103,N_19624,N_17629);
and UO_1104 (O_1104,N_19548,N_16581);
xor UO_1105 (O_1105,N_18958,N_19058);
and UO_1106 (O_1106,N_18300,N_18850);
xor UO_1107 (O_1107,N_16549,N_18739);
nand UO_1108 (O_1108,N_18050,N_17355);
xor UO_1109 (O_1109,N_17214,N_18959);
nor UO_1110 (O_1110,N_16459,N_19521);
and UO_1111 (O_1111,N_16408,N_18020);
nor UO_1112 (O_1112,N_17056,N_18706);
and UO_1113 (O_1113,N_19813,N_17047);
or UO_1114 (O_1114,N_16019,N_18570);
and UO_1115 (O_1115,N_17894,N_16201);
xor UO_1116 (O_1116,N_18895,N_19445);
nand UO_1117 (O_1117,N_17678,N_18231);
nor UO_1118 (O_1118,N_16318,N_16672);
or UO_1119 (O_1119,N_19221,N_16556);
or UO_1120 (O_1120,N_18284,N_18058);
nor UO_1121 (O_1121,N_18088,N_19339);
nand UO_1122 (O_1122,N_18049,N_18965);
or UO_1123 (O_1123,N_18213,N_17142);
nor UO_1124 (O_1124,N_19137,N_18105);
and UO_1125 (O_1125,N_18548,N_16954);
nand UO_1126 (O_1126,N_19351,N_17964);
nor UO_1127 (O_1127,N_17113,N_17765);
nand UO_1128 (O_1128,N_17664,N_19814);
or UO_1129 (O_1129,N_18162,N_18006);
and UO_1130 (O_1130,N_19294,N_17342);
or UO_1131 (O_1131,N_19083,N_18650);
nor UO_1132 (O_1132,N_18277,N_18192);
or UO_1133 (O_1133,N_18174,N_17455);
nor UO_1134 (O_1134,N_18244,N_19483);
or UO_1135 (O_1135,N_16152,N_19951);
nor UO_1136 (O_1136,N_19171,N_16171);
or UO_1137 (O_1137,N_16666,N_19424);
nand UO_1138 (O_1138,N_17474,N_16657);
nand UO_1139 (O_1139,N_19500,N_19140);
and UO_1140 (O_1140,N_17220,N_18621);
and UO_1141 (O_1141,N_19482,N_19764);
or UO_1142 (O_1142,N_16203,N_17798);
nand UO_1143 (O_1143,N_18661,N_19116);
nand UO_1144 (O_1144,N_18018,N_19710);
or UO_1145 (O_1145,N_16372,N_19869);
and UO_1146 (O_1146,N_16403,N_19405);
nor UO_1147 (O_1147,N_17065,N_19087);
nand UO_1148 (O_1148,N_18188,N_17831);
or UO_1149 (O_1149,N_19863,N_17131);
or UO_1150 (O_1150,N_16404,N_19984);
nor UO_1151 (O_1151,N_16829,N_17095);
or UO_1152 (O_1152,N_19377,N_16197);
xnor UO_1153 (O_1153,N_19964,N_17471);
nand UO_1154 (O_1154,N_18711,N_16027);
xor UO_1155 (O_1155,N_17980,N_16729);
nor UO_1156 (O_1156,N_16580,N_17025);
and UO_1157 (O_1157,N_19784,N_17548);
nor UO_1158 (O_1158,N_17972,N_17562);
nand UO_1159 (O_1159,N_18693,N_19553);
nand UO_1160 (O_1160,N_19179,N_18053);
and UO_1161 (O_1161,N_17771,N_17919);
xnor UO_1162 (O_1162,N_18139,N_16886);
and UO_1163 (O_1163,N_16057,N_18407);
xnor UO_1164 (O_1164,N_17639,N_17145);
nor UO_1165 (O_1165,N_16026,N_19689);
nor UO_1166 (O_1166,N_16796,N_18817);
or UO_1167 (O_1167,N_17935,N_17464);
or UO_1168 (O_1168,N_16150,N_16571);
or UO_1169 (O_1169,N_16478,N_16826);
and UO_1170 (O_1170,N_18330,N_16131);
nor UO_1171 (O_1171,N_16310,N_19217);
and UO_1172 (O_1172,N_19798,N_19571);
nand UO_1173 (O_1173,N_18640,N_18631);
and UO_1174 (O_1174,N_17520,N_17644);
nor UO_1175 (O_1175,N_18807,N_17224);
or UO_1176 (O_1176,N_17628,N_16517);
nand UO_1177 (O_1177,N_17176,N_16771);
or UO_1178 (O_1178,N_19052,N_19289);
nor UO_1179 (O_1179,N_17368,N_17251);
or UO_1180 (O_1180,N_16257,N_17711);
or UO_1181 (O_1181,N_19457,N_19538);
nand UO_1182 (O_1182,N_19903,N_19363);
nor UO_1183 (O_1183,N_19480,N_19793);
nand UO_1184 (O_1184,N_19659,N_16727);
xnor UO_1185 (O_1185,N_17967,N_18458);
and UO_1186 (O_1186,N_16575,N_16590);
and UO_1187 (O_1187,N_17750,N_19183);
nand UO_1188 (O_1188,N_19461,N_18001);
nand UO_1189 (O_1189,N_18986,N_17738);
nand UO_1190 (O_1190,N_18283,N_17766);
nand UO_1191 (O_1191,N_16424,N_18406);
or UO_1192 (O_1192,N_16186,N_17080);
nor UO_1193 (O_1193,N_19978,N_17836);
and UO_1194 (O_1194,N_18721,N_19943);
xnor UO_1195 (O_1195,N_17184,N_16969);
and UO_1196 (O_1196,N_19174,N_18040);
nand UO_1197 (O_1197,N_19091,N_16065);
and UO_1198 (O_1198,N_17637,N_19400);
nor UO_1199 (O_1199,N_17636,N_18000);
or UO_1200 (O_1200,N_16235,N_19321);
or UO_1201 (O_1201,N_16410,N_18576);
nand UO_1202 (O_1202,N_17312,N_19063);
and UO_1203 (O_1203,N_17208,N_19146);
xnor UO_1204 (O_1204,N_18976,N_19723);
nor UO_1205 (O_1205,N_18883,N_19410);
nand UO_1206 (O_1206,N_17583,N_18396);
nand UO_1207 (O_1207,N_17595,N_19648);
nor UO_1208 (O_1208,N_17576,N_19282);
or UO_1209 (O_1209,N_16832,N_18510);
and UO_1210 (O_1210,N_16007,N_16031);
xnor UO_1211 (O_1211,N_16795,N_16606);
nor UO_1212 (O_1212,N_16386,N_19637);
or UO_1213 (O_1213,N_16367,N_19491);
or UO_1214 (O_1214,N_18800,N_18409);
or UO_1215 (O_1215,N_18671,N_19416);
xor UO_1216 (O_1216,N_18871,N_19399);
nor UO_1217 (O_1217,N_19888,N_18586);
and UO_1218 (O_1218,N_17635,N_19641);
nor UO_1219 (O_1219,N_18674,N_17749);
nand UO_1220 (O_1220,N_16653,N_17689);
xnor UO_1221 (O_1221,N_17090,N_18897);
nand UO_1222 (O_1222,N_19668,N_19512);
or UO_1223 (O_1223,N_16977,N_17929);
or UO_1224 (O_1224,N_19875,N_16239);
nor UO_1225 (O_1225,N_19300,N_17333);
nand UO_1226 (O_1226,N_18112,N_18906);
or UO_1227 (O_1227,N_19622,N_19966);
or UO_1228 (O_1228,N_19012,N_19118);
and UO_1229 (O_1229,N_19807,N_17264);
nor UO_1230 (O_1230,N_18818,N_18589);
or UO_1231 (O_1231,N_17512,N_19699);
nor UO_1232 (O_1232,N_19085,N_16411);
nand UO_1233 (O_1233,N_17781,N_17884);
xor UO_1234 (O_1234,N_16140,N_19460);
or UO_1235 (O_1235,N_16016,N_17688);
xor UO_1236 (O_1236,N_19394,N_17579);
and UO_1237 (O_1237,N_19068,N_18560);
nor UO_1238 (O_1238,N_17690,N_17158);
or UO_1239 (O_1239,N_19433,N_16885);
or UO_1240 (O_1240,N_18044,N_19202);
and UO_1241 (O_1241,N_16698,N_16769);
nand UO_1242 (O_1242,N_16784,N_19944);
nor UO_1243 (O_1243,N_17960,N_19630);
nand UO_1244 (O_1244,N_16076,N_19683);
xnor UO_1245 (O_1245,N_16505,N_19117);
nor UO_1246 (O_1246,N_19208,N_17431);
nand UO_1247 (O_1247,N_19223,N_16808);
nor UO_1248 (O_1248,N_17412,N_19216);
nand UO_1249 (O_1249,N_16850,N_19488);
nor UO_1250 (O_1250,N_18387,N_19745);
nor UO_1251 (O_1251,N_18059,N_18779);
and UO_1252 (O_1252,N_17290,N_17276);
and UO_1253 (O_1253,N_19911,N_16687);
or UO_1254 (O_1254,N_16496,N_19629);
or UO_1255 (O_1255,N_17009,N_17233);
xnor UO_1256 (O_1256,N_18919,N_17283);
xnor UO_1257 (O_1257,N_17623,N_16810);
nor UO_1258 (O_1258,N_19720,N_18701);
nor UO_1259 (O_1259,N_18793,N_16870);
and UO_1260 (O_1260,N_18609,N_18355);
nor UO_1261 (O_1261,N_18424,N_18184);
nand UO_1262 (O_1262,N_16519,N_19722);
nand UO_1263 (O_1263,N_19933,N_17605);
nand UO_1264 (O_1264,N_19724,N_19985);
and UO_1265 (O_1265,N_17399,N_17862);
or UO_1266 (O_1266,N_16654,N_18991);
and UO_1267 (O_1267,N_19729,N_19750);
and UO_1268 (O_1268,N_16638,N_17234);
or UO_1269 (O_1269,N_19841,N_17503);
or UO_1270 (O_1270,N_18713,N_17175);
and UO_1271 (O_1271,N_18578,N_17692);
nand UO_1272 (O_1272,N_19018,N_17593);
nor UO_1273 (O_1273,N_17846,N_16630);
nand UO_1274 (O_1274,N_19565,N_16789);
nand UO_1275 (O_1275,N_16924,N_16902);
or UO_1276 (O_1276,N_19054,N_17913);
xnor UO_1277 (O_1277,N_17937,N_16263);
and UO_1278 (O_1278,N_17411,N_18055);
nand UO_1279 (O_1279,N_17117,N_18531);
nor UO_1280 (O_1280,N_16005,N_19082);
and UO_1281 (O_1281,N_18787,N_16668);
or UO_1282 (O_1282,N_18041,N_17659);
and UO_1283 (O_1283,N_16174,N_19611);
or UO_1284 (O_1284,N_16623,N_19716);
and UO_1285 (O_1285,N_18833,N_18950);
xnor UO_1286 (O_1286,N_16077,N_17488);
and UO_1287 (O_1287,N_19679,N_16996);
nor UO_1288 (O_1288,N_17821,N_18166);
nand UO_1289 (O_1289,N_18815,N_17609);
or UO_1290 (O_1290,N_18624,N_16959);
and UO_1291 (O_1291,N_17383,N_19038);
or UO_1292 (O_1292,N_16515,N_17660);
or UO_1293 (O_1293,N_18470,N_18627);
nor UO_1294 (O_1294,N_17419,N_19127);
nor UO_1295 (O_1295,N_17758,N_17619);
and UO_1296 (O_1296,N_18056,N_17400);
nor UO_1297 (O_1297,N_19631,N_18836);
nor UO_1298 (O_1298,N_17735,N_18666);
or UO_1299 (O_1299,N_18853,N_17620);
nor UO_1300 (O_1300,N_17992,N_18130);
xor UO_1301 (O_1301,N_18645,N_17669);
and UO_1302 (O_1302,N_18301,N_19780);
and UO_1303 (O_1303,N_18536,N_18709);
nand UO_1304 (O_1304,N_19053,N_19680);
and UO_1305 (O_1305,N_19688,N_16024);
nor UO_1306 (O_1306,N_17170,N_17825);
nand UO_1307 (O_1307,N_17085,N_19967);
or UO_1308 (O_1308,N_18564,N_17701);
or UO_1309 (O_1309,N_19604,N_19355);
xor UO_1310 (O_1310,N_18064,N_19252);
and UO_1311 (O_1311,N_18822,N_19487);
xnor UO_1312 (O_1312,N_16732,N_17349);
nand UO_1313 (O_1313,N_16494,N_18569);
xnor UO_1314 (O_1314,N_18023,N_16821);
nand UO_1315 (O_1315,N_16266,N_16636);
or UO_1316 (O_1316,N_17448,N_16111);
and UO_1317 (O_1317,N_17010,N_19946);
nor UO_1318 (O_1318,N_17151,N_18397);
or UO_1319 (O_1319,N_18100,N_19047);
and UO_1320 (O_1320,N_16783,N_16632);
and UO_1321 (O_1321,N_17961,N_17917);
nand UO_1322 (O_1322,N_18242,N_17129);
or UO_1323 (O_1323,N_19496,N_16163);
or UO_1324 (O_1324,N_17169,N_18608);
or UO_1325 (O_1325,N_17450,N_16717);
or UO_1326 (O_1326,N_17519,N_17557);
nor UO_1327 (O_1327,N_17883,N_18985);
or UO_1328 (O_1328,N_19003,N_19965);
or UO_1329 (O_1329,N_17424,N_19279);
or UO_1330 (O_1330,N_18468,N_16303);
and UO_1331 (O_1331,N_16819,N_17533);
nor UO_1332 (O_1332,N_16432,N_18292);
nand UO_1333 (O_1333,N_16006,N_18268);
and UO_1334 (O_1334,N_18939,N_17742);
nand UO_1335 (O_1335,N_19815,N_19102);
nor UO_1336 (O_1336,N_16956,N_18241);
nor UO_1337 (O_1337,N_17261,N_18742);
or UO_1338 (O_1338,N_19158,N_18668);
nand UO_1339 (O_1339,N_19357,N_16986);
and UO_1340 (O_1340,N_19940,N_19407);
and UO_1341 (O_1341,N_18371,N_18937);
nand UO_1342 (O_1342,N_18423,N_17786);
and UO_1343 (O_1343,N_17160,N_16576);
and UO_1344 (O_1344,N_16782,N_16207);
and UO_1345 (O_1345,N_16347,N_17229);
nor UO_1346 (O_1346,N_16901,N_17391);
xnor UO_1347 (O_1347,N_19266,N_16328);
nor UO_1348 (O_1348,N_16595,N_18238);
nand UO_1349 (O_1349,N_17590,N_19737);
and UO_1350 (O_1350,N_17288,N_18795);
nand UO_1351 (O_1351,N_16965,N_17202);
nor UO_1352 (O_1352,N_17979,N_17551);
nand UO_1353 (O_1353,N_19619,N_16961);
nand UO_1354 (O_1354,N_16541,N_18467);
or UO_1355 (O_1355,N_17885,N_18885);
and UO_1356 (O_1356,N_17873,N_16158);
nor UO_1357 (O_1357,N_16999,N_18498);
or UO_1358 (O_1358,N_19868,N_16683);
xnor UO_1359 (O_1359,N_18043,N_17058);
or UO_1360 (O_1360,N_17123,N_16736);
nor UO_1361 (O_1361,N_17463,N_19551);
or UO_1362 (O_1362,N_19979,N_17667);
xor UO_1363 (O_1363,N_19450,N_16381);
or UO_1364 (O_1364,N_19365,N_17925);
or UO_1365 (O_1365,N_19310,N_16154);
and UO_1366 (O_1366,N_16615,N_17703);
nor UO_1367 (O_1367,N_19192,N_17140);
xnor UO_1368 (O_1368,N_18081,N_18611);
or UO_1369 (O_1369,N_17524,N_18195);
and UO_1370 (O_1370,N_19231,N_18826);
or UO_1371 (O_1371,N_18390,N_16839);
nor UO_1372 (O_1372,N_16130,N_16603);
nand UO_1373 (O_1373,N_19744,N_19687);
nor UO_1374 (O_1374,N_19686,N_18326);
nand UO_1375 (O_1375,N_18859,N_17232);
or UO_1376 (O_1376,N_19633,N_19715);
nor UO_1377 (O_1377,N_19427,N_18477);
and UO_1378 (O_1378,N_19260,N_18653);
nand UO_1379 (O_1379,N_16740,N_16277);
nand UO_1380 (O_1380,N_17696,N_19655);
and UO_1381 (O_1381,N_18154,N_19684);
nand UO_1382 (O_1382,N_17209,N_16592);
nor UO_1383 (O_1383,N_19883,N_19439);
or UO_1384 (O_1384,N_19873,N_19089);
and UO_1385 (O_1385,N_17850,N_18414);
nor UO_1386 (O_1386,N_19810,N_16255);
nor UO_1387 (O_1387,N_19822,N_19961);
nand UO_1388 (O_1388,N_16327,N_19529);
nor UO_1389 (O_1389,N_16119,N_17083);
and UO_1390 (O_1390,N_19846,N_18448);
and UO_1391 (O_1391,N_17740,N_17302);
and UO_1392 (O_1392,N_16734,N_18345);
nand UO_1393 (O_1393,N_18588,N_18114);
and UO_1394 (O_1394,N_18925,N_18110);
and UO_1395 (O_1395,N_19872,N_18873);
and UO_1396 (O_1396,N_18422,N_17601);
nand UO_1397 (O_1397,N_16847,N_17881);
nand UO_1398 (O_1398,N_16516,N_18344);
and UO_1399 (O_1399,N_18385,N_17585);
and UO_1400 (O_1400,N_17483,N_16244);
and UO_1401 (O_1401,N_18574,N_16930);
nor UO_1402 (O_1402,N_19709,N_18823);
nor UO_1403 (O_1403,N_19534,N_17851);
nand UO_1404 (O_1404,N_17119,N_16894);
nor UO_1405 (O_1405,N_17712,N_16944);
and UO_1406 (O_1406,N_16052,N_16142);
nand UO_1407 (O_1407,N_16023,N_18198);
and UO_1408 (O_1408,N_17631,N_17081);
or UO_1409 (O_1409,N_17767,N_17976);
nand UO_1410 (O_1410,N_19406,N_19035);
and UO_1411 (O_1411,N_18193,N_17305);
and UO_1412 (O_1412,N_19414,N_16703);
nor UO_1413 (O_1413,N_18211,N_18200);
or UO_1414 (O_1414,N_16572,N_16365);
nand UO_1415 (O_1415,N_17449,N_18962);
and UO_1416 (O_1416,N_17694,N_16908);
nand UO_1417 (O_1417,N_17571,N_19623);
or UO_1418 (O_1418,N_18323,N_16828);
nor UO_1419 (O_1419,N_17415,N_16647);
or UO_1420 (O_1420,N_18429,N_17326);
xor UO_1421 (O_1421,N_19932,N_16262);
nand UO_1422 (O_1422,N_19077,N_17481);
xor UO_1423 (O_1423,N_17427,N_17770);
and UO_1424 (O_1424,N_18287,N_19677);
nor UO_1425 (O_1425,N_18378,N_18964);
xor UO_1426 (O_1426,N_16399,N_17791);
nand UO_1427 (O_1427,N_18928,N_18870);
or UO_1428 (O_1428,N_19387,N_19800);
or UO_1429 (O_1429,N_19021,N_17702);
or UO_1430 (O_1430,N_18104,N_16474);
nand UO_1431 (O_1431,N_17187,N_17470);
or UO_1432 (O_1432,N_16951,N_17910);
and UO_1433 (O_1433,N_16875,N_19008);
and UO_1434 (O_1434,N_16980,N_17875);
xor UO_1435 (O_1435,N_18431,N_17810);
nor UO_1436 (O_1436,N_16034,N_16370);
and UO_1437 (O_1437,N_18456,N_19222);
and UO_1438 (O_1438,N_19695,N_16761);
nor UO_1439 (O_1439,N_17107,N_18634);
nand UO_1440 (O_1440,N_16797,N_19413);
nor UO_1441 (O_1441,N_16108,N_17057);
xnor UO_1442 (O_1442,N_18532,N_17971);
nand UO_1443 (O_1443,N_19570,N_19157);
and UO_1444 (O_1444,N_16212,N_16064);
nor UO_1445 (O_1445,N_16720,N_17135);
nor UO_1446 (O_1446,N_17482,N_18781);
nand UO_1447 (O_1447,N_17691,N_17069);
nand UO_1448 (O_1448,N_19642,N_17397);
nand UO_1449 (O_1449,N_19023,N_16096);
and UO_1450 (O_1450,N_18956,N_16624);
nand UO_1451 (O_1451,N_17130,N_16584);
xor UO_1452 (O_1452,N_19770,N_16449);
or UO_1453 (O_1453,N_16062,N_17335);
nand UO_1454 (O_1454,N_18202,N_16219);
nor UO_1455 (O_1455,N_16973,N_18156);
and UO_1456 (O_1456,N_19262,N_19446);
xnor UO_1457 (O_1457,N_16612,N_18314);
and UO_1458 (O_1458,N_16221,N_17217);
nand UO_1459 (O_1459,N_17241,N_16223);
or UO_1460 (O_1460,N_17052,N_16254);
nand UO_1461 (O_1461,N_17204,N_17439);
and UO_1462 (O_1462,N_16159,N_17907);
nand UO_1463 (O_1463,N_19145,N_17934);
xor UO_1464 (O_1464,N_19834,N_18811);
and UO_1465 (O_1465,N_19156,N_18347);
nor UO_1466 (O_1466,N_16033,N_18019);
or UO_1467 (O_1467,N_18967,N_16677);
or UO_1468 (O_1468,N_17761,N_16601);
or UO_1469 (O_1469,N_19584,N_19627);
nor UO_1470 (O_1470,N_18988,N_17030);
nand UO_1471 (O_1471,N_17369,N_17497);
or UO_1472 (O_1472,N_19740,N_19056);
and UO_1473 (O_1473,N_17137,N_16331);
nor UO_1474 (O_1474,N_19073,N_17778);
or UO_1475 (O_1475,N_17947,N_17942);
or UO_1476 (O_1476,N_19292,N_19386);
nor UO_1477 (O_1477,N_19373,N_17651);
xor UO_1478 (O_1478,N_17478,N_19508);
or UO_1479 (O_1479,N_17111,N_18254);
nor UO_1480 (O_1480,N_19989,N_19276);
nand UO_1481 (O_1481,N_19207,N_19663);
or UO_1482 (O_1482,N_17300,N_17495);
and UO_1483 (O_1483,N_16867,N_18562);
nor UO_1484 (O_1484,N_19510,N_16655);
nor UO_1485 (O_1485,N_17003,N_17265);
or UO_1486 (O_1486,N_16552,N_18663);
nor UO_1487 (O_1487,N_16625,N_18443);
and UO_1488 (O_1488,N_16443,N_18842);
nor UO_1489 (O_1489,N_18605,N_16739);
or UO_1490 (O_1490,N_16987,N_17982);
nor UO_1491 (O_1491,N_18146,N_17645);
or UO_1492 (O_1492,N_17898,N_17647);
nor UO_1493 (O_1493,N_16112,N_17988);
nand UO_1494 (O_1494,N_19319,N_17141);
or UO_1495 (O_1495,N_16170,N_18517);
nand UO_1496 (O_1496,N_19275,N_17491);
and UO_1497 (O_1497,N_17521,N_16764);
nor UO_1498 (O_1498,N_18140,N_18232);
and UO_1499 (O_1499,N_19790,N_19705);
nand UO_1500 (O_1500,N_19067,N_16206);
xnor UO_1501 (O_1501,N_19818,N_16992);
nand UO_1502 (O_1502,N_16463,N_18309);
and UO_1503 (O_1503,N_16929,N_17287);
nor UO_1504 (O_1504,N_16807,N_19778);
or UO_1505 (O_1505,N_16191,N_16296);
or UO_1506 (O_1506,N_18639,N_16865);
xnor UO_1507 (O_1507,N_18575,N_18829);
xor UO_1508 (O_1508,N_16878,N_17311);
nor UO_1509 (O_1509,N_16937,N_17109);
nor UO_1510 (O_1510,N_18389,N_18285);
nand UO_1511 (O_1511,N_16236,N_16794);
nor UO_1512 (O_1512,N_18131,N_19997);
nor UO_1513 (O_1513,N_17816,N_18806);
or UO_1514 (O_1514,N_17366,N_16699);
and UO_1515 (O_1515,N_19093,N_16600);
nand UO_1516 (O_1516,N_16793,N_16582);
nand UO_1517 (O_1517,N_18410,N_19317);
nand UO_1518 (O_1518,N_16779,N_19832);
and UO_1519 (O_1519,N_19390,N_18844);
or UO_1520 (O_1520,N_18961,N_16083);
or UO_1521 (O_1521,N_18137,N_19865);
xnor UO_1522 (O_1522,N_18180,N_17414);
or UO_1523 (O_1523,N_17096,N_19607);
or UO_1524 (O_1524,N_16125,N_16087);
and UO_1525 (O_1525,N_19162,N_18745);
or UO_1526 (O_1526,N_19281,N_16440);
or UO_1527 (O_1527,N_18120,N_18274);
and UO_1528 (O_1528,N_17833,N_18905);
and UO_1529 (O_1529,N_16911,N_19981);
nor UO_1530 (O_1530,N_16196,N_18704);
nor UO_1531 (O_1531,N_19250,N_19794);
nor UO_1532 (O_1532,N_17238,N_18152);
and UO_1533 (O_1533,N_19957,N_16274);
and UO_1534 (O_1534,N_17026,N_19239);
and UO_1535 (O_1535,N_17726,N_19354);
and UO_1536 (O_1536,N_16631,N_19792);
and UO_1537 (O_1537,N_19542,N_17945);
nand UO_1538 (O_1538,N_18900,N_19240);
xor UO_1539 (O_1539,N_17806,N_17526);
xor UO_1540 (O_1540,N_17254,N_19858);
and UO_1541 (O_1541,N_19502,N_16072);
nor UO_1542 (O_1542,N_19552,N_17174);
nand UO_1543 (O_1543,N_16241,N_16814);
nor UO_1544 (O_1544,N_16534,N_17092);
nor UO_1545 (O_1545,N_16025,N_16530);
nand UO_1546 (O_1546,N_19826,N_17067);
or UO_1547 (O_1547,N_18720,N_16225);
nor UO_1548 (O_1548,N_18411,N_17996);
and UO_1549 (O_1549,N_17522,N_18430);
nand UO_1550 (O_1550,N_16696,N_17795);
nor UO_1551 (O_1551,N_18288,N_16895);
nand UO_1552 (O_1552,N_17518,N_17743);
nor UO_1553 (O_1553,N_17757,N_16960);
nor UO_1554 (O_1554,N_18864,N_19934);
nand UO_1555 (O_1555,N_19237,N_16966);
and UO_1556 (O_1556,N_17381,N_19050);
or UO_1557 (O_1557,N_19574,N_16276);
or UO_1558 (O_1558,N_18769,N_17530);
xnor UO_1559 (O_1559,N_17908,N_17024);
and UO_1560 (O_1560,N_18718,N_18316);
nand UO_1561 (O_1561,N_17154,N_17793);
and UO_1562 (O_1562,N_17768,N_16825);
xor UO_1563 (O_1563,N_17022,N_17977);
nand UO_1564 (O_1564,N_16098,N_17467);
xor UO_1565 (O_1565,N_19739,N_18628);
or UO_1566 (O_1566,N_18820,N_18909);
nor UO_1567 (O_1567,N_17473,N_19075);
or UO_1568 (O_1568,N_18598,N_17074);
or UO_1569 (O_1569,N_18481,N_18350);
nand UO_1570 (O_1570,N_16684,N_17574);
or UO_1571 (O_1571,N_17787,N_17476);
or UO_1572 (O_1572,N_16899,N_19806);
xor UO_1573 (O_1573,N_17363,N_19849);
and UO_1574 (O_1574,N_18107,N_17732);
nor UO_1575 (O_1575,N_18401,N_17541);
or UO_1576 (O_1576,N_18979,N_17773);
nand UO_1577 (O_1577,N_18340,N_19346);
nand UO_1578 (O_1578,N_17963,N_19728);
and UO_1579 (O_1579,N_19096,N_19402);
nand UO_1580 (O_1580,N_18647,N_17282);
nand UO_1581 (O_1581,N_17535,N_17016);
nand UO_1582 (O_1582,N_19768,N_18488);
and UO_1583 (O_1583,N_18688,N_17286);
nor UO_1584 (O_1584,N_17258,N_19367);
and UO_1585 (O_1585,N_16185,N_16011);
xnor UO_1586 (O_1586,N_17354,N_17809);
nor UO_1587 (O_1587,N_18453,N_17534);
and UO_1588 (O_1588,N_18464,N_18921);
nor UO_1589 (O_1589,N_17206,N_17436);
nor UO_1590 (O_1590,N_18656,N_18374);
xor UO_1591 (O_1591,N_17115,N_18881);
and UO_1592 (O_1592,N_19582,N_19499);
nand UO_1593 (O_1593,N_19702,N_18036);
nand UO_1594 (O_1594,N_16685,N_18641);
nand UO_1595 (O_1595,N_19795,N_16949);
nor UO_1596 (O_1596,N_16564,N_17432);
xnor UO_1597 (O_1597,N_18551,N_18057);
or UO_1598 (O_1598,N_19324,N_19055);
nor UO_1599 (O_1599,N_18117,N_16385);
and UO_1600 (O_1600,N_19910,N_17435);
nor UO_1601 (O_1601,N_19526,N_18882);
nand UO_1602 (O_1602,N_18446,N_16694);
or UO_1603 (O_1603,N_18266,N_18543);
nand UO_1604 (O_1604,N_18684,N_16012);
or UO_1605 (O_1605,N_19108,N_16998);
nand UO_1606 (O_1606,N_19917,N_16352);
nor UO_1607 (O_1607,N_18741,N_18648);
or UO_1608 (O_1608,N_19507,N_18804);
xnor UO_1609 (O_1609,N_16056,N_19199);
and UO_1610 (O_1610,N_16737,N_16439);
or UO_1611 (O_1611,N_17372,N_17339);
nor UO_1612 (O_1612,N_19852,N_18824);
xor UO_1613 (O_1613,N_16811,N_17602);
nor UO_1614 (O_1614,N_16697,N_18754);
or UO_1615 (O_1615,N_17505,N_18616);
xor UO_1616 (O_1616,N_16008,N_17196);
and UO_1617 (O_1617,N_17508,N_17844);
nand UO_1618 (O_1618,N_19245,N_18911);
nand UO_1619 (O_1619,N_18763,N_19532);
nor UO_1620 (O_1620,N_18737,N_16176);
xor UO_1621 (O_1621,N_19839,N_18399);
nand UO_1622 (O_1622,N_19545,N_18372);
and UO_1623 (O_1623,N_18614,N_19923);
or UO_1624 (O_1624,N_17413,N_17293);
nor UO_1625 (O_1625,N_19178,N_18673);
nand UO_1626 (O_1626,N_16281,N_16004);
xnor UO_1627 (O_1627,N_19599,N_17139);
xor UO_1628 (O_1628,N_19717,N_17416);
or UO_1629 (O_1629,N_18717,N_17193);
or UO_1630 (O_1630,N_18176,N_19603);
and UO_1631 (O_1631,N_17807,N_19986);
or UO_1632 (O_1632,N_18121,N_16003);
nor UO_1633 (O_1633,N_19742,N_19771);
xor UO_1634 (O_1634,N_16389,N_18686);
and UO_1635 (O_1635,N_17650,N_17517);
nor UO_1636 (O_1636,N_19757,N_18247);
nand UO_1637 (O_1637,N_16588,N_18194);
xnor UO_1638 (O_1638,N_19119,N_17152);
nand UO_1639 (O_1639,N_16437,N_17294);
and UO_1640 (O_1640,N_16883,N_19484);
nand UO_1641 (O_1641,N_16391,N_19752);
xnor UO_1642 (O_1642,N_18683,N_17459);
nand UO_1643 (O_1643,N_17940,N_17685);
nand UO_1644 (O_1644,N_19781,N_19897);
or UO_1645 (O_1645,N_16124,N_18747);
nor UO_1646 (O_1646,N_16117,N_17245);
xnor UO_1647 (O_1647,N_17552,N_17649);
and UO_1648 (O_1648,N_17721,N_19628);
or UO_1649 (O_1649,N_19941,N_18460);
nand UO_1650 (O_1650,N_19078,N_19098);
or UO_1651 (O_1651,N_19566,N_18173);
xnor UO_1652 (O_1652,N_18224,N_18155);
and UO_1653 (O_1653,N_16695,N_16304);
or UO_1654 (O_1654,N_18435,N_17730);
nor UO_1655 (O_1655,N_18225,N_19939);
xor UO_1656 (O_1656,N_17553,N_18702);
and UO_1657 (O_1657,N_19214,N_19632);
xor UO_1658 (O_1658,N_18762,N_17281);
nand UO_1659 (O_1659,N_17745,N_16315);
and UO_1660 (O_1660,N_17104,N_16460);
nand UO_1661 (O_1661,N_17270,N_19612);
or UO_1662 (O_1662,N_19696,N_16831);
xnor UO_1663 (O_1663,N_18580,N_16560);
nor UO_1664 (O_1664,N_19891,N_16546);
nor UO_1665 (O_1665,N_19844,N_18012);
and UO_1666 (O_1666,N_18462,N_17272);
nor UO_1667 (O_1667,N_19691,N_18359);
xnor UO_1668 (O_1668,N_16579,N_19335);
and UO_1669 (O_1669,N_19435,N_16475);
nand UO_1670 (O_1670,N_17966,N_17344);
xnor UO_1671 (O_1671,N_18115,N_19024);
and UO_1672 (O_1672,N_19651,N_17753);
nor UO_1673 (O_1673,N_17654,N_19455);
nor UO_1674 (O_1674,N_19017,N_18497);
xor UO_1675 (O_1675,N_16639,N_19066);
nand UO_1676 (O_1676,N_16169,N_16762);
and UO_1677 (O_1677,N_17812,N_18026);
nor UO_1678 (O_1678,N_17995,N_18360);
and UO_1679 (O_1679,N_19531,N_19899);
nand UO_1680 (O_1680,N_17780,N_18825);
nor UO_1681 (O_1681,N_19588,N_16661);
nor UO_1682 (O_1682,N_16705,N_17472);
nor UO_1683 (O_1683,N_16594,N_19988);
nor UO_1684 (O_1684,N_19870,N_19620);
nand UO_1685 (O_1685,N_16149,N_19931);
nand UO_1686 (O_1686,N_17887,N_19471);
nor UO_1687 (O_1687,N_18752,N_18216);
nand UO_1688 (O_1688,N_18732,N_16097);
nand UO_1689 (O_1689,N_18196,N_19808);
or UO_1690 (O_1690,N_18485,N_18509);
nor UO_1691 (O_1691,N_19995,N_16504);
and UO_1692 (O_1692,N_19444,N_19767);
nand UO_1693 (O_1693,N_16123,N_16356);
nor UO_1694 (O_1694,N_19843,N_19057);
or UO_1695 (O_1695,N_16141,N_17038);
nand UO_1696 (O_1696,N_19229,N_18934);
nand UO_1697 (O_1697,N_17584,N_18865);
nor UO_1698 (O_1698,N_18303,N_18682);
or UO_1699 (O_1699,N_16132,N_19714);
or UO_1700 (O_1700,N_18710,N_19332);
nor UO_1701 (O_1701,N_17715,N_19342);
nand UO_1702 (O_1702,N_16204,N_17611);
xor UO_1703 (O_1703,N_16679,N_19168);
nor UO_1704 (O_1704,N_19264,N_18861);
nand UO_1705 (O_1705,N_18637,N_18788);
or UO_1706 (O_1706,N_17479,N_19501);
nand UO_1707 (O_1707,N_18028,N_19949);
or UO_1708 (O_1708,N_18972,N_17744);
nand UO_1709 (O_1709,N_18553,N_19398);
nor UO_1710 (O_1710,N_18368,N_17255);
or UO_1711 (O_1711,N_18722,N_18907);
or UO_1712 (O_1712,N_16845,N_19103);
and UO_1713 (O_1713,N_16172,N_19524);
and UO_1714 (O_1714,N_16148,N_19558);
nand UO_1715 (O_1715,N_16428,N_17933);
nand UO_1716 (O_1716,N_19881,N_18103);
or UO_1717 (O_1717,N_17546,N_16246);
nor UO_1718 (O_1718,N_19148,N_16659);
and UO_1719 (O_1719,N_16284,N_16527);
and UO_1720 (O_1720,N_19555,N_19167);
nand UO_1721 (O_1721,N_19681,N_19141);
or UO_1722 (O_1722,N_16416,N_18630);
nor UO_1723 (O_1723,N_16662,N_18278);
nor UO_1724 (O_1724,N_19302,N_19597);
and UO_1725 (O_1725,N_18501,N_18109);
or UO_1726 (O_1726,N_18362,N_17155);
nand UO_1727 (O_1727,N_16237,N_16721);
or UO_1728 (O_1728,N_19866,N_19249);
and UO_1729 (O_1729,N_18957,N_16382);
and UO_1730 (O_1730,N_18659,N_16086);
nor UO_1731 (O_1731,N_17567,N_17267);
nor UO_1732 (O_1732,N_16776,N_16289);
and UO_1733 (O_1733,N_17314,N_17337);
nor UO_1734 (O_1734,N_17327,N_17792);
or UO_1735 (O_1735,N_18025,N_16433);
or UO_1736 (O_1736,N_17075,N_18408);
nand UO_1737 (O_1737,N_16842,N_18158);
nand UO_1738 (O_1738,N_18519,N_19347);
nor UO_1739 (O_1739,N_18960,N_18256);
xor UO_1740 (O_1740,N_18027,N_19019);
or UO_1741 (O_1741,N_17087,N_17079);
nand UO_1742 (O_1742,N_16597,N_19977);
nand UO_1743 (O_1743,N_19154,N_18412);
nor UO_1744 (O_1744,N_19610,N_17006);
and UO_1745 (O_1745,N_17099,N_16335);
and UO_1746 (O_1746,N_18077,N_18537);
and UO_1747 (O_1747,N_17253,N_17000);
or UO_1748 (O_1748,N_18899,N_16166);
nand UO_1749 (O_1749,N_19404,N_18014);
nand UO_1750 (O_1750,N_19020,N_17616);
and UO_1751 (O_1751,N_16053,N_17408);
nor UO_1752 (O_1752,N_19969,N_16380);
nor UO_1753 (O_1753,N_19345,N_19751);
nor UO_1754 (O_1754,N_18633,N_18566);
or UO_1755 (O_1755,N_19980,N_18472);
nor UO_1756 (O_1756,N_17922,N_17353);
and UO_1757 (O_1757,N_16915,N_16088);
nor UO_1758 (O_1758,N_18382,N_18487);
or UO_1759 (O_1759,N_18185,N_18915);
or UO_1760 (O_1760,N_16199,N_19952);
xor UO_1761 (O_1761,N_18913,N_17426);
and UO_1762 (O_1762,N_19436,N_18354);
xor UO_1763 (O_1763,N_19537,N_18626);
nor UO_1764 (O_1764,N_18113,N_19369);
nand UO_1765 (O_1765,N_16939,N_17279);
nand UO_1766 (O_1766,N_18442,N_18874);
and UO_1767 (O_1767,N_16485,N_19015);
nand UO_1768 (O_1768,N_16046,N_19830);
nor UO_1769 (O_1769,N_17221,N_19155);
nand UO_1770 (O_1770,N_19996,N_17729);
or UO_1771 (O_1771,N_17301,N_16536);
xnor UO_1772 (O_1772,N_16445,N_17120);
nand UO_1773 (O_1773,N_16248,N_19459);
nand UO_1774 (O_1774,N_16451,N_16421);
or UO_1775 (O_1775,N_17911,N_19505);
or UO_1776 (O_1776,N_17227,N_17544);
nand UO_1777 (O_1777,N_17394,N_18007);
or UO_1778 (O_1778,N_18445,N_18479);
nand UO_1779 (O_1779,N_16925,N_17879);
or UO_1780 (O_1780,N_18945,N_18230);
nand UO_1781 (O_1781,N_17536,N_17510);
or UO_1782 (O_1782,N_18331,N_18066);
and UO_1783 (O_1783,N_19235,N_17121);
and UO_1784 (O_1784,N_19466,N_17089);
or UO_1785 (O_1785,N_17138,N_19658);
xnor UO_1786 (O_1786,N_17370,N_18555);
nor UO_1787 (O_1787,N_16288,N_19397);
nand UO_1788 (O_1788,N_17059,N_17872);
or UO_1789 (O_1789,N_18383,N_18183);
and UO_1790 (O_1790,N_19613,N_19925);
nor UO_1791 (O_1791,N_17323,N_19391);
xnor UO_1792 (O_1792,N_16611,N_17226);
nand UO_1793 (O_1793,N_16778,N_18996);
or UO_1794 (O_1794,N_18356,N_17029);
nor UO_1795 (O_1795,N_19225,N_18903);
nor UO_1796 (O_1796,N_16942,N_16116);
and UO_1797 (O_1797,N_17697,N_16649);
xor UO_1798 (O_1798,N_18108,N_19203);
nand UO_1799 (O_1799,N_18106,N_16646);
nand UO_1800 (O_1800,N_19586,N_19937);
nor UO_1801 (O_1801,N_19557,N_19062);
or UO_1802 (O_1802,N_19095,N_19059);
or UO_1803 (O_1803,N_18753,N_16189);
nand UO_1804 (O_1804,N_18610,N_16947);
nor UO_1805 (O_1805,N_16602,N_17112);
nand UO_1806 (O_1806,N_16436,N_19886);
nor UO_1807 (O_1807,N_16030,N_19360);
nand UO_1808 (O_1808,N_19043,N_16665);
nand UO_1809 (O_1809,N_17900,N_19166);
xor UO_1810 (O_1810,N_17165,N_17558);
nor UO_1811 (O_1811,N_16224,N_19820);
nor UO_1812 (O_1812,N_16503,N_19805);
nor UO_1813 (O_1813,N_19590,N_16506);
nor UO_1814 (O_1814,N_19129,N_18766);
or UO_1815 (O_1815,N_19270,N_16002);
or UO_1816 (O_1816,N_18325,N_16983);
nand UO_1817 (O_1817,N_16345,N_18658);
nor UO_1818 (O_1818,N_16183,N_18172);
nand UO_1819 (O_1819,N_19585,N_16079);
and UO_1820 (O_1820,N_19876,N_16450);
nand UO_1821 (O_1821,N_17990,N_19170);
and UO_1822 (O_1822,N_19458,N_18831);
or UO_1823 (O_1823,N_16559,N_16231);
or UO_1824 (O_1824,N_19088,N_18151);
nand UO_1825 (O_1825,N_18868,N_19228);
nand UO_1826 (O_1826,N_18963,N_18901);
nand UO_1827 (O_1827,N_19259,N_19667);
and UO_1828 (O_1828,N_18315,N_16888);
xor UO_1829 (O_1829,N_19958,N_19615);
and UO_1830 (O_1830,N_18840,N_17194);
nand UO_1831 (O_1831,N_19423,N_19738);
or UO_1832 (O_1832,N_18712,N_17599);
nand UO_1833 (O_1833,N_19562,N_16044);
and UO_1834 (O_1834,N_18098,N_16311);
nor UO_1835 (O_1835,N_19343,N_18515);
nand UO_1836 (O_1836,N_19847,N_19135);
nand UO_1837 (O_1837,N_19561,N_19811);
xor UO_1838 (O_1838,N_17343,N_17362);
nor UO_1839 (O_1839,N_18248,N_16501);
xor UO_1840 (O_1840,N_17838,N_17642);
nor UO_1841 (O_1841,N_17041,N_19305);
nand UO_1842 (O_1842,N_16933,N_18417);
nor UO_1843 (O_1843,N_18297,N_18951);
nor UO_1844 (O_1844,N_16010,N_18500);
and UO_1845 (O_1845,N_19384,N_18353);
and UO_1846 (O_1846,N_17500,N_16834);
or UO_1847 (O_1847,N_19242,N_18896);
and UO_1848 (O_1848,N_16461,N_17373);
nor UO_1849 (O_1849,N_16324,N_19547);
and UO_1850 (O_1850,N_16233,N_19340);
or UO_1851 (O_1851,N_17969,N_16809);
xor UO_1852 (O_1852,N_17018,N_17359);
nor UO_1853 (O_1853,N_18346,N_19176);
xnor UO_1854 (O_1854,N_19579,N_19128);
nand UO_1855 (O_1855,N_18427,N_18927);
nand UO_1856 (O_1856,N_16054,N_18143);
and UO_1857 (O_1857,N_16178,N_19323);
nor UO_1858 (O_1858,N_18946,N_18550);
or UO_1859 (O_1859,N_17528,N_19251);
nand UO_1860 (O_1860,N_17891,N_18889);
nand UO_1861 (O_1861,N_19791,N_18999);
nor UO_1862 (O_1862,N_18667,N_18341);
nand UO_1863 (O_1863,N_16561,N_19703);
or UO_1864 (O_1864,N_16948,N_16660);
and UO_1865 (O_1865,N_18038,N_16209);
xnor UO_1866 (O_1866,N_18370,N_16768);
or UO_1867 (O_1867,N_16715,N_16493);
and UO_1868 (O_1868,N_16725,N_16941);
nor UO_1869 (O_1869,N_18119,N_16090);
or UO_1870 (O_1870,N_19131,N_18858);
nor UO_1871 (O_1871,N_16805,N_16656);
and UO_1872 (O_1872,N_17525,N_19477);
and UO_1873 (O_1873,N_19246,N_19644);
nor UO_1874 (O_1874,N_18819,N_18629);
xor UO_1875 (O_1875,N_16323,N_16017);
nor UO_1876 (O_1876,N_19550,N_19325);
or UO_1877 (O_1877,N_16489,N_18251);
nand UO_1878 (O_1878,N_19224,N_19328);
and UO_1879 (O_1879,N_19272,N_17325);
or UO_1880 (O_1880,N_16650,N_19352);
nand UO_1881 (O_1881,N_18716,N_17981);
xnor UO_1882 (O_1882,N_18890,N_19090);
or UO_1883 (O_1883,N_17077,N_18816);
nand UO_1884 (O_1884,N_16063,N_18878);
xnor UO_1885 (O_1885,N_17592,N_17219);
and UO_1886 (O_1886,N_19150,N_19609);
xnor UO_1887 (O_1887,N_19200,N_17102);
and UO_1888 (O_1888,N_18918,N_17011);
nand UO_1889 (O_1889,N_18920,N_17390);
and UO_1890 (O_1890,N_19065,N_19331);
nand UO_1891 (O_1891,N_19293,N_16988);
xnor UO_1892 (O_1892,N_18790,N_19730);
nor UO_1893 (O_1893,N_16853,N_19591);
nand UO_1894 (O_1894,N_19748,N_17824);
and UO_1895 (O_1895,N_19234,N_18493);
nor UO_1896 (O_1896,N_16028,N_19962);
nand UO_1897 (O_1897,N_16229,N_18063);
nand UO_1898 (O_1898,N_17638,N_18995);
nand UO_1899 (O_1899,N_17402,N_16029);
nand UO_1900 (O_1900,N_16127,N_16354);
or UO_1901 (O_1901,N_17049,N_16626);
nand UO_1902 (O_1902,N_16136,N_18525);
and UO_1903 (O_1903,N_18039,N_16387);
nand UO_1904 (O_1904,N_16384,N_17091);
nor UO_1905 (O_1905,N_17086,N_16547);
nand UO_1906 (O_1906,N_18311,N_17063);
and UO_1907 (O_1907,N_18636,N_18033);
xor UO_1908 (O_1908,N_18975,N_17683);
nand UO_1909 (O_1909,N_16824,N_17324);
or UO_1910 (O_1910,N_18948,N_16418);
nand UO_1911 (O_1911,N_18591,N_16589);
nor UO_1912 (O_1912,N_19675,N_16434);
nand UO_1913 (O_1913,N_18851,N_19341);
nor UO_1914 (O_1914,N_16688,N_18855);
or UO_1915 (O_1915,N_16790,N_17747);
or UO_1916 (O_1916,N_18546,N_18612);
and UO_1917 (O_1917,N_17082,N_19825);
and UO_1918 (O_1918,N_17421,N_17242);
nor UO_1919 (O_1919,N_19426,N_17797);
nand UO_1920 (O_1920,N_18740,N_17840);
and UO_1921 (O_1921,N_18492,N_19269);
nand UO_1922 (O_1922,N_18434,N_17460);
or UO_1923 (O_1923,N_18529,N_16641);
and UO_1924 (O_1924,N_18102,N_18441);
nor UO_1925 (O_1925,N_19447,N_16366);
and UO_1926 (O_1926,N_18455,N_17496);
and UO_1927 (O_1927,N_16773,N_17159);
nor UO_1928 (O_1928,N_16568,N_18955);
nand UO_1929 (O_1929,N_16061,N_18191);
or UO_1930 (O_1930,N_19401,N_16423);
or UO_1931 (O_1931,N_17060,N_17475);
and UO_1932 (O_1932,N_18724,N_18013);
nand UO_1933 (O_1933,N_19151,N_19773);
nand UO_1934 (O_1934,N_16585,N_19898);
and UO_1935 (O_1935,N_16302,N_17466);
or UO_1936 (O_1936,N_17799,N_19218);
and UO_1937 (O_1937,N_18388,N_18584);
and UO_1938 (O_1938,N_18751,N_17923);
nand UO_1939 (O_1939,N_16562,N_16483);
nand UO_1940 (O_1940,N_17725,N_18335);
and UO_1941 (O_1941,N_17434,N_18940);
xnor UO_1942 (O_1942,N_17050,N_16102);
xnor UO_1943 (O_1943,N_17814,N_16081);
nor UO_1944 (O_1944,N_17490,N_19935);
nor UO_1945 (O_1945,N_16701,N_16785);
nand UO_1946 (O_1946,N_16251,N_18542);
and UO_1947 (O_1947,N_16013,N_16073);
nand UO_1948 (O_1948,N_16388,N_18046);
and UO_1949 (O_1949,N_16468,N_17108);
nor UO_1950 (O_1950,N_18814,N_16686);
and UO_1951 (O_1951,N_17677,N_19522);
nor UO_1952 (O_1952,N_17149,N_17308);
nand UO_1953 (O_1953,N_16868,N_17643);
or UO_1954 (O_1954,N_16145,N_18405);
and UO_1955 (O_1955,N_16093,N_17384);
nor UO_1956 (O_1956,N_16754,N_19504);
and UO_1957 (O_1957,N_16091,N_19987);
nand UO_1958 (O_1958,N_18034,N_19337);
nor UO_1959 (O_1959,N_17710,N_19490);
and UO_1960 (O_1960,N_18801,N_16691);
nor UO_1961 (O_1961,N_17409,N_16802);
or UO_1962 (O_1962,N_16135,N_19330);
nor UO_1963 (O_1963,N_19743,N_18852);
nand UO_1964 (O_1964,N_19921,N_17212);
or UO_1965 (O_1965,N_19094,N_17924);
nor UO_1966 (O_1966,N_17871,N_19430);
nand UO_1967 (O_1967,N_18730,N_17101);
and UO_1968 (O_1968,N_18032,N_18126);
nand UO_1969 (O_1969,N_17974,N_19568);
and UO_1970 (O_1970,N_16678,N_16297);
nor UO_1971 (O_1971,N_16299,N_17246);
nand UO_1972 (O_1972,N_16360,N_17157);
or UO_1973 (O_1973,N_19448,N_16726);
or UO_1974 (O_1974,N_16314,N_16981);
and UO_1975 (O_1975,N_19244,N_16542);
or UO_1976 (O_1976,N_16143,N_18168);
nor UO_1977 (O_1977,N_16480,N_17128);
and UO_1978 (O_1978,N_18391,N_18971);
and UO_1979 (O_1979,N_18888,N_19520);
nand UO_1980 (O_1980,N_19564,N_19759);
and UO_1981 (O_1981,N_17899,N_16293);
nor UO_1982 (O_1982,N_19011,N_19104);
and UO_1983 (O_1983,N_16398,N_19833);
and UO_1984 (O_1984,N_19169,N_19854);
nor UO_1985 (O_1985,N_19638,N_16554);
nor UO_1986 (O_1986,N_16906,N_16935);
and UO_1987 (O_1987,N_17093,N_17722);
nand UO_1988 (O_1988,N_19646,N_16938);
and UO_1989 (O_1989,N_17215,N_19013);
nor UO_1990 (O_1990,N_16663,N_18728);
nor UO_1991 (O_1991,N_18085,N_19991);
nand UO_1992 (O_1992,N_19385,N_19928);
nand UO_1993 (O_1993,N_16069,N_17959);
and UO_1994 (O_1994,N_19028,N_19376);
nor UO_1995 (O_1995,N_18449,N_18062);
nor UO_1996 (O_1996,N_16722,N_18048);
nor UO_1997 (O_1997,N_16466,N_17675);
or UO_1998 (O_1998,N_19785,N_18904);
nand UO_1999 (O_1999,N_18502,N_16586);
and UO_2000 (O_2000,N_19314,N_16373);
and UO_2001 (O_2001,N_18397,N_18687);
and UO_2002 (O_2002,N_19968,N_18680);
or UO_2003 (O_2003,N_16587,N_19468);
xnor UO_2004 (O_2004,N_17959,N_19175);
or UO_2005 (O_2005,N_19318,N_19944);
nand UO_2006 (O_2006,N_19562,N_17248);
and UO_2007 (O_2007,N_17274,N_19008);
nand UO_2008 (O_2008,N_18652,N_18690);
and UO_2009 (O_2009,N_17498,N_19873);
xnor UO_2010 (O_2010,N_16381,N_19409);
nand UO_2011 (O_2011,N_19725,N_17907);
nand UO_2012 (O_2012,N_17913,N_17723);
and UO_2013 (O_2013,N_17572,N_17374);
and UO_2014 (O_2014,N_19700,N_18872);
xnor UO_2015 (O_2015,N_19390,N_18263);
xnor UO_2016 (O_2016,N_17291,N_18247);
nand UO_2017 (O_2017,N_16317,N_17673);
nor UO_2018 (O_2018,N_17187,N_18838);
nand UO_2019 (O_2019,N_16871,N_16141);
or UO_2020 (O_2020,N_19915,N_19938);
or UO_2021 (O_2021,N_16819,N_18155);
and UO_2022 (O_2022,N_19002,N_19601);
nand UO_2023 (O_2023,N_16333,N_18899);
nor UO_2024 (O_2024,N_17811,N_17000);
and UO_2025 (O_2025,N_19898,N_16519);
nor UO_2026 (O_2026,N_18564,N_17094);
xor UO_2027 (O_2027,N_17195,N_17537);
or UO_2028 (O_2028,N_19230,N_19641);
nor UO_2029 (O_2029,N_16184,N_16929);
nand UO_2030 (O_2030,N_17397,N_16966);
or UO_2031 (O_2031,N_17595,N_16244);
nand UO_2032 (O_2032,N_16569,N_18578);
nor UO_2033 (O_2033,N_16881,N_17505);
nand UO_2034 (O_2034,N_16829,N_17448);
nand UO_2035 (O_2035,N_19814,N_19944);
nor UO_2036 (O_2036,N_18229,N_16343);
and UO_2037 (O_2037,N_18880,N_18449);
nor UO_2038 (O_2038,N_16129,N_18661);
xnor UO_2039 (O_2039,N_18780,N_16054);
nor UO_2040 (O_2040,N_19564,N_16111);
or UO_2041 (O_2041,N_17514,N_16009);
and UO_2042 (O_2042,N_18480,N_17990);
nand UO_2043 (O_2043,N_16119,N_18399);
nor UO_2044 (O_2044,N_19415,N_19807);
or UO_2045 (O_2045,N_19702,N_17461);
xor UO_2046 (O_2046,N_18174,N_16457);
or UO_2047 (O_2047,N_16323,N_16264);
and UO_2048 (O_2048,N_16896,N_18915);
nand UO_2049 (O_2049,N_18436,N_16958);
and UO_2050 (O_2050,N_17250,N_16840);
or UO_2051 (O_2051,N_16427,N_19689);
or UO_2052 (O_2052,N_18010,N_19397);
or UO_2053 (O_2053,N_16357,N_17572);
and UO_2054 (O_2054,N_16584,N_17148);
nand UO_2055 (O_2055,N_19888,N_18820);
and UO_2056 (O_2056,N_16519,N_18980);
and UO_2057 (O_2057,N_19596,N_19216);
and UO_2058 (O_2058,N_17990,N_18711);
and UO_2059 (O_2059,N_19603,N_18493);
nor UO_2060 (O_2060,N_17489,N_19625);
and UO_2061 (O_2061,N_16534,N_19780);
nand UO_2062 (O_2062,N_17158,N_19355);
xor UO_2063 (O_2063,N_19831,N_18476);
or UO_2064 (O_2064,N_17472,N_18201);
or UO_2065 (O_2065,N_19560,N_17699);
or UO_2066 (O_2066,N_18691,N_17307);
or UO_2067 (O_2067,N_16190,N_19795);
or UO_2068 (O_2068,N_16986,N_18842);
nor UO_2069 (O_2069,N_16416,N_19473);
and UO_2070 (O_2070,N_17000,N_19628);
and UO_2071 (O_2071,N_17011,N_19561);
and UO_2072 (O_2072,N_17476,N_17393);
or UO_2073 (O_2073,N_19334,N_19168);
nand UO_2074 (O_2074,N_19267,N_17881);
and UO_2075 (O_2075,N_19945,N_19643);
and UO_2076 (O_2076,N_16211,N_18078);
xor UO_2077 (O_2077,N_17943,N_17412);
nand UO_2078 (O_2078,N_17222,N_17515);
nand UO_2079 (O_2079,N_16627,N_19660);
and UO_2080 (O_2080,N_16065,N_16212);
and UO_2081 (O_2081,N_16589,N_17319);
nor UO_2082 (O_2082,N_18787,N_19584);
nor UO_2083 (O_2083,N_19899,N_17008);
nor UO_2084 (O_2084,N_19254,N_18772);
and UO_2085 (O_2085,N_19868,N_19429);
and UO_2086 (O_2086,N_16067,N_19285);
nor UO_2087 (O_2087,N_17149,N_19264);
and UO_2088 (O_2088,N_19511,N_16033);
nand UO_2089 (O_2089,N_16910,N_16087);
or UO_2090 (O_2090,N_18854,N_19713);
nor UO_2091 (O_2091,N_18338,N_18753);
xnor UO_2092 (O_2092,N_18901,N_18802);
and UO_2093 (O_2093,N_16086,N_19550);
nor UO_2094 (O_2094,N_17137,N_17921);
and UO_2095 (O_2095,N_19758,N_19186);
and UO_2096 (O_2096,N_17390,N_19303);
nand UO_2097 (O_2097,N_18798,N_17979);
nor UO_2098 (O_2098,N_18908,N_18438);
and UO_2099 (O_2099,N_18920,N_16523);
xor UO_2100 (O_2100,N_17473,N_17619);
nor UO_2101 (O_2101,N_18584,N_18020);
nand UO_2102 (O_2102,N_16751,N_17019);
nand UO_2103 (O_2103,N_16836,N_16592);
xnor UO_2104 (O_2104,N_17660,N_17459);
nor UO_2105 (O_2105,N_19805,N_18152);
or UO_2106 (O_2106,N_16208,N_18390);
nand UO_2107 (O_2107,N_19257,N_18610);
and UO_2108 (O_2108,N_17290,N_16325);
nor UO_2109 (O_2109,N_16630,N_17583);
nor UO_2110 (O_2110,N_16428,N_17472);
nor UO_2111 (O_2111,N_19524,N_19142);
xnor UO_2112 (O_2112,N_19669,N_18527);
nand UO_2113 (O_2113,N_16705,N_18562);
or UO_2114 (O_2114,N_16381,N_18743);
nand UO_2115 (O_2115,N_16651,N_18718);
xor UO_2116 (O_2116,N_16440,N_19010);
nand UO_2117 (O_2117,N_16303,N_16285);
xnor UO_2118 (O_2118,N_17630,N_19460);
and UO_2119 (O_2119,N_16041,N_19993);
or UO_2120 (O_2120,N_19296,N_19029);
nand UO_2121 (O_2121,N_18974,N_18180);
nor UO_2122 (O_2122,N_16462,N_19268);
xor UO_2123 (O_2123,N_18122,N_17746);
nand UO_2124 (O_2124,N_18939,N_19546);
nand UO_2125 (O_2125,N_19572,N_17755);
nor UO_2126 (O_2126,N_18963,N_18703);
nor UO_2127 (O_2127,N_16960,N_18589);
nor UO_2128 (O_2128,N_17831,N_17550);
or UO_2129 (O_2129,N_19347,N_19025);
nand UO_2130 (O_2130,N_19886,N_18561);
or UO_2131 (O_2131,N_18657,N_17380);
and UO_2132 (O_2132,N_16326,N_17899);
or UO_2133 (O_2133,N_18401,N_19049);
or UO_2134 (O_2134,N_16431,N_18954);
nor UO_2135 (O_2135,N_17276,N_18248);
and UO_2136 (O_2136,N_19474,N_19655);
xor UO_2137 (O_2137,N_19146,N_18416);
nor UO_2138 (O_2138,N_19598,N_16063);
and UO_2139 (O_2139,N_16594,N_19269);
nand UO_2140 (O_2140,N_17810,N_16574);
and UO_2141 (O_2141,N_17616,N_16079);
and UO_2142 (O_2142,N_16550,N_19958);
or UO_2143 (O_2143,N_17432,N_17344);
nor UO_2144 (O_2144,N_19247,N_19949);
and UO_2145 (O_2145,N_17950,N_18542);
or UO_2146 (O_2146,N_17266,N_16641);
or UO_2147 (O_2147,N_16265,N_19923);
and UO_2148 (O_2148,N_19415,N_18124);
nor UO_2149 (O_2149,N_19573,N_18147);
and UO_2150 (O_2150,N_16131,N_18670);
nor UO_2151 (O_2151,N_16209,N_19321);
nor UO_2152 (O_2152,N_17882,N_19783);
and UO_2153 (O_2153,N_17614,N_19224);
nand UO_2154 (O_2154,N_16613,N_16915);
and UO_2155 (O_2155,N_18718,N_19497);
nor UO_2156 (O_2156,N_18901,N_17407);
and UO_2157 (O_2157,N_18649,N_17055);
and UO_2158 (O_2158,N_17187,N_16590);
or UO_2159 (O_2159,N_16694,N_17068);
or UO_2160 (O_2160,N_19866,N_17945);
nor UO_2161 (O_2161,N_18639,N_18086);
nand UO_2162 (O_2162,N_16674,N_16310);
and UO_2163 (O_2163,N_18027,N_17819);
or UO_2164 (O_2164,N_16895,N_18572);
nor UO_2165 (O_2165,N_18640,N_17101);
nand UO_2166 (O_2166,N_16737,N_19544);
nand UO_2167 (O_2167,N_19684,N_17345);
nand UO_2168 (O_2168,N_18617,N_16799);
nand UO_2169 (O_2169,N_16751,N_16102);
nor UO_2170 (O_2170,N_16839,N_16861);
nand UO_2171 (O_2171,N_17272,N_17539);
or UO_2172 (O_2172,N_18407,N_19869);
nor UO_2173 (O_2173,N_19604,N_16049);
and UO_2174 (O_2174,N_16317,N_17459);
nand UO_2175 (O_2175,N_19774,N_18393);
xnor UO_2176 (O_2176,N_19151,N_19008);
or UO_2177 (O_2177,N_16633,N_19030);
nand UO_2178 (O_2178,N_17889,N_18257);
or UO_2179 (O_2179,N_17459,N_16383);
and UO_2180 (O_2180,N_19068,N_19648);
nor UO_2181 (O_2181,N_18248,N_18901);
nor UO_2182 (O_2182,N_18811,N_17896);
or UO_2183 (O_2183,N_19608,N_19354);
nor UO_2184 (O_2184,N_18596,N_16722);
xnor UO_2185 (O_2185,N_17950,N_18355);
or UO_2186 (O_2186,N_19473,N_19695);
and UO_2187 (O_2187,N_18553,N_16936);
and UO_2188 (O_2188,N_18990,N_17155);
and UO_2189 (O_2189,N_17129,N_19082);
nand UO_2190 (O_2190,N_19975,N_16886);
nand UO_2191 (O_2191,N_18658,N_18695);
and UO_2192 (O_2192,N_19625,N_19000);
nand UO_2193 (O_2193,N_16253,N_17057);
nor UO_2194 (O_2194,N_17830,N_16901);
xor UO_2195 (O_2195,N_19791,N_19871);
nor UO_2196 (O_2196,N_16026,N_16496);
and UO_2197 (O_2197,N_17333,N_17302);
or UO_2198 (O_2198,N_18031,N_16504);
or UO_2199 (O_2199,N_16887,N_16930);
and UO_2200 (O_2200,N_16993,N_19710);
nor UO_2201 (O_2201,N_18020,N_16659);
nand UO_2202 (O_2202,N_16473,N_17849);
nor UO_2203 (O_2203,N_17356,N_16468);
or UO_2204 (O_2204,N_16828,N_18030);
or UO_2205 (O_2205,N_16133,N_17875);
or UO_2206 (O_2206,N_19711,N_19695);
or UO_2207 (O_2207,N_18364,N_19789);
and UO_2208 (O_2208,N_18151,N_17754);
nor UO_2209 (O_2209,N_18713,N_17310);
or UO_2210 (O_2210,N_16056,N_17937);
xnor UO_2211 (O_2211,N_17384,N_17093);
or UO_2212 (O_2212,N_19454,N_18448);
nand UO_2213 (O_2213,N_16212,N_19026);
nor UO_2214 (O_2214,N_18943,N_17360);
xnor UO_2215 (O_2215,N_16075,N_19315);
nand UO_2216 (O_2216,N_18701,N_16435);
nor UO_2217 (O_2217,N_19380,N_18631);
or UO_2218 (O_2218,N_19626,N_16061);
nor UO_2219 (O_2219,N_19178,N_19775);
and UO_2220 (O_2220,N_18649,N_17083);
or UO_2221 (O_2221,N_18619,N_18631);
and UO_2222 (O_2222,N_17681,N_16326);
and UO_2223 (O_2223,N_16252,N_18424);
nand UO_2224 (O_2224,N_19431,N_17286);
or UO_2225 (O_2225,N_18521,N_16235);
xnor UO_2226 (O_2226,N_17483,N_17296);
nand UO_2227 (O_2227,N_18084,N_17032);
or UO_2228 (O_2228,N_18061,N_17714);
and UO_2229 (O_2229,N_17227,N_17443);
nand UO_2230 (O_2230,N_16888,N_18029);
or UO_2231 (O_2231,N_17621,N_17469);
nand UO_2232 (O_2232,N_16093,N_16696);
or UO_2233 (O_2233,N_18097,N_17773);
and UO_2234 (O_2234,N_18559,N_17282);
nor UO_2235 (O_2235,N_19212,N_16347);
or UO_2236 (O_2236,N_16324,N_19952);
nor UO_2237 (O_2237,N_16882,N_19113);
nand UO_2238 (O_2238,N_17727,N_19322);
or UO_2239 (O_2239,N_18523,N_18468);
nor UO_2240 (O_2240,N_17641,N_19716);
nor UO_2241 (O_2241,N_16022,N_16825);
xnor UO_2242 (O_2242,N_18341,N_17952);
nand UO_2243 (O_2243,N_18295,N_17704);
or UO_2244 (O_2244,N_16648,N_18451);
or UO_2245 (O_2245,N_19098,N_18480);
xor UO_2246 (O_2246,N_19928,N_19253);
or UO_2247 (O_2247,N_17509,N_19720);
or UO_2248 (O_2248,N_18807,N_17291);
nor UO_2249 (O_2249,N_19368,N_17659);
nor UO_2250 (O_2250,N_17757,N_16868);
xnor UO_2251 (O_2251,N_16452,N_18367);
and UO_2252 (O_2252,N_16124,N_19890);
xnor UO_2253 (O_2253,N_19846,N_18754);
and UO_2254 (O_2254,N_19928,N_18441);
and UO_2255 (O_2255,N_18804,N_16652);
or UO_2256 (O_2256,N_16562,N_16853);
and UO_2257 (O_2257,N_18281,N_17357);
nand UO_2258 (O_2258,N_17064,N_16653);
and UO_2259 (O_2259,N_17350,N_19602);
or UO_2260 (O_2260,N_17985,N_19770);
nor UO_2261 (O_2261,N_16891,N_17653);
nor UO_2262 (O_2262,N_19273,N_16222);
and UO_2263 (O_2263,N_19134,N_18655);
or UO_2264 (O_2264,N_18001,N_16379);
nor UO_2265 (O_2265,N_17424,N_18607);
nand UO_2266 (O_2266,N_18252,N_19261);
nor UO_2267 (O_2267,N_18589,N_19718);
and UO_2268 (O_2268,N_17905,N_17396);
nor UO_2269 (O_2269,N_17572,N_19499);
and UO_2270 (O_2270,N_19761,N_16544);
xnor UO_2271 (O_2271,N_18087,N_16782);
xnor UO_2272 (O_2272,N_17526,N_17397);
and UO_2273 (O_2273,N_18740,N_19635);
and UO_2274 (O_2274,N_17920,N_16888);
nand UO_2275 (O_2275,N_17626,N_17531);
xor UO_2276 (O_2276,N_16493,N_19365);
nand UO_2277 (O_2277,N_17999,N_18596);
and UO_2278 (O_2278,N_19262,N_18068);
nand UO_2279 (O_2279,N_16532,N_17394);
nand UO_2280 (O_2280,N_16391,N_17232);
nor UO_2281 (O_2281,N_19759,N_16466);
or UO_2282 (O_2282,N_19477,N_17321);
xnor UO_2283 (O_2283,N_19440,N_17853);
nor UO_2284 (O_2284,N_16404,N_16481);
nor UO_2285 (O_2285,N_19544,N_16395);
or UO_2286 (O_2286,N_17493,N_17616);
or UO_2287 (O_2287,N_19498,N_19560);
nor UO_2288 (O_2288,N_19043,N_17454);
nand UO_2289 (O_2289,N_16474,N_17899);
nor UO_2290 (O_2290,N_17493,N_16482);
and UO_2291 (O_2291,N_17613,N_16587);
nand UO_2292 (O_2292,N_16963,N_18454);
nor UO_2293 (O_2293,N_16387,N_18566);
nand UO_2294 (O_2294,N_18026,N_16881);
xnor UO_2295 (O_2295,N_17781,N_19045);
nor UO_2296 (O_2296,N_16127,N_18510);
or UO_2297 (O_2297,N_18817,N_19723);
and UO_2298 (O_2298,N_17664,N_18772);
nand UO_2299 (O_2299,N_18732,N_16123);
xnor UO_2300 (O_2300,N_17723,N_16062);
nor UO_2301 (O_2301,N_19781,N_16137);
and UO_2302 (O_2302,N_16154,N_16270);
nand UO_2303 (O_2303,N_17599,N_16016);
nand UO_2304 (O_2304,N_17748,N_17190);
nand UO_2305 (O_2305,N_16575,N_19191);
nor UO_2306 (O_2306,N_18762,N_18934);
and UO_2307 (O_2307,N_18111,N_16166);
xor UO_2308 (O_2308,N_17505,N_19367);
or UO_2309 (O_2309,N_18353,N_16794);
nand UO_2310 (O_2310,N_18629,N_19542);
nand UO_2311 (O_2311,N_17244,N_19716);
xnor UO_2312 (O_2312,N_17237,N_19014);
and UO_2313 (O_2313,N_19258,N_19221);
nand UO_2314 (O_2314,N_19402,N_19455);
nand UO_2315 (O_2315,N_19331,N_18561);
nand UO_2316 (O_2316,N_16683,N_16002);
nor UO_2317 (O_2317,N_19135,N_16160);
and UO_2318 (O_2318,N_16668,N_18812);
nand UO_2319 (O_2319,N_17341,N_18021);
nand UO_2320 (O_2320,N_17894,N_18562);
nor UO_2321 (O_2321,N_18931,N_16397);
xnor UO_2322 (O_2322,N_17332,N_19991);
or UO_2323 (O_2323,N_19958,N_17528);
nor UO_2324 (O_2324,N_18395,N_18310);
or UO_2325 (O_2325,N_16855,N_17131);
nor UO_2326 (O_2326,N_18669,N_18632);
and UO_2327 (O_2327,N_18508,N_17955);
nand UO_2328 (O_2328,N_17863,N_17811);
or UO_2329 (O_2329,N_17545,N_19968);
or UO_2330 (O_2330,N_18851,N_17040);
or UO_2331 (O_2331,N_17650,N_16637);
nand UO_2332 (O_2332,N_19490,N_19074);
nor UO_2333 (O_2333,N_16393,N_18065);
nor UO_2334 (O_2334,N_17515,N_16220);
xnor UO_2335 (O_2335,N_17653,N_19903);
nand UO_2336 (O_2336,N_16485,N_16072);
or UO_2337 (O_2337,N_17923,N_16091);
nand UO_2338 (O_2338,N_18831,N_16907);
nor UO_2339 (O_2339,N_16474,N_18597);
nand UO_2340 (O_2340,N_19576,N_16435);
or UO_2341 (O_2341,N_16696,N_16905);
nor UO_2342 (O_2342,N_16128,N_18096);
nor UO_2343 (O_2343,N_19624,N_16359);
nand UO_2344 (O_2344,N_17835,N_17660);
nor UO_2345 (O_2345,N_17995,N_16143);
nand UO_2346 (O_2346,N_18309,N_19109);
xor UO_2347 (O_2347,N_17208,N_19584);
nand UO_2348 (O_2348,N_18240,N_19850);
xor UO_2349 (O_2349,N_19690,N_19348);
and UO_2350 (O_2350,N_19253,N_16831);
nand UO_2351 (O_2351,N_18667,N_18000);
or UO_2352 (O_2352,N_19539,N_16473);
and UO_2353 (O_2353,N_16358,N_18342);
and UO_2354 (O_2354,N_18136,N_19739);
and UO_2355 (O_2355,N_19122,N_16356);
or UO_2356 (O_2356,N_18961,N_18853);
nand UO_2357 (O_2357,N_16617,N_19916);
nand UO_2358 (O_2358,N_18443,N_16688);
or UO_2359 (O_2359,N_16633,N_16447);
nand UO_2360 (O_2360,N_16229,N_19744);
or UO_2361 (O_2361,N_18308,N_18560);
xor UO_2362 (O_2362,N_19940,N_17005);
nand UO_2363 (O_2363,N_16589,N_18070);
and UO_2364 (O_2364,N_16599,N_17527);
or UO_2365 (O_2365,N_17278,N_17924);
xor UO_2366 (O_2366,N_16648,N_16815);
nor UO_2367 (O_2367,N_19158,N_19846);
nand UO_2368 (O_2368,N_17773,N_18863);
or UO_2369 (O_2369,N_19631,N_19879);
xor UO_2370 (O_2370,N_16883,N_17078);
nor UO_2371 (O_2371,N_18056,N_16414);
xnor UO_2372 (O_2372,N_16687,N_16435);
or UO_2373 (O_2373,N_16811,N_19513);
or UO_2374 (O_2374,N_17036,N_18354);
and UO_2375 (O_2375,N_18446,N_19406);
xnor UO_2376 (O_2376,N_18254,N_19343);
nand UO_2377 (O_2377,N_18745,N_17617);
nand UO_2378 (O_2378,N_19439,N_16175);
nand UO_2379 (O_2379,N_17366,N_17178);
nor UO_2380 (O_2380,N_18155,N_18804);
nor UO_2381 (O_2381,N_17701,N_19621);
nand UO_2382 (O_2382,N_16536,N_18516);
nand UO_2383 (O_2383,N_19790,N_17389);
and UO_2384 (O_2384,N_19542,N_17864);
or UO_2385 (O_2385,N_16513,N_18643);
nand UO_2386 (O_2386,N_17171,N_18252);
nor UO_2387 (O_2387,N_18338,N_18922);
nor UO_2388 (O_2388,N_18537,N_17463);
xnor UO_2389 (O_2389,N_16390,N_19499);
nand UO_2390 (O_2390,N_17287,N_19570);
and UO_2391 (O_2391,N_19074,N_19268);
nor UO_2392 (O_2392,N_16767,N_16970);
nand UO_2393 (O_2393,N_19129,N_18678);
nand UO_2394 (O_2394,N_16384,N_19871);
and UO_2395 (O_2395,N_19395,N_18836);
nand UO_2396 (O_2396,N_19184,N_16363);
or UO_2397 (O_2397,N_18934,N_16295);
nand UO_2398 (O_2398,N_18652,N_17670);
nand UO_2399 (O_2399,N_18598,N_19096);
nor UO_2400 (O_2400,N_19534,N_16386);
nand UO_2401 (O_2401,N_17572,N_18025);
nor UO_2402 (O_2402,N_17342,N_17132);
xnor UO_2403 (O_2403,N_17184,N_19028);
nor UO_2404 (O_2404,N_18898,N_16128);
nor UO_2405 (O_2405,N_16155,N_17680);
nand UO_2406 (O_2406,N_17180,N_16964);
nor UO_2407 (O_2407,N_19545,N_19807);
or UO_2408 (O_2408,N_16929,N_17543);
or UO_2409 (O_2409,N_16146,N_18357);
nand UO_2410 (O_2410,N_18391,N_16775);
nand UO_2411 (O_2411,N_17203,N_16927);
and UO_2412 (O_2412,N_18801,N_19367);
nand UO_2413 (O_2413,N_18763,N_19039);
or UO_2414 (O_2414,N_19577,N_17042);
nand UO_2415 (O_2415,N_18120,N_19741);
or UO_2416 (O_2416,N_19011,N_16025);
nor UO_2417 (O_2417,N_19307,N_19389);
nand UO_2418 (O_2418,N_17613,N_17445);
nor UO_2419 (O_2419,N_19109,N_16285);
nor UO_2420 (O_2420,N_16737,N_16465);
and UO_2421 (O_2421,N_16260,N_18475);
or UO_2422 (O_2422,N_16393,N_16670);
or UO_2423 (O_2423,N_17780,N_18506);
nor UO_2424 (O_2424,N_18155,N_18468);
or UO_2425 (O_2425,N_19742,N_18861);
or UO_2426 (O_2426,N_19035,N_19782);
nand UO_2427 (O_2427,N_16177,N_18062);
or UO_2428 (O_2428,N_18414,N_17381);
nor UO_2429 (O_2429,N_18159,N_16462);
nand UO_2430 (O_2430,N_16722,N_18060);
nand UO_2431 (O_2431,N_19993,N_19666);
and UO_2432 (O_2432,N_19911,N_17810);
nor UO_2433 (O_2433,N_19845,N_18702);
xnor UO_2434 (O_2434,N_18028,N_16641);
or UO_2435 (O_2435,N_16941,N_19286);
nor UO_2436 (O_2436,N_17971,N_19397);
nor UO_2437 (O_2437,N_16768,N_19296);
nor UO_2438 (O_2438,N_19399,N_18194);
and UO_2439 (O_2439,N_19995,N_17592);
and UO_2440 (O_2440,N_18996,N_18039);
nand UO_2441 (O_2441,N_17081,N_19777);
xor UO_2442 (O_2442,N_16754,N_17540);
and UO_2443 (O_2443,N_18926,N_19247);
or UO_2444 (O_2444,N_18017,N_19207);
or UO_2445 (O_2445,N_16483,N_18710);
nor UO_2446 (O_2446,N_16703,N_16442);
nand UO_2447 (O_2447,N_17882,N_19865);
or UO_2448 (O_2448,N_18298,N_19151);
and UO_2449 (O_2449,N_18665,N_18305);
nor UO_2450 (O_2450,N_17596,N_19165);
or UO_2451 (O_2451,N_17434,N_17128);
nor UO_2452 (O_2452,N_18135,N_17537);
or UO_2453 (O_2453,N_19037,N_16352);
or UO_2454 (O_2454,N_16368,N_19214);
or UO_2455 (O_2455,N_18403,N_17600);
nor UO_2456 (O_2456,N_17323,N_19365);
or UO_2457 (O_2457,N_19132,N_16517);
or UO_2458 (O_2458,N_17708,N_17479);
or UO_2459 (O_2459,N_19505,N_19899);
and UO_2460 (O_2460,N_19313,N_18316);
and UO_2461 (O_2461,N_18458,N_19386);
or UO_2462 (O_2462,N_17613,N_18743);
and UO_2463 (O_2463,N_19318,N_17535);
or UO_2464 (O_2464,N_19245,N_17477);
xor UO_2465 (O_2465,N_19056,N_17149);
or UO_2466 (O_2466,N_17089,N_16243);
nor UO_2467 (O_2467,N_17352,N_19102);
nor UO_2468 (O_2468,N_18166,N_19004);
nand UO_2469 (O_2469,N_17534,N_17317);
or UO_2470 (O_2470,N_17650,N_17755);
nand UO_2471 (O_2471,N_16424,N_16000);
and UO_2472 (O_2472,N_17150,N_17853);
or UO_2473 (O_2473,N_16302,N_17152);
or UO_2474 (O_2474,N_17232,N_16879);
nand UO_2475 (O_2475,N_18562,N_16439);
or UO_2476 (O_2476,N_18295,N_16247);
xnor UO_2477 (O_2477,N_17229,N_19155);
and UO_2478 (O_2478,N_18228,N_19371);
nor UO_2479 (O_2479,N_16187,N_16239);
nand UO_2480 (O_2480,N_17150,N_18888);
xor UO_2481 (O_2481,N_18084,N_18327);
xor UO_2482 (O_2482,N_18776,N_18927);
nor UO_2483 (O_2483,N_19222,N_18569);
or UO_2484 (O_2484,N_17588,N_18540);
nor UO_2485 (O_2485,N_18379,N_16716);
and UO_2486 (O_2486,N_18167,N_19675);
nor UO_2487 (O_2487,N_18471,N_17205);
xnor UO_2488 (O_2488,N_17492,N_19207);
nor UO_2489 (O_2489,N_19696,N_16449);
and UO_2490 (O_2490,N_17864,N_17785);
nand UO_2491 (O_2491,N_16231,N_16259);
nor UO_2492 (O_2492,N_17828,N_19891);
or UO_2493 (O_2493,N_16243,N_16414);
or UO_2494 (O_2494,N_19043,N_17894);
or UO_2495 (O_2495,N_18716,N_19260);
nand UO_2496 (O_2496,N_18442,N_19689);
and UO_2497 (O_2497,N_16904,N_16266);
or UO_2498 (O_2498,N_19752,N_19657);
nand UO_2499 (O_2499,N_19438,N_17262);
endmodule