module basic_2000_20000_2500_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1840,In_1105);
and U1 (N_1,In_1398,In_279);
nand U2 (N_2,In_1873,In_108);
nand U3 (N_3,In_605,In_857);
nor U4 (N_4,In_1715,In_1075);
or U5 (N_5,In_706,In_596);
nand U6 (N_6,In_906,In_157);
xnor U7 (N_7,In_1851,In_213);
or U8 (N_8,In_328,In_1215);
nor U9 (N_9,In_936,In_426);
nand U10 (N_10,In_1405,In_69);
or U11 (N_11,In_1511,In_1368);
xor U12 (N_12,In_1196,In_1136);
and U13 (N_13,In_1123,In_1596);
nor U14 (N_14,In_1619,In_9);
and U15 (N_15,In_1327,In_1239);
nand U16 (N_16,In_1080,In_948);
or U17 (N_17,In_761,In_1953);
nand U18 (N_18,In_1412,In_1231);
and U19 (N_19,In_1346,In_577);
or U20 (N_20,In_1127,In_172);
nor U21 (N_21,In_560,In_124);
or U22 (N_22,In_477,In_1950);
nand U23 (N_23,In_767,In_280);
nand U24 (N_24,In_1340,In_23);
or U25 (N_25,In_1587,In_1021);
xor U26 (N_26,In_1498,In_620);
nand U27 (N_27,In_1278,In_915);
or U28 (N_28,In_1572,In_1833);
nand U29 (N_29,In_1914,In_87);
nand U30 (N_30,In_917,In_104);
nor U31 (N_31,In_229,In_292);
xnor U32 (N_32,In_1975,In_1118);
nor U33 (N_33,In_1857,In_1148);
and U34 (N_34,In_960,In_750);
xor U35 (N_35,In_1053,In_1030);
nor U36 (N_36,In_600,In_497);
or U37 (N_37,In_595,In_447);
xor U38 (N_38,In_552,In_1515);
nand U39 (N_39,In_1439,In_914);
nor U40 (N_40,In_296,In_766);
nor U41 (N_41,In_13,In_51);
xor U42 (N_42,In_524,In_663);
or U43 (N_43,In_291,In_347);
xnor U44 (N_44,In_1742,In_772);
xor U45 (N_45,In_176,In_238);
xnor U46 (N_46,In_1437,In_697);
and U47 (N_47,In_308,In_476);
and U48 (N_48,In_1130,In_617);
xnor U49 (N_49,In_145,In_516);
nand U50 (N_50,In_1977,In_470);
nor U51 (N_51,In_488,In_660);
and U52 (N_52,In_437,In_1777);
xor U53 (N_53,In_775,In_231);
or U54 (N_54,In_1804,In_1828);
nor U55 (N_55,In_1948,In_1556);
nor U56 (N_56,In_537,In_1124);
nor U57 (N_57,In_1653,In_1473);
xnor U58 (N_58,In_679,In_1012);
or U59 (N_59,In_1680,In_1481);
and U60 (N_60,In_1815,In_34);
nor U61 (N_61,In_1630,In_1474);
and U62 (N_62,In_127,In_216);
or U63 (N_63,In_668,In_55);
nand U64 (N_64,In_763,In_546);
nor U65 (N_65,In_746,In_743);
nand U66 (N_66,In_727,In_1378);
nor U67 (N_67,In_1035,In_922);
or U68 (N_68,In_634,In_1272);
nor U69 (N_69,In_1218,In_1013);
nand U70 (N_70,In_1959,In_155);
and U71 (N_71,In_30,In_959);
nor U72 (N_72,In_1343,In_1791);
nand U73 (N_73,In_1536,In_1158);
nor U74 (N_74,In_1685,In_318);
and U75 (N_75,In_1911,In_616);
xor U76 (N_76,In_764,In_1312);
nand U77 (N_77,In_554,In_1357);
or U78 (N_78,In_1877,In_412);
nand U79 (N_79,In_1837,In_645);
nand U80 (N_80,In_359,In_869);
xor U81 (N_81,In_952,In_1902);
nor U82 (N_82,In_1812,In_1388);
nor U83 (N_83,In_496,In_838);
or U84 (N_84,In_1037,In_1734);
and U85 (N_85,In_1025,In_378);
xor U86 (N_86,In_1475,In_1095);
xnor U87 (N_87,In_726,In_452);
and U88 (N_88,In_1187,In_1735);
nor U89 (N_89,In_950,In_1930);
nor U90 (N_90,In_626,In_1903);
xnor U91 (N_91,In_1768,In_1623);
or U92 (N_92,In_1248,In_137);
or U93 (N_93,In_1585,In_29);
nand U94 (N_94,In_1334,In_326);
nor U95 (N_95,In_1070,In_1298);
and U96 (N_96,In_286,In_1329);
nand U97 (N_97,In_1604,In_1979);
xor U98 (N_98,In_938,In_47);
or U99 (N_99,In_1933,In_994);
and U100 (N_100,In_1874,In_1721);
xnor U101 (N_101,In_1602,In_1171);
and U102 (N_102,In_1484,In_141);
nor U103 (N_103,In_411,In_539);
or U104 (N_104,In_1699,In_93);
and U105 (N_105,In_1214,In_1417);
or U106 (N_106,In_1045,In_1076);
nor U107 (N_107,In_268,In_1956);
and U108 (N_108,In_1390,In_1251);
xor U109 (N_109,In_1372,In_1918);
and U110 (N_110,In_1011,In_1269);
xnor U111 (N_111,In_1254,In_1594);
or U112 (N_112,In_1686,In_1925);
nand U113 (N_113,In_841,In_888);
or U114 (N_114,In_895,In_196);
or U115 (N_115,In_712,In_345);
nor U116 (N_116,In_757,In_1164);
nor U117 (N_117,In_1018,In_250);
and U118 (N_118,In_852,In_1490);
xnor U119 (N_119,In_1938,In_981);
nor U120 (N_120,In_1794,In_442);
xor U121 (N_121,In_774,In_1769);
nand U122 (N_122,In_1816,In_1692);
nor U123 (N_123,In_1316,In_165);
nand U124 (N_124,In_581,In_957);
or U125 (N_125,In_1611,In_1170);
or U126 (N_126,In_1762,In_622);
xor U127 (N_127,In_1448,In_1726);
xor U128 (N_128,In_1173,In_1360);
xnor U129 (N_129,In_1972,In_86);
nand U130 (N_130,In_717,In_1431);
nand U131 (N_131,In_1188,In_843);
xnor U132 (N_132,In_222,In_803);
and U133 (N_133,In_203,In_457);
and U134 (N_134,In_1322,In_110);
or U135 (N_135,In_1121,In_502);
nor U136 (N_136,In_850,In_1951);
xnor U137 (N_137,In_10,In_1072);
or U138 (N_138,In_694,In_787);
or U139 (N_139,In_673,In_313);
xnor U140 (N_140,In_773,In_1210);
xor U141 (N_141,In_1748,In_1798);
nor U142 (N_142,In_1666,In_354);
nand U143 (N_143,In_1182,In_640);
xnor U144 (N_144,In_220,In_1954);
xor U145 (N_145,In_830,In_603);
nor U146 (N_146,In_1440,In_372);
nor U147 (N_147,In_1042,In_1132);
or U148 (N_148,In_1553,In_342);
nor U149 (N_149,In_1016,In_1510);
nor U150 (N_150,In_814,In_1443);
nor U151 (N_151,In_1714,In_1701);
xor U152 (N_152,In_1051,In_1201);
or U153 (N_153,In_885,In_333);
nor U154 (N_154,In_43,In_1356);
xnor U155 (N_155,In_1819,In_659);
nand U156 (N_156,In_919,In_1420);
nand U157 (N_157,In_60,In_541);
nor U158 (N_158,In_1458,In_1811);
xor U159 (N_159,In_1563,In_1947);
nor U160 (N_160,In_262,In_1307);
and U161 (N_161,In_863,In_64);
xnor U162 (N_162,In_718,In_271);
xor U163 (N_163,In_45,In_37);
nor U164 (N_164,In_584,In_930);
xor U165 (N_165,In_1221,In_1174);
nand U166 (N_166,In_283,In_968);
xor U167 (N_167,In_287,In_1236);
nor U168 (N_168,In_1415,In_954);
and U169 (N_169,In_369,In_877);
nand U170 (N_170,In_479,In_884);
nor U171 (N_171,In_218,In_1999);
nand U172 (N_172,In_1424,In_1371);
nor U173 (N_173,In_1129,In_1891);
nand U174 (N_174,In_682,In_484);
nand U175 (N_175,In_591,In_1617);
nor U176 (N_176,In_1382,In_490);
nand U177 (N_177,In_1491,In_251);
nand U178 (N_178,In_1416,In_1883);
xor U179 (N_179,In_1281,In_1758);
xnor U180 (N_180,In_740,In_818);
nor U181 (N_181,In_1419,In_851);
or U182 (N_182,In_953,In_1019);
nor U183 (N_183,In_1880,In_6);
or U184 (N_184,In_1519,In_1684);
nand U185 (N_185,In_168,In_1659);
and U186 (N_186,In_1471,In_1761);
xnor U187 (N_187,In_1559,In_97);
nor U188 (N_188,In_1286,In_1526);
nand U189 (N_189,In_1125,In_1493);
nor U190 (N_190,In_192,In_445);
nand U191 (N_191,In_1856,In_329);
or U192 (N_192,In_17,In_1425);
nand U193 (N_193,In_901,In_1632);
and U194 (N_194,In_1647,In_1151);
nor U195 (N_195,In_257,In_471);
and U196 (N_196,In_1970,In_711);
or U197 (N_197,In_702,In_1482);
nor U198 (N_198,In_1,In_710);
and U199 (N_199,In_1079,In_1780);
and U200 (N_200,In_31,In_1292);
nand U201 (N_201,In_1932,In_1328);
xnor U202 (N_202,In_294,In_80);
and U203 (N_203,In_654,In_1900);
and U204 (N_204,In_1504,In_21);
and U205 (N_205,In_1062,In_847);
or U206 (N_206,In_902,In_1213);
and U207 (N_207,In_1314,In_1789);
and U208 (N_208,In_1983,In_241);
nand U209 (N_209,In_74,In_138);
nor U210 (N_210,In_782,In_462);
and U211 (N_211,In_1919,In_1108);
nand U212 (N_212,In_1285,In_1376);
and U213 (N_213,In_252,In_1598);
or U214 (N_214,In_1595,In_995);
and U215 (N_215,In_453,In_664);
and U216 (N_216,In_908,In_201);
nor U217 (N_217,In_234,In_1884);
or U218 (N_218,In_842,In_236);
xnor U219 (N_219,In_1797,In_1060);
xor U220 (N_220,In_864,In_182);
or U221 (N_221,In_628,In_1090);
and U222 (N_222,In_449,In_1696);
xnor U223 (N_223,In_1428,In_481);
or U224 (N_224,In_1176,In_428);
nand U225 (N_225,In_184,In_824);
nor U226 (N_226,In_1896,In_1909);
or U227 (N_227,In_1367,In_1112);
nor U228 (N_228,In_941,In_39);
and U229 (N_229,In_78,In_886);
nor U230 (N_230,In_71,In_121);
or U231 (N_231,In_612,In_1955);
or U232 (N_232,In_415,In_945);
nor U233 (N_233,In_1636,In_1853);
nand U234 (N_234,In_473,In_1374);
nand U235 (N_235,In_1237,In_1200);
nor U236 (N_236,In_1331,In_105);
and U237 (N_237,In_375,In_1655);
and U238 (N_238,In_1134,In_1245);
or U239 (N_239,In_1971,In_1624);
xor U240 (N_240,In_1878,In_912);
nor U241 (N_241,In_247,In_1897);
xor U242 (N_242,In_320,In_1033);
and U243 (N_243,In_114,In_808);
or U244 (N_244,In_707,In_1578);
nand U245 (N_245,In_1640,In_1059);
and U246 (N_246,In_1841,In_1973);
or U247 (N_247,In_1233,In_230);
and U248 (N_248,In_1399,In_1820);
or U249 (N_249,In_1675,In_671);
nor U250 (N_250,In_716,In_466);
and U251 (N_251,In_1238,In_278);
nor U252 (N_252,In_1434,In_243);
and U253 (N_253,In_469,In_204);
nor U254 (N_254,In_1609,In_1226);
nand U255 (N_255,In_1538,In_1864);
and U256 (N_256,In_1993,In_1353);
nand U257 (N_257,In_1147,In_1994);
nand U258 (N_258,In_357,In_1302);
nor U259 (N_259,In_1224,In_1806);
or U260 (N_260,In_753,In_1673);
and U261 (N_261,In_1778,In_1802);
nand U262 (N_262,In_625,In_579);
xnor U263 (N_263,In_878,In_391);
nor U264 (N_264,In_1184,In_510);
nand U265 (N_265,In_1261,In_633);
xnor U266 (N_266,In_139,In_529);
xor U267 (N_267,In_747,In_1501);
nor U268 (N_268,In_742,In_33);
nand U269 (N_269,In_1592,In_572);
and U270 (N_270,In_1093,In_1092);
nor U271 (N_271,In_304,In_190);
nand U272 (N_272,In_170,In_1427);
nor U273 (N_273,In_18,In_444);
or U274 (N_274,In_822,In_223);
or U275 (N_275,In_768,In_1839);
nand U276 (N_276,In_565,In_991);
xnor U277 (N_277,In_260,In_638);
and U278 (N_278,In_1986,In_131);
nor U279 (N_279,In_1257,In_1629);
or U280 (N_280,In_1370,In_62);
nor U281 (N_281,In_228,In_1264);
nor U282 (N_282,In_25,In_563);
nand U283 (N_283,In_376,In_732);
and U284 (N_284,In_478,In_429);
nand U285 (N_285,In_1890,In_217);
nor U286 (N_286,In_609,In_1268);
or U287 (N_287,In_1892,In_387);
nand U288 (N_288,In_530,In_424);
nor U289 (N_289,In_158,In_19);
nand U290 (N_290,In_235,In_1697);
xor U291 (N_291,In_1143,In_1985);
nand U292 (N_292,In_1205,In_129);
nand U293 (N_293,In_371,In_1198);
or U294 (N_294,In_334,In_474);
and U295 (N_295,In_1410,In_1438);
nor U296 (N_296,In_1209,In_993);
xor U297 (N_297,In_1273,In_1430);
or U298 (N_298,In_1028,In_343);
or U299 (N_299,In_1140,In_14);
nand U300 (N_300,In_1854,In_1262);
nor U301 (N_301,In_1404,In_367);
xor U302 (N_302,In_1117,In_1267);
or U303 (N_303,In_1863,In_1083);
nand U304 (N_304,In_1392,In_1024);
nor U305 (N_305,In_1679,In_951);
nand U306 (N_306,In_643,In_338);
xnor U307 (N_307,In_1451,In_933);
nand U308 (N_308,In_403,In_1470);
nand U309 (N_309,In_430,In_789);
or U310 (N_310,In_737,In_1097);
nor U311 (N_311,In_544,In_7);
or U312 (N_312,In_748,In_422);
xor U313 (N_313,In_1779,In_1861);
and U314 (N_314,In_1512,In_866);
xor U315 (N_315,In_739,In_1494);
nand U316 (N_316,In_1645,In_658);
nand U317 (N_317,In_862,In_558);
or U318 (N_318,In_698,In_734);
or U319 (N_319,In_1313,In_881);
and U320 (N_320,In_94,In_794);
and U321 (N_321,In_1687,In_1620);
and U322 (N_322,In_175,In_1691);
and U323 (N_323,In_984,In_588);
or U324 (N_324,In_1287,In_185);
nand U325 (N_325,In_368,In_570);
nor U326 (N_326,In_22,In_248);
or U327 (N_327,In_1227,In_1128);
and U328 (N_328,In_1365,In_1270);
and U329 (N_329,In_1581,In_1107);
nand U330 (N_330,In_880,In_1713);
nand U331 (N_331,In_233,In_819);
or U332 (N_332,In_382,In_249);
nor U333 (N_333,In_162,In_290);
nor U334 (N_334,In_237,In_282);
or U335 (N_335,In_1646,In_340);
or U336 (N_336,In_1846,In_1384);
xnor U337 (N_337,In_298,In_1867);
and U338 (N_338,In_1961,In_1457);
or U339 (N_339,In_780,In_518);
or U340 (N_340,In_788,In_1468);
nor U341 (N_341,In_344,In_538);
and U342 (N_342,In_613,In_578);
nor U343 (N_343,In_562,In_551);
or U344 (N_344,In_594,In_1608);
nand U345 (N_345,In_1586,In_111);
nor U346 (N_346,In_1488,In_762);
xnor U347 (N_347,In_1177,In_977);
and U348 (N_348,In_684,In_611);
nor U349 (N_349,In_446,In_1064);
nor U350 (N_350,In_920,In_511);
nor U351 (N_351,In_1936,In_1913);
or U352 (N_352,In_784,In_1981);
xnor U353 (N_353,In_1393,In_1926);
and U354 (N_354,In_983,In_642);
nor U355 (N_355,In_132,In_149);
or U356 (N_356,In_691,In_173);
xor U357 (N_357,In_635,In_1517);
nor U358 (N_358,In_1263,In_1858);
nand U359 (N_359,In_962,In_1391);
nand U360 (N_360,In_76,In_1319);
or U361 (N_361,In_1989,In_1690);
or U362 (N_362,In_3,In_831);
or U363 (N_363,In_1271,In_1736);
nor U364 (N_364,In_83,In_1234);
nor U365 (N_365,In_353,In_1014);
nor U366 (N_366,In_1760,In_1605);
xor U367 (N_367,In_1157,In_724);
and U368 (N_368,In_1664,In_365);
nor U369 (N_369,In_1300,In_1545);
nand U370 (N_370,In_845,In_409);
nor U371 (N_371,In_319,In_148);
or U372 (N_372,In_704,In_624);
and U373 (N_373,In_1669,In_1834);
or U374 (N_374,In_1242,In_1991);
nor U375 (N_375,In_1461,In_987);
nor U376 (N_376,In_1688,In_180);
or U377 (N_377,In_1875,In_1813);
xor U378 (N_378,In_692,In_259);
nand U379 (N_379,In_1848,In_1560);
and U380 (N_380,In_373,In_341);
nand U381 (N_381,In_1027,In_85);
nand U382 (N_382,In_736,In_1650);
nand U383 (N_383,In_1787,In_1554);
nor U384 (N_384,In_580,In_508);
nor U385 (N_385,In_536,In_651);
and U386 (N_386,In_1100,In_307);
nor U387 (N_387,In_515,In_499);
nand U388 (N_388,In_1321,In_63);
or U389 (N_389,In_1400,In_1723);
nand U390 (N_390,In_42,In_53);
nand U391 (N_391,In_1114,In_1421);
xnor U392 (N_392,In_1980,In_1386);
and U393 (N_393,In_1463,In_41);
xor U394 (N_394,In_1192,In_905);
nand U395 (N_395,In_1509,In_1749);
or U396 (N_396,In_72,In_534);
nand U397 (N_397,In_1244,In_1557);
nor U398 (N_398,In_1852,In_1898);
nor U399 (N_399,In_1197,In_1901);
and U400 (N_400,In_191,In_1574);
and U401 (N_401,In_463,In_1912);
and U402 (N_402,In_160,In_1558);
nand U403 (N_403,In_1453,In_576);
or U404 (N_404,In_1150,In_1822);
xor U405 (N_405,In_777,In_336);
and U406 (N_406,In_289,In_1580);
or U407 (N_407,In_815,In_1739);
nand U408 (N_408,In_586,In_126);
nor U409 (N_409,In_1710,In_1389);
nand U410 (N_410,In_1223,In_1654);
and U411 (N_411,In_1774,In_1061);
nor U412 (N_412,In_1110,In_350);
or U413 (N_413,In_1102,In_632);
xor U414 (N_414,In_892,In_1454);
and U415 (N_415,In_791,In_1396);
nor U416 (N_416,In_687,In_285);
and U417 (N_417,In_1499,In_1309);
nand U418 (N_418,In_221,In_1330);
nand U419 (N_419,In_1626,In_956);
nand U420 (N_420,In_370,In_194);
or U421 (N_421,In_1698,In_924);
or U422 (N_422,In_639,In_939);
and U423 (N_423,In_1905,In_275);
nor U424 (N_424,In_1922,In_1591);
nor U425 (N_425,In_1403,In_269);
xnor U426 (N_426,In_441,In_1700);
nor U427 (N_427,In_535,In_1377);
and U428 (N_428,In_1135,In_1310);
or U429 (N_429,In_1601,In_1916);
and U430 (N_430,In_672,In_879);
nand U431 (N_431,In_493,In_186);
nor U432 (N_432,In_744,In_1450);
xor U433 (N_433,In_505,In_1823);
nand U434 (N_434,In_487,In_629);
nor U435 (N_435,In_1502,In_1153);
nor U436 (N_436,In_91,In_1831);
nor U437 (N_437,In_693,In_662);
xor U438 (N_438,In_918,In_450);
xnor U439 (N_439,In_550,In_460);
nor U440 (N_440,In_1478,In_873);
or U441 (N_441,In_1432,In_1159);
nand U442 (N_442,In_677,In_1906);
nand U443 (N_443,In_1167,In_756);
nor U444 (N_444,In_1345,In_246);
xnor U445 (N_445,In_1639,In_475);
nor U446 (N_446,In_730,In_929);
nor U447 (N_447,In_388,In_829);
xor U448 (N_448,In_1467,In_1219);
and U449 (N_449,In_1843,In_1612);
nor U450 (N_450,In_708,In_164);
and U451 (N_451,In_1705,In_1116);
and U452 (N_452,In_1422,In_1743);
nand U453 (N_453,In_623,In_870);
and U454 (N_454,In_408,In_200);
or U455 (N_455,In_823,In_1476);
and U456 (N_456,In_1879,In_1282);
and U457 (N_457,In_506,In_1336);
or U458 (N_458,In_295,In_1308);
xor U459 (N_459,In_655,In_618);
xnor U460 (N_460,In_1614,In_899);
nor U461 (N_461,In_1208,In_385);
or U462 (N_462,In_758,In_942);
or U463 (N_463,In_75,In_1695);
and U464 (N_464,In_1589,In_982);
and U465 (N_465,In_1962,In_733);
nor U466 (N_466,In_549,In_58);
or U467 (N_467,In_573,In_1369);
xor U468 (N_468,In_32,In_1941);
or U469 (N_469,In_1304,In_1104);
or U470 (N_470,In_1288,In_1395);
or U471 (N_471,In_1541,In_66);
or U472 (N_472,In_90,In_514);
nand U473 (N_473,In_410,In_1644);
nor U474 (N_474,In_178,In_384);
nor U475 (N_475,In_1363,In_1078);
and U476 (N_476,In_1339,In_1455);
and U477 (N_477,In_1155,In_79);
nor U478 (N_478,In_1615,In_1163);
xor U479 (N_479,In_1923,In_1976);
or U480 (N_480,In_871,In_431);
and U481 (N_481,In_1480,In_486);
and U482 (N_482,In_383,In_1034);
nand U483 (N_483,In_1741,In_330);
xor U484 (N_484,In_1759,In_472);
nand U485 (N_485,In_900,In_807);
xnor U486 (N_486,In_210,In_421);
or U487 (N_487,In_875,In_1069);
nor U488 (N_488,In_1446,In_1436);
nand U489 (N_489,In_142,In_377);
nor U490 (N_490,In_783,In_440);
nor U491 (N_491,In_597,In_20);
nor U492 (N_492,In_1284,In_1801);
nor U493 (N_493,In_1521,In_494);
nand U494 (N_494,In_1290,In_1529);
or U495 (N_495,In_1677,In_752);
nor U496 (N_496,In_1862,In_1842);
nor U497 (N_497,In_381,In_1401);
nand U498 (N_498,In_1067,In_315);
and U499 (N_499,In_24,In_57);
and U500 (N_500,In_454,In_363);
nor U501 (N_501,In_1007,In_1500);
nand U502 (N_502,In_614,In_1711);
or U503 (N_503,In_1662,In_1566);
and U504 (N_504,In_1332,In_1216);
nor U505 (N_505,In_909,In_1656);
xnor U506 (N_506,In_206,In_351);
or U507 (N_507,In_503,In_1888);
xnor U508 (N_508,In_1773,In_1895);
nor U509 (N_509,In_1719,In_827);
nor U510 (N_510,In_751,In_755);
xor U511 (N_511,In_1516,In_171);
xnor U512 (N_512,In_1546,In_1411);
xnor U513 (N_513,In_1567,In_574);
nor U514 (N_514,In_1483,In_1138);
or U515 (N_515,In_242,In_1131);
and U516 (N_516,In_1505,In_427);
and U517 (N_517,In_599,In_1256);
nor U518 (N_518,In_1023,In_927);
nor U519 (N_519,In_1660,In_48);
nor U520 (N_520,In_627,In_1046);
xnor U521 (N_521,In_154,In_1995);
xor U522 (N_522,In_680,In_281);
nand U523 (N_523,In_676,In_1693);
or U524 (N_524,In_1533,In_1049);
xnor U525 (N_525,In_100,In_1212);
xor U526 (N_526,In_1709,In_865);
nor U527 (N_527,In_593,In_1496);
xnor U528 (N_528,In_199,In_891);
xnor U529 (N_529,In_826,In_1775);
xor U530 (N_530,In_876,In_1810);
and U531 (N_531,In_1670,In_56);
nor U532 (N_532,In_1265,In_272);
nand U533 (N_533,In_433,In_1530);
nor U534 (N_534,In_1259,In_1094);
or U535 (N_535,In_1185,In_719);
nor U536 (N_536,In_921,In_940);
nand U537 (N_537,In_1988,In_1426);
and U538 (N_538,In_1232,In_972);
and U539 (N_539,In_652,In_973);
or U540 (N_540,In_999,In_1038);
nand U541 (N_541,In_1997,In_193);
or U542 (N_542,In_361,In_735);
or U543 (N_543,In_1893,In_455);
nand U544 (N_544,In_816,In_1156);
or U545 (N_545,In_181,In_386);
or U546 (N_546,In_1456,In_1531);
or U547 (N_547,In_1358,In_1689);
nand U548 (N_548,In_209,In_1850);
and U549 (N_549,In_1133,In_1729);
and U550 (N_550,In_971,In_1166);
and U551 (N_551,In_1335,In_346);
nor U552 (N_552,In_113,In_226);
xnor U553 (N_553,In_837,In_797);
or U554 (N_554,In_1180,In_723);
and U555 (N_555,In_545,In_1235);
or U556 (N_556,In_16,In_1766);
xnor U557 (N_557,In_1738,In_848);
nor U558 (N_558,In_1829,In_187);
and U559 (N_559,In_1073,In_1648);
or U560 (N_560,In_1459,In_699);
and U561 (N_561,In_1631,In_348);
xnor U562 (N_562,In_1931,In_582);
xnor U563 (N_563,In_443,In_49);
or U564 (N_564,In_219,In_1280);
nor U565 (N_565,In_504,In_1354);
and U566 (N_566,In_465,In_1295);
xor U567 (N_567,In_1071,In_1996);
nand U568 (N_568,In_1489,In_1755);
and U569 (N_569,In_1561,In_1004);
and U570 (N_570,In_156,In_270);
and U571 (N_571,In_986,In_1055);
nand U572 (N_572,In_907,In_860);
nor U573 (N_573,In_1296,In_1730);
nand U574 (N_574,In_1579,In_398);
or U575 (N_575,In_805,In_1757);
nor U576 (N_576,In_1003,In_1838);
xor U577 (N_577,In_557,In_480);
and U578 (N_578,In_1676,In_713);
or U579 (N_579,In_277,In_1022);
and U580 (N_580,In_189,In_1402);
nand U581 (N_581,In_1945,In_1712);
xor U582 (N_582,In_1939,In_1246);
and U583 (N_583,In_224,In_1041);
nor U584 (N_584,In_1814,In_571);
nor U585 (N_585,In_1935,In_1009);
nor U586 (N_586,In_1347,In_397);
nor U587 (N_587,In_267,In_998);
and U588 (N_588,In_1825,In_512);
nand U589 (N_589,In_1725,In_1366);
nor U590 (N_590,In_396,In_1460);
or U591 (N_591,In_811,In_932);
nor U592 (N_592,In_1548,In_1781);
or U593 (N_593,In_520,In_770);
nand U594 (N_594,In_745,In_1341);
or U595 (N_595,In_1894,In_358);
or U596 (N_596,In_641,In_1006);
nor U597 (N_597,In_1885,In_405);
nand U598 (N_598,In_1904,In_253);
or U599 (N_599,In_1058,In_547);
nor U600 (N_600,In_720,In_1344);
xor U601 (N_601,In_1048,In_975);
nand U602 (N_602,In_54,In_1266);
nor U603 (N_603,In_653,In_867);
or U604 (N_604,In_1942,In_1817);
and U605 (N_605,In_1717,In_321);
nor U606 (N_606,In_1086,In_1379);
nand U607 (N_607,In_167,In_468);
nand U608 (N_608,In_1407,In_1462);
or U609 (N_609,In_1667,In_261);
xor U610 (N_610,In_73,In_81);
nand U611 (N_611,In_1628,In_1178);
xor U612 (N_612,In_725,In_681);
nor U613 (N_613,In_650,In_232);
or U614 (N_614,In_309,In_135);
nand U615 (N_615,In_1576,In_1968);
or U616 (N_616,In_1657,In_451);
or U617 (N_617,In_389,In_1291);
nor U618 (N_618,In_482,In_26);
xor U619 (N_619,In_799,In_1969);
and U620 (N_620,In_785,In_134);
xnor U621 (N_621,In_1486,In_1303);
or U622 (N_622,In_670,In_125);
nor U623 (N_623,In_1274,In_311);
and U624 (N_624,In_528,In_1724);
nor U625 (N_625,In_1606,In_935);
nor U626 (N_626,In_214,In_314);
or U627 (N_627,In_1479,In_517);
or U628 (N_628,In_107,In_1017);
and U629 (N_629,In_1145,In_1137);
or U630 (N_630,In_798,In_273);
or U631 (N_631,In_1179,In_1527);
nor U632 (N_632,In_1194,In_1767);
and U633 (N_633,In_65,In_1008);
nor U634 (N_634,In_1211,In_898);
and U635 (N_635,In_637,In_116);
xnor U636 (N_636,In_585,In_256);
and U637 (N_637,In_1562,In_1949);
and U638 (N_638,In_1506,In_395);
or U639 (N_639,In_606,In_925);
or U640 (N_640,In_136,In_1668);
xor U641 (N_641,In_1065,In_832);
or U642 (N_642,In_501,In_159);
or U643 (N_643,In_910,In_1722);
nor U644 (N_644,In_364,In_587);
or U645 (N_645,In_406,In_1348);
xor U646 (N_646,In_1564,In_118);
nor U647 (N_647,In_1169,In_1015);
or U648 (N_648,In_1435,In_619);
or U649 (N_649,In_1441,In_568);
and U650 (N_650,In_996,In_84);
xnor U651 (N_651,In_934,In_417);
nor U652 (N_652,In_1241,In_543);
xnor U653 (N_653,In_1613,In_456);
and U654 (N_654,In_1087,In_931);
and U655 (N_655,In_117,In_317);
nor U656 (N_656,In_555,In_400);
nor U657 (N_657,In_112,In_448);
or U658 (N_658,In_1731,In_965);
and U659 (N_659,In_631,In_1325);
xor U660 (N_660,In_1109,In_781);
and U661 (N_661,In_1020,In_1277);
xnor U662 (N_662,In_331,In_263);
xor U663 (N_663,In_106,In_1373);
or U664 (N_664,In_542,In_608);
and U665 (N_665,In_52,In_1297);
nand U666 (N_666,In_1694,In_109);
xnor U667 (N_667,In_1750,In_592);
nand U668 (N_668,In_1495,In_1418);
nor U669 (N_669,In_647,In_435);
and U670 (N_670,In_1101,In_1957);
xor U671 (N_671,In_1835,In_1570);
and U672 (N_672,In_1799,In_402);
nor U673 (N_673,In_1671,In_1665);
or U674 (N_674,In_1836,In_92);
xor U675 (N_675,In_1790,In_38);
xor U676 (N_676,In_46,In_1872);
and U677 (N_677,In_325,In_1318);
nand U678 (N_678,In_904,In_1276);
or U679 (N_679,In_150,In_1543);
xor U680 (N_680,In_882,In_1849);
nand U681 (N_681,In_759,In_715);
nor U682 (N_682,In_868,In_946);
nor U683 (N_683,In_569,In_1206);
nand U684 (N_684,In_1152,In_754);
or U685 (N_685,In_1634,In_1868);
and U686 (N_686,In_792,In_489);
xor U687 (N_687,In_35,In_1915);
xnor U688 (N_688,In_1754,In_796);
nor U689 (N_689,In_590,In_1740);
or U690 (N_690,In_1784,In_1727);
or U691 (N_691,In_299,In_961);
or U692 (N_692,In_853,In_1098);
and U693 (N_693,In_564,In_656);
nand U694 (N_694,In_1681,In_360);
or U695 (N_695,In_846,In_779);
nand U696 (N_696,In_894,In_1786);
or U697 (N_697,In_202,In_211);
nor U698 (N_698,In_1607,In_355);
or U699 (N_699,In_1824,In_1040);
nor U700 (N_700,In_1575,In_1139);
nor U701 (N_701,In_976,In_1122);
nand U702 (N_702,In_1091,In_1940);
nand U703 (N_703,In_306,In_1785);
xnor U704 (N_704,In_467,In_327);
nand U705 (N_705,In_140,In_696);
or U706 (N_706,In_1126,In_1068);
and U707 (N_707,In_1333,In_820);
nor U708 (N_708,In_872,In_163);
nand U709 (N_709,In_1752,In_1141);
nand U710 (N_710,In_559,In_1283);
xnor U711 (N_711,In_1503,In_1990);
xnor U712 (N_712,In_1381,In_362);
or U713 (N_713,In_1532,In_1472);
xor U714 (N_714,In_1658,In_1364);
nand U715 (N_715,In_258,In_1044);
and U716 (N_716,In_366,In_1523);
or U717 (N_717,In_1753,In_459);
nor U718 (N_718,In_1444,In_1886);
nand U719 (N_719,In_1583,In_533);
nand U720 (N_720,In_1518,In_1776);
xnor U721 (N_721,In_1445,In_337);
or U722 (N_722,In_896,In_305);
nand U723 (N_723,In_721,In_1889);
or U724 (N_724,In_390,In_1099);
xnor U725 (N_725,In_1002,In_1920);
nor U726 (N_726,In_1584,In_119);
nor U727 (N_727,In_1525,In_130);
or U728 (N_728,In_1796,In_1204);
and U729 (N_729,In_1899,In_1442);
nor U730 (N_730,In_1464,In_1818);
or U731 (N_731,In_1514,In_507);
nor U732 (N_732,In_1550,In_1908);
xor U733 (N_733,In_1089,In_1821);
and U734 (N_734,In_1433,In_1641);
xor U735 (N_735,In_1728,In_1255);
nor U736 (N_736,In_601,In_963);
nand U737 (N_737,In_776,In_1096);
xor U738 (N_738,In_1301,In_1183);
nor U739 (N_739,In_301,In_1361);
or U740 (N_740,In_1952,In_913);
and U741 (N_741,In_1084,In_1937);
and U742 (N_742,In_1230,In_302);
nand U743 (N_743,In_649,In_1855);
or U744 (N_744,In_1610,In_1637);
and U745 (N_745,In_840,In_70);
nor U746 (N_746,In_1189,In_1119);
and U747 (N_747,In_667,In_36);
and U748 (N_748,In_700,In_434);
and U749 (N_749,In_404,In_1805);
nor U750 (N_750,In_1944,In_88);
and U751 (N_751,In_531,In_335);
or U752 (N_752,In_903,In_1409);
and U753 (N_753,In_1465,In_771);
and U754 (N_754,In_276,In_985);
nor U755 (N_755,In_1186,In_1001);
nor U756 (N_756,In_1678,In_856);
xor U757 (N_757,In_964,In_1763);
and U758 (N_758,In_1565,In_523);
and U759 (N_759,In_115,In_103);
nor U760 (N_760,In_461,In_790);
xnor U761 (N_761,In_197,In_1039);
or U762 (N_762,In_169,In_1537);
or U763 (N_763,In_1764,In_1387);
nand U764 (N_764,In_661,In_491);
nand U765 (N_765,In_188,In_1599);
xor U766 (N_766,In_665,In_1871);
xnor U767 (N_767,In_1771,In_974);
or U768 (N_768,In_1674,In_817);
nor U769 (N_769,In_1921,In_207);
or U770 (N_770,In_323,In_1965);
and U771 (N_771,In_1770,In_310);
nand U772 (N_772,In_288,In_1643);
nor U773 (N_773,In_1887,In_1520);
nand U774 (N_774,In_1252,In_1032);
and U775 (N_775,In_215,In_1088);
xnor U776 (N_776,In_1998,In_198);
and U777 (N_777,In_666,In_1844);
or U778 (N_778,In_1746,In_152);
or U779 (N_779,In_532,In_648);
or U780 (N_780,In_1633,In_858);
or U781 (N_781,In_1191,In_1247);
nand U782 (N_782,In_205,In_1549);
nor U783 (N_783,In_1555,In_566);
or U784 (N_784,In_28,In_1847);
and U785 (N_785,In_266,In_399);
nand U786 (N_786,In_1010,In_1958);
nand U787 (N_787,In_265,In_1337);
nor U788 (N_788,In_183,In_1449);
and U789 (N_789,In_1663,In_1324);
nor U790 (N_790,In_825,In_61);
xnor U791 (N_791,In_8,In_133);
nor U792 (N_792,In_245,In_967);
nor U793 (N_793,In_1342,In_1146);
or U794 (N_794,In_498,In_978);
nor U795 (N_795,In_804,In_701);
or U796 (N_796,In_1106,In_2);
nor U797 (N_797,In_689,In_1547);
xnor U798 (N_798,In_1240,In_495);
and U799 (N_799,In_208,In_1026);
nor U800 (N_800,In_1881,In_485);
nand U801 (N_801,In_407,In_423);
xnor U802 (N_802,In_1702,In_1782);
xnor U803 (N_803,In_1826,In_68);
nor U804 (N_804,In_1508,In_1228);
and U805 (N_805,In_312,In_897);
nor U806 (N_806,In_1162,In_1907);
nor U807 (N_807,In_1111,In_1524);
xor U808 (N_808,In_177,In_303);
or U809 (N_809,In_1807,In_1984);
or U810 (N_810,In_1528,In_144);
or U811 (N_811,In_749,In_436);
and U812 (N_812,In_413,In_174);
nand U813 (N_813,In_1279,In_800);
or U814 (N_814,In_77,In_1732);
nand U815 (N_815,In_1452,In_1974);
nand U816 (N_816,In_1651,In_1963);
nor U817 (N_817,In_821,In_769);
nor U818 (N_818,In_128,In_1414);
nor U819 (N_819,In_244,In_890);
nor U820 (N_820,In_1783,In_44);
nand U821 (N_821,In_1803,In_50);
and U822 (N_822,In_1293,In_5);
xnor U823 (N_823,In_526,In_1160);
xor U824 (N_824,In_1845,In_1737);
or U825 (N_825,In_1193,In_630);
and U826 (N_826,In_1720,In_1869);
xor U827 (N_827,In_1161,In_1413);
xnor U828 (N_828,In_11,In_1394);
or U829 (N_829,In_1258,In_1120);
and U830 (N_830,In_1144,In_225);
xnor U831 (N_831,In_143,In_464);
and U832 (N_832,In_380,In_1029);
and U833 (N_833,In_548,In_1306);
nor U834 (N_834,In_607,In_855);
and U835 (N_835,In_264,In_760);
nand U836 (N_836,In_212,In_1927);
nand U837 (N_837,In_195,In_82);
and U838 (N_838,In_1793,In_688);
nor U839 (N_839,In_99,In_1243);
nand U840 (N_840,In_835,In_1573);
and U841 (N_841,In_1652,In_1054);
xor U842 (N_842,In_1317,In_432);
xor U843 (N_843,In_1638,In_657);
nand U844 (N_844,In_522,In_356);
nor U845 (N_845,In_293,In_439);
xnor U846 (N_846,In_854,In_741);
xnor U847 (N_847,In_1703,In_166);
nor U848 (N_848,In_1220,In_1338);
nor U849 (N_849,In_604,In_420);
or U850 (N_850,In_556,In_1222);
and U851 (N_851,In_1172,In_1149);
nand U852 (N_852,In_1081,In_674);
nand U853 (N_853,In_970,In_40);
xnor U854 (N_854,In_1622,In_521);
xnor U855 (N_855,In_95,In_1311);
nand U856 (N_856,In_1000,In_795);
xor U857 (N_857,In_1469,In_874);
and U858 (N_858,In_4,In_1704);
nor U859 (N_859,In_1052,In_1362);
xnor U860 (N_860,In_1751,In_1964);
and U861 (N_861,In_1349,In_1588);
nand U862 (N_862,In_1056,In_1795);
xnor U863 (N_863,In_1934,In_1047);
nand U864 (N_864,In_988,In_1305);
and U865 (N_865,In_1217,In_1577);
xnor U866 (N_866,In_254,In_1756);
xnor U867 (N_867,In_1005,In_1827);
and U868 (N_868,In_284,In_1616);
and U869 (N_869,In_1203,In_1326);
or U870 (N_870,In_1649,In_300);
and U871 (N_871,In_861,In_1582);
nor U872 (N_872,In_322,In_889);
xor U873 (N_873,In_1195,In_1551);
xnor U874 (N_874,In_1672,In_1207);
or U875 (N_875,In_509,In_393);
nor U876 (N_876,In_683,In_1154);
or U877 (N_877,In_1350,In_1618);
xor U878 (N_878,In_1168,In_12);
xnor U879 (N_879,In_1423,In_1074);
nand U880 (N_880,In_1978,In_1323);
and U881 (N_881,In_1635,In_1539);
nand U882 (N_882,In_379,In_893);
and U883 (N_883,In_1487,In_1765);
or U884 (N_884,In_602,In_1355);
and U885 (N_885,In_1593,In_778);
nand U886 (N_886,In_392,In_1190);
and U887 (N_887,In_1115,In_1181);
nor U888 (N_888,In_1603,In_1987);
xnor U889 (N_889,In_122,In_1866);
or U890 (N_890,In_27,In_1800);
and U891 (N_891,In_793,In_0);
xnor U892 (N_892,In_1661,In_911);
nand U893 (N_893,In_1966,In_1809);
and U894 (N_894,In_483,In_926);
or U895 (N_895,In_703,In_1352);
nand U896 (N_896,In_1375,In_1063);
nand U897 (N_897,In_997,In_709);
xnor U898 (N_898,In_1621,In_738);
nand U899 (N_899,In_1477,In_943);
and U900 (N_900,In_1036,In_1250);
xnor U901 (N_901,In_1299,In_1568);
xnor U902 (N_902,In_806,In_1772);
nor U903 (N_903,In_1466,In_349);
nand U904 (N_904,In_646,In_928);
or U905 (N_905,In_1625,In_416);
or U906 (N_906,In_1385,In_836);
and U907 (N_907,In_179,In_1683);
nand U908 (N_908,In_15,In_123);
nor U909 (N_909,In_1860,In_458);
xor U910 (N_910,In_120,In_1544);
nand U911 (N_911,In_316,In_969);
nand U912 (N_912,In_1383,In_966);
or U913 (N_913,In_1535,In_1943);
or U914 (N_914,In_227,In_685);
nor U915 (N_915,In_813,In_274);
xor U916 (N_916,In_990,In_802);
and U917 (N_917,In_1788,In_1992);
xnor U918 (N_918,In_1967,In_669);
nor U919 (N_919,In_598,In_1910);
nor U920 (N_920,In_1552,In_1569);
nor U921 (N_921,In_675,In_394);
and U922 (N_922,In_1359,In_883);
or U923 (N_923,In_621,In_1103);
xnor U924 (N_924,In_1447,In_1113);
nor U925 (N_925,In_947,In_1946);
nor U926 (N_926,In_615,In_636);
nand U927 (N_927,In_419,In_1929);
nand U928 (N_928,In_610,In_1744);
or U929 (N_929,In_553,In_839);
or U930 (N_930,In_1597,In_401);
or U931 (N_931,In_1249,In_102);
nor U932 (N_932,In_352,In_1882);
xor U933 (N_933,In_786,In_1716);
and U934 (N_934,In_1522,In_1043);
xnor U935 (N_935,In_1747,In_1706);
nand U936 (N_936,In_705,In_1859);
xor U937 (N_937,In_513,In_722);
nor U938 (N_938,In_992,In_89);
nand U939 (N_939,In_1085,In_1351);
or U940 (N_940,In_1865,In_1627);
xnor U941 (N_941,In_153,In_519);
and U942 (N_942,In_1492,In_1590);
and U943 (N_943,In_1485,In_1718);
nand U944 (N_944,In_240,In_887);
xnor U945 (N_945,In_1057,In_332);
and U946 (N_946,In_1600,In_1199);
nor U947 (N_947,In_418,In_101);
nor U948 (N_948,In_678,In_765);
xor U949 (N_949,In_810,In_1960);
and U950 (N_950,In_1408,In_1870);
nor U951 (N_951,In_1534,In_438);
nand U952 (N_952,In_374,In_980);
nand U953 (N_953,In_809,In_1642);
nand U954 (N_954,In_686,In_728);
nand U955 (N_955,In_833,In_492);
nand U956 (N_956,In_1982,In_1513);
and U957 (N_957,In_151,In_1066);
and U958 (N_958,In_1294,In_414);
nand U959 (N_959,In_1142,In_1050);
nand U960 (N_960,In_1406,In_844);
and U961 (N_961,In_944,In_828);
nor U962 (N_962,In_644,In_98);
nor U963 (N_963,In_1202,In_958);
or U964 (N_964,In_1745,In_1830);
nand U965 (N_965,In_989,In_1808);
nand U966 (N_966,In_1275,In_1082);
nand U967 (N_967,In_583,In_690);
and U968 (N_968,In_729,In_425);
nor U969 (N_969,In_527,In_1542);
nor U970 (N_970,In_1571,In_812);
nor U971 (N_971,In_1253,In_1031);
and U972 (N_972,In_1320,In_1924);
nand U973 (N_973,In_859,In_1429);
or U974 (N_974,In_1175,In_949);
or U975 (N_975,In_1260,In_561);
nor U976 (N_976,In_801,In_1707);
nand U977 (N_977,In_937,In_1733);
and U978 (N_978,In_500,In_540);
xor U979 (N_979,In_324,In_1876);
or U980 (N_980,In_1380,In_589);
and U981 (N_981,In_1682,In_916);
nor U982 (N_982,In_1289,In_147);
xnor U983 (N_983,In_255,In_1077);
nor U984 (N_984,In_955,In_239);
nand U985 (N_985,In_1507,In_834);
xnor U986 (N_986,In_1225,In_1315);
nor U987 (N_987,In_849,In_1397);
and U988 (N_988,In_1832,In_297);
nand U989 (N_989,In_1708,In_575);
or U990 (N_990,In_1928,In_1229);
nand U991 (N_991,In_1497,In_67);
nand U992 (N_992,In_339,In_1540);
xor U993 (N_993,In_525,In_146);
nor U994 (N_994,In_731,In_59);
and U995 (N_995,In_979,In_923);
nand U996 (N_996,In_96,In_1792);
or U997 (N_997,In_1165,In_567);
nand U998 (N_998,In_714,In_1917);
and U999 (N_999,In_161,In_695);
nand U1000 (N_1000,In_535,In_655);
and U1001 (N_1001,In_1006,In_53);
and U1002 (N_1002,In_1611,In_370);
nand U1003 (N_1003,In_246,In_1600);
nor U1004 (N_1004,In_47,In_815);
nor U1005 (N_1005,In_1306,In_1896);
nand U1006 (N_1006,In_1125,In_254);
nor U1007 (N_1007,In_316,In_1468);
nand U1008 (N_1008,In_1861,In_1767);
xnor U1009 (N_1009,In_1608,In_1990);
and U1010 (N_1010,In_100,In_129);
xnor U1011 (N_1011,In_1503,In_1499);
and U1012 (N_1012,In_1584,In_1228);
xnor U1013 (N_1013,In_1297,In_1119);
nand U1014 (N_1014,In_47,In_1736);
xnor U1015 (N_1015,In_962,In_1396);
and U1016 (N_1016,In_1438,In_258);
nand U1017 (N_1017,In_712,In_1071);
nand U1018 (N_1018,In_223,In_1561);
nand U1019 (N_1019,In_1726,In_123);
nand U1020 (N_1020,In_412,In_118);
or U1021 (N_1021,In_1190,In_1311);
or U1022 (N_1022,In_1024,In_1989);
or U1023 (N_1023,In_1269,In_158);
nor U1024 (N_1024,In_1784,In_1285);
or U1025 (N_1025,In_1984,In_605);
and U1026 (N_1026,In_488,In_629);
or U1027 (N_1027,In_554,In_1394);
xnor U1028 (N_1028,In_768,In_815);
xnor U1029 (N_1029,In_27,In_1159);
nor U1030 (N_1030,In_1376,In_1535);
nand U1031 (N_1031,In_419,In_834);
xor U1032 (N_1032,In_333,In_1479);
and U1033 (N_1033,In_1557,In_1232);
or U1034 (N_1034,In_1160,In_362);
and U1035 (N_1035,In_1674,In_619);
nand U1036 (N_1036,In_100,In_1558);
and U1037 (N_1037,In_158,In_733);
nand U1038 (N_1038,In_372,In_957);
or U1039 (N_1039,In_1965,In_741);
and U1040 (N_1040,In_930,In_739);
or U1041 (N_1041,In_584,In_572);
xnor U1042 (N_1042,In_23,In_1415);
nor U1043 (N_1043,In_65,In_1053);
and U1044 (N_1044,In_242,In_1834);
xor U1045 (N_1045,In_174,In_1241);
and U1046 (N_1046,In_1644,In_581);
nand U1047 (N_1047,In_1280,In_757);
nand U1048 (N_1048,In_1054,In_1585);
nand U1049 (N_1049,In_1119,In_1644);
nor U1050 (N_1050,In_1244,In_1869);
or U1051 (N_1051,In_1459,In_463);
nor U1052 (N_1052,In_1259,In_1052);
and U1053 (N_1053,In_1561,In_283);
nand U1054 (N_1054,In_1241,In_877);
nand U1055 (N_1055,In_773,In_887);
xor U1056 (N_1056,In_980,In_1443);
nand U1057 (N_1057,In_4,In_992);
xnor U1058 (N_1058,In_1769,In_1084);
nand U1059 (N_1059,In_1988,In_873);
or U1060 (N_1060,In_1882,In_743);
nand U1061 (N_1061,In_434,In_1956);
nand U1062 (N_1062,In_1197,In_507);
or U1063 (N_1063,In_232,In_367);
xnor U1064 (N_1064,In_868,In_1863);
xor U1065 (N_1065,In_1150,In_1601);
nor U1066 (N_1066,In_1888,In_957);
xor U1067 (N_1067,In_1361,In_869);
or U1068 (N_1068,In_452,In_179);
xnor U1069 (N_1069,In_1834,In_1991);
and U1070 (N_1070,In_339,In_470);
nand U1071 (N_1071,In_631,In_209);
and U1072 (N_1072,In_1933,In_1503);
xor U1073 (N_1073,In_1978,In_594);
and U1074 (N_1074,In_1837,In_432);
nand U1075 (N_1075,In_1674,In_493);
and U1076 (N_1076,In_680,In_1970);
nand U1077 (N_1077,In_1928,In_404);
nand U1078 (N_1078,In_541,In_1920);
nand U1079 (N_1079,In_491,In_604);
xnor U1080 (N_1080,In_576,In_1783);
nor U1081 (N_1081,In_1431,In_339);
nand U1082 (N_1082,In_47,In_416);
xnor U1083 (N_1083,In_415,In_656);
nor U1084 (N_1084,In_1688,In_1782);
or U1085 (N_1085,In_1607,In_1301);
and U1086 (N_1086,In_544,In_1542);
nand U1087 (N_1087,In_585,In_1358);
and U1088 (N_1088,In_1739,In_346);
or U1089 (N_1089,In_1341,In_1042);
and U1090 (N_1090,In_1740,In_1776);
nor U1091 (N_1091,In_898,In_1604);
nand U1092 (N_1092,In_1750,In_508);
nor U1093 (N_1093,In_162,In_102);
nor U1094 (N_1094,In_1902,In_1720);
xnor U1095 (N_1095,In_1764,In_889);
nand U1096 (N_1096,In_1723,In_1783);
nand U1097 (N_1097,In_601,In_4);
or U1098 (N_1098,In_1958,In_1352);
nor U1099 (N_1099,In_160,In_100);
nor U1100 (N_1100,In_637,In_1570);
and U1101 (N_1101,In_898,In_518);
and U1102 (N_1102,In_126,In_415);
nand U1103 (N_1103,In_184,In_735);
and U1104 (N_1104,In_618,In_192);
xnor U1105 (N_1105,In_451,In_285);
nand U1106 (N_1106,In_383,In_186);
or U1107 (N_1107,In_437,In_276);
nor U1108 (N_1108,In_1220,In_603);
nand U1109 (N_1109,In_866,In_1761);
nor U1110 (N_1110,In_1708,In_1527);
nand U1111 (N_1111,In_274,In_1132);
xnor U1112 (N_1112,In_519,In_305);
nor U1113 (N_1113,In_189,In_1890);
and U1114 (N_1114,In_1131,In_691);
or U1115 (N_1115,In_1972,In_23);
nand U1116 (N_1116,In_1738,In_1348);
nor U1117 (N_1117,In_1467,In_444);
xor U1118 (N_1118,In_672,In_844);
xnor U1119 (N_1119,In_553,In_956);
nand U1120 (N_1120,In_600,In_807);
xor U1121 (N_1121,In_1096,In_1015);
or U1122 (N_1122,In_860,In_1183);
xnor U1123 (N_1123,In_1567,In_988);
xor U1124 (N_1124,In_1223,In_765);
nand U1125 (N_1125,In_799,In_887);
xnor U1126 (N_1126,In_35,In_1310);
and U1127 (N_1127,In_1701,In_30);
xnor U1128 (N_1128,In_1120,In_1509);
xnor U1129 (N_1129,In_661,In_1144);
nor U1130 (N_1130,In_1105,In_1791);
nor U1131 (N_1131,In_1772,In_153);
nand U1132 (N_1132,In_1900,In_44);
or U1133 (N_1133,In_1435,In_1478);
or U1134 (N_1134,In_79,In_503);
xnor U1135 (N_1135,In_1726,In_992);
nor U1136 (N_1136,In_1546,In_1518);
xnor U1137 (N_1137,In_1058,In_1168);
xnor U1138 (N_1138,In_1275,In_372);
nor U1139 (N_1139,In_1435,In_1176);
xnor U1140 (N_1140,In_677,In_683);
nor U1141 (N_1141,In_478,In_230);
and U1142 (N_1142,In_1252,In_1807);
and U1143 (N_1143,In_802,In_958);
xnor U1144 (N_1144,In_1142,In_24);
nand U1145 (N_1145,In_388,In_1119);
or U1146 (N_1146,In_786,In_1427);
xor U1147 (N_1147,In_718,In_532);
and U1148 (N_1148,In_1589,In_301);
nand U1149 (N_1149,In_463,In_840);
xor U1150 (N_1150,In_13,In_238);
and U1151 (N_1151,In_1353,In_627);
nand U1152 (N_1152,In_1679,In_500);
xnor U1153 (N_1153,In_1880,In_429);
or U1154 (N_1154,In_1617,In_533);
or U1155 (N_1155,In_152,In_456);
and U1156 (N_1156,In_1005,In_1187);
xor U1157 (N_1157,In_879,In_1342);
or U1158 (N_1158,In_423,In_1276);
and U1159 (N_1159,In_1670,In_770);
nor U1160 (N_1160,In_887,In_1752);
nand U1161 (N_1161,In_1683,In_1615);
nand U1162 (N_1162,In_1547,In_1709);
xnor U1163 (N_1163,In_1445,In_1756);
xnor U1164 (N_1164,In_111,In_1873);
nor U1165 (N_1165,In_1397,In_294);
xor U1166 (N_1166,In_397,In_264);
and U1167 (N_1167,In_1154,In_1765);
or U1168 (N_1168,In_1129,In_1339);
nor U1169 (N_1169,In_1608,In_417);
and U1170 (N_1170,In_1697,In_1727);
nand U1171 (N_1171,In_910,In_558);
nand U1172 (N_1172,In_156,In_982);
xor U1173 (N_1173,In_451,In_740);
or U1174 (N_1174,In_85,In_1784);
nor U1175 (N_1175,In_633,In_1387);
and U1176 (N_1176,In_565,In_5);
and U1177 (N_1177,In_560,In_408);
nand U1178 (N_1178,In_1365,In_1290);
and U1179 (N_1179,In_1001,In_1675);
xnor U1180 (N_1180,In_856,In_1235);
nand U1181 (N_1181,In_1592,In_1880);
xnor U1182 (N_1182,In_23,In_1729);
nand U1183 (N_1183,In_1123,In_1447);
or U1184 (N_1184,In_1819,In_1526);
nand U1185 (N_1185,In_1331,In_1823);
xor U1186 (N_1186,In_637,In_1340);
nand U1187 (N_1187,In_693,In_1562);
and U1188 (N_1188,In_371,In_1481);
nor U1189 (N_1189,In_1398,In_427);
and U1190 (N_1190,In_610,In_1660);
and U1191 (N_1191,In_1962,In_1738);
or U1192 (N_1192,In_1351,In_1300);
or U1193 (N_1193,In_752,In_1479);
and U1194 (N_1194,In_1672,In_535);
xor U1195 (N_1195,In_758,In_1727);
nor U1196 (N_1196,In_928,In_1678);
nand U1197 (N_1197,In_1153,In_1947);
xnor U1198 (N_1198,In_633,In_1042);
and U1199 (N_1199,In_431,In_1016);
or U1200 (N_1200,In_392,In_1115);
xor U1201 (N_1201,In_932,In_1004);
and U1202 (N_1202,In_621,In_1647);
and U1203 (N_1203,In_712,In_653);
nor U1204 (N_1204,In_1073,In_1733);
xor U1205 (N_1205,In_977,In_508);
nand U1206 (N_1206,In_391,In_532);
nand U1207 (N_1207,In_1205,In_1909);
or U1208 (N_1208,In_688,In_627);
and U1209 (N_1209,In_1944,In_1237);
nand U1210 (N_1210,In_1196,In_1623);
xor U1211 (N_1211,In_1729,In_181);
and U1212 (N_1212,In_1534,In_321);
nor U1213 (N_1213,In_1280,In_529);
xor U1214 (N_1214,In_1849,In_419);
nor U1215 (N_1215,In_1581,In_715);
nand U1216 (N_1216,In_686,In_882);
nand U1217 (N_1217,In_831,In_477);
nand U1218 (N_1218,In_429,In_1732);
xnor U1219 (N_1219,In_1494,In_1817);
nor U1220 (N_1220,In_1150,In_1376);
nor U1221 (N_1221,In_1071,In_1889);
nor U1222 (N_1222,In_313,In_342);
nand U1223 (N_1223,In_1398,In_1154);
nor U1224 (N_1224,In_1276,In_1596);
nand U1225 (N_1225,In_2,In_310);
nand U1226 (N_1226,In_1461,In_547);
xor U1227 (N_1227,In_99,In_1807);
and U1228 (N_1228,In_1473,In_1479);
or U1229 (N_1229,In_225,In_1293);
and U1230 (N_1230,In_1061,In_947);
and U1231 (N_1231,In_1748,In_826);
and U1232 (N_1232,In_1916,In_1578);
or U1233 (N_1233,In_1534,In_947);
nand U1234 (N_1234,In_1716,In_1812);
or U1235 (N_1235,In_38,In_1892);
or U1236 (N_1236,In_1167,In_987);
nand U1237 (N_1237,In_882,In_1990);
or U1238 (N_1238,In_642,In_1888);
nand U1239 (N_1239,In_197,In_1993);
nor U1240 (N_1240,In_1995,In_1657);
xor U1241 (N_1241,In_454,In_1586);
and U1242 (N_1242,In_1475,In_1494);
or U1243 (N_1243,In_149,In_461);
and U1244 (N_1244,In_75,In_1805);
or U1245 (N_1245,In_1442,In_122);
or U1246 (N_1246,In_947,In_979);
nand U1247 (N_1247,In_1910,In_449);
xor U1248 (N_1248,In_1005,In_1022);
or U1249 (N_1249,In_555,In_1296);
nand U1250 (N_1250,In_1676,In_104);
and U1251 (N_1251,In_1276,In_1084);
nor U1252 (N_1252,In_1524,In_209);
nand U1253 (N_1253,In_1746,In_1465);
or U1254 (N_1254,In_857,In_1146);
and U1255 (N_1255,In_999,In_1881);
nand U1256 (N_1256,In_753,In_999);
or U1257 (N_1257,In_331,In_655);
and U1258 (N_1258,In_579,In_742);
nor U1259 (N_1259,In_1503,In_646);
or U1260 (N_1260,In_714,In_305);
and U1261 (N_1261,In_543,In_481);
and U1262 (N_1262,In_797,In_1261);
nor U1263 (N_1263,In_254,In_1567);
or U1264 (N_1264,In_1585,In_1000);
nor U1265 (N_1265,In_123,In_314);
or U1266 (N_1266,In_1212,In_1725);
or U1267 (N_1267,In_682,In_726);
nor U1268 (N_1268,In_1712,In_244);
nor U1269 (N_1269,In_524,In_676);
xor U1270 (N_1270,In_1543,In_1346);
nand U1271 (N_1271,In_1471,In_813);
and U1272 (N_1272,In_1692,In_497);
and U1273 (N_1273,In_33,In_1394);
or U1274 (N_1274,In_1424,In_1807);
and U1275 (N_1275,In_1218,In_808);
or U1276 (N_1276,In_1826,In_1384);
and U1277 (N_1277,In_1066,In_274);
or U1278 (N_1278,In_1578,In_1659);
and U1279 (N_1279,In_1936,In_1975);
or U1280 (N_1280,In_880,In_545);
nand U1281 (N_1281,In_762,In_1109);
and U1282 (N_1282,In_1888,In_1107);
and U1283 (N_1283,In_1196,In_1102);
nand U1284 (N_1284,In_996,In_1604);
nand U1285 (N_1285,In_1350,In_1829);
and U1286 (N_1286,In_409,In_1326);
and U1287 (N_1287,In_1180,In_530);
nand U1288 (N_1288,In_431,In_1338);
and U1289 (N_1289,In_651,In_1265);
xnor U1290 (N_1290,In_789,In_1599);
or U1291 (N_1291,In_809,In_800);
nand U1292 (N_1292,In_728,In_872);
nor U1293 (N_1293,In_1128,In_761);
and U1294 (N_1294,In_106,In_418);
and U1295 (N_1295,In_303,In_1885);
nor U1296 (N_1296,In_381,In_255);
or U1297 (N_1297,In_1073,In_1143);
and U1298 (N_1298,In_1044,In_123);
or U1299 (N_1299,In_1056,In_769);
xor U1300 (N_1300,In_1779,In_1322);
and U1301 (N_1301,In_437,In_1659);
nand U1302 (N_1302,In_412,In_318);
xor U1303 (N_1303,In_1925,In_683);
and U1304 (N_1304,In_1842,In_1025);
xnor U1305 (N_1305,In_1871,In_67);
nand U1306 (N_1306,In_527,In_851);
and U1307 (N_1307,In_1871,In_902);
and U1308 (N_1308,In_113,In_1957);
xnor U1309 (N_1309,In_579,In_567);
and U1310 (N_1310,In_1964,In_1238);
xnor U1311 (N_1311,In_617,In_165);
and U1312 (N_1312,In_968,In_415);
and U1313 (N_1313,In_1713,In_1334);
or U1314 (N_1314,In_1889,In_408);
or U1315 (N_1315,In_474,In_1564);
nor U1316 (N_1316,In_1296,In_1593);
and U1317 (N_1317,In_1812,In_836);
nor U1318 (N_1318,In_1176,In_1040);
or U1319 (N_1319,In_1768,In_1284);
or U1320 (N_1320,In_1863,In_846);
nor U1321 (N_1321,In_1805,In_1358);
xor U1322 (N_1322,In_525,In_1148);
nand U1323 (N_1323,In_1807,In_118);
nand U1324 (N_1324,In_325,In_393);
nor U1325 (N_1325,In_1390,In_801);
xnor U1326 (N_1326,In_1383,In_1547);
xor U1327 (N_1327,In_1034,In_1325);
and U1328 (N_1328,In_69,In_634);
xnor U1329 (N_1329,In_1699,In_1929);
or U1330 (N_1330,In_597,In_1533);
xor U1331 (N_1331,In_1105,In_1661);
or U1332 (N_1332,In_1920,In_1413);
or U1333 (N_1333,In_1588,In_458);
and U1334 (N_1334,In_1648,In_1782);
xor U1335 (N_1335,In_397,In_406);
or U1336 (N_1336,In_701,In_1490);
or U1337 (N_1337,In_924,In_1050);
or U1338 (N_1338,In_1768,In_1235);
xnor U1339 (N_1339,In_208,In_1039);
and U1340 (N_1340,In_89,In_1075);
and U1341 (N_1341,In_529,In_99);
xor U1342 (N_1342,In_864,In_1459);
or U1343 (N_1343,In_1766,In_1382);
or U1344 (N_1344,In_562,In_1682);
nor U1345 (N_1345,In_850,In_1198);
and U1346 (N_1346,In_1178,In_1814);
nor U1347 (N_1347,In_359,In_6);
nor U1348 (N_1348,In_936,In_1958);
or U1349 (N_1349,In_255,In_395);
and U1350 (N_1350,In_1242,In_1240);
nor U1351 (N_1351,In_864,In_995);
and U1352 (N_1352,In_1939,In_1344);
nand U1353 (N_1353,In_1630,In_1653);
and U1354 (N_1354,In_1956,In_567);
nor U1355 (N_1355,In_996,In_629);
and U1356 (N_1356,In_91,In_1614);
or U1357 (N_1357,In_830,In_75);
and U1358 (N_1358,In_1493,In_1065);
xor U1359 (N_1359,In_878,In_243);
nand U1360 (N_1360,In_1726,In_1866);
nor U1361 (N_1361,In_1985,In_1520);
and U1362 (N_1362,In_597,In_1658);
nor U1363 (N_1363,In_330,In_970);
and U1364 (N_1364,In_833,In_72);
nand U1365 (N_1365,In_701,In_246);
xnor U1366 (N_1366,In_43,In_767);
and U1367 (N_1367,In_91,In_1156);
or U1368 (N_1368,In_733,In_121);
xnor U1369 (N_1369,In_1864,In_619);
nand U1370 (N_1370,In_753,In_1063);
or U1371 (N_1371,In_429,In_1952);
nand U1372 (N_1372,In_1624,In_1466);
and U1373 (N_1373,In_1867,In_1265);
and U1374 (N_1374,In_1147,In_515);
or U1375 (N_1375,In_150,In_785);
nand U1376 (N_1376,In_140,In_856);
or U1377 (N_1377,In_1860,In_1007);
xnor U1378 (N_1378,In_1732,In_1612);
and U1379 (N_1379,In_1515,In_1309);
and U1380 (N_1380,In_919,In_1135);
nor U1381 (N_1381,In_1525,In_1117);
nand U1382 (N_1382,In_923,In_220);
and U1383 (N_1383,In_452,In_1910);
and U1384 (N_1384,In_472,In_447);
nor U1385 (N_1385,In_879,In_7);
and U1386 (N_1386,In_1540,In_1841);
xor U1387 (N_1387,In_842,In_1592);
xor U1388 (N_1388,In_1250,In_1707);
xnor U1389 (N_1389,In_1973,In_835);
and U1390 (N_1390,In_1821,In_1685);
nand U1391 (N_1391,In_1346,In_347);
and U1392 (N_1392,In_644,In_1354);
nor U1393 (N_1393,In_1731,In_1392);
and U1394 (N_1394,In_1910,In_1755);
and U1395 (N_1395,In_403,In_1519);
and U1396 (N_1396,In_1606,In_380);
nor U1397 (N_1397,In_1443,In_1691);
nor U1398 (N_1398,In_860,In_1915);
nand U1399 (N_1399,In_1463,In_417);
and U1400 (N_1400,In_1707,In_1813);
and U1401 (N_1401,In_5,In_1731);
nand U1402 (N_1402,In_1096,In_1423);
nor U1403 (N_1403,In_304,In_1984);
or U1404 (N_1404,In_307,In_1212);
nand U1405 (N_1405,In_1785,In_740);
or U1406 (N_1406,In_386,In_1591);
or U1407 (N_1407,In_1797,In_1605);
and U1408 (N_1408,In_142,In_1353);
nor U1409 (N_1409,In_1105,In_1727);
xor U1410 (N_1410,In_122,In_1895);
nor U1411 (N_1411,In_706,In_1187);
nand U1412 (N_1412,In_1742,In_1857);
and U1413 (N_1413,In_1969,In_1690);
nor U1414 (N_1414,In_869,In_1564);
or U1415 (N_1415,In_176,In_746);
xor U1416 (N_1416,In_1200,In_921);
xnor U1417 (N_1417,In_1985,In_1428);
or U1418 (N_1418,In_975,In_1193);
nor U1419 (N_1419,In_713,In_881);
nor U1420 (N_1420,In_1691,In_412);
or U1421 (N_1421,In_1173,In_508);
or U1422 (N_1422,In_1938,In_1717);
and U1423 (N_1423,In_816,In_875);
nor U1424 (N_1424,In_1428,In_68);
or U1425 (N_1425,In_710,In_1534);
xnor U1426 (N_1426,In_1993,In_548);
nor U1427 (N_1427,In_728,In_1604);
or U1428 (N_1428,In_1117,In_90);
xnor U1429 (N_1429,In_988,In_1660);
nor U1430 (N_1430,In_1433,In_1643);
nor U1431 (N_1431,In_1973,In_822);
or U1432 (N_1432,In_948,In_1760);
nand U1433 (N_1433,In_650,In_1191);
nor U1434 (N_1434,In_1719,In_545);
nor U1435 (N_1435,In_1754,In_1361);
and U1436 (N_1436,In_655,In_1896);
xor U1437 (N_1437,In_1146,In_1897);
nand U1438 (N_1438,In_156,In_1880);
or U1439 (N_1439,In_674,In_315);
nand U1440 (N_1440,In_265,In_566);
nor U1441 (N_1441,In_627,In_1150);
nand U1442 (N_1442,In_248,In_1416);
and U1443 (N_1443,In_1734,In_155);
nand U1444 (N_1444,In_189,In_1921);
xor U1445 (N_1445,In_66,In_1343);
xnor U1446 (N_1446,In_134,In_858);
nor U1447 (N_1447,In_840,In_584);
nor U1448 (N_1448,In_739,In_92);
xnor U1449 (N_1449,In_625,In_876);
nand U1450 (N_1450,In_960,In_990);
xnor U1451 (N_1451,In_272,In_693);
nand U1452 (N_1452,In_1016,In_275);
nor U1453 (N_1453,In_147,In_1121);
xor U1454 (N_1454,In_906,In_1606);
xnor U1455 (N_1455,In_1111,In_1786);
xor U1456 (N_1456,In_1926,In_316);
and U1457 (N_1457,In_996,In_1214);
or U1458 (N_1458,In_256,In_1697);
or U1459 (N_1459,In_1738,In_234);
or U1460 (N_1460,In_926,In_1899);
or U1461 (N_1461,In_896,In_1775);
nand U1462 (N_1462,In_810,In_990);
or U1463 (N_1463,In_13,In_694);
nor U1464 (N_1464,In_945,In_791);
nand U1465 (N_1465,In_994,In_1355);
or U1466 (N_1466,In_1076,In_1834);
nand U1467 (N_1467,In_455,In_733);
and U1468 (N_1468,In_1064,In_66);
xor U1469 (N_1469,In_1599,In_1310);
nor U1470 (N_1470,In_1091,In_703);
xnor U1471 (N_1471,In_761,In_721);
or U1472 (N_1472,In_599,In_1980);
nor U1473 (N_1473,In_210,In_138);
xor U1474 (N_1474,In_161,In_746);
xor U1475 (N_1475,In_829,In_1035);
and U1476 (N_1476,In_1374,In_1531);
or U1477 (N_1477,In_351,In_1610);
nand U1478 (N_1478,In_1166,In_605);
and U1479 (N_1479,In_735,In_387);
or U1480 (N_1480,In_36,In_1932);
xor U1481 (N_1481,In_685,In_126);
or U1482 (N_1482,In_115,In_877);
nor U1483 (N_1483,In_161,In_1472);
nand U1484 (N_1484,In_1456,In_50);
or U1485 (N_1485,In_370,In_315);
nor U1486 (N_1486,In_845,In_1994);
or U1487 (N_1487,In_1056,In_1287);
or U1488 (N_1488,In_377,In_1643);
nand U1489 (N_1489,In_144,In_1957);
and U1490 (N_1490,In_1516,In_1599);
or U1491 (N_1491,In_1427,In_802);
xnor U1492 (N_1492,In_645,In_1336);
xnor U1493 (N_1493,In_1107,In_665);
or U1494 (N_1494,In_1252,In_1014);
and U1495 (N_1495,In_1770,In_605);
xnor U1496 (N_1496,In_467,In_1543);
or U1497 (N_1497,In_1511,In_519);
nor U1498 (N_1498,In_175,In_340);
xor U1499 (N_1499,In_935,In_1926);
xnor U1500 (N_1500,In_1669,In_1923);
nor U1501 (N_1501,In_1060,In_128);
xnor U1502 (N_1502,In_1190,In_1166);
nand U1503 (N_1503,In_734,In_837);
nor U1504 (N_1504,In_341,In_1463);
and U1505 (N_1505,In_1675,In_1942);
xnor U1506 (N_1506,In_1706,In_363);
and U1507 (N_1507,In_1016,In_1628);
nor U1508 (N_1508,In_668,In_288);
or U1509 (N_1509,In_78,In_725);
and U1510 (N_1510,In_1928,In_1914);
nor U1511 (N_1511,In_655,In_332);
xnor U1512 (N_1512,In_316,In_1068);
xor U1513 (N_1513,In_155,In_1651);
nand U1514 (N_1514,In_567,In_1445);
xnor U1515 (N_1515,In_1841,In_1837);
xor U1516 (N_1516,In_1798,In_1614);
xor U1517 (N_1517,In_1451,In_143);
and U1518 (N_1518,In_1831,In_810);
nand U1519 (N_1519,In_102,In_299);
xnor U1520 (N_1520,In_1882,In_380);
and U1521 (N_1521,In_982,In_1806);
or U1522 (N_1522,In_633,In_1039);
xnor U1523 (N_1523,In_578,In_1338);
xnor U1524 (N_1524,In_133,In_651);
and U1525 (N_1525,In_367,In_95);
nor U1526 (N_1526,In_1534,In_115);
nor U1527 (N_1527,In_1274,In_1080);
and U1528 (N_1528,In_116,In_301);
xnor U1529 (N_1529,In_156,In_474);
and U1530 (N_1530,In_80,In_584);
nand U1531 (N_1531,In_1749,In_1069);
nand U1532 (N_1532,In_155,In_157);
nor U1533 (N_1533,In_966,In_1050);
xor U1534 (N_1534,In_1673,In_688);
xor U1535 (N_1535,In_181,In_1485);
nor U1536 (N_1536,In_319,In_287);
xnor U1537 (N_1537,In_1223,In_1977);
or U1538 (N_1538,In_1548,In_1865);
and U1539 (N_1539,In_116,In_1500);
and U1540 (N_1540,In_175,In_1534);
and U1541 (N_1541,In_1195,In_788);
xor U1542 (N_1542,In_1105,In_1576);
or U1543 (N_1543,In_1771,In_1714);
nor U1544 (N_1544,In_1139,In_1348);
nor U1545 (N_1545,In_1647,In_1639);
nand U1546 (N_1546,In_1540,In_1903);
or U1547 (N_1547,In_1618,In_1175);
or U1548 (N_1548,In_605,In_154);
xnor U1549 (N_1549,In_808,In_823);
nor U1550 (N_1550,In_1199,In_1419);
xor U1551 (N_1551,In_549,In_499);
xor U1552 (N_1552,In_862,In_1014);
or U1553 (N_1553,In_1384,In_1709);
nand U1554 (N_1554,In_1370,In_1757);
or U1555 (N_1555,In_1,In_1136);
nand U1556 (N_1556,In_822,In_1795);
or U1557 (N_1557,In_1447,In_11);
or U1558 (N_1558,In_1438,In_1188);
xor U1559 (N_1559,In_1210,In_1645);
nor U1560 (N_1560,In_653,In_1827);
and U1561 (N_1561,In_84,In_265);
and U1562 (N_1562,In_877,In_1582);
nand U1563 (N_1563,In_1375,In_1755);
and U1564 (N_1564,In_520,In_1026);
nand U1565 (N_1565,In_1978,In_1164);
nor U1566 (N_1566,In_729,In_1490);
nand U1567 (N_1567,In_1793,In_856);
and U1568 (N_1568,In_612,In_1237);
nand U1569 (N_1569,In_1626,In_1667);
nand U1570 (N_1570,In_1214,In_1158);
or U1571 (N_1571,In_872,In_502);
nand U1572 (N_1572,In_922,In_756);
nor U1573 (N_1573,In_556,In_1832);
xnor U1574 (N_1574,In_1978,In_1089);
nand U1575 (N_1575,In_929,In_1058);
and U1576 (N_1576,In_549,In_1229);
nor U1577 (N_1577,In_40,In_371);
nor U1578 (N_1578,In_90,In_667);
or U1579 (N_1579,In_760,In_1709);
nand U1580 (N_1580,In_1873,In_1100);
nand U1581 (N_1581,In_1541,In_1743);
and U1582 (N_1582,In_1285,In_1617);
xor U1583 (N_1583,In_444,In_346);
nand U1584 (N_1584,In_1564,In_295);
nand U1585 (N_1585,In_1582,In_14);
nor U1586 (N_1586,In_1166,In_1195);
and U1587 (N_1587,In_569,In_426);
and U1588 (N_1588,In_1900,In_927);
nor U1589 (N_1589,In_65,In_1855);
nor U1590 (N_1590,In_1941,In_771);
nand U1591 (N_1591,In_1557,In_1023);
or U1592 (N_1592,In_1842,In_1329);
and U1593 (N_1593,In_1449,In_1937);
or U1594 (N_1594,In_1752,In_1501);
xor U1595 (N_1595,In_168,In_1456);
or U1596 (N_1596,In_1422,In_701);
and U1597 (N_1597,In_454,In_13);
xor U1598 (N_1598,In_1068,In_796);
or U1599 (N_1599,In_162,In_1960);
and U1600 (N_1600,In_1186,In_107);
nor U1601 (N_1601,In_1433,In_1);
nand U1602 (N_1602,In_1302,In_845);
and U1603 (N_1603,In_778,In_398);
nor U1604 (N_1604,In_1889,In_933);
xnor U1605 (N_1605,In_653,In_679);
nand U1606 (N_1606,In_1744,In_1850);
nor U1607 (N_1607,In_507,In_1884);
or U1608 (N_1608,In_1534,In_420);
nand U1609 (N_1609,In_72,In_1025);
xnor U1610 (N_1610,In_1251,In_758);
nor U1611 (N_1611,In_615,In_916);
or U1612 (N_1612,In_221,In_1897);
xor U1613 (N_1613,In_915,In_320);
and U1614 (N_1614,In_1233,In_36);
nand U1615 (N_1615,In_104,In_1971);
and U1616 (N_1616,In_1223,In_1940);
or U1617 (N_1617,In_332,In_1582);
nand U1618 (N_1618,In_62,In_1769);
nor U1619 (N_1619,In_414,In_695);
or U1620 (N_1620,In_1967,In_684);
nor U1621 (N_1621,In_1532,In_382);
and U1622 (N_1622,In_1585,In_1620);
and U1623 (N_1623,In_1195,In_1606);
xor U1624 (N_1624,In_1897,In_95);
xor U1625 (N_1625,In_869,In_296);
nor U1626 (N_1626,In_582,In_1887);
and U1627 (N_1627,In_1139,In_1871);
or U1628 (N_1628,In_1233,In_396);
and U1629 (N_1629,In_1827,In_1526);
xor U1630 (N_1630,In_1553,In_694);
xor U1631 (N_1631,In_1060,In_1569);
or U1632 (N_1632,In_1728,In_1622);
or U1633 (N_1633,In_953,In_1716);
or U1634 (N_1634,In_927,In_1401);
nand U1635 (N_1635,In_599,In_212);
or U1636 (N_1636,In_698,In_220);
nand U1637 (N_1637,In_624,In_1560);
nand U1638 (N_1638,In_1365,In_1643);
nand U1639 (N_1639,In_148,In_582);
nand U1640 (N_1640,In_1337,In_160);
nand U1641 (N_1641,In_842,In_380);
nor U1642 (N_1642,In_717,In_1187);
or U1643 (N_1643,In_840,In_462);
and U1644 (N_1644,In_1979,In_407);
nor U1645 (N_1645,In_1333,In_1794);
or U1646 (N_1646,In_1439,In_874);
or U1647 (N_1647,In_724,In_1544);
xnor U1648 (N_1648,In_1963,In_60);
nand U1649 (N_1649,In_1261,In_668);
xor U1650 (N_1650,In_1001,In_536);
or U1651 (N_1651,In_221,In_865);
or U1652 (N_1652,In_723,In_1046);
nor U1653 (N_1653,In_244,In_951);
xor U1654 (N_1654,In_1597,In_1157);
nor U1655 (N_1655,In_398,In_1991);
or U1656 (N_1656,In_1758,In_1924);
nand U1657 (N_1657,In_964,In_744);
nand U1658 (N_1658,In_184,In_584);
nor U1659 (N_1659,In_1241,In_1064);
nand U1660 (N_1660,In_1611,In_1003);
or U1661 (N_1661,In_489,In_1092);
nor U1662 (N_1662,In_719,In_1341);
nand U1663 (N_1663,In_168,In_703);
xor U1664 (N_1664,In_271,In_1869);
nand U1665 (N_1665,In_147,In_259);
nand U1666 (N_1666,In_1878,In_129);
xnor U1667 (N_1667,In_1174,In_253);
or U1668 (N_1668,In_60,In_267);
and U1669 (N_1669,In_361,In_1688);
nand U1670 (N_1670,In_1854,In_90);
xnor U1671 (N_1671,In_1695,In_1807);
or U1672 (N_1672,In_1255,In_307);
and U1673 (N_1673,In_802,In_933);
xnor U1674 (N_1674,In_102,In_1197);
and U1675 (N_1675,In_582,In_1807);
nor U1676 (N_1676,In_82,In_1133);
or U1677 (N_1677,In_1323,In_15);
and U1678 (N_1678,In_1803,In_1500);
and U1679 (N_1679,In_681,In_1648);
and U1680 (N_1680,In_559,In_639);
nor U1681 (N_1681,In_48,In_1466);
nor U1682 (N_1682,In_695,In_1597);
or U1683 (N_1683,In_152,In_1401);
xnor U1684 (N_1684,In_1214,In_947);
and U1685 (N_1685,In_525,In_372);
or U1686 (N_1686,In_1187,In_147);
and U1687 (N_1687,In_878,In_1208);
and U1688 (N_1688,In_1307,In_1722);
and U1689 (N_1689,In_929,In_1403);
xnor U1690 (N_1690,In_370,In_387);
and U1691 (N_1691,In_1437,In_458);
nor U1692 (N_1692,In_830,In_1220);
nand U1693 (N_1693,In_970,In_1500);
xor U1694 (N_1694,In_563,In_547);
nand U1695 (N_1695,In_1885,In_760);
nand U1696 (N_1696,In_1341,In_491);
and U1697 (N_1697,In_666,In_1144);
and U1698 (N_1698,In_1818,In_860);
and U1699 (N_1699,In_1361,In_744);
and U1700 (N_1700,In_1984,In_782);
nor U1701 (N_1701,In_116,In_1828);
nand U1702 (N_1702,In_656,In_464);
or U1703 (N_1703,In_1934,In_1205);
xnor U1704 (N_1704,In_264,In_651);
nand U1705 (N_1705,In_1831,In_737);
or U1706 (N_1706,In_1847,In_1472);
and U1707 (N_1707,In_1059,In_910);
or U1708 (N_1708,In_996,In_294);
and U1709 (N_1709,In_925,In_1964);
xnor U1710 (N_1710,In_793,In_458);
xor U1711 (N_1711,In_653,In_1864);
xor U1712 (N_1712,In_852,In_1367);
and U1713 (N_1713,In_56,In_1974);
or U1714 (N_1714,In_742,In_1690);
or U1715 (N_1715,In_340,In_826);
or U1716 (N_1716,In_138,In_1225);
nor U1717 (N_1717,In_1056,In_113);
or U1718 (N_1718,In_1769,In_1424);
or U1719 (N_1719,In_1606,In_1106);
and U1720 (N_1720,In_1518,In_978);
and U1721 (N_1721,In_706,In_1047);
and U1722 (N_1722,In_1527,In_834);
or U1723 (N_1723,In_1782,In_1207);
nor U1724 (N_1724,In_571,In_26);
nor U1725 (N_1725,In_136,In_1733);
nor U1726 (N_1726,In_1821,In_1727);
or U1727 (N_1727,In_213,In_1870);
or U1728 (N_1728,In_1230,In_1949);
or U1729 (N_1729,In_1796,In_584);
nor U1730 (N_1730,In_1188,In_1644);
nor U1731 (N_1731,In_496,In_808);
xor U1732 (N_1732,In_1054,In_1193);
nand U1733 (N_1733,In_127,In_384);
or U1734 (N_1734,In_104,In_1472);
or U1735 (N_1735,In_680,In_1154);
nand U1736 (N_1736,In_647,In_481);
and U1737 (N_1737,In_707,In_1243);
xor U1738 (N_1738,In_283,In_1108);
nor U1739 (N_1739,In_1447,In_206);
and U1740 (N_1740,In_1686,In_1613);
or U1741 (N_1741,In_1080,In_639);
nor U1742 (N_1742,In_233,In_996);
nor U1743 (N_1743,In_62,In_1359);
nand U1744 (N_1744,In_1996,In_890);
nor U1745 (N_1745,In_694,In_1371);
nor U1746 (N_1746,In_1554,In_437);
nand U1747 (N_1747,In_448,In_84);
and U1748 (N_1748,In_853,In_544);
and U1749 (N_1749,In_1779,In_383);
nand U1750 (N_1750,In_903,In_363);
xnor U1751 (N_1751,In_1209,In_1734);
nand U1752 (N_1752,In_688,In_1839);
nor U1753 (N_1753,In_1143,In_1706);
xnor U1754 (N_1754,In_642,In_206);
or U1755 (N_1755,In_165,In_643);
nand U1756 (N_1756,In_1241,In_1152);
and U1757 (N_1757,In_1443,In_178);
nand U1758 (N_1758,In_1379,In_1403);
nor U1759 (N_1759,In_633,In_1217);
or U1760 (N_1760,In_948,In_744);
or U1761 (N_1761,In_426,In_965);
nand U1762 (N_1762,In_757,In_1689);
or U1763 (N_1763,In_1603,In_746);
and U1764 (N_1764,In_651,In_1113);
and U1765 (N_1765,In_1685,In_1813);
nor U1766 (N_1766,In_1315,In_1894);
and U1767 (N_1767,In_1738,In_401);
nand U1768 (N_1768,In_217,In_1409);
and U1769 (N_1769,In_302,In_1346);
and U1770 (N_1770,In_1902,In_199);
or U1771 (N_1771,In_1248,In_1400);
nor U1772 (N_1772,In_1629,In_727);
xnor U1773 (N_1773,In_1368,In_563);
and U1774 (N_1774,In_748,In_202);
xnor U1775 (N_1775,In_167,In_1392);
nor U1776 (N_1776,In_1004,In_1994);
or U1777 (N_1777,In_208,In_556);
and U1778 (N_1778,In_1196,In_1628);
or U1779 (N_1779,In_718,In_1181);
and U1780 (N_1780,In_282,In_1171);
nand U1781 (N_1781,In_116,In_1736);
or U1782 (N_1782,In_1847,In_1941);
nor U1783 (N_1783,In_487,In_1006);
or U1784 (N_1784,In_802,In_1702);
and U1785 (N_1785,In_965,In_1780);
or U1786 (N_1786,In_184,In_1712);
nand U1787 (N_1787,In_1283,In_681);
xnor U1788 (N_1788,In_1782,In_972);
nor U1789 (N_1789,In_936,In_1160);
or U1790 (N_1790,In_207,In_683);
nor U1791 (N_1791,In_1413,In_385);
nor U1792 (N_1792,In_599,In_278);
and U1793 (N_1793,In_33,In_405);
or U1794 (N_1794,In_1921,In_1136);
nor U1795 (N_1795,In_771,In_939);
xor U1796 (N_1796,In_1140,In_766);
or U1797 (N_1797,In_1583,In_1569);
and U1798 (N_1798,In_101,In_353);
or U1799 (N_1799,In_403,In_1953);
or U1800 (N_1800,In_708,In_1109);
and U1801 (N_1801,In_1455,In_1878);
xor U1802 (N_1802,In_938,In_631);
or U1803 (N_1803,In_661,In_27);
nand U1804 (N_1804,In_322,In_1038);
or U1805 (N_1805,In_966,In_401);
xnor U1806 (N_1806,In_804,In_819);
nand U1807 (N_1807,In_833,In_499);
or U1808 (N_1808,In_1103,In_1437);
or U1809 (N_1809,In_1177,In_1711);
or U1810 (N_1810,In_1493,In_1023);
or U1811 (N_1811,In_842,In_1473);
xor U1812 (N_1812,In_1971,In_1094);
and U1813 (N_1813,In_1934,In_611);
nor U1814 (N_1814,In_462,In_1887);
nand U1815 (N_1815,In_1917,In_1885);
xnor U1816 (N_1816,In_1430,In_1738);
and U1817 (N_1817,In_435,In_1056);
nand U1818 (N_1818,In_1853,In_596);
nand U1819 (N_1819,In_832,In_1830);
nor U1820 (N_1820,In_776,In_1007);
and U1821 (N_1821,In_594,In_593);
nand U1822 (N_1822,In_1868,In_1461);
xnor U1823 (N_1823,In_1660,In_204);
or U1824 (N_1824,In_852,In_1826);
or U1825 (N_1825,In_264,In_518);
nor U1826 (N_1826,In_273,In_1457);
and U1827 (N_1827,In_630,In_1139);
xnor U1828 (N_1828,In_1061,In_295);
nor U1829 (N_1829,In_1784,In_1658);
xnor U1830 (N_1830,In_1757,In_401);
or U1831 (N_1831,In_1964,In_1570);
nor U1832 (N_1832,In_70,In_1456);
nor U1833 (N_1833,In_749,In_1985);
nor U1834 (N_1834,In_1629,In_1121);
xnor U1835 (N_1835,In_1277,In_729);
xnor U1836 (N_1836,In_440,In_1908);
or U1837 (N_1837,In_1142,In_1425);
nor U1838 (N_1838,In_712,In_1577);
and U1839 (N_1839,In_1271,In_789);
nand U1840 (N_1840,In_1197,In_1281);
or U1841 (N_1841,In_687,In_1530);
xnor U1842 (N_1842,In_809,In_518);
and U1843 (N_1843,In_1275,In_441);
nand U1844 (N_1844,In_1014,In_700);
xnor U1845 (N_1845,In_1452,In_1007);
xor U1846 (N_1846,In_1483,In_561);
xor U1847 (N_1847,In_836,In_1137);
nor U1848 (N_1848,In_888,In_1504);
nor U1849 (N_1849,In_216,In_1142);
xor U1850 (N_1850,In_860,In_112);
and U1851 (N_1851,In_111,In_1546);
nand U1852 (N_1852,In_1888,In_234);
nor U1853 (N_1853,In_405,In_1097);
or U1854 (N_1854,In_1790,In_1455);
nand U1855 (N_1855,In_1155,In_876);
or U1856 (N_1856,In_1463,In_257);
and U1857 (N_1857,In_1671,In_1105);
and U1858 (N_1858,In_1438,In_1698);
and U1859 (N_1859,In_912,In_1934);
nor U1860 (N_1860,In_1496,In_354);
and U1861 (N_1861,In_1051,In_862);
nor U1862 (N_1862,In_418,In_27);
nand U1863 (N_1863,In_635,In_95);
nand U1864 (N_1864,In_1595,In_896);
xor U1865 (N_1865,In_1853,In_1167);
and U1866 (N_1866,In_353,In_52);
nor U1867 (N_1867,In_1246,In_1520);
or U1868 (N_1868,In_1516,In_1785);
nand U1869 (N_1869,In_1616,In_644);
or U1870 (N_1870,In_1654,In_1301);
nand U1871 (N_1871,In_544,In_1951);
or U1872 (N_1872,In_1271,In_1623);
or U1873 (N_1873,In_1416,In_1591);
or U1874 (N_1874,In_1418,In_1291);
or U1875 (N_1875,In_711,In_19);
nor U1876 (N_1876,In_1184,In_459);
xnor U1877 (N_1877,In_358,In_633);
xnor U1878 (N_1878,In_407,In_49);
nand U1879 (N_1879,In_1011,In_8);
or U1880 (N_1880,In_888,In_285);
or U1881 (N_1881,In_5,In_1);
nor U1882 (N_1882,In_1434,In_1832);
nor U1883 (N_1883,In_1610,In_313);
nor U1884 (N_1884,In_392,In_785);
xor U1885 (N_1885,In_1069,In_804);
or U1886 (N_1886,In_1376,In_1109);
nor U1887 (N_1887,In_100,In_10);
or U1888 (N_1888,In_1080,In_120);
and U1889 (N_1889,In_818,In_460);
nor U1890 (N_1890,In_1678,In_1077);
or U1891 (N_1891,In_338,In_636);
or U1892 (N_1892,In_1035,In_1930);
xnor U1893 (N_1893,In_44,In_673);
xnor U1894 (N_1894,In_96,In_160);
and U1895 (N_1895,In_1512,In_455);
nor U1896 (N_1896,In_1935,In_1671);
or U1897 (N_1897,In_1101,In_1558);
nand U1898 (N_1898,In_1695,In_508);
and U1899 (N_1899,In_1996,In_269);
nor U1900 (N_1900,In_233,In_1205);
or U1901 (N_1901,In_1115,In_1196);
nand U1902 (N_1902,In_435,In_706);
or U1903 (N_1903,In_1131,In_1446);
and U1904 (N_1904,In_1082,In_1647);
nor U1905 (N_1905,In_1423,In_1949);
xor U1906 (N_1906,In_116,In_1430);
nand U1907 (N_1907,In_54,In_1947);
and U1908 (N_1908,In_392,In_1936);
xor U1909 (N_1909,In_698,In_695);
xor U1910 (N_1910,In_1440,In_1348);
nor U1911 (N_1911,In_1202,In_1637);
and U1912 (N_1912,In_1354,In_1188);
or U1913 (N_1913,In_1056,In_1756);
nand U1914 (N_1914,In_716,In_1457);
nand U1915 (N_1915,In_773,In_1222);
or U1916 (N_1916,In_1226,In_970);
nor U1917 (N_1917,In_1266,In_809);
or U1918 (N_1918,In_1515,In_751);
or U1919 (N_1919,In_246,In_61);
nor U1920 (N_1920,In_443,In_1376);
or U1921 (N_1921,In_1260,In_555);
nand U1922 (N_1922,In_156,In_1644);
nor U1923 (N_1923,In_1890,In_107);
nor U1924 (N_1924,In_1145,In_26);
nand U1925 (N_1925,In_1594,In_1660);
nor U1926 (N_1926,In_775,In_1587);
and U1927 (N_1927,In_121,In_1840);
or U1928 (N_1928,In_1109,In_111);
nor U1929 (N_1929,In_1919,In_1564);
nor U1930 (N_1930,In_113,In_1510);
nand U1931 (N_1931,In_1831,In_1258);
or U1932 (N_1932,In_1537,In_536);
nor U1933 (N_1933,In_1520,In_1472);
nor U1934 (N_1934,In_1879,In_942);
and U1935 (N_1935,In_942,In_1404);
xnor U1936 (N_1936,In_1464,In_1859);
nor U1937 (N_1937,In_1471,In_418);
nand U1938 (N_1938,In_214,In_1431);
and U1939 (N_1939,In_346,In_1658);
xnor U1940 (N_1940,In_306,In_1725);
nand U1941 (N_1941,In_801,In_951);
and U1942 (N_1942,In_1858,In_1876);
or U1943 (N_1943,In_1434,In_1287);
nor U1944 (N_1944,In_687,In_1438);
xor U1945 (N_1945,In_1252,In_1750);
xor U1946 (N_1946,In_203,In_1577);
nand U1947 (N_1947,In_846,In_471);
and U1948 (N_1948,In_391,In_1297);
nand U1949 (N_1949,In_73,In_1802);
nand U1950 (N_1950,In_205,In_1090);
and U1951 (N_1951,In_1114,In_1785);
or U1952 (N_1952,In_744,In_488);
xor U1953 (N_1953,In_1037,In_754);
nand U1954 (N_1954,In_1269,In_602);
nand U1955 (N_1955,In_1940,In_253);
nand U1956 (N_1956,In_659,In_475);
nand U1957 (N_1957,In_1954,In_1000);
or U1958 (N_1958,In_953,In_768);
or U1959 (N_1959,In_1441,In_1117);
xor U1960 (N_1960,In_1976,In_1772);
nand U1961 (N_1961,In_1779,In_1991);
nor U1962 (N_1962,In_1268,In_458);
nand U1963 (N_1963,In_1171,In_1380);
or U1964 (N_1964,In_1451,In_525);
nand U1965 (N_1965,In_379,In_97);
nand U1966 (N_1966,In_882,In_245);
and U1967 (N_1967,In_665,In_439);
nor U1968 (N_1968,In_262,In_1069);
nor U1969 (N_1969,In_740,In_416);
nor U1970 (N_1970,In_1017,In_165);
and U1971 (N_1971,In_927,In_555);
xor U1972 (N_1972,In_907,In_1000);
or U1973 (N_1973,In_132,In_514);
and U1974 (N_1974,In_421,In_516);
and U1975 (N_1975,In_1257,In_962);
or U1976 (N_1976,In_1213,In_1470);
and U1977 (N_1977,In_241,In_709);
and U1978 (N_1978,In_1857,In_718);
or U1979 (N_1979,In_274,In_1146);
nor U1980 (N_1980,In_884,In_31);
nand U1981 (N_1981,In_1778,In_989);
xnor U1982 (N_1982,In_988,In_914);
nand U1983 (N_1983,In_1416,In_1344);
or U1984 (N_1984,In_201,In_347);
and U1985 (N_1985,In_1252,In_1022);
nor U1986 (N_1986,In_1643,In_1649);
or U1987 (N_1987,In_23,In_817);
and U1988 (N_1988,In_522,In_937);
nand U1989 (N_1989,In_1358,In_779);
and U1990 (N_1990,In_1918,In_432);
and U1991 (N_1991,In_1402,In_507);
nor U1992 (N_1992,In_1570,In_1621);
xor U1993 (N_1993,In_611,In_1941);
nor U1994 (N_1994,In_1908,In_165);
xnor U1995 (N_1995,In_761,In_1118);
or U1996 (N_1996,In_311,In_1822);
and U1997 (N_1997,In_1529,In_183);
nor U1998 (N_1998,In_1235,In_790);
xnor U1999 (N_1999,In_1595,In_1542);
xor U2000 (N_2000,In_1301,In_1287);
nor U2001 (N_2001,In_1926,In_1179);
and U2002 (N_2002,In_1454,In_189);
nand U2003 (N_2003,In_1230,In_966);
or U2004 (N_2004,In_828,In_1986);
and U2005 (N_2005,In_671,In_250);
and U2006 (N_2006,In_269,In_220);
nand U2007 (N_2007,In_265,In_1590);
nor U2008 (N_2008,In_1082,In_1686);
and U2009 (N_2009,In_1819,In_789);
nand U2010 (N_2010,In_1761,In_1930);
nor U2011 (N_2011,In_1237,In_1793);
and U2012 (N_2012,In_983,In_1657);
nor U2013 (N_2013,In_41,In_1368);
and U2014 (N_2014,In_103,In_1290);
nor U2015 (N_2015,In_230,In_1976);
nor U2016 (N_2016,In_1215,In_1087);
and U2017 (N_2017,In_1670,In_807);
nor U2018 (N_2018,In_130,In_1294);
nor U2019 (N_2019,In_77,In_1060);
xnor U2020 (N_2020,In_1993,In_1523);
nand U2021 (N_2021,In_1291,In_186);
nand U2022 (N_2022,In_1461,In_560);
and U2023 (N_2023,In_1482,In_908);
nand U2024 (N_2024,In_980,In_611);
nand U2025 (N_2025,In_446,In_219);
or U2026 (N_2026,In_1281,In_97);
nor U2027 (N_2027,In_1684,In_258);
or U2028 (N_2028,In_835,In_23);
xor U2029 (N_2029,In_1325,In_282);
xnor U2030 (N_2030,In_1741,In_1759);
and U2031 (N_2031,In_1248,In_1192);
and U2032 (N_2032,In_1227,In_198);
nor U2033 (N_2033,In_633,In_1660);
nor U2034 (N_2034,In_421,In_956);
and U2035 (N_2035,In_716,In_541);
nand U2036 (N_2036,In_1331,In_1019);
and U2037 (N_2037,In_1892,In_586);
nor U2038 (N_2038,In_1749,In_987);
nor U2039 (N_2039,In_1467,In_144);
xnor U2040 (N_2040,In_973,In_1386);
nand U2041 (N_2041,In_1884,In_1414);
or U2042 (N_2042,In_535,In_14);
nor U2043 (N_2043,In_1142,In_629);
or U2044 (N_2044,In_849,In_1852);
nor U2045 (N_2045,In_891,In_227);
nand U2046 (N_2046,In_1138,In_1796);
and U2047 (N_2047,In_1447,In_1736);
nand U2048 (N_2048,In_1494,In_989);
or U2049 (N_2049,In_474,In_133);
and U2050 (N_2050,In_1549,In_1854);
and U2051 (N_2051,In_1204,In_752);
nor U2052 (N_2052,In_1477,In_667);
and U2053 (N_2053,In_610,In_1898);
nand U2054 (N_2054,In_1144,In_238);
or U2055 (N_2055,In_54,In_1703);
and U2056 (N_2056,In_1041,In_116);
and U2057 (N_2057,In_1864,In_348);
nor U2058 (N_2058,In_310,In_1515);
xnor U2059 (N_2059,In_113,In_1190);
or U2060 (N_2060,In_16,In_882);
and U2061 (N_2061,In_671,In_672);
nor U2062 (N_2062,In_1520,In_1824);
or U2063 (N_2063,In_416,In_1272);
nand U2064 (N_2064,In_811,In_86);
nand U2065 (N_2065,In_808,In_425);
nor U2066 (N_2066,In_624,In_657);
xnor U2067 (N_2067,In_1958,In_392);
or U2068 (N_2068,In_1376,In_1950);
xnor U2069 (N_2069,In_572,In_753);
or U2070 (N_2070,In_1035,In_1043);
nor U2071 (N_2071,In_1514,In_193);
and U2072 (N_2072,In_1245,In_893);
nor U2073 (N_2073,In_662,In_1986);
and U2074 (N_2074,In_1918,In_1287);
nand U2075 (N_2075,In_364,In_1695);
nand U2076 (N_2076,In_1098,In_49);
and U2077 (N_2077,In_951,In_1764);
and U2078 (N_2078,In_508,In_587);
xnor U2079 (N_2079,In_1618,In_191);
and U2080 (N_2080,In_1424,In_539);
or U2081 (N_2081,In_1734,In_29);
and U2082 (N_2082,In_711,In_1780);
nand U2083 (N_2083,In_1801,In_910);
nand U2084 (N_2084,In_297,In_1215);
xor U2085 (N_2085,In_680,In_506);
and U2086 (N_2086,In_1584,In_1902);
or U2087 (N_2087,In_1837,In_379);
xor U2088 (N_2088,In_637,In_455);
nor U2089 (N_2089,In_83,In_1558);
nor U2090 (N_2090,In_1658,In_1930);
or U2091 (N_2091,In_1569,In_1755);
or U2092 (N_2092,In_1066,In_1708);
or U2093 (N_2093,In_339,In_1572);
nor U2094 (N_2094,In_1945,In_1802);
xnor U2095 (N_2095,In_214,In_641);
or U2096 (N_2096,In_1371,In_268);
xnor U2097 (N_2097,In_5,In_1474);
nand U2098 (N_2098,In_1832,In_894);
or U2099 (N_2099,In_1335,In_109);
xor U2100 (N_2100,In_1976,In_1834);
or U2101 (N_2101,In_1372,In_100);
and U2102 (N_2102,In_547,In_1402);
or U2103 (N_2103,In_1205,In_143);
or U2104 (N_2104,In_1166,In_882);
and U2105 (N_2105,In_1384,In_1287);
or U2106 (N_2106,In_861,In_1429);
nand U2107 (N_2107,In_249,In_278);
nand U2108 (N_2108,In_51,In_1326);
and U2109 (N_2109,In_1885,In_1941);
and U2110 (N_2110,In_1045,In_238);
and U2111 (N_2111,In_57,In_76);
nand U2112 (N_2112,In_352,In_129);
or U2113 (N_2113,In_507,In_1969);
nand U2114 (N_2114,In_752,In_1113);
or U2115 (N_2115,In_1480,In_429);
nor U2116 (N_2116,In_1644,In_1805);
nand U2117 (N_2117,In_360,In_299);
nor U2118 (N_2118,In_1795,In_570);
xnor U2119 (N_2119,In_298,In_881);
and U2120 (N_2120,In_935,In_247);
nand U2121 (N_2121,In_1451,In_270);
and U2122 (N_2122,In_1813,In_534);
and U2123 (N_2123,In_1768,In_1800);
nand U2124 (N_2124,In_596,In_191);
xnor U2125 (N_2125,In_795,In_1471);
nor U2126 (N_2126,In_1423,In_529);
xnor U2127 (N_2127,In_173,In_685);
nand U2128 (N_2128,In_714,In_807);
or U2129 (N_2129,In_342,In_142);
nand U2130 (N_2130,In_1536,In_655);
and U2131 (N_2131,In_794,In_197);
xnor U2132 (N_2132,In_1968,In_205);
or U2133 (N_2133,In_1303,In_711);
xor U2134 (N_2134,In_1585,In_1251);
or U2135 (N_2135,In_198,In_1986);
or U2136 (N_2136,In_1829,In_1748);
and U2137 (N_2137,In_810,In_1185);
xor U2138 (N_2138,In_1735,In_1976);
xnor U2139 (N_2139,In_393,In_936);
and U2140 (N_2140,In_1749,In_895);
nand U2141 (N_2141,In_1204,In_1475);
xnor U2142 (N_2142,In_23,In_1362);
nor U2143 (N_2143,In_592,In_1111);
nor U2144 (N_2144,In_1262,In_286);
nor U2145 (N_2145,In_1701,In_1983);
or U2146 (N_2146,In_1677,In_1543);
nand U2147 (N_2147,In_1752,In_538);
or U2148 (N_2148,In_1714,In_1400);
nand U2149 (N_2149,In_1515,In_521);
nand U2150 (N_2150,In_17,In_1552);
nand U2151 (N_2151,In_1523,In_1007);
xnor U2152 (N_2152,In_1603,In_1245);
nand U2153 (N_2153,In_1244,In_701);
nand U2154 (N_2154,In_291,In_1177);
nand U2155 (N_2155,In_536,In_743);
nand U2156 (N_2156,In_1886,In_1576);
nor U2157 (N_2157,In_409,In_1334);
nor U2158 (N_2158,In_655,In_469);
or U2159 (N_2159,In_1417,In_1351);
nand U2160 (N_2160,In_1579,In_1172);
nor U2161 (N_2161,In_1846,In_1764);
nor U2162 (N_2162,In_269,In_1530);
nor U2163 (N_2163,In_456,In_1972);
nor U2164 (N_2164,In_1666,In_1595);
nor U2165 (N_2165,In_184,In_678);
nand U2166 (N_2166,In_1662,In_1086);
or U2167 (N_2167,In_1897,In_1447);
nand U2168 (N_2168,In_53,In_279);
xnor U2169 (N_2169,In_1077,In_36);
nand U2170 (N_2170,In_1518,In_1977);
or U2171 (N_2171,In_473,In_1097);
nand U2172 (N_2172,In_502,In_1585);
or U2173 (N_2173,In_1853,In_43);
and U2174 (N_2174,In_1598,In_215);
xor U2175 (N_2175,In_674,In_502);
or U2176 (N_2176,In_1807,In_983);
xnor U2177 (N_2177,In_1248,In_1505);
or U2178 (N_2178,In_1732,In_1138);
and U2179 (N_2179,In_1610,In_314);
nor U2180 (N_2180,In_1338,In_1951);
xor U2181 (N_2181,In_1626,In_1305);
nor U2182 (N_2182,In_593,In_1588);
and U2183 (N_2183,In_209,In_258);
nand U2184 (N_2184,In_1188,In_1240);
or U2185 (N_2185,In_1722,In_1793);
and U2186 (N_2186,In_45,In_1533);
and U2187 (N_2187,In_225,In_181);
or U2188 (N_2188,In_1219,In_1013);
and U2189 (N_2189,In_189,In_198);
and U2190 (N_2190,In_502,In_692);
nor U2191 (N_2191,In_355,In_1198);
or U2192 (N_2192,In_1954,In_1210);
nor U2193 (N_2193,In_693,In_1990);
xnor U2194 (N_2194,In_1081,In_137);
xnor U2195 (N_2195,In_1271,In_1748);
or U2196 (N_2196,In_1220,In_994);
or U2197 (N_2197,In_626,In_834);
and U2198 (N_2198,In_1671,In_1241);
nor U2199 (N_2199,In_1855,In_407);
or U2200 (N_2200,In_1886,In_1979);
nand U2201 (N_2201,In_1511,In_189);
and U2202 (N_2202,In_798,In_1909);
xnor U2203 (N_2203,In_1211,In_452);
xor U2204 (N_2204,In_1756,In_433);
or U2205 (N_2205,In_678,In_908);
xor U2206 (N_2206,In_1606,In_1675);
and U2207 (N_2207,In_919,In_1106);
xnor U2208 (N_2208,In_1863,In_954);
nor U2209 (N_2209,In_1225,In_1436);
nand U2210 (N_2210,In_199,In_204);
nand U2211 (N_2211,In_1415,In_1206);
nor U2212 (N_2212,In_1094,In_1185);
and U2213 (N_2213,In_942,In_873);
and U2214 (N_2214,In_1388,In_536);
nor U2215 (N_2215,In_1570,In_103);
xor U2216 (N_2216,In_1330,In_241);
or U2217 (N_2217,In_1646,In_1272);
or U2218 (N_2218,In_394,In_1963);
nor U2219 (N_2219,In_626,In_299);
nor U2220 (N_2220,In_496,In_1021);
or U2221 (N_2221,In_756,In_974);
or U2222 (N_2222,In_213,In_111);
or U2223 (N_2223,In_1719,In_836);
nor U2224 (N_2224,In_1854,In_1005);
nor U2225 (N_2225,In_1478,In_846);
nand U2226 (N_2226,In_511,In_585);
or U2227 (N_2227,In_23,In_1794);
and U2228 (N_2228,In_1344,In_383);
nand U2229 (N_2229,In_1332,In_1586);
and U2230 (N_2230,In_1429,In_1311);
nand U2231 (N_2231,In_1857,In_1817);
xnor U2232 (N_2232,In_519,In_1829);
nand U2233 (N_2233,In_544,In_1070);
xnor U2234 (N_2234,In_184,In_1978);
xnor U2235 (N_2235,In_216,In_1911);
and U2236 (N_2236,In_190,In_5);
nor U2237 (N_2237,In_340,In_1634);
nand U2238 (N_2238,In_1482,In_1442);
nor U2239 (N_2239,In_1193,In_1645);
nand U2240 (N_2240,In_560,In_829);
and U2241 (N_2241,In_1978,In_1829);
xor U2242 (N_2242,In_39,In_1499);
nor U2243 (N_2243,In_748,In_1327);
and U2244 (N_2244,In_521,In_777);
and U2245 (N_2245,In_1809,In_1608);
nor U2246 (N_2246,In_967,In_928);
nand U2247 (N_2247,In_482,In_1833);
and U2248 (N_2248,In_906,In_481);
nand U2249 (N_2249,In_715,In_1681);
nor U2250 (N_2250,In_1504,In_682);
xnor U2251 (N_2251,In_1924,In_806);
nor U2252 (N_2252,In_1202,In_1952);
or U2253 (N_2253,In_303,In_1600);
and U2254 (N_2254,In_1700,In_230);
nor U2255 (N_2255,In_239,In_345);
or U2256 (N_2256,In_1329,In_67);
and U2257 (N_2257,In_1485,In_49);
nand U2258 (N_2258,In_383,In_1393);
nand U2259 (N_2259,In_1084,In_1110);
nor U2260 (N_2260,In_992,In_1748);
and U2261 (N_2261,In_907,In_1981);
or U2262 (N_2262,In_1882,In_309);
and U2263 (N_2263,In_1889,In_1433);
nand U2264 (N_2264,In_415,In_446);
and U2265 (N_2265,In_969,In_97);
and U2266 (N_2266,In_678,In_1635);
nand U2267 (N_2267,In_1164,In_1655);
and U2268 (N_2268,In_1992,In_1330);
and U2269 (N_2269,In_72,In_1659);
nand U2270 (N_2270,In_1317,In_641);
and U2271 (N_2271,In_445,In_1386);
nand U2272 (N_2272,In_174,In_937);
or U2273 (N_2273,In_1355,In_1840);
xnor U2274 (N_2274,In_594,In_1291);
nor U2275 (N_2275,In_1536,In_481);
nand U2276 (N_2276,In_1546,In_317);
xnor U2277 (N_2277,In_1237,In_269);
or U2278 (N_2278,In_777,In_1632);
nor U2279 (N_2279,In_1333,In_376);
nor U2280 (N_2280,In_1686,In_560);
nor U2281 (N_2281,In_1014,In_1746);
xor U2282 (N_2282,In_75,In_676);
nand U2283 (N_2283,In_213,In_1199);
xor U2284 (N_2284,In_542,In_1389);
xor U2285 (N_2285,In_65,In_1318);
nor U2286 (N_2286,In_1083,In_779);
nor U2287 (N_2287,In_1324,In_506);
or U2288 (N_2288,In_667,In_277);
or U2289 (N_2289,In_1469,In_1704);
and U2290 (N_2290,In_73,In_1543);
nor U2291 (N_2291,In_1769,In_1822);
nor U2292 (N_2292,In_159,In_701);
xnor U2293 (N_2293,In_1092,In_1515);
nor U2294 (N_2294,In_1,In_249);
or U2295 (N_2295,In_770,In_1446);
and U2296 (N_2296,In_694,In_1615);
nor U2297 (N_2297,In_652,In_153);
nand U2298 (N_2298,In_741,In_20);
and U2299 (N_2299,In_774,In_1688);
nand U2300 (N_2300,In_523,In_168);
nand U2301 (N_2301,In_1551,In_221);
and U2302 (N_2302,In_1459,In_1864);
or U2303 (N_2303,In_1764,In_78);
and U2304 (N_2304,In_1270,In_1752);
nor U2305 (N_2305,In_873,In_1713);
xnor U2306 (N_2306,In_1066,In_1960);
xor U2307 (N_2307,In_1599,In_141);
nand U2308 (N_2308,In_1950,In_890);
and U2309 (N_2309,In_712,In_1363);
or U2310 (N_2310,In_69,In_1754);
nor U2311 (N_2311,In_1636,In_1792);
nor U2312 (N_2312,In_17,In_1565);
nor U2313 (N_2313,In_542,In_1175);
nand U2314 (N_2314,In_151,In_972);
or U2315 (N_2315,In_1383,In_983);
nand U2316 (N_2316,In_648,In_1912);
and U2317 (N_2317,In_1967,In_1775);
nand U2318 (N_2318,In_579,In_1531);
xnor U2319 (N_2319,In_882,In_69);
or U2320 (N_2320,In_307,In_271);
and U2321 (N_2321,In_1364,In_63);
and U2322 (N_2322,In_28,In_1137);
xor U2323 (N_2323,In_435,In_1863);
xnor U2324 (N_2324,In_569,In_1912);
nand U2325 (N_2325,In_1142,In_1724);
or U2326 (N_2326,In_921,In_949);
or U2327 (N_2327,In_205,In_746);
and U2328 (N_2328,In_1342,In_511);
nor U2329 (N_2329,In_33,In_1384);
nand U2330 (N_2330,In_1108,In_1198);
xnor U2331 (N_2331,In_151,In_1778);
xnor U2332 (N_2332,In_327,In_24);
or U2333 (N_2333,In_1062,In_1030);
and U2334 (N_2334,In_868,In_1634);
or U2335 (N_2335,In_1161,In_148);
xor U2336 (N_2336,In_622,In_1402);
nand U2337 (N_2337,In_45,In_1307);
nor U2338 (N_2338,In_1090,In_1699);
nor U2339 (N_2339,In_1545,In_372);
or U2340 (N_2340,In_1414,In_1578);
and U2341 (N_2341,In_1627,In_1829);
and U2342 (N_2342,In_27,In_1114);
or U2343 (N_2343,In_1913,In_193);
and U2344 (N_2344,In_365,In_1517);
nor U2345 (N_2345,In_304,In_14);
xor U2346 (N_2346,In_1309,In_811);
nand U2347 (N_2347,In_203,In_1018);
and U2348 (N_2348,In_685,In_1448);
or U2349 (N_2349,In_1380,In_692);
xor U2350 (N_2350,In_761,In_1273);
nand U2351 (N_2351,In_723,In_1316);
nor U2352 (N_2352,In_1464,In_1361);
xnor U2353 (N_2353,In_619,In_640);
nand U2354 (N_2354,In_1783,In_1422);
nand U2355 (N_2355,In_407,In_1514);
xnor U2356 (N_2356,In_196,In_123);
nand U2357 (N_2357,In_1573,In_1057);
nor U2358 (N_2358,In_1736,In_114);
nand U2359 (N_2359,In_1431,In_1022);
nor U2360 (N_2360,In_1487,In_1799);
and U2361 (N_2361,In_1052,In_1241);
and U2362 (N_2362,In_1561,In_61);
and U2363 (N_2363,In_1284,In_1002);
and U2364 (N_2364,In_1304,In_1837);
xnor U2365 (N_2365,In_1745,In_979);
nand U2366 (N_2366,In_292,In_379);
or U2367 (N_2367,In_1661,In_259);
nand U2368 (N_2368,In_322,In_1362);
xnor U2369 (N_2369,In_1096,In_205);
nor U2370 (N_2370,In_698,In_1234);
and U2371 (N_2371,In_754,In_1234);
or U2372 (N_2372,In_1508,In_1891);
nor U2373 (N_2373,In_1693,In_1042);
nor U2374 (N_2374,In_635,In_959);
and U2375 (N_2375,In_582,In_1524);
nand U2376 (N_2376,In_1904,In_1741);
nor U2377 (N_2377,In_1910,In_342);
or U2378 (N_2378,In_1204,In_71);
nand U2379 (N_2379,In_512,In_1289);
nand U2380 (N_2380,In_1747,In_1081);
or U2381 (N_2381,In_696,In_293);
nor U2382 (N_2382,In_1625,In_1647);
xor U2383 (N_2383,In_731,In_1481);
and U2384 (N_2384,In_250,In_1888);
and U2385 (N_2385,In_691,In_718);
and U2386 (N_2386,In_801,In_1790);
xnor U2387 (N_2387,In_1736,In_802);
xnor U2388 (N_2388,In_887,In_952);
nor U2389 (N_2389,In_384,In_308);
xor U2390 (N_2390,In_1280,In_413);
nand U2391 (N_2391,In_1682,In_589);
nor U2392 (N_2392,In_1073,In_1138);
xnor U2393 (N_2393,In_74,In_1105);
and U2394 (N_2394,In_768,In_1426);
nand U2395 (N_2395,In_596,In_878);
nor U2396 (N_2396,In_148,In_957);
nand U2397 (N_2397,In_1660,In_857);
xnor U2398 (N_2398,In_1107,In_1041);
xnor U2399 (N_2399,In_1690,In_745);
nand U2400 (N_2400,In_1090,In_1851);
or U2401 (N_2401,In_203,In_1921);
and U2402 (N_2402,In_1059,In_1171);
xnor U2403 (N_2403,In_1347,In_1651);
nor U2404 (N_2404,In_106,In_1531);
and U2405 (N_2405,In_1093,In_11);
nand U2406 (N_2406,In_1367,In_1989);
or U2407 (N_2407,In_799,In_1105);
nand U2408 (N_2408,In_643,In_930);
xor U2409 (N_2409,In_848,In_1359);
or U2410 (N_2410,In_842,In_1644);
nand U2411 (N_2411,In_1100,In_915);
xor U2412 (N_2412,In_626,In_91);
xnor U2413 (N_2413,In_1575,In_1714);
xor U2414 (N_2414,In_1764,In_1952);
or U2415 (N_2415,In_460,In_1770);
xor U2416 (N_2416,In_1513,In_1415);
and U2417 (N_2417,In_1925,In_170);
xor U2418 (N_2418,In_1320,In_843);
nor U2419 (N_2419,In_1379,In_1897);
nor U2420 (N_2420,In_1171,In_1428);
xnor U2421 (N_2421,In_1846,In_1879);
xor U2422 (N_2422,In_1484,In_1154);
xnor U2423 (N_2423,In_1356,In_1548);
nor U2424 (N_2424,In_1385,In_978);
nor U2425 (N_2425,In_1443,In_113);
or U2426 (N_2426,In_78,In_1378);
xnor U2427 (N_2427,In_913,In_1434);
nand U2428 (N_2428,In_1532,In_458);
or U2429 (N_2429,In_814,In_227);
nor U2430 (N_2430,In_45,In_339);
nand U2431 (N_2431,In_1614,In_1725);
xnor U2432 (N_2432,In_305,In_1419);
nor U2433 (N_2433,In_1833,In_1826);
and U2434 (N_2434,In_274,In_908);
nor U2435 (N_2435,In_1119,In_76);
or U2436 (N_2436,In_335,In_1432);
nand U2437 (N_2437,In_499,In_1693);
nor U2438 (N_2438,In_660,In_725);
nor U2439 (N_2439,In_1606,In_330);
or U2440 (N_2440,In_179,In_1336);
or U2441 (N_2441,In_904,In_923);
or U2442 (N_2442,In_1210,In_1321);
and U2443 (N_2443,In_690,In_620);
nand U2444 (N_2444,In_529,In_493);
xor U2445 (N_2445,In_46,In_234);
nor U2446 (N_2446,In_438,In_615);
xnor U2447 (N_2447,In_1976,In_1140);
and U2448 (N_2448,In_353,In_1658);
xnor U2449 (N_2449,In_1918,In_1282);
nor U2450 (N_2450,In_1937,In_1154);
xor U2451 (N_2451,In_1319,In_899);
xnor U2452 (N_2452,In_47,In_1947);
xor U2453 (N_2453,In_489,In_1676);
xnor U2454 (N_2454,In_290,In_938);
and U2455 (N_2455,In_1890,In_1469);
xor U2456 (N_2456,In_531,In_1851);
xnor U2457 (N_2457,In_764,In_435);
and U2458 (N_2458,In_614,In_1091);
or U2459 (N_2459,In_540,In_847);
nor U2460 (N_2460,In_172,In_1780);
and U2461 (N_2461,In_48,In_1440);
and U2462 (N_2462,In_931,In_1026);
or U2463 (N_2463,In_1784,In_1090);
or U2464 (N_2464,In_554,In_349);
and U2465 (N_2465,In_182,In_1389);
xnor U2466 (N_2466,In_631,In_847);
and U2467 (N_2467,In_911,In_1204);
and U2468 (N_2468,In_1929,In_1153);
nand U2469 (N_2469,In_120,In_1950);
nand U2470 (N_2470,In_1783,In_1509);
xor U2471 (N_2471,In_1929,In_69);
nor U2472 (N_2472,In_1704,In_1641);
and U2473 (N_2473,In_1307,In_1524);
nand U2474 (N_2474,In_47,In_633);
nand U2475 (N_2475,In_681,In_815);
or U2476 (N_2476,In_174,In_1667);
nand U2477 (N_2477,In_344,In_1328);
nand U2478 (N_2478,In_806,In_723);
or U2479 (N_2479,In_55,In_1153);
and U2480 (N_2480,In_43,In_1451);
xnor U2481 (N_2481,In_403,In_76);
xnor U2482 (N_2482,In_1683,In_1178);
or U2483 (N_2483,In_741,In_1123);
xnor U2484 (N_2484,In_354,In_1383);
and U2485 (N_2485,In_175,In_1736);
nor U2486 (N_2486,In_1921,In_453);
nand U2487 (N_2487,In_1692,In_276);
nand U2488 (N_2488,In_755,In_1168);
xnor U2489 (N_2489,In_707,In_1637);
or U2490 (N_2490,In_1123,In_578);
and U2491 (N_2491,In_1428,In_797);
xnor U2492 (N_2492,In_348,In_556);
or U2493 (N_2493,In_1645,In_1254);
nor U2494 (N_2494,In_940,In_827);
xnor U2495 (N_2495,In_1192,In_323);
or U2496 (N_2496,In_774,In_156);
nor U2497 (N_2497,In_1487,In_1817);
nor U2498 (N_2498,In_450,In_1065);
and U2499 (N_2499,In_92,In_1572);
or U2500 (N_2500,In_525,In_1454);
and U2501 (N_2501,In_1286,In_418);
xnor U2502 (N_2502,In_431,In_1627);
and U2503 (N_2503,In_1046,In_659);
xnor U2504 (N_2504,In_823,In_890);
or U2505 (N_2505,In_741,In_72);
nor U2506 (N_2506,In_148,In_1239);
or U2507 (N_2507,In_1049,In_662);
nand U2508 (N_2508,In_1492,In_516);
or U2509 (N_2509,In_1575,In_1870);
xor U2510 (N_2510,In_1822,In_1296);
or U2511 (N_2511,In_343,In_1687);
nor U2512 (N_2512,In_1601,In_202);
nand U2513 (N_2513,In_1354,In_1391);
nand U2514 (N_2514,In_1320,In_321);
xor U2515 (N_2515,In_1387,In_1813);
nor U2516 (N_2516,In_1303,In_1383);
nor U2517 (N_2517,In_1178,In_1246);
and U2518 (N_2518,In_520,In_1663);
or U2519 (N_2519,In_313,In_302);
nand U2520 (N_2520,In_192,In_1757);
xor U2521 (N_2521,In_1048,In_1362);
nand U2522 (N_2522,In_1953,In_1287);
xor U2523 (N_2523,In_1614,In_1101);
nor U2524 (N_2524,In_344,In_1666);
nor U2525 (N_2525,In_932,In_1178);
nand U2526 (N_2526,In_558,In_1636);
and U2527 (N_2527,In_1374,In_1304);
or U2528 (N_2528,In_1041,In_29);
nor U2529 (N_2529,In_188,In_222);
or U2530 (N_2530,In_992,In_1857);
nand U2531 (N_2531,In_1706,In_530);
xnor U2532 (N_2532,In_1894,In_185);
or U2533 (N_2533,In_253,In_972);
or U2534 (N_2534,In_829,In_664);
and U2535 (N_2535,In_1855,In_720);
nor U2536 (N_2536,In_1559,In_1211);
or U2537 (N_2537,In_860,In_32);
nand U2538 (N_2538,In_1976,In_580);
nor U2539 (N_2539,In_1737,In_1666);
xor U2540 (N_2540,In_1678,In_1730);
or U2541 (N_2541,In_231,In_931);
and U2542 (N_2542,In_322,In_713);
nor U2543 (N_2543,In_261,In_508);
or U2544 (N_2544,In_1894,In_1665);
or U2545 (N_2545,In_989,In_623);
nor U2546 (N_2546,In_1539,In_1940);
and U2547 (N_2547,In_1487,In_1674);
or U2548 (N_2548,In_717,In_1504);
nand U2549 (N_2549,In_1148,In_1774);
and U2550 (N_2550,In_18,In_15);
nor U2551 (N_2551,In_977,In_43);
nor U2552 (N_2552,In_1958,In_538);
nor U2553 (N_2553,In_262,In_1018);
xor U2554 (N_2554,In_1175,In_346);
and U2555 (N_2555,In_1204,In_132);
nor U2556 (N_2556,In_151,In_1046);
nand U2557 (N_2557,In_1182,In_64);
or U2558 (N_2558,In_17,In_118);
nand U2559 (N_2559,In_762,In_500);
nand U2560 (N_2560,In_1854,In_225);
nor U2561 (N_2561,In_1437,In_631);
and U2562 (N_2562,In_740,In_703);
nand U2563 (N_2563,In_1790,In_1149);
nor U2564 (N_2564,In_1493,In_743);
nand U2565 (N_2565,In_192,In_119);
and U2566 (N_2566,In_1516,In_1952);
or U2567 (N_2567,In_1251,In_483);
xnor U2568 (N_2568,In_1336,In_1692);
xnor U2569 (N_2569,In_1902,In_457);
nand U2570 (N_2570,In_1257,In_1339);
and U2571 (N_2571,In_1697,In_560);
nand U2572 (N_2572,In_1469,In_1962);
or U2573 (N_2573,In_1087,In_1094);
xnor U2574 (N_2574,In_1910,In_1636);
nand U2575 (N_2575,In_1099,In_1572);
xnor U2576 (N_2576,In_1357,In_1883);
xnor U2577 (N_2577,In_862,In_1693);
and U2578 (N_2578,In_284,In_1336);
or U2579 (N_2579,In_1460,In_1637);
or U2580 (N_2580,In_661,In_1893);
or U2581 (N_2581,In_557,In_1042);
and U2582 (N_2582,In_776,In_1162);
nand U2583 (N_2583,In_1921,In_741);
xor U2584 (N_2584,In_1203,In_455);
nor U2585 (N_2585,In_1110,In_1498);
and U2586 (N_2586,In_1858,In_874);
nand U2587 (N_2587,In_1080,In_1898);
nand U2588 (N_2588,In_116,In_695);
or U2589 (N_2589,In_69,In_1150);
xor U2590 (N_2590,In_1589,In_544);
xor U2591 (N_2591,In_1448,In_1740);
or U2592 (N_2592,In_1467,In_407);
nor U2593 (N_2593,In_357,In_1487);
nand U2594 (N_2594,In_428,In_1343);
and U2595 (N_2595,In_1783,In_906);
nand U2596 (N_2596,In_1423,In_1379);
or U2597 (N_2597,In_271,In_1417);
or U2598 (N_2598,In_1243,In_228);
and U2599 (N_2599,In_1041,In_763);
xor U2600 (N_2600,In_1708,In_404);
nor U2601 (N_2601,In_1259,In_616);
or U2602 (N_2602,In_1834,In_492);
and U2603 (N_2603,In_309,In_1520);
xnor U2604 (N_2604,In_671,In_1168);
xnor U2605 (N_2605,In_1923,In_1968);
and U2606 (N_2606,In_1218,In_648);
or U2607 (N_2607,In_1301,In_1594);
nor U2608 (N_2608,In_1013,In_745);
xnor U2609 (N_2609,In_1649,In_245);
and U2610 (N_2610,In_1903,In_569);
nand U2611 (N_2611,In_1896,In_1358);
nand U2612 (N_2612,In_1580,In_1600);
xor U2613 (N_2613,In_1758,In_1982);
or U2614 (N_2614,In_1517,In_1316);
or U2615 (N_2615,In_1288,In_119);
and U2616 (N_2616,In_632,In_342);
and U2617 (N_2617,In_1922,In_1864);
nor U2618 (N_2618,In_1305,In_1296);
or U2619 (N_2619,In_1021,In_1409);
xnor U2620 (N_2620,In_1233,In_680);
or U2621 (N_2621,In_492,In_405);
nor U2622 (N_2622,In_987,In_1333);
xor U2623 (N_2623,In_664,In_789);
or U2624 (N_2624,In_131,In_634);
or U2625 (N_2625,In_665,In_206);
nor U2626 (N_2626,In_1155,In_1733);
nand U2627 (N_2627,In_651,In_1201);
or U2628 (N_2628,In_1890,In_1356);
nand U2629 (N_2629,In_1204,In_671);
xnor U2630 (N_2630,In_1946,In_1304);
nand U2631 (N_2631,In_851,In_900);
or U2632 (N_2632,In_1999,In_1495);
and U2633 (N_2633,In_1118,In_1478);
or U2634 (N_2634,In_939,In_208);
nand U2635 (N_2635,In_1475,In_162);
nand U2636 (N_2636,In_946,In_1394);
xnor U2637 (N_2637,In_1677,In_215);
nand U2638 (N_2638,In_825,In_929);
nand U2639 (N_2639,In_127,In_1790);
or U2640 (N_2640,In_87,In_1754);
nand U2641 (N_2641,In_1691,In_952);
nand U2642 (N_2642,In_169,In_843);
xor U2643 (N_2643,In_732,In_1937);
nor U2644 (N_2644,In_1261,In_1771);
or U2645 (N_2645,In_1452,In_162);
and U2646 (N_2646,In_663,In_616);
nand U2647 (N_2647,In_651,In_1203);
nand U2648 (N_2648,In_384,In_1413);
and U2649 (N_2649,In_1987,In_908);
or U2650 (N_2650,In_1344,In_402);
xnor U2651 (N_2651,In_957,In_1500);
and U2652 (N_2652,In_1115,In_1575);
and U2653 (N_2653,In_704,In_1017);
nand U2654 (N_2654,In_255,In_1281);
or U2655 (N_2655,In_1377,In_1924);
and U2656 (N_2656,In_95,In_1508);
nand U2657 (N_2657,In_1042,In_1572);
and U2658 (N_2658,In_1444,In_79);
xnor U2659 (N_2659,In_392,In_1163);
nand U2660 (N_2660,In_1818,In_947);
nor U2661 (N_2661,In_637,In_531);
or U2662 (N_2662,In_1402,In_1580);
xor U2663 (N_2663,In_1965,In_1938);
nand U2664 (N_2664,In_1270,In_949);
nand U2665 (N_2665,In_1338,In_491);
and U2666 (N_2666,In_1393,In_1603);
and U2667 (N_2667,In_24,In_1825);
xnor U2668 (N_2668,In_595,In_293);
and U2669 (N_2669,In_734,In_323);
nand U2670 (N_2670,In_1732,In_262);
nand U2671 (N_2671,In_596,In_1908);
nor U2672 (N_2672,In_1936,In_849);
xnor U2673 (N_2673,In_739,In_194);
or U2674 (N_2674,In_546,In_718);
xor U2675 (N_2675,In_1493,In_1797);
or U2676 (N_2676,In_250,In_1056);
or U2677 (N_2677,In_1770,In_1553);
and U2678 (N_2678,In_1144,In_1676);
nand U2679 (N_2679,In_1082,In_137);
nand U2680 (N_2680,In_881,In_1090);
nor U2681 (N_2681,In_405,In_184);
nand U2682 (N_2682,In_808,In_1457);
nand U2683 (N_2683,In_698,In_435);
nand U2684 (N_2684,In_653,In_472);
nand U2685 (N_2685,In_22,In_309);
and U2686 (N_2686,In_861,In_1501);
nand U2687 (N_2687,In_1699,In_1934);
xor U2688 (N_2688,In_747,In_151);
and U2689 (N_2689,In_298,In_1089);
nor U2690 (N_2690,In_866,In_295);
nor U2691 (N_2691,In_1693,In_328);
xor U2692 (N_2692,In_557,In_611);
nor U2693 (N_2693,In_784,In_626);
and U2694 (N_2694,In_1405,In_1370);
nand U2695 (N_2695,In_1528,In_397);
or U2696 (N_2696,In_829,In_1842);
xnor U2697 (N_2697,In_1804,In_566);
or U2698 (N_2698,In_990,In_1522);
nand U2699 (N_2699,In_909,In_990);
nand U2700 (N_2700,In_1499,In_1621);
or U2701 (N_2701,In_1280,In_1959);
or U2702 (N_2702,In_187,In_1963);
or U2703 (N_2703,In_225,In_1519);
or U2704 (N_2704,In_1309,In_1720);
and U2705 (N_2705,In_519,In_1028);
or U2706 (N_2706,In_904,In_1304);
xor U2707 (N_2707,In_378,In_954);
nand U2708 (N_2708,In_998,In_758);
nor U2709 (N_2709,In_555,In_823);
nor U2710 (N_2710,In_694,In_465);
nor U2711 (N_2711,In_921,In_1645);
nand U2712 (N_2712,In_1350,In_268);
nand U2713 (N_2713,In_1232,In_1416);
and U2714 (N_2714,In_1259,In_115);
xor U2715 (N_2715,In_1337,In_1575);
and U2716 (N_2716,In_1377,In_1523);
or U2717 (N_2717,In_1733,In_670);
nand U2718 (N_2718,In_1198,In_38);
nand U2719 (N_2719,In_1590,In_1532);
nand U2720 (N_2720,In_1173,In_371);
xnor U2721 (N_2721,In_1469,In_934);
or U2722 (N_2722,In_788,In_89);
nor U2723 (N_2723,In_470,In_137);
nand U2724 (N_2724,In_1538,In_1959);
or U2725 (N_2725,In_1308,In_309);
nand U2726 (N_2726,In_1367,In_72);
nand U2727 (N_2727,In_122,In_1900);
or U2728 (N_2728,In_1810,In_1187);
xor U2729 (N_2729,In_1887,In_356);
or U2730 (N_2730,In_1321,In_561);
or U2731 (N_2731,In_682,In_1038);
or U2732 (N_2732,In_1649,In_702);
xor U2733 (N_2733,In_475,In_76);
or U2734 (N_2734,In_174,In_614);
nor U2735 (N_2735,In_1010,In_554);
or U2736 (N_2736,In_615,In_1449);
xor U2737 (N_2737,In_252,In_1815);
nor U2738 (N_2738,In_1650,In_673);
xnor U2739 (N_2739,In_672,In_958);
and U2740 (N_2740,In_1377,In_549);
nand U2741 (N_2741,In_1251,In_1714);
nor U2742 (N_2742,In_69,In_565);
or U2743 (N_2743,In_1082,In_1704);
nand U2744 (N_2744,In_484,In_880);
and U2745 (N_2745,In_332,In_1745);
xor U2746 (N_2746,In_602,In_1925);
nand U2747 (N_2747,In_730,In_1972);
and U2748 (N_2748,In_1168,In_1190);
xnor U2749 (N_2749,In_1183,In_1015);
or U2750 (N_2750,In_666,In_1951);
and U2751 (N_2751,In_1687,In_1013);
nor U2752 (N_2752,In_143,In_1629);
xor U2753 (N_2753,In_1507,In_210);
or U2754 (N_2754,In_158,In_1696);
xor U2755 (N_2755,In_136,In_812);
xor U2756 (N_2756,In_703,In_1315);
xor U2757 (N_2757,In_1563,In_618);
nand U2758 (N_2758,In_1698,In_1547);
xnor U2759 (N_2759,In_55,In_1998);
nor U2760 (N_2760,In_1653,In_15);
nand U2761 (N_2761,In_941,In_233);
or U2762 (N_2762,In_97,In_1960);
and U2763 (N_2763,In_1305,In_1018);
nand U2764 (N_2764,In_788,In_203);
and U2765 (N_2765,In_906,In_762);
nor U2766 (N_2766,In_988,In_1555);
and U2767 (N_2767,In_1084,In_1163);
and U2768 (N_2768,In_1707,In_333);
nor U2769 (N_2769,In_1975,In_817);
and U2770 (N_2770,In_372,In_46);
and U2771 (N_2771,In_1841,In_790);
nand U2772 (N_2772,In_1272,In_356);
or U2773 (N_2773,In_385,In_1652);
nor U2774 (N_2774,In_1761,In_1229);
nor U2775 (N_2775,In_1136,In_194);
nand U2776 (N_2776,In_1892,In_1169);
nand U2777 (N_2777,In_1209,In_377);
xnor U2778 (N_2778,In_661,In_1282);
or U2779 (N_2779,In_1817,In_691);
nor U2780 (N_2780,In_1626,In_459);
xor U2781 (N_2781,In_375,In_1719);
nand U2782 (N_2782,In_962,In_543);
xor U2783 (N_2783,In_1052,In_783);
or U2784 (N_2784,In_1165,In_582);
nand U2785 (N_2785,In_1093,In_602);
nor U2786 (N_2786,In_207,In_1753);
nand U2787 (N_2787,In_1252,In_523);
and U2788 (N_2788,In_1484,In_1851);
nor U2789 (N_2789,In_1898,In_1843);
nand U2790 (N_2790,In_1258,In_92);
or U2791 (N_2791,In_1334,In_32);
nand U2792 (N_2792,In_1752,In_468);
nand U2793 (N_2793,In_375,In_197);
nand U2794 (N_2794,In_1525,In_1457);
or U2795 (N_2795,In_307,In_1172);
nor U2796 (N_2796,In_1585,In_8);
or U2797 (N_2797,In_529,In_1276);
nand U2798 (N_2798,In_1021,In_50);
nand U2799 (N_2799,In_1500,In_1071);
nor U2800 (N_2800,In_930,In_95);
or U2801 (N_2801,In_50,In_863);
xor U2802 (N_2802,In_285,In_1329);
xnor U2803 (N_2803,In_1512,In_416);
nor U2804 (N_2804,In_1724,In_735);
and U2805 (N_2805,In_905,In_1795);
and U2806 (N_2806,In_1288,In_174);
nor U2807 (N_2807,In_1072,In_1037);
nand U2808 (N_2808,In_1337,In_1817);
xor U2809 (N_2809,In_1497,In_350);
and U2810 (N_2810,In_1269,In_1176);
and U2811 (N_2811,In_1866,In_1222);
or U2812 (N_2812,In_1942,In_1709);
xor U2813 (N_2813,In_470,In_1969);
and U2814 (N_2814,In_421,In_699);
and U2815 (N_2815,In_1016,In_350);
xnor U2816 (N_2816,In_544,In_139);
nor U2817 (N_2817,In_833,In_171);
xnor U2818 (N_2818,In_1465,In_605);
nand U2819 (N_2819,In_1359,In_177);
or U2820 (N_2820,In_1220,In_1564);
xnor U2821 (N_2821,In_1380,In_224);
nand U2822 (N_2822,In_253,In_931);
or U2823 (N_2823,In_520,In_400);
nor U2824 (N_2824,In_1158,In_213);
or U2825 (N_2825,In_1122,In_1449);
and U2826 (N_2826,In_1575,In_158);
nand U2827 (N_2827,In_1220,In_1612);
nor U2828 (N_2828,In_1018,In_1422);
xnor U2829 (N_2829,In_14,In_227);
nand U2830 (N_2830,In_1950,In_1245);
nor U2831 (N_2831,In_335,In_1502);
or U2832 (N_2832,In_760,In_1014);
nor U2833 (N_2833,In_784,In_594);
nand U2834 (N_2834,In_657,In_974);
or U2835 (N_2835,In_379,In_592);
and U2836 (N_2836,In_1350,In_836);
xor U2837 (N_2837,In_1374,In_1297);
nor U2838 (N_2838,In_1864,In_665);
nor U2839 (N_2839,In_296,In_1585);
and U2840 (N_2840,In_1703,In_1800);
or U2841 (N_2841,In_283,In_1666);
nor U2842 (N_2842,In_1733,In_1204);
xnor U2843 (N_2843,In_315,In_1654);
or U2844 (N_2844,In_628,In_1505);
or U2845 (N_2845,In_436,In_1348);
or U2846 (N_2846,In_1565,In_541);
nor U2847 (N_2847,In_1014,In_1476);
nand U2848 (N_2848,In_1996,In_974);
or U2849 (N_2849,In_267,In_1607);
or U2850 (N_2850,In_1957,In_632);
and U2851 (N_2851,In_1464,In_1577);
and U2852 (N_2852,In_1947,In_291);
xnor U2853 (N_2853,In_1358,In_1793);
xor U2854 (N_2854,In_177,In_726);
and U2855 (N_2855,In_1269,In_386);
nor U2856 (N_2856,In_1298,In_108);
xor U2857 (N_2857,In_990,In_733);
nand U2858 (N_2858,In_340,In_1584);
nand U2859 (N_2859,In_1360,In_620);
or U2860 (N_2860,In_58,In_912);
or U2861 (N_2861,In_196,In_623);
xor U2862 (N_2862,In_372,In_541);
nand U2863 (N_2863,In_409,In_1850);
nor U2864 (N_2864,In_1827,In_1420);
xnor U2865 (N_2865,In_486,In_1234);
nand U2866 (N_2866,In_1930,In_1938);
nand U2867 (N_2867,In_1468,In_1629);
nor U2868 (N_2868,In_1358,In_822);
and U2869 (N_2869,In_1957,In_1403);
nand U2870 (N_2870,In_458,In_13);
nor U2871 (N_2871,In_1733,In_301);
and U2872 (N_2872,In_1892,In_396);
nor U2873 (N_2873,In_108,In_1797);
nand U2874 (N_2874,In_107,In_1312);
nand U2875 (N_2875,In_1978,In_59);
and U2876 (N_2876,In_830,In_849);
and U2877 (N_2877,In_1778,In_961);
nand U2878 (N_2878,In_1636,In_956);
nand U2879 (N_2879,In_1730,In_292);
nand U2880 (N_2880,In_1090,In_692);
nand U2881 (N_2881,In_1366,In_697);
nand U2882 (N_2882,In_209,In_1983);
or U2883 (N_2883,In_1,In_1969);
xor U2884 (N_2884,In_119,In_207);
nand U2885 (N_2885,In_1083,In_1377);
or U2886 (N_2886,In_306,In_823);
xor U2887 (N_2887,In_1801,In_1732);
and U2888 (N_2888,In_599,In_37);
xnor U2889 (N_2889,In_138,In_482);
xor U2890 (N_2890,In_1671,In_33);
or U2891 (N_2891,In_9,In_856);
and U2892 (N_2892,In_1928,In_1296);
nor U2893 (N_2893,In_1589,In_108);
nand U2894 (N_2894,In_1852,In_504);
or U2895 (N_2895,In_441,In_902);
nand U2896 (N_2896,In_130,In_1843);
nand U2897 (N_2897,In_1089,In_1347);
xnor U2898 (N_2898,In_990,In_600);
xor U2899 (N_2899,In_580,In_1443);
and U2900 (N_2900,In_121,In_1571);
or U2901 (N_2901,In_1673,In_349);
nor U2902 (N_2902,In_1955,In_903);
or U2903 (N_2903,In_863,In_1223);
or U2904 (N_2904,In_1289,In_906);
and U2905 (N_2905,In_1017,In_102);
and U2906 (N_2906,In_1373,In_484);
nor U2907 (N_2907,In_1490,In_663);
nor U2908 (N_2908,In_1846,In_1414);
nand U2909 (N_2909,In_1601,In_752);
xnor U2910 (N_2910,In_1606,In_197);
and U2911 (N_2911,In_1027,In_1105);
and U2912 (N_2912,In_1274,In_1450);
or U2913 (N_2913,In_846,In_1871);
or U2914 (N_2914,In_1476,In_1368);
nor U2915 (N_2915,In_1959,In_31);
or U2916 (N_2916,In_489,In_921);
nand U2917 (N_2917,In_1094,In_844);
and U2918 (N_2918,In_19,In_199);
xnor U2919 (N_2919,In_1896,In_293);
or U2920 (N_2920,In_1448,In_1703);
and U2921 (N_2921,In_1809,In_1469);
or U2922 (N_2922,In_331,In_728);
nor U2923 (N_2923,In_1078,In_882);
or U2924 (N_2924,In_880,In_128);
xor U2925 (N_2925,In_1442,In_1639);
and U2926 (N_2926,In_476,In_1581);
or U2927 (N_2927,In_1812,In_1898);
or U2928 (N_2928,In_10,In_928);
nand U2929 (N_2929,In_723,In_906);
or U2930 (N_2930,In_1630,In_666);
xnor U2931 (N_2931,In_863,In_495);
nand U2932 (N_2932,In_1934,In_764);
nor U2933 (N_2933,In_1971,In_902);
and U2934 (N_2934,In_1101,In_1088);
and U2935 (N_2935,In_1749,In_14);
and U2936 (N_2936,In_1787,In_1430);
xor U2937 (N_2937,In_1632,In_580);
xor U2938 (N_2938,In_1813,In_1708);
or U2939 (N_2939,In_1319,In_782);
or U2940 (N_2940,In_334,In_250);
nor U2941 (N_2941,In_611,In_1696);
nor U2942 (N_2942,In_701,In_459);
and U2943 (N_2943,In_1982,In_355);
or U2944 (N_2944,In_194,In_545);
and U2945 (N_2945,In_609,In_276);
and U2946 (N_2946,In_1285,In_274);
nand U2947 (N_2947,In_489,In_684);
or U2948 (N_2948,In_1043,In_1384);
and U2949 (N_2949,In_959,In_676);
xor U2950 (N_2950,In_1514,In_672);
xnor U2951 (N_2951,In_183,In_571);
nor U2952 (N_2952,In_553,In_751);
xnor U2953 (N_2953,In_186,In_1089);
xnor U2954 (N_2954,In_142,In_814);
nor U2955 (N_2955,In_187,In_320);
xor U2956 (N_2956,In_228,In_852);
nor U2957 (N_2957,In_1355,In_218);
nor U2958 (N_2958,In_370,In_333);
xor U2959 (N_2959,In_595,In_601);
nor U2960 (N_2960,In_56,In_1361);
and U2961 (N_2961,In_1725,In_1796);
nand U2962 (N_2962,In_126,In_1649);
xor U2963 (N_2963,In_1281,In_1070);
xnor U2964 (N_2964,In_1042,In_550);
xor U2965 (N_2965,In_1868,In_793);
xnor U2966 (N_2966,In_1134,In_1100);
and U2967 (N_2967,In_1940,In_1373);
xor U2968 (N_2968,In_869,In_1138);
and U2969 (N_2969,In_1290,In_1996);
and U2970 (N_2970,In_779,In_1802);
and U2971 (N_2971,In_1221,In_1714);
and U2972 (N_2972,In_1084,In_1331);
nor U2973 (N_2973,In_1116,In_92);
xnor U2974 (N_2974,In_3,In_326);
xor U2975 (N_2975,In_909,In_1327);
nand U2976 (N_2976,In_828,In_574);
xnor U2977 (N_2977,In_1540,In_1252);
nor U2978 (N_2978,In_1190,In_11);
or U2979 (N_2979,In_1909,In_431);
and U2980 (N_2980,In_1354,In_1654);
xnor U2981 (N_2981,In_1812,In_1534);
nand U2982 (N_2982,In_573,In_878);
xnor U2983 (N_2983,In_903,In_744);
nand U2984 (N_2984,In_1821,In_1456);
nand U2985 (N_2985,In_619,In_1319);
or U2986 (N_2986,In_1347,In_1708);
nand U2987 (N_2987,In_815,In_1575);
nor U2988 (N_2988,In_1656,In_982);
and U2989 (N_2989,In_167,In_1989);
xnor U2990 (N_2990,In_1890,In_82);
xnor U2991 (N_2991,In_684,In_1593);
nor U2992 (N_2992,In_1647,In_1426);
nand U2993 (N_2993,In_894,In_954);
xor U2994 (N_2994,In_1529,In_1428);
nor U2995 (N_2995,In_488,In_844);
xor U2996 (N_2996,In_624,In_983);
and U2997 (N_2997,In_158,In_1309);
nor U2998 (N_2998,In_269,In_841);
xor U2999 (N_2999,In_763,In_1903);
nor U3000 (N_3000,In_1329,In_209);
nand U3001 (N_3001,In_1704,In_1994);
xor U3002 (N_3002,In_459,In_723);
nand U3003 (N_3003,In_1147,In_257);
nand U3004 (N_3004,In_69,In_585);
xnor U3005 (N_3005,In_1317,In_861);
nand U3006 (N_3006,In_1788,In_891);
and U3007 (N_3007,In_789,In_6);
nor U3008 (N_3008,In_237,In_528);
or U3009 (N_3009,In_1407,In_1692);
nand U3010 (N_3010,In_1474,In_1452);
nor U3011 (N_3011,In_19,In_539);
xor U3012 (N_3012,In_87,In_1134);
nand U3013 (N_3013,In_1573,In_689);
nor U3014 (N_3014,In_1083,In_1410);
nand U3015 (N_3015,In_1313,In_1225);
or U3016 (N_3016,In_322,In_1570);
or U3017 (N_3017,In_847,In_144);
nand U3018 (N_3018,In_983,In_535);
or U3019 (N_3019,In_670,In_1017);
and U3020 (N_3020,In_425,In_286);
or U3021 (N_3021,In_535,In_1872);
nand U3022 (N_3022,In_1967,In_968);
or U3023 (N_3023,In_21,In_1522);
or U3024 (N_3024,In_1865,In_1463);
and U3025 (N_3025,In_887,In_1814);
and U3026 (N_3026,In_126,In_1953);
nand U3027 (N_3027,In_1023,In_266);
and U3028 (N_3028,In_1728,In_1230);
xnor U3029 (N_3029,In_174,In_377);
nor U3030 (N_3030,In_1267,In_901);
nand U3031 (N_3031,In_1863,In_1096);
nor U3032 (N_3032,In_781,In_1977);
or U3033 (N_3033,In_1615,In_908);
or U3034 (N_3034,In_350,In_980);
and U3035 (N_3035,In_1092,In_1830);
or U3036 (N_3036,In_1486,In_789);
nand U3037 (N_3037,In_1715,In_1906);
and U3038 (N_3038,In_1870,In_1108);
and U3039 (N_3039,In_990,In_1683);
xor U3040 (N_3040,In_1001,In_214);
nor U3041 (N_3041,In_1602,In_1590);
or U3042 (N_3042,In_1986,In_770);
and U3043 (N_3043,In_71,In_193);
and U3044 (N_3044,In_1756,In_402);
xnor U3045 (N_3045,In_596,In_1441);
and U3046 (N_3046,In_345,In_1042);
nor U3047 (N_3047,In_169,In_74);
nor U3048 (N_3048,In_516,In_1227);
nand U3049 (N_3049,In_1344,In_978);
nor U3050 (N_3050,In_1046,In_536);
and U3051 (N_3051,In_63,In_574);
xor U3052 (N_3052,In_1868,In_1085);
and U3053 (N_3053,In_1806,In_1461);
xnor U3054 (N_3054,In_404,In_1981);
xor U3055 (N_3055,In_1813,In_11);
xnor U3056 (N_3056,In_1450,In_1908);
nand U3057 (N_3057,In_686,In_3);
nor U3058 (N_3058,In_1289,In_1092);
xnor U3059 (N_3059,In_812,In_1159);
nand U3060 (N_3060,In_1839,In_244);
xnor U3061 (N_3061,In_1597,In_682);
and U3062 (N_3062,In_1352,In_202);
xor U3063 (N_3063,In_1992,In_1920);
xor U3064 (N_3064,In_1743,In_1626);
or U3065 (N_3065,In_777,In_1987);
nand U3066 (N_3066,In_1513,In_1742);
nor U3067 (N_3067,In_1491,In_1205);
and U3068 (N_3068,In_1470,In_103);
nor U3069 (N_3069,In_621,In_95);
xor U3070 (N_3070,In_1034,In_1801);
nor U3071 (N_3071,In_663,In_216);
and U3072 (N_3072,In_348,In_974);
xor U3073 (N_3073,In_1239,In_969);
nand U3074 (N_3074,In_1573,In_1838);
and U3075 (N_3075,In_1673,In_1962);
xnor U3076 (N_3076,In_49,In_1865);
nor U3077 (N_3077,In_128,In_1749);
nor U3078 (N_3078,In_1110,In_1555);
xor U3079 (N_3079,In_664,In_1504);
nand U3080 (N_3080,In_818,In_884);
or U3081 (N_3081,In_504,In_93);
xnor U3082 (N_3082,In_1323,In_1826);
and U3083 (N_3083,In_241,In_1029);
and U3084 (N_3084,In_1505,In_1452);
nand U3085 (N_3085,In_1055,In_723);
xnor U3086 (N_3086,In_114,In_1047);
nand U3087 (N_3087,In_608,In_1515);
and U3088 (N_3088,In_95,In_186);
nand U3089 (N_3089,In_239,In_1290);
and U3090 (N_3090,In_963,In_1728);
and U3091 (N_3091,In_1932,In_1150);
or U3092 (N_3092,In_1921,In_1832);
nor U3093 (N_3093,In_601,In_1651);
nand U3094 (N_3094,In_906,In_1989);
nor U3095 (N_3095,In_1909,In_655);
or U3096 (N_3096,In_483,In_905);
xnor U3097 (N_3097,In_1406,In_229);
or U3098 (N_3098,In_204,In_1811);
nand U3099 (N_3099,In_999,In_110);
and U3100 (N_3100,In_1680,In_454);
and U3101 (N_3101,In_1764,In_1398);
and U3102 (N_3102,In_1344,In_191);
xnor U3103 (N_3103,In_205,In_1738);
and U3104 (N_3104,In_725,In_972);
xor U3105 (N_3105,In_976,In_21);
and U3106 (N_3106,In_3,In_1162);
nand U3107 (N_3107,In_1648,In_493);
nand U3108 (N_3108,In_1142,In_108);
xor U3109 (N_3109,In_1197,In_1775);
nor U3110 (N_3110,In_1862,In_1571);
nand U3111 (N_3111,In_1793,In_1230);
and U3112 (N_3112,In_820,In_76);
nand U3113 (N_3113,In_1958,In_1858);
or U3114 (N_3114,In_817,In_374);
xor U3115 (N_3115,In_1638,In_89);
and U3116 (N_3116,In_1121,In_818);
nor U3117 (N_3117,In_865,In_1628);
and U3118 (N_3118,In_1031,In_985);
nand U3119 (N_3119,In_1244,In_902);
nor U3120 (N_3120,In_626,In_770);
and U3121 (N_3121,In_1285,In_1901);
nand U3122 (N_3122,In_287,In_1439);
xnor U3123 (N_3123,In_20,In_1089);
and U3124 (N_3124,In_423,In_1068);
nand U3125 (N_3125,In_533,In_1837);
xnor U3126 (N_3126,In_1000,In_1150);
xor U3127 (N_3127,In_1143,In_1083);
and U3128 (N_3128,In_1795,In_932);
nor U3129 (N_3129,In_1079,In_1526);
nand U3130 (N_3130,In_1582,In_603);
nand U3131 (N_3131,In_1186,In_1410);
and U3132 (N_3132,In_1800,In_1312);
xor U3133 (N_3133,In_1429,In_1793);
xor U3134 (N_3134,In_1250,In_1355);
or U3135 (N_3135,In_1135,In_943);
nand U3136 (N_3136,In_795,In_320);
nor U3137 (N_3137,In_755,In_658);
and U3138 (N_3138,In_993,In_1905);
or U3139 (N_3139,In_1540,In_692);
or U3140 (N_3140,In_1693,In_1021);
nand U3141 (N_3141,In_1746,In_950);
xnor U3142 (N_3142,In_1151,In_1059);
nand U3143 (N_3143,In_1328,In_1461);
nor U3144 (N_3144,In_23,In_1805);
xor U3145 (N_3145,In_1432,In_489);
and U3146 (N_3146,In_24,In_1082);
xnor U3147 (N_3147,In_728,In_1109);
nor U3148 (N_3148,In_1334,In_254);
nand U3149 (N_3149,In_1290,In_1408);
xnor U3150 (N_3150,In_1687,In_1191);
or U3151 (N_3151,In_164,In_853);
and U3152 (N_3152,In_1115,In_532);
xnor U3153 (N_3153,In_832,In_1023);
nor U3154 (N_3154,In_1381,In_1620);
nand U3155 (N_3155,In_1971,In_300);
or U3156 (N_3156,In_916,In_1892);
and U3157 (N_3157,In_1072,In_1040);
or U3158 (N_3158,In_1400,In_1349);
and U3159 (N_3159,In_33,In_1937);
nand U3160 (N_3160,In_737,In_715);
xnor U3161 (N_3161,In_1729,In_573);
xnor U3162 (N_3162,In_473,In_873);
or U3163 (N_3163,In_1130,In_1567);
xnor U3164 (N_3164,In_1242,In_650);
or U3165 (N_3165,In_1786,In_622);
and U3166 (N_3166,In_722,In_1328);
or U3167 (N_3167,In_680,In_1383);
nor U3168 (N_3168,In_77,In_552);
and U3169 (N_3169,In_788,In_1509);
xor U3170 (N_3170,In_521,In_1586);
nand U3171 (N_3171,In_418,In_8);
or U3172 (N_3172,In_1621,In_1195);
or U3173 (N_3173,In_1257,In_140);
and U3174 (N_3174,In_787,In_1479);
or U3175 (N_3175,In_1144,In_817);
nor U3176 (N_3176,In_599,In_1869);
nand U3177 (N_3177,In_916,In_1600);
nor U3178 (N_3178,In_1939,In_1050);
nor U3179 (N_3179,In_17,In_689);
xnor U3180 (N_3180,In_490,In_1291);
or U3181 (N_3181,In_1665,In_1491);
nand U3182 (N_3182,In_766,In_1814);
nand U3183 (N_3183,In_1765,In_1373);
xor U3184 (N_3184,In_490,In_846);
nor U3185 (N_3185,In_600,In_242);
xnor U3186 (N_3186,In_916,In_337);
or U3187 (N_3187,In_1111,In_840);
and U3188 (N_3188,In_1187,In_356);
and U3189 (N_3189,In_1752,In_1114);
xnor U3190 (N_3190,In_1073,In_1270);
or U3191 (N_3191,In_1934,In_207);
nand U3192 (N_3192,In_748,In_1673);
nor U3193 (N_3193,In_1874,In_128);
nor U3194 (N_3194,In_237,In_683);
or U3195 (N_3195,In_1153,In_1314);
or U3196 (N_3196,In_1631,In_1680);
and U3197 (N_3197,In_762,In_871);
and U3198 (N_3198,In_30,In_1390);
xnor U3199 (N_3199,In_1979,In_1779);
or U3200 (N_3200,In_1678,In_1742);
xnor U3201 (N_3201,In_1753,In_990);
xnor U3202 (N_3202,In_1771,In_686);
xnor U3203 (N_3203,In_51,In_24);
and U3204 (N_3204,In_1040,In_1466);
nand U3205 (N_3205,In_778,In_1483);
nor U3206 (N_3206,In_1393,In_487);
or U3207 (N_3207,In_1674,In_1642);
nand U3208 (N_3208,In_866,In_1133);
and U3209 (N_3209,In_775,In_1184);
nand U3210 (N_3210,In_793,In_1978);
or U3211 (N_3211,In_1972,In_392);
and U3212 (N_3212,In_523,In_1002);
nor U3213 (N_3213,In_147,In_72);
nand U3214 (N_3214,In_1390,In_1095);
and U3215 (N_3215,In_1334,In_1211);
nand U3216 (N_3216,In_1055,In_774);
xor U3217 (N_3217,In_1296,In_1150);
and U3218 (N_3218,In_517,In_234);
or U3219 (N_3219,In_529,In_1329);
or U3220 (N_3220,In_1947,In_1118);
and U3221 (N_3221,In_1505,In_1937);
nor U3222 (N_3222,In_1736,In_336);
xor U3223 (N_3223,In_915,In_1837);
nand U3224 (N_3224,In_515,In_187);
or U3225 (N_3225,In_1844,In_780);
nor U3226 (N_3226,In_975,In_1544);
and U3227 (N_3227,In_1039,In_1801);
nand U3228 (N_3228,In_873,In_724);
and U3229 (N_3229,In_1157,In_1293);
or U3230 (N_3230,In_1126,In_364);
or U3231 (N_3231,In_298,In_256);
xor U3232 (N_3232,In_1392,In_1919);
and U3233 (N_3233,In_1610,In_880);
xnor U3234 (N_3234,In_1577,In_835);
nand U3235 (N_3235,In_557,In_1637);
xnor U3236 (N_3236,In_197,In_1370);
or U3237 (N_3237,In_813,In_277);
and U3238 (N_3238,In_523,In_673);
or U3239 (N_3239,In_945,In_1991);
nand U3240 (N_3240,In_1790,In_553);
nand U3241 (N_3241,In_1341,In_1736);
nand U3242 (N_3242,In_559,In_1625);
xor U3243 (N_3243,In_1013,In_1612);
nor U3244 (N_3244,In_523,In_1695);
nor U3245 (N_3245,In_425,In_1518);
xnor U3246 (N_3246,In_370,In_77);
xor U3247 (N_3247,In_1050,In_773);
nor U3248 (N_3248,In_130,In_631);
or U3249 (N_3249,In_1858,In_640);
and U3250 (N_3250,In_298,In_79);
nor U3251 (N_3251,In_1422,In_1987);
or U3252 (N_3252,In_1859,In_735);
nand U3253 (N_3253,In_349,In_1292);
nand U3254 (N_3254,In_1817,In_767);
xor U3255 (N_3255,In_817,In_1112);
xor U3256 (N_3256,In_749,In_284);
nor U3257 (N_3257,In_197,In_534);
xor U3258 (N_3258,In_1955,In_501);
xnor U3259 (N_3259,In_793,In_1394);
and U3260 (N_3260,In_1632,In_799);
and U3261 (N_3261,In_1430,In_1777);
or U3262 (N_3262,In_1963,In_1130);
or U3263 (N_3263,In_1070,In_290);
and U3264 (N_3264,In_1156,In_856);
and U3265 (N_3265,In_221,In_992);
nand U3266 (N_3266,In_473,In_570);
nor U3267 (N_3267,In_1619,In_1061);
xnor U3268 (N_3268,In_1677,In_1560);
nor U3269 (N_3269,In_1513,In_710);
xor U3270 (N_3270,In_169,In_1408);
nand U3271 (N_3271,In_1255,In_1643);
or U3272 (N_3272,In_1181,In_467);
xnor U3273 (N_3273,In_691,In_1858);
nor U3274 (N_3274,In_1927,In_1190);
nor U3275 (N_3275,In_53,In_94);
xnor U3276 (N_3276,In_1682,In_1079);
or U3277 (N_3277,In_348,In_1967);
and U3278 (N_3278,In_1995,In_159);
nand U3279 (N_3279,In_1709,In_386);
and U3280 (N_3280,In_327,In_1317);
xnor U3281 (N_3281,In_1724,In_404);
or U3282 (N_3282,In_680,In_269);
nand U3283 (N_3283,In_1598,In_1488);
or U3284 (N_3284,In_1306,In_1787);
nand U3285 (N_3285,In_98,In_1617);
nor U3286 (N_3286,In_940,In_1294);
or U3287 (N_3287,In_462,In_861);
nor U3288 (N_3288,In_137,In_520);
nand U3289 (N_3289,In_319,In_1148);
xnor U3290 (N_3290,In_509,In_838);
and U3291 (N_3291,In_1160,In_1462);
or U3292 (N_3292,In_302,In_28);
nor U3293 (N_3293,In_641,In_941);
and U3294 (N_3294,In_54,In_325);
xnor U3295 (N_3295,In_448,In_1467);
xnor U3296 (N_3296,In_1393,In_384);
nand U3297 (N_3297,In_369,In_898);
and U3298 (N_3298,In_104,In_1322);
xnor U3299 (N_3299,In_398,In_898);
or U3300 (N_3300,In_46,In_1873);
or U3301 (N_3301,In_568,In_534);
and U3302 (N_3302,In_112,In_955);
and U3303 (N_3303,In_1172,In_1980);
nand U3304 (N_3304,In_1051,In_587);
or U3305 (N_3305,In_957,In_369);
or U3306 (N_3306,In_1699,In_541);
xor U3307 (N_3307,In_1374,In_88);
nand U3308 (N_3308,In_705,In_146);
xnor U3309 (N_3309,In_1561,In_1980);
and U3310 (N_3310,In_224,In_618);
nand U3311 (N_3311,In_588,In_573);
or U3312 (N_3312,In_1110,In_1848);
nor U3313 (N_3313,In_1939,In_653);
and U3314 (N_3314,In_1649,In_1235);
and U3315 (N_3315,In_1619,In_851);
and U3316 (N_3316,In_1447,In_877);
and U3317 (N_3317,In_181,In_716);
and U3318 (N_3318,In_1764,In_1996);
and U3319 (N_3319,In_1211,In_395);
or U3320 (N_3320,In_1049,In_1152);
xor U3321 (N_3321,In_1907,In_1487);
nand U3322 (N_3322,In_1855,In_248);
nor U3323 (N_3323,In_579,In_764);
or U3324 (N_3324,In_471,In_1743);
and U3325 (N_3325,In_1959,In_1180);
or U3326 (N_3326,In_1731,In_183);
xnor U3327 (N_3327,In_642,In_1553);
and U3328 (N_3328,In_1230,In_505);
nand U3329 (N_3329,In_1695,In_847);
nor U3330 (N_3330,In_261,In_915);
or U3331 (N_3331,In_1443,In_1131);
nand U3332 (N_3332,In_1857,In_1703);
or U3333 (N_3333,In_801,In_624);
nand U3334 (N_3334,In_1143,In_1536);
or U3335 (N_3335,In_646,In_1795);
nand U3336 (N_3336,In_206,In_51);
or U3337 (N_3337,In_1891,In_230);
xor U3338 (N_3338,In_827,In_1099);
nor U3339 (N_3339,In_404,In_543);
or U3340 (N_3340,In_1734,In_282);
or U3341 (N_3341,In_1884,In_36);
or U3342 (N_3342,In_280,In_1028);
or U3343 (N_3343,In_1264,In_333);
xnor U3344 (N_3344,In_905,In_1288);
or U3345 (N_3345,In_1238,In_370);
nand U3346 (N_3346,In_1983,In_1953);
nor U3347 (N_3347,In_615,In_1517);
nor U3348 (N_3348,In_1631,In_91);
and U3349 (N_3349,In_1299,In_1850);
nor U3350 (N_3350,In_268,In_1505);
xnor U3351 (N_3351,In_46,In_195);
nand U3352 (N_3352,In_1286,In_825);
or U3353 (N_3353,In_1342,In_1401);
nor U3354 (N_3354,In_175,In_287);
nor U3355 (N_3355,In_795,In_1330);
or U3356 (N_3356,In_1963,In_505);
xor U3357 (N_3357,In_29,In_1970);
and U3358 (N_3358,In_1184,In_93);
and U3359 (N_3359,In_466,In_1335);
nor U3360 (N_3360,In_411,In_556);
nor U3361 (N_3361,In_588,In_562);
xor U3362 (N_3362,In_814,In_1092);
and U3363 (N_3363,In_1762,In_1125);
or U3364 (N_3364,In_307,In_1941);
nor U3365 (N_3365,In_1895,In_428);
and U3366 (N_3366,In_825,In_1315);
xnor U3367 (N_3367,In_843,In_1575);
nand U3368 (N_3368,In_975,In_827);
nor U3369 (N_3369,In_288,In_746);
xnor U3370 (N_3370,In_820,In_1148);
nor U3371 (N_3371,In_716,In_619);
or U3372 (N_3372,In_281,In_236);
and U3373 (N_3373,In_124,In_1782);
and U3374 (N_3374,In_678,In_924);
or U3375 (N_3375,In_1594,In_987);
or U3376 (N_3376,In_1000,In_278);
or U3377 (N_3377,In_1766,In_1031);
nor U3378 (N_3378,In_468,In_1368);
and U3379 (N_3379,In_1866,In_351);
xor U3380 (N_3380,In_1825,In_11);
and U3381 (N_3381,In_1735,In_623);
and U3382 (N_3382,In_1984,In_1261);
xnor U3383 (N_3383,In_613,In_1308);
nand U3384 (N_3384,In_1329,In_254);
nand U3385 (N_3385,In_188,In_822);
xor U3386 (N_3386,In_365,In_1303);
nor U3387 (N_3387,In_1275,In_1056);
or U3388 (N_3388,In_838,In_1688);
and U3389 (N_3389,In_746,In_741);
xnor U3390 (N_3390,In_1394,In_1338);
xnor U3391 (N_3391,In_997,In_265);
or U3392 (N_3392,In_1273,In_593);
nand U3393 (N_3393,In_622,In_1218);
and U3394 (N_3394,In_1315,In_526);
or U3395 (N_3395,In_186,In_1104);
xnor U3396 (N_3396,In_317,In_35);
xor U3397 (N_3397,In_1580,In_1870);
nor U3398 (N_3398,In_1995,In_662);
and U3399 (N_3399,In_1015,In_1401);
xnor U3400 (N_3400,In_235,In_41);
nor U3401 (N_3401,In_407,In_778);
nor U3402 (N_3402,In_836,In_1476);
nand U3403 (N_3403,In_728,In_1498);
and U3404 (N_3404,In_1318,In_912);
xor U3405 (N_3405,In_1448,In_512);
and U3406 (N_3406,In_740,In_819);
nor U3407 (N_3407,In_1444,In_602);
nand U3408 (N_3408,In_424,In_1769);
nand U3409 (N_3409,In_165,In_500);
or U3410 (N_3410,In_1669,In_628);
nor U3411 (N_3411,In_411,In_1193);
nor U3412 (N_3412,In_313,In_1935);
xnor U3413 (N_3413,In_942,In_350);
xor U3414 (N_3414,In_410,In_1317);
xor U3415 (N_3415,In_42,In_1784);
xnor U3416 (N_3416,In_1501,In_151);
and U3417 (N_3417,In_1821,In_859);
or U3418 (N_3418,In_1072,In_1428);
xnor U3419 (N_3419,In_196,In_1687);
or U3420 (N_3420,In_1620,In_1883);
nor U3421 (N_3421,In_313,In_788);
nor U3422 (N_3422,In_1676,In_1414);
nand U3423 (N_3423,In_461,In_1509);
and U3424 (N_3424,In_1961,In_704);
and U3425 (N_3425,In_1772,In_1471);
or U3426 (N_3426,In_1995,In_1813);
nand U3427 (N_3427,In_1019,In_1641);
xnor U3428 (N_3428,In_1649,In_1341);
nand U3429 (N_3429,In_1101,In_1971);
and U3430 (N_3430,In_823,In_1420);
and U3431 (N_3431,In_461,In_761);
and U3432 (N_3432,In_61,In_156);
nand U3433 (N_3433,In_1500,In_1029);
or U3434 (N_3434,In_267,In_1898);
xor U3435 (N_3435,In_1986,In_62);
or U3436 (N_3436,In_1214,In_1690);
nand U3437 (N_3437,In_1279,In_1045);
nand U3438 (N_3438,In_1296,In_71);
nand U3439 (N_3439,In_1184,In_1772);
nand U3440 (N_3440,In_1213,In_553);
or U3441 (N_3441,In_1211,In_1090);
nor U3442 (N_3442,In_812,In_1247);
nand U3443 (N_3443,In_1420,In_53);
xnor U3444 (N_3444,In_42,In_546);
or U3445 (N_3445,In_482,In_1217);
nor U3446 (N_3446,In_1110,In_1623);
or U3447 (N_3447,In_674,In_1682);
and U3448 (N_3448,In_1132,In_112);
xor U3449 (N_3449,In_1352,In_74);
or U3450 (N_3450,In_1443,In_994);
xor U3451 (N_3451,In_1031,In_1575);
nor U3452 (N_3452,In_223,In_877);
nand U3453 (N_3453,In_125,In_1442);
nor U3454 (N_3454,In_88,In_827);
nor U3455 (N_3455,In_1082,In_536);
nand U3456 (N_3456,In_698,In_901);
and U3457 (N_3457,In_755,In_915);
and U3458 (N_3458,In_151,In_512);
or U3459 (N_3459,In_1193,In_389);
or U3460 (N_3460,In_818,In_403);
or U3461 (N_3461,In_932,In_1249);
nand U3462 (N_3462,In_470,In_11);
nor U3463 (N_3463,In_1707,In_1799);
or U3464 (N_3464,In_920,In_1366);
nor U3465 (N_3465,In_1377,In_1814);
or U3466 (N_3466,In_553,In_425);
nand U3467 (N_3467,In_1991,In_51);
or U3468 (N_3468,In_1500,In_850);
and U3469 (N_3469,In_1835,In_599);
nand U3470 (N_3470,In_1046,In_407);
xor U3471 (N_3471,In_315,In_253);
nand U3472 (N_3472,In_552,In_1357);
or U3473 (N_3473,In_386,In_1949);
or U3474 (N_3474,In_9,In_872);
or U3475 (N_3475,In_535,In_480);
nand U3476 (N_3476,In_1774,In_935);
and U3477 (N_3477,In_454,In_21);
and U3478 (N_3478,In_1759,In_1214);
and U3479 (N_3479,In_1307,In_1429);
or U3480 (N_3480,In_288,In_1748);
xor U3481 (N_3481,In_1079,In_267);
and U3482 (N_3482,In_1605,In_1693);
xor U3483 (N_3483,In_393,In_625);
nor U3484 (N_3484,In_1746,In_1837);
and U3485 (N_3485,In_1946,In_1408);
nor U3486 (N_3486,In_1207,In_165);
and U3487 (N_3487,In_134,In_504);
or U3488 (N_3488,In_824,In_1372);
or U3489 (N_3489,In_947,In_412);
nor U3490 (N_3490,In_600,In_1464);
xor U3491 (N_3491,In_1667,In_1400);
and U3492 (N_3492,In_1789,In_1165);
xnor U3493 (N_3493,In_724,In_616);
or U3494 (N_3494,In_1303,In_1871);
nor U3495 (N_3495,In_46,In_455);
and U3496 (N_3496,In_880,In_1326);
or U3497 (N_3497,In_827,In_1583);
or U3498 (N_3498,In_1692,In_399);
and U3499 (N_3499,In_169,In_1153);
nor U3500 (N_3500,In_1178,In_1261);
nor U3501 (N_3501,In_226,In_1763);
nor U3502 (N_3502,In_1443,In_544);
and U3503 (N_3503,In_1446,In_134);
xor U3504 (N_3504,In_1787,In_1224);
nand U3505 (N_3505,In_432,In_825);
or U3506 (N_3506,In_828,In_683);
nand U3507 (N_3507,In_913,In_1309);
or U3508 (N_3508,In_1263,In_773);
or U3509 (N_3509,In_999,In_1714);
or U3510 (N_3510,In_692,In_1655);
and U3511 (N_3511,In_1110,In_1058);
nor U3512 (N_3512,In_314,In_85);
xor U3513 (N_3513,In_85,In_1637);
and U3514 (N_3514,In_538,In_810);
and U3515 (N_3515,In_520,In_232);
nand U3516 (N_3516,In_1217,In_1502);
xnor U3517 (N_3517,In_1933,In_1953);
or U3518 (N_3518,In_1917,In_445);
nand U3519 (N_3519,In_1405,In_199);
xor U3520 (N_3520,In_1396,In_1714);
and U3521 (N_3521,In_1310,In_279);
nor U3522 (N_3522,In_1611,In_1869);
nand U3523 (N_3523,In_1856,In_1167);
nor U3524 (N_3524,In_1133,In_553);
and U3525 (N_3525,In_1488,In_766);
nand U3526 (N_3526,In_1910,In_805);
or U3527 (N_3527,In_1911,In_1225);
nor U3528 (N_3528,In_1160,In_1368);
nand U3529 (N_3529,In_750,In_1553);
nand U3530 (N_3530,In_1165,In_429);
and U3531 (N_3531,In_1189,In_1968);
or U3532 (N_3532,In_1032,In_773);
nand U3533 (N_3533,In_126,In_1983);
nand U3534 (N_3534,In_405,In_880);
nand U3535 (N_3535,In_1950,In_54);
and U3536 (N_3536,In_302,In_568);
xnor U3537 (N_3537,In_658,In_1421);
nor U3538 (N_3538,In_751,In_966);
nand U3539 (N_3539,In_801,In_48);
xnor U3540 (N_3540,In_802,In_558);
nor U3541 (N_3541,In_302,In_1283);
and U3542 (N_3542,In_1160,In_1394);
nand U3543 (N_3543,In_648,In_164);
nand U3544 (N_3544,In_1059,In_939);
nor U3545 (N_3545,In_1452,In_1248);
nor U3546 (N_3546,In_1371,In_1295);
or U3547 (N_3547,In_104,In_1446);
xnor U3548 (N_3548,In_1159,In_259);
xor U3549 (N_3549,In_1519,In_95);
nand U3550 (N_3550,In_1243,In_705);
nand U3551 (N_3551,In_1349,In_579);
nor U3552 (N_3552,In_331,In_1500);
xnor U3553 (N_3553,In_315,In_1379);
or U3554 (N_3554,In_1716,In_992);
or U3555 (N_3555,In_1060,In_991);
nand U3556 (N_3556,In_674,In_1539);
xor U3557 (N_3557,In_519,In_1173);
and U3558 (N_3558,In_1847,In_649);
nor U3559 (N_3559,In_1290,In_1088);
nor U3560 (N_3560,In_1701,In_1025);
and U3561 (N_3561,In_1173,In_1281);
xor U3562 (N_3562,In_169,In_1714);
nand U3563 (N_3563,In_944,In_1519);
xnor U3564 (N_3564,In_1628,In_1060);
or U3565 (N_3565,In_315,In_1130);
nand U3566 (N_3566,In_1236,In_961);
and U3567 (N_3567,In_1910,In_1009);
or U3568 (N_3568,In_1969,In_637);
nor U3569 (N_3569,In_1041,In_914);
nand U3570 (N_3570,In_1671,In_1338);
nand U3571 (N_3571,In_69,In_1822);
xnor U3572 (N_3572,In_1912,In_1558);
nor U3573 (N_3573,In_537,In_1750);
or U3574 (N_3574,In_314,In_833);
nor U3575 (N_3575,In_1432,In_1805);
and U3576 (N_3576,In_972,In_1605);
nor U3577 (N_3577,In_1699,In_60);
nor U3578 (N_3578,In_471,In_630);
nand U3579 (N_3579,In_770,In_1740);
and U3580 (N_3580,In_1661,In_62);
nand U3581 (N_3581,In_1444,In_1684);
nor U3582 (N_3582,In_175,In_598);
xor U3583 (N_3583,In_0,In_151);
xnor U3584 (N_3584,In_462,In_1030);
xor U3585 (N_3585,In_1284,In_1089);
and U3586 (N_3586,In_300,In_1093);
xnor U3587 (N_3587,In_69,In_83);
nor U3588 (N_3588,In_418,In_902);
or U3589 (N_3589,In_1438,In_1737);
nor U3590 (N_3590,In_1124,In_944);
and U3591 (N_3591,In_957,In_107);
xnor U3592 (N_3592,In_1299,In_1656);
nor U3593 (N_3593,In_699,In_1483);
or U3594 (N_3594,In_395,In_222);
nor U3595 (N_3595,In_5,In_716);
nand U3596 (N_3596,In_1389,In_1447);
nand U3597 (N_3597,In_1814,In_1871);
or U3598 (N_3598,In_175,In_721);
or U3599 (N_3599,In_1697,In_1538);
xor U3600 (N_3600,In_1839,In_455);
xnor U3601 (N_3601,In_1586,In_1980);
and U3602 (N_3602,In_205,In_1434);
and U3603 (N_3603,In_476,In_739);
or U3604 (N_3604,In_613,In_85);
and U3605 (N_3605,In_100,In_1170);
and U3606 (N_3606,In_275,In_1659);
nand U3607 (N_3607,In_1379,In_1270);
nand U3608 (N_3608,In_223,In_395);
xor U3609 (N_3609,In_834,In_872);
xnor U3610 (N_3610,In_43,In_387);
or U3611 (N_3611,In_981,In_1655);
nand U3612 (N_3612,In_116,In_203);
nor U3613 (N_3613,In_1563,In_1967);
or U3614 (N_3614,In_1028,In_426);
or U3615 (N_3615,In_866,In_973);
nand U3616 (N_3616,In_86,In_1417);
xnor U3617 (N_3617,In_636,In_1991);
or U3618 (N_3618,In_1238,In_1944);
or U3619 (N_3619,In_641,In_783);
or U3620 (N_3620,In_1198,In_1110);
and U3621 (N_3621,In_1002,In_1176);
and U3622 (N_3622,In_377,In_432);
and U3623 (N_3623,In_243,In_1713);
nor U3624 (N_3624,In_16,In_1284);
and U3625 (N_3625,In_670,In_749);
nor U3626 (N_3626,In_1899,In_491);
xor U3627 (N_3627,In_1315,In_1926);
nand U3628 (N_3628,In_1637,In_1449);
and U3629 (N_3629,In_1942,In_562);
nand U3630 (N_3630,In_115,In_606);
or U3631 (N_3631,In_338,In_1174);
or U3632 (N_3632,In_1317,In_258);
and U3633 (N_3633,In_1836,In_521);
nor U3634 (N_3634,In_445,In_1617);
or U3635 (N_3635,In_1286,In_657);
xor U3636 (N_3636,In_1278,In_1525);
and U3637 (N_3637,In_1790,In_1571);
nor U3638 (N_3638,In_1911,In_1866);
nand U3639 (N_3639,In_1462,In_834);
nand U3640 (N_3640,In_1317,In_1233);
nor U3641 (N_3641,In_1946,In_1084);
nor U3642 (N_3642,In_1145,In_118);
and U3643 (N_3643,In_110,In_131);
and U3644 (N_3644,In_420,In_930);
and U3645 (N_3645,In_1234,In_1354);
or U3646 (N_3646,In_1767,In_428);
and U3647 (N_3647,In_803,In_885);
nand U3648 (N_3648,In_1120,In_1340);
or U3649 (N_3649,In_978,In_1239);
nor U3650 (N_3650,In_15,In_718);
and U3651 (N_3651,In_342,In_678);
and U3652 (N_3652,In_232,In_484);
nor U3653 (N_3653,In_457,In_1462);
and U3654 (N_3654,In_490,In_153);
or U3655 (N_3655,In_921,In_117);
or U3656 (N_3656,In_1539,In_1885);
or U3657 (N_3657,In_464,In_1777);
or U3658 (N_3658,In_1651,In_1265);
nand U3659 (N_3659,In_1104,In_1525);
nand U3660 (N_3660,In_100,In_1420);
nor U3661 (N_3661,In_434,In_401);
nand U3662 (N_3662,In_709,In_1045);
nand U3663 (N_3663,In_1805,In_477);
nand U3664 (N_3664,In_258,In_342);
nand U3665 (N_3665,In_613,In_27);
xnor U3666 (N_3666,In_513,In_726);
nand U3667 (N_3667,In_876,In_932);
and U3668 (N_3668,In_1123,In_1609);
or U3669 (N_3669,In_6,In_1272);
and U3670 (N_3670,In_1648,In_1645);
or U3671 (N_3671,In_656,In_755);
xor U3672 (N_3672,In_709,In_544);
and U3673 (N_3673,In_870,In_1971);
xor U3674 (N_3674,In_1517,In_1073);
or U3675 (N_3675,In_1616,In_1894);
and U3676 (N_3676,In_1829,In_1125);
xor U3677 (N_3677,In_1810,In_1687);
or U3678 (N_3678,In_1363,In_1219);
or U3679 (N_3679,In_1162,In_506);
and U3680 (N_3680,In_795,In_1333);
xor U3681 (N_3681,In_1571,In_939);
nor U3682 (N_3682,In_596,In_674);
or U3683 (N_3683,In_276,In_1693);
xor U3684 (N_3684,In_1954,In_1695);
nor U3685 (N_3685,In_1385,In_334);
nand U3686 (N_3686,In_730,In_317);
and U3687 (N_3687,In_413,In_1482);
xnor U3688 (N_3688,In_1079,In_145);
or U3689 (N_3689,In_584,In_1274);
xor U3690 (N_3690,In_663,In_41);
nand U3691 (N_3691,In_1751,In_797);
or U3692 (N_3692,In_1858,In_1407);
nand U3693 (N_3693,In_531,In_1805);
nand U3694 (N_3694,In_897,In_29);
and U3695 (N_3695,In_1627,In_294);
nor U3696 (N_3696,In_1578,In_1966);
nor U3697 (N_3697,In_613,In_1217);
nand U3698 (N_3698,In_206,In_1938);
or U3699 (N_3699,In_1319,In_559);
xor U3700 (N_3700,In_1237,In_680);
nand U3701 (N_3701,In_1657,In_1845);
nor U3702 (N_3702,In_318,In_1117);
and U3703 (N_3703,In_1965,In_992);
xor U3704 (N_3704,In_311,In_1294);
nand U3705 (N_3705,In_1359,In_1321);
and U3706 (N_3706,In_1245,In_1496);
nor U3707 (N_3707,In_1412,In_850);
and U3708 (N_3708,In_1947,In_948);
nor U3709 (N_3709,In_1487,In_879);
and U3710 (N_3710,In_1003,In_102);
nand U3711 (N_3711,In_1388,In_695);
nand U3712 (N_3712,In_766,In_1208);
xor U3713 (N_3713,In_18,In_970);
nand U3714 (N_3714,In_1250,In_733);
xor U3715 (N_3715,In_199,In_1832);
xor U3716 (N_3716,In_1536,In_681);
nor U3717 (N_3717,In_1632,In_1743);
nand U3718 (N_3718,In_966,In_770);
nand U3719 (N_3719,In_1125,In_199);
nand U3720 (N_3720,In_1225,In_60);
nand U3721 (N_3721,In_1321,In_1432);
or U3722 (N_3722,In_612,In_19);
xor U3723 (N_3723,In_1703,In_84);
xor U3724 (N_3724,In_1258,In_1860);
and U3725 (N_3725,In_304,In_1719);
or U3726 (N_3726,In_1408,In_484);
or U3727 (N_3727,In_144,In_1226);
nand U3728 (N_3728,In_1209,In_335);
nand U3729 (N_3729,In_1283,In_608);
nor U3730 (N_3730,In_1336,In_780);
xor U3731 (N_3731,In_1472,In_1623);
nor U3732 (N_3732,In_980,In_115);
xor U3733 (N_3733,In_1290,In_254);
or U3734 (N_3734,In_396,In_1969);
or U3735 (N_3735,In_1792,In_730);
nor U3736 (N_3736,In_1113,In_1578);
or U3737 (N_3737,In_27,In_1779);
nand U3738 (N_3738,In_113,In_1614);
nand U3739 (N_3739,In_953,In_215);
or U3740 (N_3740,In_565,In_1606);
nor U3741 (N_3741,In_1193,In_206);
nor U3742 (N_3742,In_1565,In_151);
or U3743 (N_3743,In_596,In_1579);
or U3744 (N_3744,In_1021,In_332);
and U3745 (N_3745,In_1251,In_931);
xnor U3746 (N_3746,In_379,In_1456);
nand U3747 (N_3747,In_1409,In_908);
nor U3748 (N_3748,In_283,In_1749);
and U3749 (N_3749,In_740,In_233);
or U3750 (N_3750,In_127,In_1702);
and U3751 (N_3751,In_567,In_1648);
and U3752 (N_3752,In_296,In_1088);
and U3753 (N_3753,In_1828,In_77);
nand U3754 (N_3754,In_1253,In_559);
xnor U3755 (N_3755,In_1844,In_278);
nor U3756 (N_3756,In_847,In_159);
nand U3757 (N_3757,In_1595,In_1576);
and U3758 (N_3758,In_1069,In_752);
and U3759 (N_3759,In_1358,In_325);
or U3760 (N_3760,In_1766,In_1944);
nor U3761 (N_3761,In_1739,In_1445);
nand U3762 (N_3762,In_868,In_690);
nor U3763 (N_3763,In_1403,In_275);
or U3764 (N_3764,In_827,In_3);
nor U3765 (N_3765,In_1135,In_1445);
xor U3766 (N_3766,In_394,In_1143);
xor U3767 (N_3767,In_1640,In_1765);
or U3768 (N_3768,In_536,In_1216);
nand U3769 (N_3769,In_422,In_1341);
xor U3770 (N_3770,In_963,In_527);
and U3771 (N_3771,In_453,In_33);
xor U3772 (N_3772,In_129,In_275);
xor U3773 (N_3773,In_767,In_1151);
nor U3774 (N_3774,In_854,In_1113);
and U3775 (N_3775,In_1575,In_913);
nor U3776 (N_3776,In_889,In_1526);
nand U3777 (N_3777,In_1743,In_113);
xnor U3778 (N_3778,In_561,In_545);
or U3779 (N_3779,In_999,In_1113);
and U3780 (N_3780,In_1385,In_354);
nand U3781 (N_3781,In_1536,In_1728);
nand U3782 (N_3782,In_585,In_1963);
nand U3783 (N_3783,In_105,In_1455);
nand U3784 (N_3784,In_85,In_75);
and U3785 (N_3785,In_886,In_1007);
or U3786 (N_3786,In_475,In_1837);
nand U3787 (N_3787,In_1932,In_43);
or U3788 (N_3788,In_223,In_1996);
and U3789 (N_3789,In_1440,In_1988);
xnor U3790 (N_3790,In_1831,In_1038);
and U3791 (N_3791,In_191,In_1880);
or U3792 (N_3792,In_73,In_4);
nand U3793 (N_3793,In_1858,In_1937);
nor U3794 (N_3794,In_823,In_1911);
or U3795 (N_3795,In_443,In_1170);
nor U3796 (N_3796,In_74,In_822);
nor U3797 (N_3797,In_1255,In_803);
nor U3798 (N_3798,In_1271,In_992);
nor U3799 (N_3799,In_1558,In_1149);
xor U3800 (N_3800,In_1326,In_1545);
nor U3801 (N_3801,In_1744,In_1405);
and U3802 (N_3802,In_1528,In_1374);
or U3803 (N_3803,In_56,In_1620);
or U3804 (N_3804,In_1699,In_1860);
nor U3805 (N_3805,In_394,In_1417);
or U3806 (N_3806,In_1183,In_1801);
or U3807 (N_3807,In_965,In_1460);
xor U3808 (N_3808,In_412,In_1531);
nor U3809 (N_3809,In_1038,In_969);
nand U3810 (N_3810,In_1120,In_635);
and U3811 (N_3811,In_900,In_399);
or U3812 (N_3812,In_478,In_89);
or U3813 (N_3813,In_1519,In_300);
nand U3814 (N_3814,In_1728,In_387);
or U3815 (N_3815,In_1509,In_1732);
and U3816 (N_3816,In_944,In_1192);
nand U3817 (N_3817,In_1829,In_1586);
xor U3818 (N_3818,In_1114,In_1932);
xnor U3819 (N_3819,In_1752,In_338);
nor U3820 (N_3820,In_1698,In_1634);
xnor U3821 (N_3821,In_738,In_1591);
and U3822 (N_3822,In_352,In_1259);
nand U3823 (N_3823,In_288,In_1379);
or U3824 (N_3824,In_1169,In_1091);
nand U3825 (N_3825,In_151,In_269);
or U3826 (N_3826,In_1023,In_51);
nor U3827 (N_3827,In_1516,In_1855);
xor U3828 (N_3828,In_209,In_577);
nor U3829 (N_3829,In_1437,In_832);
nor U3830 (N_3830,In_197,In_782);
nor U3831 (N_3831,In_1910,In_1648);
nor U3832 (N_3832,In_294,In_1228);
xnor U3833 (N_3833,In_1433,In_1505);
or U3834 (N_3834,In_515,In_146);
nor U3835 (N_3835,In_180,In_1461);
nand U3836 (N_3836,In_1229,In_939);
and U3837 (N_3837,In_401,In_1186);
nor U3838 (N_3838,In_1600,In_747);
or U3839 (N_3839,In_1308,In_1142);
nor U3840 (N_3840,In_1052,In_471);
or U3841 (N_3841,In_1737,In_1471);
nor U3842 (N_3842,In_1165,In_773);
or U3843 (N_3843,In_873,In_519);
or U3844 (N_3844,In_1023,In_1631);
or U3845 (N_3845,In_1243,In_497);
nand U3846 (N_3846,In_1922,In_398);
or U3847 (N_3847,In_967,In_425);
nand U3848 (N_3848,In_1517,In_924);
nor U3849 (N_3849,In_1263,In_1747);
or U3850 (N_3850,In_570,In_992);
and U3851 (N_3851,In_896,In_1159);
and U3852 (N_3852,In_876,In_1517);
xor U3853 (N_3853,In_1139,In_409);
nand U3854 (N_3854,In_354,In_1208);
nand U3855 (N_3855,In_287,In_1725);
and U3856 (N_3856,In_381,In_907);
or U3857 (N_3857,In_80,In_1380);
or U3858 (N_3858,In_936,In_1790);
and U3859 (N_3859,In_626,In_1089);
and U3860 (N_3860,In_1766,In_1255);
nor U3861 (N_3861,In_1048,In_447);
nand U3862 (N_3862,In_812,In_1679);
and U3863 (N_3863,In_1031,In_1314);
and U3864 (N_3864,In_406,In_1443);
nand U3865 (N_3865,In_1811,In_1682);
nor U3866 (N_3866,In_924,In_488);
nand U3867 (N_3867,In_1669,In_877);
nor U3868 (N_3868,In_1051,In_1381);
or U3869 (N_3869,In_1508,In_920);
and U3870 (N_3870,In_670,In_559);
xnor U3871 (N_3871,In_405,In_798);
nand U3872 (N_3872,In_1266,In_542);
xnor U3873 (N_3873,In_1231,In_1843);
xor U3874 (N_3874,In_232,In_218);
and U3875 (N_3875,In_1353,In_1450);
or U3876 (N_3876,In_1374,In_1285);
or U3877 (N_3877,In_1258,In_1927);
nand U3878 (N_3878,In_373,In_268);
nor U3879 (N_3879,In_914,In_261);
and U3880 (N_3880,In_141,In_1685);
xor U3881 (N_3881,In_620,In_1346);
or U3882 (N_3882,In_93,In_7);
or U3883 (N_3883,In_1755,In_264);
nand U3884 (N_3884,In_946,In_1204);
nor U3885 (N_3885,In_373,In_464);
nand U3886 (N_3886,In_588,In_279);
xor U3887 (N_3887,In_655,In_1606);
or U3888 (N_3888,In_896,In_289);
and U3889 (N_3889,In_885,In_1051);
or U3890 (N_3890,In_808,In_387);
nand U3891 (N_3891,In_417,In_654);
and U3892 (N_3892,In_165,In_1347);
xor U3893 (N_3893,In_1023,In_555);
and U3894 (N_3894,In_335,In_1650);
nor U3895 (N_3895,In_261,In_97);
nor U3896 (N_3896,In_1967,In_29);
xnor U3897 (N_3897,In_1991,In_736);
xor U3898 (N_3898,In_617,In_903);
nand U3899 (N_3899,In_600,In_1383);
nand U3900 (N_3900,In_231,In_1747);
xnor U3901 (N_3901,In_733,In_230);
xor U3902 (N_3902,In_1445,In_1363);
and U3903 (N_3903,In_550,In_1972);
or U3904 (N_3904,In_1575,In_471);
or U3905 (N_3905,In_1172,In_76);
xnor U3906 (N_3906,In_1460,In_1726);
xor U3907 (N_3907,In_1035,In_339);
nor U3908 (N_3908,In_1700,In_427);
nor U3909 (N_3909,In_793,In_1449);
nor U3910 (N_3910,In_111,In_1762);
xor U3911 (N_3911,In_1207,In_1329);
or U3912 (N_3912,In_1108,In_844);
xor U3913 (N_3913,In_128,In_1016);
or U3914 (N_3914,In_1775,In_869);
or U3915 (N_3915,In_1059,In_772);
xor U3916 (N_3916,In_1181,In_689);
nand U3917 (N_3917,In_441,In_141);
xnor U3918 (N_3918,In_496,In_488);
xor U3919 (N_3919,In_1244,In_110);
and U3920 (N_3920,In_579,In_308);
or U3921 (N_3921,In_1066,In_543);
nor U3922 (N_3922,In_1093,In_209);
xor U3923 (N_3923,In_142,In_1780);
and U3924 (N_3924,In_1413,In_1335);
nand U3925 (N_3925,In_1669,In_992);
or U3926 (N_3926,In_821,In_695);
and U3927 (N_3927,In_1634,In_1423);
nand U3928 (N_3928,In_1851,In_668);
nand U3929 (N_3929,In_724,In_773);
or U3930 (N_3930,In_873,In_1081);
xnor U3931 (N_3931,In_1917,In_1835);
nand U3932 (N_3932,In_274,In_890);
or U3933 (N_3933,In_242,In_1394);
nand U3934 (N_3934,In_338,In_265);
nand U3935 (N_3935,In_28,In_786);
nor U3936 (N_3936,In_1632,In_1376);
or U3937 (N_3937,In_924,In_1867);
or U3938 (N_3938,In_839,In_1160);
or U3939 (N_3939,In_371,In_1535);
nand U3940 (N_3940,In_844,In_1343);
nor U3941 (N_3941,In_444,In_1704);
or U3942 (N_3942,In_488,In_1265);
and U3943 (N_3943,In_812,In_189);
or U3944 (N_3944,In_21,In_507);
nand U3945 (N_3945,In_942,In_928);
xor U3946 (N_3946,In_195,In_285);
nor U3947 (N_3947,In_649,In_1814);
nor U3948 (N_3948,In_1860,In_995);
and U3949 (N_3949,In_1970,In_1446);
or U3950 (N_3950,In_142,In_1822);
and U3951 (N_3951,In_1713,In_1272);
nand U3952 (N_3952,In_740,In_89);
nand U3953 (N_3953,In_1899,In_1745);
and U3954 (N_3954,In_222,In_679);
or U3955 (N_3955,In_1681,In_9);
xor U3956 (N_3956,In_1218,In_131);
or U3957 (N_3957,In_606,In_247);
xor U3958 (N_3958,In_1353,In_1557);
nor U3959 (N_3959,In_947,In_886);
nand U3960 (N_3960,In_157,In_1281);
and U3961 (N_3961,In_801,In_1062);
nor U3962 (N_3962,In_1047,In_1149);
and U3963 (N_3963,In_1515,In_1265);
xnor U3964 (N_3964,In_1280,In_1549);
nor U3965 (N_3965,In_537,In_1738);
or U3966 (N_3966,In_677,In_1989);
and U3967 (N_3967,In_1680,In_1411);
xnor U3968 (N_3968,In_1780,In_600);
or U3969 (N_3969,In_1897,In_1997);
nor U3970 (N_3970,In_1719,In_1435);
or U3971 (N_3971,In_1252,In_1702);
or U3972 (N_3972,In_573,In_1847);
and U3973 (N_3973,In_801,In_1161);
nand U3974 (N_3974,In_908,In_905);
or U3975 (N_3975,In_260,In_987);
nand U3976 (N_3976,In_1862,In_1296);
nand U3977 (N_3977,In_1338,In_780);
nor U3978 (N_3978,In_1587,In_1733);
xor U3979 (N_3979,In_220,In_1916);
or U3980 (N_3980,In_1259,In_1498);
or U3981 (N_3981,In_422,In_403);
nand U3982 (N_3982,In_51,In_451);
xor U3983 (N_3983,In_1493,In_1284);
nand U3984 (N_3984,In_962,In_611);
xnor U3985 (N_3985,In_687,In_1373);
and U3986 (N_3986,In_1593,In_1461);
nor U3987 (N_3987,In_1572,In_1491);
nand U3988 (N_3988,In_1784,In_382);
and U3989 (N_3989,In_1209,In_1227);
nand U3990 (N_3990,In_1646,In_591);
nor U3991 (N_3991,In_422,In_242);
nor U3992 (N_3992,In_1430,In_458);
or U3993 (N_3993,In_575,In_697);
nor U3994 (N_3994,In_346,In_1153);
xnor U3995 (N_3995,In_244,In_1172);
and U3996 (N_3996,In_1724,In_1511);
and U3997 (N_3997,In_545,In_1133);
nor U3998 (N_3998,In_1083,In_1998);
nand U3999 (N_3999,In_1815,In_1875);
and U4000 (N_4000,N_2046,N_3202);
nand U4001 (N_4001,N_770,N_3598);
xnor U4002 (N_4002,N_1698,N_3137);
xor U4003 (N_4003,N_3778,N_298);
nand U4004 (N_4004,N_3392,N_1821);
xnor U4005 (N_4005,N_419,N_1769);
nand U4006 (N_4006,N_3053,N_3200);
nand U4007 (N_4007,N_3352,N_923);
nand U4008 (N_4008,N_1619,N_1621);
or U4009 (N_4009,N_3817,N_228);
nand U4010 (N_4010,N_807,N_728);
and U4011 (N_4011,N_1606,N_37);
and U4012 (N_4012,N_992,N_1797);
xor U4013 (N_4013,N_2480,N_9);
or U4014 (N_4014,N_3286,N_3579);
nor U4015 (N_4015,N_945,N_3015);
nand U4016 (N_4016,N_3561,N_3198);
xor U4017 (N_4017,N_2958,N_2922);
xor U4018 (N_4018,N_237,N_3270);
xnor U4019 (N_4019,N_638,N_3495);
nand U4020 (N_4020,N_3390,N_2780);
and U4021 (N_4021,N_69,N_2696);
xnor U4022 (N_4022,N_3965,N_3010);
nand U4023 (N_4023,N_1939,N_2019);
xor U4024 (N_4024,N_1135,N_3224);
nor U4025 (N_4025,N_3570,N_959);
nor U4026 (N_4026,N_1720,N_2106);
xor U4027 (N_4027,N_1782,N_3100);
xnor U4028 (N_4028,N_2527,N_304);
or U4029 (N_4029,N_2458,N_2886);
xnor U4030 (N_4030,N_1214,N_2490);
and U4031 (N_4031,N_3321,N_1902);
xnor U4032 (N_4032,N_2836,N_3958);
nand U4033 (N_4033,N_1272,N_825);
nand U4034 (N_4034,N_3109,N_3765);
or U4035 (N_4035,N_2436,N_3768);
and U4036 (N_4036,N_198,N_649);
xor U4037 (N_4037,N_1943,N_3758);
or U4038 (N_4038,N_2028,N_197);
and U4039 (N_4039,N_3003,N_2113);
nor U4040 (N_4040,N_3948,N_2277);
or U4041 (N_4041,N_2292,N_1058);
or U4042 (N_4042,N_3252,N_3411);
nor U4043 (N_4043,N_173,N_35);
and U4044 (N_4044,N_3833,N_3050);
nor U4045 (N_4045,N_3950,N_312);
nor U4046 (N_4046,N_1642,N_1008);
or U4047 (N_4047,N_1830,N_2086);
xnor U4048 (N_4048,N_2718,N_3464);
or U4049 (N_4049,N_2099,N_1278);
nor U4050 (N_4050,N_3282,N_1450);
or U4051 (N_4051,N_518,N_2395);
or U4052 (N_4052,N_3344,N_1504);
xor U4053 (N_4053,N_915,N_1861);
xor U4054 (N_4054,N_3697,N_2469);
nor U4055 (N_4055,N_3964,N_365);
and U4056 (N_4056,N_3077,N_2830);
nor U4057 (N_4057,N_1670,N_3361);
nor U4058 (N_4058,N_405,N_3215);
nor U4059 (N_4059,N_3481,N_2342);
nor U4060 (N_4060,N_2363,N_3770);
nand U4061 (N_4061,N_804,N_1481);
nand U4062 (N_4062,N_3438,N_2392);
xor U4063 (N_4063,N_495,N_3811);
nor U4064 (N_4064,N_2597,N_3025);
nor U4065 (N_4065,N_508,N_700);
xor U4066 (N_4066,N_307,N_596);
and U4067 (N_4067,N_1182,N_835);
nand U4068 (N_4068,N_2297,N_3850);
xnor U4069 (N_4069,N_1100,N_3550);
or U4070 (N_4070,N_3514,N_3253);
nor U4071 (N_4071,N_347,N_1498);
nand U4072 (N_4072,N_3216,N_2984);
or U4073 (N_4073,N_824,N_1665);
nand U4074 (N_4074,N_3158,N_3991);
nand U4075 (N_4075,N_3276,N_633);
nand U4076 (N_4076,N_2837,N_3132);
and U4077 (N_4077,N_1890,N_1886);
nor U4078 (N_4078,N_3445,N_366);
nor U4079 (N_4079,N_3803,N_568);
and U4080 (N_4080,N_3799,N_3838);
and U4081 (N_4081,N_3298,N_2358);
or U4082 (N_4082,N_11,N_3559);
or U4083 (N_4083,N_2758,N_1839);
xor U4084 (N_4084,N_3394,N_1571);
nor U4085 (N_4085,N_609,N_3002);
nor U4086 (N_4086,N_3869,N_2692);
nand U4087 (N_4087,N_2932,N_3296);
nor U4088 (N_4088,N_3939,N_190);
nand U4089 (N_4089,N_2821,N_3779);
xnor U4090 (N_4090,N_806,N_89);
nor U4091 (N_4091,N_2265,N_3750);
and U4092 (N_4092,N_1049,N_2471);
xor U4093 (N_4093,N_60,N_2771);
nand U4094 (N_4094,N_561,N_3035);
or U4095 (N_4095,N_1757,N_206);
xnor U4096 (N_4096,N_3447,N_2309);
or U4097 (N_4097,N_2041,N_484);
nand U4098 (N_4098,N_2670,N_3754);
nor U4099 (N_4099,N_2738,N_3805);
nor U4100 (N_4100,N_2484,N_290);
or U4101 (N_4101,N_3075,N_2854);
or U4102 (N_4102,N_1525,N_178);
nor U4103 (N_4103,N_1427,N_332);
xor U4104 (N_4104,N_2027,N_61);
or U4105 (N_4105,N_3551,N_1880);
and U4106 (N_4106,N_8,N_2699);
xnor U4107 (N_4107,N_1169,N_3111);
nor U4108 (N_4108,N_971,N_975);
nand U4109 (N_4109,N_3846,N_2721);
nor U4110 (N_4110,N_1967,N_665);
or U4111 (N_4111,N_3466,N_3162);
nor U4112 (N_4112,N_995,N_2675);
xnor U4113 (N_4113,N_2452,N_2900);
and U4114 (N_4114,N_1108,N_353);
nand U4115 (N_4115,N_3874,N_2439);
or U4116 (N_4116,N_3099,N_780);
nor U4117 (N_4117,N_3458,N_1065);
nand U4118 (N_4118,N_2250,N_182);
and U4119 (N_4119,N_1148,N_1739);
and U4120 (N_4120,N_2038,N_3440);
xor U4121 (N_4121,N_585,N_3266);
nand U4122 (N_4122,N_2034,N_3530);
or U4123 (N_4123,N_2919,N_1628);
xor U4124 (N_4124,N_1255,N_1671);
xnor U4125 (N_4125,N_2295,N_3297);
and U4126 (N_4126,N_604,N_1177);
or U4127 (N_4127,N_3804,N_556);
nand U4128 (N_4128,N_2056,N_472);
or U4129 (N_4129,N_2101,N_1848);
and U4130 (N_4130,N_2216,N_2559);
or U4131 (N_4131,N_2181,N_99);
nand U4132 (N_4132,N_1716,N_3292);
and U4133 (N_4133,N_2194,N_0);
nor U4134 (N_4134,N_1356,N_3364);
or U4135 (N_4135,N_3400,N_3090);
and U4136 (N_4136,N_2136,N_1057);
nor U4137 (N_4137,N_1770,N_3715);
xnor U4138 (N_4138,N_1324,N_758);
and U4139 (N_4139,N_1857,N_3316);
nor U4140 (N_4140,N_1660,N_3365);
or U4141 (N_4141,N_1611,N_1156);
nor U4142 (N_4142,N_1672,N_2831);
nor U4143 (N_4143,N_3726,N_1134);
and U4144 (N_4144,N_176,N_3903);
or U4145 (N_4145,N_1973,N_1876);
xnor U4146 (N_4146,N_608,N_1413);
nand U4147 (N_4147,N_1154,N_3139);
xnor U4148 (N_4148,N_3335,N_2115);
nand U4149 (N_4149,N_2648,N_787);
nand U4150 (N_4150,N_3027,N_558);
xor U4151 (N_4151,N_1003,N_1898);
nor U4152 (N_4152,N_640,N_1728);
nor U4153 (N_4153,N_1888,N_2207);
or U4154 (N_4154,N_2196,N_2201);
and U4155 (N_4155,N_626,N_2506);
xnor U4156 (N_4156,N_792,N_2734);
xnor U4157 (N_4157,N_3360,N_49);
xnor U4158 (N_4158,N_3247,N_3349);
nor U4159 (N_4159,N_3023,N_3152);
or U4160 (N_4160,N_3556,N_413);
nand U4161 (N_4161,N_3615,N_1909);
xor U4162 (N_4162,N_2915,N_1925);
and U4163 (N_4163,N_468,N_2347);
xnor U4164 (N_4164,N_1483,N_1569);
and U4165 (N_4165,N_1480,N_2379);
xnor U4166 (N_4166,N_149,N_3240);
and U4167 (N_4167,N_2977,N_186);
or U4168 (N_4168,N_1692,N_1865);
and U4169 (N_4169,N_3171,N_3467);
nand U4170 (N_4170,N_3572,N_3573);
and U4171 (N_4171,N_3944,N_256);
nor U4172 (N_4172,N_2609,N_907);
nand U4173 (N_4173,N_255,N_2645);
xnor U4174 (N_4174,N_1624,N_727);
nand U4175 (N_4175,N_3119,N_3674);
or U4176 (N_4176,N_76,N_863);
and U4177 (N_4177,N_2271,N_1731);
nor U4178 (N_4178,N_3117,N_2328);
or U4179 (N_4179,N_831,N_2822);
or U4180 (N_4180,N_2377,N_3694);
nand U4181 (N_4181,N_2291,N_3338);
nor U4182 (N_4182,N_766,N_1500);
or U4183 (N_4183,N_1445,N_3806);
xnor U4184 (N_4184,N_2501,N_2555);
xnor U4185 (N_4185,N_465,N_1572);
and U4186 (N_4186,N_3876,N_2708);
and U4187 (N_4187,N_3657,N_2422);
or U4188 (N_4188,N_1603,N_1538);
xnor U4189 (N_4189,N_762,N_2685);
xor U4190 (N_4190,N_1393,N_53);
nand U4191 (N_4191,N_185,N_381);
nand U4192 (N_4192,N_1249,N_319);
or U4193 (N_4193,N_254,N_3990);
xor U4194 (N_4194,N_2170,N_3340);
and U4195 (N_4195,N_1798,N_965);
nand U4196 (N_4196,N_1547,N_1335);
or U4197 (N_4197,N_2499,N_3502);
nand U4198 (N_4198,N_1027,N_2402);
or U4199 (N_4199,N_3695,N_899);
xor U4200 (N_4200,N_1284,N_2596);
and U4201 (N_4201,N_3433,N_1106);
nand U4202 (N_4202,N_3016,N_1144);
and U4203 (N_4203,N_1792,N_269);
nand U4204 (N_4204,N_94,N_2902);
nor U4205 (N_4205,N_36,N_768);
xnor U4206 (N_4206,N_257,N_3672);
xor U4207 (N_4207,N_2512,N_3047);
nand U4208 (N_4208,N_1173,N_889);
or U4209 (N_4209,N_826,N_2391);
xnor U4210 (N_4210,N_1537,N_554);
or U4211 (N_4211,N_3531,N_2001);
and U4212 (N_4212,N_3148,N_3135);
and U4213 (N_4213,N_3260,N_3037);
nor U4214 (N_4214,N_494,N_1062);
and U4215 (N_4215,N_2239,N_3866);
xnor U4216 (N_4216,N_3059,N_1655);
or U4217 (N_4217,N_1127,N_1205);
xnor U4218 (N_4218,N_675,N_2053);
nand U4219 (N_4219,N_3346,N_2209);
and U4220 (N_4220,N_1392,N_2128);
or U4221 (N_4221,N_643,N_1153);
and U4222 (N_4222,N_1286,N_1662);
xor U4223 (N_4223,N_2202,N_2278);
and U4224 (N_4224,N_3490,N_2470);
or U4225 (N_4225,N_2500,N_1970);
xnor U4226 (N_4226,N_349,N_86);
nand U4227 (N_4227,N_773,N_3051);
xor U4228 (N_4228,N_3147,N_2937);
or U4229 (N_4229,N_3107,N_1942);
nor U4230 (N_4230,N_3217,N_3317);
and U4231 (N_4231,N_3853,N_2116);
nor U4232 (N_4232,N_2762,N_286);
xor U4233 (N_4233,N_2330,N_2518);
or U4234 (N_4234,N_877,N_93);
xor U4235 (N_4235,N_3620,N_1453);
and U4236 (N_4236,N_430,N_1311);
nor U4237 (N_4237,N_3542,N_2917);
nor U4238 (N_4238,N_2816,N_1800);
and U4239 (N_4239,N_576,N_3771);
nor U4240 (N_4240,N_1962,N_2415);
nand U4241 (N_4241,N_3309,N_2087);
xor U4242 (N_4242,N_1685,N_1227);
nand U4243 (N_4243,N_418,N_315);
xnor U4244 (N_4244,N_2749,N_815);
nor U4245 (N_4245,N_865,N_2554);
and U4246 (N_4246,N_2051,N_1410);
nor U4247 (N_4247,N_1400,N_450);
xnor U4248 (N_4248,N_2560,N_2097);
or U4249 (N_4249,N_1610,N_3566);
nand U4250 (N_4250,N_2066,N_3156);
nor U4251 (N_4251,N_2033,N_2705);
xor U4252 (N_4252,N_2127,N_3505);
nand U4253 (N_4253,N_1763,N_3391);
nor U4254 (N_4254,N_1122,N_226);
nand U4255 (N_4255,N_1318,N_3623);
or U4256 (N_4256,N_978,N_3702);
nand U4257 (N_4257,N_326,N_2174);
nand U4258 (N_4258,N_1308,N_1023);
nand U4259 (N_4259,N_617,N_3794);
and U4260 (N_4260,N_1162,N_3412);
xor U4261 (N_4261,N_1194,N_632);
and U4262 (N_4262,N_125,N_3060);
nor U4263 (N_4263,N_3870,N_1218);
or U4264 (N_4264,N_3508,N_208);
nor U4265 (N_4265,N_1588,N_3863);
nor U4266 (N_4266,N_920,N_876);
or U4267 (N_4267,N_657,N_1353);
xnor U4268 (N_4268,N_1653,N_778);
nand U4269 (N_4269,N_732,N_793);
xor U4270 (N_4270,N_730,N_3783);
nand U4271 (N_4271,N_2859,N_2600);
nor U4272 (N_4272,N_33,N_1337);
nand U4273 (N_4273,N_387,N_1639);
nor U4274 (N_4274,N_1586,N_3905);
and U4275 (N_4275,N_1248,N_3048);
or U4276 (N_4276,N_954,N_3528);
or U4277 (N_4277,N_3320,N_2766);
and U4278 (N_4278,N_1854,N_1747);
and U4279 (N_4279,N_3359,N_3040);
or U4280 (N_4280,N_3256,N_588);
or U4281 (N_4281,N_3115,N_127);
nor U4282 (N_4282,N_3402,N_3933);
nor U4283 (N_4283,N_3473,N_1447);
nand U4284 (N_4284,N_1836,N_227);
nand U4285 (N_4285,N_151,N_1107);
nor U4286 (N_4286,N_2048,N_2121);
nand U4287 (N_4287,N_2643,N_1405);
and U4288 (N_4288,N_489,N_1046);
or U4289 (N_4289,N_48,N_195);
or U4290 (N_4290,N_3153,N_1222);
nand U4291 (N_4291,N_962,N_2994);
and U4292 (N_4292,N_2795,N_2975);
and U4293 (N_4293,N_1828,N_21);
xnor U4294 (N_4294,N_3666,N_647);
xnor U4295 (N_4295,N_1364,N_1109);
or U4296 (N_4296,N_2599,N_1919);
xnor U4297 (N_4297,N_467,N_458);
nor U4298 (N_4298,N_2695,N_1256);
or U4299 (N_4299,N_1784,N_648);
and U4300 (N_4300,N_2140,N_3746);
xnor U4301 (N_4301,N_1564,N_2388);
xnor U4302 (N_4302,N_2163,N_398);
nor U4303 (N_4303,N_2578,N_2535);
nor U4304 (N_4304,N_565,N_2827);
or U4305 (N_4305,N_2063,N_2025);
nand U4306 (N_4306,N_1972,N_2934);
and U4307 (N_4307,N_423,N_2938);
and U4308 (N_4308,N_1893,N_3303);
xor U4309 (N_4309,N_2857,N_878);
and U4310 (N_4310,N_1831,N_321);
and U4311 (N_4311,N_2117,N_618);
nor U4312 (N_4312,N_305,N_331);
nand U4313 (N_4313,N_998,N_1391);
xor U4314 (N_4314,N_2335,N_3136);
or U4315 (N_4315,N_531,N_1724);
xnor U4316 (N_4316,N_901,N_989);
nand U4317 (N_4317,N_1577,N_1645);
xor U4318 (N_4318,N_3498,N_1971);
nor U4319 (N_4319,N_1323,N_2299);
nand U4320 (N_4320,N_3398,N_1551);
or U4321 (N_4321,N_3149,N_1584);
nand U4322 (N_4322,N_3534,N_3722);
or U4323 (N_4323,N_402,N_2050);
nand U4324 (N_4324,N_3062,N_3920);
nand U4325 (N_4325,N_1138,N_2185);
and U4326 (N_4326,N_2214,N_893);
nand U4327 (N_4327,N_2767,N_1515);
xor U4328 (N_4328,N_3367,N_3204);
nand U4329 (N_4329,N_1600,N_1799);
xor U4330 (N_4330,N_3506,N_352);
nor U4331 (N_4331,N_1633,N_246);
or U4332 (N_4332,N_1403,N_3713);
nand U4333 (N_4333,N_2594,N_1191);
or U4334 (N_4334,N_1220,N_533);
and U4335 (N_4335,N_2962,N_371);
and U4336 (N_4336,N_1167,N_859);
and U4337 (N_4337,N_983,N_911);
nand U4338 (N_4338,N_3834,N_3717);
or U4339 (N_4339,N_3568,N_1917);
xor U4340 (N_4340,N_2589,N_3668);
and U4341 (N_4341,N_3503,N_80);
nand U4342 (N_4342,N_902,N_1711);
or U4343 (N_4343,N_1047,N_2088);
nor U4344 (N_4344,N_1729,N_1690);
nor U4345 (N_4345,N_2445,N_2444);
nor U4346 (N_4346,N_1612,N_215);
or U4347 (N_4347,N_504,N_2825);
and U4348 (N_4348,N_1873,N_3789);
and U4349 (N_4349,N_3667,N_20);
nor U4350 (N_4350,N_2591,N_38);
or U4351 (N_4351,N_3245,N_433);
nand U4352 (N_4352,N_275,N_216);
xor U4353 (N_4353,N_137,N_1691);
nor U4354 (N_4354,N_2475,N_2243);
xnor U4355 (N_4355,N_3486,N_2944);
nor U4356 (N_4356,N_392,N_1037);
or U4357 (N_4357,N_3329,N_3214);
xnor U4358 (N_4358,N_1123,N_3688);
nand U4359 (N_4359,N_3238,N_887);
nor U4360 (N_4360,N_442,N_761);
nand U4361 (N_4361,N_3819,N_3138);
nand U4362 (N_4362,N_3773,N_3234);
nor U4363 (N_4363,N_3686,N_2376);
xor U4364 (N_4364,N_3425,N_3922);
or U4365 (N_4365,N_3629,N_2720);
xnor U4366 (N_4366,N_2964,N_2782);
nor U4367 (N_4367,N_2809,N_654);
and U4368 (N_4368,N_473,N_2636);
and U4369 (N_4369,N_2907,N_1228);
and U4370 (N_4370,N_1843,N_710);
xor U4371 (N_4371,N_2344,N_1964);
nand U4372 (N_4372,N_129,N_1811);
xnor U4373 (N_4373,N_2916,N_1847);
and U4374 (N_4374,N_1579,N_747);
or U4375 (N_4375,N_2109,N_621);
or U4376 (N_4376,N_2089,N_1735);
xor U4377 (N_4377,N_3720,N_2306);
and U4378 (N_4378,N_1221,N_302);
nor U4379 (N_4379,N_1915,N_3463);
xor U4380 (N_4380,N_2218,N_1315);
or U4381 (N_4381,N_281,N_2204);
and U4382 (N_4382,N_1506,N_2808);
nand U4383 (N_4383,N_2725,N_3314);
nor U4384 (N_4384,N_3019,N_2175);
and U4385 (N_4385,N_2419,N_557);
xnor U4386 (N_4386,N_1926,N_1781);
nand U4387 (N_4387,N_2006,N_469);
nand U4388 (N_4388,N_3818,N_2715);
nand U4389 (N_4389,N_84,N_2741);
xor U4390 (N_4390,N_1486,N_2910);
nand U4391 (N_4391,N_1912,N_1754);
nor U4392 (N_4392,N_2093,N_2264);
and U4393 (N_4393,N_3843,N_429);
or U4394 (N_4394,N_2655,N_2681);
xnor U4395 (N_4395,N_1009,N_1869);
nor U4396 (N_4396,N_3327,N_2346);
nand U4397 (N_4397,N_1072,N_2684);
and U4398 (N_4398,N_2287,N_3821);
nand U4399 (N_4399,N_1230,N_1945);
nor U4400 (N_4400,N_847,N_3350);
nor U4401 (N_4401,N_2094,N_3943);
nand U4402 (N_4402,N_3949,N_879);
nand U4403 (N_4403,N_3637,N_2270);
xnor U4404 (N_4404,N_2550,N_355);
and U4405 (N_4405,N_3413,N_91);
and U4406 (N_4406,N_662,N_313);
nor U4407 (N_4407,N_3927,N_3093);
nand U4408 (N_4408,N_1197,N_3646);
and U4409 (N_4409,N_250,N_703);
nor U4410 (N_4410,N_3801,N_3606);
nor U4411 (N_4411,N_2482,N_3822);
nor U4412 (N_4412,N_2068,N_722);
nor U4413 (N_4413,N_56,N_3553);
and U4414 (N_4414,N_264,N_1712);
nor U4415 (N_4415,N_800,N_763);
nand U4416 (N_4416,N_3507,N_2325);
or U4417 (N_4417,N_2768,N_976);
and U4418 (N_4418,N_201,N_134);
nand U4419 (N_4419,N_897,N_303);
and U4420 (N_4420,N_165,N_1914);
and U4421 (N_4421,N_933,N_414);
xnor U4422 (N_4422,N_2014,N_3258);
nand U4423 (N_4423,N_2362,N_1702);
nand U4424 (N_4424,N_3068,N_2814);
nand U4425 (N_4425,N_1402,N_559);
xnor U4426 (N_4426,N_691,N_2933);
and U4427 (N_4427,N_2948,N_2032);
and U4428 (N_4428,N_1257,N_271);
and U4429 (N_4429,N_1432,N_2940);
and U4430 (N_4430,N_2774,N_2081);
nand U4431 (N_4431,N_1786,N_1576);
or U4432 (N_4432,N_374,N_2205);
and U4433 (N_4433,N_2778,N_3181);
nand U4434 (N_4434,N_2273,N_3194);
nand U4435 (N_4435,N_492,N_335);
and U4436 (N_4436,N_1526,N_3431);
xnor U4437 (N_4437,N_1442,N_2030);
xnor U4438 (N_4438,N_291,N_1259);
nand U4439 (N_4439,N_836,N_3174);
nor U4440 (N_4440,N_2074,N_3435);
or U4441 (N_4441,N_1170,N_1916);
nor U4442 (N_4442,N_3867,N_3848);
nor U4443 (N_4443,N_148,N_2083);
nand U4444 (N_4444,N_994,N_3523);
xnor U4445 (N_4445,N_3893,N_2612);
and U4446 (N_4446,N_2252,N_759);
nand U4447 (N_4447,N_2256,N_1598);
and U4448 (N_4448,N_3705,N_3081);
xor U4449 (N_4449,N_1592,N_3800);
nand U4450 (N_4450,N_39,N_3222);
xor U4451 (N_4451,N_2073,N_3696);
or U4452 (N_4452,N_2798,N_2105);
or U4453 (N_4453,N_90,N_3179);
nand U4454 (N_4454,N_767,N_2790);
xnor U4455 (N_4455,N_2451,N_112);
or U4456 (N_4456,N_1495,N_580);
or U4457 (N_4457,N_3225,N_2625);
nor U4458 (N_4458,N_1505,N_3756);
nor U4459 (N_4459,N_1264,N_2572);
xnor U4460 (N_4460,N_510,N_3041);
nor U4461 (N_4461,N_3061,N_168);
nand U4462 (N_4462,N_1549,N_1140);
xor U4463 (N_4463,N_1431,N_3393);
or U4464 (N_4464,N_2453,N_3069);
nand U4465 (N_4465,N_1136,N_29);
nand U4466 (N_4466,N_2693,N_3462);
nor U4467 (N_4467,N_1285,N_2383);
and U4468 (N_4468,N_3760,N_1275);
nor U4469 (N_4469,N_3894,N_30);
and U4470 (N_4470,N_1082,N_622);
nor U4471 (N_4471,N_288,N_3299);
xor U4472 (N_4472,N_1244,N_2180);
nor U4473 (N_4473,N_200,N_328);
and U4474 (N_4474,N_1950,N_699);
and U4475 (N_4475,N_3759,N_635);
xor U4476 (N_4476,N_1802,N_3951);
nor U4477 (N_4477,N_1790,N_1198);
or U4478 (N_4478,N_3628,N_3246);
nor U4479 (N_4479,N_2435,N_1440);
or U4480 (N_4480,N_2421,N_2161);
nor U4481 (N_4481,N_1000,N_470);
xor U4482 (N_4482,N_3786,N_2844);
and U4483 (N_4483,N_726,N_986);
nor U4484 (N_4484,N_3112,N_2040);
nor U4485 (N_4485,N_3029,N_2381);
nand U4486 (N_4486,N_2761,N_1556);
nand U4487 (N_4487,N_2903,N_3558);
nor U4488 (N_4488,N_3187,N_3422);
and U4489 (N_4489,N_3900,N_1852);
nand U4490 (N_4490,N_393,N_1605);
and U4491 (N_4491,N_3382,N_2158);
or U4492 (N_4492,N_1988,N_3362);
nand U4493 (N_4493,N_3691,N_2748);
nand U4494 (N_4494,N_2246,N_1710);
and U4495 (N_4495,N_929,N_3969);
or U4496 (N_4496,N_1089,N_1636);
xor U4497 (N_4497,N_2261,N_420);
xor U4498 (N_4498,N_3459,N_3782);
nand U4499 (N_4499,N_612,N_925);
and U4500 (N_4500,N_3342,N_3923);
and U4501 (N_4501,N_1246,N_322);
xor U4502 (N_4502,N_904,N_1087);
nor U4503 (N_4503,N_528,N_388);
nand U4504 (N_4504,N_3525,N_2495);
or U4505 (N_4505,N_2448,N_886);
xnor U4506 (N_4506,N_3496,N_2614);
xnor U4507 (N_4507,N_2449,N_752);
nor U4508 (N_4508,N_2662,N_2062);
xor U4509 (N_4509,N_583,N_3043);
nand U4510 (N_4510,N_564,N_3988);
nand U4511 (N_4511,N_297,N_28);
nand U4512 (N_4512,N_1996,N_3840);
or U4513 (N_4513,N_2356,N_3243);
xnor U4514 (N_4514,N_2232,N_3529);
or U4515 (N_4515,N_3512,N_1938);
and U4516 (N_4516,N_1143,N_2921);
or U4517 (N_4517,N_285,N_3065);
nor U4518 (N_4518,N_3913,N_299);
and U4519 (N_4519,N_3910,N_812);
nor U4520 (N_4520,N_1680,N_2286);
nor U4521 (N_4521,N_713,N_3374);
nand U4522 (N_4522,N_1497,N_3960);
and U4523 (N_4523,N_610,N_1560);
and U4524 (N_4524,N_2710,N_3595);
or U4525 (N_4525,N_2258,N_1150);
xor U4526 (N_4526,N_530,N_3419);
nand U4527 (N_4527,N_241,N_2031);
xnor U4528 (N_4528,N_1425,N_2301);
or U4529 (N_4529,N_1312,N_895);
nand U4530 (N_4530,N_2698,N_3571);
nand U4531 (N_4531,N_720,N_3828);
nand U4532 (N_4532,N_1266,N_3544);
or U4533 (N_4533,N_1086,N_3254);
nand U4534 (N_4534,N_2103,N_2314);
nand U4535 (N_4535,N_2037,N_1382);
and U4536 (N_4536,N_1409,N_3926);
or U4537 (N_4537,N_2085,N_1322);
xnor U4538 (N_4538,N_1163,N_356);
xnor U4539 (N_4539,N_3968,N_1243);
xor U4540 (N_4540,N_2259,N_2724);
nand U4541 (N_4541,N_3873,N_3429);
nor U4542 (N_4542,N_278,N_3678);
nor U4543 (N_4543,N_62,N_2626);
nor U4544 (N_4544,N_2678,N_1271);
xnor U4545 (N_4545,N_3120,N_2642);
nand U4546 (N_4546,N_688,N_1548);
nor U4547 (N_4547,N_3574,N_2169);
nor U4548 (N_4548,N_218,N_639);
xnor U4549 (N_4549,N_3956,N_619);
nand U4550 (N_4550,N_3347,N_829);
xnor U4551 (N_4551,N_3835,N_1454);
and U4552 (N_4552,N_2289,N_2015);
or U4553 (N_4553,N_3640,N_982);
nand U4554 (N_4554,N_2888,N_3231);
xor U4555 (N_4555,N_2928,N_858);
or U4556 (N_4556,N_1567,N_3094);
nor U4557 (N_4557,N_3679,N_3963);
and U4558 (N_4558,N_1963,N_2987);
or U4559 (N_4559,N_2564,N_799);
or U4560 (N_4560,N_1407,N_1826);
or U4561 (N_4561,N_344,N_891);
xor U4562 (N_4562,N_1738,N_1935);
and U4563 (N_4563,N_104,N_3934);
and U4564 (N_4564,N_2873,N_2389);
nor U4565 (N_4565,N_2714,N_2473);
xor U4566 (N_4566,N_1542,N_1471);
nor U4567 (N_4567,N_514,N_1517);
or U4568 (N_4568,N_3165,N_3781);
nor U4569 (N_4569,N_1727,N_2820);
xor U4570 (N_4570,N_2755,N_2998);
nand U4571 (N_4571,N_2082,N_1119);
or U4572 (N_4572,N_947,N_716);
nor U4573 (N_4573,N_2497,N_2503);
nand U4574 (N_4574,N_1607,N_2401);
and U4575 (N_4575,N_3849,N_123);
xor U4576 (N_4576,N_1806,N_1386);
xor U4577 (N_4577,N_935,N_293);
and U4578 (N_4578,N_362,N_2533);
nor U4579 (N_4579,N_3698,N_1184);
xnor U4580 (N_4580,N_1827,N_138);
xor U4581 (N_4581,N_2340,N_677);
xor U4582 (N_4582,N_2861,N_3711);
xor U4583 (N_4583,N_1260,N_2268);
xor U4584 (N_4584,N_2851,N_549);
nand U4585 (N_4585,N_3184,N_3066);
and U4586 (N_4586,N_2542,N_1530);
nor U4587 (N_4587,N_1820,N_3197);
nand U4588 (N_4588,N_1928,N_1956);
nor U4589 (N_4589,N_880,N_1487);
or U4590 (N_4590,N_2474,N_813);
and U4591 (N_4591,N_551,N_2858);
xor U4592 (N_4592,N_1024,N_3743);
nand U4593 (N_4593,N_2212,N_2164);
or U4594 (N_4594,N_2187,N_1390);
nor U4595 (N_4595,N_3159,N_2717);
nor U4596 (N_4596,N_705,N_3740);
nor U4597 (N_4597,N_1299,N_811);
nand U4598 (N_4598,N_435,N_3106);
nand U4599 (N_4599,N_211,N_2162);
or U4600 (N_4600,N_2586,N_1875);
nand U4601 (N_4601,N_2551,N_2241);
xnor U4602 (N_4602,N_2323,N_3470);
xor U4603 (N_4603,N_399,N_3889);
or U4604 (N_4604,N_707,N_213);
xnor U4605 (N_4605,N_3975,N_3414);
nand U4606 (N_4606,N_159,N_2864);
xnor U4607 (N_4607,N_2628,N_3141);
xor U4608 (N_4608,N_242,N_196);
nor U4609 (N_4609,N_3005,N_3288);
and U4610 (N_4610,N_243,N_2337);
nand U4611 (N_4611,N_2157,N_3239);
or U4612 (N_4612,N_1200,N_3383);
and U4613 (N_4613,N_888,N_3912);
and U4614 (N_4614,N_1051,N_575);
nand U4615 (N_4615,N_2333,N_2407);
or U4616 (N_4616,N_327,N_3052);
nand U4617 (N_4617,N_2566,N_330);
xnor U4618 (N_4618,N_3888,N_3565);
nor U4619 (N_4619,N_1080,N_1726);
nor U4620 (N_4620,N_323,N_124);
nand U4621 (N_4621,N_1937,N_1036);
xor U4622 (N_4622,N_3205,N_3264);
or U4623 (N_4623,N_3929,N_1889);
and U4624 (N_4624,N_1289,N_2787);
and U4625 (N_4625,N_809,N_1626);
nor U4626 (N_4626,N_956,N_436);
nor U4627 (N_4627,N_320,N_267);
or U4628 (N_4628,N_2284,N_477);
and U4629 (N_4629,N_3710,N_2438);
nand U4630 (N_4630,N_1947,N_1578);
xor U4631 (N_4631,N_3476,N_1021);
nor U4632 (N_4632,N_1306,N_3203);
nor U4633 (N_4633,N_1554,N_2549);
or U4634 (N_4634,N_1294,N_854);
and U4635 (N_4635,N_2478,N_2382);
or U4636 (N_4636,N_3725,N_3585);
nand U4637 (N_4637,N_2236,N_3259);
and U4638 (N_4638,N_3954,N_2305);
and U4639 (N_4639,N_3182,N_3931);
and U4640 (N_4640,N_574,N_1536);
and U4641 (N_4641,N_903,N_1860);
nand U4642 (N_4642,N_937,N_2024);
nor U4643 (N_4643,N_2508,N_140);
xnor U4644 (N_4644,N_2529,N_2702);
nand U4645 (N_4645,N_1235,N_1809);
and U4646 (N_4646,N_1979,N_2889);
nor U4647 (N_4647,N_3644,N_2627);
and U4648 (N_4648,N_2983,N_3864);
xnor U4649 (N_4649,N_1539,N_3911);
and U4650 (N_4650,N_1434,N_1514);
xnor U4651 (N_4651,N_2908,N_1261);
and U4652 (N_4652,N_287,N_95);
nand U4653 (N_4653,N_2806,N_2640);
xor U4654 (N_4654,N_2331,N_2226);
or U4655 (N_4655,N_3377,N_1749);
xor U4656 (N_4656,N_2080,N_1076);
and U4657 (N_4657,N_221,N_194);
xor U4658 (N_4658,N_3937,N_1531);
and U4659 (N_4659,N_1348,N_731);
nand U4660 (N_4660,N_2192,N_1638);
or U4661 (N_4661,N_3169,N_788);
and U4662 (N_4662,N_2429,N_2968);
xor U4663 (N_4663,N_2131,N_3897);
or U4664 (N_4664,N_2709,N_2035);
xor U4665 (N_4665,N_993,N_1631);
and U4666 (N_4666,N_3714,N_1849);
xnor U4667 (N_4667,N_1778,N_3124);
and U4668 (N_4668,N_3488,N_1387);
or U4669 (N_4669,N_3191,N_2369);
and U4670 (N_4670,N_1213,N_3524);
xor U4671 (N_4671,N_3677,N_1438);
or U4672 (N_4672,N_63,N_2133);
nor U4673 (N_4673,N_894,N_1361);
nor U4674 (N_4674,N_2052,N_1053);
and U4675 (N_4675,N_220,N_1006);
nor U4676 (N_4676,N_443,N_1030);
nand U4677 (N_4677,N_1635,N_2623);
nand U4678 (N_4678,N_2641,N_2293);
and U4679 (N_4679,N_361,N_3596);
nand U4680 (N_4680,N_3302,N_3510);
xnor U4681 (N_4681,N_1813,N_916);
and U4682 (N_4682,N_1367,N_1597);
nor U4683 (N_4683,N_1941,N_3334);
nand U4684 (N_4684,N_3177,N_512);
nor U4685 (N_4685,N_3955,N_2279);
nor U4686 (N_4686,N_3830,N_3031);
and U4687 (N_4687,N_2716,N_437);
nor U4688 (N_4688,N_1667,N_3178);
xnor U4689 (N_4689,N_2510,N_279);
or U4690 (N_4690,N_2598,N_629);
nand U4691 (N_4691,N_997,N_1519);
and U4692 (N_4692,N_350,N_3454);
xor U4693 (N_4693,N_2991,N_3736);
xor U4694 (N_4694,N_571,N_3526);
and U4695 (N_4695,N_2091,N_3557);
xor U4696 (N_4696,N_542,N_2124);
xnor U4697 (N_4697,N_708,N_1630);
nand U4698 (N_4698,N_1301,N_1679);
and U4699 (N_4699,N_2880,N_1242);
nand U4700 (N_4700,N_1359,N_742);
nor U4701 (N_4701,N_3121,N_2426);
nor U4702 (N_4702,N_1274,N_2217);
and U4703 (N_4703,N_2156,N_292);
xnor U4704 (N_4704,N_623,N_77);
and U4705 (N_4705,N_1507,N_3586);
or U4706 (N_4706,N_1974,N_3267);
or U4707 (N_4707,N_3129,N_2777);
and U4708 (N_4708,N_1095,N_680);
and U4709 (N_4709,N_454,N_2459);
and U4710 (N_4710,N_3064,N_434);
and U4711 (N_4711,N_1899,N_2573);
xnor U4712 (N_4712,N_1472,N_50);
nor U4713 (N_4713,N_1159,N_2483);
xor U4714 (N_4714,N_2899,N_2894);
nor U4715 (N_4715,N_615,N_2315);
and U4716 (N_4716,N_3265,N_1022);
xor U4717 (N_4717,N_1373,N_3658);
and U4718 (N_4718,N_2498,N_1817);
nor U4719 (N_4719,N_797,N_209);
or U4720 (N_4720,N_3013,N_2727);
nor U4721 (N_4721,N_1965,N_2875);
or U4722 (N_4722,N_2002,N_306);
nor U4723 (N_4723,N_2186,N_2447);
and U4724 (N_4724,N_1350,N_464);
nand U4725 (N_4725,N_3289,N_1279);
nor U4726 (N_4726,N_1887,N_1146);
nor U4727 (N_4727,N_3718,N_2350);
or U4728 (N_4728,N_3815,N_3537);
xor U4729 (N_4729,N_3663,N_967);
and U4730 (N_4730,N_485,N_3883);
or U4731 (N_4731,N_3724,N_689);
xor U4732 (N_4732,N_2905,N_2607);
and U4733 (N_4733,N_1424,N_1559);
or U4734 (N_4734,N_1396,N_1878);
nand U4735 (N_4735,N_3639,N_2078);
xor U4736 (N_4736,N_1034,N_2847);
or U4737 (N_4737,N_2819,N_3981);
or U4738 (N_4738,N_336,N_1874);
and U4739 (N_4739,N_3483,N_3244);
or U4740 (N_4740,N_3599,N_1705);
xor U4741 (N_4741,N_658,N_1978);
or U4742 (N_4742,N_2865,N_274);
nand U4743 (N_4743,N_3113,N_169);
or U4744 (N_4744,N_202,N_1094);
and U4745 (N_4745,N_534,N_3076);
and U4746 (N_4746,N_2581,N_2828);
or U4747 (N_4747,N_2047,N_2011);
nand U4748 (N_4748,N_2108,N_862);
nand U4749 (N_4749,N_1940,N_318);
nand U4750 (N_4750,N_3511,N_1565);
nor U4751 (N_4751,N_3940,N_1871);
xor U4752 (N_4752,N_3520,N_592);
nand U4753 (N_4753,N_972,N_3032);
nand U4754 (N_4754,N_3622,N_1052);
xnor U4755 (N_4755,N_3536,N_1742);
and U4756 (N_4756,N_425,N_2676);
nand U4757 (N_4757,N_97,N_309);
and U4758 (N_4758,N_2059,N_296);
nand U4759 (N_4759,N_341,N_2332);
or U4760 (N_4760,N_1439,N_553);
nand U4761 (N_4761,N_1112,N_3499);
nor U4762 (N_4762,N_146,N_1994);
xnor U4763 (N_4763,N_709,N_2810);
nor U4764 (N_4764,N_391,N_3154);
xnor U4765 (N_4765,N_415,N_1589);
nand U4766 (N_4766,N_3318,N_711);
nor U4767 (N_4767,N_440,N_1268);
nand U4768 (N_4768,N_3729,N_987);
xor U4769 (N_4769,N_3494,N_3020);
nand U4770 (N_4770,N_1263,N_2479);
nand U4771 (N_4771,N_2970,N_1171);
nor U4772 (N_4772,N_1683,N_3410);
nor U4773 (N_4773,N_2235,N_1510);
nand U4774 (N_4774,N_3407,N_961);
nand U4775 (N_4775,N_1341,N_1302);
xnor U4776 (N_4776,N_1574,N_2060);
nor U4777 (N_4777,N_3906,N_3581);
xnor U4778 (N_4778,N_363,N_408);
nand U4779 (N_4779,N_3868,N_1656);
or U4780 (N_4780,N_2244,N_2366);
or U4781 (N_4781,N_3627,N_2606);
or U4782 (N_4782,N_1345,N_34);
or U4783 (N_4783,N_3368,N_1428);
nand U4784 (N_4784,N_3301,N_1099);
nand U4785 (N_4785,N_2148,N_1709);
nand U4786 (N_4786,N_900,N_2743);
and U4787 (N_4787,N_3823,N_3567);
nand U4788 (N_4788,N_1856,N_3827);
and U4789 (N_4789,N_3313,N_644);
and U4790 (N_4790,N_2871,N_1474);
and U4791 (N_4791,N_3993,N_3237);
nor U4792 (N_4792,N_452,N_785);
nor U4793 (N_4793,N_938,N_397);
and U4794 (N_4794,N_3034,N_2657);
nand U4795 (N_4795,N_1659,N_3208);
nand U4796 (N_4796,N_3996,N_2496);
nand U4797 (N_4797,N_1193,N_3408);
and U4798 (N_4798,N_345,N_466);
and U4799 (N_4799,N_833,N_502);
and U4800 (N_4800,N_3279,N_655);
or U4801 (N_4801,N_2206,N_1459);
nor U4802 (N_4802,N_842,N_1657);
nor U4803 (N_4803,N_1835,N_2633);
nor U4804 (N_4804,N_1165,N_2579);
or U4805 (N_4805,N_1241,N_1297);
nand U4806 (N_4806,N_798,N_1011);
nand U4807 (N_4807,N_3693,N_1756);
nor U4808 (N_4808,N_3332,N_3485);
xnor U4809 (N_4809,N_192,N_3212);
xor U4810 (N_4810,N_1552,N_808);
and U4811 (N_4811,N_3641,N_3004);
or U4812 (N_4812,N_934,N_2319);
xnor U4813 (N_4813,N_1029,N_3095);
xnor U4814 (N_4814,N_3130,N_1103);
and U4815 (N_4815,N_2141,N_3102);
nor U4816 (N_4816,N_2803,N_1216);
or U4817 (N_4817,N_74,N_2711);
or U4818 (N_4818,N_2815,N_2920);
or U4819 (N_4819,N_2208,N_24);
nand U4820 (N_4820,N_980,N_3085);
nand U4821 (N_4821,N_1287,N_2923);
or U4822 (N_4822,N_653,N_3997);
xnor U4823 (N_4823,N_411,N_550);
or U4824 (N_4824,N_579,N_1277);
nor U4825 (N_4825,N_1070,N_142);
or U4826 (N_4826,N_184,N_2008);
nand U4827 (N_4827,N_757,N_2513);
and U4828 (N_4828,N_2147,N_776);
and U4829 (N_4829,N_1897,N_3946);
nor U4830 (N_4830,N_2511,N_2872);
xnor U4831 (N_4831,N_2621,N_3189);
xnor U4832 (N_4832,N_147,N_2488);
nor U4833 (N_4833,N_188,N_3457);
nand U4834 (N_4834,N_3844,N_2849);
or U4835 (N_4835,N_2493,N_1766);
nand U4836 (N_4836,N_3763,N_2114);
nand U4837 (N_4837,N_734,N_131);
xor U4838 (N_4838,N_1952,N_3480);
nand U4839 (N_4839,N_1535,N_6);
xor U4840 (N_4840,N_1933,N_791);
nor U4841 (N_4841,N_2839,N_1824);
nor U4842 (N_4842,N_1147,N_1291);
or U4843 (N_4843,N_2745,N_339);
nor U4844 (N_4844,N_1999,N_2067);
xnor U4845 (N_4845,N_3635,N_3366);
nor U4846 (N_4846,N_1696,N_3209);
or U4847 (N_4847,N_1805,N_2225);
or U4848 (N_4848,N_3578,N_917);
and U4849 (N_4849,N_3469,N_317);
or U4850 (N_4850,N_2142,N_3907);
and U4851 (N_4851,N_15,N_2992);
nand U4852 (N_4852,N_130,N_3896);
or U4853 (N_4853,N_3613,N_3183);
xnor U4854 (N_4854,N_2656,N_2637);
nor U4855 (N_4855,N_171,N_2957);
nor U4856 (N_4856,N_1236,N_912);
xor U4857 (N_4857,N_244,N_3028);
or U4858 (N_4858,N_522,N_2238);
and U4859 (N_4859,N_3087,N_2739);
and U4860 (N_4860,N_3734,N_781);
xor U4861 (N_4861,N_2913,N_1695);
nor U4862 (N_4862,N_1295,N_2914);
or U4863 (N_4863,N_2742,N_1238);
or U4864 (N_4864,N_3477,N_167);
or U4865 (N_4865,N_277,N_2995);
or U4866 (N_4866,N_750,N_1478);
nand U4867 (N_4867,N_2075,N_1783);
and U4868 (N_4868,N_3180,N_482);
or U4869 (N_4869,N_1634,N_3088);
nand U4870 (N_4870,N_942,N_1460);
xor U4871 (N_4871,N_3448,N_3653);
nand U4872 (N_4872,N_3426,N_3648);
xnor U4873 (N_4873,N_3744,N_1896);
and U4874 (N_4874,N_1793,N_3116);
nand U4875 (N_4875,N_43,N_3739);
or U4876 (N_4876,N_2516,N_1580);
nor U4877 (N_4877,N_496,N_1563);
nor U4878 (N_4878,N_3521,N_3624);
nand U4879 (N_4879,N_2020,N_890);
or U4880 (N_4880,N_686,N_2390);
and U4881 (N_4881,N_1644,N_2582);
xor U4882 (N_4882,N_873,N_1374);
or U4883 (N_4883,N_2746,N_310);
xor U4884 (N_4884,N_2950,N_73);
and U4885 (N_4885,N_2414,N_910);
or U4886 (N_4886,N_1853,N_3860);
or U4887 (N_4887,N_2895,N_3386);
or U4888 (N_4888,N_1841,N_2489);
or U4889 (N_4889,N_3131,N_3957);
xor U4890 (N_4890,N_2321,N_162);
xor U4891 (N_4891,N_394,N_535);
and U4892 (N_4892,N_3767,N_1251);
and U4893 (N_4893,N_2841,N_2049);
and U4894 (N_4894,N_844,N_3861);
and U4895 (N_4895,N_3044,N_463);
and U4896 (N_4896,N_2647,N_544);
and U4897 (N_4897,N_821,N_985);
nor U4898 (N_4898,N_3058,N_3038);
and U4899 (N_4899,N_1900,N_1550);
nor U4900 (N_4900,N_3757,N_1250);
or U4901 (N_4901,N_490,N_3);
nand U4902 (N_4902,N_1771,N_740);
xor U4903 (N_4903,N_204,N_2690);
or U4904 (N_4904,N_3337,N_2341);
nand U4905 (N_4905,N_3151,N_2431);
nor U4906 (N_4906,N_2165,N_2021);
nand U4907 (N_4907,N_424,N_3974);
nand U4908 (N_4908,N_1433,N_1186);
nand U4909 (N_4909,N_2371,N_1762);
and U4910 (N_4910,N_3315,N_2679);
and U4911 (N_4911,N_802,N_3953);
nor U4912 (N_4912,N_2359,N_174);
xor U4913 (N_4913,N_1518,N_2373);
nor U4914 (N_4914,N_673,N_2461);
and U4915 (N_4915,N_1025,N_2349);
and U4916 (N_4916,N_2791,N_1594);
and U4917 (N_4917,N_3700,N_581);
nor U4918 (N_4918,N_695,N_3269);
nand U4919 (N_4919,N_1288,N_1948);
nor U4920 (N_4920,N_1485,N_822);
or U4921 (N_4921,N_2409,N_1815);
and U4922 (N_4922,N_18,N_1960);
nor U4923 (N_4923,N_3369,N_2786);
nand U4924 (N_4924,N_1157,N_1758);
xor U4925 (N_4925,N_507,N_2355);
nor U4926 (N_4926,N_2945,N_1048);
nand U4927 (N_4927,N_2769,N_3935);
xnor U4928 (N_4928,N_2044,N_3895);
and U4929 (N_4929,N_3007,N_1892);
or U4930 (N_4930,N_2665,N_3540);
xor U4931 (N_4931,N_2736,N_2152);
xnor U4932 (N_4932,N_2191,N_795);
nand U4933 (N_4933,N_3928,N_1491);
and U4934 (N_4934,N_316,N_3793);
nand U4935 (N_4935,N_2846,N_3952);
or U4936 (N_4936,N_682,N_1252);
nor U4937 (N_4937,N_3082,N_71);
or U4938 (N_4938,N_3484,N_3170);
or U4939 (N_4939,N_1975,N_1609);
nor U4940 (N_4940,N_1151,N_3798);
or U4941 (N_4941,N_569,N_3727);
or U4942 (N_4942,N_3932,N_745);
and U4943 (N_4943,N_1355,N_3446);
and U4944 (N_4944,N_1686,N_2956);
or U4945 (N_4945,N_1469,N_3638);
nand U4946 (N_4946,N_2732,N_1044);
nand U4947 (N_4947,N_1317,N_3914);
nand U4948 (N_4948,N_2965,N_1903);
and U4949 (N_4949,N_2215,N_1944);
xor U4950 (N_4950,N_2118,N_2491);
and U4951 (N_4951,N_1045,N_1591);
or U4952 (N_4952,N_2862,N_453);
nand U4953 (N_4953,N_3898,N_3882);
nand U4954 (N_4954,N_748,N_372);
or U4955 (N_4955,N_2013,N_547);
xor U4956 (N_4956,N_1842,N_1617);
nand U4957 (N_4957,N_3664,N_953);
xor U4958 (N_4958,N_3938,N_3608);
and U4959 (N_4959,N_3632,N_765);
and U4960 (N_4960,N_2666,N_2303);
xor U4961 (N_4961,N_428,N_2272);
nor U4962 (N_4962,N_3468,N_2986);
nor U4963 (N_4963,N_2735,N_2661);
nor U4964 (N_4964,N_2310,N_3432);
nor U4965 (N_4965,N_1697,N_54);
nor U4966 (N_4966,N_805,N_1767);
or U4967 (N_4967,N_943,N_2800);
xnor U4968 (N_4968,N_970,N_3885);
or U4969 (N_4969,N_3322,N_656);
or U4970 (N_4970,N_782,N_2781);
nand U4971 (N_4971,N_3795,N_1521);
nor U4972 (N_4972,N_1613,N_3777);
and U4973 (N_4973,N_1444,N_3406);
nor U4974 (N_4974,N_2396,N_1601);
nor U4975 (N_4975,N_135,N_590);
nand U4976 (N_4976,N_1622,N_921);
nand U4977 (N_4977,N_627,N_1895);
nand U4978 (N_4978,N_2601,N_2567);
nor U4979 (N_4979,N_2885,N_1868);
and U4980 (N_4980,N_3396,N_1422);
nand U4981 (N_4981,N_2320,N_2797);
xor U4982 (N_4982,N_294,N_2547);
nor U4983 (N_4983,N_2988,N_1223);
and U4984 (N_4984,N_3341,N_295);
or U4985 (N_4985,N_624,N_1614);
xor U4986 (N_4986,N_1233,N_1283);
and U4987 (N_4987,N_2763,N_2911);
nand U4988 (N_4988,N_3775,N_1932);
nand U4989 (N_4989,N_1366,N_616);
nand U4990 (N_4990,N_3552,N_455);
or U4991 (N_4991,N_1362,N_3336);
or U4992 (N_4992,N_395,N_1059);
nor U4993 (N_4993,N_3605,N_1343);
nor U4994 (N_4994,N_101,N_3792);
and U4995 (N_4995,N_2884,N_301);
xor U4996 (N_4996,N_3461,N_715);
or U4997 (N_4997,N_852,N_905);
and U4998 (N_4998,N_1629,N_3331);
and U4999 (N_4999,N_280,N_2248);
nor U5000 (N_5000,N_1389,N_2652);
nand U5001 (N_5001,N_446,N_918);
and U5002 (N_5002,N_932,N_885);
nand U5003 (N_5003,N_247,N_2255);
xnor U5004 (N_5004,N_1399,N_1553);
or U5005 (N_5005,N_2274,N_1473);
or U5006 (N_5006,N_1936,N_537);
or U5007 (N_5007,N_1152,N_111);
nor U5008 (N_5008,N_1694,N_2775);
or U5009 (N_5009,N_2804,N_1467);
and U5010 (N_5010,N_3324,N_2230);
and U5011 (N_5011,N_526,N_2697);
and U5012 (N_5012,N_1412,N_1395);
and U5013 (N_5013,N_1093,N_83);
nor U5014 (N_5014,N_270,N_2004);
xnor U5015 (N_5015,N_1934,N_3421);
and U5016 (N_5016,N_268,N_818);
xor U5017 (N_5017,N_3636,N_3616);
nand U5018 (N_5018,N_2779,N_1673);
nand U5019 (N_5019,N_1137,N_2622);
or U5020 (N_5020,N_827,N_3825);
or U5021 (N_5021,N_1906,N_483);
nor U5022 (N_5022,N_3692,N_801);
or U5023 (N_5023,N_908,N_2294);
and U5024 (N_5024,N_774,N_2410);
and U5025 (N_5025,N_928,N_1713);
nand U5026 (N_5026,N_2651,N_1736);
xnor U5027 (N_5027,N_756,N_2562);
and U5028 (N_5028,N_2605,N_1351);
nor U5029 (N_5029,N_3443,N_1209);
or U5030 (N_5030,N_487,N_3497);
nor U5031 (N_5031,N_589,N_2686);
or U5032 (N_5032,N_2701,N_2632);
or U5033 (N_5033,N_1901,N_3199);
and U5034 (N_5034,N_1785,N_3591);
nor U5035 (N_5035,N_755,N_276);
nor U5036 (N_5036,N_1040,N_687);
nor U5037 (N_5037,N_2486,N_1954);
and U5038 (N_5038,N_342,N_2959);
and U5039 (N_5039,N_3554,N_160);
and U5040 (N_5040,N_2850,N_1812);
or U5041 (N_5041,N_2892,N_1981);
xor U5042 (N_5042,N_1085,N_1078);
nor U5043 (N_5043,N_2989,N_3442);
and U5044 (N_5044,N_217,N_2437);
and U5045 (N_5045,N_2288,N_560);
nor U5046 (N_5046,N_251,N_3826);
nor U5047 (N_5047,N_3097,N_41);
nand U5048 (N_5048,N_2556,N_1232);
nand U5049 (N_5049,N_523,N_164);
or U5050 (N_5050,N_1419,N_3749);
nand U5051 (N_5051,N_1748,N_2153);
and U5052 (N_5052,N_1074,N_1075);
and U5053 (N_5053,N_212,N_3163);
or U5054 (N_5054,N_3086,N_1570);
or U5055 (N_5055,N_3741,N_1540);
xor U5056 (N_5056,N_2689,N_1620);
nor U5057 (N_5057,N_2454,N_1930);
xnor U5058 (N_5058,N_3856,N_224);
and U5059 (N_5059,N_1682,N_427);
or U5060 (N_5060,N_3229,N_2634);
nand U5061 (N_5061,N_3862,N_3437);
nand U5062 (N_5062,N_2951,N_1032);
nor U5063 (N_5063,N_219,N_830);
nor U5064 (N_5064,N_132,N_1002);
nor U5065 (N_5065,N_460,N_1648);
nor U5066 (N_5066,N_2540,N_2275);
and U5067 (N_5067,N_3858,N_2007);
nand U5068 (N_5068,N_325,N_2367);
and U5069 (N_5069,N_68,N_229);
and U5070 (N_5070,N_3607,N_1207);
or U5071 (N_5071,N_143,N_3802);
or U5072 (N_5072,N_1016,N_3073);
and U5073 (N_5073,N_1484,N_3127);
nor U5074 (N_5074,N_1114,N_2668);
nor U5075 (N_5075,N_2065,N_2231);
or U5076 (N_5076,N_1270,N_1533);
xor U5077 (N_5077,N_739,N_1850);
or U5078 (N_5078,N_3033,N_404);
nand U5079 (N_5079,N_3353,N_3017);
or U5080 (N_5080,N_1746,N_591);
or U5081 (N_5081,N_45,N_3319);
xor U5082 (N_5082,N_1544,N_1522);
or U5083 (N_5083,N_3812,N_1913);
xnor U5084 (N_5084,N_2683,N_1372);
and U5085 (N_5085,N_284,N_3681);
nand U5086 (N_5086,N_1379,N_115);
nand U5087 (N_5087,N_1832,N_2906);
nor U5088 (N_5088,N_820,N_519);
and U5089 (N_5089,N_1625,N_2963);
and U5090 (N_5090,N_3101,N_2061);
or U5091 (N_5091,N_1573,N_3271);
nor U5092 (N_5092,N_343,N_940);
and U5093 (N_5093,N_1993,N_546);
nand U5094 (N_5094,N_2311,N_1166);
and U5095 (N_5095,N_3660,N_2863);
and U5096 (N_5096,N_2183,N_1503);
nor U5097 (N_5097,N_2941,N_3709);
or U5098 (N_5098,N_205,N_152);
nor U5099 (N_5099,N_529,N_729);
and U5100 (N_5100,N_2897,N_116);
nor U5101 (N_5101,N_1398,N_679);
nor U5102 (N_5102,N_57,N_678);
and U5103 (N_5103,N_2752,N_1035);
nand U5104 (N_5104,N_3375,N_1124);
and U5105 (N_5105,N_2896,N_81);
and U5106 (N_5106,N_949,N_1921);
nor U5107 (N_5107,N_2468,N_459);
xor U5108 (N_5108,N_1587,N_3328);
nor U5109 (N_5109,N_3277,N_2565);
and U5110 (N_5110,N_2102,N_2523);
xor U5111 (N_5111,N_5,N_694);
or U5112 (N_5112,N_3072,N_1822);
or U5113 (N_5113,N_1489,N_1381);
xnor U5114 (N_5114,N_150,N_1759);
nor U5115 (N_5115,N_1254,N_1041);
or U5116 (N_5116,N_1304,N_3621);
or U5117 (N_5117,N_796,N_541);
nand U5118 (N_5118,N_2417,N_3966);
nor U5119 (N_5119,N_2430,N_1258);
xor U5120 (N_5120,N_333,N_936);
and U5121 (N_5121,N_475,N_2588);
nand U5122 (N_5122,N_3423,N_3547);
nand U5123 (N_5123,N_2663,N_3814);
or U5124 (N_5124,N_2502,N_769);
xor U5125 (N_5125,N_3223,N_3228);
and U5126 (N_5126,N_2197,N_2339);
or U5127 (N_5127,N_1649,N_3420);
xor U5128 (N_5128,N_2744,N_3904);
nand U5129 (N_5129,N_536,N_2829);
and U5130 (N_5130,N_2624,N_3186);
or U5131 (N_5131,N_3600,N_2802);
or U5132 (N_5132,N_2195,N_527);
or U5133 (N_5133,N_2982,N_1744);
or U5134 (N_5134,N_1310,N_410);
or U5135 (N_5135,N_2487,N_2090);
or U5136 (N_5136,N_1385,N_3925);
xor U5137 (N_5137,N_58,N_988);
or U5138 (N_5138,N_1520,N_1745);
nor U5139 (N_5139,N_1363,N_1884);
or U5140 (N_5140,N_735,N_3472);
nor U5141 (N_5141,N_2813,N_630);
nand U5142 (N_5142,N_1019,N_3592);
and U5143 (N_5143,N_1980,N_674);
xnor U5144 (N_5144,N_1524,N_2918);
xnor U5145 (N_5145,N_2240,N_2003);
nand U5146 (N_5146,N_2485,N_289);
nand U5147 (N_5147,N_1224,N_2893);
nor U5148 (N_5148,N_950,N_1807);
and U5149 (N_5149,N_1292,N_1293);
or U5150 (N_5150,N_2307,N_384);
nor U5151 (N_5151,N_1632,N_1219);
and U5152 (N_5152,N_499,N_1924);
and U5153 (N_5153,N_3839,N_520);
nor U5154 (N_5154,N_3249,N_3532);
and U5155 (N_5155,N_3465,N_563);
nor U5156 (N_5156,N_1862,N_2281);
or U5157 (N_5157,N_3001,N_1814);
nor U5158 (N_5158,N_3651,N_595);
and U5159 (N_5159,N_1545,N_2608);
nor U5160 (N_5160,N_3670,N_3478);
xor U5161 (N_5161,N_1911,N_2558);
nand U5162 (N_5162,N_47,N_2282);
or U5163 (N_5163,N_79,N_1927);
and U5164 (N_5164,N_1446,N_106);
nand U5165 (N_5165,N_733,N_2525);
xor U5166 (N_5166,N_1583,N_2351);
and U5167 (N_5167,N_263,N_2104);
xor U5168 (N_5168,N_1368,N_3915);
xnor U5169 (N_5169,N_1998,N_3381);
nor U5170 (N_5170,N_3728,N_2096);
nand U5171 (N_5171,N_283,N_2481);
xnor U5172 (N_5172,N_3647,N_3614);
or U5173 (N_5173,N_1267,N_1833);
or U5174 (N_5174,N_1031,N_704);
nand U5175 (N_5175,N_128,N_2138);
xnor U5176 (N_5176,N_1397,N_3851);
and U5177 (N_5177,N_552,N_2891);
and U5178 (N_5178,N_2650,N_31);
and U5179 (N_5179,N_1795,N_794);
and U5180 (N_5180,N_1042,N_1825);
and U5181 (N_5181,N_1305,N_2357);
nor U5182 (N_5182,N_3430,N_2343);
or U5183 (N_5183,N_1116,N_671);
nand U5184 (N_5184,N_2269,N_1253);
or U5185 (N_5185,N_2673,N_814);
xnor U5186 (N_5186,N_13,N_22);
or U5187 (N_5187,N_66,N_3409);
and U5188 (N_5188,N_2980,N_199);
xnor U5189 (N_5189,N_2385,N_1066);
nand U5190 (N_5190,N_1834,N_2524);
nand U5191 (N_5191,N_1966,N_2602);
xor U5192 (N_5192,N_1039,N_3242);
and U5193 (N_5193,N_2200,N_1989);
or U5194 (N_5194,N_2111,N_2380);
and U5195 (N_5195,N_2856,N_2203);
nand U5196 (N_5196,N_2018,N_2386);
nand U5197 (N_5197,N_232,N_874);
or U5198 (N_5198,N_1185,N_476);
nand U5199 (N_5199,N_2413,N_3982);
nor U5200 (N_5200,N_351,N_3945);
and U5201 (N_5201,N_3871,N_3395);
and U5202 (N_5202,N_3009,N_1992);
nand U5203 (N_5203,N_1298,N_64);
nand U5204 (N_5204,N_1723,N_850);
xnor U5205 (N_5205,N_2026,N_2455);
nand U5206 (N_5206,N_1179,N_577);
nand U5207 (N_5207,N_1017,N_1885);
nor U5208 (N_5208,N_1908,N_119);
or U5209 (N_5209,N_2193,N_1646);
nor U5210 (N_5210,N_1608,N_1693);
and U5211 (N_5211,N_690,N_2504);
and U5212 (N_5212,N_2969,N_2210);
nor U5213 (N_5213,N_3987,N_3509);
xnor U5214 (N_5214,N_2860,N_3742);
xnor U5215 (N_5215,N_605,N_210);
nand U5216 (N_5216,N_1202,N_845);
and U5217 (N_5217,N_1751,N_272);
or U5218 (N_5218,N_2167,N_871);
and U5219 (N_5219,N_1463,N_1730);
and U5220 (N_5220,N_3887,N_1325);
nor U5221 (N_5221,N_2427,N_416);
xnor U5222 (N_5222,N_368,N_2644);
or U5223 (N_5223,N_3358,N_2811);
and U5224 (N_5224,N_701,N_1905);
and U5225 (N_5225,N_1501,N_1376);
nand U5226 (N_5226,N_2833,N_1566);
and U5227 (N_5227,N_3733,N_1982);
and U5228 (N_5228,N_273,N_958);
nand U5229 (N_5229,N_2077,N_3601);
nor U5230 (N_5230,N_358,N_3436);
nand U5231 (N_5231,N_1568,N_1870);
and U5232 (N_5232,N_702,N_2546);
or U5233 (N_5233,N_1661,N_1753);
nor U5234 (N_5234,N_979,N_105);
xnor U5235 (N_5235,N_1721,N_417);
nand U5236 (N_5236,N_3356,N_1449);
or U5237 (N_5237,N_3333,N_3339);
nor U5238 (N_5238,N_357,N_32);
or U5239 (N_5239,N_3884,N_3455);
xor U5240 (N_5240,N_2318,N_3685);
nor U5241 (N_5241,N_3753,N_3577);
and U5242 (N_5242,N_2397,N_25);
or U5243 (N_5243,N_3290,N_1976);
nand U5244 (N_5244,N_628,N_1596);
or U5245 (N_5245,N_1358,N_2610);
and U5246 (N_5246,N_240,N_2704);
or U5247 (N_5247,N_2728,N_2070);
and U5248 (N_5248,N_1319,N_2719);
nor U5249 (N_5249,N_3971,N_3859);
xnor U5250 (N_5250,N_144,N_439);
nor U5251 (N_5251,N_567,N_2394);
xor U5252 (N_5252,N_1206,N_753);
or U5253 (N_5253,N_1990,N_2184);
nand U5254 (N_5254,N_1787,N_1946);
and U5255 (N_5255,N_2999,N_2370);
xor U5256 (N_5256,N_3128,N_1451);
xnor U5257 (N_5257,N_70,N_2304);
or U5258 (N_5258,N_1532,N_1534);
xnor U5259 (N_5259,N_1776,N_3281);
nand U5260 (N_5260,N_1752,N_751);
and U5261 (N_5261,N_1791,N_977);
or U5262 (N_5262,N_1212,N_2317);
nor U5263 (N_5263,N_2234,N_1429);
and U5264 (N_5264,N_817,N_996);
and U5265 (N_5265,N_3188,N_2936);
nand U5266 (N_5266,N_2729,N_3941);
and U5267 (N_5267,N_1437,N_207);
xnor U5268 (N_5268,N_1918,N_3312);
nand U5269 (N_5269,N_3796,N_3976);
and U5270 (N_5270,N_126,N_2751);
xnor U5271 (N_5271,N_2877,N_1768);
and U5272 (N_5272,N_3676,N_744);
or U5273 (N_5273,N_1240,N_1007);
or U5274 (N_5274,N_88,N_2776);
nor U5275 (N_5275,N_2467,N_2465);
and U5276 (N_5276,N_3841,N_3345);
and U5277 (N_5277,N_3235,N_2667);
xnor U5278 (N_5278,N_337,N_3014);
and U5279 (N_5279,N_3227,N_3546);
or U5280 (N_5280,N_163,N_1247);
and U5281 (N_5281,N_2677,N_2682);
nor U5282 (N_5282,N_2420,N_3500);
nand U5283 (N_5283,N_2927,N_2443);
or U5284 (N_5284,N_1430,N_2909);
and U5285 (N_5285,N_1012,N_3842);
xor U5286 (N_5286,N_2517,N_2505);
and U5287 (N_5287,N_1541,N_3213);
or U5288 (N_5288,N_1327,N_189);
nor U5289 (N_5289,N_1336,N_203);
and U5290 (N_5290,N_1855,N_3748);
xor U5291 (N_5291,N_1590,N_2154);
xor U5292 (N_5292,N_187,N_1923);
nand U5293 (N_5293,N_1172,N_3745);
nand U5294 (N_5294,N_1804,N_685);
xor U5295 (N_5295,N_3583,N_2179);
or U5296 (N_5296,N_973,N_1161);
or U5297 (N_5297,N_926,N_3354);
and U5298 (N_5298,N_449,N_3603);
or U5299 (N_5299,N_1650,N_1717);
or U5300 (N_5300,N_3157,N_78);
nor U5301 (N_5301,N_1226,N_1281);
nand U5302 (N_5302,N_1276,N_3293);
or U5303 (N_5303,N_2569,N_1675);
or U5304 (N_5304,N_642,N_3492);
or U5305 (N_5305,N_3972,N_3045);
nand U5306 (N_5306,N_3983,N_1838);
or U5307 (N_5307,N_1599,N_2952);
or U5308 (N_5308,N_2384,N_3877);
and U5309 (N_5309,N_1018,N_3219);
and U5310 (N_5310,N_2353,N_3441);
nand U5311 (N_5311,N_2784,N_100);
xor U5312 (N_5312,N_7,N_2613);
or U5313 (N_5313,N_1421,N_2387);
and U5314 (N_5314,N_3787,N_1664);
nor U5315 (N_5315,N_3563,N_3735);
and U5316 (N_5316,N_1764,N_1365);
nand U5317 (N_5317,N_3936,N_193);
xnor U5318 (N_5318,N_3192,N_2536);
nor U5319 (N_5319,N_2929,N_3291);
and U5320 (N_5320,N_2424,N_1615);
xor U5321 (N_5321,N_968,N_2796);
xnor U5322 (N_5322,N_225,N_2534);
nand U5323 (N_5323,N_2760,N_2079);
and U5324 (N_5324,N_108,N_1678);
xnor U5325 (N_5325,N_2477,N_3307);
xor U5326 (N_5326,N_1701,N_3308);
or U5327 (N_5327,N_664,N_3924);
xor U5328 (N_5328,N_2262,N_1004);
nand U5329 (N_5329,N_3533,N_2901);
xnor U5330 (N_5330,N_3036,N_75);
and U5331 (N_5331,N_1309,N_521);
and U5332 (N_5332,N_3764,N_1050);
or U5333 (N_5333,N_1623,N_2659);
or U5334 (N_5334,N_3535,N_2433);
or U5335 (N_5335,N_2961,N_1508);
nor U5336 (N_5336,N_999,N_1703);
and U5337 (N_5337,N_3979,N_3405);
and U5338 (N_5338,N_2563,N_3305);
and U5339 (N_5339,N_3784,N_1203);
xnor U5340 (N_5340,N_3909,N_1217);
xor U5341 (N_5341,N_3807,N_3018);
or U5342 (N_5342,N_816,N_2029);
nor U5343 (N_5343,N_1557,N_717);
xor U5344 (N_5344,N_2457,N_3576);
nor U5345 (N_5345,N_843,N_841);
and U5346 (N_5346,N_1105,N_1840);
nor U5347 (N_5347,N_3879,N_3886);
xnor U5348 (N_5348,N_2593,N_1931);
xnor U5349 (N_5349,N_461,N_3994);
nor U5350 (N_5350,N_2233,N_3092);
nor U5351 (N_5351,N_819,N_2112);
nor U5352 (N_5352,N_1779,N_2590);
and U5353 (N_5353,N_3776,N_1415);
nand U5354 (N_5354,N_1418,N_3201);
xor U5355 (N_5355,N_1872,N_2146);
and U5356 (N_5356,N_2631,N_1388);
nor U5357 (N_5357,N_2071,N_3096);
or U5358 (N_5358,N_2283,N_258);
and U5359 (N_5359,N_3326,N_1801);
and U5360 (N_5360,N_1546,N_1401);
nand U5361 (N_5361,N_431,N_3167);
nand U5362 (N_5362,N_3855,N_2772);
and U5363 (N_5363,N_1851,N_2817);
and U5364 (N_5364,N_1020,N_1715);
and U5365 (N_5365,N_2793,N_2526);
or U5366 (N_5366,N_245,N_3504);
xor U5367 (N_5367,N_2160,N_3230);
or U5368 (N_5368,N_1071,N_2260);
nor U5369 (N_5369,N_1741,N_1330);
nor U5370 (N_5370,N_2000,N_2213);
or U5371 (N_5371,N_1010,N_2361);
xnor U5372 (N_5372,N_181,N_1225);
xor U5373 (N_5373,N_2423,N_2730);
or U5374 (N_5374,N_614,N_1977);
and U5375 (N_5375,N_2039,N_260);
or U5376 (N_5376,N_3388,N_2706);
xnor U5377 (N_5377,N_1384,N_1462);
xnor U5378 (N_5378,N_1269,N_359);
nor U5379 (N_5379,N_3587,N_3808);
and U5380 (N_5380,N_2017,N_2100);
nor U5381 (N_5381,N_1174,N_3538);
or U5382 (N_5382,N_2834,N_1618);
nand U5383 (N_5383,N_1344,N_872);
or U5384 (N_5384,N_1328,N_2177);
nand U5385 (N_5385,N_2425,N_810);
xor U5386 (N_5386,N_1196,N_2583);
nand U5387 (N_5387,N_120,N_3134);
nor U5388 (N_5388,N_3351,N_16);
xor U5389 (N_5389,N_2440,N_26);
nor U5390 (N_5390,N_3207,N_2224);
xor U5391 (N_5391,N_3716,N_898);
and U5392 (N_5392,N_2219,N_1674);
nor U5393 (N_5393,N_2552,N_389);
xnor U5394 (N_5394,N_501,N_1761);
nand U5395 (N_5395,N_524,N_1516);
nor U5396 (N_5396,N_1991,N_1468);
or U5397 (N_5397,N_823,N_3039);
nor U5398 (N_5398,N_3160,N_1643);
or U5399 (N_5399,N_1061,N_3917);
nand U5400 (N_5400,N_42,N_1654);
xor U5401 (N_5401,N_55,N_3493);
or U5402 (N_5402,N_3652,N_1013);
and U5403 (N_5403,N_103,N_2978);
xor U5404 (N_5404,N_1416,N_3248);
xor U5405 (N_5405,N_3625,N_1816);
or U5406 (N_5406,N_2853,N_741);
xor U5407 (N_5407,N_1466,N_548);
nor U5408 (N_5408,N_133,N_2570);
nand U5409 (N_5409,N_944,N_3452);
nor U5410 (N_5410,N_1616,N_2881);
or U5411 (N_5411,N_249,N_1819);
and U5412 (N_5412,N_1700,N_516);
and U5413 (N_5413,N_3978,N_2326);
nor U5414 (N_5414,N_17,N_2528);
xor U5415 (N_5415,N_2223,N_1718);
nand U5416 (N_5416,N_14,N_2400);
and U5417 (N_5417,N_2267,N_1780);
nand U5418 (N_5418,N_3146,N_253);
nand U5419 (N_5419,N_3766,N_403);
nor U5420 (N_5420,N_1986,N_1755);
or U5421 (N_5421,N_789,N_3083);
and U5422 (N_5422,N_1479,N_2842);
nand U5423 (N_5423,N_1475,N_3057);
nand U5424 (N_5424,N_2620,N_223);
nor U5425 (N_5425,N_3837,N_1929);
nor U5426 (N_5426,N_175,N_236);
nand U5427 (N_5427,N_1329,N_3210);
nand U5428 (N_5428,N_2649,N_3785);
and U5429 (N_5429,N_3854,N_107);
nor U5430 (N_5430,N_1722,N_3098);
and U5431 (N_5431,N_513,N_2022);
and U5432 (N_5432,N_96,N_486);
xnor U5433 (N_5433,N_3730,N_1707);
or U5434 (N_5434,N_3011,N_3453);
and U5435 (N_5435,N_2023,N_3211);
xnor U5436 (N_5436,N_170,N_570);
nand U5437 (N_5437,N_3797,N_1423);
xor U5438 (N_5438,N_2532,N_432);
nand U5439 (N_5439,N_719,N_1211);
nand U5440 (N_5440,N_3719,N_1488);
nor U5441 (N_5441,N_3703,N_1015);
xor U5442 (N_5442,N_1117,N_2939);
or U5443 (N_5443,N_2123,N_1132);
xor U5444 (N_5444,N_2399,N_3145);
or U5445 (N_5445,N_582,N_2955);
nand U5446 (N_5446,N_1088,N_1687);
or U5447 (N_5447,N_3809,N_183);
nand U5448 (N_5448,N_3519,N_1110);
nor U5449 (N_5449,N_471,N_2054);
xor U5450 (N_5450,N_3022,N_2450);
nand U5451 (N_5451,N_1864,N_114);
nor U5452 (N_5452,N_1331,N_631);
or U5453 (N_5453,N_1773,N_3857);
xnor U5454 (N_5454,N_1273,N_1346);
xnor U5455 (N_5455,N_346,N_2553);
nor U5456 (N_5456,N_3721,N_1858);
xor U5457 (N_5457,N_1699,N_1126);
xor U5458 (N_5458,N_3304,N_1456);
or U5459 (N_5459,N_607,N_2688);
nand U5460 (N_5460,N_3820,N_2687);
and U5461 (N_5461,N_1290,N_2171);
and U5462 (N_5462,N_3403,N_749);
and U5463 (N_5463,N_1435,N_1158);
xor U5464 (N_5464,N_3712,N_2799);
xnor U5465 (N_5465,N_832,N_360);
nor U5466 (N_5466,N_3921,N_790);
or U5467 (N_5467,N_2981,N_3195);
or U5468 (N_5468,N_1907,N_3575);
and U5469 (N_5469,N_914,N_1490);
nor U5470 (N_5470,N_2312,N_1406);
or U5471 (N_5471,N_2300,N_2522);
and U5472 (N_5472,N_139,N_1737);
and U5473 (N_5473,N_300,N_3829);
nand U5474 (N_5474,N_2095,N_974);
and U5475 (N_5475,N_3372,N_2794);
and U5476 (N_5476,N_1005,N_3908);
or U5477 (N_5477,N_909,N_828);
nand U5478 (N_5478,N_4,N_2199);
xor U5479 (N_5479,N_1995,N_1968);
or U5480 (N_5480,N_683,N_3080);
nand U5481 (N_5481,N_2867,N_377);
xor U5482 (N_5482,N_2890,N_2723);
nand U5483 (N_5483,N_1725,N_2010);
or U5484 (N_5484,N_991,N_866);
xor U5485 (N_5485,N_3973,N_952);
xnor U5486 (N_5486,N_3962,N_2954);
nand U5487 (N_5487,N_641,N_2406);
nand U5488 (N_5488,N_1750,N_1477);
and U5489 (N_5489,N_1069,N_441);
xor U5490 (N_5490,N_1823,N_2009);
xnor U5491 (N_5491,N_2611,N_2151);
and U5492 (N_5492,N_3761,N_2092);
or U5493 (N_5493,N_1502,N_2016);
nor U5494 (N_5494,N_775,N_3030);
and U5495 (N_5495,N_2122,N_984);
nand U5496 (N_5496,N_3175,N_3650);
and U5497 (N_5497,N_230,N_2514);
and U5498 (N_5498,N_340,N_444);
xor U5499 (N_5499,N_2946,N_1229);
xor U5500 (N_5500,N_2144,N_3371);
or U5501 (N_5501,N_1668,N_3380);
xor U5502 (N_5502,N_1168,N_3232);
nor U5503 (N_5503,N_2765,N_2561);
nor U5504 (N_5504,N_868,N_407);
nand U5505 (N_5505,N_2155,N_1113);
nor U5506 (N_5506,N_2126,N_2188);
or U5507 (N_5507,N_875,N_736);
nand U5508 (N_5508,N_1604,N_1371);
nand U5509 (N_5509,N_3852,N_2971);
xor U5510 (N_5510,N_3618,N_1987);
xnor U5511 (N_5511,N_3656,N_511);
xnor U5512 (N_5512,N_922,N_3610);
nor U5513 (N_5513,N_447,N_697);
nor U5514 (N_5514,N_498,N_488);
nor U5515 (N_5515,N_2398,N_2134);
and U5516 (N_5516,N_1881,N_3370);
xor U5517 (N_5517,N_566,N_3918);
nand U5518 (N_5518,N_2036,N_725);
nand U5519 (N_5519,N_651,N_1338);
or U5520 (N_5520,N_2129,N_1296);
xor U5521 (N_5521,N_955,N_3063);
nor U5522 (N_5522,N_3633,N_2178);
nor U5523 (N_5523,N_1139,N_2773);
nor U5524 (N_5524,N_646,N_3597);
xnor U5525 (N_5525,N_3919,N_2630);
or U5526 (N_5526,N_1313,N_92);
xnor U5527 (N_5527,N_1201,N_1320);
nand U5528 (N_5528,N_2263,N_1789);
nand U5529 (N_5529,N_1420,N_2788);
nor U5530 (N_5530,N_2785,N_1951);
and U5531 (N_5531,N_712,N_2408);
xor U5532 (N_5532,N_3836,N_2336);
nand U5533 (N_5533,N_2587,N_2462);
xnor U5534 (N_5534,N_122,N_951);
or U5535 (N_5535,N_1997,N_40);
nand U5536 (N_5536,N_2548,N_1090);
or U5537 (N_5537,N_157,N_603);
nand U5538 (N_5538,N_378,N_663);
and U5539 (N_5539,N_1064,N_2840);
nor U5540 (N_5540,N_1457,N_2338);
nor U5541 (N_5541,N_946,N_3630);
and U5542 (N_5542,N_3589,N_586);
and U5543 (N_5543,N_2672,N_3218);
or U5544 (N_5544,N_385,N_2372);
xor U5545 (N_5545,N_594,N_1262);
nand U5546 (N_5546,N_892,N_2603);
and U5547 (N_5547,N_2254,N_597);
xor U5548 (N_5548,N_539,N_746);
or U5549 (N_5549,N_2638,N_3980);
nor U5550 (N_5550,N_1408,N_506);
nand U5551 (N_5551,N_1326,N_1681);
and U5552 (N_5552,N_1130,N_2575);
or U5553 (N_5553,N_3737,N_3513);
and U5554 (N_5554,N_3612,N_1234);
or U5555 (N_5555,N_1528,N_1195);
xnor U5556 (N_5556,N_660,N_3545);
and U5557 (N_5557,N_2211,N_1178);
nand U5558 (N_5558,N_1237,N_2507);
xor U5559 (N_5559,N_2365,N_2942);
and U5560 (N_5560,N_3143,N_698);
or U5561 (N_5561,N_1142,N_1332);
nor U5562 (N_5562,N_966,N_1775);
xnor U5563 (N_5563,N_803,N_2324);
nor U5564 (N_5564,N_2887,N_3257);
xor U5565 (N_5565,N_2416,N_3089);
xnor U5566 (N_5566,N_764,N_1092);
nand U5567 (N_5567,N_3173,N_2198);
and U5568 (N_5568,N_3284,N_1060);
xnor U5569 (N_5569,N_760,N_3233);
or U5570 (N_5570,N_3594,N_456);
xnor U5571 (N_5571,N_1512,N_233);
or U5572 (N_5572,N_3042,N_3684);
nor U5573 (N_5573,N_2904,N_3751);
nand U5574 (N_5574,N_2543,N_156);
nor U5575 (N_5575,N_234,N_1055);
nand U5576 (N_5576,N_957,N_1282);
nor U5577 (N_5577,N_2855,N_1511);
xnor U5578 (N_5578,N_855,N_2466);
nor U5579 (N_5579,N_1104,N_1448);
or U5580 (N_5580,N_2374,N_3970);
or U5581 (N_5581,N_669,N_3560);
nand U5582 (N_5582,N_515,N_2280);
nand U5583 (N_5583,N_1529,N_525);
and U5584 (N_5584,N_3790,N_1708);
nand U5585 (N_5585,N_1492,N_1357);
and U5586 (N_5586,N_2005,N_3881);
or U5587 (N_5587,N_3275,N_1719);
nor U5588 (N_5588,N_3306,N_3144);
nand U5589 (N_5589,N_1026,N_2935);
xor U5590 (N_5590,N_1575,N_3172);
and U5591 (N_5591,N_1637,N_3103);
or U5592 (N_5592,N_329,N_1001);
and U5593 (N_5593,N_3590,N_672);
and U5594 (N_5594,N_562,N_3845);
and U5595 (N_5595,N_969,N_2253);
and U5596 (N_5596,N_1111,N_3959);
and U5597 (N_5597,N_3662,N_584);
nand U5598 (N_5598,N_3699,N_1558);
nor U5599 (N_5599,N_2990,N_659);
nand U5600 (N_5600,N_3071,N_3527);
or U5601 (N_5601,N_1101,N_3046);
and U5602 (N_5602,N_2947,N_1882);
nand U5603 (N_5603,N_625,N_180);
nor U5604 (N_5604,N_3995,N_334);
nor U5605 (N_5605,N_3378,N_3220);
nor U5606 (N_5606,N_51,N_2176);
nand U5607 (N_5607,N_3155,N_3865);
or U5608 (N_5608,N_338,N_2615);
nor U5609 (N_5609,N_1788,N_2472);
nor U5610 (N_5610,N_1063,N_2119);
nor U5611 (N_5611,N_1128,N_3788);
nor U5612 (N_5612,N_491,N_1985);
xor U5613 (N_5613,N_1188,N_2064);
nor U5614 (N_5614,N_1280,N_3006);
xnor U5615 (N_5615,N_931,N_462);
xnor U5616 (N_5616,N_2329,N_3515);
and U5617 (N_5617,N_1133,N_1883);
nor U5618 (N_5618,N_849,N_3985);
nor U5619 (N_5619,N_3168,N_27);
nand U5620 (N_5620,N_2845,N_1180);
nor U5621 (N_5621,N_2931,N_540);
nor U5622 (N_5622,N_3074,N_1347);
nor U5623 (N_5623,N_696,N_2055);
or U5624 (N_5624,N_2898,N_602);
and U5625 (N_5625,N_2930,N_2364);
nor U5626 (N_5626,N_2824,N_2538);
and U5627 (N_5627,N_3661,N_3427);
nand U5628 (N_5628,N_158,N_1582);
nand U5629 (N_5629,N_754,N_259);
nor U5630 (N_5630,N_2617,N_2354);
or U5631 (N_5631,N_867,N_2759);
and U5632 (N_5632,N_721,N_3140);
or U5633 (N_5633,N_1118,N_383);
or U5634 (N_5634,N_593,N_3285);
xor U5635 (N_5635,N_451,N_426);
and U5636 (N_5636,N_3847,N_3294);
nand U5637 (N_5637,N_2832,N_1470);
xnor U5638 (N_5638,N_98,N_2876);
or U5639 (N_5639,N_1455,N_2753);
nor U5640 (N_5640,N_1321,N_3384);
or U5641 (N_5641,N_3482,N_2042);
xor U5642 (N_5642,N_1714,N_2352);
nand U5643 (N_5643,N_834,N_154);
nor U5644 (N_5644,N_23,N_600);
or U5645 (N_5645,N_2076,N_3125);
nand U5646 (N_5646,N_2520,N_1844);
nand U5647 (N_5647,N_846,N_906);
or U5648 (N_5648,N_611,N_3104);
xor U5649 (N_5649,N_3325,N_1417);
nor U5650 (N_5650,N_155,N_2973);
nand U5651 (N_5651,N_2852,N_3989);
nand U5652 (N_5652,N_3892,N_3348);
nand U5653 (N_5653,N_3471,N_2012);
or U5654 (N_5654,N_474,N_3604);
xnor U5655 (N_5655,N_2826,N_3385);
nand U5656 (N_5656,N_1863,N_1414);
nand U5657 (N_5657,N_2058,N_1866);
nor U5658 (N_5658,N_172,N_1581);
xnor U5659 (N_5659,N_2460,N_3673);
and U5660 (N_5660,N_1265,N_1342);
or U5661 (N_5661,N_3449,N_2658);
and U5662 (N_5662,N_2792,N_493);
nor U5663 (N_5663,N_2120,N_3133);
or U5664 (N_5664,N_354,N_265);
or U5665 (N_5665,N_3479,N_3236);
nand U5666 (N_5666,N_2290,N_2360);
nor U5667 (N_5667,N_2072,N_3631);
or U5668 (N_5668,N_3278,N_1652);
and U5669 (N_5669,N_2492,N_1096);
nand U5670 (N_5670,N_3791,N_941);
nor U5671 (N_5671,N_3539,N_1953);
xnor U5672 (N_5672,N_1056,N_2874);
nand U5673 (N_5673,N_1380,N_248);
and U5674 (N_5674,N_1215,N_1663);
or U5675 (N_5675,N_1378,N_1145);
nand U5676 (N_5676,N_964,N_2997);
nand U5677 (N_5677,N_3399,N_1772);
xor U5678 (N_5678,N_421,N_457);
or U5679 (N_5679,N_3569,N_3992);
xnor U5680 (N_5680,N_2463,N_3682);
and U5681 (N_5681,N_670,N_3891);
nor U5682 (N_5682,N_2285,N_545);
nand U5683 (N_5683,N_136,N_743);
and U5684 (N_5684,N_1120,N_2604);
xor U5685 (N_5685,N_3967,N_2882);
nand U5686 (N_5686,N_2592,N_3118);
nor U5687 (N_5687,N_1706,N_2664);
nor U5688 (N_5688,N_3549,N_3272);
or U5689 (N_5689,N_1704,N_261);
xor U5690 (N_5690,N_3397,N_1794);
and U5691 (N_5691,N_231,N_2434);
nand U5692 (N_5692,N_882,N_2541);
xor U5693 (N_5693,N_153,N_3491);
nor U5694 (N_5694,N_367,N_2189);
xnor U5695 (N_5695,N_2412,N_645);
and U5696 (N_5696,N_400,N_3562);
or U5697 (N_5697,N_3708,N_2712);
or U5698 (N_5698,N_737,N_3687);
and U5699 (N_5699,N_2545,N_869);
nor U5700 (N_5700,N_445,N_44);
nand U5701 (N_5701,N_401,N_2726);
nor U5702 (N_5702,N_620,N_1585);
nand U5703 (N_5703,N_3161,N_1190);
nor U5704 (N_5704,N_2949,N_3024);
xnor U5705 (N_5705,N_1543,N_72);
or U5706 (N_5706,N_2750,N_1129);
or U5707 (N_5707,N_2979,N_87);
nor U5708 (N_5708,N_3274,N_370);
nand U5709 (N_5709,N_102,N_1121);
xor U5710 (N_5710,N_1955,N_503);
or U5711 (N_5711,N_2883,N_1239);
nand U5712 (N_5712,N_1199,N_2130);
xor U5713 (N_5713,N_1210,N_587);
and U5714 (N_5714,N_214,N_2585);
or U5715 (N_5715,N_3517,N_3196);
or U5716 (N_5716,N_2296,N_3832);
nand U5717 (N_5717,N_1796,N_3626);
or U5718 (N_5718,N_2618,N_1091);
xnor U5719 (N_5719,N_3878,N_1859);
or U5720 (N_5720,N_3689,N_3643);
and U5721 (N_5721,N_856,N_1054);
xnor U5722 (N_5722,N_3091,N_1561);
xor U5723 (N_5723,N_939,N_2691);
xnor U5724 (N_5724,N_448,N_1676);
or U5725 (N_5725,N_2057,N_668);
nor U5726 (N_5726,N_262,N_3999);
or U5727 (N_5727,N_1920,N_3872);
or U5728 (N_5728,N_2045,N_1810);
and U5729 (N_5729,N_3283,N_1647);
xor U5730 (N_5730,N_1891,N_376);
and U5731 (N_5731,N_1523,N_141);
nand U5732 (N_5732,N_1452,N_1067);
nand U5733 (N_5733,N_1732,N_266);
xor U5734 (N_5734,N_2393,N_606);
or U5735 (N_5735,N_375,N_1877);
nor U5736 (N_5736,N_1333,N_2173);
and U5737 (N_5737,N_2996,N_538);
or U5738 (N_5738,N_2403,N_927);
or U5739 (N_5739,N_2149,N_1808);
nor U5740 (N_5740,N_1307,N_2432);
and U5741 (N_5741,N_3683,N_1846);
nand U5742 (N_5742,N_2870,N_1375);
nor U5743 (N_5743,N_3611,N_118);
and U5744 (N_5744,N_2,N_3930);
nand U5745 (N_5745,N_1043,N_870);
or U5746 (N_5746,N_2069,N_2671);
nand U5747 (N_5747,N_252,N_1509);
nand U5748 (N_5748,N_3475,N_2544);
nand U5749 (N_5749,N_2783,N_2866);
and U5750 (N_5750,N_1879,N_3769);
or U5751 (N_5751,N_2098,N_1959);
nand U5752 (N_5752,N_2571,N_1957);
xor U5753 (N_5753,N_1961,N_2159);
nor U5754 (N_5754,N_1303,N_3723);
and U5755 (N_5755,N_1314,N_692);
nor U5756 (N_5756,N_1651,N_667);
or U5757 (N_5757,N_1164,N_3193);
nand U5758 (N_5758,N_3241,N_2322);
nor U5759 (N_5759,N_861,N_422);
xnor U5760 (N_5760,N_3450,N_718);
xnor U5761 (N_5761,N_3300,N_179);
nand U5762 (N_5762,N_3706,N_3774);
or U5763 (N_5763,N_1684,N_2428);
or U5764 (N_5764,N_1669,N_369);
xor U5765 (N_5765,N_3049,N_2298);
nand U5766 (N_5766,N_1658,N_3489);
nand U5767 (N_5767,N_1354,N_3655);
xnor U5768 (N_5768,N_500,N_2818);
and U5769 (N_5769,N_2494,N_1189);
or U5770 (N_5770,N_2166,N_1339);
or U5771 (N_5771,N_2654,N_3451);
and U5772 (N_5772,N_784,N_2993);
xnor U5773 (N_5773,N_3268,N_1115);
and U5774 (N_5774,N_3387,N_2313);
xor U5775 (N_5775,N_2441,N_2220);
nor U5776 (N_5776,N_3522,N_2669);
and U5777 (N_5777,N_771,N_714);
nor U5778 (N_5778,N_2976,N_1818);
nand U5779 (N_5779,N_3645,N_2446);
or U5780 (N_5780,N_145,N_2530);
or U5781 (N_5781,N_3747,N_2139);
nor U5782 (N_5782,N_838,N_1183);
nor U5783 (N_5783,N_348,N_1482);
and U5784 (N_5784,N_2635,N_1641);
and U5785 (N_5785,N_2257,N_2674);
xor U5786 (N_5786,N_3311,N_1155);
nand U5787 (N_5787,N_1640,N_3263);
and U5788 (N_5788,N_783,N_3998);
nand U5789 (N_5789,N_1394,N_2245);
xnor U5790 (N_5790,N_2308,N_1688);
nand U5791 (N_5791,N_2249,N_3255);
nand U5792 (N_5792,N_2276,N_1443);
xnor U5793 (N_5793,N_3593,N_896);
nand U5794 (N_5794,N_2764,N_2515);
nor U5795 (N_5795,N_3287,N_1845);
or U5796 (N_5796,N_2107,N_113);
and U5797 (N_5797,N_1149,N_3439);
nor U5798 (N_5798,N_948,N_599);
and U5799 (N_5799,N_2411,N_860);
nor U5800 (N_5800,N_373,N_2509);
nor U5801 (N_5801,N_3323,N_1476);
xnor U5802 (N_5802,N_637,N_3122);
xor U5803 (N_5803,N_3418,N_3376);
or U5804 (N_5804,N_1829,N_2584);
nor U5805 (N_5805,N_3880,N_555);
nor U5806 (N_5806,N_3126,N_772);
xor U5807 (N_5807,N_1595,N_1436);
xor U5808 (N_5808,N_3416,N_1910);
xor U5809 (N_5809,N_3690,N_919);
or U5810 (N_5810,N_3659,N_2974);
or U5811 (N_5811,N_2442,N_239);
nand U5812 (N_5812,N_517,N_1562);
nand U5813 (N_5813,N_3634,N_3642);
nand U5814 (N_5814,N_2740,N_777);
or U5815 (N_5815,N_2619,N_1733);
or U5816 (N_5816,N_990,N_3669);
nor U5817 (N_5817,N_497,N_3295);
nor U5818 (N_5818,N_2132,N_2125);
nor U5819 (N_5819,N_2985,N_3460);
or U5820 (N_5820,N_532,N_666);
nor U5821 (N_5821,N_786,N_738);
nor U5822 (N_5822,N_161,N_601);
or U5823 (N_5823,N_2805,N_3110);
xor U5824 (N_5824,N_3185,N_308);
nor U5825 (N_5825,N_3357,N_2722);
nand U5826 (N_5826,N_2770,N_2747);
nand U5827 (N_5827,N_1984,N_3813);
and U5828 (N_5828,N_884,N_3150);
xor U5829 (N_5829,N_2731,N_3588);
nand U5830 (N_5830,N_3078,N_314);
and U5831 (N_5831,N_1404,N_881);
and U5832 (N_5832,N_2616,N_3114);
nor U5833 (N_5833,N_3251,N_2879);
nand U5834 (N_5834,N_2694,N_3123);
nor U5835 (N_5835,N_1131,N_382);
nand U5836 (N_5836,N_3680,N_1334);
and U5837 (N_5837,N_59,N_1014);
nand U5838 (N_5838,N_1370,N_1689);
nand U5839 (N_5839,N_117,N_2568);
nand U5840 (N_5840,N_1740,N_2378);
nor U5841 (N_5841,N_1774,N_3401);
or U5842 (N_5842,N_2537,N_1602);
xor U5843 (N_5843,N_65,N_1527);
nor U5844 (N_5844,N_364,N_1426);
and U5845 (N_5845,N_3899,N_481);
or U5846 (N_5846,N_379,N_2953);
xnor U5847 (N_5847,N_2580,N_380);
nand U5848 (N_5848,N_2707,N_3986);
and U5849 (N_5849,N_913,N_3665);
or U5850 (N_5850,N_3619,N_3707);
nor U5851 (N_5851,N_3108,N_2713);
nor U5852 (N_5852,N_2135,N_1969);
nor U5853 (N_5853,N_3070,N_3890);
nor U5854 (N_5854,N_1028,N_681);
nor U5855 (N_5855,N_2228,N_1033);
xnor U5856 (N_5856,N_1038,N_509);
xor U5857 (N_5857,N_3675,N_676);
xnor U5858 (N_5858,N_2221,N_2972);
nor U5859 (N_5859,N_3580,N_2835);
and U5860 (N_5860,N_3518,N_2869);
nand U5861 (N_5861,N_1461,N_3732);
nor U5862 (N_5862,N_480,N_837);
nor U5863 (N_5863,N_2229,N_3582);
nor U5864 (N_5864,N_12,N_1068);
and U5865 (N_5865,N_3701,N_1125);
or U5866 (N_5866,N_3704,N_1369);
and U5867 (N_5867,N_2084,N_3772);
nand U5868 (N_5868,N_3026,N_3084);
or U5869 (N_5869,N_2680,N_3280);
nor U5870 (N_5870,N_636,N_2577);
nand U5871 (N_5871,N_3261,N_1160);
nand U5872 (N_5872,N_1083,N_3516);
nor U5873 (N_5873,N_2801,N_3273);
nor U5874 (N_5874,N_2237,N_2348);
nand U5875 (N_5875,N_2754,N_864);
nor U5876 (N_5876,N_1513,N_121);
or U5877 (N_5877,N_1411,N_3831);
xor U5878 (N_5878,N_1677,N_3373);
nor U5879 (N_5879,N_2327,N_1300);
xor U5880 (N_5880,N_2926,N_3176);
and U5881 (N_5881,N_3166,N_2660);
nor U5882 (N_5882,N_1141,N_1627);
and U5883 (N_5883,N_3810,N_1666);
or U5884 (N_5884,N_613,N_3961);
nor U5885 (N_5885,N_851,N_3330);
xor U5886 (N_5886,N_2912,N_1803);
xor U5887 (N_5887,N_1377,N_2823);
nor U5888 (N_5888,N_3731,N_1077);
or U5889 (N_5889,N_2639,N_2756);
and U5890 (N_5890,N_981,N_1208);
nor U5891 (N_5891,N_3824,N_1);
or U5892 (N_5892,N_1465,N_1493);
or U5893 (N_5893,N_3379,N_3543);
nand U5894 (N_5894,N_650,N_1458);
nand U5895 (N_5895,N_2700,N_110);
nand U5896 (N_5896,N_1734,N_661);
xor U5897 (N_5897,N_2703,N_1867);
xnor U5898 (N_5898,N_853,N_191);
nor U5899 (N_5899,N_3456,N_3056);
xor U5900 (N_5900,N_1441,N_3816);
xor U5901 (N_5901,N_2574,N_3262);
or U5902 (N_5902,N_85,N_2595);
nor U5903 (N_5903,N_2737,N_3250);
and U5904 (N_5904,N_3310,N_779);
or U5905 (N_5905,N_1192,N_3000);
and U5906 (N_5906,N_839,N_572);
and U5907 (N_5907,N_963,N_2375);
and U5908 (N_5908,N_3142,N_1102);
nor U5909 (N_5909,N_706,N_2925);
nor U5910 (N_5910,N_2757,N_2789);
or U5911 (N_5911,N_2404,N_3487);
xnor U5912 (N_5912,N_1176,N_1743);
nand U5913 (N_5913,N_2807,N_438);
or U5914 (N_5914,N_2960,N_2539);
nand U5915 (N_5915,N_3942,N_1777);
and U5916 (N_5916,N_2966,N_2316);
or U5917 (N_5917,N_2143,N_1352);
nor U5918 (N_5918,N_478,N_724);
nor U5919 (N_5919,N_3474,N_1081);
nor U5920 (N_5920,N_2043,N_2110);
or U5921 (N_5921,N_3355,N_2182);
nor U5922 (N_5922,N_238,N_693);
or U5923 (N_5923,N_2967,N_3902);
nor U5924 (N_5924,N_634,N_3343);
or U5925 (N_5925,N_222,N_723);
and U5926 (N_5926,N_1175,N_386);
and U5927 (N_5927,N_3079,N_3363);
or U5928 (N_5928,N_1494,N_3548);
or U5929 (N_5929,N_3105,N_1316);
nor U5930 (N_5930,N_3541,N_3404);
nand U5931 (N_5931,N_3755,N_1837);
and U5932 (N_5932,N_1383,N_2247);
nand U5933 (N_5933,N_1983,N_46);
xor U5934 (N_5934,N_3434,N_235);
nor U5935 (N_5935,N_3501,N_19);
and U5936 (N_5936,N_2733,N_82);
or U5937 (N_5937,N_2943,N_2418);
xnor U5938 (N_5938,N_3654,N_2843);
nor U5939 (N_5939,N_3875,N_3609);
xor U5940 (N_5940,N_1360,N_409);
and U5941 (N_5941,N_1245,N_857);
and U5942 (N_5942,N_3752,N_2222);
xnor U5943 (N_5943,N_2172,N_109);
xnor U5944 (N_5944,N_1904,N_3564);
xnor U5945 (N_5945,N_2251,N_1958);
or U5946 (N_5946,N_1231,N_3738);
nor U5947 (N_5947,N_3190,N_652);
and U5948 (N_5948,N_1084,N_598);
xor U5949 (N_5949,N_282,N_3221);
nand U5950 (N_5950,N_3916,N_3012);
and U5951 (N_5951,N_406,N_2334);
xnor U5952 (N_5952,N_479,N_2368);
nand U5953 (N_5953,N_1765,N_2924);
or U5954 (N_5954,N_2168,N_1593);
or U5955 (N_5955,N_3584,N_3617);
nand U5956 (N_5956,N_573,N_2150);
and U5957 (N_5957,N_2345,N_2646);
nor U5958 (N_5958,N_1922,N_2456);
xnor U5959 (N_5959,N_3762,N_1894);
nor U5960 (N_5960,N_3008,N_2405);
nor U5961 (N_5961,N_1097,N_1349);
and U5962 (N_5962,N_3444,N_3164);
nor U5963 (N_5963,N_311,N_2242);
nor U5964 (N_5964,N_1760,N_2145);
or U5965 (N_5965,N_324,N_1187);
nand U5966 (N_5966,N_2848,N_2476);
and U5967 (N_5967,N_543,N_3602);
or U5968 (N_5968,N_3984,N_3415);
or U5969 (N_5969,N_3389,N_67);
nor U5970 (N_5970,N_177,N_3428);
xor U5971 (N_5971,N_2878,N_2812);
nand U5972 (N_5972,N_412,N_3226);
nand U5973 (N_5973,N_3021,N_1073);
nor U5974 (N_5974,N_883,N_3671);
and U5975 (N_5975,N_396,N_1555);
xnor U5976 (N_5976,N_2464,N_3417);
nand U5977 (N_5977,N_166,N_3054);
nand U5978 (N_5978,N_2519,N_3649);
nor U5979 (N_5979,N_848,N_2868);
xnor U5980 (N_5980,N_930,N_2227);
xor U5981 (N_5981,N_2629,N_3780);
nor U5982 (N_5982,N_2557,N_2190);
xnor U5983 (N_5983,N_2653,N_2521);
or U5984 (N_5984,N_1079,N_3947);
or U5985 (N_5985,N_3424,N_3055);
and U5986 (N_5986,N_2576,N_2302);
and U5987 (N_5987,N_3067,N_1098);
nor U5988 (N_5988,N_1464,N_2838);
nand U5989 (N_5989,N_1499,N_10);
nand U5990 (N_5990,N_684,N_578);
xnor U5991 (N_5991,N_3901,N_1204);
or U5992 (N_5992,N_2137,N_960);
or U5993 (N_5993,N_1340,N_3555);
xor U5994 (N_5994,N_52,N_1496);
xnor U5995 (N_5995,N_3206,N_924);
or U5996 (N_5996,N_1949,N_3977);
nand U5997 (N_5997,N_840,N_1181);
and U5998 (N_5998,N_505,N_2531);
and U5999 (N_5999,N_2266,N_390);
xnor U6000 (N_6000,N_903,N_1280);
or U6001 (N_6001,N_3707,N_895);
nor U6002 (N_6002,N_1298,N_126);
and U6003 (N_6003,N_2565,N_2902);
xnor U6004 (N_6004,N_269,N_3322);
nand U6005 (N_6005,N_1270,N_1357);
or U6006 (N_6006,N_1210,N_1647);
or U6007 (N_6007,N_1271,N_3544);
nor U6008 (N_6008,N_1983,N_3096);
or U6009 (N_6009,N_1545,N_3200);
nand U6010 (N_6010,N_1282,N_2125);
nand U6011 (N_6011,N_258,N_1703);
nor U6012 (N_6012,N_417,N_3215);
and U6013 (N_6013,N_3430,N_3796);
or U6014 (N_6014,N_441,N_1374);
nand U6015 (N_6015,N_1363,N_1111);
xnor U6016 (N_6016,N_1572,N_1529);
and U6017 (N_6017,N_190,N_477);
and U6018 (N_6018,N_1156,N_3009);
and U6019 (N_6019,N_439,N_2598);
nor U6020 (N_6020,N_28,N_1074);
or U6021 (N_6021,N_1959,N_862);
nand U6022 (N_6022,N_3808,N_3814);
xnor U6023 (N_6023,N_2618,N_1969);
and U6024 (N_6024,N_1615,N_2090);
and U6025 (N_6025,N_2374,N_1501);
xor U6026 (N_6026,N_3118,N_2498);
or U6027 (N_6027,N_2450,N_3954);
nand U6028 (N_6028,N_361,N_2488);
or U6029 (N_6029,N_2630,N_1413);
or U6030 (N_6030,N_1945,N_2661);
nor U6031 (N_6031,N_3272,N_693);
xnor U6032 (N_6032,N_916,N_849);
nand U6033 (N_6033,N_259,N_3937);
nand U6034 (N_6034,N_2351,N_3850);
and U6035 (N_6035,N_2131,N_3416);
nor U6036 (N_6036,N_2711,N_3770);
or U6037 (N_6037,N_93,N_2340);
or U6038 (N_6038,N_1300,N_1199);
and U6039 (N_6039,N_3111,N_2172);
nor U6040 (N_6040,N_487,N_1576);
and U6041 (N_6041,N_2923,N_665);
and U6042 (N_6042,N_2291,N_333);
nand U6043 (N_6043,N_1503,N_1242);
and U6044 (N_6044,N_274,N_609);
and U6045 (N_6045,N_3493,N_1899);
or U6046 (N_6046,N_1144,N_1513);
nor U6047 (N_6047,N_2089,N_3507);
nand U6048 (N_6048,N_2887,N_2669);
nand U6049 (N_6049,N_1839,N_3090);
nor U6050 (N_6050,N_311,N_393);
or U6051 (N_6051,N_719,N_3054);
and U6052 (N_6052,N_3881,N_3739);
nand U6053 (N_6053,N_3698,N_3666);
xor U6054 (N_6054,N_2950,N_2659);
nand U6055 (N_6055,N_2007,N_2691);
or U6056 (N_6056,N_1151,N_1849);
and U6057 (N_6057,N_1816,N_3096);
nor U6058 (N_6058,N_1962,N_2699);
xnor U6059 (N_6059,N_2707,N_1421);
nor U6060 (N_6060,N_1212,N_1373);
nand U6061 (N_6061,N_1547,N_2134);
xnor U6062 (N_6062,N_2333,N_81);
or U6063 (N_6063,N_3915,N_247);
and U6064 (N_6064,N_714,N_3942);
or U6065 (N_6065,N_1162,N_3737);
xor U6066 (N_6066,N_209,N_2012);
xor U6067 (N_6067,N_3498,N_2389);
or U6068 (N_6068,N_3214,N_1221);
nand U6069 (N_6069,N_995,N_898);
and U6070 (N_6070,N_884,N_439);
nor U6071 (N_6071,N_2491,N_1977);
and U6072 (N_6072,N_340,N_1390);
or U6073 (N_6073,N_764,N_3471);
nand U6074 (N_6074,N_3647,N_2502);
and U6075 (N_6075,N_1969,N_124);
and U6076 (N_6076,N_745,N_3240);
nand U6077 (N_6077,N_776,N_3670);
xnor U6078 (N_6078,N_2108,N_2396);
nand U6079 (N_6079,N_2349,N_1615);
or U6080 (N_6080,N_3442,N_935);
and U6081 (N_6081,N_2752,N_592);
xor U6082 (N_6082,N_1350,N_718);
xor U6083 (N_6083,N_2623,N_3101);
nand U6084 (N_6084,N_3551,N_2672);
and U6085 (N_6085,N_3587,N_1992);
nor U6086 (N_6086,N_2353,N_1006);
nor U6087 (N_6087,N_3470,N_3211);
xor U6088 (N_6088,N_3971,N_1294);
or U6089 (N_6089,N_437,N_3957);
or U6090 (N_6090,N_2826,N_3852);
or U6091 (N_6091,N_1965,N_1293);
xor U6092 (N_6092,N_613,N_2933);
and U6093 (N_6093,N_372,N_2837);
or U6094 (N_6094,N_830,N_3024);
nor U6095 (N_6095,N_275,N_2111);
xnor U6096 (N_6096,N_3445,N_2792);
and U6097 (N_6097,N_888,N_3675);
nor U6098 (N_6098,N_3883,N_1859);
and U6099 (N_6099,N_2328,N_160);
and U6100 (N_6100,N_860,N_2083);
or U6101 (N_6101,N_2238,N_3300);
xnor U6102 (N_6102,N_2815,N_3806);
or U6103 (N_6103,N_106,N_2613);
and U6104 (N_6104,N_2654,N_3509);
or U6105 (N_6105,N_3557,N_1609);
nand U6106 (N_6106,N_1713,N_814);
xor U6107 (N_6107,N_3903,N_2792);
xor U6108 (N_6108,N_2990,N_502);
nor U6109 (N_6109,N_2884,N_445);
nand U6110 (N_6110,N_376,N_2018);
xnor U6111 (N_6111,N_500,N_3519);
or U6112 (N_6112,N_529,N_2393);
and U6113 (N_6113,N_280,N_2073);
nand U6114 (N_6114,N_357,N_1258);
and U6115 (N_6115,N_2995,N_802);
nand U6116 (N_6116,N_2513,N_1148);
or U6117 (N_6117,N_3728,N_1589);
xnor U6118 (N_6118,N_3625,N_2991);
nor U6119 (N_6119,N_2878,N_1449);
or U6120 (N_6120,N_2627,N_1577);
or U6121 (N_6121,N_1374,N_1516);
nand U6122 (N_6122,N_1626,N_2079);
and U6123 (N_6123,N_2258,N_877);
xnor U6124 (N_6124,N_1114,N_2174);
xor U6125 (N_6125,N_3161,N_1342);
nor U6126 (N_6126,N_3565,N_1855);
xnor U6127 (N_6127,N_1015,N_1768);
or U6128 (N_6128,N_360,N_2530);
or U6129 (N_6129,N_2062,N_2823);
and U6130 (N_6130,N_1607,N_3070);
or U6131 (N_6131,N_1804,N_2090);
or U6132 (N_6132,N_3902,N_2271);
and U6133 (N_6133,N_1292,N_2714);
xor U6134 (N_6134,N_1399,N_842);
nor U6135 (N_6135,N_574,N_494);
or U6136 (N_6136,N_202,N_2989);
and U6137 (N_6137,N_3022,N_272);
or U6138 (N_6138,N_115,N_2944);
nor U6139 (N_6139,N_3569,N_1711);
xor U6140 (N_6140,N_3415,N_1282);
or U6141 (N_6141,N_1829,N_2379);
nand U6142 (N_6142,N_3143,N_3953);
and U6143 (N_6143,N_1794,N_1703);
xnor U6144 (N_6144,N_2805,N_2747);
nor U6145 (N_6145,N_2757,N_3724);
and U6146 (N_6146,N_78,N_2786);
or U6147 (N_6147,N_2498,N_2563);
and U6148 (N_6148,N_3448,N_2409);
xor U6149 (N_6149,N_2805,N_3045);
and U6150 (N_6150,N_844,N_766);
or U6151 (N_6151,N_299,N_2247);
xor U6152 (N_6152,N_8,N_2497);
and U6153 (N_6153,N_3898,N_1298);
or U6154 (N_6154,N_335,N_3617);
and U6155 (N_6155,N_1937,N_3786);
xnor U6156 (N_6156,N_3405,N_3095);
or U6157 (N_6157,N_2693,N_1072);
nor U6158 (N_6158,N_1420,N_2960);
and U6159 (N_6159,N_2760,N_1036);
nor U6160 (N_6160,N_2731,N_1431);
nand U6161 (N_6161,N_1363,N_2524);
nand U6162 (N_6162,N_1479,N_484);
nor U6163 (N_6163,N_2580,N_1376);
nor U6164 (N_6164,N_436,N_3474);
and U6165 (N_6165,N_2200,N_1813);
nor U6166 (N_6166,N_2925,N_2046);
and U6167 (N_6167,N_667,N_2808);
or U6168 (N_6168,N_764,N_3440);
nand U6169 (N_6169,N_3418,N_946);
xor U6170 (N_6170,N_1423,N_2211);
nor U6171 (N_6171,N_183,N_583);
or U6172 (N_6172,N_3388,N_778);
nand U6173 (N_6173,N_733,N_3532);
xnor U6174 (N_6174,N_1023,N_3507);
nand U6175 (N_6175,N_385,N_1967);
xor U6176 (N_6176,N_3610,N_1817);
and U6177 (N_6177,N_2009,N_1886);
nor U6178 (N_6178,N_2116,N_611);
nor U6179 (N_6179,N_2450,N_410);
and U6180 (N_6180,N_2341,N_583);
xnor U6181 (N_6181,N_3274,N_3236);
and U6182 (N_6182,N_569,N_2612);
xor U6183 (N_6183,N_2109,N_1924);
nand U6184 (N_6184,N_2286,N_808);
xor U6185 (N_6185,N_119,N_2427);
xnor U6186 (N_6186,N_1337,N_1612);
xnor U6187 (N_6187,N_1771,N_2738);
xor U6188 (N_6188,N_825,N_3010);
nand U6189 (N_6189,N_3552,N_3917);
xnor U6190 (N_6190,N_210,N_2666);
xor U6191 (N_6191,N_95,N_1571);
xor U6192 (N_6192,N_2776,N_2673);
nand U6193 (N_6193,N_2257,N_998);
nor U6194 (N_6194,N_2562,N_2743);
and U6195 (N_6195,N_3423,N_2670);
nand U6196 (N_6196,N_2836,N_1749);
or U6197 (N_6197,N_542,N_2997);
and U6198 (N_6198,N_1659,N_2628);
xor U6199 (N_6199,N_1012,N_3030);
and U6200 (N_6200,N_2803,N_3414);
nand U6201 (N_6201,N_1625,N_2577);
nor U6202 (N_6202,N_2020,N_235);
nand U6203 (N_6203,N_997,N_1008);
nor U6204 (N_6204,N_1900,N_3472);
nand U6205 (N_6205,N_117,N_1216);
and U6206 (N_6206,N_401,N_3673);
nand U6207 (N_6207,N_3492,N_3594);
nor U6208 (N_6208,N_3320,N_1916);
nor U6209 (N_6209,N_795,N_82);
nand U6210 (N_6210,N_3469,N_3356);
and U6211 (N_6211,N_592,N_671);
nor U6212 (N_6212,N_795,N_222);
xor U6213 (N_6213,N_901,N_2984);
or U6214 (N_6214,N_2650,N_1757);
nor U6215 (N_6215,N_3978,N_2747);
or U6216 (N_6216,N_1801,N_1439);
xor U6217 (N_6217,N_1130,N_1479);
nand U6218 (N_6218,N_2438,N_3371);
and U6219 (N_6219,N_468,N_1166);
xnor U6220 (N_6220,N_1467,N_82);
xnor U6221 (N_6221,N_3201,N_2450);
nand U6222 (N_6222,N_3924,N_832);
or U6223 (N_6223,N_1704,N_3750);
and U6224 (N_6224,N_2440,N_1982);
nand U6225 (N_6225,N_2107,N_11);
nor U6226 (N_6226,N_1045,N_1599);
xor U6227 (N_6227,N_2326,N_3855);
nand U6228 (N_6228,N_396,N_1207);
or U6229 (N_6229,N_1402,N_1233);
nand U6230 (N_6230,N_2582,N_3874);
xor U6231 (N_6231,N_2414,N_1727);
and U6232 (N_6232,N_1929,N_3939);
xnor U6233 (N_6233,N_613,N_1571);
nand U6234 (N_6234,N_1622,N_370);
or U6235 (N_6235,N_3312,N_1959);
nand U6236 (N_6236,N_1588,N_125);
nand U6237 (N_6237,N_1206,N_1482);
nor U6238 (N_6238,N_2857,N_983);
xor U6239 (N_6239,N_1354,N_3815);
and U6240 (N_6240,N_2714,N_3008);
and U6241 (N_6241,N_3199,N_1930);
nor U6242 (N_6242,N_570,N_3539);
or U6243 (N_6243,N_3278,N_1795);
xor U6244 (N_6244,N_2805,N_1628);
nand U6245 (N_6245,N_3283,N_2610);
nand U6246 (N_6246,N_2691,N_3131);
nand U6247 (N_6247,N_2536,N_872);
or U6248 (N_6248,N_3986,N_2851);
or U6249 (N_6249,N_3436,N_382);
nor U6250 (N_6250,N_2223,N_2494);
xnor U6251 (N_6251,N_2613,N_2031);
nor U6252 (N_6252,N_3411,N_3997);
xor U6253 (N_6253,N_3532,N_3100);
xnor U6254 (N_6254,N_1180,N_2980);
nor U6255 (N_6255,N_3172,N_856);
or U6256 (N_6256,N_3989,N_848);
and U6257 (N_6257,N_475,N_1196);
and U6258 (N_6258,N_86,N_2015);
nor U6259 (N_6259,N_2151,N_1209);
nand U6260 (N_6260,N_899,N_361);
and U6261 (N_6261,N_1562,N_1966);
nand U6262 (N_6262,N_3925,N_3025);
xor U6263 (N_6263,N_3678,N_2158);
xnor U6264 (N_6264,N_2867,N_2616);
and U6265 (N_6265,N_2681,N_75);
xor U6266 (N_6266,N_1321,N_580);
nand U6267 (N_6267,N_1529,N_1894);
nor U6268 (N_6268,N_546,N_1786);
or U6269 (N_6269,N_2367,N_288);
or U6270 (N_6270,N_3529,N_3727);
and U6271 (N_6271,N_2795,N_1768);
xnor U6272 (N_6272,N_2475,N_1081);
nand U6273 (N_6273,N_908,N_3047);
or U6274 (N_6274,N_3341,N_1785);
xor U6275 (N_6275,N_2748,N_3621);
nand U6276 (N_6276,N_1329,N_2798);
nand U6277 (N_6277,N_343,N_3133);
or U6278 (N_6278,N_545,N_3531);
xor U6279 (N_6279,N_2621,N_821);
and U6280 (N_6280,N_262,N_3376);
or U6281 (N_6281,N_1117,N_437);
nor U6282 (N_6282,N_794,N_2600);
or U6283 (N_6283,N_1383,N_2390);
or U6284 (N_6284,N_3492,N_1221);
or U6285 (N_6285,N_915,N_2939);
xnor U6286 (N_6286,N_2368,N_3122);
nor U6287 (N_6287,N_3342,N_2591);
nor U6288 (N_6288,N_2988,N_2774);
or U6289 (N_6289,N_1551,N_631);
nor U6290 (N_6290,N_1196,N_2839);
nor U6291 (N_6291,N_1529,N_1843);
nand U6292 (N_6292,N_1594,N_1992);
and U6293 (N_6293,N_2272,N_1207);
or U6294 (N_6294,N_652,N_1876);
nor U6295 (N_6295,N_727,N_1478);
or U6296 (N_6296,N_3097,N_1711);
nor U6297 (N_6297,N_186,N_331);
nand U6298 (N_6298,N_888,N_1421);
xnor U6299 (N_6299,N_3055,N_2504);
or U6300 (N_6300,N_1174,N_2150);
or U6301 (N_6301,N_790,N_2444);
and U6302 (N_6302,N_2508,N_3946);
nand U6303 (N_6303,N_1987,N_1337);
or U6304 (N_6304,N_2321,N_3270);
or U6305 (N_6305,N_904,N_481);
nor U6306 (N_6306,N_3440,N_524);
or U6307 (N_6307,N_1143,N_563);
and U6308 (N_6308,N_3060,N_2353);
nand U6309 (N_6309,N_3097,N_3520);
nor U6310 (N_6310,N_3793,N_164);
or U6311 (N_6311,N_3952,N_3955);
or U6312 (N_6312,N_3597,N_455);
nor U6313 (N_6313,N_1510,N_497);
or U6314 (N_6314,N_3276,N_16);
xnor U6315 (N_6315,N_2763,N_263);
nor U6316 (N_6316,N_2337,N_1980);
or U6317 (N_6317,N_1157,N_3995);
xnor U6318 (N_6318,N_46,N_1196);
xor U6319 (N_6319,N_1431,N_363);
nor U6320 (N_6320,N_2868,N_2020);
nand U6321 (N_6321,N_2401,N_2743);
and U6322 (N_6322,N_21,N_1649);
xnor U6323 (N_6323,N_1188,N_3593);
nand U6324 (N_6324,N_1972,N_2545);
nand U6325 (N_6325,N_1587,N_630);
or U6326 (N_6326,N_3964,N_1390);
nor U6327 (N_6327,N_2242,N_967);
xor U6328 (N_6328,N_1114,N_704);
and U6329 (N_6329,N_1389,N_400);
or U6330 (N_6330,N_2061,N_3740);
or U6331 (N_6331,N_3874,N_1696);
xor U6332 (N_6332,N_3972,N_2233);
and U6333 (N_6333,N_2041,N_314);
and U6334 (N_6334,N_512,N_3157);
nand U6335 (N_6335,N_3238,N_2793);
xnor U6336 (N_6336,N_1917,N_789);
and U6337 (N_6337,N_2374,N_2878);
or U6338 (N_6338,N_3241,N_1156);
and U6339 (N_6339,N_2007,N_510);
nor U6340 (N_6340,N_1860,N_1484);
nor U6341 (N_6341,N_3008,N_3422);
nand U6342 (N_6342,N_1520,N_276);
nand U6343 (N_6343,N_3505,N_1040);
nor U6344 (N_6344,N_145,N_534);
and U6345 (N_6345,N_2974,N_3660);
or U6346 (N_6346,N_2094,N_3721);
or U6347 (N_6347,N_658,N_101);
xnor U6348 (N_6348,N_3223,N_3884);
nor U6349 (N_6349,N_847,N_1576);
nand U6350 (N_6350,N_3393,N_2698);
nor U6351 (N_6351,N_1941,N_537);
nand U6352 (N_6352,N_2795,N_2492);
nor U6353 (N_6353,N_2318,N_2035);
or U6354 (N_6354,N_560,N_1666);
nand U6355 (N_6355,N_1139,N_1721);
nand U6356 (N_6356,N_2123,N_1534);
xnor U6357 (N_6357,N_121,N_2140);
or U6358 (N_6358,N_1647,N_2460);
nand U6359 (N_6359,N_3253,N_953);
or U6360 (N_6360,N_1005,N_395);
and U6361 (N_6361,N_716,N_133);
nand U6362 (N_6362,N_168,N_448);
and U6363 (N_6363,N_1899,N_3741);
or U6364 (N_6364,N_3923,N_531);
xnor U6365 (N_6365,N_312,N_3230);
xnor U6366 (N_6366,N_1457,N_2566);
nor U6367 (N_6367,N_2012,N_1394);
xor U6368 (N_6368,N_395,N_582);
and U6369 (N_6369,N_2917,N_1580);
nor U6370 (N_6370,N_502,N_95);
nand U6371 (N_6371,N_1814,N_3478);
xor U6372 (N_6372,N_297,N_3823);
nand U6373 (N_6373,N_3876,N_2948);
and U6374 (N_6374,N_863,N_542);
nor U6375 (N_6375,N_32,N_3068);
xnor U6376 (N_6376,N_319,N_2391);
and U6377 (N_6377,N_3589,N_1729);
xnor U6378 (N_6378,N_50,N_1033);
nor U6379 (N_6379,N_2959,N_2161);
or U6380 (N_6380,N_1901,N_3709);
or U6381 (N_6381,N_650,N_3769);
nor U6382 (N_6382,N_2862,N_3717);
xor U6383 (N_6383,N_2628,N_636);
or U6384 (N_6384,N_651,N_1114);
nand U6385 (N_6385,N_2759,N_342);
nand U6386 (N_6386,N_3853,N_3175);
or U6387 (N_6387,N_1452,N_1165);
xnor U6388 (N_6388,N_1736,N_2923);
xnor U6389 (N_6389,N_83,N_943);
nor U6390 (N_6390,N_3559,N_3629);
nor U6391 (N_6391,N_161,N_1204);
nor U6392 (N_6392,N_2091,N_670);
xor U6393 (N_6393,N_580,N_1308);
and U6394 (N_6394,N_2240,N_292);
and U6395 (N_6395,N_1072,N_2744);
and U6396 (N_6396,N_2104,N_1940);
or U6397 (N_6397,N_1920,N_3356);
nor U6398 (N_6398,N_2278,N_1760);
nor U6399 (N_6399,N_2795,N_245);
or U6400 (N_6400,N_839,N_3075);
and U6401 (N_6401,N_1535,N_3189);
nand U6402 (N_6402,N_1759,N_3475);
nor U6403 (N_6403,N_2493,N_263);
nor U6404 (N_6404,N_1607,N_2876);
nor U6405 (N_6405,N_1967,N_2198);
xnor U6406 (N_6406,N_2810,N_2670);
and U6407 (N_6407,N_3951,N_1831);
and U6408 (N_6408,N_2135,N_1113);
nor U6409 (N_6409,N_1858,N_2877);
or U6410 (N_6410,N_867,N_3169);
nor U6411 (N_6411,N_2105,N_1684);
and U6412 (N_6412,N_1128,N_1928);
and U6413 (N_6413,N_2489,N_2712);
nand U6414 (N_6414,N_3866,N_3518);
nand U6415 (N_6415,N_169,N_3891);
and U6416 (N_6416,N_1213,N_684);
xor U6417 (N_6417,N_989,N_1931);
nand U6418 (N_6418,N_1782,N_2021);
nand U6419 (N_6419,N_3656,N_1835);
or U6420 (N_6420,N_3152,N_3284);
xnor U6421 (N_6421,N_12,N_2866);
and U6422 (N_6422,N_452,N_814);
xor U6423 (N_6423,N_1695,N_3412);
and U6424 (N_6424,N_2424,N_1441);
xnor U6425 (N_6425,N_2894,N_3136);
nand U6426 (N_6426,N_1321,N_845);
and U6427 (N_6427,N_3796,N_3714);
and U6428 (N_6428,N_3655,N_2454);
and U6429 (N_6429,N_2440,N_2390);
nor U6430 (N_6430,N_444,N_2160);
xnor U6431 (N_6431,N_497,N_344);
nor U6432 (N_6432,N_1647,N_2683);
nand U6433 (N_6433,N_1314,N_895);
and U6434 (N_6434,N_271,N_2015);
xor U6435 (N_6435,N_952,N_545);
nor U6436 (N_6436,N_2369,N_1355);
nor U6437 (N_6437,N_3984,N_3862);
and U6438 (N_6438,N_2321,N_1817);
or U6439 (N_6439,N_3150,N_2173);
or U6440 (N_6440,N_461,N_3415);
nand U6441 (N_6441,N_2832,N_549);
nor U6442 (N_6442,N_2354,N_1422);
xnor U6443 (N_6443,N_3320,N_540);
or U6444 (N_6444,N_801,N_2387);
and U6445 (N_6445,N_127,N_2923);
nor U6446 (N_6446,N_2586,N_3151);
or U6447 (N_6447,N_858,N_2003);
nand U6448 (N_6448,N_3748,N_3802);
nand U6449 (N_6449,N_3903,N_2433);
and U6450 (N_6450,N_1951,N_987);
and U6451 (N_6451,N_3289,N_551);
or U6452 (N_6452,N_3759,N_1766);
nor U6453 (N_6453,N_1039,N_2582);
nand U6454 (N_6454,N_2243,N_2112);
xor U6455 (N_6455,N_1963,N_1861);
nand U6456 (N_6456,N_2155,N_720);
nand U6457 (N_6457,N_1603,N_1944);
and U6458 (N_6458,N_1712,N_859);
and U6459 (N_6459,N_1489,N_1819);
and U6460 (N_6460,N_2250,N_3466);
and U6461 (N_6461,N_3741,N_316);
or U6462 (N_6462,N_2445,N_2237);
nor U6463 (N_6463,N_1082,N_1557);
or U6464 (N_6464,N_2989,N_747);
xor U6465 (N_6465,N_3894,N_407);
nand U6466 (N_6466,N_3193,N_3682);
or U6467 (N_6467,N_2814,N_1045);
xor U6468 (N_6468,N_3883,N_1154);
nor U6469 (N_6469,N_1434,N_165);
xor U6470 (N_6470,N_286,N_3730);
nand U6471 (N_6471,N_641,N_2378);
nor U6472 (N_6472,N_3247,N_3755);
nand U6473 (N_6473,N_1356,N_3120);
or U6474 (N_6474,N_412,N_771);
and U6475 (N_6475,N_9,N_2881);
or U6476 (N_6476,N_1648,N_230);
and U6477 (N_6477,N_944,N_1926);
and U6478 (N_6478,N_909,N_2607);
nor U6479 (N_6479,N_2342,N_3614);
and U6480 (N_6480,N_732,N_408);
or U6481 (N_6481,N_3370,N_3340);
and U6482 (N_6482,N_1497,N_3689);
xnor U6483 (N_6483,N_883,N_485);
nor U6484 (N_6484,N_2950,N_1233);
nor U6485 (N_6485,N_2711,N_2086);
or U6486 (N_6486,N_1099,N_3383);
or U6487 (N_6487,N_2810,N_1096);
or U6488 (N_6488,N_1530,N_2295);
xnor U6489 (N_6489,N_3556,N_2540);
or U6490 (N_6490,N_3703,N_344);
and U6491 (N_6491,N_1553,N_2430);
nand U6492 (N_6492,N_2489,N_1575);
nand U6493 (N_6493,N_867,N_2666);
and U6494 (N_6494,N_1217,N_3323);
nand U6495 (N_6495,N_2637,N_2982);
nor U6496 (N_6496,N_2854,N_1452);
nor U6497 (N_6497,N_1231,N_824);
or U6498 (N_6498,N_1192,N_3713);
nand U6499 (N_6499,N_3473,N_3579);
or U6500 (N_6500,N_649,N_1378);
nand U6501 (N_6501,N_2307,N_2079);
nor U6502 (N_6502,N_765,N_845);
nand U6503 (N_6503,N_2851,N_3444);
nand U6504 (N_6504,N_3984,N_2676);
xor U6505 (N_6505,N_1453,N_147);
or U6506 (N_6506,N_1380,N_3896);
and U6507 (N_6507,N_913,N_2909);
nand U6508 (N_6508,N_974,N_3836);
or U6509 (N_6509,N_1160,N_2825);
and U6510 (N_6510,N_2532,N_2457);
and U6511 (N_6511,N_3083,N_1119);
or U6512 (N_6512,N_1817,N_3723);
or U6513 (N_6513,N_3312,N_3734);
nand U6514 (N_6514,N_3651,N_1451);
nor U6515 (N_6515,N_3375,N_2262);
and U6516 (N_6516,N_3110,N_3605);
or U6517 (N_6517,N_943,N_2326);
and U6518 (N_6518,N_2494,N_2156);
and U6519 (N_6519,N_3257,N_651);
or U6520 (N_6520,N_1661,N_2935);
nand U6521 (N_6521,N_3439,N_3388);
or U6522 (N_6522,N_2372,N_1289);
nand U6523 (N_6523,N_170,N_3575);
xor U6524 (N_6524,N_2632,N_247);
xnor U6525 (N_6525,N_3952,N_3860);
xnor U6526 (N_6526,N_3315,N_1274);
xnor U6527 (N_6527,N_1678,N_374);
nor U6528 (N_6528,N_1320,N_3547);
and U6529 (N_6529,N_1283,N_864);
nand U6530 (N_6530,N_556,N_3136);
nor U6531 (N_6531,N_2316,N_3487);
or U6532 (N_6532,N_3066,N_361);
and U6533 (N_6533,N_3290,N_3707);
and U6534 (N_6534,N_2660,N_599);
and U6535 (N_6535,N_3874,N_684);
or U6536 (N_6536,N_660,N_677);
and U6537 (N_6537,N_3486,N_1779);
or U6538 (N_6538,N_760,N_328);
and U6539 (N_6539,N_3011,N_3266);
xor U6540 (N_6540,N_2482,N_1965);
nor U6541 (N_6541,N_699,N_1658);
or U6542 (N_6542,N_2292,N_1566);
or U6543 (N_6543,N_1114,N_181);
or U6544 (N_6544,N_2167,N_1251);
xnor U6545 (N_6545,N_2418,N_2795);
or U6546 (N_6546,N_2818,N_1885);
xor U6547 (N_6547,N_2807,N_3467);
or U6548 (N_6548,N_1401,N_3233);
xnor U6549 (N_6549,N_3244,N_1473);
and U6550 (N_6550,N_2813,N_3030);
and U6551 (N_6551,N_1679,N_3004);
nor U6552 (N_6552,N_401,N_2353);
or U6553 (N_6553,N_3540,N_669);
or U6554 (N_6554,N_3872,N_2373);
and U6555 (N_6555,N_2339,N_1959);
xnor U6556 (N_6556,N_2436,N_2205);
xnor U6557 (N_6557,N_1196,N_2602);
nand U6558 (N_6558,N_2611,N_444);
nor U6559 (N_6559,N_2385,N_91);
nand U6560 (N_6560,N_3216,N_1176);
or U6561 (N_6561,N_1016,N_1671);
xnor U6562 (N_6562,N_650,N_294);
xor U6563 (N_6563,N_3568,N_1360);
nand U6564 (N_6564,N_3001,N_2241);
or U6565 (N_6565,N_687,N_1192);
or U6566 (N_6566,N_3932,N_867);
and U6567 (N_6567,N_1308,N_1706);
nor U6568 (N_6568,N_1348,N_567);
xor U6569 (N_6569,N_55,N_3999);
xnor U6570 (N_6570,N_698,N_1993);
xnor U6571 (N_6571,N_862,N_333);
nor U6572 (N_6572,N_1230,N_949);
xnor U6573 (N_6573,N_3464,N_2393);
and U6574 (N_6574,N_853,N_2264);
and U6575 (N_6575,N_3530,N_90);
or U6576 (N_6576,N_2521,N_544);
or U6577 (N_6577,N_2168,N_2054);
xor U6578 (N_6578,N_1099,N_1335);
or U6579 (N_6579,N_2503,N_1706);
nand U6580 (N_6580,N_2161,N_1459);
xor U6581 (N_6581,N_2425,N_336);
and U6582 (N_6582,N_3879,N_2435);
or U6583 (N_6583,N_2975,N_1493);
xor U6584 (N_6584,N_3841,N_3501);
nor U6585 (N_6585,N_765,N_3985);
nand U6586 (N_6586,N_247,N_3796);
and U6587 (N_6587,N_2808,N_2931);
or U6588 (N_6588,N_3341,N_3964);
xnor U6589 (N_6589,N_3606,N_1372);
and U6590 (N_6590,N_3387,N_324);
nand U6591 (N_6591,N_332,N_359);
xnor U6592 (N_6592,N_2148,N_2962);
or U6593 (N_6593,N_3476,N_286);
nand U6594 (N_6594,N_1640,N_576);
nand U6595 (N_6595,N_3542,N_3978);
nor U6596 (N_6596,N_2140,N_1741);
and U6597 (N_6597,N_3189,N_2564);
xor U6598 (N_6598,N_955,N_1746);
xor U6599 (N_6599,N_96,N_1439);
nor U6600 (N_6600,N_1436,N_2346);
xor U6601 (N_6601,N_2791,N_3000);
or U6602 (N_6602,N_3693,N_469);
xor U6603 (N_6603,N_3832,N_964);
nand U6604 (N_6604,N_1899,N_2210);
nand U6605 (N_6605,N_2687,N_537);
nand U6606 (N_6606,N_1146,N_1761);
and U6607 (N_6607,N_2213,N_2946);
xnor U6608 (N_6608,N_1988,N_3482);
nor U6609 (N_6609,N_294,N_2113);
nor U6610 (N_6610,N_1169,N_952);
or U6611 (N_6611,N_3203,N_2415);
and U6612 (N_6612,N_2578,N_1722);
or U6613 (N_6613,N_802,N_2175);
or U6614 (N_6614,N_568,N_1039);
nor U6615 (N_6615,N_1123,N_875);
xor U6616 (N_6616,N_1034,N_571);
xnor U6617 (N_6617,N_3429,N_3828);
and U6618 (N_6618,N_2542,N_2521);
or U6619 (N_6619,N_2982,N_1688);
xor U6620 (N_6620,N_3665,N_172);
nand U6621 (N_6621,N_2967,N_2819);
and U6622 (N_6622,N_2400,N_1818);
or U6623 (N_6623,N_3103,N_2806);
nand U6624 (N_6624,N_2916,N_134);
nand U6625 (N_6625,N_1103,N_2143);
nand U6626 (N_6626,N_3172,N_3779);
or U6627 (N_6627,N_2383,N_3832);
xor U6628 (N_6628,N_3532,N_2646);
nand U6629 (N_6629,N_2682,N_1531);
nor U6630 (N_6630,N_2357,N_912);
and U6631 (N_6631,N_1344,N_3704);
nand U6632 (N_6632,N_3729,N_984);
xnor U6633 (N_6633,N_1709,N_73);
nand U6634 (N_6634,N_2510,N_3289);
nor U6635 (N_6635,N_995,N_3902);
and U6636 (N_6636,N_3708,N_3836);
xnor U6637 (N_6637,N_2772,N_521);
or U6638 (N_6638,N_815,N_2586);
nand U6639 (N_6639,N_3514,N_3394);
and U6640 (N_6640,N_185,N_1263);
or U6641 (N_6641,N_1142,N_346);
nand U6642 (N_6642,N_3074,N_1182);
nand U6643 (N_6643,N_2146,N_3949);
and U6644 (N_6644,N_3378,N_710);
and U6645 (N_6645,N_3254,N_3127);
and U6646 (N_6646,N_1001,N_529);
or U6647 (N_6647,N_2630,N_2564);
nor U6648 (N_6648,N_3184,N_3835);
nor U6649 (N_6649,N_1740,N_1274);
xnor U6650 (N_6650,N_3626,N_1616);
and U6651 (N_6651,N_1361,N_3819);
nor U6652 (N_6652,N_1658,N_841);
nand U6653 (N_6653,N_699,N_1860);
and U6654 (N_6654,N_715,N_139);
or U6655 (N_6655,N_3095,N_3868);
and U6656 (N_6656,N_3305,N_1513);
xnor U6657 (N_6657,N_3042,N_3691);
and U6658 (N_6658,N_2447,N_586);
and U6659 (N_6659,N_2768,N_3099);
nand U6660 (N_6660,N_3345,N_2463);
or U6661 (N_6661,N_1123,N_3909);
nor U6662 (N_6662,N_1572,N_3267);
nand U6663 (N_6663,N_2382,N_2533);
nand U6664 (N_6664,N_574,N_2993);
or U6665 (N_6665,N_494,N_1958);
xnor U6666 (N_6666,N_752,N_1225);
nand U6667 (N_6667,N_1081,N_2347);
or U6668 (N_6668,N_3721,N_2469);
and U6669 (N_6669,N_1282,N_375);
nand U6670 (N_6670,N_2445,N_770);
xnor U6671 (N_6671,N_1362,N_3806);
and U6672 (N_6672,N_2626,N_1099);
xnor U6673 (N_6673,N_2312,N_5);
xor U6674 (N_6674,N_3676,N_3013);
nand U6675 (N_6675,N_3836,N_3000);
and U6676 (N_6676,N_651,N_3653);
xnor U6677 (N_6677,N_457,N_3310);
nand U6678 (N_6678,N_1277,N_3074);
or U6679 (N_6679,N_711,N_1701);
nor U6680 (N_6680,N_2476,N_1871);
and U6681 (N_6681,N_1402,N_1105);
xor U6682 (N_6682,N_1290,N_494);
nand U6683 (N_6683,N_1680,N_2167);
xnor U6684 (N_6684,N_1172,N_3831);
or U6685 (N_6685,N_2186,N_2962);
and U6686 (N_6686,N_350,N_2185);
and U6687 (N_6687,N_2347,N_990);
and U6688 (N_6688,N_298,N_1243);
and U6689 (N_6689,N_1030,N_2324);
nor U6690 (N_6690,N_3197,N_192);
nor U6691 (N_6691,N_1978,N_3332);
nand U6692 (N_6692,N_268,N_3018);
nand U6693 (N_6693,N_3488,N_218);
nand U6694 (N_6694,N_2615,N_738);
xor U6695 (N_6695,N_2631,N_879);
and U6696 (N_6696,N_729,N_3768);
nor U6697 (N_6697,N_3064,N_3661);
or U6698 (N_6698,N_1299,N_1988);
nand U6699 (N_6699,N_402,N_1562);
xor U6700 (N_6700,N_1456,N_3402);
nand U6701 (N_6701,N_2748,N_3623);
or U6702 (N_6702,N_836,N_1575);
and U6703 (N_6703,N_247,N_53);
or U6704 (N_6704,N_449,N_3072);
or U6705 (N_6705,N_2570,N_402);
and U6706 (N_6706,N_3883,N_145);
nor U6707 (N_6707,N_422,N_1936);
xnor U6708 (N_6708,N_3373,N_536);
nor U6709 (N_6709,N_667,N_1976);
and U6710 (N_6710,N_1270,N_2264);
and U6711 (N_6711,N_3518,N_2621);
and U6712 (N_6712,N_965,N_1810);
nor U6713 (N_6713,N_3892,N_828);
nor U6714 (N_6714,N_3427,N_1189);
and U6715 (N_6715,N_250,N_1499);
nor U6716 (N_6716,N_1887,N_1397);
xnor U6717 (N_6717,N_1660,N_3243);
and U6718 (N_6718,N_321,N_3417);
nand U6719 (N_6719,N_1102,N_3450);
and U6720 (N_6720,N_3418,N_2198);
and U6721 (N_6721,N_2312,N_2902);
or U6722 (N_6722,N_1788,N_645);
or U6723 (N_6723,N_3169,N_3400);
nor U6724 (N_6724,N_3528,N_2616);
or U6725 (N_6725,N_3459,N_2855);
xor U6726 (N_6726,N_232,N_1178);
nor U6727 (N_6727,N_3378,N_1562);
nor U6728 (N_6728,N_3061,N_166);
xor U6729 (N_6729,N_37,N_3820);
nor U6730 (N_6730,N_1064,N_3268);
nor U6731 (N_6731,N_3699,N_3052);
nor U6732 (N_6732,N_145,N_2877);
nor U6733 (N_6733,N_2918,N_704);
nor U6734 (N_6734,N_512,N_371);
nand U6735 (N_6735,N_1377,N_656);
and U6736 (N_6736,N_560,N_1360);
nand U6737 (N_6737,N_2756,N_2018);
nand U6738 (N_6738,N_106,N_3475);
nand U6739 (N_6739,N_1234,N_3382);
or U6740 (N_6740,N_2369,N_2217);
nor U6741 (N_6741,N_2615,N_1310);
nor U6742 (N_6742,N_2323,N_1267);
and U6743 (N_6743,N_3576,N_3427);
and U6744 (N_6744,N_3779,N_112);
xor U6745 (N_6745,N_372,N_3215);
nor U6746 (N_6746,N_2504,N_971);
nand U6747 (N_6747,N_2656,N_1844);
and U6748 (N_6748,N_534,N_3051);
nor U6749 (N_6749,N_3953,N_2545);
xnor U6750 (N_6750,N_3490,N_710);
nor U6751 (N_6751,N_1910,N_3206);
nor U6752 (N_6752,N_941,N_1236);
nand U6753 (N_6753,N_166,N_2801);
nor U6754 (N_6754,N_810,N_2368);
or U6755 (N_6755,N_736,N_1483);
and U6756 (N_6756,N_3610,N_3250);
and U6757 (N_6757,N_1890,N_2527);
nand U6758 (N_6758,N_993,N_3697);
nand U6759 (N_6759,N_1790,N_2265);
xor U6760 (N_6760,N_3159,N_1686);
nor U6761 (N_6761,N_2759,N_1823);
or U6762 (N_6762,N_1330,N_1361);
or U6763 (N_6763,N_1859,N_1528);
and U6764 (N_6764,N_1936,N_2160);
nor U6765 (N_6765,N_2791,N_1603);
nand U6766 (N_6766,N_201,N_712);
or U6767 (N_6767,N_468,N_1156);
and U6768 (N_6768,N_2743,N_1566);
xnor U6769 (N_6769,N_526,N_167);
nor U6770 (N_6770,N_377,N_2614);
nor U6771 (N_6771,N_2904,N_2752);
and U6772 (N_6772,N_380,N_1763);
nor U6773 (N_6773,N_3454,N_2545);
nand U6774 (N_6774,N_2866,N_3428);
nand U6775 (N_6775,N_3634,N_3146);
nand U6776 (N_6776,N_412,N_1534);
nor U6777 (N_6777,N_1396,N_3800);
or U6778 (N_6778,N_2855,N_1406);
or U6779 (N_6779,N_3508,N_1125);
and U6780 (N_6780,N_50,N_717);
nand U6781 (N_6781,N_730,N_1362);
and U6782 (N_6782,N_3415,N_2553);
or U6783 (N_6783,N_2695,N_821);
or U6784 (N_6784,N_1160,N_900);
nor U6785 (N_6785,N_2976,N_380);
or U6786 (N_6786,N_646,N_699);
nand U6787 (N_6787,N_1065,N_1021);
nor U6788 (N_6788,N_2171,N_734);
nor U6789 (N_6789,N_666,N_2125);
nand U6790 (N_6790,N_1282,N_1020);
nor U6791 (N_6791,N_1890,N_2257);
xor U6792 (N_6792,N_2460,N_2075);
nor U6793 (N_6793,N_2385,N_2841);
nor U6794 (N_6794,N_3761,N_2300);
and U6795 (N_6795,N_1465,N_1617);
xnor U6796 (N_6796,N_143,N_2790);
xor U6797 (N_6797,N_1076,N_1127);
and U6798 (N_6798,N_825,N_487);
or U6799 (N_6799,N_3313,N_1534);
and U6800 (N_6800,N_1067,N_1774);
or U6801 (N_6801,N_3059,N_1353);
xnor U6802 (N_6802,N_2247,N_844);
nand U6803 (N_6803,N_3927,N_1864);
or U6804 (N_6804,N_1961,N_1566);
nand U6805 (N_6805,N_957,N_3857);
nor U6806 (N_6806,N_3344,N_1014);
and U6807 (N_6807,N_1314,N_3199);
or U6808 (N_6808,N_3555,N_3434);
nand U6809 (N_6809,N_3585,N_1955);
and U6810 (N_6810,N_2811,N_2673);
or U6811 (N_6811,N_3875,N_2929);
or U6812 (N_6812,N_3887,N_3175);
and U6813 (N_6813,N_32,N_1066);
or U6814 (N_6814,N_25,N_2018);
nor U6815 (N_6815,N_3879,N_3940);
and U6816 (N_6816,N_2228,N_655);
xor U6817 (N_6817,N_3807,N_1452);
nor U6818 (N_6818,N_341,N_2845);
nor U6819 (N_6819,N_1207,N_3508);
nand U6820 (N_6820,N_3827,N_60);
and U6821 (N_6821,N_3060,N_668);
nand U6822 (N_6822,N_704,N_3103);
or U6823 (N_6823,N_3609,N_3869);
nand U6824 (N_6824,N_554,N_3185);
or U6825 (N_6825,N_1211,N_2446);
or U6826 (N_6826,N_3933,N_2049);
or U6827 (N_6827,N_1535,N_119);
xor U6828 (N_6828,N_2521,N_2492);
or U6829 (N_6829,N_2468,N_2500);
or U6830 (N_6830,N_961,N_2851);
xor U6831 (N_6831,N_2501,N_2695);
xor U6832 (N_6832,N_3240,N_3794);
and U6833 (N_6833,N_1745,N_2498);
xnor U6834 (N_6834,N_3535,N_47);
xnor U6835 (N_6835,N_177,N_1997);
xor U6836 (N_6836,N_3335,N_3271);
nor U6837 (N_6837,N_3386,N_1625);
xnor U6838 (N_6838,N_3325,N_3822);
xor U6839 (N_6839,N_2083,N_2142);
nor U6840 (N_6840,N_3293,N_891);
nand U6841 (N_6841,N_2372,N_1070);
or U6842 (N_6842,N_1310,N_1985);
or U6843 (N_6843,N_2025,N_949);
xnor U6844 (N_6844,N_2066,N_3707);
nand U6845 (N_6845,N_1277,N_1854);
xor U6846 (N_6846,N_1566,N_367);
nor U6847 (N_6847,N_589,N_2362);
xor U6848 (N_6848,N_118,N_244);
nor U6849 (N_6849,N_1388,N_3637);
xor U6850 (N_6850,N_2021,N_927);
and U6851 (N_6851,N_3404,N_2781);
or U6852 (N_6852,N_2678,N_3814);
nor U6853 (N_6853,N_2994,N_1586);
or U6854 (N_6854,N_3111,N_2324);
nor U6855 (N_6855,N_302,N_1595);
or U6856 (N_6856,N_1412,N_2203);
nand U6857 (N_6857,N_156,N_269);
and U6858 (N_6858,N_1062,N_1675);
and U6859 (N_6859,N_2018,N_1079);
nand U6860 (N_6860,N_3596,N_1622);
nand U6861 (N_6861,N_901,N_3054);
nand U6862 (N_6862,N_1190,N_982);
and U6863 (N_6863,N_1694,N_1536);
nor U6864 (N_6864,N_3850,N_626);
nor U6865 (N_6865,N_3058,N_2028);
and U6866 (N_6866,N_1860,N_3260);
nand U6867 (N_6867,N_2850,N_181);
and U6868 (N_6868,N_1104,N_415);
or U6869 (N_6869,N_746,N_444);
nand U6870 (N_6870,N_1140,N_3884);
xor U6871 (N_6871,N_77,N_3797);
xnor U6872 (N_6872,N_182,N_2819);
or U6873 (N_6873,N_973,N_918);
and U6874 (N_6874,N_983,N_1694);
xnor U6875 (N_6875,N_1976,N_57);
and U6876 (N_6876,N_2886,N_620);
and U6877 (N_6877,N_1069,N_503);
xnor U6878 (N_6878,N_2178,N_1685);
or U6879 (N_6879,N_1366,N_3637);
nor U6880 (N_6880,N_3686,N_717);
xor U6881 (N_6881,N_3130,N_449);
nor U6882 (N_6882,N_64,N_228);
and U6883 (N_6883,N_1590,N_3474);
xnor U6884 (N_6884,N_1434,N_2188);
nor U6885 (N_6885,N_1260,N_2839);
xor U6886 (N_6886,N_3406,N_693);
and U6887 (N_6887,N_1237,N_3152);
xnor U6888 (N_6888,N_3537,N_879);
and U6889 (N_6889,N_976,N_277);
and U6890 (N_6890,N_3475,N_3856);
xnor U6891 (N_6891,N_1006,N_1985);
xor U6892 (N_6892,N_2183,N_1884);
nor U6893 (N_6893,N_678,N_3763);
nor U6894 (N_6894,N_2258,N_3061);
nand U6895 (N_6895,N_3535,N_3231);
xor U6896 (N_6896,N_2524,N_2218);
and U6897 (N_6897,N_2060,N_2523);
xnor U6898 (N_6898,N_1877,N_1369);
nand U6899 (N_6899,N_2703,N_1444);
nor U6900 (N_6900,N_78,N_2867);
nor U6901 (N_6901,N_1455,N_3793);
nand U6902 (N_6902,N_2961,N_1349);
or U6903 (N_6903,N_2560,N_2183);
and U6904 (N_6904,N_3099,N_90);
and U6905 (N_6905,N_2952,N_833);
xor U6906 (N_6906,N_456,N_1355);
nand U6907 (N_6907,N_512,N_2562);
nor U6908 (N_6908,N_529,N_3319);
nand U6909 (N_6909,N_983,N_1881);
nand U6910 (N_6910,N_651,N_1702);
nand U6911 (N_6911,N_2819,N_577);
xnor U6912 (N_6912,N_1847,N_3273);
or U6913 (N_6913,N_1593,N_3805);
or U6914 (N_6914,N_3640,N_1463);
xnor U6915 (N_6915,N_1122,N_2461);
or U6916 (N_6916,N_287,N_2587);
nor U6917 (N_6917,N_931,N_2853);
nand U6918 (N_6918,N_2816,N_747);
or U6919 (N_6919,N_1355,N_697);
nand U6920 (N_6920,N_3323,N_1435);
or U6921 (N_6921,N_2091,N_2024);
and U6922 (N_6922,N_1037,N_1133);
nor U6923 (N_6923,N_3146,N_1396);
nand U6924 (N_6924,N_2186,N_1975);
nor U6925 (N_6925,N_2171,N_718);
or U6926 (N_6926,N_2842,N_2019);
nand U6927 (N_6927,N_1468,N_2869);
xor U6928 (N_6928,N_1005,N_3561);
and U6929 (N_6929,N_1640,N_1564);
xnor U6930 (N_6930,N_1961,N_1694);
or U6931 (N_6931,N_338,N_1479);
nor U6932 (N_6932,N_61,N_2584);
or U6933 (N_6933,N_2111,N_558);
nand U6934 (N_6934,N_3697,N_2422);
or U6935 (N_6935,N_551,N_951);
nor U6936 (N_6936,N_2378,N_2177);
and U6937 (N_6937,N_2135,N_1465);
xor U6938 (N_6938,N_542,N_2252);
nor U6939 (N_6939,N_1889,N_2217);
or U6940 (N_6940,N_125,N_831);
nand U6941 (N_6941,N_393,N_1856);
or U6942 (N_6942,N_2844,N_3878);
nor U6943 (N_6943,N_1135,N_3669);
nand U6944 (N_6944,N_981,N_3905);
and U6945 (N_6945,N_2642,N_159);
or U6946 (N_6946,N_1109,N_1108);
and U6947 (N_6947,N_2679,N_2148);
and U6948 (N_6948,N_1793,N_3410);
nand U6949 (N_6949,N_1461,N_3058);
nor U6950 (N_6950,N_714,N_409);
or U6951 (N_6951,N_739,N_1155);
and U6952 (N_6952,N_1815,N_9);
nor U6953 (N_6953,N_3317,N_2640);
xnor U6954 (N_6954,N_592,N_2657);
nand U6955 (N_6955,N_1862,N_2565);
or U6956 (N_6956,N_473,N_3694);
or U6957 (N_6957,N_1901,N_2404);
nor U6958 (N_6958,N_2952,N_2447);
nor U6959 (N_6959,N_1822,N_2610);
or U6960 (N_6960,N_2560,N_1247);
nand U6961 (N_6961,N_2945,N_134);
and U6962 (N_6962,N_95,N_3007);
or U6963 (N_6963,N_3791,N_2014);
nor U6964 (N_6964,N_1020,N_3293);
nand U6965 (N_6965,N_1952,N_335);
or U6966 (N_6966,N_173,N_2366);
nand U6967 (N_6967,N_1990,N_2043);
or U6968 (N_6968,N_1347,N_2978);
nor U6969 (N_6969,N_545,N_627);
nand U6970 (N_6970,N_2274,N_674);
nor U6971 (N_6971,N_2711,N_596);
or U6972 (N_6972,N_1665,N_637);
nor U6973 (N_6973,N_1736,N_1587);
nand U6974 (N_6974,N_902,N_1294);
xnor U6975 (N_6975,N_2908,N_3430);
nand U6976 (N_6976,N_843,N_3140);
nand U6977 (N_6977,N_1771,N_1362);
nand U6978 (N_6978,N_1309,N_3426);
nor U6979 (N_6979,N_649,N_2706);
nand U6980 (N_6980,N_1525,N_3398);
or U6981 (N_6981,N_3259,N_3350);
xnor U6982 (N_6982,N_383,N_2042);
xor U6983 (N_6983,N_3566,N_1753);
nor U6984 (N_6984,N_3831,N_2192);
nand U6985 (N_6985,N_993,N_915);
xor U6986 (N_6986,N_1817,N_3979);
or U6987 (N_6987,N_3285,N_41);
nand U6988 (N_6988,N_2197,N_3653);
nor U6989 (N_6989,N_3302,N_3856);
and U6990 (N_6990,N_1893,N_834);
nand U6991 (N_6991,N_344,N_2575);
nand U6992 (N_6992,N_66,N_1293);
nand U6993 (N_6993,N_1273,N_3058);
or U6994 (N_6994,N_3475,N_3585);
nand U6995 (N_6995,N_3408,N_3734);
xor U6996 (N_6996,N_1357,N_3293);
and U6997 (N_6997,N_398,N_3958);
or U6998 (N_6998,N_1019,N_302);
or U6999 (N_6999,N_3321,N_713);
nor U7000 (N_7000,N_3260,N_2320);
xnor U7001 (N_7001,N_3502,N_485);
and U7002 (N_7002,N_1723,N_2903);
and U7003 (N_7003,N_2926,N_699);
nand U7004 (N_7004,N_1749,N_1781);
and U7005 (N_7005,N_110,N_2344);
xor U7006 (N_7006,N_2065,N_3495);
nand U7007 (N_7007,N_996,N_1956);
or U7008 (N_7008,N_3396,N_2018);
nor U7009 (N_7009,N_925,N_1507);
nor U7010 (N_7010,N_1229,N_1864);
xor U7011 (N_7011,N_1952,N_2458);
and U7012 (N_7012,N_1417,N_1728);
nor U7013 (N_7013,N_832,N_1005);
or U7014 (N_7014,N_2009,N_3674);
nor U7015 (N_7015,N_1301,N_733);
and U7016 (N_7016,N_1003,N_801);
nand U7017 (N_7017,N_719,N_1753);
or U7018 (N_7018,N_2012,N_2525);
and U7019 (N_7019,N_2139,N_3822);
or U7020 (N_7020,N_2259,N_3024);
or U7021 (N_7021,N_2092,N_106);
xor U7022 (N_7022,N_2302,N_3649);
xnor U7023 (N_7023,N_706,N_2802);
xnor U7024 (N_7024,N_1196,N_1342);
nor U7025 (N_7025,N_3801,N_2965);
xor U7026 (N_7026,N_3083,N_1509);
and U7027 (N_7027,N_3035,N_1909);
or U7028 (N_7028,N_3026,N_2582);
nor U7029 (N_7029,N_228,N_2485);
nand U7030 (N_7030,N_3548,N_454);
xor U7031 (N_7031,N_2961,N_3049);
and U7032 (N_7032,N_29,N_1346);
or U7033 (N_7033,N_762,N_811);
xor U7034 (N_7034,N_1744,N_13);
and U7035 (N_7035,N_1265,N_2562);
and U7036 (N_7036,N_3586,N_3650);
xnor U7037 (N_7037,N_1980,N_928);
nor U7038 (N_7038,N_1033,N_2868);
xor U7039 (N_7039,N_3656,N_3588);
or U7040 (N_7040,N_2069,N_1082);
and U7041 (N_7041,N_2394,N_2799);
nor U7042 (N_7042,N_3604,N_419);
xor U7043 (N_7043,N_1945,N_431);
and U7044 (N_7044,N_2494,N_593);
and U7045 (N_7045,N_67,N_3574);
xnor U7046 (N_7046,N_3234,N_3520);
nor U7047 (N_7047,N_3366,N_3820);
xor U7048 (N_7048,N_2840,N_691);
nand U7049 (N_7049,N_1627,N_2446);
xnor U7050 (N_7050,N_194,N_653);
xnor U7051 (N_7051,N_120,N_2688);
nor U7052 (N_7052,N_410,N_964);
or U7053 (N_7053,N_1910,N_77);
nor U7054 (N_7054,N_1888,N_1086);
or U7055 (N_7055,N_42,N_2395);
nor U7056 (N_7056,N_825,N_3835);
xnor U7057 (N_7057,N_1283,N_1429);
or U7058 (N_7058,N_1672,N_3886);
or U7059 (N_7059,N_3394,N_1464);
or U7060 (N_7060,N_1808,N_40);
xnor U7061 (N_7061,N_171,N_1943);
or U7062 (N_7062,N_982,N_2306);
nor U7063 (N_7063,N_208,N_91);
xnor U7064 (N_7064,N_1634,N_3276);
and U7065 (N_7065,N_3169,N_3120);
and U7066 (N_7066,N_2361,N_2826);
xor U7067 (N_7067,N_2047,N_1707);
and U7068 (N_7068,N_2284,N_3655);
nand U7069 (N_7069,N_147,N_3433);
nand U7070 (N_7070,N_2979,N_1084);
xor U7071 (N_7071,N_2559,N_297);
and U7072 (N_7072,N_3905,N_37);
xnor U7073 (N_7073,N_3083,N_1922);
or U7074 (N_7074,N_3206,N_1295);
and U7075 (N_7075,N_3950,N_3088);
nand U7076 (N_7076,N_3315,N_1527);
and U7077 (N_7077,N_1924,N_3837);
xnor U7078 (N_7078,N_3579,N_2401);
nand U7079 (N_7079,N_2983,N_2392);
or U7080 (N_7080,N_1026,N_2940);
nor U7081 (N_7081,N_3826,N_1200);
xnor U7082 (N_7082,N_786,N_1387);
and U7083 (N_7083,N_1311,N_1254);
nand U7084 (N_7084,N_1127,N_2207);
nor U7085 (N_7085,N_365,N_3282);
xnor U7086 (N_7086,N_3156,N_907);
nor U7087 (N_7087,N_2064,N_559);
xnor U7088 (N_7088,N_1976,N_1457);
nand U7089 (N_7089,N_751,N_3715);
nand U7090 (N_7090,N_1405,N_482);
or U7091 (N_7091,N_2331,N_1520);
xor U7092 (N_7092,N_3558,N_136);
nand U7093 (N_7093,N_3502,N_211);
or U7094 (N_7094,N_212,N_3782);
nand U7095 (N_7095,N_3621,N_1191);
or U7096 (N_7096,N_685,N_1368);
xor U7097 (N_7097,N_2137,N_1893);
nor U7098 (N_7098,N_1983,N_2984);
nand U7099 (N_7099,N_2671,N_1790);
and U7100 (N_7100,N_1181,N_3712);
and U7101 (N_7101,N_2032,N_585);
nand U7102 (N_7102,N_2569,N_2996);
nor U7103 (N_7103,N_1492,N_1764);
xor U7104 (N_7104,N_1932,N_3452);
xor U7105 (N_7105,N_3601,N_3045);
nand U7106 (N_7106,N_3264,N_3719);
and U7107 (N_7107,N_1789,N_1638);
and U7108 (N_7108,N_3121,N_3065);
and U7109 (N_7109,N_1980,N_823);
and U7110 (N_7110,N_619,N_1111);
or U7111 (N_7111,N_1377,N_3482);
and U7112 (N_7112,N_1071,N_1222);
and U7113 (N_7113,N_922,N_3627);
xor U7114 (N_7114,N_1847,N_1166);
nand U7115 (N_7115,N_1601,N_1950);
nor U7116 (N_7116,N_2300,N_1056);
and U7117 (N_7117,N_2547,N_2832);
nand U7118 (N_7118,N_1576,N_2054);
or U7119 (N_7119,N_990,N_1216);
and U7120 (N_7120,N_2334,N_447);
nor U7121 (N_7121,N_2831,N_2818);
nand U7122 (N_7122,N_2242,N_1965);
nor U7123 (N_7123,N_3735,N_2706);
xor U7124 (N_7124,N_3303,N_1673);
and U7125 (N_7125,N_755,N_1568);
nor U7126 (N_7126,N_3413,N_2875);
and U7127 (N_7127,N_2353,N_3613);
xnor U7128 (N_7128,N_2316,N_1881);
xor U7129 (N_7129,N_3655,N_690);
or U7130 (N_7130,N_2457,N_134);
and U7131 (N_7131,N_3471,N_2116);
or U7132 (N_7132,N_500,N_2832);
nand U7133 (N_7133,N_972,N_3247);
nand U7134 (N_7134,N_694,N_2784);
xor U7135 (N_7135,N_1079,N_1016);
and U7136 (N_7136,N_1208,N_2088);
or U7137 (N_7137,N_306,N_1189);
and U7138 (N_7138,N_1985,N_3494);
or U7139 (N_7139,N_3346,N_958);
and U7140 (N_7140,N_3003,N_2271);
and U7141 (N_7141,N_2153,N_1807);
xor U7142 (N_7142,N_3397,N_3094);
nor U7143 (N_7143,N_2926,N_2349);
and U7144 (N_7144,N_3468,N_2031);
nor U7145 (N_7145,N_1499,N_3378);
xnor U7146 (N_7146,N_2379,N_851);
or U7147 (N_7147,N_1773,N_2543);
nor U7148 (N_7148,N_3863,N_106);
xnor U7149 (N_7149,N_3512,N_2554);
xnor U7150 (N_7150,N_3962,N_872);
and U7151 (N_7151,N_3102,N_558);
nor U7152 (N_7152,N_755,N_3266);
or U7153 (N_7153,N_1265,N_107);
and U7154 (N_7154,N_3397,N_3606);
nand U7155 (N_7155,N_3823,N_3710);
nor U7156 (N_7156,N_2805,N_1629);
and U7157 (N_7157,N_2681,N_901);
nor U7158 (N_7158,N_133,N_1821);
nor U7159 (N_7159,N_1336,N_1386);
or U7160 (N_7160,N_3659,N_2280);
and U7161 (N_7161,N_2463,N_704);
and U7162 (N_7162,N_291,N_2948);
or U7163 (N_7163,N_850,N_3707);
nor U7164 (N_7164,N_1502,N_809);
nor U7165 (N_7165,N_3134,N_2986);
xnor U7166 (N_7166,N_144,N_3384);
nand U7167 (N_7167,N_844,N_1969);
xnor U7168 (N_7168,N_47,N_1315);
nor U7169 (N_7169,N_1742,N_1931);
nor U7170 (N_7170,N_1380,N_907);
and U7171 (N_7171,N_2269,N_3196);
or U7172 (N_7172,N_3318,N_1295);
nor U7173 (N_7173,N_3047,N_3068);
nand U7174 (N_7174,N_411,N_2077);
or U7175 (N_7175,N_866,N_925);
or U7176 (N_7176,N_3412,N_2543);
nand U7177 (N_7177,N_2831,N_2965);
or U7178 (N_7178,N_612,N_260);
nor U7179 (N_7179,N_1843,N_3431);
and U7180 (N_7180,N_2029,N_2620);
nor U7181 (N_7181,N_3022,N_860);
xor U7182 (N_7182,N_1424,N_3787);
xor U7183 (N_7183,N_891,N_36);
nand U7184 (N_7184,N_2439,N_1655);
xnor U7185 (N_7185,N_2478,N_2110);
and U7186 (N_7186,N_2355,N_2012);
nand U7187 (N_7187,N_57,N_1546);
nand U7188 (N_7188,N_3558,N_2101);
nor U7189 (N_7189,N_650,N_271);
xor U7190 (N_7190,N_3464,N_2349);
or U7191 (N_7191,N_1423,N_386);
and U7192 (N_7192,N_1593,N_385);
and U7193 (N_7193,N_3570,N_482);
nand U7194 (N_7194,N_2411,N_105);
xor U7195 (N_7195,N_176,N_2496);
and U7196 (N_7196,N_2872,N_1195);
and U7197 (N_7197,N_2089,N_2436);
or U7198 (N_7198,N_1015,N_3502);
or U7199 (N_7199,N_2085,N_2887);
xnor U7200 (N_7200,N_3926,N_3878);
or U7201 (N_7201,N_247,N_1863);
or U7202 (N_7202,N_2486,N_2339);
xor U7203 (N_7203,N_2494,N_254);
nand U7204 (N_7204,N_2836,N_243);
and U7205 (N_7205,N_3990,N_854);
and U7206 (N_7206,N_2399,N_3831);
xor U7207 (N_7207,N_3124,N_2146);
nor U7208 (N_7208,N_163,N_1167);
and U7209 (N_7209,N_536,N_501);
or U7210 (N_7210,N_1107,N_33);
xor U7211 (N_7211,N_1673,N_236);
or U7212 (N_7212,N_3620,N_274);
or U7213 (N_7213,N_1960,N_1796);
and U7214 (N_7214,N_890,N_3676);
xor U7215 (N_7215,N_29,N_1549);
or U7216 (N_7216,N_723,N_1312);
nand U7217 (N_7217,N_535,N_216);
nand U7218 (N_7218,N_3076,N_3931);
nor U7219 (N_7219,N_3211,N_798);
or U7220 (N_7220,N_1765,N_304);
nand U7221 (N_7221,N_84,N_3325);
or U7222 (N_7222,N_1472,N_1657);
and U7223 (N_7223,N_2533,N_3742);
or U7224 (N_7224,N_3259,N_1855);
nand U7225 (N_7225,N_1136,N_2817);
xor U7226 (N_7226,N_196,N_31);
nand U7227 (N_7227,N_1817,N_1595);
xnor U7228 (N_7228,N_850,N_2638);
xor U7229 (N_7229,N_1912,N_3349);
and U7230 (N_7230,N_3019,N_1712);
xor U7231 (N_7231,N_2003,N_1765);
xnor U7232 (N_7232,N_3800,N_3553);
or U7233 (N_7233,N_2481,N_2824);
xnor U7234 (N_7234,N_2587,N_1764);
and U7235 (N_7235,N_3565,N_2466);
xnor U7236 (N_7236,N_1719,N_756);
xnor U7237 (N_7237,N_565,N_1259);
or U7238 (N_7238,N_809,N_2891);
nand U7239 (N_7239,N_1546,N_3768);
xnor U7240 (N_7240,N_429,N_1913);
nand U7241 (N_7241,N_634,N_101);
or U7242 (N_7242,N_359,N_649);
and U7243 (N_7243,N_3145,N_1833);
and U7244 (N_7244,N_3850,N_1373);
and U7245 (N_7245,N_3029,N_122);
or U7246 (N_7246,N_3499,N_652);
nand U7247 (N_7247,N_2347,N_1505);
and U7248 (N_7248,N_3294,N_3337);
and U7249 (N_7249,N_3214,N_637);
xnor U7250 (N_7250,N_3427,N_3226);
and U7251 (N_7251,N_1012,N_3058);
or U7252 (N_7252,N_3075,N_1974);
nand U7253 (N_7253,N_139,N_2293);
xor U7254 (N_7254,N_606,N_551);
or U7255 (N_7255,N_3740,N_3425);
or U7256 (N_7256,N_65,N_934);
and U7257 (N_7257,N_666,N_1236);
nor U7258 (N_7258,N_2545,N_2591);
and U7259 (N_7259,N_643,N_3887);
xor U7260 (N_7260,N_1053,N_90);
nand U7261 (N_7261,N_1541,N_3676);
xnor U7262 (N_7262,N_344,N_3259);
nand U7263 (N_7263,N_1043,N_2894);
xnor U7264 (N_7264,N_882,N_746);
nor U7265 (N_7265,N_2383,N_1340);
nand U7266 (N_7266,N_971,N_52);
and U7267 (N_7267,N_1747,N_485);
xnor U7268 (N_7268,N_2033,N_207);
nand U7269 (N_7269,N_2510,N_3311);
or U7270 (N_7270,N_2730,N_152);
nand U7271 (N_7271,N_1389,N_2304);
nand U7272 (N_7272,N_1652,N_3538);
and U7273 (N_7273,N_3252,N_479);
and U7274 (N_7274,N_619,N_2006);
nor U7275 (N_7275,N_3549,N_2523);
and U7276 (N_7276,N_3487,N_31);
or U7277 (N_7277,N_3416,N_1810);
and U7278 (N_7278,N_2860,N_1650);
xnor U7279 (N_7279,N_3903,N_1181);
nand U7280 (N_7280,N_3349,N_3048);
nand U7281 (N_7281,N_3965,N_1587);
nand U7282 (N_7282,N_68,N_1243);
nand U7283 (N_7283,N_1059,N_1868);
xnor U7284 (N_7284,N_1859,N_1296);
or U7285 (N_7285,N_1142,N_1459);
nor U7286 (N_7286,N_1899,N_2641);
xnor U7287 (N_7287,N_1468,N_2651);
and U7288 (N_7288,N_736,N_2927);
and U7289 (N_7289,N_2451,N_1319);
nor U7290 (N_7290,N_1506,N_2942);
and U7291 (N_7291,N_854,N_588);
or U7292 (N_7292,N_366,N_2114);
or U7293 (N_7293,N_2982,N_9);
or U7294 (N_7294,N_2402,N_2123);
nor U7295 (N_7295,N_3958,N_1055);
nand U7296 (N_7296,N_2338,N_174);
nand U7297 (N_7297,N_1532,N_1878);
and U7298 (N_7298,N_2882,N_3748);
xnor U7299 (N_7299,N_3827,N_1406);
and U7300 (N_7300,N_1605,N_3453);
nand U7301 (N_7301,N_3206,N_683);
or U7302 (N_7302,N_224,N_3938);
and U7303 (N_7303,N_2200,N_8);
xor U7304 (N_7304,N_3687,N_673);
nor U7305 (N_7305,N_1894,N_135);
or U7306 (N_7306,N_1811,N_3957);
nand U7307 (N_7307,N_2011,N_3678);
and U7308 (N_7308,N_675,N_3195);
xnor U7309 (N_7309,N_2956,N_2412);
nand U7310 (N_7310,N_2531,N_1391);
xnor U7311 (N_7311,N_3671,N_1646);
and U7312 (N_7312,N_3247,N_3512);
nand U7313 (N_7313,N_1789,N_3789);
nor U7314 (N_7314,N_3833,N_785);
or U7315 (N_7315,N_1209,N_1443);
nor U7316 (N_7316,N_3119,N_803);
xor U7317 (N_7317,N_1964,N_3653);
nand U7318 (N_7318,N_1483,N_2504);
nor U7319 (N_7319,N_879,N_3385);
or U7320 (N_7320,N_170,N_3175);
or U7321 (N_7321,N_1338,N_2247);
xor U7322 (N_7322,N_2118,N_2009);
nor U7323 (N_7323,N_1926,N_3210);
or U7324 (N_7324,N_2837,N_3030);
nand U7325 (N_7325,N_710,N_2716);
nor U7326 (N_7326,N_341,N_2832);
or U7327 (N_7327,N_390,N_3719);
nand U7328 (N_7328,N_3822,N_358);
or U7329 (N_7329,N_1427,N_2720);
nor U7330 (N_7330,N_1364,N_336);
xor U7331 (N_7331,N_1633,N_1497);
nor U7332 (N_7332,N_1509,N_746);
nand U7333 (N_7333,N_1326,N_2469);
or U7334 (N_7334,N_2306,N_620);
and U7335 (N_7335,N_1841,N_3506);
nand U7336 (N_7336,N_2970,N_291);
nor U7337 (N_7337,N_2014,N_379);
or U7338 (N_7338,N_2532,N_3359);
and U7339 (N_7339,N_209,N_227);
nor U7340 (N_7340,N_1656,N_1879);
xor U7341 (N_7341,N_1879,N_690);
nand U7342 (N_7342,N_3616,N_2811);
and U7343 (N_7343,N_454,N_182);
xor U7344 (N_7344,N_224,N_3053);
xnor U7345 (N_7345,N_1691,N_3576);
nor U7346 (N_7346,N_2510,N_2749);
nand U7347 (N_7347,N_485,N_2728);
nor U7348 (N_7348,N_2413,N_176);
nor U7349 (N_7349,N_3030,N_1780);
and U7350 (N_7350,N_2182,N_2330);
or U7351 (N_7351,N_3150,N_3567);
or U7352 (N_7352,N_1748,N_2232);
nand U7353 (N_7353,N_2728,N_2993);
and U7354 (N_7354,N_3837,N_1759);
and U7355 (N_7355,N_2977,N_3777);
and U7356 (N_7356,N_2344,N_3068);
nand U7357 (N_7357,N_527,N_3382);
or U7358 (N_7358,N_912,N_3621);
or U7359 (N_7359,N_2077,N_589);
nand U7360 (N_7360,N_2835,N_2485);
and U7361 (N_7361,N_2888,N_3003);
nor U7362 (N_7362,N_3693,N_689);
xnor U7363 (N_7363,N_1832,N_2343);
nand U7364 (N_7364,N_624,N_2605);
xor U7365 (N_7365,N_667,N_3565);
or U7366 (N_7366,N_727,N_63);
and U7367 (N_7367,N_3307,N_1113);
and U7368 (N_7368,N_2021,N_1542);
and U7369 (N_7369,N_1188,N_2332);
and U7370 (N_7370,N_19,N_3847);
or U7371 (N_7371,N_306,N_1961);
nand U7372 (N_7372,N_1654,N_2907);
xor U7373 (N_7373,N_1589,N_540);
xor U7374 (N_7374,N_710,N_2254);
nand U7375 (N_7375,N_2409,N_3076);
and U7376 (N_7376,N_1329,N_2411);
or U7377 (N_7377,N_2337,N_1103);
nand U7378 (N_7378,N_3095,N_3075);
xnor U7379 (N_7379,N_2536,N_3601);
or U7380 (N_7380,N_1771,N_3886);
nand U7381 (N_7381,N_3471,N_2436);
nand U7382 (N_7382,N_3339,N_137);
and U7383 (N_7383,N_356,N_1787);
or U7384 (N_7384,N_3040,N_1306);
or U7385 (N_7385,N_3160,N_2891);
and U7386 (N_7386,N_1961,N_3680);
xnor U7387 (N_7387,N_880,N_2220);
xor U7388 (N_7388,N_635,N_2858);
or U7389 (N_7389,N_150,N_876);
nand U7390 (N_7390,N_1136,N_3932);
nor U7391 (N_7391,N_3965,N_884);
or U7392 (N_7392,N_1139,N_772);
or U7393 (N_7393,N_2677,N_1957);
nor U7394 (N_7394,N_2691,N_1456);
and U7395 (N_7395,N_2720,N_458);
or U7396 (N_7396,N_2972,N_3969);
nor U7397 (N_7397,N_484,N_3433);
xnor U7398 (N_7398,N_1534,N_398);
nand U7399 (N_7399,N_3976,N_1666);
xor U7400 (N_7400,N_1610,N_813);
and U7401 (N_7401,N_508,N_1232);
nor U7402 (N_7402,N_3677,N_879);
and U7403 (N_7403,N_2126,N_940);
and U7404 (N_7404,N_2711,N_2319);
xor U7405 (N_7405,N_291,N_2333);
nand U7406 (N_7406,N_3074,N_2760);
or U7407 (N_7407,N_1078,N_1241);
nor U7408 (N_7408,N_1033,N_1334);
and U7409 (N_7409,N_2410,N_720);
xnor U7410 (N_7410,N_141,N_3575);
or U7411 (N_7411,N_800,N_3125);
nor U7412 (N_7412,N_206,N_3819);
and U7413 (N_7413,N_1529,N_468);
and U7414 (N_7414,N_3512,N_1175);
nor U7415 (N_7415,N_2593,N_1963);
nor U7416 (N_7416,N_3949,N_1459);
xor U7417 (N_7417,N_1353,N_3579);
nor U7418 (N_7418,N_2214,N_461);
nand U7419 (N_7419,N_3140,N_429);
xnor U7420 (N_7420,N_1947,N_1619);
nor U7421 (N_7421,N_2248,N_3685);
or U7422 (N_7422,N_1533,N_2785);
nand U7423 (N_7423,N_1540,N_2193);
and U7424 (N_7424,N_362,N_3827);
or U7425 (N_7425,N_3755,N_3133);
and U7426 (N_7426,N_1847,N_654);
or U7427 (N_7427,N_3058,N_182);
nor U7428 (N_7428,N_2518,N_2173);
nor U7429 (N_7429,N_2799,N_2573);
nand U7430 (N_7430,N_32,N_1967);
and U7431 (N_7431,N_818,N_3805);
nor U7432 (N_7432,N_1921,N_2442);
nor U7433 (N_7433,N_872,N_594);
xnor U7434 (N_7434,N_1124,N_1581);
or U7435 (N_7435,N_1230,N_1374);
and U7436 (N_7436,N_3602,N_614);
or U7437 (N_7437,N_3105,N_1446);
xnor U7438 (N_7438,N_3840,N_2068);
nand U7439 (N_7439,N_2873,N_3709);
or U7440 (N_7440,N_248,N_295);
nand U7441 (N_7441,N_140,N_2013);
or U7442 (N_7442,N_2972,N_209);
nand U7443 (N_7443,N_2608,N_3854);
xnor U7444 (N_7444,N_2185,N_1329);
and U7445 (N_7445,N_421,N_2539);
and U7446 (N_7446,N_3390,N_73);
nand U7447 (N_7447,N_3164,N_991);
nor U7448 (N_7448,N_1569,N_2009);
nand U7449 (N_7449,N_1545,N_3270);
nand U7450 (N_7450,N_2302,N_3541);
xnor U7451 (N_7451,N_3507,N_1874);
xor U7452 (N_7452,N_155,N_473);
nor U7453 (N_7453,N_3211,N_3809);
and U7454 (N_7454,N_56,N_3012);
nor U7455 (N_7455,N_1778,N_2146);
nand U7456 (N_7456,N_1463,N_2185);
xnor U7457 (N_7457,N_1988,N_15);
nor U7458 (N_7458,N_2486,N_3064);
nand U7459 (N_7459,N_488,N_1329);
nand U7460 (N_7460,N_2019,N_2641);
and U7461 (N_7461,N_429,N_2625);
nand U7462 (N_7462,N_2103,N_2972);
or U7463 (N_7463,N_2949,N_1065);
nor U7464 (N_7464,N_221,N_1808);
nand U7465 (N_7465,N_472,N_3722);
xnor U7466 (N_7466,N_68,N_1109);
xnor U7467 (N_7467,N_911,N_863);
and U7468 (N_7468,N_1519,N_1278);
or U7469 (N_7469,N_3629,N_1888);
or U7470 (N_7470,N_3681,N_1631);
and U7471 (N_7471,N_793,N_2665);
xor U7472 (N_7472,N_1949,N_3023);
nand U7473 (N_7473,N_3448,N_3536);
or U7474 (N_7474,N_2034,N_3574);
or U7475 (N_7475,N_1057,N_3779);
xnor U7476 (N_7476,N_2046,N_1202);
nor U7477 (N_7477,N_853,N_56);
nor U7478 (N_7478,N_1402,N_885);
nor U7479 (N_7479,N_1832,N_1209);
or U7480 (N_7480,N_2095,N_1677);
nand U7481 (N_7481,N_3164,N_556);
xor U7482 (N_7482,N_88,N_2202);
xnor U7483 (N_7483,N_945,N_810);
or U7484 (N_7484,N_2969,N_3383);
xnor U7485 (N_7485,N_2162,N_1453);
nor U7486 (N_7486,N_3223,N_1738);
nand U7487 (N_7487,N_2931,N_537);
nand U7488 (N_7488,N_1481,N_3963);
or U7489 (N_7489,N_385,N_2574);
nor U7490 (N_7490,N_421,N_390);
nor U7491 (N_7491,N_658,N_1563);
nor U7492 (N_7492,N_116,N_2713);
xor U7493 (N_7493,N_3361,N_2737);
and U7494 (N_7494,N_1360,N_1674);
and U7495 (N_7495,N_3536,N_3540);
xor U7496 (N_7496,N_3895,N_3241);
xor U7497 (N_7497,N_573,N_1009);
or U7498 (N_7498,N_3868,N_2240);
nand U7499 (N_7499,N_1813,N_2772);
or U7500 (N_7500,N_1744,N_949);
and U7501 (N_7501,N_1858,N_306);
or U7502 (N_7502,N_3147,N_3798);
nor U7503 (N_7503,N_2175,N_2793);
nor U7504 (N_7504,N_1499,N_286);
nor U7505 (N_7505,N_1781,N_1924);
nand U7506 (N_7506,N_3145,N_2854);
nor U7507 (N_7507,N_2087,N_661);
nand U7508 (N_7508,N_2343,N_3479);
nor U7509 (N_7509,N_0,N_2991);
or U7510 (N_7510,N_237,N_763);
or U7511 (N_7511,N_1074,N_300);
and U7512 (N_7512,N_3438,N_1524);
and U7513 (N_7513,N_3913,N_1110);
and U7514 (N_7514,N_3425,N_1743);
xnor U7515 (N_7515,N_2164,N_2107);
or U7516 (N_7516,N_1735,N_998);
nand U7517 (N_7517,N_57,N_3254);
nor U7518 (N_7518,N_1724,N_2480);
nand U7519 (N_7519,N_1013,N_2199);
and U7520 (N_7520,N_3173,N_2792);
and U7521 (N_7521,N_3513,N_1234);
and U7522 (N_7522,N_2917,N_3367);
or U7523 (N_7523,N_3402,N_1018);
or U7524 (N_7524,N_707,N_3994);
or U7525 (N_7525,N_3470,N_886);
nor U7526 (N_7526,N_322,N_147);
or U7527 (N_7527,N_1055,N_2784);
nand U7528 (N_7528,N_3181,N_3742);
nand U7529 (N_7529,N_1931,N_1314);
nand U7530 (N_7530,N_1706,N_2043);
or U7531 (N_7531,N_1487,N_2895);
or U7532 (N_7532,N_1513,N_2606);
or U7533 (N_7533,N_2673,N_339);
or U7534 (N_7534,N_3081,N_3815);
xor U7535 (N_7535,N_430,N_3289);
and U7536 (N_7536,N_1649,N_2174);
or U7537 (N_7537,N_2783,N_913);
nand U7538 (N_7538,N_3174,N_1247);
xor U7539 (N_7539,N_3594,N_131);
nor U7540 (N_7540,N_3237,N_1555);
nand U7541 (N_7541,N_3375,N_1376);
nor U7542 (N_7542,N_2141,N_2677);
nor U7543 (N_7543,N_301,N_2291);
or U7544 (N_7544,N_2863,N_3218);
nand U7545 (N_7545,N_1469,N_2308);
nor U7546 (N_7546,N_1889,N_2601);
nand U7547 (N_7547,N_3014,N_1644);
nor U7548 (N_7548,N_2500,N_3322);
nand U7549 (N_7549,N_2642,N_2511);
nor U7550 (N_7550,N_949,N_61);
xnor U7551 (N_7551,N_438,N_3204);
and U7552 (N_7552,N_99,N_3270);
nor U7553 (N_7553,N_2773,N_3573);
or U7554 (N_7554,N_628,N_1711);
nand U7555 (N_7555,N_1529,N_211);
and U7556 (N_7556,N_524,N_97);
nor U7557 (N_7557,N_895,N_358);
or U7558 (N_7558,N_2174,N_3592);
nand U7559 (N_7559,N_2231,N_2543);
xor U7560 (N_7560,N_1935,N_3528);
xor U7561 (N_7561,N_3811,N_3195);
nand U7562 (N_7562,N_3512,N_804);
nor U7563 (N_7563,N_1937,N_1944);
nor U7564 (N_7564,N_465,N_1359);
or U7565 (N_7565,N_875,N_2661);
xnor U7566 (N_7566,N_3923,N_2148);
xor U7567 (N_7567,N_15,N_232);
or U7568 (N_7568,N_3085,N_817);
and U7569 (N_7569,N_821,N_3246);
nand U7570 (N_7570,N_1933,N_103);
and U7571 (N_7571,N_467,N_283);
xor U7572 (N_7572,N_2117,N_2798);
and U7573 (N_7573,N_2812,N_3892);
or U7574 (N_7574,N_909,N_654);
nand U7575 (N_7575,N_3682,N_2338);
and U7576 (N_7576,N_1458,N_3326);
nand U7577 (N_7577,N_3737,N_3680);
and U7578 (N_7578,N_3641,N_181);
nand U7579 (N_7579,N_938,N_1683);
nor U7580 (N_7580,N_312,N_2739);
nor U7581 (N_7581,N_512,N_3766);
xnor U7582 (N_7582,N_2407,N_524);
nand U7583 (N_7583,N_3232,N_3127);
nor U7584 (N_7584,N_485,N_2644);
and U7585 (N_7585,N_2944,N_2079);
or U7586 (N_7586,N_2728,N_268);
nand U7587 (N_7587,N_2193,N_77);
and U7588 (N_7588,N_1470,N_1793);
nor U7589 (N_7589,N_3730,N_3818);
and U7590 (N_7590,N_2282,N_2047);
or U7591 (N_7591,N_1845,N_2945);
nand U7592 (N_7592,N_1331,N_879);
xor U7593 (N_7593,N_2266,N_585);
and U7594 (N_7594,N_2530,N_3835);
xnor U7595 (N_7595,N_473,N_1805);
xnor U7596 (N_7596,N_218,N_2708);
or U7597 (N_7597,N_3192,N_3365);
or U7598 (N_7598,N_2197,N_3634);
nor U7599 (N_7599,N_3376,N_131);
xnor U7600 (N_7600,N_779,N_619);
nand U7601 (N_7601,N_1297,N_2513);
and U7602 (N_7602,N_443,N_1590);
nand U7603 (N_7603,N_265,N_1489);
and U7604 (N_7604,N_2823,N_1634);
nand U7605 (N_7605,N_653,N_3812);
xnor U7606 (N_7606,N_3961,N_2416);
nand U7607 (N_7607,N_2348,N_1875);
nand U7608 (N_7608,N_2446,N_45);
nor U7609 (N_7609,N_3474,N_3199);
nor U7610 (N_7610,N_3318,N_3447);
nand U7611 (N_7611,N_3945,N_3201);
xnor U7612 (N_7612,N_3731,N_2787);
nor U7613 (N_7613,N_882,N_3740);
or U7614 (N_7614,N_931,N_582);
nand U7615 (N_7615,N_3701,N_1168);
nand U7616 (N_7616,N_696,N_3666);
or U7617 (N_7617,N_548,N_3127);
xor U7618 (N_7618,N_1729,N_3080);
xnor U7619 (N_7619,N_321,N_505);
nand U7620 (N_7620,N_3460,N_2494);
or U7621 (N_7621,N_3506,N_1730);
and U7622 (N_7622,N_739,N_2560);
and U7623 (N_7623,N_1856,N_795);
nor U7624 (N_7624,N_1144,N_1517);
nor U7625 (N_7625,N_2819,N_2788);
or U7626 (N_7626,N_877,N_2151);
or U7627 (N_7627,N_2790,N_357);
nand U7628 (N_7628,N_2392,N_452);
nor U7629 (N_7629,N_3121,N_26);
and U7630 (N_7630,N_212,N_1189);
xor U7631 (N_7631,N_2613,N_1659);
nor U7632 (N_7632,N_2814,N_2998);
xor U7633 (N_7633,N_3000,N_1889);
nor U7634 (N_7634,N_3368,N_1818);
xnor U7635 (N_7635,N_2686,N_3093);
nand U7636 (N_7636,N_1190,N_2789);
nor U7637 (N_7637,N_3875,N_2241);
nand U7638 (N_7638,N_3160,N_847);
nand U7639 (N_7639,N_2537,N_1870);
or U7640 (N_7640,N_1153,N_492);
xnor U7641 (N_7641,N_1356,N_3588);
nand U7642 (N_7642,N_2559,N_3730);
nand U7643 (N_7643,N_2838,N_1554);
and U7644 (N_7644,N_3241,N_3297);
xnor U7645 (N_7645,N_1092,N_3485);
xor U7646 (N_7646,N_1835,N_1802);
nor U7647 (N_7647,N_350,N_2684);
and U7648 (N_7648,N_3470,N_986);
or U7649 (N_7649,N_1223,N_3386);
or U7650 (N_7650,N_1374,N_711);
and U7651 (N_7651,N_3449,N_3252);
nand U7652 (N_7652,N_983,N_2784);
nor U7653 (N_7653,N_1549,N_2837);
nor U7654 (N_7654,N_1406,N_727);
xor U7655 (N_7655,N_1115,N_1153);
nand U7656 (N_7656,N_923,N_2822);
xnor U7657 (N_7657,N_1442,N_823);
nor U7658 (N_7658,N_506,N_2898);
xor U7659 (N_7659,N_1147,N_2788);
nor U7660 (N_7660,N_342,N_3480);
or U7661 (N_7661,N_2949,N_880);
and U7662 (N_7662,N_2982,N_1052);
nor U7663 (N_7663,N_911,N_1171);
or U7664 (N_7664,N_2281,N_2199);
nand U7665 (N_7665,N_2154,N_3142);
nor U7666 (N_7666,N_1406,N_2132);
nand U7667 (N_7667,N_1647,N_1905);
xnor U7668 (N_7668,N_1567,N_2822);
and U7669 (N_7669,N_3414,N_1760);
nor U7670 (N_7670,N_142,N_3834);
or U7671 (N_7671,N_1433,N_3901);
xor U7672 (N_7672,N_198,N_3989);
and U7673 (N_7673,N_3196,N_499);
or U7674 (N_7674,N_3247,N_1574);
and U7675 (N_7675,N_1804,N_2392);
xor U7676 (N_7676,N_2875,N_2696);
or U7677 (N_7677,N_2346,N_1198);
or U7678 (N_7678,N_849,N_2900);
nand U7679 (N_7679,N_1567,N_945);
and U7680 (N_7680,N_2868,N_112);
nand U7681 (N_7681,N_2901,N_2943);
and U7682 (N_7682,N_1434,N_3751);
xor U7683 (N_7683,N_102,N_126);
or U7684 (N_7684,N_199,N_3032);
xor U7685 (N_7685,N_1376,N_1577);
and U7686 (N_7686,N_1146,N_754);
xor U7687 (N_7687,N_3128,N_450);
and U7688 (N_7688,N_1018,N_119);
or U7689 (N_7689,N_1719,N_1926);
nand U7690 (N_7690,N_2674,N_523);
xnor U7691 (N_7691,N_469,N_3829);
or U7692 (N_7692,N_82,N_3544);
nand U7693 (N_7693,N_2574,N_2655);
nand U7694 (N_7694,N_2487,N_2878);
xor U7695 (N_7695,N_2203,N_3758);
and U7696 (N_7696,N_3652,N_2468);
xnor U7697 (N_7697,N_2041,N_3098);
or U7698 (N_7698,N_2875,N_3389);
and U7699 (N_7699,N_2439,N_3590);
nand U7700 (N_7700,N_3506,N_1280);
nor U7701 (N_7701,N_3844,N_2352);
or U7702 (N_7702,N_1941,N_1650);
and U7703 (N_7703,N_1111,N_262);
nor U7704 (N_7704,N_2145,N_1758);
or U7705 (N_7705,N_2566,N_2299);
nor U7706 (N_7706,N_3856,N_3985);
nor U7707 (N_7707,N_3741,N_1042);
nor U7708 (N_7708,N_1055,N_3088);
or U7709 (N_7709,N_2629,N_494);
nand U7710 (N_7710,N_2508,N_1903);
nand U7711 (N_7711,N_2835,N_790);
nand U7712 (N_7712,N_2997,N_3511);
or U7713 (N_7713,N_353,N_162);
and U7714 (N_7714,N_2151,N_1830);
xnor U7715 (N_7715,N_2019,N_1219);
nand U7716 (N_7716,N_480,N_2522);
or U7717 (N_7717,N_3849,N_1017);
or U7718 (N_7718,N_3906,N_3373);
xor U7719 (N_7719,N_2737,N_3900);
nand U7720 (N_7720,N_3013,N_2732);
and U7721 (N_7721,N_1324,N_2438);
or U7722 (N_7722,N_3231,N_2012);
nand U7723 (N_7723,N_402,N_3361);
xnor U7724 (N_7724,N_1411,N_1280);
and U7725 (N_7725,N_584,N_1004);
xnor U7726 (N_7726,N_611,N_387);
nor U7727 (N_7727,N_3358,N_740);
nand U7728 (N_7728,N_3812,N_2160);
nor U7729 (N_7729,N_867,N_936);
xor U7730 (N_7730,N_2485,N_2986);
nor U7731 (N_7731,N_1184,N_3770);
xor U7732 (N_7732,N_1525,N_1209);
xnor U7733 (N_7733,N_3362,N_451);
and U7734 (N_7734,N_1829,N_2640);
and U7735 (N_7735,N_3942,N_3094);
or U7736 (N_7736,N_603,N_1100);
nand U7737 (N_7737,N_301,N_2605);
or U7738 (N_7738,N_9,N_1613);
or U7739 (N_7739,N_2364,N_2154);
xor U7740 (N_7740,N_1689,N_2602);
nand U7741 (N_7741,N_3904,N_2431);
nand U7742 (N_7742,N_3705,N_770);
and U7743 (N_7743,N_3904,N_1788);
nor U7744 (N_7744,N_2736,N_36);
or U7745 (N_7745,N_506,N_1210);
nor U7746 (N_7746,N_2237,N_2990);
or U7747 (N_7747,N_1653,N_186);
nand U7748 (N_7748,N_498,N_2950);
xnor U7749 (N_7749,N_546,N_1423);
xor U7750 (N_7750,N_351,N_3588);
and U7751 (N_7751,N_3892,N_2792);
or U7752 (N_7752,N_2698,N_1190);
xnor U7753 (N_7753,N_870,N_503);
nor U7754 (N_7754,N_2864,N_120);
or U7755 (N_7755,N_927,N_3805);
xnor U7756 (N_7756,N_3968,N_2638);
nand U7757 (N_7757,N_1190,N_1449);
and U7758 (N_7758,N_3196,N_653);
or U7759 (N_7759,N_3015,N_1712);
xnor U7760 (N_7760,N_629,N_1609);
and U7761 (N_7761,N_819,N_153);
xor U7762 (N_7762,N_2206,N_2754);
and U7763 (N_7763,N_333,N_2220);
and U7764 (N_7764,N_668,N_3792);
or U7765 (N_7765,N_1489,N_297);
nand U7766 (N_7766,N_1539,N_1488);
nand U7767 (N_7767,N_2304,N_2306);
or U7768 (N_7768,N_3040,N_1895);
or U7769 (N_7769,N_2124,N_3045);
or U7770 (N_7770,N_2328,N_1211);
nand U7771 (N_7771,N_1223,N_1484);
and U7772 (N_7772,N_169,N_1226);
or U7773 (N_7773,N_2056,N_638);
xnor U7774 (N_7774,N_2391,N_3506);
nor U7775 (N_7775,N_3908,N_590);
xor U7776 (N_7776,N_3271,N_2685);
or U7777 (N_7777,N_688,N_1113);
and U7778 (N_7778,N_2501,N_1287);
nand U7779 (N_7779,N_854,N_1393);
nor U7780 (N_7780,N_1348,N_2688);
or U7781 (N_7781,N_811,N_3561);
or U7782 (N_7782,N_1328,N_3673);
xor U7783 (N_7783,N_3867,N_2412);
and U7784 (N_7784,N_1057,N_3071);
nor U7785 (N_7785,N_2969,N_48);
xor U7786 (N_7786,N_1374,N_3654);
nor U7787 (N_7787,N_1611,N_2417);
xnor U7788 (N_7788,N_1514,N_983);
nand U7789 (N_7789,N_961,N_2476);
nor U7790 (N_7790,N_3036,N_1094);
nor U7791 (N_7791,N_991,N_63);
nor U7792 (N_7792,N_1871,N_3891);
or U7793 (N_7793,N_1978,N_1102);
xor U7794 (N_7794,N_1123,N_1801);
nand U7795 (N_7795,N_537,N_298);
nor U7796 (N_7796,N_476,N_2104);
or U7797 (N_7797,N_2785,N_1);
nor U7798 (N_7798,N_2880,N_2971);
and U7799 (N_7799,N_1314,N_3596);
or U7800 (N_7800,N_2217,N_749);
nor U7801 (N_7801,N_434,N_1475);
xor U7802 (N_7802,N_2619,N_3928);
nand U7803 (N_7803,N_3552,N_2695);
nand U7804 (N_7804,N_1186,N_584);
xnor U7805 (N_7805,N_1464,N_2574);
xor U7806 (N_7806,N_1067,N_2498);
xnor U7807 (N_7807,N_1233,N_1842);
and U7808 (N_7808,N_2696,N_1571);
nor U7809 (N_7809,N_381,N_454);
nor U7810 (N_7810,N_3614,N_3374);
or U7811 (N_7811,N_3400,N_3490);
or U7812 (N_7812,N_472,N_3582);
xnor U7813 (N_7813,N_1631,N_1428);
or U7814 (N_7814,N_3306,N_2761);
nand U7815 (N_7815,N_1030,N_3524);
and U7816 (N_7816,N_1263,N_3787);
or U7817 (N_7817,N_2134,N_1937);
nand U7818 (N_7818,N_3318,N_276);
nor U7819 (N_7819,N_213,N_1058);
and U7820 (N_7820,N_2583,N_2428);
xor U7821 (N_7821,N_1920,N_2115);
and U7822 (N_7822,N_633,N_2402);
or U7823 (N_7823,N_3225,N_2065);
or U7824 (N_7824,N_286,N_363);
xor U7825 (N_7825,N_1813,N_3141);
xor U7826 (N_7826,N_1602,N_1629);
xnor U7827 (N_7827,N_231,N_576);
nor U7828 (N_7828,N_680,N_2947);
xor U7829 (N_7829,N_1034,N_2717);
and U7830 (N_7830,N_1891,N_848);
and U7831 (N_7831,N_1419,N_3565);
xor U7832 (N_7832,N_372,N_3226);
nand U7833 (N_7833,N_1457,N_338);
and U7834 (N_7834,N_1777,N_2636);
xnor U7835 (N_7835,N_1998,N_663);
xor U7836 (N_7836,N_1314,N_1334);
nor U7837 (N_7837,N_1420,N_2074);
xor U7838 (N_7838,N_2235,N_3938);
nand U7839 (N_7839,N_662,N_2227);
nand U7840 (N_7840,N_3501,N_3156);
and U7841 (N_7841,N_1131,N_3995);
or U7842 (N_7842,N_1961,N_1310);
and U7843 (N_7843,N_1967,N_2047);
nor U7844 (N_7844,N_3425,N_3781);
nor U7845 (N_7845,N_1078,N_1980);
xor U7846 (N_7846,N_3606,N_889);
nor U7847 (N_7847,N_2556,N_2712);
or U7848 (N_7848,N_2374,N_1997);
nand U7849 (N_7849,N_3935,N_3702);
and U7850 (N_7850,N_1452,N_3992);
and U7851 (N_7851,N_444,N_778);
nor U7852 (N_7852,N_1252,N_780);
and U7853 (N_7853,N_3467,N_3295);
and U7854 (N_7854,N_1841,N_3682);
and U7855 (N_7855,N_2157,N_2090);
or U7856 (N_7856,N_888,N_2819);
and U7857 (N_7857,N_1684,N_1504);
xnor U7858 (N_7858,N_2115,N_83);
xor U7859 (N_7859,N_1209,N_2362);
nor U7860 (N_7860,N_14,N_1928);
xor U7861 (N_7861,N_974,N_3004);
xor U7862 (N_7862,N_2107,N_1204);
and U7863 (N_7863,N_1113,N_2120);
nand U7864 (N_7864,N_2754,N_525);
and U7865 (N_7865,N_1528,N_3412);
nor U7866 (N_7866,N_28,N_2183);
nand U7867 (N_7867,N_3345,N_3121);
nor U7868 (N_7868,N_3149,N_1113);
or U7869 (N_7869,N_2411,N_3564);
and U7870 (N_7870,N_2726,N_123);
nor U7871 (N_7871,N_1262,N_3505);
xnor U7872 (N_7872,N_1556,N_3176);
nor U7873 (N_7873,N_2521,N_1767);
nor U7874 (N_7874,N_3115,N_814);
nor U7875 (N_7875,N_984,N_3049);
nand U7876 (N_7876,N_2656,N_1141);
nand U7877 (N_7877,N_2052,N_1999);
nand U7878 (N_7878,N_2604,N_2831);
or U7879 (N_7879,N_3905,N_3416);
or U7880 (N_7880,N_704,N_1750);
or U7881 (N_7881,N_765,N_3584);
nor U7882 (N_7882,N_1027,N_808);
and U7883 (N_7883,N_198,N_1912);
nor U7884 (N_7884,N_2905,N_1824);
or U7885 (N_7885,N_2165,N_3877);
and U7886 (N_7886,N_2256,N_1338);
and U7887 (N_7887,N_850,N_2799);
nor U7888 (N_7888,N_568,N_2579);
nor U7889 (N_7889,N_2662,N_1479);
xnor U7890 (N_7890,N_1803,N_3619);
nor U7891 (N_7891,N_2480,N_3848);
nor U7892 (N_7892,N_2118,N_3634);
nor U7893 (N_7893,N_3905,N_2659);
nor U7894 (N_7894,N_306,N_3658);
xor U7895 (N_7895,N_1452,N_569);
xor U7896 (N_7896,N_321,N_350);
xnor U7897 (N_7897,N_279,N_2672);
xnor U7898 (N_7898,N_905,N_3921);
xnor U7899 (N_7899,N_221,N_2589);
nand U7900 (N_7900,N_1097,N_1556);
or U7901 (N_7901,N_3907,N_1809);
xnor U7902 (N_7902,N_2417,N_2427);
or U7903 (N_7903,N_1903,N_2711);
nand U7904 (N_7904,N_1462,N_2667);
xnor U7905 (N_7905,N_2993,N_1007);
and U7906 (N_7906,N_431,N_3399);
or U7907 (N_7907,N_1803,N_1119);
nand U7908 (N_7908,N_2822,N_3224);
xnor U7909 (N_7909,N_358,N_62);
and U7910 (N_7910,N_3810,N_1364);
or U7911 (N_7911,N_1804,N_2115);
nand U7912 (N_7912,N_3361,N_3465);
nor U7913 (N_7913,N_3538,N_3567);
xnor U7914 (N_7914,N_398,N_618);
and U7915 (N_7915,N_474,N_2585);
and U7916 (N_7916,N_772,N_3204);
nor U7917 (N_7917,N_3035,N_2184);
nor U7918 (N_7918,N_3696,N_1111);
or U7919 (N_7919,N_564,N_3690);
or U7920 (N_7920,N_1881,N_1085);
xnor U7921 (N_7921,N_3161,N_2216);
xor U7922 (N_7922,N_1398,N_2017);
nor U7923 (N_7923,N_1271,N_158);
xor U7924 (N_7924,N_2556,N_3836);
and U7925 (N_7925,N_1073,N_3338);
or U7926 (N_7926,N_2544,N_2196);
nand U7927 (N_7927,N_3252,N_1156);
xnor U7928 (N_7928,N_866,N_2025);
xnor U7929 (N_7929,N_951,N_2824);
and U7930 (N_7930,N_573,N_1485);
nand U7931 (N_7931,N_2433,N_3013);
nor U7932 (N_7932,N_3315,N_2043);
nand U7933 (N_7933,N_3677,N_1041);
and U7934 (N_7934,N_1600,N_2220);
or U7935 (N_7935,N_3279,N_2079);
xnor U7936 (N_7936,N_3793,N_198);
or U7937 (N_7937,N_929,N_2364);
nor U7938 (N_7938,N_3448,N_2703);
or U7939 (N_7939,N_1592,N_2954);
xnor U7940 (N_7940,N_3296,N_568);
nand U7941 (N_7941,N_1541,N_2286);
nand U7942 (N_7942,N_32,N_888);
or U7943 (N_7943,N_2729,N_3973);
or U7944 (N_7944,N_875,N_3175);
or U7945 (N_7945,N_196,N_831);
and U7946 (N_7946,N_279,N_3689);
and U7947 (N_7947,N_177,N_1070);
or U7948 (N_7948,N_826,N_503);
xnor U7949 (N_7949,N_3399,N_1417);
nand U7950 (N_7950,N_863,N_2669);
nor U7951 (N_7951,N_3697,N_3590);
xor U7952 (N_7952,N_1893,N_874);
xor U7953 (N_7953,N_3338,N_517);
and U7954 (N_7954,N_2099,N_1747);
and U7955 (N_7955,N_39,N_1034);
nand U7956 (N_7956,N_2423,N_3524);
nand U7957 (N_7957,N_3478,N_2139);
xor U7958 (N_7958,N_465,N_3731);
nand U7959 (N_7959,N_1240,N_3448);
nor U7960 (N_7960,N_3547,N_3280);
nor U7961 (N_7961,N_958,N_2296);
nand U7962 (N_7962,N_2153,N_1104);
nor U7963 (N_7963,N_2958,N_491);
and U7964 (N_7964,N_2958,N_1380);
and U7965 (N_7965,N_1643,N_1891);
and U7966 (N_7966,N_2175,N_2421);
nor U7967 (N_7967,N_2985,N_3962);
nand U7968 (N_7968,N_3582,N_290);
and U7969 (N_7969,N_3073,N_1623);
and U7970 (N_7970,N_2385,N_257);
nor U7971 (N_7971,N_1689,N_3714);
or U7972 (N_7972,N_1431,N_1566);
and U7973 (N_7973,N_3660,N_350);
or U7974 (N_7974,N_2308,N_2832);
nand U7975 (N_7975,N_3539,N_773);
nor U7976 (N_7976,N_3523,N_697);
or U7977 (N_7977,N_3102,N_1531);
or U7978 (N_7978,N_170,N_2231);
nor U7979 (N_7979,N_2285,N_2382);
and U7980 (N_7980,N_3763,N_2605);
xnor U7981 (N_7981,N_2312,N_1713);
nor U7982 (N_7982,N_217,N_10);
nor U7983 (N_7983,N_992,N_3901);
nand U7984 (N_7984,N_1813,N_495);
nor U7985 (N_7985,N_461,N_35);
nor U7986 (N_7986,N_3895,N_2907);
nand U7987 (N_7987,N_2911,N_3118);
or U7988 (N_7988,N_1587,N_2227);
nor U7989 (N_7989,N_3797,N_1052);
or U7990 (N_7990,N_2868,N_784);
nor U7991 (N_7991,N_1618,N_669);
nand U7992 (N_7992,N_3715,N_466);
xnor U7993 (N_7993,N_2905,N_2654);
and U7994 (N_7994,N_2624,N_2929);
and U7995 (N_7995,N_1202,N_1951);
nand U7996 (N_7996,N_3977,N_1605);
or U7997 (N_7997,N_3367,N_1851);
and U7998 (N_7998,N_3364,N_2224);
xnor U7999 (N_7999,N_217,N_160);
or U8000 (N_8000,N_7941,N_5295);
and U8001 (N_8001,N_7215,N_7739);
and U8002 (N_8002,N_7338,N_6657);
or U8003 (N_8003,N_5839,N_6928);
nor U8004 (N_8004,N_5886,N_6620);
or U8005 (N_8005,N_4590,N_5760);
nor U8006 (N_8006,N_5904,N_5527);
nor U8007 (N_8007,N_4743,N_4558);
or U8008 (N_8008,N_7637,N_4937);
nor U8009 (N_8009,N_5436,N_5265);
xor U8010 (N_8010,N_4854,N_6636);
and U8011 (N_8011,N_7270,N_4389);
nand U8012 (N_8012,N_4894,N_5506);
or U8013 (N_8013,N_7575,N_5223);
xnor U8014 (N_8014,N_4981,N_4461);
and U8015 (N_8015,N_6836,N_5144);
and U8016 (N_8016,N_4507,N_6607);
nand U8017 (N_8017,N_5484,N_6659);
nand U8018 (N_8018,N_7461,N_6751);
or U8019 (N_8019,N_7572,N_7694);
or U8020 (N_8020,N_6197,N_7036);
nand U8021 (N_8021,N_5642,N_6989);
xor U8022 (N_8022,N_7828,N_5028);
and U8023 (N_8023,N_4178,N_4960);
nor U8024 (N_8024,N_4306,N_7288);
and U8025 (N_8025,N_4046,N_6641);
and U8026 (N_8026,N_5941,N_7237);
nor U8027 (N_8027,N_5174,N_4391);
nor U8028 (N_8028,N_4101,N_4739);
nand U8029 (N_8029,N_4261,N_6480);
and U8030 (N_8030,N_5188,N_4893);
xnor U8031 (N_8031,N_6418,N_7540);
and U8032 (N_8032,N_6972,N_5947);
xor U8033 (N_8033,N_5725,N_7538);
nor U8034 (N_8034,N_7160,N_7188);
nor U8035 (N_8035,N_4526,N_6211);
and U8036 (N_8036,N_5175,N_7300);
nor U8037 (N_8037,N_6360,N_7184);
and U8038 (N_8038,N_4976,N_4621);
and U8039 (N_8039,N_6679,N_5117);
or U8040 (N_8040,N_6115,N_6578);
nand U8041 (N_8041,N_4239,N_5385);
nor U8042 (N_8042,N_7445,N_4544);
and U8043 (N_8043,N_4768,N_4908);
and U8044 (N_8044,N_6473,N_4518);
or U8045 (N_8045,N_7214,N_7938);
xor U8046 (N_8046,N_7335,N_5804);
xnor U8047 (N_8047,N_6483,N_4123);
and U8048 (N_8048,N_7043,N_6967);
nor U8049 (N_8049,N_6630,N_4554);
xnor U8050 (N_8050,N_4111,N_5923);
and U8051 (N_8051,N_6691,N_5944);
nor U8052 (N_8052,N_5940,N_7217);
or U8053 (N_8053,N_5691,N_5663);
xor U8054 (N_8054,N_5353,N_6390);
nor U8055 (N_8055,N_6112,N_4135);
xnor U8056 (N_8056,N_6367,N_7148);
nor U8057 (N_8057,N_6369,N_6275);
nand U8058 (N_8058,N_5890,N_7407);
nor U8059 (N_8059,N_6507,N_7636);
nand U8060 (N_8060,N_7859,N_5039);
or U8061 (N_8061,N_6032,N_5778);
and U8062 (N_8062,N_7910,N_5560);
nor U8063 (N_8063,N_4596,N_6531);
or U8064 (N_8064,N_4760,N_4051);
and U8065 (N_8065,N_5370,N_5795);
nor U8066 (N_8066,N_4232,N_7187);
xor U8067 (N_8067,N_5312,N_7563);
nor U8068 (N_8068,N_7852,N_6355);
nand U8069 (N_8069,N_4424,N_5178);
nand U8070 (N_8070,N_6464,N_4578);
nor U8071 (N_8071,N_4494,N_4673);
nand U8072 (N_8072,N_5897,N_4680);
nor U8073 (N_8073,N_5917,N_5196);
nand U8074 (N_8074,N_5679,N_7109);
nand U8075 (N_8075,N_4863,N_7626);
and U8076 (N_8076,N_4065,N_7957);
or U8077 (N_8077,N_7441,N_6109);
nand U8078 (N_8078,N_7380,N_4284);
xnor U8079 (N_8079,N_6138,N_6811);
nand U8080 (N_8080,N_5049,N_4022);
or U8081 (N_8081,N_7586,N_5596);
nor U8082 (N_8082,N_7582,N_7659);
nand U8083 (N_8083,N_5009,N_4551);
or U8084 (N_8084,N_4789,N_6207);
and U8085 (N_8085,N_5414,N_6568);
or U8086 (N_8086,N_5422,N_7012);
nand U8087 (N_8087,N_5038,N_6626);
or U8088 (N_8088,N_7974,N_6297);
xnor U8089 (N_8089,N_7256,N_4514);
xnor U8090 (N_8090,N_6341,N_6669);
xor U8091 (N_8091,N_5936,N_5666);
or U8092 (N_8092,N_4331,N_6897);
or U8093 (N_8093,N_7312,N_7071);
nor U8094 (N_8094,N_7097,N_6218);
or U8095 (N_8095,N_4358,N_5584);
nor U8096 (N_8096,N_7352,N_5930);
nor U8097 (N_8097,N_6075,N_5182);
or U8098 (N_8098,N_4822,N_5736);
nor U8099 (N_8099,N_6071,N_6344);
and U8100 (N_8100,N_5798,N_4546);
and U8101 (N_8101,N_5772,N_4279);
or U8102 (N_8102,N_4699,N_6447);
xnor U8103 (N_8103,N_4532,N_4539);
or U8104 (N_8104,N_5927,N_7499);
xnor U8105 (N_8105,N_7462,N_7606);
nand U8106 (N_8106,N_5045,N_5373);
or U8107 (N_8107,N_6263,N_7922);
nor U8108 (N_8108,N_6181,N_7894);
xor U8109 (N_8109,N_5728,N_5632);
nand U8110 (N_8110,N_7918,N_4502);
nor U8111 (N_8111,N_4865,N_6183);
xnor U8112 (N_8112,N_4687,N_7720);
or U8113 (N_8113,N_7113,N_7088);
and U8114 (N_8114,N_6978,N_7559);
nor U8115 (N_8115,N_6948,N_4052);
nand U8116 (N_8116,N_7459,N_6717);
nand U8117 (N_8117,N_6366,N_7676);
xnor U8118 (N_8118,N_6853,N_6221);
xnor U8119 (N_8119,N_4847,N_4165);
or U8120 (N_8120,N_7703,N_5700);
nor U8121 (N_8121,N_4393,N_7501);
or U8122 (N_8122,N_5483,N_6844);
nand U8123 (N_8123,N_5746,N_4094);
xnor U8124 (N_8124,N_4282,N_4626);
and U8125 (N_8125,N_5456,N_5915);
nand U8126 (N_8126,N_5518,N_4764);
and U8127 (N_8127,N_7610,N_7044);
or U8128 (N_8128,N_7170,N_5934);
nor U8129 (N_8129,N_5368,N_6414);
nand U8130 (N_8130,N_6637,N_6767);
or U8131 (N_8131,N_7144,N_5545);
nand U8132 (N_8132,N_6623,N_5571);
and U8133 (N_8133,N_5163,N_4054);
and U8134 (N_8134,N_4450,N_4812);
and U8135 (N_8135,N_4696,N_6590);
or U8136 (N_8136,N_5346,N_6465);
nand U8137 (N_8137,N_6925,N_6909);
xnor U8138 (N_8138,N_4770,N_5693);
and U8139 (N_8139,N_7701,N_7764);
nor U8140 (N_8140,N_7756,N_6514);
nor U8141 (N_8141,N_7363,N_4669);
or U8142 (N_8142,N_6544,N_6865);
nand U8143 (N_8143,N_5744,N_6233);
xor U8144 (N_8144,N_7372,N_7588);
and U8145 (N_8145,N_7106,N_6765);
xnor U8146 (N_8146,N_6770,N_4096);
and U8147 (N_8147,N_6795,N_5379);
nor U8148 (N_8148,N_7203,N_4308);
nand U8149 (N_8149,N_6371,N_7506);
nand U8150 (N_8150,N_4614,N_6290);
and U8151 (N_8151,N_4221,N_4707);
nor U8152 (N_8152,N_6158,N_4242);
xnor U8153 (N_8153,N_5745,N_6692);
and U8154 (N_8154,N_6908,N_7924);
nor U8155 (N_8155,N_5149,N_5645);
or U8156 (N_8156,N_6624,N_5334);
or U8157 (N_8157,N_5910,N_6838);
nor U8158 (N_8158,N_6815,N_6431);
nor U8159 (N_8159,N_7598,N_7503);
nor U8160 (N_8160,N_6437,N_4993);
nand U8161 (N_8161,N_5701,N_6672);
or U8162 (N_8162,N_5043,N_7241);
xor U8163 (N_8163,N_7309,N_7679);
xnor U8164 (N_8164,N_6269,N_7193);
or U8165 (N_8165,N_5329,N_6884);
xor U8166 (N_8166,N_5668,N_4975);
or U8167 (N_8167,N_5870,N_5986);
nor U8168 (N_8168,N_4860,N_7081);
nand U8169 (N_8169,N_6634,N_4664);
nor U8170 (N_8170,N_7509,N_5249);
xnor U8171 (N_8171,N_7933,N_5577);
or U8172 (N_8172,N_5699,N_5828);
or U8173 (N_8173,N_5046,N_6809);
or U8174 (N_8174,N_4767,N_7954);
xnor U8175 (N_8175,N_5869,N_6089);
xnor U8176 (N_8176,N_7593,N_6270);
nand U8177 (N_8177,N_6654,N_4800);
or U8178 (N_8178,N_4160,N_7020);
xnor U8179 (N_8179,N_5352,N_7349);
nand U8180 (N_8180,N_6528,N_4721);
and U8181 (N_8181,N_4161,N_5752);
xor U8182 (N_8182,N_7523,N_5620);
nor U8183 (N_8183,N_7452,N_6594);
xor U8184 (N_8184,N_5789,N_4697);
or U8185 (N_8185,N_6043,N_7706);
xor U8186 (N_8186,N_7988,N_4049);
or U8187 (N_8187,N_6087,N_5720);
xnor U8188 (N_8188,N_6920,N_4489);
or U8189 (N_8189,N_4216,N_5335);
nand U8190 (N_8190,N_4106,N_7913);
xor U8191 (N_8191,N_7478,N_6813);
nand U8192 (N_8192,N_5777,N_7823);
nand U8193 (N_8193,N_5326,N_5238);
or U8194 (N_8194,N_5523,N_7026);
and U8195 (N_8195,N_5261,N_6790);
xor U8196 (N_8196,N_4375,N_5774);
nand U8197 (N_8197,N_6200,N_4006);
or U8198 (N_8198,N_7614,N_5511);
nand U8199 (N_8199,N_7769,N_6354);
xor U8200 (N_8200,N_4271,N_6533);
nand U8201 (N_8201,N_7695,N_6247);
or U8202 (N_8202,N_5347,N_5431);
nor U8203 (N_8203,N_6176,N_4373);
nor U8204 (N_8204,N_5776,N_5737);
nand U8205 (N_8205,N_5631,N_6913);
and U8206 (N_8206,N_5847,N_6093);
nor U8207 (N_8207,N_4058,N_5874);
or U8208 (N_8208,N_5228,N_5125);
nor U8209 (N_8209,N_5758,N_4897);
xor U8210 (N_8210,N_4370,N_7140);
or U8211 (N_8211,N_7630,N_7060);
nor U8212 (N_8212,N_5389,N_5582);
nor U8213 (N_8213,N_6651,N_7632);
nor U8214 (N_8214,N_7024,N_7644);
nor U8215 (N_8215,N_5189,N_7476);
xnor U8216 (N_8216,N_5826,N_5973);
xnor U8217 (N_8217,N_5980,N_6031);
nand U8218 (N_8218,N_5367,N_4986);
xnor U8219 (N_8219,N_4119,N_4785);
xnor U8220 (N_8220,N_5094,N_6614);
or U8221 (N_8221,N_7774,N_4678);
nand U8222 (N_8222,N_4200,N_5735);
nand U8223 (N_8223,N_4952,N_7866);
or U8224 (N_8224,N_4451,N_4182);
xnor U8225 (N_8225,N_6165,N_4132);
or U8226 (N_8226,N_6723,N_5920);
xnor U8227 (N_8227,N_4835,N_6585);
or U8228 (N_8228,N_4074,N_4333);
and U8229 (N_8229,N_7935,N_7623);
xor U8230 (N_8230,N_5573,N_5697);
xnor U8231 (N_8231,N_5661,N_6021);
and U8232 (N_8232,N_5985,N_5900);
or U8233 (N_8233,N_7487,N_6244);
or U8234 (N_8234,N_6224,N_6264);
xnor U8235 (N_8235,N_5682,N_7277);
nor U8236 (N_8236,N_7420,N_7273);
nand U8237 (N_8237,N_6326,N_4433);
xor U8238 (N_8238,N_4662,N_7987);
nor U8239 (N_8239,N_5893,N_5921);
or U8240 (N_8240,N_5868,N_5112);
nand U8241 (N_8241,N_6532,N_4979);
xor U8242 (N_8242,N_7732,N_6294);
or U8243 (N_8243,N_5763,N_7443);
and U8244 (N_8244,N_5757,N_7371);
or U8245 (N_8245,N_4076,N_6364);
nor U8246 (N_8246,N_4268,N_7154);
nor U8247 (N_8247,N_7504,N_4519);
nand U8248 (N_8248,N_7816,N_5124);
nor U8249 (N_8249,N_4487,N_7172);
and U8250 (N_8250,N_6508,N_5686);
nor U8251 (N_8251,N_5994,N_6822);
xnor U8252 (N_8252,N_7591,N_4517);
and U8253 (N_8253,N_7661,N_4215);
xnor U8254 (N_8254,N_4134,N_6454);
nor U8255 (N_8255,N_7440,N_4043);
nor U8256 (N_8256,N_4350,N_5954);
or U8257 (N_8257,N_4409,N_6420);
and U8258 (N_8258,N_7307,N_6864);
nand U8259 (N_8259,N_4326,N_5794);
nand U8260 (N_8260,N_5041,N_7920);
nand U8261 (N_8261,N_5628,N_6322);
nor U8262 (N_8262,N_7495,N_6889);
xor U8263 (N_8263,N_5327,N_4925);
and U8264 (N_8264,N_5190,N_6100);
nor U8265 (N_8265,N_7693,N_6567);
or U8266 (N_8266,N_5222,N_7683);
nor U8267 (N_8267,N_6756,N_6504);
and U8268 (N_8268,N_7233,N_6803);
nor U8269 (N_8269,N_6015,N_5572);
or U8270 (N_8270,N_6764,N_4116);
or U8271 (N_8271,N_5110,N_4412);
nor U8272 (N_8272,N_6379,N_6957);
nand U8273 (N_8273,N_5416,N_6539);
or U8274 (N_8274,N_5053,N_5226);
xnor U8275 (N_8275,N_4066,N_7386);
and U8276 (N_8276,N_7391,N_5817);
nor U8277 (N_8277,N_7865,N_6748);
and U8278 (N_8278,N_6951,N_4668);
nor U8279 (N_8279,N_7361,N_5204);
or U8280 (N_8280,N_7677,N_5215);
xor U8281 (N_8281,N_6314,N_7741);
xnor U8282 (N_8282,N_5294,N_4813);
xnor U8283 (N_8283,N_7378,N_6313);
nand U8284 (N_8284,N_5998,N_5296);
nand U8285 (N_8285,N_7670,N_7547);
nand U8286 (N_8286,N_7416,N_5280);
xor U8287 (N_8287,N_7156,N_4646);
xor U8288 (N_8288,N_5165,N_5195);
nand U8289 (N_8289,N_4024,N_7743);
nand U8290 (N_8290,N_5221,N_4900);
nor U8291 (N_8291,N_6148,N_4228);
nand U8292 (N_8292,N_7903,N_4613);
and U8293 (N_8293,N_5270,N_4862);
and U8294 (N_8294,N_5621,N_4769);
xor U8295 (N_8295,N_4458,N_6052);
nor U8296 (N_8296,N_4164,N_4851);
nor U8297 (N_8297,N_4432,N_7771);
and U8298 (N_8298,N_4725,N_6734);
nor U8299 (N_8299,N_7834,N_5486);
or U8300 (N_8300,N_5465,N_4758);
xnor U8301 (N_8301,N_5820,N_6240);
xnor U8302 (N_8302,N_6016,N_7004);
xor U8303 (N_8303,N_6582,N_4513);
and U8304 (N_8304,N_4700,N_4062);
or U8305 (N_8305,N_7114,N_6094);
nor U8306 (N_8306,N_5521,N_5922);
or U8307 (N_8307,N_7736,N_5888);
or U8308 (N_8308,N_5674,N_5318);
nor U8309 (N_8309,N_5611,N_4766);
xor U8310 (N_8310,N_5528,N_6296);
nor U8311 (N_8311,N_5997,N_5481);
nor U8312 (N_8312,N_7993,N_5304);
and U8313 (N_8313,N_5533,N_4332);
nor U8314 (N_8314,N_5770,N_5390);
nor U8315 (N_8315,N_6556,N_4014);
xor U8316 (N_8316,N_4837,N_4434);
nor U8317 (N_8317,N_6571,N_5931);
xor U8318 (N_8318,N_4886,N_5371);
or U8319 (N_8319,N_4728,N_5507);
nor U8320 (N_8320,N_4522,N_7339);
nor U8321 (N_8321,N_7464,N_7931);
and U8322 (N_8322,N_4418,N_7327);
nand U8323 (N_8323,N_5741,N_7139);
or U8324 (N_8324,N_4642,N_7009);
or U8325 (N_8325,N_7599,N_4070);
and U8326 (N_8326,N_5858,N_4152);
and U8327 (N_8327,N_6226,N_6061);
xor U8328 (N_8328,N_7134,N_6219);
and U8329 (N_8329,N_4500,N_6635);
nand U8330 (N_8330,N_4672,N_4984);
xnor U8331 (N_8331,N_7342,N_6416);
nand U8332 (N_8332,N_4419,N_4638);
or U8333 (N_8333,N_7448,N_4644);
or U8334 (N_8334,N_6168,N_4968);
nand U8335 (N_8335,N_4238,N_4328);
xnor U8336 (N_8336,N_7098,N_5076);
and U8337 (N_8337,N_4869,N_4653);
and U8338 (N_8338,N_7246,N_4749);
xor U8339 (N_8339,N_6410,N_7212);
and U8340 (N_8340,N_4220,N_7616);
or U8341 (N_8341,N_5199,N_4751);
or U8342 (N_8342,N_6698,N_6793);
nand U8343 (N_8343,N_7486,N_7287);
xnor U8344 (N_8344,N_4969,N_4225);
or U8345 (N_8345,N_7209,N_6388);
nand U8346 (N_8346,N_6317,N_6505);
nand U8347 (N_8347,N_4151,N_7469);
nand U8348 (N_8348,N_7734,N_4741);
nor U8349 (N_8349,N_4942,N_4137);
nor U8350 (N_8350,N_6337,N_6118);
xor U8351 (N_8351,N_5830,N_6543);
and U8352 (N_8352,N_4531,N_7123);
and U8353 (N_8353,N_7992,N_4097);
or U8354 (N_8354,N_6991,N_6586);
or U8355 (N_8355,N_6903,N_7733);
nor U8356 (N_8356,N_5365,N_7620);
nor U8357 (N_8357,N_5877,N_5609);
nor U8358 (N_8358,N_6904,N_5970);
or U8359 (N_8359,N_5495,N_6816);
and U8360 (N_8360,N_6945,N_6716);
nor U8361 (N_8361,N_5432,N_7658);
nor U8362 (N_8362,N_4559,N_4223);
nand U8363 (N_8363,N_7375,N_4730);
nand U8364 (N_8364,N_6339,N_7937);
nand U8365 (N_8365,N_6194,N_6984);
or U8366 (N_8366,N_5861,N_7249);
nor U8367 (N_8367,N_6861,N_7169);
xnor U8368 (N_8368,N_5756,N_4472);
nor U8369 (N_8369,N_5767,N_4501);
or U8370 (N_8370,N_6246,N_5059);
nor U8371 (N_8371,N_5077,N_6882);
and U8372 (N_8372,N_6996,N_4219);
and U8373 (N_8373,N_7498,N_4368);
nor U8374 (N_8374,N_5148,N_6726);
nand U8375 (N_8375,N_4427,N_7612);
xnor U8376 (N_8376,N_6936,N_6135);
and U8377 (N_8377,N_6029,N_6564);
and U8378 (N_8378,N_7773,N_4192);
xor U8379 (N_8379,N_4950,N_6085);
nor U8380 (N_8380,N_6137,N_6126);
or U8381 (N_8381,N_5090,N_7532);
and U8382 (N_8382,N_6092,N_7345);
nand U8383 (N_8383,N_6959,N_5082);
nand U8384 (N_8384,N_6640,N_7735);
xnor U8385 (N_8385,N_6828,N_6417);
and U8386 (N_8386,N_5173,N_5616);
and U8387 (N_8387,N_5372,N_5843);
xor U8388 (N_8388,N_7709,N_7867);
nand U8389 (N_8389,N_5299,N_6274);
and U8390 (N_8390,N_4019,N_5286);
and U8391 (N_8391,N_4631,N_7171);
or U8392 (N_8392,N_6729,N_6325);
or U8393 (N_8393,N_5999,N_6592);
xor U8394 (N_8394,N_7979,N_6744);
xor U8395 (N_8395,N_6549,N_7763);
nor U8396 (N_8396,N_6724,N_4297);
nand U8397 (N_8397,N_5171,N_4480);
and U8398 (N_8398,N_4289,N_4752);
or U8399 (N_8399,N_6699,N_6358);
or U8400 (N_8400,N_7853,N_7124);
nand U8401 (N_8401,N_5780,N_6057);
nor U8402 (N_8402,N_6214,N_6099);
or U8403 (N_8403,N_5988,N_5054);
nand U8404 (N_8404,N_4740,N_7267);
nand U8405 (N_8405,N_6587,N_6510);
or U8406 (N_8406,N_5557,N_7727);
or U8407 (N_8407,N_4444,N_6456);
nand U8408 (N_8408,N_4157,N_7365);
xor U8409 (N_8409,N_4233,N_7279);
and U8410 (N_8410,N_7211,N_5946);
and U8411 (N_8411,N_5751,N_4658);
nor U8412 (N_8412,N_6799,N_7989);
nand U8413 (N_8413,N_5978,N_7624);
nand U8414 (N_8414,N_4612,N_4719);
and U8415 (N_8415,N_5233,N_6164);
and U8416 (N_8416,N_7467,N_5979);
nor U8417 (N_8417,N_4711,N_5241);
xnor U8418 (N_8418,N_4938,N_7404);
nand U8419 (N_8419,N_4247,N_7149);
nand U8420 (N_8420,N_5837,N_7016);
xor U8421 (N_8421,N_6067,N_4523);
or U8422 (N_8422,N_5383,N_5969);
nand U8423 (N_8423,N_7596,N_5738);
xnor U8424 (N_8424,N_7565,N_5101);
nand U8425 (N_8425,N_7711,N_4377);
nor U8426 (N_8426,N_6139,N_5502);
nor U8427 (N_8427,N_6956,N_4727);
or U8428 (N_8428,N_7500,N_4540);
and U8429 (N_8429,N_7055,N_7647);
or U8430 (N_8430,N_7994,N_4398);
xor U8431 (N_8431,N_6848,N_6445);
nand U8432 (N_8432,N_7765,N_7655);
nand U8433 (N_8433,N_4899,N_7179);
xnor U8434 (N_8434,N_7900,N_7873);
nor U8435 (N_8435,N_5583,N_4557);
nand U8436 (N_8436,N_6080,N_5659);
nand U8437 (N_8437,N_7602,N_7926);
and U8438 (N_8438,N_7454,N_6512);
nand U8439 (N_8439,N_4748,N_5435);
or U8440 (N_8440,N_7529,N_5032);
xor U8441 (N_8441,N_4124,N_4805);
xnor U8442 (N_8442,N_6715,N_6804);
xor U8443 (N_8443,N_5578,N_7904);
xor U8444 (N_8444,N_5865,N_4195);
nor U8445 (N_8445,N_4277,N_5179);
xnor U8446 (N_8446,N_6867,N_5643);
and U8447 (N_8447,N_6312,N_4920);
xor U8448 (N_8448,N_4294,N_5216);
or U8449 (N_8449,N_4599,N_6947);
nand U8450 (N_8450,N_4484,N_5575);
or U8451 (N_8451,N_5727,N_4462);
or U8452 (N_8452,N_4831,N_6642);
nand U8453 (N_8453,N_5587,N_6428);
nor U8454 (N_8454,N_6849,N_7493);
or U8455 (N_8455,N_4230,N_5321);
or U8456 (N_8456,N_5162,N_7609);
and U8457 (N_8457,N_4428,N_4413);
nor U8458 (N_8458,N_6045,N_7811);
nand U8459 (N_8459,N_5311,N_6072);
xnor U8460 (N_8460,N_4144,N_6459);
nor U8461 (N_8461,N_6468,N_4998);
nand U8462 (N_8462,N_4488,N_5717);
xnor U8463 (N_8463,N_5463,N_4804);
nand U8464 (N_8464,N_6593,N_5272);
nor U8465 (N_8465,N_5333,N_5019);
nand U8466 (N_8466,N_5884,N_7185);
and U8467 (N_8467,N_4840,N_7668);
nand U8468 (N_8468,N_5879,N_5419);
nand U8469 (N_8469,N_4643,N_6040);
nor U8470 (N_8470,N_4198,N_5702);
nor U8471 (N_8471,N_6887,N_4781);
nand U8472 (N_8472,N_7052,N_7408);
nor U8473 (N_8473,N_4009,N_5906);
nand U8474 (N_8474,N_4112,N_5601);
nand U8475 (N_8475,N_7178,N_6303);
nand U8476 (N_8476,N_4218,N_4909);
nor U8477 (N_8477,N_4545,N_4262);
nand U8478 (N_8478,N_5395,N_6345);
or U8479 (N_8479,N_6186,N_6022);
xor U8480 (N_8480,N_5084,N_4567);
xor U8481 (N_8481,N_4628,N_4846);
or U8482 (N_8482,N_6287,N_4237);
nor U8483 (N_8483,N_5651,N_5867);
and U8484 (N_8484,N_6150,N_5472);
nand U8485 (N_8485,N_6814,N_6631);
and U8486 (N_8486,N_4275,N_7022);
nand U8487 (N_8487,N_4026,N_5662);
nand U8488 (N_8488,N_7562,N_5950);
xor U8489 (N_8489,N_4285,N_4324);
and U8490 (N_8490,N_5277,N_7791);
nand U8491 (N_8491,N_5812,N_5600);
nor U8492 (N_8492,N_6033,N_7250);
nor U8493 (N_8493,N_7990,N_4746);
nor U8494 (N_8494,N_7227,N_6788);
and U8495 (N_8495,N_4129,N_5547);
nor U8496 (N_8496,N_5857,N_4474);
nand U8497 (N_8497,N_5656,N_5871);
nand U8498 (N_8498,N_4027,N_7438);
nor U8499 (N_8499,N_5360,N_7162);
nor U8500 (N_8500,N_7949,N_4961);
or U8501 (N_8501,N_7389,N_5166);
nand U8502 (N_8502,N_5153,N_6857);
nor U8503 (N_8503,N_4053,N_4372);
and U8504 (N_8504,N_7678,N_7087);
xor U8505 (N_8505,N_7387,N_6516);
or U8506 (N_8506,N_4390,N_4356);
xnor U8507 (N_8507,N_4603,N_7611);
and U8508 (N_8508,N_6190,N_4803);
xnor U8509 (N_8509,N_4127,N_7810);
and U8510 (N_8510,N_7056,N_4498);
and U8511 (N_8511,N_4826,N_7579);
nor U8512 (N_8512,N_7671,N_7700);
and U8513 (N_8513,N_6271,N_4924);
or U8514 (N_8514,N_6036,N_6488);
xnor U8515 (N_8515,N_6173,N_6975);
and U8516 (N_8516,N_5018,N_6565);
and U8517 (N_8517,N_5485,N_6937);
xnor U8518 (N_8518,N_6854,N_5989);
or U8519 (N_8519,N_4139,N_4455);
nand U8520 (N_8520,N_4061,N_6604);
nand U8521 (N_8521,N_5325,N_6230);
xor U8522 (N_8522,N_6704,N_4943);
or U8523 (N_8523,N_4177,N_5551);
and U8524 (N_8524,N_4354,N_6974);
xnor U8525 (N_8525,N_5909,N_4257);
nor U8526 (N_8526,N_5191,N_5493);
nor U8527 (N_8527,N_4429,N_6621);
xor U8528 (N_8528,N_7639,N_6633);
nand U8529 (N_8529,N_5681,N_5302);
nand U8530 (N_8530,N_7437,N_6537);
or U8531 (N_8531,N_7278,N_5017);
xor U8532 (N_8532,N_5324,N_4399);
or U8533 (N_8533,N_7833,N_7463);
and U8534 (N_8534,N_5480,N_4890);
and U8535 (N_8535,N_4003,N_6761);
nor U8536 (N_8536,N_7061,N_5487);
or U8537 (N_8537,N_4184,N_7234);
and U8538 (N_8538,N_6665,N_4888);
nand U8539 (N_8539,N_5550,N_5088);
xnor U8540 (N_8540,N_5791,N_6935);
xnor U8541 (N_8541,N_4449,N_6353);
and U8542 (N_8542,N_4201,N_4337);
xnor U8543 (N_8543,N_6840,N_7003);
nand U8544 (N_8544,N_6824,N_7785);
xor U8545 (N_8545,N_7316,N_5391);
or U8546 (N_8546,N_5186,N_7550);
xor U8547 (N_8547,N_6306,N_5743);
and U8548 (N_8548,N_6966,N_6286);
and U8549 (N_8549,N_7294,N_4892);
nor U8550 (N_8550,N_4168,N_4880);
nand U8551 (N_8551,N_4755,N_4330);
nor U8552 (N_8552,N_4577,N_6215);
xnor U8553 (N_8553,N_4042,N_7450);
or U8554 (N_8554,N_5846,N_4790);
nand U8555 (N_8555,N_7073,N_6132);
or U8556 (N_8556,N_7830,N_7397);
or U8557 (N_8557,N_7128,N_5114);
and U8558 (N_8558,N_6442,N_6602);
nor U8559 (N_8559,N_5349,N_5409);
xor U8560 (N_8560,N_6953,N_7761);
and U8561 (N_8561,N_7323,N_4542);
and U8562 (N_8562,N_4876,N_6900);
and U8563 (N_8563,N_6648,N_4296);
xor U8564 (N_8564,N_4564,N_7680);
and U8565 (N_8565,N_4176,N_7719);
nand U8566 (N_8566,N_4798,N_6285);
or U8567 (N_8567,N_5818,N_7266);
nand U8568 (N_8568,N_5508,N_5517);
and U8569 (N_8569,N_5627,N_5853);
and U8570 (N_8570,N_4447,N_4110);
or U8571 (N_8571,N_6359,N_7152);
and U8572 (N_8572,N_7320,N_7977);
nand U8573 (N_8573,N_6450,N_5119);
xnor U8574 (N_8574,N_4606,N_7164);
xnor U8575 (N_8575,N_6127,N_6791);
nand U8576 (N_8576,N_6128,N_5712);
nor U8577 (N_8577,N_6477,N_7130);
or U8578 (N_8578,N_5862,N_4410);
xor U8579 (N_8579,N_4479,N_5561);
xnor U8580 (N_8580,N_5929,N_7191);
nand U8581 (N_8581,N_7804,N_4553);
xor U8582 (N_8582,N_6969,N_4154);
or U8583 (N_8583,N_4015,N_6346);
or U8584 (N_8584,N_5714,N_4209);
nor U8585 (N_8585,N_6710,N_4990);
or U8586 (N_8586,N_5845,N_4885);
and U8587 (N_8587,N_5881,N_4425);
nor U8588 (N_8588,N_7228,N_4273);
and U8589 (N_8589,N_7400,N_7888);
nand U8590 (N_8590,N_6676,N_6013);
and U8591 (N_8591,N_4274,N_7255);
nand U8592 (N_8592,N_7673,N_5255);
and U8593 (N_8593,N_4955,N_4105);
xor U8594 (N_8594,N_6235,N_7293);
nor U8595 (N_8595,N_5058,N_7886);
nand U8596 (N_8596,N_7812,N_7784);
nand U8597 (N_8597,N_6812,N_5694);
nor U8598 (N_8598,N_5821,N_6147);
nor U8599 (N_8599,N_5220,N_7264);
nand U8600 (N_8600,N_4204,N_4102);
nor U8601 (N_8601,N_4689,N_4555);
xnor U8602 (N_8602,N_6133,N_6035);
or U8603 (N_8603,N_5548,N_6740);
nand U8604 (N_8604,N_4276,N_6088);
nor U8605 (N_8605,N_5636,N_6911);
xnor U8606 (N_8606,N_6509,N_5438);
or U8607 (N_8607,N_5317,N_6662);
nand U8608 (N_8608,N_4453,N_7502);
and U8609 (N_8609,N_6149,N_4683);
or U8610 (N_8610,N_6577,N_5254);
or U8611 (N_8611,N_5382,N_7813);
nand U8612 (N_8612,N_7961,N_6860);
nor U8613 (N_8613,N_4763,N_5585);
or U8614 (N_8614,N_7135,N_7567);
or U8615 (N_8615,N_4343,N_4670);
and U8616 (N_8616,N_7200,N_5309);
xnor U8617 (N_8617,N_5671,N_4923);
and U8618 (N_8618,N_6178,N_7433);
and U8619 (N_8619,N_5555,N_6649);
or U8620 (N_8620,N_7369,N_4988);
or U8621 (N_8621,N_6439,N_6919);
nor U8622 (N_8622,N_5423,N_4903);
nor U8623 (N_8623,N_4688,N_7229);
nand U8624 (N_8624,N_5398,N_6627);
or U8625 (N_8625,N_5048,N_6167);
xnor U8626 (N_8626,N_4948,N_4619);
xor U8627 (N_8627,N_7986,N_7422);
xor U8628 (N_8628,N_4383,N_5181);
nor U8629 (N_8629,N_6695,N_6111);
xor U8630 (N_8630,N_5568,N_6489);
xor U8631 (N_8631,N_6288,N_7645);
and U8632 (N_8632,N_6625,N_7295);
nand U8633 (N_8633,N_4405,N_5943);
nand U8634 (N_8634,N_5099,N_4156);
and U8635 (N_8635,N_6688,N_5851);
or U8636 (N_8636,N_7402,N_7984);
nor U8637 (N_8637,N_6758,N_5836);
nand U8638 (N_8638,N_4910,N_7482);
and U8639 (N_8639,N_7945,N_4008);
nand U8640 (N_8640,N_7274,N_4874);
nor U8641 (N_8641,N_6242,N_6229);
xor U8642 (N_8642,N_7790,N_7808);
xnor U8643 (N_8643,N_7651,N_4757);
nor U8644 (N_8644,N_7181,N_4547);
nand U8645 (N_8645,N_6192,N_5580);
and U8646 (N_8646,N_7410,N_6693);
or U8647 (N_8647,N_6024,N_5429);
nor U8648 (N_8648,N_6171,N_5381);
xnor U8649 (N_8649,N_6601,N_7231);
nor U8650 (N_8650,N_6332,N_4591);
nor U8651 (N_8651,N_5130,N_5460);
nor U8652 (N_8652,N_5338,N_5387);
nor U8653 (N_8653,N_6628,N_7822);
or U8654 (N_8654,N_4293,N_6960);
nand U8655 (N_8655,N_7068,N_6703);
or U8656 (N_8656,N_4717,N_5342);
nand U8657 (N_8657,N_6284,N_5499);
and U8658 (N_8658,N_6709,N_5875);
xor U8659 (N_8659,N_7199,N_7507);
nor U8660 (N_8660,N_6182,N_5003);
and U8661 (N_8661,N_5469,N_5301);
nand U8662 (N_8662,N_4824,N_6058);
xnor U8663 (N_8663,N_5996,N_5503);
nor U8664 (N_8664,N_7515,N_6906);
xnor U8665 (N_8665,N_4287,N_6892);
nor U8666 (N_8666,N_4944,N_6478);
nor U8667 (N_8667,N_6546,N_6689);
nand U8668 (N_8668,N_5337,N_7561);
xor U8669 (N_8669,N_4213,N_5993);
nor U8670 (N_8670,N_4845,N_7749);
xor U8671 (N_8671,N_5313,N_5602);
and U8672 (N_8672,N_7334,N_5284);
nor U8673 (N_8673,N_5765,N_5995);
and U8674 (N_8674,N_6774,N_5723);
or U8675 (N_8675,N_5402,N_5650);
nand U8676 (N_8676,N_4774,N_6259);
and U8677 (N_8677,N_7017,N_4067);
nand U8678 (N_8678,N_6434,N_7354);
and U8679 (N_8679,N_6658,N_5732);
xnor U8680 (N_8680,N_5375,N_5087);
nand U8681 (N_8681,N_5914,N_6277);
xor U8682 (N_8682,N_5913,N_5004);
or U8683 (N_8683,N_4045,N_5844);
or U8684 (N_8684,N_5462,N_5142);
and U8685 (N_8685,N_7432,N_7014);
nor U8686 (N_8686,N_4964,N_7878);
xor U8687 (N_8687,N_6159,N_4448);
nand U8688 (N_8688,N_5677,N_4347);
xor U8689 (N_8689,N_6515,N_6881);
nor U8690 (N_8690,N_4159,N_6090);
nand U8691 (N_8691,N_4972,N_6706);
or U8692 (N_8692,N_7091,N_4821);
nor U8693 (N_8693,N_7348,N_7254);
nand U8694 (N_8694,N_7667,N_6548);
nand U8695 (N_8695,N_6643,N_5007);
nand U8696 (N_8696,N_5433,N_7782);
and U8697 (N_8697,N_5137,N_4457);
nor U8698 (N_8698,N_7556,N_5690);
xnor U8699 (N_8699,N_7663,N_4303);
xor U8700 (N_8700,N_7455,N_5399);
xnor U8701 (N_8701,N_7851,N_7326);
xnor U8702 (N_8702,N_5589,N_4878);
nand U8703 (N_8703,N_7196,N_4208);
xor U8704 (N_8704,N_5451,N_6843);
nand U8705 (N_8705,N_7689,N_5707);
and U8706 (N_8706,N_6771,N_6850);
and U8707 (N_8707,N_7662,N_6941);
nand U8708 (N_8708,N_6597,N_7037);
and U8709 (N_8709,N_4153,N_4166);
and U8710 (N_8710,N_5626,N_6255);
and U8711 (N_8711,N_6405,N_7789);
nand U8712 (N_8712,N_4364,N_5939);
and U8713 (N_8713,N_5143,N_4666);
nor U8714 (N_8714,N_7265,N_4468);
xnor U8715 (N_8715,N_5885,N_6191);
nand U8716 (N_8716,N_6839,N_7724);
nand U8717 (N_8717,N_5273,N_4568);
or U8718 (N_8718,N_5247,N_7893);
xor U8719 (N_8719,N_7872,N_6102);
nor U8720 (N_8720,N_6361,N_4205);
and U8721 (N_8721,N_6595,N_4870);
and U8722 (N_8722,N_7831,N_5544);
nand U8723 (N_8723,N_4508,N_4315);
nor U8724 (N_8724,N_5648,N_7390);
and U8725 (N_8725,N_7141,N_5948);
xnor U8726 (N_8726,N_4100,N_6712);
nor U8727 (N_8727,N_6097,N_7373);
and U8728 (N_8728,N_5298,N_7634);
nand U8729 (N_8729,N_7580,N_6964);
xor U8730 (N_8730,N_5030,N_7111);
nor U8731 (N_8731,N_4973,N_4141);
and U8732 (N_8732,N_7600,N_4772);
xor U8733 (N_8733,N_7018,N_6566);
nor U8734 (N_8734,N_5721,N_6939);
and U8735 (N_8735,N_4320,N_5020);
and U8736 (N_8736,N_4685,N_7403);
nand U8737 (N_8737,N_4260,N_6776);
nor U8738 (N_8738,N_7031,N_5932);
nand U8739 (N_8739,N_7105,N_4575);
nand U8740 (N_8740,N_5768,N_5849);
nand U8741 (N_8741,N_5805,N_7934);
xor U8742 (N_8742,N_5305,N_5797);
nor U8743 (N_8743,N_7521,N_4828);
nand U8744 (N_8744,N_6012,N_7082);
nor U8745 (N_8745,N_4207,N_6462);
nand U8746 (N_8746,N_6823,N_5957);
or U8747 (N_8747,N_6307,N_4871);
and U8748 (N_8748,N_6797,N_4630);
xor U8749 (N_8749,N_6563,N_6146);
nor U8750 (N_8750,N_4313,N_6476);
xnor U8751 (N_8751,N_5928,N_6081);
and U8752 (N_8752,N_6293,N_4736);
xnor U8753 (N_8753,N_4570,N_4524);
xnor U8754 (N_8754,N_6372,N_4556);
xnor U8755 (N_8755,N_4742,N_5467);
nor U8756 (N_8756,N_6260,N_4637);
nand U8757 (N_8757,N_5477,N_6409);
nand U8758 (N_8758,N_4902,N_5831);
nand U8759 (N_8759,N_6030,N_6373);
nor U8760 (N_8760,N_7447,N_5376);
xor U8761 (N_8761,N_6407,N_7589);
xnor U8762 (N_8762,N_5308,N_5185);
xnor U8763 (N_8763,N_4808,N_5673);
nor U8764 (N_8764,N_5581,N_5066);
or U8765 (N_8765,N_4629,N_7535);
xor U8766 (N_8766,N_4675,N_7158);
or U8767 (N_8767,N_7282,N_5275);
xnor U8768 (N_8768,N_4471,N_5095);
nand U8769 (N_8769,N_4565,N_5633);
or U8770 (N_8770,N_7877,N_4396);
nor U8771 (N_8771,N_4401,N_4493);
nor U8772 (N_8772,N_7622,N_4844);
nor U8773 (N_8773,N_6223,N_5734);
or U8774 (N_8774,N_5242,N_5443);
or U8775 (N_8775,N_7021,N_7836);
and U8776 (N_8776,N_6647,N_5647);
and U8777 (N_8777,N_5310,N_5688);
nand U8778 (N_8778,N_4784,N_6042);
nand U8779 (N_8779,N_7898,N_4175);
xor U8780 (N_8780,N_6119,N_5963);
xnor U8781 (N_8781,N_7190,N_4187);
nor U8782 (N_8782,N_7496,N_5106);
nand U8783 (N_8783,N_5013,N_5990);
nand U8784 (N_8784,N_4702,N_7511);
or U8785 (N_8785,N_5501,N_6847);
xor U8786 (N_8786,N_4416,N_7649);
xnor U8787 (N_8787,N_5078,N_4252);
nor U8788 (N_8788,N_4316,N_6385);
or U8789 (N_8789,N_7965,N_5512);
and U8790 (N_8790,N_5854,N_4958);
xnor U8791 (N_8791,N_7223,N_6261);
nand U8792 (N_8792,N_7051,N_7730);
or U8793 (N_8793,N_5992,N_7078);
and U8794 (N_8794,N_6440,N_7539);
or U8795 (N_8795,N_5590,N_4934);
or U8796 (N_8796,N_5113,N_4953);
and U8797 (N_8797,N_5239,N_6041);
and U8798 (N_8798,N_7120,N_7850);
xnor U8799 (N_8799,N_4810,N_6541);
xnor U8800 (N_8800,N_6965,N_5654);
and U8801 (N_8801,N_5937,N_5695);
xnor U8802 (N_8802,N_6561,N_5665);
nand U8803 (N_8803,N_7869,N_4657);
nor U8804 (N_8804,N_7409,N_4534);
nor U8805 (N_8805,N_5307,N_4317);
or U8806 (N_8806,N_4283,N_6156);
xnor U8807 (N_8807,N_7122,N_4704);
and U8808 (N_8808,N_6513,N_5724);
xor U8809 (N_8809,N_7543,N_5634);
nand U8810 (N_8810,N_5361,N_7980);
nor U8811 (N_8811,N_7881,N_6963);
or U8812 (N_8812,N_5593,N_4801);
xnor U8813 (N_8813,N_6324,N_7220);
xnor U8814 (N_8814,N_4571,N_6023);
nand U8815 (N_8815,N_4510,N_5675);
nand U8816 (N_8816,N_6020,N_6955);
or U8817 (N_8817,N_5172,N_6392);
or U8818 (N_8818,N_4486,N_6694);
nor U8819 (N_8819,N_4005,N_6001);
xnor U8820 (N_8820,N_4466,N_7396);
and U8821 (N_8821,N_4980,N_4623);
nor U8822 (N_8822,N_7685,N_7202);
xnor U8823 (N_8823,N_6588,N_6292);
nor U8824 (N_8824,N_4355,N_5448);
nor U8825 (N_8825,N_4738,N_7174);
or U8826 (N_8826,N_5863,N_6419);
or U8827 (N_8827,N_6808,N_6603);
nor U8828 (N_8828,N_5594,N_7062);
and U8829 (N_8829,N_6754,N_4476);
or U8830 (N_8830,N_7479,N_4610);
xor U8831 (N_8831,N_6819,N_7716);
xnor U8832 (N_8832,N_6291,N_5121);
and U8833 (N_8833,N_6926,N_6212);
nor U8834 (N_8834,N_5678,N_7385);
or U8835 (N_8835,N_5800,N_6116);
nor U8836 (N_8836,N_5079,N_6027);
and U8837 (N_8837,N_6310,N_7757);
and U8838 (N_8838,N_4852,N_5878);
nor U8839 (N_8839,N_6901,N_7737);
xor U8840 (N_8840,N_4314,N_4633);
or U8841 (N_8841,N_4971,N_7858);
nand U8842 (N_8842,N_5413,N_5546);
or U8843 (N_8843,N_5187,N_7466);
or U8844 (N_8844,N_5440,N_5345);
or U8845 (N_8845,N_6069,N_5050);
and U8846 (N_8846,N_4475,N_7417);
nor U8847 (N_8847,N_4431,N_7558);
nand U8848 (N_8848,N_7377,N_7715);
xor U8849 (N_8849,N_4085,N_4415);
and U8850 (N_8850,N_7194,N_5025);
nor U8851 (N_8851,N_4440,N_4983);
xnor U8852 (N_8852,N_5977,N_6395);
and U8853 (N_8853,N_4833,N_4839);
nor U8854 (N_8854,N_5864,N_7182);
xnor U8855 (N_8855,N_7401,N_7257);
or U8856 (N_8856,N_6251,N_6482);
or U8857 (N_8857,N_6902,N_4645);
nand U8858 (N_8858,N_7337,N_5014);
and U8859 (N_8859,N_7748,N_6617);
nor U8860 (N_8860,N_4723,N_7592);
nor U8861 (N_8861,N_5441,N_7578);
nand U8862 (N_8862,N_4965,N_7488);
nor U8863 (N_8863,N_7657,N_6832);
nor U8864 (N_8864,N_6535,N_6738);
nor U8865 (N_8865,N_6893,N_4864);
nor U8866 (N_8866,N_5206,N_4263);
xor U8867 (N_8867,N_6461,N_5027);
and U8868 (N_8868,N_5494,N_6378);
nand U8869 (N_8869,N_6743,N_4654);
xnor U8870 (N_8870,N_5848,N_7847);
or U8871 (N_8871,N_7161,N_7355);
nand U8872 (N_8872,N_4792,N_4191);
nor U8873 (N_8873,N_7070,N_5975);
xor U8874 (N_8874,N_6856,N_7713);
nand U8875 (N_8875,N_6855,N_4146);
nor U8876 (N_8876,N_6249,N_4363);
nor U8877 (N_8877,N_5128,N_4196);
nor U8878 (N_8878,N_5607,N_6068);
or U8879 (N_8879,N_7546,N_7522);
and U8880 (N_8880,N_6121,N_7034);
and U8881 (N_8881,N_6368,N_6912);
or U8882 (N_8882,N_6475,N_6404);
nor U8883 (N_8883,N_5248,N_5924);
and U8884 (N_8884,N_7251,N_6382);
or U8885 (N_8885,N_6558,N_4716);
or U8886 (N_8886,N_4023,N_4172);
and U8887 (N_8887,N_7364,N_4174);
and U8888 (N_8888,N_4750,N_5819);
nor U8889 (N_8889,N_4709,N_6618);
or U8890 (N_8890,N_5827,N_6425);
or U8891 (N_8891,N_4075,N_4214);
nand U8892 (N_8892,N_7195,N_5256);
and U8893 (N_8893,N_4078,N_6938);
nor U8894 (N_8894,N_4125,N_6503);
xnor U8895 (N_8895,N_7571,N_7414);
or U8896 (N_8896,N_7650,N_7762);
nor U8897 (N_8897,N_6550,N_6466);
nor U8898 (N_8898,N_7826,N_5168);
nand U8899 (N_8899,N_5364,N_4245);
and U8900 (N_8900,N_7032,N_6309);
xor U8901 (N_8901,N_5538,N_4585);
or U8902 (N_8902,N_5730,N_7943);
xnor U8903 (N_8903,N_4818,N_7206);
and U8904 (N_8904,N_6666,N_7321);
or U8905 (N_8905,N_6655,N_5579);
nand U8906 (N_8906,N_4339,N_4982);
nand U8907 (N_8907,N_7125,N_7374);
or U8908 (N_8908,N_5420,N_7242);
xnor U8909 (N_8909,N_7457,N_6281);
xor U8910 (N_8910,N_6423,N_5540);
and U8911 (N_8911,N_5252,N_7040);
nand U8912 (N_8912,N_6495,N_4855);
or U8913 (N_8913,N_5588,N_6467);
or U8914 (N_8914,N_5698,N_5618);
xnor U8915 (N_8915,N_4241,N_7236);
xor U8916 (N_8916,N_4478,N_7340);
nand U8917 (N_8917,N_4470,N_5711);
nor U8918 (N_8918,N_4905,N_5926);
nand U8919 (N_8919,N_6096,N_4650);
nand U8920 (N_8920,N_5638,N_6834);
xnor U8921 (N_8921,N_4036,N_6841);
nand U8922 (N_8922,N_6485,N_4002);
nand U8923 (N_8923,N_5667,N_4795);
and U8924 (N_8924,N_4148,N_6411);
and U8925 (N_8925,N_6615,N_7411);
nor U8926 (N_8926,N_6330,N_4380);
nor U8927 (N_8927,N_7093,N_6980);
xnor U8928 (N_8928,N_6348,N_5563);
nor U8929 (N_8929,N_7792,N_5891);
xnor U8930 (N_8930,N_5916,N_5531);
nand U8931 (N_8931,N_7568,N_6098);
xnor U8932 (N_8932,N_7767,N_6837);
and U8933 (N_8933,N_4710,N_7076);
nand U8934 (N_8934,N_6562,N_6526);
xnor U8935 (N_8935,N_6254,N_6725);
nor U8936 (N_8936,N_7094,N_7198);
xor U8937 (N_8937,N_6258,N_6144);
and U8938 (N_8938,N_6399,N_4734);
xor U8939 (N_8939,N_7524,N_4149);
and U8940 (N_8940,N_7039,N_6352);
and U8941 (N_8941,N_7848,N_6078);
and U8942 (N_8942,N_4823,N_5630);
nand U8943 (N_8943,N_4080,N_7615);
and U8944 (N_8944,N_5293,N_4891);
and U8945 (N_8945,N_7281,N_7168);
xnor U8946 (N_8946,N_4099,N_4422);
nor U8947 (N_8947,N_4254,N_6047);
xnor U8948 (N_8948,N_7490,N_7077);
nor U8949 (N_8949,N_4622,N_5290);
nor U8950 (N_8950,N_4407,N_6319);
xor U8951 (N_8951,N_4692,N_7699);
and U8952 (N_8952,N_7069,N_5091);
nor U8953 (N_8953,N_6004,N_5670);
nor U8954 (N_8954,N_4499,N_4485);
or U8955 (N_8955,N_5889,N_4465);
nor U8956 (N_8956,N_7726,N_7947);
or U8957 (N_8957,N_6172,N_5155);
xor U8958 (N_8958,N_4873,N_7322);
and U8959 (N_8959,N_4592,N_5489);
and U8960 (N_8960,N_6193,N_7827);
xnor U8961 (N_8961,N_5894,N_7292);
and U8962 (N_8962,N_4301,N_4140);
xor U8963 (N_8963,N_5224,N_7095);
xor U8964 (N_8964,N_7912,N_4020);
xor U8965 (N_8965,N_5459,N_5592);
nand U8966 (N_8966,N_6879,N_6396);
or U8967 (N_8967,N_6511,N_4318);
xnor U8968 (N_8968,N_4035,N_7005);
and U8969 (N_8969,N_7429,N_6106);
nor U8970 (N_8970,N_7008,N_4512);
or U8971 (N_8971,N_6228,N_6873);
xor U8972 (N_8972,N_6412,N_4807);
and U8973 (N_8973,N_4030,N_6632);
xor U8974 (N_8974,N_5209,N_4552);
xnor U8975 (N_8975,N_6968,N_4872);
nand U8976 (N_8976,N_4820,N_4367);
and U8977 (N_8977,N_4684,N_5396);
nor U8978 (N_8978,N_7729,N_7314);
nand U8979 (N_8979,N_6667,N_5852);
xor U8980 (N_8980,N_4095,N_5029);
nand U8981 (N_8981,N_6166,N_6608);
and U8982 (N_8982,N_6720,N_5539);
nor U8983 (N_8983,N_6161,N_7057);
nor U8984 (N_8984,N_7183,N_6470);
nand U8985 (N_8985,N_5193,N_7315);
nor U8986 (N_8986,N_6930,N_6598);
xor U8987 (N_8987,N_4705,N_6424);
and U8988 (N_8988,N_6721,N_6343);
xor U8989 (N_8989,N_6988,N_4608);
or U8990 (N_8990,N_6973,N_7110);
nand U8991 (N_8991,N_7204,N_7173);
or U8992 (N_8992,N_7103,N_6806);
nor U8993 (N_8993,N_7697,N_6835);
or U8994 (N_8994,N_6773,N_5062);
and U8995 (N_8995,N_7413,N_7841);
xnor U8996 (N_8996,N_4194,N_7796);
or U8997 (N_8997,N_6304,N_4832);
nor U8998 (N_8998,N_4724,N_6363);
xnor U8999 (N_8999,N_7885,N_7394);
or U9000 (N_9000,N_4473,N_7516);
nor U9001 (N_9001,N_7770,N_5250);
xnor U9002 (N_9002,N_4562,N_6668);
xor U9003 (N_9003,N_4681,N_7857);
nand U9004 (N_9004,N_6569,N_5968);
xor U9005 (N_9005,N_4659,N_4113);
or U9006 (N_9006,N_5362,N_4060);
nand U9007 (N_9007,N_6737,N_5586);
nor U9008 (N_9008,N_7189,N_5983);
xnor U9009 (N_9009,N_4917,N_6766);
and U9010 (N_9010,N_5903,N_4706);
nor U9011 (N_9011,N_5052,N_7358);
xnor U9012 (N_9012,N_5873,N_5401);
or U9013 (N_9013,N_6609,N_4584);
nand U9014 (N_9014,N_7460,N_7772);
nand U9015 (N_9015,N_5047,N_7165);
nand U9016 (N_9016,N_4616,N_6870);
or U9017 (N_9017,N_5509,N_6213);
or U9018 (N_9018,N_4515,N_5984);
xnor U9019 (N_9019,N_6136,N_7384);
xnor U9020 (N_9020,N_4454,N_6054);
or U9021 (N_9021,N_5033,N_6877);
nor U9022 (N_9022,N_4932,N_4304);
xnor U9023 (N_9023,N_5447,N_6852);
and U9024 (N_9024,N_6859,N_7760);
or U9025 (N_9025,N_6318,N_4647);
or U9026 (N_9026,N_5444,N_7936);
and U9027 (N_9027,N_7818,N_4460);
nand U9028 (N_9028,N_4939,N_6262);
nor U9029 (N_9029,N_7219,N_7518);
or U9030 (N_9030,N_6987,N_6394);
and U9031 (N_9031,N_7007,N_7643);
xor U9032 (N_9032,N_5676,N_7783);
nor U9033 (N_9033,N_6243,N_4761);
and U9034 (N_9034,N_4509,N_6914);
xnor U9035 (N_9035,N_6646,N_4248);
xor U9036 (N_9036,N_7909,N_6798);
and U9037 (N_9037,N_6559,N_7481);
and U9038 (N_9038,N_4010,N_4536);
nor U9039 (N_9039,N_6645,N_5446);
or U9040 (N_9040,N_5603,N_5057);
nor U9041 (N_9041,N_5971,N_6753);
xnor U9042 (N_9042,N_4255,N_7976);
and U9043 (N_9043,N_5473,N_7041);
xnor U9044 (N_9044,N_5392,N_4034);
nand U9045 (N_9045,N_6236,N_7664);
nor U9046 (N_9046,N_4530,N_4802);
and U9047 (N_9047,N_7310,N_7921);
nor U9048 (N_9048,N_5322,N_6874);
nor U9049 (N_9049,N_6498,N_5554);
xnor U9050 (N_9050,N_7906,N_4342);
and U9051 (N_9051,N_5288,N_7080);
nand U9052 (N_9052,N_7127,N_6443);
xor U9053 (N_9053,N_4348,N_6302);
or U9054 (N_9054,N_5766,N_4091);
nand U9055 (N_9055,N_7108,N_7451);
and U9056 (N_9056,N_7053,N_7356);
xor U9057 (N_9057,N_5945,N_7628);
or U9058 (N_9058,N_7752,N_4901);
xor U9059 (N_9059,N_4443,N_4264);
or U9060 (N_9060,N_7406,N_4686);
or U9061 (N_9061,N_4904,N_7489);
and U9062 (N_9062,N_4809,N_5492);
nor U9063 (N_9063,N_4921,N_7453);
or U9064 (N_9064,N_5504,N_6347);
xor U9065 (N_9065,N_5842,N_7740);
and U9066 (N_9066,N_4031,N_5194);
nand U9067 (N_9067,N_5108,N_6141);
xor U9068 (N_9068,N_6555,N_7601);
nor U9069 (N_9069,N_7192,N_7159);
xnor U9070 (N_9070,N_4779,N_6519);
or U9071 (N_9071,N_4050,N_4056);
or U9072 (N_9072,N_6789,N_4092);
nand U9073 (N_9073,N_6003,N_7138);
nand U9074 (N_9074,N_5907,N_6484);
nor U9075 (N_9075,N_4922,N_7075);
nor U9076 (N_9076,N_7029,N_5558);
and U9077 (N_9077,N_5267,N_6189);
or U9078 (N_9078,N_6446,N_6398);
or U9079 (N_9079,N_5475,N_4841);
and U9080 (N_9080,N_6315,N_6421);
or U9081 (N_9081,N_5214,N_5689);
or U9082 (N_9082,N_4093,N_6117);
or U9083 (N_9083,N_5790,N_4676);
xor U9084 (N_9084,N_5966,N_4830);
and U9085 (N_9085,N_4780,N_6851);
nor U9086 (N_9086,N_5748,N_6129);
and U9087 (N_9087,N_6145,N_4838);
nor U9088 (N_9088,N_4762,N_4071);
nand U9089 (N_9089,N_7392,N_5958);
and U9090 (N_9090,N_7870,N_5715);
and U9091 (N_9091,N_5859,N_6506);
nor U9092 (N_9092,N_4441,N_5529);
nor U9093 (N_9093,N_5464,N_6331);
xor U9094 (N_9094,N_4087,N_7970);
nor U9095 (N_9095,N_4572,N_6660);
nor U9096 (N_9096,N_4962,N_5685);
or U9097 (N_9097,N_6629,N_4305);
and U9098 (N_9098,N_4516,N_7285);
nand U9099 (N_9099,N_4799,N_4639);
nand U9100 (N_9100,N_6573,N_6583);
xor U9101 (N_9101,N_7896,N_7684);
nor U9102 (N_9102,N_4037,N_6534);
and U9103 (N_9103,N_7554,N_6444);
and U9104 (N_9104,N_5306,N_7399);
nor U9105 (N_9105,N_4941,N_4996);
and U9106 (N_9106,N_4945,N_5067);
nand U9107 (N_9107,N_5292,N_4351);
or U9108 (N_9108,N_4786,N_7698);
and U9109 (N_9109,N_4978,N_7325);
and U9110 (N_9110,N_7962,N_7940);
xnor U9111 (N_9111,N_6206,N_6784);
xor U9112 (N_9112,N_4463,N_4423);
nand U9113 (N_9113,N_5835,N_6082);
nor U9114 (N_9114,N_4883,N_6494);
or U9115 (N_9115,N_4677,N_6638);
nand U9116 (N_9116,N_7484,N_5264);
nor U9117 (N_9117,N_6622,N_6518);
and U9118 (N_9118,N_7682,N_5608);
nand U9119 (N_9119,N_5176,N_7809);
nor U9120 (N_9120,N_5016,N_6073);
nand U9121 (N_9121,N_6397,N_7751);
nor U9122 (N_9122,N_6350,N_5063);
or U9123 (N_9123,N_5722,N_7150);
nand U9124 (N_9124,N_4469,N_6025);
and U9125 (N_9125,N_5141,N_6179);
nor U9126 (N_9126,N_5598,N_6888);
xor U9127 (N_9127,N_6408,N_4298);
xor U9128 (N_9128,N_5437,N_7262);
xnor U9129 (N_9129,N_4898,N_4064);
xnor U9130 (N_9130,N_7815,N_5962);
xor U9131 (N_9131,N_6891,N_4118);
or U9132 (N_9132,N_5964,N_4167);
or U9133 (N_9133,N_4940,N_4661);
or U9134 (N_9134,N_4607,N_6177);
and U9135 (N_9135,N_7333,N_4667);
xnor U9136 (N_9136,N_6522,N_6038);
nand U9137 (N_9137,N_4384,N_5624);
nand U9138 (N_9138,N_5775,N_4319);
nor U9139 (N_9139,N_6241,N_6705);
and U9140 (N_9140,N_4492,N_5967);
nand U9141 (N_9141,N_6007,N_6878);
nand U9142 (N_9142,N_7063,N_7425);
and U9143 (N_9143,N_6547,N_4032);
or U9144 (N_9144,N_6866,N_5833);
and U9145 (N_9145,N_7519,N_6846);
and U9146 (N_9146,N_6907,N_6521);
nand U9147 (N_9147,N_4088,N_4708);
nand U9148 (N_9148,N_7446,N_4641);
and U9149 (N_9149,N_7838,N_5131);
or U9150 (N_9150,N_5243,N_5169);
xnor U9151 (N_9151,N_7927,N_6376);
nor U9152 (N_9152,N_4402,N_4185);
or U9153 (N_9153,N_5145,N_4875);
or U9154 (N_9154,N_5832,N_5450);
or U9155 (N_9155,N_6383,N_6611);
xnor U9156 (N_9156,N_6091,N_6542);
or U9157 (N_9157,N_6557,N_6365);
xnor U9158 (N_9158,N_4256,N_5107);
or U9159 (N_9159,N_6108,N_6934);
and U9160 (N_9160,N_6077,N_6017);
nand U9161 (N_9161,N_6553,N_5565);
nand U9162 (N_9162,N_5933,N_4117);
xor U9163 (N_9163,N_7999,N_5949);
and U9164 (N_9164,N_7427,N_5074);
nand U9165 (N_9165,N_4266,N_4991);
nand U9166 (N_9166,N_5823,N_4290);
and U9167 (N_9167,N_5519,N_5482);
xnor U9168 (N_9168,N_7197,N_6619);
and U9169 (N_9169,N_7541,N_6606);
nand U9170 (N_9170,N_7555,N_6923);
or U9171 (N_9171,N_5072,N_7902);
or U9172 (N_9172,N_4292,N_7806);
and U9173 (N_9173,N_5180,N_5543);
or U9174 (N_9174,N_4543,N_7248);
nor U9175 (N_9175,N_7820,N_6684);
nor U9176 (N_9176,N_5035,N_5386);
and U9177 (N_9177,N_5323,N_5856);
nand U9178 (N_9178,N_4179,N_6104);
and U9179 (N_9179,N_6238,N_5786);
nor U9180 (N_9180,N_4197,N_7619);
nand U9181 (N_9181,N_7038,N_6105);
nor U9182 (N_9182,N_7654,N_5031);
nor U9183 (N_9183,N_7627,N_7672);
nor U9184 (N_9184,N_4907,N_4445);
and U9185 (N_9185,N_4222,N_5866);
or U9186 (N_9186,N_4636,N_5227);
nor U9187 (N_9187,N_4210,N_7324);
xor U9188 (N_9188,N_6971,N_5655);
nor U9189 (N_9189,N_6472,N_7932);
nor U9190 (N_9190,N_6123,N_6321);
nor U9191 (N_9191,N_5491,N_7239);
nand U9192 (N_9192,N_7534,N_7742);
or U9193 (N_9193,N_5476,N_5122);
or U9194 (N_9194,N_7028,N_5625);
nor U9195 (N_9195,N_6055,N_5559);
nand U9196 (N_9196,N_4819,N_5524);
xnor U9197 (N_9197,N_6066,N_7595);
xnor U9198 (N_9198,N_6086,N_5534);
or U9199 (N_9199,N_4713,N_5350);
nand U9200 (N_9200,N_5201,N_4966);
or U9201 (N_9201,N_7553,N_7996);
nand U9202 (N_9202,N_5454,N_7431);
xnor U9203 (N_9203,N_4989,N_7268);
nand U9204 (N_9204,N_4084,N_7542);
or U9205 (N_9205,N_5303,N_5742);
nand U9206 (N_9206,N_4299,N_6328);
xor U9207 (N_9207,N_5908,N_6733);
xor U9208 (N_9208,N_5458,N_4369);
and U9209 (N_9209,N_5773,N_7718);
xor U9210 (N_9210,N_5541,N_6719);
nor U9211 (N_9211,N_6492,N_4291);
and U9212 (N_9212,N_6524,N_4374);
nor U9213 (N_9213,N_7968,N_7045);
and U9214 (N_9214,N_5771,N_4853);
nor U9215 (N_9215,N_7641,N_5192);
and U9216 (N_9216,N_7793,N_7423);
nor U9217 (N_9217,N_7383,N_4550);
and U9218 (N_9218,N_7696,N_7712);
or U9219 (N_9219,N_6048,N_4029);
and U9220 (N_9220,N_7911,N_6441);
xnor U9221 (N_9221,N_5759,N_6779);
xor U9222 (N_9222,N_4103,N_7240);
xor U9223 (N_9223,N_6202,N_5784);
or U9224 (N_9224,N_6781,N_5918);
and U9225 (N_9225,N_5704,N_7271);
nor U9226 (N_9226,N_4267,N_7033);
xor U9227 (N_9227,N_5955,N_4496);
nand U9228 (N_9228,N_4814,N_7840);
or U9229 (N_9229,N_4403,N_5404);
nand U9230 (N_9230,N_7311,N_7835);
xnor U9231 (N_9231,N_6685,N_5251);
nand U9232 (N_9232,N_6752,N_4574);
nor U9233 (N_9233,N_4956,N_4366);
or U9234 (N_9234,N_6184,N_7258);
or U9235 (N_9235,N_6239,N_6157);
nand U9236 (N_9236,N_7738,N_5405);
nand U9237 (N_9237,N_7759,N_6064);
nor U9238 (N_9238,N_5716,N_4911);
nand U9239 (N_9239,N_4963,N_7329);
nor U9240 (N_9240,N_5705,N_5532);
or U9241 (N_9241,N_5901,N_5680);
or U9242 (N_9242,N_7607,N_6195);
xor U9243 (N_9243,N_5073,N_6800);
or U9244 (N_9244,N_4866,N_7890);
nor U9245 (N_9245,N_6393,N_4021);
nand U9246 (N_9246,N_4089,N_4114);
and U9247 (N_9247,N_7465,N_7525);
or U9248 (N_9248,N_4323,N_6232);
or U9249 (N_9249,N_7112,N_4341);
or U9250 (N_9250,N_6018,N_7629);
xor U9251 (N_9251,N_5081,N_6777);
nor U9252 (N_9252,N_6079,N_7702);
nand U9253 (N_9253,N_6276,N_6153);
and U9254 (N_9254,N_4481,N_6256);
nor U9255 (N_9255,N_5418,N_4718);
xnor U9256 (N_9256,N_5234,N_6677);
nor U9257 (N_9257,N_5972,N_5217);
xor U9258 (N_9258,N_6334,N_5340);
nor U9259 (N_9259,N_4357,N_5080);
nor U9260 (N_9260,N_5344,N_6552);
xor U9261 (N_9261,N_6661,N_7449);
xnor U9262 (N_9262,N_5246,N_5154);
or U9263 (N_9263,N_7854,N_7721);
and U9264 (N_9264,N_4243,N_6389);
and U9265 (N_9265,N_6801,N_5787);
or U9266 (N_9266,N_6886,N_6210);
xnor U9267 (N_9267,N_7283,N_7814);
and U9268 (N_9268,N_6435,N_5331);
or U9269 (N_9269,N_6896,N_5466);
nor U9270 (N_9270,N_5872,N_4234);
nand U9271 (N_9271,N_7879,N_6786);
nand U9272 (N_9272,N_4226,N_5100);
xor U9273 (N_9273,N_5516,N_4609);
xnor U9274 (N_9274,N_5535,N_7946);
or U9275 (N_9275,N_7863,N_4224);
nor U9276 (N_9276,N_7224,N_6970);
nor U9277 (N_9277,N_6992,N_7966);
xor U9278 (N_9278,N_4655,N_7982);
nand U9279 (N_9279,N_7983,N_7477);
or U9280 (N_9280,N_5801,N_5316);
nand U9281 (N_9281,N_4731,N_5177);
nand U9282 (N_9282,N_7573,N_5026);
xor U9283 (N_9283,N_6357,N_7745);
xnor U9284 (N_9284,N_7786,N_7618);
or U9285 (N_9285,N_4360,N_4082);
and U9286 (N_9286,N_7245,N_5262);
nand U9287 (N_9287,N_4206,N_7981);
or U9288 (N_9288,N_5426,N_7590);
nand U9289 (N_9289,N_7975,N_5105);
and U9290 (N_9290,N_7548,N_5514);
nand U9291 (N_9291,N_7991,N_4081);
or U9292 (N_9292,N_5127,N_4143);
xor U9293 (N_9293,N_4951,N_4528);
nor U9294 (N_9294,N_7025,N_4312);
nor U9295 (N_9295,N_7907,N_6895);
and U9296 (N_9296,N_7533,N_4145);
xor U9297 (N_9297,N_4381,N_7849);
nor U9298 (N_9298,N_4295,N_4916);
nor U9299 (N_9299,N_6299,N_4270);
nand U9300 (N_9300,N_4504,N_5453);
and U9301 (N_9301,N_4618,N_6829);
or U9302 (N_9302,N_4349,N_6845);
or U9303 (N_9303,N_7566,N_5257);
and U9304 (N_9304,N_6487,N_7107);
nor U9305 (N_9305,N_5606,N_6433);
or U9306 (N_9306,N_5133,N_6169);
and U9307 (N_9307,N_5354,N_7690);
nand U9308 (N_9308,N_4914,N_6982);
nand U9309 (N_9309,N_6162,N_4307);
nor U9310 (N_9310,N_6876,N_6644);
xor U9311 (N_9311,N_6083,N_6650);
nor U9312 (N_9312,N_7583,N_7030);
nand U9313 (N_9313,N_5140,N_4579);
and U9314 (N_9314,N_6794,N_5407);
nor U9315 (N_9315,N_5556,N_7419);
xor U9316 (N_9316,N_4712,N_5566);
nand U9317 (N_9317,N_4745,N_6034);
or U9318 (N_9318,N_5960,N_4756);
and U9319 (N_9319,N_5120,N_4827);
xor U9320 (N_9320,N_4850,N_5591);
nor U9321 (N_9321,N_4665,N_7691);
xnor U9322 (N_9322,N_4788,N_5010);
xnor U9323 (N_9323,N_7398,N_4600);
nor U9324 (N_9324,N_6006,N_5285);
xnor U9325 (N_9325,N_6713,N_5351);
or U9326 (N_9326,N_6560,N_7585);
nand U9327 (N_9327,N_6037,N_5092);
nor U9328 (N_9328,N_7260,N_5024);
nor U9329 (N_9329,N_7366,N_4593);
nor U9330 (N_9330,N_4028,N_7930);
xnor U9331 (N_9331,N_6810,N_4211);
nand U9332 (N_9332,N_4811,N_4889);
nor U9333 (N_9333,N_4927,N_7067);
nand U9334 (N_9334,N_4371,N_4817);
and U9335 (N_9335,N_6990,N_6046);
xnor U9336 (N_9336,N_7513,N_7929);
nor U9337 (N_9337,N_5834,N_7919);
nand U9338 (N_9338,N_7415,N_5799);
or U9339 (N_9339,N_4163,N_4437);
or U9340 (N_9340,N_7717,N_5898);
and U9341 (N_9341,N_5008,N_7304);
nand U9342 (N_9342,N_5384,N_7780);
and U9343 (N_9343,N_4849,N_4967);
or U9344 (N_9344,N_5613,N_7126);
and U9345 (N_9345,N_7969,N_6049);
and U9346 (N_9346,N_4217,N_5982);
and U9347 (N_9347,N_6950,N_7343);
nand U9348 (N_9348,N_6491,N_6880);
xor U9349 (N_9349,N_5731,N_7247);
xnor U9350 (N_9350,N_6538,N_7536);
xnor U9351 (N_9351,N_6599,N_4682);
xnor U9352 (N_9352,N_4272,N_5892);
and U9353 (N_9353,N_7951,N_4632);
and U9354 (N_9354,N_6002,N_4387);
nand U9355 (N_9355,N_4069,N_7115);
or U9356 (N_9356,N_7121,N_6175);
nand U9357 (N_9357,N_6787,N_5278);
xor U9358 (N_9358,N_4759,N_7960);
and U9359 (N_9359,N_7471,N_5424);
nor U9360 (N_9360,N_7638,N_5287);
nor U9361 (N_9361,N_6134,N_7376);
xor U9362 (N_9362,N_7013,N_7084);
nand U9363 (N_9363,N_7552,N_5452);
and U9364 (N_9364,N_5549,N_4439);
xnor U9365 (N_9365,N_4671,N_4674);
nor U9366 (N_9366,N_5788,N_5513);
or U9367 (N_9367,N_4240,N_7359);
xor U9368 (N_9368,N_6940,N_5729);
nand U9369 (N_9369,N_7439,N_6386);
nor U9370 (N_9370,N_4949,N_5576);
and U9371 (N_9371,N_7528,N_4913);
and U9372 (N_9372,N_7205,N_5281);
or U9373 (N_9373,N_4538,N_5807);
nand U9374 (N_9374,N_4627,N_7576);
nor U9375 (N_9375,N_7344,N_6469);
xnor U9376 (N_9376,N_7083,N_4482);
or U9377 (N_9377,N_5488,N_7725);
and U9378 (N_9378,N_5537,N_5822);
nor U9379 (N_9379,N_4456,N_6225);
nand U9380 (N_9380,N_7666,N_7117);
nor U9381 (N_9381,N_5428,N_6160);
nor U9382 (N_9382,N_7430,N_4753);
or U9383 (N_9383,N_4505,N_6502);
nor U9384 (N_9384,N_5883,N_6780);
or U9385 (N_9385,N_5266,N_6683);
and U9386 (N_9386,N_6474,N_5230);
nor U9387 (N_9387,N_7681,N_5060);
nand U9388 (N_9388,N_5319,N_4703);
or U9389 (N_9389,N_7754,N_7880);
nand U9390 (N_9390,N_6222,N_7584);
or U9391 (N_9391,N_7891,N_6124);
nand U9392 (N_9392,N_7570,N_5434);
and U9393 (N_9393,N_7208,N_6742);
or U9394 (N_9394,N_5953,N_5236);
and U9395 (N_9395,N_4771,N_4426);
nand U9396 (N_9396,N_6530,N_6501);
nor U9397 (N_9397,N_5104,N_4013);
nor U9398 (N_9398,N_5415,N_5703);
or U9399 (N_9399,N_7942,N_5781);
or U9400 (N_9400,N_6283,N_4246);
nand U9401 (N_9401,N_7497,N_5470);
nor U9402 (N_9402,N_5664,N_5397);
and U9403 (N_9403,N_5976,N_5393);
nand U9404 (N_9404,N_5840,N_5779);
nand U9405 (N_9405,N_4288,N_6298);
nand U9406 (N_9406,N_6110,N_6113);
or U9407 (N_9407,N_4936,N_7512);
xnor U9408 (N_9408,N_5279,N_6605);
nand U9409 (N_9409,N_7381,N_4977);
xor U9410 (N_9410,N_6929,N_4881);
nand U9411 (N_9411,N_6529,N_6727);
xor U9412 (N_9412,N_6245,N_6351);
nand U9413 (N_9413,N_7603,N_6697);
or U9414 (N_9414,N_7395,N_7747);
xnor U9415 (N_9415,N_4992,N_6986);
xor U9416 (N_9416,N_5002,N_4417);
xnor U9417 (N_9417,N_4017,N_4001);
xor U9418 (N_9418,N_5855,N_6875);
and U9419 (N_9419,N_6422,N_4404);
nor U9420 (N_9420,N_4581,N_7864);
or U9421 (N_9421,N_6458,N_7213);
and U9422 (N_9422,N_7795,N_5164);
or U9423 (N_9423,N_4954,N_6871);
xnor U9424 (N_9424,N_5158,N_5753);
or U9425 (N_9425,N_5330,N_6237);
nor U9426 (N_9426,N_4040,N_7346);
nor U9427 (N_9427,N_7875,N_5905);
xor U9428 (N_9428,N_6406,N_4776);
or U9429 (N_9429,N_5652,N_4895);
or U9430 (N_9430,N_7350,N_5762);
nor U9431 (N_9431,N_4806,N_6103);
xor U9432 (N_9432,N_5498,N_5260);
nor U9433 (N_9433,N_5510,N_7483);
or U9434 (N_9434,N_7839,N_7035);
nor U9435 (N_9435,N_7261,N_6279);
or U9436 (N_9436,N_4625,N_4128);
xor U9437 (N_9437,N_5761,N_7332);
xnor U9438 (N_9438,N_6311,N_7347);
or U9439 (N_9439,N_5071,N_5622);
nor U9440 (N_9440,N_7587,N_5377);
and U9441 (N_9441,N_6663,N_6209);
xor U9442 (N_9442,N_7442,N_7577);
and U9443 (N_9443,N_4231,N_4797);
nor U9444 (N_9444,N_6185,N_4189);
nor U9445 (N_9445,N_7952,N_5111);
nor U9446 (N_9446,N_4778,N_5412);
and U9447 (N_9447,N_7505,N_4928);
and U9448 (N_9448,N_7370,N_5612);
nand U9449 (N_9449,N_4138,N_4136);
xor U9450 (N_9450,N_7985,N_7794);
or U9451 (N_9451,N_6954,N_6993);
and U9452 (N_9452,N_5641,N_5782);
and U9453 (N_9453,N_7147,N_4340);
or U9454 (N_9454,N_6401,N_4483);
nor U9455 (N_9455,N_5536,N_5055);
or U9456 (N_9456,N_6451,N_6749);
nor U9457 (N_9457,N_4527,N_7275);
nor U9458 (N_9458,N_4506,N_7175);
nor U9459 (N_9459,N_5750,N_6114);
nand U9460 (N_9460,N_6946,N_4193);
and U9461 (N_9461,N_5219,N_4594);
or U9462 (N_9462,N_4589,N_5525);
xor U9463 (N_9463,N_4737,N_5520);
or U9464 (N_9464,N_7263,N_5619);
xor U9465 (N_9465,N_5034,N_6574);
or U9466 (N_9466,N_5644,N_5783);
or U9467 (N_9467,N_5646,N_7928);
nand U9468 (N_9468,N_7527,N_7313);
xnor U9469 (N_9469,N_4580,N_4933);
nor U9470 (N_9470,N_7631,N_5001);
and U9471 (N_9471,N_6438,N_4620);
xor U9472 (N_9472,N_4336,N_4777);
and U9473 (N_9473,N_5297,N_7551);
or U9474 (N_9474,N_5208,N_5739);
xor U9475 (N_9475,N_6308,N_7207);
nor U9476 (N_9476,N_6932,N_4155);
and U9477 (N_9477,N_7104,N_6576);
nand U9478 (N_9478,N_6711,N_6610);
nor U9479 (N_9479,N_6728,N_6481);
or U9480 (N_9480,N_4359,N_7674);
nand U9481 (N_9481,N_5089,N_4586);
xnor U9482 (N_9482,N_6342,N_7837);
nor U9483 (N_9483,N_4278,N_5069);
nor U9484 (N_9484,N_4548,N_6785);
and U9485 (N_9485,N_5274,N_6757);
and U9486 (N_9486,N_7468,N_7297);
or U9487 (N_9487,N_7362,N_4495);
and U9488 (N_9488,N_5496,N_6403);
or U9489 (N_9489,N_5526,N_5749);
or U9490 (N_9490,N_7967,N_4503);
nand U9491 (N_9491,N_5569,N_5147);
and U9492 (N_9492,N_7100,N_7331);
nand U9493 (N_9493,N_6204,N_6775);
nor U9494 (N_9494,N_7341,N_4090);
and U9495 (N_9495,N_5406,N_4836);
or U9496 (N_9496,N_7494,N_4856);
nor U9497 (N_9497,N_5315,N_6333);
nand U9498 (N_9498,N_5952,N_4327);
nand U9499 (N_9499,N_6883,N_6885);
nand U9500 (N_9500,N_4735,N_7531);
nand U9501 (N_9501,N_6196,N_5268);
nand U9502 (N_9502,N_4906,N_5461);
nand U9503 (N_9503,N_6143,N_4018);
nand U9504 (N_9504,N_5838,N_4617);
or U9505 (N_9505,N_5408,N_6231);
nand U9506 (N_9506,N_7291,N_4072);
nor U9507 (N_9507,N_6266,N_6415);
and U9508 (N_9508,N_7019,N_5615);
xnor U9509 (N_9509,N_5378,N_7146);
and U9510 (N_9510,N_6131,N_4987);
nand U9511 (N_9511,N_7272,N_7305);
nor U9512 (N_9512,N_4997,N_6872);
and U9513 (N_9513,N_5336,N_5445);
and U9514 (N_9514,N_5098,N_4382);
xnor U9515 (N_9515,N_6076,N_7074);
and U9516 (N_9516,N_7143,N_5887);
xnor U9517 (N_9517,N_4732,N_6120);
nand U9518 (N_9518,N_4791,N_4715);
nand U9519 (N_9519,N_4025,N_4162);
nand U9520 (N_9520,N_6958,N_6591);
and U9521 (N_9521,N_6336,N_4477);
and U9522 (N_9522,N_7874,N_6979);
nand U9523 (N_9523,N_4595,N_4199);
or U9524 (N_9524,N_7821,N_5425);
and U9525 (N_9525,N_7861,N_4648);
and U9526 (N_9526,N_7944,N_4660);
and U9527 (N_9527,N_7475,N_4857);
xnor U9528 (N_9528,N_5938,N_7101);
xnor U9529 (N_9529,N_7855,N_4073);
nor U9530 (N_9530,N_6755,N_5011);
or U9531 (N_9531,N_4322,N_5150);
or U9532 (N_9532,N_6180,N_4310);
and U9533 (N_9533,N_4825,N_4362);
xnor U9534 (N_9534,N_7079,N_5332);
or U9535 (N_9535,N_7472,N_7086);
or U9536 (N_9536,N_5672,N_4104);
and U9537 (N_9537,N_7728,N_5919);
nand U9538 (N_9538,N_5244,N_4947);
nor U9539 (N_9539,N_4325,N_5253);
xor U9540 (N_9540,N_4537,N_7844);
nand U9541 (N_9541,N_6273,N_4083);
or U9542 (N_9542,N_4329,N_4929);
nor U9543 (N_9543,N_4926,N_7633);
nor U9544 (N_9544,N_7646,N_7301);
or U9545 (N_9545,N_7330,N_5809);
and U9546 (N_9546,N_7710,N_4346);
or U9547 (N_9547,N_4848,N_4131);
nand U9548 (N_9548,N_4438,N_5713);
nand U9549 (N_9549,N_4253,N_7948);
or U9550 (N_9550,N_5042,N_7956);
nor U9551 (N_9551,N_5116,N_5956);
xnor U9552 (N_9552,N_6374,N_4120);
and U9553 (N_9553,N_5036,N_7089);
or U9554 (N_9554,N_4190,N_4115);
nor U9555 (N_9555,N_5156,N_4535);
or U9556 (N_9556,N_5912,N_6589);
xnor U9557 (N_9557,N_7151,N_4566);
nor U9558 (N_9558,N_6217,N_4520);
or U9559 (N_9559,N_5259,N_5355);
nor U9560 (N_9560,N_7303,N_4378);
or U9561 (N_9561,N_5044,N_4345);
xor U9562 (N_9562,N_7648,N_4994);
nand U9563 (N_9563,N_7537,N_5442);
xor U9564 (N_9564,N_4754,N_5271);
xnor U9565 (N_9565,N_7216,N_6690);
nand U9566 (N_9566,N_4435,N_4815);
xnor U9567 (N_9567,N_6818,N_5542);
nor U9568 (N_9568,N_4511,N_7306);
nand U9569 (N_9569,N_6250,N_7157);
xnor U9570 (N_9570,N_6455,N_4970);
nor U9571 (N_9571,N_4265,N_4859);
and U9572 (N_9572,N_7118,N_4281);
xnor U9573 (N_9573,N_5925,N_6994);
or U9574 (N_9574,N_4286,N_6453);
nor U9575 (N_9575,N_5841,N_7597);
nor U9576 (N_9576,N_4394,N_4884);
and U9577 (N_9577,N_4079,N_4701);
or U9578 (N_9578,N_6014,N_5103);
or U9579 (N_9579,N_7011,N_4549);
nand U9580 (N_9580,N_4877,N_6596);
xnor U9581 (N_9581,N_6949,N_6154);
nand U9582 (N_9582,N_7564,N_7799);
or U9583 (N_9583,N_6523,N_5793);
nor U9584 (N_9584,N_7000,N_5269);
nand U9585 (N_9585,N_7269,N_7015);
nor U9586 (N_9586,N_7569,N_4044);
nor U9587 (N_9587,N_4459,N_4063);
xor U9588 (N_9588,N_7971,N_7801);
nand U9589 (N_9589,N_7357,N_4919);
nor U9590 (N_9590,N_6656,N_7905);
or U9591 (N_9591,N_5430,N_7652);
nand U9592 (N_9592,N_4912,N_5200);
or U9593 (N_9593,N_7137,N_7608);
nor U9594 (N_9594,N_5614,N_6527);
or U9595 (N_9595,N_6051,N_5245);
nor U9596 (N_9596,N_5300,N_7787);
and U9597 (N_9597,N_4235,N_4816);
nor U9598 (N_9598,N_6151,N_7001);
xnor U9599 (N_9599,N_6140,N_4605);
xnor U9600 (N_9600,N_6700,N_6570);
nor U9601 (N_9601,N_6687,N_4411);
and U9602 (N_9602,N_7995,N_7798);
and U9603 (N_9603,N_5109,N_5314);
nand U9604 (N_9604,N_6981,N_6323);
nor U9605 (N_9605,N_4249,N_6257);
xor U9606 (N_9606,N_4698,N_5829);
nor U9607 (N_9607,N_4995,N_6335);
nand U9608 (N_9608,N_5006,N_5605);
nand U9609 (N_9609,N_4935,N_6377);
xnor U9610 (N_9610,N_5085,N_6278);
or U9611 (N_9611,N_5410,N_7099);
and U9612 (N_9612,N_5449,N_6817);
nand U9613 (N_9613,N_7973,N_6028);
or U9614 (N_9614,N_5126,N_7544);
or U9615 (N_9615,N_7776,N_4868);
nand U9616 (N_9616,N_7163,N_5709);
nand U9617 (N_9617,N_4414,N_5198);
nand U9618 (N_9618,N_5902,N_5421);
and U9619 (N_9619,N_7132,N_6927);
or U9620 (N_9620,N_5202,N_5553);
and U9621 (N_9621,N_6525,N_6807);
nand U9622 (N_9622,N_5225,N_5567);
nor U9623 (N_9623,N_4068,N_5339);
nor U9624 (N_9624,N_7530,N_5123);
and U9625 (N_9625,N_6731,N_5574);
xnor U9626 (N_9626,N_7027,N_6019);
and U9627 (N_9627,N_7803,N_6493);
or U9628 (N_9628,N_4133,N_7997);
and U9629 (N_9629,N_5417,N_4690);
or U9630 (N_9630,N_6391,N_7775);
and U9631 (N_9631,N_4108,N_6778);
nand U9632 (N_9632,N_6387,N_4879);
xnor U9633 (N_9633,N_6985,N_4300);
nand U9634 (N_9634,N_7049,N_4541);
or U9635 (N_9635,N_6678,N_6905);
nand U9636 (N_9636,N_5213,N_5159);
or U9637 (N_9637,N_6338,N_7660);
xor U9638 (N_9638,N_4931,N_4843);
xnor U9639 (N_9639,N_7705,N_7805);
nor U9640 (N_9640,N_5394,N_6381);
xnor U9641 (N_9641,N_5942,N_4656);
xnor U9642 (N_9642,N_5037,N_4280);
or U9643 (N_9643,N_5657,N_6107);
and U9644 (N_9644,N_5726,N_4930);
xnor U9645 (N_9645,N_5358,N_4227);
and U9646 (N_9646,N_4400,N_6497);
nor U9647 (N_9647,N_7421,N_7925);
nand U9648 (N_9648,N_6101,N_6670);
nor U9649 (N_9649,N_4086,N_6616);
and U9650 (N_9650,N_5083,N_6059);
nand U9651 (N_9651,N_6545,N_7914);
xnor U9652 (N_9652,N_7899,N_6961);
nand U9653 (N_9653,N_6295,N_4946);
or U9654 (N_9654,N_4783,N_5899);
and U9655 (N_9655,N_5343,N_4533);
and U9656 (N_9656,N_7876,N_6536);
nand U9657 (N_9657,N_4395,N_5961);
nand U9658 (N_9658,N_4169,N_5708);
xnor U9659 (N_9659,N_5500,N_6600);
nand U9660 (N_9660,N_4635,N_6471);
or U9661 (N_9661,N_7230,N_4726);
and U9662 (N_9662,N_6205,N_5439);
nand U9663 (N_9663,N_4039,N_4244);
or U9664 (N_9664,N_4744,N_6520);
or U9665 (N_9665,N_5341,N_4181);
xnor U9666 (N_9666,N_4693,N_6830);
xnor U9667 (N_9667,N_4467,N_7064);
xnor U9668 (N_9668,N_6122,N_5320);
or U9669 (N_9669,N_5806,N_6268);
and U9670 (N_9670,N_6267,N_4376);
and U9671 (N_9671,N_6792,N_7621);
xnor U9672 (N_9672,N_6050,N_5184);
and U9673 (N_9673,N_5599,N_5692);
and U9674 (N_9674,N_4882,N_5530);
xnor U9675 (N_9675,N_4634,N_7692);
xnor U9676 (N_9676,N_4624,N_5570);
or U9677 (N_9677,N_7252,N_5455);
or U9678 (N_9678,N_7688,N_5959);
nor U9679 (N_9679,N_7360,N_7006);
and U9680 (N_9680,N_5115,N_6300);
nand U9681 (N_9681,N_6805,N_5719);
nor U9682 (N_9682,N_7243,N_7860);
nand U9683 (N_9683,N_7514,N_4033);
nand U9684 (N_9684,N_5097,N_7744);
nand U9685 (N_9685,N_5132,N_5660);
nand U9686 (N_9686,N_7319,N_5152);
nor U9687 (N_9687,N_5051,N_7581);
and U9688 (N_9688,N_6745,N_7046);
nand U9689 (N_9689,N_4361,N_6868);
or U9690 (N_9690,N_4782,N_4335);
nor U9691 (N_9691,N_6952,N_5138);
and U9692 (N_9692,N_7832,N_7845);
xnor U9693 (N_9693,N_4311,N_6933);
and U9694 (N_9694,N_7978,N_7526);
or U9695 (N_9695,N_7964,N_7456);
nor U9696 (N_9696,N_7418,N_4334);
nor U9697 (N_9697,N_7862,N_7704);
or U9698 (N_9698,N_7308,N_5658);
nor U9699 (N_9699,N_6430,N_4186);
nor U9700 (N_9700,N_4861,N_5981);
nor U9701 (N_9701,N_7829,N_6674);
and U9702 (N_9702,N_6898,N_5237);
and U9703 (N_9703,N_6380,N_4446);
nand U9704 (N_9704,N_4601,N_7298);
xor U9705 (N_9705,N_4365,N_4421);
or U9706 (N_9706,N_6827,N_6613);
nor U9707 (N_9707,N_5813,N_5747);
or U9708 (N_9708,N_5400,N_5610);
nor U9709 (N_9709,N_4171,N_6739);
xnor U9710 (N_9710,N_5935,N_5710);
xnor U9711 (N_9711,N_7296,N_7714);
and U9712 (N_9712,N_6735,N_6457);
xnor U9713 (N_9713,N_7915,N_4188);
xnor U9714 (N_9714,N_4583,N_5380);
or U9715 (N_9715,N_6316,N_4147);
xor U9716 (N_9716,N_6998,N_4158);
and U9717 (N_9717,N_4126,N_6289);
or U9718 (N_9718,N_6580,N_6203);
or U9719 (N_9719,N_4408,N_5733);
nand U9720 (N_9720,N_6802,N_7042);
nand U9721 (N_9721,N_5706,N_7750);
xor U9722 (N_9722,N_5282,N_7868);
nor U9723 (N_9723,N_4867,N_7895);
nor U9724 (N_9724,N_5562,N_4309);
nor U9725 (N_9725,N_4765,N_4722);
xnor U9726 (N_9726,N_6999,N_4598);
nand U9727 (N_9727,N_6825,N_5205);
nor U9728 (N_9728,N_5479,N_7153);
and U9729 (N_9729,N_5754,N_4047);
and U9730 (N_9730,N_6142,N_7802);
nand U9731 (N_9731,N_7656,N_4170);
nor U9732 (N_9732,N_7473,N_5218);
nand U9733 (N_9733,N_7560,N_6463);
nor U9734 (N_9734,N_4385,N_6199);
xnor U9735 (N_9735,N_5796,N_4142);
xor U9736 (N_9736,N_7010,N_7653);
nand U9737 (N_9737,N_7485,N_5328);
and U9738 (N_9738,N_6768,N_6063);
xor U9739 (N_9739,N_7825,N_7972);
nand U9740 (N_9740,N_4563,N_6783);
and U9741 (N_9741,N_5792,N_7722);
nand U9742 (N_9742,N_7102,N_7871);
nor U9743 (N_9743,N_7259,N_6664);
and U9744 (N_9744,N_5811,N_4392);
or U9745 (N_9745,N_5471,N_6863);
or U9746 (N_9746,N_6708,N_7491);
or U9747 (N_9747,N_4150,N_7807);
nand U9748 (N_9748,N_7635,N_6479);
nand U9749 (N_9749,N_7963,N_7781);
nor U9750 (N_9750,N_4714,N_6427);
and U9751 (N_9751,N_5065,N_7318);
xnor U9752 (N_9752,N_6696,N_4353);
nand U9753 (N_9753,N_5135,N_5951);
xor U9754 (N_9754,N_5240,N_6009);
nor U9755 (N_9755,N_7758,N_4569);
or U9756 (N_9756,N_4793,N_7889);
nand U9757 (N_9757,N_7958,N_6448);
nand U9758 (N_9758,N_7066,N_4122);
xor U9759 (N_9759,N_5061,N_6772);
nand U9760 (N_9760,N_7092,N_7155);
nand U9761 (N_9761,N_5882,N_6746);
xnor U9762 (N_9762,N_6915,N_6436);
nor U9763 (N_9763,N_5850,N_5474);
nand U9764 (N_9764,N_4430,N_7096);
and U9765 (N_9765,N_7549,N_7883);
and U9766 (N_9766,N_7090,N_6163);
and U9767 (N_9767,N_6821,N_7133);
and U9768 (N_9768,N_4057,N_5374);
xnor U9769 (N_9769,N_6460,N_6349);
nor U9770 (N_9770,N_5880,N_7788);
nand U9771 (N_9771,N_5136,N_6681);
nand U9772 (N_9772,N_4957,N_6763);
or U9773 (N_9773,N_4258,N_5359);
nor U9774 (N_9774,N_4729,N_5824);
and U9775 (N_9775,N_6432,N_6362);
xor U9776 (N_9776,N_4048,N_5232);
nand U9777 (N_9777,N_4733,N_5212);
xor U9778 (N_9778,N_6152,N_4858);
and U9779 (N_9779,N_7136,N_5987);
xor U9780 (N_9780,N_6890,N_7186);
nor U9781 (N_9781,N_7917,N_6762);
and U9782 (N_9782,N_5235,N_4576);
xor U9783 (N_9783,N_4587,N_7336);
nand U9784 (N_9784,N_5896,N_5056);
nand U9785 (N_9785,N_7882,N_7755);
or U9786 (N_9786,N_6680,N_7480);
nor U9787 (N_9787,N_4203,N_5167);
and U9788 (N_9788,N_5640,N_7594);
xor U9789 (N_9789,N_4747,N_5096);
xnor U9790 (N_9790,N_6551,N_5276);
or U9791 (N_9791,N_7843,N_6554);
and U9792 (N_9792,N_5411,N_4679);
xnor U9793 (N_9793,N_5515,N_6320);
nor U9794 (N_9794,N_4999,N_6095);
nor U9795 (N_9795,N_4663,N_6174);
and U9796 (N_9796,N_6010,N_7887);
or U9797 (N_9797,N_7856,N_6581);
nor U9798 (N_9798,N_6671,N_5687);
nand U9799 (N_9799,N_4787,N_7353);
xnor U9800 (N_9800,N_5755,N_5564);
or U9801 (N_9801,N_6995,N_4041);
xnor U9802 (N_9802,N_7176,N_7351);
xor U9803 (N_9803,N_5000,N_6125);
or U9804 (N_9804,N_6862,N_5769);
nor U9805 (N_9805,N_7047,N_7604);
and U9806 (N_9806,N_7065,N_4651);
nand U9807 (N_9807,N_5040,N_7177);
or U9808 (N_9808,N_4202,N_5403);
and U9809 (N_9809,N_4887,N_6675);
or U9810 (N_9810,N_7299,N_6011);
xnor U9811 (N_9811,N_4352,N_7166);
nor U9812 (N_9812,N_6584,N_7131);
and U9813 (N_9813,N_5068,N_5617);
and U9814 (N_9814,N_6026,N_4388);
xor U9815 (N_9815,N_6452,N_7617);
xnor U9816 (N_9816,N_7201,N_4615);
or U9817 (N_9817,N_5478,N_4173);
nand U9818 (N_9818,N_5808,N_7605);
nor U9819 (N_9819,N_7238,N_6682);
nor U9820 (N_9820,N_7707,N_6496);
xnor U9821 (N_9821,N_5810,N_5139);
nor U9822 (N_9822,N_5522,N_6540);
nand U9823 (N_9823,N_6842,N_4098);
xor U9824 (N_9824,N_7884,N_6070);
nor U9825 (N_9825,N_7746,N_7613);
nor U9826 (N_9826,N_5490,N_4834);
or U9827 (N_9827,N_6253,N_5814);
nand U9828 (N_9828,N_5505,N_6370);
nor U9829 (N_9829,N_7129,N_5102);
and U9830 (N_9830,N_6917,N_6074);
nor U9831 (N_9831,N_7424,N_6983);
nor U9832 (N_9832,N_5911,N_7145);
or U9833 (N_9833,N_4397,N_6282);
and U9834 (N_9834,N_5718,N_6707);
xnor U9835 (N_9835,N_7388,N_6305);
nand U9836 (N_9836,N_6340,N_6796);
or U9837 (N_9837,N_7054,N_4604);
nor U9838 (N_9838,N_5357,N_7708);
nand U9839 (N_9839,N_4406,N_4251);
nand U9840 (N_9840,N_4338,N_7434);
nand U9841 (N_9841,N_6248,N_7405);
xnor U9842 (N_9842,N_6429,N_5764);
nor U9843 (N_9843,N_5974,N_4180);
nor U9844 (N_9844,N_7901,N_5263);
and U9845 (N_9845,N_7180,N_5860);
or U9846 (N_9846,N_4842,N_6922);
and U9847 (N_9847,N_7939,N_7059);
nand U9848 (N_9848,N_6831,N_4004);
and U9849 (N_9849,N_7458,N_4386);
nor U9850 (N_9850,N_6486,N_4597);
xor U9851 (N_9851,N_7517,N_7085);
and U9852 (N_9852,N_6426,N_7048);
and U9853 (N_9853,N_7002,N_4011);
or U9854 (N_9854,N_7142,N_6612);
nor U9855 (N_9855,N_4796,N_7470);
xor U9856 (N_9856,N_6673,N_5595);
or U9857 (N_9857,N_5134,N_6402);
nand U9858 (N_9858,N_7302,N_5369);
nand U9859 (N_9859,N_6265,N_4077);
nand U9860 (N_9860,N_7669,N_7686);
or U9861 (N_9861,N_4985,N_7210);
or U9862 (N_9862,N_5803,N_4183);
nor U9863 (N_9863,N_5965,N_7819);
nor U9864 (N_9864,N_7766,N_6234);
xnor U9865 (N_9865,N_4560,N_6065);
nor U9866 (N_9866,N_6858,N_7731);
nor U9867 (N_9867,N_5129,N_4259);
nor U9868 (N_9868,N_5283,N_6702);
or U9869 (N_9869,N_6732,N_6060);
nand U9870 (N_9870,N_4521,N_5991);
nor U9871 (N_9871,N_5231,N_6869);
nand U9872 (N_9872,N_7317,N_7023);
nand U9873 (N_9873,N_7119,N_6188);
xnor U9874 (N_9874,N_7557,N_4344);
and U9875 (N_9875,N_5291,N_4442);
xnor U9876 (N_9876,N_7235,N_6747);
nand U9877 (N_9877,N_4497,N_6652);
or U9878 (N_9878,N_7817,N_6005);
and U9879 (N_9879,N_4109,N_4773);
nor U9880 (N_9880,N_6329,N_4640);
nand U9881 (N_9881,N_6916,N_6039);
and U9882 (N_9882,N_7520,N_6977);
or U9883 (N_9883,N_5497,N_6741);
nand U9884 (N_9884,N_6216,N_7892);
or U9885 (N_9885,N_7753,N_4302);
or U9886 (N_9886,N_5207,N_4269);
xnor U9887 (N_9887,N_6062,N_7218);
and U9888 (N_9888,N_6499,N_7276);
or U9889 (N_9889,N_4691,N_7492);
or U9890 (N_9890,N_7777,N_5653);
xor U9891 (N_9891,N_7379,N_4829);
nand U9892 (N_9892,N_5604,N_5649);
and U9893 (N_9893,N_6130,N_7474);
and U9894 (N_9894,N_4588,N_4420);
xor U9895 (N_9895,N_5637,N_5635);
or U9896 (N_9896,N_6000,N_5086);
or U9897 (N_9897,N_7232,N_7916);
nand U9898 (N_9898,N_6639,N_6942);
nor U9899 (N_9899,N_7435,N_5816);
or U9900 (N_9900,N_6201,N_4130);
xor U9901 (N_9901,N_4573,N_6931);
nor U9902 (N_9902,N_4794,N_6579);
nand U9903 (N_9903,N_6220,N_5015);
xor U9904 (N_9904,N_5118,N_7368);
nor U9905 (N_9905,N_7955,N_4491);
nand U9906 (N_9906,N_6053,N_7222);
xnor U9907 (N_9907,N_7800,N_7286);
or U9908 (N_9908,N_5021,N_5457);
nor U9909 (N_9909,N_5211,N_6833);
xnor U9910 (N_9910,N_4121,N_6976);
and U9911 (N_9911,N_7058,N_4611);
xnor U9912 (N_9912,N_5348,N_5684);
and U9913 (N_9913,N_4436,N_7675);
and U9914 (N_9914,N_6750,N_5070);
or U9915 (N_9915,N_7846,N_7510);
nand U9916 (N_9916,N_6575,N_7280);
nor U9917 (N_9917,N_7167,N_6400);
or U9918 (N_9918,N_7382,N_7723);
nand U9919 (N_9919,N_7908,N_5093);
nor U9920 (N_9920,N_4694,N_6008);
nor U9921 (N_9921,N_6084,N_7393);
xor U9922 (N_9922,N_4229,N_7642);
nor U9923 (N_9923,N_6449,N_6918);
nand U9924 (N_9924,N_5427,N_5146);
nand U9925 (N_9925,N_7779,N_7574);
nor U9926 (N_9926,N_6301,N_5151);
nand U9927 (N_9927,N_6718,N_4250);
xnor U9928 (N_9928,N_7367,N_6714);
nor U9929 (N_9929,N_7998,N_6759);
nor U9930 (N_9930,N_4379,N_7444);
xnor U9931 (N_9931,N_4490,N_5740);
nor U9932 (N_9932,N_6943,N_4000);
and U9933 (N_9933,N_6413,N_5183);
nand U9934 (N_9934,N_7284,N_5064);
xnor U9935 (N_9935,N_6686,N_5639);
xor U9936 (N_9936,N_6910,N_5552);
nor U9937 (N_9937,N_6198,N_5289);
xnor U9938 (N_9938,N_7436,N_6272);
nor U9939 (N_9939,N_6921,N_5683);
nand U9940 (N_9940,N_7824,N_4007);
or U9941 (N_9941,N_4016,N_5366);
nand U9942 (N_9942,N_6500,N_7897);
and U9943 (N_9943,N_5160,N_5696);
or U9944 (N_9944,N_4775,N_6736);
nand U9945 (N_9945,N_5258,N_6769);
or U9946 (N_9946,N_7508,N_7797);
nand U9947 (N_9947,N_4107,N_4652);
nand U9948 (N_9948,N_7923,N_5005);
and U9949 (N_9949,N_6384,N_6375);
or U9950 (N_9950,N_6208,N_6653);
nand U9951 (N_9951,N_5785,N_5815);
nor U9952 (N_9952,N_6490,N_4602);
nor U9953 (N_9953,N_5023,N_7226);
xor U9954 (N_9954,N_5356,N_7778);
and U9955 (N_9955,N_5895,N_5197);
or U9956 (N_9956,N_5170,N_4918);
nor U9957 (N_9957,N_5629,N_6356);
and U9958 (N_9958,N_7289,N_4561);
nor U9959 (N_9959,N_7545,N_6701);
or U9960 (N_9960,N_4012,N_7428);
or U9961 (N_9961,N_6782,N_7665);
or U9962 (N_9962,N_6722,N_5229);
nor U9963 (N_9963,N_7412,N_6056);
nand U9964 (N_9964,N_4582,N_4959);
nor U9965 (N_9965,N_4212,N_5203);
nor U9966 (N_9966,N_5876,N_7950);
or U9967 (N_9967,N_7072,N_5161);
nor U9968 (N_9968,N_4321,N_6997);
nor U9969 (N_9969,N_6044,N_7687);
nor U9970 (N_9970,N_6327,N_6820);
nand U9971 (N_9971,N_6826,N_7221);
and U9972 (N_9972,N_5669,N_5022);
and U9973 (N_9973,N_6227,N_7225);
xnor U9974 (N_9974,N_7959,N_7328);
and U9975 (N_9975,N_5363,N_6899);
nand U9976 (N_9976,N_7625,N_4055);
nor U9977 (N_9977,N_7640,N_7842);
and U9978 (N_9978,N_7953,N_5157);
or U9979 (N_9979,N_4896,N_4915);
or U9980 (N_9980,N_6517,N_5012);
nor U9981 (N_9981,N_6944,N_6894);
nand U9982 (N_9982,N_7244,N_6572);
and U9983 (N_9983,N_5468,N_5075);
xor U9984 (N_9984,N_5825,N_4464);
xnor U9985 (N_9985,N_4529,N_4038);
xor U9986 (N_9986,N_5802,N_7768);
and U9987 (N_9987,N_7050,N_5623);
nor U9988 (N_9988,N_6924,N_6280);
or U9989 (N_9989,N_6252,N_7253);
nand U9990 (N_9990,N_6155,N_4059);
and U9991 (N_9991,N_6962,N_4720);
and U9992 (N_9992,N_5210,N_5597);
and U9993 (N_9993,N_4525,N_5388);
and U9994 (N_9994,N_4695,N_4649);
xnor U9995 (N_9995,N_6760,N_6187);
and U9996 (N_9996,N_4974,N_4236);
xnor U9997 (N_9997,N_6170,N_7116);
or U9998 (N_9998,N_6730,N_7290);
nand U9999 (N_9999,N_4452,N_7426);
xnor U10000 (N_10000,N_7743,N_4607);
nand U10001 (N_10001,N_7363,N_6353);
and U10002 (N_10002,N_4497,N_7527);
xnor U10003 (N_10003,N_7365,N_4769);
xor U10004 (N_10004,N_5249,N_4195);
xor U10005 (N_10005,N_6496,N_7597);
or U10006 (N_10006,N_6561,N_4870);
xnor U10007 (N_10007,N_5800,N_7465);
nor U10008 (N_10008,N_6045,N_5851);
nand U10009 (N_10009,N_4283,N_5951);
nand U10010 (N_10010,N_6332,N_5744);
nand U10011 (N_10011,N_7809,N_5057);
or U10012 (N_10012,N_5400,N_5451);
or U10013 (N_10013,N_4305,N_4532);
xor U10014 (N_10014,N_7214,N_4909);
or U10015 (N_10015,N_4944,N_6806);
or U10016 (N_10016,N_6102,N_4022);
nor U10017 (N_10017,N_4731,N_4972);
nand U10018 (N_10018,N_5092,N_6958);
xnor U10019 (N_10019,N_4005,N_7518);
nor U10020 (N_10020,N_5174,N_6509);
and U10021 (N_10021,N_6153,N_5506);
xnor U10022 (N_10022,N_6344,N_6259);
nand U10023 (N_10023,N_6875,N_4690);
or U10024 (N_10024,N_6605,N_5026);
xnor U10025 (N_10025,N_6166,N_6951);
and U10026 (N_10026,N_4248,N_5608);
nor U10027 (N_10027,N_6651,N_6628);
and U10028 (N_10028,N_5713,N_4513);
nand U10029 (N_10029,N_7126,N_6340);
nand U10030 (N_10030,N_4542,N_6383);
or U10031 (N_10031,N_4545,N_5380);
nor U10032 (N_10032,N_4557,N_4085);
nor U10033 (N_10033,N_4836,N_6864);
xor U10034 (N_10034,N_4636,N_5612);
nand U10035 (N_10035,N_5195,N_5788);
and U10036 (N_10036,N_7958,N_4207);
nor U10037 (N_10037,N_6438,N_4956);
nor U10038 (N_10038,N_4420,N_7129);
nand U10039 (N_10039,N_7711,N_5724);
and U10040 (N_10040,N_4945,N_6056);
nor U10041 (N_10041,N_5575,N_7306);
xor U10042 (N_10042,N_4615,N_4298);
or U10043 (N_10043,N_7991,N_6780);
nor U10044 (N_10044,N_7843,N_4473);
and U10045 (N_10045,N_6088,N_6227);
or U10046 (N_10046,N_7221,N_4494);
and U10047 (N_10047,N_7389,N_7883);
or U10048 (N_10048,N_5614,N_6039);
xor U10049 (N_10049,N_5068,N_7217);
nand U10050 (N_10050,N_6024,N_7326);
and U10051 (N_10051,N_5507,N_7105);
nor U10052 (N_10052,N_6497,N_6680);
nand U10053 (N_10053,N_6334,N_7591);
nand U10054 (N_10054,N_6434,N_5019);
nor U10055 (N_10055,N_7109,N_7562);
nand U10056 (N_10056,N_4606,N_6232);
xnor U10057 (N_10057,N_7500,N_5552);
and U10058 (N_10058,N_4264,N_6476);
nor U10059 (N_10059,N_7109,N_4681);
or U10060 (N_10060,N_6790,N_7216);
nor U10061 (N_10061,N_4797,N_5830);
and U10062 (N_10062,N_4837,N_7201);
xor U10063 (N_10063,N_7838,N_6319);
or U10064 (N_10064,N_4834,N_6266);
nor U10065 (N_10065,N_6741,N_5813);
nand U10066 (N_10066,N_4431,N_4367);
xnor U10067 (N_10067,N_5963,N_6174);
nor U10068 (N_10068,N_6064,N_4195);
or U10069 (N_10069,N_4448,N_7331);
or U10070 (N_10070,N_4379,N_7112);
nand U10071 (N_10071,N_7786,N_7601);
and U10072 (N_10072,N_5417,N_7635);
and U10073 (N_10073,N_7184,N_7412);
and U10074 (N_10074,N_5324,N_5727);
or U10075 (N_10075,N_4603,N_4009);
or U10076 (N_10076,N_7032,N_4074);
or U10077 (N_10077,N_6426,N_4663);
nand U10078 (N_10078,N_6341,N_5608);
and U10079 (N_10079,N_5480,N_7347);
or U10080 (N_10080,N_6381,N_6884);
or U10081 (N_10081,N_4446,N_7831);
and U10082 (N_10082,N_5205,N_5822);
nand U10083 (N_10083,N_6599,N_7231);
and U10084 (N_10084,N_5097,N_7283);
xor U10085 (N_10085,N_7616,N_5657);
or U10086 (N_10086,N_5097,N_5601);
or U10087 (N_10087,N_4639,N_7053);
nor U10088 (N_10088,N_4175,N_7476);
nand U10089 (N_10089,N_6766,N_7309);
and U10090 (N_10090,N_4226,N_7853);
or U10091 (N_10091,N_6268,N_5938);
xnor U10092 (N_10092,N_4792,N_6724);
xnor U10093 (N_10093,N_5553,N_7849);
nand U10094 (N_10094,N_5608,N_4569);
and U10095 (N_10095,N_5921,N_7908);
xnor U10096 (N_10096,N_4771,N_6970);
xnor U10097 (N_10097,N_5702,N_4021);
or U10098 (N_10098,N_6005,N_6029);
nand U10099 (N_10099,N_5541,N_6549);
nor U10100 (N_10100,N_5063,N_7396);
xnor U10101 (N_10101,N_6806,N_5166);
nor U10102 (N_10102,N_5038,N_7318);
and U10103 (N_10103,N_4453,N_4277);
xnor U10104 (N_10104,N_6997,N_4180);
nor U10105 (N_10105,N_6913,N_5497);
or U10106 (N_10106,N_6061,N_5172);
and U10107 (N_10107,N_6448,N_5264);
xnor U10108 (N_10108,N_6333,N_6070);
or U10109 (N_10109,N_7780,N_4527);
or U10110 (N_10110,N_7009,N_7711);
nand U10111 (N_10111,N_7455,N_5676);
nor U10112 (N_10112,N_6172,N_5305);
nor U10113 (N_10113,N_4393,N_7661);
nand U10114 (N_10114,N_5168,N_4895);
or U10115 (N_10115,N_4454,N_5322);
or U10116 (N_10116,N_4090,N_7192);
nor U10117 (N_10117,N_4462,N_4015);
xor U10118 (N_10118,N_7319,N_5197);
and U10119 (N_10119,N_5111,N_6530);
nand U10120 (N_10120,N_5149,N_5301);
xor U10121 (N_10121,N_5179,N_6935);
and U10122 (N_10122,N_5763,N_6885);
xnor U10123 (N_10123,N_6215,N_6567);
nor U10124 (N_10124,N_5798,N_7241);
xor U10125 (N_10125,N_6071,N_4654);
and U10126 (N_10126,N_7768,N_4746);
nor U10127 (N_10127,N_5855,N_5275);
xor U10128 (N_10128,N_4400,N_6046);
and U10129 (N_10129,N_5237,N_6753);
xor U10130 (N_10130,N_6973,N_6690);
nor U10131 (N_10131,N_5814,N_5657);
nand U10132 (N_10132,N_5445,N_4148);
xnor U10133 (N_10133,N_5617,N_5647);
and U10134 (N_10134,N_4438,N_5854);
and U10135 (N_10135,N_7166,N_6833);
xor U10136 (N_10136,N_6332,N_5527);
xor U10137 (N_10137,N_7041,N_7164);
and U10138 (N_10138,N_5985,N_7247);
nor U10139 (N_10139,N_5645,N_4108);
nand U10140 (N_10140,N_6993,N_6937);
nand U10141 (N_10141,N_4691,N_5562);
or U10142 (N_10142,N_4720,N_5802);
and U10143 (N_10143,N_7104,N_5039);
and U10144 (N_10144,N_7712,N_4850);
or U10145 (N_10145,N_5138,N_5116);
and U10146 (N_10146,N_4957,N_5899);
nand U10147 (N_10147,N_7534,N_6149);
nor U10148 (N_10148,N_5914,N_7461);
or U10149 (N_10149,N_6500,N_7680);
nor U10150 (N_10150,N_5387,N_6150);
nor U10151 (N_10151,N_4460,N_6380);
xnor U10152 (N_10152,N_4115,N_6044);
and U10153 (N_10153,N_7647,N_7407);
nor U10154 (N_10154,N_5617,N_6957);
xnor U10155 (N_10155,N_6664,N_6815);
nand U10156 (N_10156,N_5555,N_6048);
xnor U10157 (N_10157,N_4476,N_5293);
or U10158 (N_10158,N_5564,N_5276);
nand U10159 (N_10159,N_7299,N_5766);
nand U10160 (N_10160,N_5815,N_5952);
xor U10161 (N_10161,N_7588,N_7881);
or U10162 (N_10162,N_5630,N_7443);
and U10163 (N_10163,N_4312,N_6182);
xor U10164 (N_10164,N_6282,N_4791);
xnor U10165 (N_10165,N_7864,N_6250);
and U10166 (N_10166,N_5906,N_5919);
and U10167 (N_10167,N_6787,N_4483);
nand U10168 (N_10168,N_6847,N_6199);
xnor U10169 (N_10169,N_7935,N_7447);
nand U10170 (N_10170,N_4735,N_4068);
nor U10171 (N_10171,N_7812,N_5227);
or U10172 (N_10172,N_6676,N_6812);
nor U10173 (N_10173,N_5477,N_4768);
and U10174 (N_10174,N_4828,N_4479);
xnor U10175 (N_10175,N_5210,N_7061);
xor U10176 (N_10176,N_4703,N_5577);
xor U10177 (N_10177,N_5337,N_6579);
nor U10178 (N_10178,N_6107,N_6125);
xnor U10179 (N_10179,N_7279,N_4547);
or U10180 (N_10180,N_7793,N_6400);
nor U10181 (N_10181,N_4572,N_5074);
nand U10182 (N_10182,N_4732,N_6646);
and U10183 (N_10183,N_6211,N_6061);
nor U10184 (N_10184,N_4005,N_5640);
xnor U10185 (N_10185,N_6568,N_5519);
or U10186 (N_10186,N_5825,N_4687);
nand U10187 (N_10187,N_5022,N_4270);
nand U10188 (N_10188,N_5614,N_4287);
or U10189 (N_10189,N_5746,N_7266);
and U10190 (N_10190,N_5922,N_6829);
xnor U10191 (N_10191,N_5173,N_5900);
nor U10192 (N_10192,N_6514,N_7577);
or U10193 (N_10193,N_5833,N_7471);
xnor U10194 (N_10194,N_6948,N_6989);
or U10195 (N_10195,N_4807,N_4281);
xnor U10196 (N_10196,N_7471,N_4398);
nand U10197 (N_10197,N_5005,N_7897);
and U10198 (N_10198,N_7108,N_7144);
nand U10199 (N_10199,N_5700,N_5689);
and U10200 (N_10200,N_4863,N_7964);
xor U10201 (N_10201,N_4749,N_7244);
and U10202 (N_10202,N_5693,N_5395);
nand U10203 (N_10203,N_4144,N_5126);
xor U10204 (N_10204,N_5797,N_4244);
or U10205 (N_10205,N_6358,N_6411);
xnor U10206 (N_10206,N_5244,N_5800);
xnor U10207 (N_10207,N_6792,N_6703);
nand U10208 (N_10208,N_7944,N_5289);
and U10209 (N_10209,N_6121,N_4631);
and U10210 (N_10210,N_6169,N_4262);
nand U10211 (N_10211,N_5535,N_7055);
xnor U10212 (N_10212,N_4133,N_7036);
xnor U10213 (N_10213,N_4737,N_6325);
and U10214 (N_10214,N_4883,N_5496);
or U10215 (N_10215,N_7565,N_6293);
and U10216 (N_10216,N_5696,N_5859);
nor U10217 (N_10217,N_6749,N_7986);
and U10218 (N_10218,N_6845,N_5414);
and U10219 (N_10219,N_4160,N_7673);
xor U10220 (N_10220,N_4124,N_6146);
nor U10221 (N_10221,N_4884,N_7135);
nand U10222 (N_10222,N_7580,N_4975);
or U10223 (N_10223,N_4526,N_5886);
xor U10224 (N_10224,N_5293,N_4112);
xor U10225 (N_10225,N_5072,N_4138);
nor U10226 (N_10226,N_4137,N_7526);
nor U10227 (N_10227,N_4498,N_7931);
xor U10228 (N_10228,N_5853,N_7033);
and U10229 (N_10229,N_7796,N_5616);
nand U10230 (N_10230,N_4651,N_7418);
or U10231 (N_10231,N_4439,N_4751);
and U10232 (N_10232,N_7259,N_6296);
nand U10233 (N_10233,N_4663,N_4174);
nor U10234 (N_10234,N_5798,N_4583);
and U10235 (N_10235,N_7487,N_6522);
and U10236 (N_10236,N_5329,N_4171);
nand U10237 (N_10237,N_5367,N_7771);
xnor U10238 (N_10238,N_7010,N_4481);
and U10239 (N_10239,N_4845,N_6953);
or U10240 (N_10240,N_6853,N_5211);
or U10241 (N_10241,N_7848,N_4620);
nand U10242 (N_10242,N_7448,N_4314);
xor U10243 (N_10243,N_5894,N_4037);
nor U10244 (N_10244,N_6862,N_5262);
or U10245 (N_10245,N_7368,N_5274);
xor U10246 (N_10246,N_6606,N_4796);
and U10247 (N_10247,N_7436,N_5265);
xnor U10248 (N_10248,N_7341,N_6200);
and U10249 (N_10249,N_6875,N_5998);
nand U10250 (N_10250,N_7797,N_6314);
or U10251 (N_10251,N_5142,N_5759);
nand U10252 (N_10252,N_5315,N_7296);
or U10253 (N_10253,N_7108,N_5157);
xor U10254 (N_10254,N_6871,N_5392);
or U10255 (N_10255,N_7121,N_7221);
nor U10256 (N_10256,N_7484,N_4732);
and U10257 (N_10257,N_5407,N_7436);
or U10258 (N_10258,N_4779,N_7639);
nand U10259 (N_10259,N_7722,N_5655);
nor U10260 (N_10260,N_5263,N_5589);
xor U10261 (N_10261,N_5817,N_4689);
and U10262 (N_10262,N_4599,N_4701);
nand U10263 (N_10263,N_5110,N_6669);
nand U10264 (N_10264,N_6835,N_5420);
or U10265 (N_10265,N_6204,N_7857);
nand U10266 (N_10266,N_7384,N_5938);
or U10267 (N_10267,N_6590,N_6991);
xor U10268 (N_10268,N_4156,N_4464);
or U10269 (N_10269,N_5238,N_7011);
xor U10270 (N_10270,N_6085,N_5264);
xnor U10271 (N_10271,N_7987,N_4716);
nand U10272 (N_10272,N_6056,N_7738);
nor U10273 (N_10273,N_5493,N_5389);
xor U10274 (N_10274,N_5205,N_5463);
nand U10275 (N_10275,N_6864,N_4070);
nand U10276 (N_10276,N_5430,N_7073);
nand U10277 (N_10277,N_7559,N_6652);
xor U10278 (N_10278,N_6661,N_4874);
or U10279 (N_10279,N_7160,N_7916);
xor U10280 (N_10280,N_4902,N_4322);
nor U10281 (N_10281,N_6443,N_6705);
xnor U10282 (N_10282,N_7173,N_4350);
nand U10283 (N_10283,N_6641,N_5843);
and U10284 (N_10284,N_6147,N_4475);
nand U10285 (N_10285,N_6520,N_7479);
or U10286 (N_10286,N_6999,N_4884);
or U10287 (N_10287,N_5380,N_7363);
or U10288 (N_10288,N_4958,N_4815);
and U10289 (N_10289,N_7766,N_4815);
xor U10290 (N_10290,N_5136,N_7040);
xnor U10291 (N_10291,N_5535,N_7149);
or U10292 (N_10292,N_5252,N_6227);
nor U10293 (N_10293,N_7954,N_5307);
nand U10294 (N_10294,N_5457,N_5612);
and U10295 (N_10295,N_6017,N_4944);
nand U10296 (N_10296,N_5743,N_7791);
nand U10297 (N_10297,N_6850,N_4178);
nand U10298 (N_10298,N_7341,N_6193);
nor U10299 (N_10299,N_6180,N_6007);
or U10300 (N_10300,N_4858,N_6842);
or U10301 (N_10301,N_6836,N_6873);
or U10302 (N_10302,N_6313,N_7785);
nor U10303 (N_10303,N_7032,N_7167);
nand U10304 (N_10304,N_4005,N_6584);
or U10305 (N_10305,N_4299,N_7682);
and U10306 (N_10306,N_5030,N_6290);
nand U10307 (N_10307,N_7553,N_7001);
and U10308 (N_10308,N_5135,N_5339);
nor U10309 (N_10309,N_4536,N_7101);
nand U10310 (N_10310,N_4291,N_6595);
xor U10311 (N_10311,N_5560,N_7140);
nor U10312 (N_10312,N_6570,N_4134);
nor U10313 (N_10313,N_6919,N_6807);
nor U10314 (N_10314,N_5050,N_5528);
xnor U10315 (N_10315,N_4408,N_7062);
and U10316 (N_10316,N_7186,N_4959);
or U10317 (N_10317,N_7226,N_4653);
xnor U10318 (N_10318,N_5779,N_5448);
or U10319 (N_10319,N_5637,N_6860);
nor U10320 (N_10320,N_6301,N_7825);
nand U10321 (N_10321,N_7549,N_5885);
nor U10322 (N_10322,N_7532,N_7992);
and U10323 (N_10323,N_6980,N_6862);
nand U10324 (N_10324,N_5382,N_4974);
nor U10325 (N_10325,N_6662,N_5305);
or U10326 (N_10326,N_7128,N_7760);
or U10327 (N_10327,N_6334,N_7209);
and U10328 (N_10328,N_4960,N_7121);
or U10329 (N_10329,N_6916,N_5997);
and U10330 (N_10330,N_7393,N_7067);
nor U10331 (N_10331,N_5815,N_6488);
and U10332 (N_10332,N_4861,N_4569);
and U10333 (N_10333,N_6343,N_5389);
nand U10334 (N_10334,N_6900,N_6742);
or U10335 (N_10335,N_6888,N_6601);
and U10336 (N_10336,N_7860,N_6705);
nand U10337 (N_10337,N_5417,N_4981);
xnor U10338 (N_10338,N_5516,N_7079);
and U10339 (N_10339,N_7971,N_6344);
or U10340 (N_10340,N_6722,N_7790);
or U10341 (N_10341,N_6484,N_6315);
xor U10342 (N_10342,N_7104,N_5922);
nor U10343 (N_10343,N_5485,N_6914);
nand U10344 (N_10344,N_5229,N_5186);
xor U10345 (N_10345,N_5265,N_6718);
and U10346 (N_10346,N_5025,N_7041);
nor U10347 (N_10347,N_5062,N_6820);
xor U10348 (N_10348,N_6242,N_7315);
xor U10349 (N_10349,N_7785,N_6228);
xor U10350 (N_10350,N_5602,N_5011);
and U10351 (N_10351,N_7933,N_6804);
or U10352 (N_10352,N_5372,N_7172);
and U10353 (N_10353,N_6014,N_7205);
and U10354 (N_10354,N_4561,N_7854);
and U10355 (N_10355,N_4452,N_5318);
nor U10356 (N_10356,N_6176,N_5560);
and U10357 (N_10357,N_5325,N_6276);
nand U10358 (N_10358,N_6658,N_7660);
xnor U10359 (N_10359,N_4099,N_6707);
and U10360 (N_10360,N_7772,N_7095);
xnor U10361 (N_10361,N_7727,N_5712);
and U10362 (N_10362,N_7567,N_7460);
or U10363 (N_10363,N_6229,N_4875);
nand U10364 (N_10364,N_7720,N_6328);
or U10365 (N_10365,N_5185,N_4804);
nand U10366 (N_10366,N_5759,N_5900);
xor U10367 (N_10367,N_4066,N_7384);
or U10368 (N_10368,N_6901,N_4902);
xor U10369 (N_10369,N_4142,N_5101);
nor U10370 (N_10370,N_4011,N_7623);
nand U10371 (N_10371,N_7759,N_7934);
xor U10372 (N_10372,N_5837,N_4625);
nand U10373 (N_10373,N_5637,N_7983);
xnor U10374 (N_10374,N_4965,N_6274);
nand U10375 (N_10375,N_6153,N_4012);
nor U10376 (N_10376,N_5509,N_6504);
and U10377 (N_10377,N_5920,N_6640);
and U10378 (N_10378,N_4976,N_5869);
nand U10379 (N_10379,N_4102,N_4571);
xnor U10380 (N_10380,N_7927,N_6467);
nor U10381 (N_10381,N_7730,N_4093);
nor U10382 (N_10382,N_5070,N_5358);
nand U10383 (N_10383,N_6730,N_6292);
nand U10384 (N_10384,N_4581,N_7262);
and U10385 (N_10385,N_6096,N_4076);
and U10386 (N_10386,N_4502,N_5398);
nor U10387 (N_10387,N_5906,N_5229);
or U10388 (N_10388,N_5705,N_4551);
and U10389 (N_10389,N_5790,N_7174);
xnor U10390 (N_10390,N_6097,N_7776);
nor U10391 (N_10391,N_4024,N_5965);
xnor U10392 (N_10392,N_7510,N_5232);
and U10393 (N_10393,N_5995,N_7464);
nor U10394 (N_10394,N_5599,N_4417);
nor U10395 (N_10395,N_6779,N_7181);
xnor U10396 (N_10396,N_5771,N_6088);
or U10397 (N_10397,N_6140,N_6525);
nor U10398 (N_10398,N_4743,N_7764);
and U10399 (N_10399,N_4630,N_5588);
nor U10400 (N_10400,N_7068,N_4151);
and U10401 (N_10401,N_7963,N_5293);
and U10402 (N_10402,N_5010,N_7023);
or U10403 (N_10403,N_4104,N_4113);
xnor U10404 (N_10404,N_5298,N_5029);
xnor U10405 (N_10405,N_5411,N_6782);
xnor U10406 (N_10406,N_5101,N_5240);
and U10407 (N_10407,N_4161,N_7022);
xor U10408 (N_10408,N_6540,N_5246);
xnor U10409 (N_10409,N_5297,N_4108);
nor U10410 (N_10410,N_5136,N_4180);
and U10411 (N_10411,N_6202,N_7403);
or U10412 (N_10412,N_4156,N_7027);
nor U10413 (N_10413,N_7094,N_6128);
or U10414 (N_10414,N_5211,N_4204);
and U10415 (N_10415,N_6334,N_6174);
and U10416 (N_10416,N_7607,N_6227);
nand U10417 (N_10417,N_5699,N_4884);
or U10418 (N_10418,N_6464,N_6962);
nand U10419 (N_10419,N_6436,N_4897);
nand U10420 (N_10420,N_4278,N_4294);
or U10421 (N_10421,N_5279,N_7003);
or U10422 (N_10422,N_6323,N_7634);
nand U10423 (N_10423,N_6805,N_6448);
xor U10424 (N_10424,N_5580,N_7180);
xor U10425 (N_10425,N_5328,N_4365);
nand U10426 (N_10426,N_4118,N_7745);
and U10427 (N_10427,N_7387,N_7827);
and U10428 (N_10428,N_7995,N_4281);
nand U10429 (N_10429,N_7396,N_5833);
or U10430 (N_10430,N_6966,N_4437);
or U10431 (N_10431,N_5177,N_6127);
xnor U10432 (N_10432,N_6803,N_5285);
or U10433 (N_10433,N_6196,N_5886);
xor U10434 (N_10434,N_6926,N_5535);
xnor U10435 (N_10435,N_7834,N_6080);
or U10436 (N_10436,N_5961,N_4593);
and U10437 (N_10437,N_7705,N_5491);
xnor U10438 (N_10438,N_5707,N_5591);
nor U10439 (N_10439,N_6031,N_4397);
xor U10440 (N_10440,N_7467,N_5499);
and U10441 (N_10441,N_7978,N_4790);
nand U10442 (N_10442,N_7359,N_6062);
or U10443 (N_10443,N_4687,N_6666);
or U10444 (N_10444,N_7096,N_5209);
or U10445 (N_10445,N_4605,N_4187);
nand U10446 (N_10446,N_5316,N_5364);
nand U10447 (N_10447,N_7781,N_6924);
xor U10448 (N_10448,N_4167,N_4407);
nor U10449 (N_10449,N_6129,N_6889);
or U10450 (N_10450,N_5991,N_6018);
and U10451 (N_10451,N_6756,N_6604);
nor U10452 (N_10452,N_7373,N_5162);
nand U10453 (N_10453,N_5251,N_7959);
or U10454 (N_10454,N_5789,N_7591);
xor U10455 (N_10455,N_5230,N_7557);
xor U10456 (N_10456,N_7909,N_6241);
or U10457 (N_10457,N_7302,N_4850);
xor U10458 (N_10458,N_7502,N_7996);
and U10459 (N_10459,N_5752,N_5953);
and U10460 (N_10460,N_5871,N_7771);
xor U10461 (N_10461,N_7482,N_5451);
or U10462 (N_10462,N_4729,N_6545);
xor U10463 (N_10463,N_5565,N_4261);
and U10464 (N_10464,N_6601,N_5013);
xor U10465 (N_10465,N_4920,N_4312);
or U10466 (N_10466,N_7979,N_6857);
and U10467 (N_10467,N_4652,N_7700);
nand U10468 (N_10468,N_4958,N_4980);
and U10469 (N_10469,N_4449,N_7114);
nor U10470 (N_10470,N_4265,N_5268);
nor U10471 (N_10471,N_7630,N_4496);
and U10472 (N_10472,N_4752,N_4998);
or U10473 (N_10473,N_4098,N_7899);
or U10474 (N_10474,N_4709,N_5866);
and U10475 (N_10475,N_4258,N_7946);
and U10476 (N_10476,N_7690,N_6597);
and U10477 (N_10477,N_6496,N_6583);
and U10478 (N_10478,N_5042,N_7957);
nor U10479 (N_10479,N_7677,N_6326);
or U10480 (N_10480,N_5629,N_7027);
nor U10481 (N_10481,N_7036,N_5555);
xnor U10482 (N_10482,N_4063,N_5468);
xor U10483 (N_10483,N_4020,N_5456);
nor U10484 (N_10484,N_7032,N_4527);
and U10485 (N_10485,N_7989,N_6681);
xnor U10486 (N_10486,N_4918,N_6366);
xor U10487 (N_10487,N_6033,N_5970);
nand U10488 (N_10488,N_6554,N_7743);
or U10489 (N_10489,N_7358,N_5537);
xor U10490 (N_10490,N_4546,N_7452);
or U10491 (N_10491,N_4894,N_6169);
and U10492 (N_10492,N_4405,N_5773);
nand U10493 (N_10493,N_4967,N_4737);
nand U10494 (N_10494,N_4544,N_4886);
nor U10495 (N_10495,N_7134,N_7389);
nor U10496 (N_10496,N_7629,N_7371);
nand U10497 (N_10497,N_4781,N_6737);
and U10498 (N_10498,N_4038,N_4628);
nor U10499 (N_10499,N_5897,N_7387);
xnor U10500 (N_10500,N_6579,N_5219);
and U10501 (N_10501,N_4231,N_5417);
or U10502 (N_10502,N_5036,N_4668);
or U10503 (N_10503,N_4777,N_6714);
and U10504 (N_10504,N_5066,N_4241);
and U10505 (N_10505,N_7484,N_6606);
nand U10506 (N_10506,N_4434,N_4439);
and U10507 (N_10507,N_7139,N_5870);
or U10508 (N_10508,N_5712,N_7971);
nor U10509 (N_10509,N_5286,N_5899);
and U10510 (N_10510,N_5919,N_4776);
nor U10511 (N_10511,N_4351,N_5659);
nand U10512 (N_10512,N_4089,N_7963);
nor U10513 (N_10513,N_5023,N_5865);
or U10514 (N_10514,N_7833,N_5457);
and U10515 (N_10515,N_4330,N_5821);
or U10516 (N_10516,N_5817,N_5163);
or U10517 (N_10517,N_4345,N_7028);
nor U10518 (N_10518,N_7871,N_5435);
xor U10519 (N_10519,N_7859,N_6820);
and U10520 (N_10520,N_6352,N_6793);
and U10521 (N_10521,N_7724,N_4431);
xnor U10522 (N_10522,N_6658,N_6565);
and U10523 (N_10523,N_4532,N_6667);
nand U10524 (N_10524,N_4880,N_6118);
or U10525 (N_10525,N_6464,N_7948);
or U10526 (N_10526,N_5293,N_4012);
nor U10527 (N_10527,N_4041,N_6552);
and U10528 (N_10528,N_4693,N_4912);
nand U10529 (N_10529,N_4894,N_6843);
nor U10530 (N_10530,N_7609,N_6534);
nor U10531 (N_10531,N_7084,N_4265);
nand U10532 (N_10532,N_5270,N_7907);
nand U10533 (N_10533,N_4070,N_6514);
and U10534 (N_10534,N_7293,N_5258);
xor U10535 (N_10535,N_6545,N_4809);
xor U10536 (N_10536,N_7529,N_7443);
and U10537 (N_10537,N_7388,N_4786);
or U10538 (N_10538,N_4361,N_7388);
and U10539 (N_10539,N_4530,N_6272);
nand U10540 (N_10540,N_6260,N_4434);
or U10541 (N_10541,N_6369,N_5995);
xor U10542 (N_10542,N_7774,N_6957);
xor U10543 (N_10543,N_6811,N_6148);
nand U10544 (N_10544,N_7478,N_4298);
nor U10545 (N_10545,N_6716,N_7418);
xnor U10546 (N_10546,N_5269,N_5153);
xnor U10547 (N_10547,N_6841,N_6783);
and U10548 (N_10548,N_5030,N_4093);
xor U10549 (N_10549,N_5072,N_4625);
nand U10550 (N_10550,N_7197,N_7589);
xor U10551 (N_10551,N_5065,N_6206);
or U10552 (N_10552,N_4649,N_7115);
nand U10553 (N_10553,N_7641,N_7428);
nor U10554 (N_10554,N_7964,N_5345);
or U10555 (N_10555,N_6195,N_5425);
and U10556 (N_10556,N_5956,N_6034);
nor U10557 (N_10557,N_4131,N_4627);
xnor U10558 (N_10558,N_4895,N_6581);
and U10559 (N_10559,N_4352,N_6185);
and U10560 (N_10560,N_4798,N_7205);
or U10561 (N_10561,N_4113,N_4465);
or U10562 (N_10562,N_6100,N_4940);
or U10563 (N_10563,N_7040,N_4191);
and U10564 (N_10564,N_6366,N_4725);
nand U10565 (N_10565,N_7250,N_6933);
nand U10566 (N_10566,N_7218,N_7157);
nor U10567 (N_10567,N_5178,N_4128);
or U10568 (N_10568,N_5811,N_5376);
nand U10569 (N_10569,N_5023,N_5633);
nand U10570 (N_10570,N_4317,N_6710);
xnor U10571 (N_10571,N_7510,N_5352);
or U10572 (N_10572,N_6320,N_4305);
nor U10573 (N_10573,N_5126,N_7492);
nor U10574 (N_10574,N_5158,N_5284);
nand U10575 (N_10575,N_6392,N_6597);
or U10576 (N_10576,N_6136,N_4473);
nor U10577 (N_10577,N_7599,N_5038);
and U10578 (N_10578,N_6023,N_4346);
nor U10579 (N_10579,N_6855,N_6464);
xor U10580 (N_10580,N_4626,N_7336);
nand U10581 (N_10581,N_5401,N_6640);
nand U10582 (N_10582,N_6576,N_6884);
nand U10583 (N_10583,N_5405,N_7295);
and U10584 (N_10584,N_5152,N_6165);
nand U10585 (N_10585,N_4506,N_4397);
or U10586 (N_10586,N_4239,N_4691);
nor U10587 (N_10587,N_5413,N_5801);
and U10588 (N_10588,N_5959,N_5270);
and U10589 (N_10589,N_5559,N_6980);
xnor U10590 (N_10590,N_4322,N_4703);
xor U10591 (N_10591,N_6512,N_6588);
and U10592 (N_10592,N_7050,N_6793);
nand U10593 (N_10593,N_4447,N_6420);
nor U10594 (N_10594,N_4991,N_5925);
nand U10595 (N_10595,N_5813,N_5022);
or U10596 (N_10596,N_7811,N_5493);
xor U10597 (N_10597,N_5183,N_6836);
or U10598 (N_10598,N_6519,N_6942);
nand U10599 (N_10599,N_7002,N_7350);
nor U10600 (N_10600,N_5289,N_6360);
and U10601 (N_10601,N_4928,N_6157);
nand U10602 (N_10602,N_7588,N_7224);
and U10603 (N_10603,N_6815,N_6915);
xnor U10604 (N_10604,N_4759,N_6853);
or U10605 (N_10605,N_7939,N_5589);
nor U10606 (N_10606,N_6667,N_4918);
or U10607 (N_10607,N_6625,N_6628);
nand U10608 (N_10608,N_7609,N_6010);
or U10609 (N_10609,N_6147,N_6451);
or U10610 (N_10610,N_5728,N_5607);
and U10611 (N_10611,N_4231,N_6578);
nand U10612 (N_10612,N_5145,N_5746);
nor U10613 (N_10613,N_5600,N_7652);
nor U10614 (N_10614,N_5226,N_6361);
nand U10615 (N_10615,N_4508,N_6560);
nand U10616 (N_10616,N_6088,N_4598);
xnor U10617 (N_10617,N_6912,N_7847);
nand U10618 (N_10618,N_7787,N_7465);
nand U10619 (N_10619,N_6926,N_7137);
nor U10620 (N_10620,N_6731,N_6050);
nor U10621 (N_10621,N_7360,N_5033);
nor U10622 (N_10622,N_5832,N_6260);
nand U10623 (N_10623,N_6721,N_4593);
nor U10624 (N_10624,N_4308,N_5945);
or U10625 (N_10625,N_5603,N_4366);
and U10626 (N_10626,N_4832,N_5925);
and U10627 (N_10627,N_7412,N_4530);
xor U10628 (N_10628,N_5901,N_5479);
or U10629 (N_10629,N_4586,N_5555);
and U10630 (N_10630,N_6535,N_5586);
nand U10631 (N_10631,N_7504,N_5305);
nand U10632 (N_10632,N_5878,N_6272);
and U10633 (N_10633,N_7931,N_4572);
or U10634 (N_10634,N_4385,N_4263);
xor U10635 (N_10635,N_7210,N_5953);
xor U10636 (N_10636,N_6573,N_4190);
xnor U10637 (N_10637,N_6155,N_6452);
xor U10638 (N_10638,N_6413,N_4169);
xnor U10639 (N_10639,N_6200,N_6622);
nor U10640 (N_10640,N_6237,N_6886);
and U10641 (N_10641,N_7616,N_6437);
xor U10642 (N_10642,N_4093,N_7001);
and U10643 (N_10643,N_6649,N_6613);
xor U10644 (N_10644,N_7308,N_6310);
nand U10645 (N_10645,N_5435,N_7333);
xor U10646 (N_10646,N_7647,N_5212);
or U10647 (N_10647,N_5957,N_7985);
nand U10648 (N_10648,N_6138,N_7436);
or U10649 (N_10649,N_6116,N_4091);
or U10650 (N_10650,N_7453,N_6323);
xor U10651 (N_10651,N_4483,N_4155);
nand U10652 (N_10652,N_7965,N_4690);
xor U10653 (N_10653,N_7830,N_5782);
and U10654 (N_10654,N_6559,N_5551);
and U10655 (N_10655,N_6104,N_7407);
nor U10656 (N_10656,N_4849,N_7608);
xor U10657 (N_10657,N_4340,N_6786);
nor U10658 (N_10658,N_6644,N_7706);
and U10659 (N_10659,N_7604,N_4553);
nand U10660 (N_10660,N_7092,N_5943);
or U10661 (N_10661,N_7249,N_6934);
nand U10662 (N_10662,N_7733,N_4421);
xnor U10663 (N_10663,N_4943,N_7702);
or U10664 (N_10664,N_5326,N_6171);
or U10665 (N_10665,N_7886,N_4767);
xnor U10666 (N_10666,N_5734,N_7898);
and U10667 (N_10667,N_4020,N_6983);
or U10668 (N_10668,N_4186,N_4558);
nor U10669 (N_10669,N_7500,N_4072);
nand U10670 (N_10670,N_4041,N_7062);
and U10671 (N_10671,N_5057,N_4558);
or U10672 (N_10672,N_4075,N_4213);
xnor U10673 (N_10673,N_4048,N_6266);
and U10674 (N_10674,N_5436,N_4340);
nand U10675 (N_10675,N_5338,N_5843);
nand U10676 (N_10676,N_7321,N_4009);
and U10677 (N_10677,N_5878,N_5622);
or U10678 (N_10678,N_4314,N_7557);
and U10679 (N_10679,N_7372,N_4113);
or U10680 (N_10680,N_6072,N_6745);
or U10681 (N_10681,N_5714,N_4543);
xor U10682 (N_10682,N_6627,N_6950);
nand U10683 (N_10683,N_7541,N_7977);
nand U10684 (N_10684,N_7669,N_5787);
or U10685 (N_10685,N_7672,N_5522);
nor U10686 (N_10686,N_4990,N_5586);
and U10687 (N_10687,N_4168,N_5317);
nor U10688 (N_10688,N_4010,N_6486);
xnor U10689 (N_10689,N_4946,N_5019);
and U10690 (N_10690,N_5229,N_4372);
xor U10691 (N_10691,N_6882,N_4359);
xor U10692 (N_10692,N_7485,N_4591);
nor U10693 (N_10693,N_4997,N_4190);
nand U10694 (N_10694,N_7530,N_7278);
nor U10695 (N_10695,N_5590,N_4439);
nand U10696 (N_10696,N_7045,N_4279);
nand U10697 (N_10697,N_6947,N_6913);
nor U10698 (N_10698,N_4183,N_5430);
xor U10699 (N_10699,N_6096,N_5535);
and U10700 (N_10700,N_4146,N_7883);
nand U10701 (N_10701,N_4546,N_5652);
nor U10702 (N_10702,N_6722,N_4443);
and U10703 (N_10703,N_4765,N_7595);
nand U10704 (N_10704,N_6631,N_5963);
and U10705 (N_10705,N_7840,N_6551);
or U10706 (N_10706,N_6301,N_7419);
nand U10707 (N_10707,N_4457,N_5374);
nor U10708 (N_10708,N_7308,N_6702);
xnor U10709 (N_10709,N_7405,N_5083);
nor U10710 (N_10710,N_5085,N_5919);
and U10711 (N_10711,N_4776,N_4259);
or U10712 (N_10712,N_6241,N_7573);
xnor U10713 (N_10713,N_5757,N_4179);
nand U10714 (N_10714,N_4044,N_7110);
nor U10715 (N_10715,N_4552,N_4323);
and U10716 (N_10716,N_4224,N_5824);
xor U10717 (N_10717,N_7653,N_7609);
xor U10718 (N_10718,N_5083,N_6543);
nor U10719 (N_10719,N_7221,N_7912);
nor U10720 (N_10720,N_7012,N_5183);
nand U10721 (N_10721,N_4880,N_6815);
nand U10722 (N_10722,N_6391,N_4177);
nand U10723 (N_10723,N_6562,N_6587);
xnor U10724 (N_10724,N_6799,N_4677);
xnor U10725 (N_10725,N_7194,N_4525);
or U10726 (N_10726,N_7948,N_7185);
nand U10727 (N_10727,N_6616,N_4137);
nor U10728 (N_10728,N_6083,N_4925);
xnor U10729 (N_10729,N_7021,N_5433);
xor U10730 (N_10730,N_6209,N_5703);
and U10731 (N_10731,N_7262,N_7795);
and U10732 (N_10732,N_4005,N_6201);
nor U10733 (N_10733,N_5650,N_4806);
nand U10734 (N_10734,N_6958,N_6132);
xor U10735 (N_10735,N_5735,N_7547);
or U10736 (N_10736,N_7878,N_4676);
and U10737 (N_10737,N_5607,N_4018);
and U10738 (N_10738,N_4172,N_7060);
or U10739 (N_10739,N_7673,N_6154);
nand U10740 (N_10740,N_7202,N_7178);
xor U10741 (N_10741,N_6938,N_4979);
and U10742 (N_10742,N_6314,N_6471);
nor U10743 (N_10743,N_7380,N_5648);
or U10744 (N_10744,N_6151,N_4619);
xor U10745 (N_10745,N_6120,N_5526);
xnor U10746 (N_10746,N_6358,N_6185);
or U10747 (N_10747,N_4433,N_5440);
xnor U10748 (N_10748,N_7029,N_4176);
xnor U10749 (N_10749,N_5187,N_7598);
nand U10750 (N_10750,N_6470,N_5345);
xor U10751 (N_10751,N_5259,N_5898);
or U10752 (N_10752,N_4752,N_5184);
or U10753 (N_10753,N_7857,N_6240);
nor U10754 (N_10754,N_6302,N_7801);
nand U10755 (N_10755,N_7334,N_6217);
nor U10756 (N_10756,N_6300,N_6843);
xnor U10757 (N_10757,N_7248,N_4592);
or U10758 (N_10758,N_5603,N_7484);
and U10759 (N_10759,N_5044,N_6007);
and U10760 (N_10760,N_6228,N_5286);
nor U10761 (N_10761,N_6037,N_4284);
nor U10762 (N_10762,N_6449,N_5732);
nand U10763 (N_10763,N_5640,N_6937);
nor U10764 (N_10764,N_6146,N_7816);
nor U10765 (N_10765,N_4041,N_4419);
or U10766 (N_10766,N_4978,N_7419);
or U10767 (N_10767,N_4941,N_4263);
xnor U10768 (N_10768,N_4277,N_5682);
xnor U10769 (N_10769,N_4223,N_6797);
nand U10770 (N_10770,N_6255,N_4170);
xnor U10771 (N_10771,N_6640,N_5634);
or U10772 (N_10772,N_7259,N_5102);
xor U10773 (N_10773,N_7519,N_4751);
nand U10774 (N_10774,N_6070,N_6052);
or U10775 (N_10775,N_7922,N_7355);
nor U10776 (N_10776,N_5884,N_4766);
and U10777 (N_10777,N_6567,N_4143);
nand U10778 (N_10778,N_6879,N_4099);
xnor U10779 (N_10779,N_5090,N_5243);
and U10780 (N_10780,N_5665,N_5633);
or U10781 (N_10781,N_7021,N_4817);
or U10782 (N_10782,N_4405,N_7459);
nor U10783 (N_10783,N_7327,N_4403);
nor U10784 (N_10784,N_7256,N_4013);
and U10785 (N_10785,N_5266,N_7671);
nor U10786 (N_10786,N_4449,N_7401);
and U10787 (N_10787,N_4480,N_4020);
xor U10788 (N_10788,N_5341,N_5665);
and U10789 (N_10789,N_4456,N_7764);
nand U10790 (N_10790,N_4856,N_5103);
and U10791 (N_10791,N_7350,N_5086);
and U10792 (N_10792,N_6316,N_4879);
nor U10793 (N_10793,N_4108,N_5729);
and U10794 (N_10794,N_6368,N_5435);
nand U10795 (N_10795,N_6795,N_4503);
nand U10796 (N_10796,N_7997,N_4171);
and U10797 (N_10797,N_6751,N_5747);
nor U10798 (N_10798,N_5190,N_4881);
or U10799 (N_10799,N_6531,N_7759);
xnor U10800 (N_10800,N_4111,N_5068);
nand U10801 (N_10801,N_6004,N_6091);
xor U10802 (N_10802,N_6470,N_4093);
nor U10803 (N_10803,N_6106,N_5643);
xor U10804 (N_10804,N_6214,N_5185);
xnor U10805 (N_10805,N_5828,N_5246);
and U10806 (N_10806,N_6613,N_5459);
nand U10807 (N_10807,N_6212,N_6208);
nor U10808 (N_10808,N_4941,N_4089);
nand U10809 (N_10809,N_7233,N_7146);
nor U10810 (N_10810,N_6738,N_4123);
nand U10811 (N_10811,N_5012,N_7963);
and U10812 (N_10812,N_6717,N_7464);
nor U10813 (N_10813,N_5001,N_6595);
xnor U10814 (N_10814,N_4493,N_6956);
or U10815 (N_10815,N_6059,N_6886);
and U10816 (N_10816,N_4494,N_6721);
or U10817 (N_10817,N_4478,N_5145);
and U10818 (N_10818,N_7228,N_4189);
or U10819 (N_10819,N_5532,N_7069);
or U10820 (N_10820,N_7044,N_5583);
nand U10821 (N_10821,N_4716,N_5738);
nand U10822 (N_10822,N_6549,N_7024);
or U10823 (N_10823,N_7078,N_4207);
xor U10824 (N_10824,N_5232,N_4707);
and U10825 (N_10825,N_5643,N_7652);
nand U10826 (N_10826,N_7276,N_4710);
xor U10827 (N_10827,N_4992,N_4871);
or U10828 (N_10828,N_4434,N_6748);
nor U10829 (N_10829,N_7658,N_6398);
nand U10830 (N_10830,N_5853,N_4313);
nor U10831 (N_10831,N_5323,N_5388);
nand U10832 (N_10832,N_4345,N_7317);
or U10833 (N_10833,N_6360,N_6092);
nand U10834 (N_10834,N_6811,N_5717);
xor U10835 (N_10835,N_6277,N_5643);
or U10836 (N_10836,N_7584,N_6574);
and U10837 (N_10837,N_6337,N_5783);
xor U10838 (N_10838,N_5868,N_5275);
and U10839 (N_10839,N_5560,N_7121);
nand U10840 (N_10840,N_5316,N_4565);
nor U10841 (N_10841,N_5920,N_7478);
nor U10842 (N_10842,N_7690,N_4830);
or U10843 (N_10843,N_4674,N_5780);
nand U10844 (N_10844,N_4226,N_5324);
xor U10845 (N_10845,N_7762,N_6877);
nor U10846 (N_10846,N_4437,N_6236);
and U10847 (N_10847,N_4283,N_7552);
nor U10848 (N_10848,N_4289,N_7850);
and U10849 (N_10849,N_7086,N_5380);
and U10850 (N_10850,N_6314,N_4760);
nor U10851 (N_10851,N_6548,N_6945);
nand U10852 (N_10852,N_6178,N_7871);
nor U10853 (N_10853,N_7277,N_6666);
and U10854 (N_10854,N_4270,N_5778);
or U10855 (N_10855,N_4861,N_6676);
or U10856 (N_10856,N_4952,N_7071);
and U10857 (N_10857,N_7601,N_7169);
xor U10858 (N_10858,N_7462,N_5513);
xor U10859 (N_10859,N_7489,N_5447);
nand U10860 (N_10860,N_7585,N_7869);
xnor U10861 (N_10861,N_7294,N_4009);
or U10862 (N_10862,N_5388,N_4598);
nor U10863 (N_10863,N_7221,N_7424);
nand U10864 (N_10864,N_5958,N_4286);
or U10865 (N_10865,N_4564,N_5091);
xor U10866 (N_10866,N_6365,N_6745);
or U10867 (N_10867,N_6415,N_7514);
and U10868 (N_10868,N_6431,N_6981);
xor U10869 (N_10869,N_4824,N_6745);
nor U10870 (N_10870,N_5341,N_4001);
nand U10871 (N_10871,N_5167,N_5262);
nor U10872 (N_10872,N_4989,N_7019);
xor U10873 (N_10873,N_4778,N_7203);
and U10874 (N_10874,N_7226,N_6279);
and U10875 (N_10875,N_7928,N_6682);
xnor U10876 (N_10876,N_7768,N_7493);
and U10877 (N_10877,N_5467,N_6712);
nor U10878 (N_10878,N_7036,N_4082);
or U10879 (N_10879,N_6379,N_6110);
or U10880 (N_10880,N_6596,N_6722);
nand U10881 (N_10881,N_5218,N_7704);
xor U10882 (N_10882,N_4697,N_6448);
xnor U10883 (N_10883,N_5999,N_6715);
or U10884 (N_10884,N_4342,N_6250);
and U10885 (N_10885,N_4077,N_6005);
or U10886 (N_10886,N_7293,N_4197);
xnor U10887 (N_10887,N_5865,N_7074);
xor U10888 (N_10888,N_5516,N_5466);
and U10889 (N_10889,N_6893,N_7667);
nand U10890 (N_10890,N_7142,N_6940);
and U10891 (N_10891,N_5306,N_6455);
nor U10892 (N_10892,N_4223,N_6191);
xor U10893 (N_10893,N_5615,N_5677);
or U10894 (N_10894,N_4210,N_4097);
and U10895 (N_10895,N_5395,N_5090);
or U10896 (N_10896,N_6180,N_5175);
and U10897 (N_10897,N_7209,N_7933);
and U10898 (N_10898,N_6046,N_4580);
and U10899 (N_10899,N_6288,N_4395);
xnor U10900 (N_10900,N_4164,N_7749);
xnor U10901 (N_10901,N_5097,N_4953);
nand U10902 (N_10902,N_6625,N_6064);
xnor U10903 (N_10903,N_4988,N_6988);
nand U10904 (N_10904,N_7878,N_6599);
nand U10905 (N_10905,N_5469,N_6387);
and U10906 (N_10906,N_4263,N_5609);
xor U10907 (N_10907,N_4525,N_5074);
nor U10908 (N_10908,N_5759,N_5637);
nand U10909 (N_10909,N_6106,N_7517);
and U10910 (N_10910,N_4700,N_5406);
nand U10911 (N_10911,N_4565,N_4924);
nor U10912 (N_10912,N_7103,N_7847);
xor U10913 (N_10913,N_5561,N_6634);
and U10914 (N_10914,N_4678,N_6284);
nand U10915 (N_10915,N_4267,N_5960);
xnor U10916 (N_10916,N_7604,N_7117);
nor U10917 (N_10917,N_7278,N_5156);
nor U10918 (N_10918,N_7958,N_4841);
or U10919 (N_10919,N_7008,N_6171);
nor U10920 (N_10920,N_6859,N_7787);
or U10921 (N_10921,N_6467,N_6655);
xnor U10922 (N_10922,N_5973,N_5997);
or U10923 (N_10923,N_4009,N_6435);
or U10924 (N_10924,N_6439,N_7093);
xnor U10925 (N_10925,N_7719,N_5118);
nor U10926 (N_10926,N_5621,N_7831);
nand U10927 (N_10927,N_6973,N_5342);
or U10928 (N_10928,N_7655,N_4527);
and U10929 (N_10929,N_7650,N_6795);
or U10930 (N_10930,N_5885,N_4387);
or U10931 (N_10931,N_6845,N_6136);
and U10932 (N_10932,N_4000,N_7772);
nand U10933 (N_10933,N_6601,N_5022);
nor U10934 (N_10934,N_6945,N_5476);
or U10935 (N_10935,N_4110,N_5714);
xor U10936 (N_10936,N_5327,N_6753);
nor U10937 (N_10937,N_6085,N_7881);
or U10938 (N_10938,N_6554,N_5251);
xnor U10939 (N_10939,N_5960,N_4357);
xor U10940 (N_10940,N_6399,N_7297);
nor U10941 (N_10941,N_7394,N_6241);
nand U10942 (N_10942,N_7656,N_4366);
nand U10943 (N_10943,N_7098,N_5210);
nand U10944 (N_10944,N_5053,N_4546);
nor U10945 (N_10945,N_5408,N_6990);
nor U10946 (N_10946,N_7045,N_4894);
and U10947 (N_10947,N_7503,N_5517);
nand U10948 (N_10948,N_4253,N_5229);
nor U10949 (N_10949,N_5325,N_6250);
or U10950 (N_10950,N_6467,N_5031);
nand U10951 (N_10951,N_7901,N_5408);
nand U10952 (N_10952,N_5695,N_6447);
nor U10953 (N_10953,N_7238,N_6503);
nand U10954 (N_10954,N_5801,N_7813);
nor U10955 (N_10955,N_4402,N_6559);
and U10956 (N_10956,N_4539,N_7846);
nand U10957 (N_10957,N_6095,N_5814);
nand U10958 (N_10958,N_6841,N_6905);
nand U10959 (N_10959,N_5478,N_7949);
and U10960 (N_10960,N_5459,N_6623);
nor U10961 (N_10961,N_7994,N_5448);
nand U10962 (N_10962,N_6326,N_4386);
xor U10963 (N_10963,N_4720,N_6999);
nand U10964 (N_10964,N_4651,N_6558);
nand U10965 (N_10965,N_7614,N_6896);
or U10966 (N_10966,N_5150,N_5220);
and U10967 (N_10967,N_4697,N_7406);
nor U10968 (N_10968,N_6484,N_4261);
or U10969 (N_10969,N_4593,N_4860);
nand U10970 (N_10970,N_5359,N_6889);
xor U10971 (N_10971,N_7234,N_5863);
nand U10972 (N_10972,N_7256,N_6906);
xor U10973 (N_10973,N_4814,N_6547);
nand U10974 (N_10974,N_7000,N_4635);
nor U10975 (N_10975,N_7596,N_7232);
or U10976 (N_10976,N_5563,N_5580);
and U10977 (N_10977,N_4490,N_7438);
xnor U10978 (N_10978,N_6082,N_4557);
xnor U10979 (N_10979,N_5929,N_6782);
xnor U10980 (N_10980,N_7969,N_7550);
and U10981 (N_10981,N_4075,N_5617);
and U10982 (N_10982,N_6739,N_7210);
or U10983 (N_10983,N_6089,N_7838);
nor U10984 (N_10984,N_7980,N_5295);
xor U10985 (N_10985,N_6188,N_4286);
or U10986 (N_10986,N_7104,N_4070);
nand U10987 (N_10987,N_7027,N_5270);
and U10988 (N_10988,N_4530,N_4622);
and U10989 (N_10989,N_6941,N_4071);
xnor U10990 (N_10990,N_7371,N_5925);
or U10991 (N_10991,N_6443,N_4848);
nor U10992 (N_10992,N_7887,N_7891);
nand U10993 (N_10993,N_6358,N_6553);
nand U10994 (N_10994,N_5773,N_5940);
nand U10995 (N_10995,N_6357,N_4401);
xnor U10996 (N_10996,N_4492,N_6942);
nand U10997 (N_10997,N_5346,N_5364);
nor U10998 (N_10998,N_6902,N_6066);
xor U10999 (N_10999,N_7807,N_6878);
or U11000 (N_11000,N_5899,N_4544);
nand U11001 (N_11001,N_7153,N_5244);
xor U11002 (N_11002,N_6078,N_5056);
xor U11003 (N_11003,N_7598,N_6292);
xor U11004 (N_11004,N_5798,N_5187);
and U11005 (N_11005,N_6239,N_4173);
and U11006 (N_11006,N_7659,N_4100);
nor U11007 (N_11007,N_6357,N_7149);
or U11008 (N_11008,N_6468,N_4944);
and U11009 (N_11009,N_4092,N_6505);
or U11010 (N_11010,N_4607,N_4118);
or U11011 (N_11011,N_7601,N_5176);
xor U11012 (N_11012,N_7461,N_4692);
and U11013 (N_11013,N_5698,N_4867);
nor U11014 (N_11014,N_7289,N_5936);
nor U11015 (N_11015,N_5199,N_4470);
nor U11016 (N_11016,N_4287,N_4144);
xnor U11017 (N_11017,N_5591,N_7256);
nand U11018 (N_11018,N_6282,N_7603);
xnor U11019 (N_11019,N_4534,N_5841);
nor U11020 (N_11020,N_7018,N_5049);
nand U11021 (N_11021,N_6794,N_4840);
and U11022 (N_11022,N_4818,N_6719);
nor U11023 (N_11023,N_5622,N_6741);
nor U11024 (N_11024,N_4666,N_7656);
or U11025 (N_11025,N_5696,N_5387);
nand U11026 (N_11026,N_7689,N_7656);
and U11027 (N_11027,N_5084,N_5462);
nand U11028 (N_11028,N_6578,N_5290);
and U11029 (N_11029,N_4145,N_6348);
or U11030 (N_11030,N_4120,N_7372);
or U11031 (N_11031,N_6828,N_7696);
nand U11032 (N_11032,N_7705,N_7496);
and U11033 (N_11033,N_5005,N_6836);
and U11034 (N_11034,N_5735,N_7001);
nor U11035 (N_11035,N_4538,N_6782);
nand U11036 (N_11036,N_5821,N_4763);
or U11037 (N_11037,N_6349,N_6436);
nand U11038 (N_11038,N_7881,N_5727);
nand U11039 (N_11039,N_6738,N_7768);
nor U11040 (N_11040,N_5998,N_6022);
nor U11041 (N_11041,N_7723,N_4924);
and U11042 (N_11042,N_6227,N_4530);
nand U11043 (N_11043,N_5001,N_4104);
or U11044 (N_11044,N_4128,N_7094);
or U11045 (N_11045,N_4662,N_7788);
and U11046 (N_11046,N_7965,N_5924);
xnor U11047 (N_11047,N_5561,N_7576);
or U11048 (N_11048,N_6890,N_4865);
or U11049 (N_11049,N_5802,N_4753);
nand U11050 (N_11050,N_4145,N_4163);
and U11051 (N_11051,N_7312,N_5102);
nor U11052 (N_11052,N_4312,N_7546);
or U11053 (N_11053,N_4063,N_5951);
nor U11054 (N_11054,N_4584,N_5581);
and U11055 (N_11055,N_6814,N_6301);
xor U11056 (N_11056,N_4630,N_7821);
or U11057 (N_11057,N_6360,N_4592);
or U11058 (N_11058,N_5297,N_6787);
xnor U11059 (N_11059,N_5745,N_7341);
xnor U11060 (N_11060,N_6226,N_4060);
or U11061 (N_11061,N_5840,N_7723);
xor U11062 (N_11062,N_6392,N_6768);
nor U11063 (N_11063,N_6154,N_4037);
and U11064 (N_11064,N_6994,N_6142);
and U11065 (N_11065,N_7727,N_5936);
nand U11066 (N_11066,N_4900,N_6379);
nand U11067 (N_11067,N_6122,N_7747);
xnor U11068 (N_11068,N_7457,N_7010);
and U11069 (N_11069,N_4034,N_7719);
and U11070 (N_11070,N_7465,N_5622);
xnor U11071 (N_11071,N_4374,N_4099);
nand U11072 (N_11072,N_6384,N_6564);
nand U11073 (N_11073,N_7179,N_6324);
nand U11074 (N_11074,N_6768,N_5857);
nand U11075 (N_11075,N_4395,N_7218);
nor U11076 (N_11076,N_5971,N_7421);
nor U11077 (N_11077,N_6498,N_6869);
or U11078 (N_11078,N_5358,N_4994);
and U11079 (N_11079,N_5983,N_7731);
nand U11080 (N_11080,N_5384,N_6854);
and U11081 (N_11081,N_7005,N_6212);
and U11082 (N_11082,N_4973,N_7985);
or U11083 (N_11083,N_5015,N_7909);
and U11084 (N_11084,N_4341,N_5700);
nor U11085 (N_11085,N_5239,N_4699);
nor U11086 (N_11086,N_5845,N_5162);
and U11087 (N_11087,N_7560,N_4028);
nand U11088 (N_11088,N_4585,N_6139);
xnor U11089 (N_11089,N_5632,N_7010);
nand U11090 (N_11090,N_4519,N_4891);
xnor U11091 (N_11091,N_7392,N_7240);
nor U11092 (N_11092,N_5253,N_5987);
nand U11093 (N_11093,N_7590,N_4778);
nor U11094 (N_11094,N_4137,N_7477);
nand U11095 (N_11095,N_7369,N_6696);
xnor U11096 (N_11096,N_5150,N_6631);
xnor U11097 (N_11097,N_5029,N_5459);
and U11098 (N_11098,N_5943,N_7973);
or U11099 (N_11099,N_6503,N_6931);
or U11100 (N_11100,N_5233,N_5554);
and U11101 (N_11101,N_4133,N_4559);
xnor U11102 (N_11102,N_7316,N_6532);
nor U11103 (N_11103,N_5619,N_4851);
nor U11104 (N_11104,N_5126,N_5445);
nor U11105 (N_11105,N_7031,N_5597);
nand U11106 (N_11106,N_6786,N_4222);
and U11107 (N_11107,N_6010,N_4742);
nor U11108 (N_11108,N_6266,N_5798);
nor U11109 (N_11109,N_4099,N_7905);
xor U11110 (N_11110,N_4406,N_6122);
nor U11111 (N_11111,N_7823,N_7625);
nor U11112 (N_11112,N_7043,N_5181);
nor U11113 (N_11113,N_6754,N_7492);
and U11114 (N_11114,N_6532,N_6706);
nand U11115 (N_11115,N_5741,N_5348);
xor U11116 (N_11116,N_5772,N_4998);
nand U11117 (N_11117,N_5484,N_6940);
and U11118 (N_11118,N_5095,N_6254);
nor U11119 (N_11119,N_5419,N_7022);
nor U11120 (N_11120,N_7258,N_4920);
nand U11121 (N_11121,N_5993,N_7011);
or U11122 (N_11122,N_7019,N_4437);
xor U11123 (N_11123,N_4378,N_4170);
nand U11124 (N_11124,N_7735,N_5591);
and U11125 (N_11125,N_5970,N_6430);
nand U11126 (N_11126,N_4769,N_6642);
nor U11127 (N_11127,N_7941,N_4029);
nand U11128 (N_11128,N_6284,N_6886);
nand U11129 (N_11129,N_5832,N_7435);
xnor U11130 (N_11130,N_7581,N_4828);
nor U11131 (N_11131,N_6239,N_7732);
nor U11132 (N_11132,N_5443,N_6756);
nor U11133 (N_11133,N_7530,N_5130);
or U11134 (N_11134,N_4037,N_6987);
xnor U11135 (N_11135,N_6574,N_7512);
nand U11136 (N_11136,N_5021,N_5952);
nor U11137 (N_11137,N_7459,N_7088);
nor U11138 (N_11138,N_7517,N_5977);
nor U11139 (N_11139,N_6647,N_5361);
or U11140 (N_11140,N_6691,N_5776);
nor U11141 (N_11141,N_6213,N_6081);
and U11142 (N_11142,N_4450,N_6859);
or U11143 (N_11143,N_6197,N_7721);
nand U11144 (N_11144,N_6444,N_7718);
nor U11145 (N_11145,N_7954,N_7268);
xnor U11146 (N_11146,N_5619,N_7471);
nor U11147 (N_11147,N_4087,N_7829);
and U11148 (N_11148,N_7867,N_6292);
nor U11149 (N_11149,N_4795,N_6854);
and U11150 (N_11150,N_4138,N_5055);
xnor U11151 (N_11151,N_7921,N_7670);
nand U11152 (N_11152,N_7021,N_7012);
nor U11153 (N_11153,N_7437,N_5848);
nand U11154 (N_11154,N_6838,N_4037);
xnor U11155 (N_11155,N_4783,N_5506);
and U11156 (N_11156,N_4071,N_7271);
or U11157 (N_11157,N_7098,N_5021);
nand U11158 (N_11158,N_7769,N_7062);
xor U11159 (N_11159,N_7899,N_6644);
xnor U11160 (N_11160,N_4742,N_5054);
nand U11161 (N_11161,N_5481,N_7757);
nand U11162 (N_11162,N_7249,N_5992);
nand U11163 (N_11163,N_6141,N_5280);
xnor U11164 (N_11164,N_4548,N_6141);
nor U11165 (N_11165,N_4808,N_7030);
or U11166 (N_11166,N_5560,N_4393);
or U11167 (N_11167,N_6928,N_7760);
or U11168 (N_11168,N_6517,N_5037);
or U11169 (N_11169,N_7020,N_5565);
or U11170 (N_11170,N_5942,N_4042);
nand U11171 (N_11171,N_6911,N_6149);
and U11172 (N_11172,N_6116,N_7819);
or U11173 (N_11173,N_7319,N_7187);
xor U11174 (N_11174,N_4723,N_7958);
and U11175 (N_11175,N_5259,N_5331);
or U11176 (N_11176,N_5199,N_4657);
nand U11177 (N_11177,N_4890,N_5587);
xor U11178 (N_11178,N_5300,N_4952);
or U11179 (N_11179,N_5613,N_5240);
nand U11180 (N_11180,N_7300,N_7642);
or U11181 (N_11181,N_6715,N_5209);
nand U11182 (N_11182,N_4387,N_4331);
xnor U11183 (N_11183,N_4097,N_6145);
nor U11184 (N_11184,N_6429,N_5484);
nand U11185 (N_11185,N_5164,N_5182);
and U11186 (N_11186,N_4299,N_5880);
xnor U11187 (N_11187,N_4827,N_7931);
xor U11188 (N_11188,N_7159,N_6411);
and U11189 (N_11189,N_6786,N_4177);
nand U11190 (N_11190,N_4749,N_6081);
nor U11191 (N_11191,N_4031,N_7457);
or U11192 (N_11192,N_7145,N_7481);
nor U11193 (N_11193,N_4382,N_7545);
and U11194 (N_11194,N_7709,N_5424);
xnor U11195 (N_11195,N_5455,N_6331);
nand U11196 (N_11196,N_4302,N_4696);
or U11197 (N_11197,N_6587,N_4056);
xnor U11198 (N_11198,N_4543,N_4905);
xor U11199 (N_11199,N_7436,N_5658);
or U11200 (N_11200,N_7189,N_4174);
xor U11201 (N_11201,N_4405,N_6525);
nor U11202 (N_11202,N_5453,N_6348);
or U11203 (N_11203,N_4952,N_5423);
or U11204 (N_11204,N_6200,N_4276);
nand U11205 (N_11205,N_7900,N_6751);
nand U11206 (N_11206,N_4842,N_7846);
xnor U11207 (N_11207,N_6303,N_4341);
nand U11208 (N_11208,N_6547,N_7551);
and U11209 (N_11209,N_5494,N_4486);
xor U11210 (N_11210,N_4654,N_6058);
xor U11211 (N_11211,N_4650,N_4499);
or U11212 (N_11212,N_5332,N_6011);
xnor U11213 (N_11213,N_4701,N_7213);
or U11214 (N_11214,N_7348,N_6392);
nand U11215 (N_11215,N_7371,N_6790);
xnor U11216 (N_11216,N_4710,N_5780);
and U11217 (N_11217,N_7203,N_4484);
xnor U11218 (N_11218,N_4355,N_7727);
xnor U11219 (N_11219,N_5505,N_6504);
and U11220 (N_11220,N_4151,N_7964);
nand U11221 (N_11221,N_4617,N_7706);
or U11222 (N_11222,N_7580,N_6891);
xor U11223 (N_11223,N_6004,N_7766);
nand U11224 (N_11224,N_7677,N_4927);
nor U11225 (N_11225,N_7140,N_6530);
xnor U11226 (N_11226,N_5567,N_7919);
or U11227 (N_11227,N_6700,N_5090);
nor U11228 (N_11228,N_6499,N_6326);
xor U11229 (N_11229,N_7244,N_4172);
nand U11230 (N_11230,N_4126,N_5101);
nor U11231 (N_11231,N_5436,N_7045);
and U11232 (N_11232,N_5674,N_4299);
and U11233 (N_11233,N_7692,N_7716);
nor U11234 (N_11234,N_5310,N_6941);
or U11235 (N_11235,N_6616,N_4195);
nand U11236 (N_11236,N_5440,N_6564);
nand U11237 (N_11237,N_6402,N_5142);
nor U11238 (N_11238,N_7275,N_7110);
or U11239 (N_11239,N_5383,N_4175);
nor U11240 (N_11240,N_6603,N_7794);
nand U11241 (N_11241,N_5104,N_5785);
xnor U11242 (N_11242,N_6464,N_7422);
or U11243 (N_11243,N_6774,N_6577);
xnor U11244 (N_11244,N_7568,N_5184);
xnor U11245 (N_11245,N_4692,N_6856);
or U11246 (N_11246,N_5830,N_7345);
and U11247 (N_11247,N_4595,N_7061);
nand U11248 (N_11248,N_4835,N_7950);
nand U11249 (N_11249,N_7421,N_5877);
nand U11250 (N_11250,N_6655,N_4334);
xnor U11251 (N_11251,N_7249,N_5427);
xor U11252 (N_11252,N_7141,N_6806);
nor U11253 (N_11253,N_4931,N_7276);
xor U11254 (N_11254,N_5699,N_6253);
xor U11255 (N_11255,N_4815,N_5040);
nand U11256 (N_11256,N_5342,N_6956);
nor U11257 (N_11257,N_7023,N_6426);
or U11258 (N_11258,N_7775,N_5331);
nor U11259 (N_11259,N_7115,N_5280);
nand U11260 (N_11260,N_4974,N_7618);
nor U11261 (N_11261,N_7447,N_7747);
nand U11262 (N_11262,N_7990,N_7732);
or U11263 (N_11263,N_4954,N_5989);
nand U11264 (N_11264,N_4469,N_6553);
and U11265 (N_11265,N_5466,N_6686);
xnor U11266 (N_11266,N_4961,N_4299);
xnor U11267 (N_11267,N_5509,N_4193);
nor U11268 (N_11268,N_7673,N_7068);
nor U11269 (N_11269,N_7350,N_4070);
or U11270 (N_11270,N_4784,N_4927);
or U11271 (N_11271,N_7898,N_6336);
nor U11272 (N_11272,N_4499,N_5116);
nand U11273 (N_11273,N_5761,N_6044);
nor U11274 (N_11274,N_4957,N_7065);
and U11275 (N_11275,N_6577,N_7559);
nand U11276 (N_11276,N_7816,N_6770);
xor U11277 (N_11277,N_5237,N_5783);
nor U11278 (N_11278,N_6643,N_5095);
nor U11279 (N_11279,N_7782,N_6425);
nand U11280 (N_11280,N_7915,N_6484);
nand U11281 (N_11281,N_6189,N_5668);
nand U11282 (N_11282,N_5513,N_4322);
or U11283 (N_11283,N_7603,N_5086);
nor U11284 (N_11284,N_7864,N_6959);
and U11285 (N_11285,N_5428,N_6120);
nor U11286 (N_11286,N_6153,N_5089);
and U11287 (N_11287,N_7222,N_7625);
nand U11288 (N_11288,N_6446,N_6994);
or U11289 (N_11289,N_5430,N_6792);
nand U11290 (N_11290,N_6444,N_6550);
and U11291 (N_11291,N_4983,N_7760);
or U11292 (N_11292,N_4451,N_5678);
nand U11293 (N_11293,N_7587,N_6080);
and U11294 (N_11294,N_5254,N_7007);
nor U11295 (N_11295,N_4495,N_5847);
and U11296 (N_11296,N_7544,N_4067);
nand U11297 (N_11297,N_7007,N_4341);
and U11298 (N_11298,N_4846,N_4256);
nor U11299 (N_11299,N_7830,N_4722);
and U11300 (N_11300,N_7854,N_4183);
nor U11301 (N_11301,N_6704,N_4442);
xor U11302 (N_11302,N_5683,N_4765);
nor U11303 (N_11303,N_4250,N_5459);
nor U11304 (N_11304,N_7722,N_4317);
nand U11305 (N_11305,N_5271,N_4868);
nand U11306 (N_11306,N_5823,N_6415);
xnor U11307 (N_11307,N_7388,N_4098);
and U11308 (N_11308,N_4131,N_7331);
xnor U11309 (N_11309,N_6823,N_7506);
xnor U11310 (N_11310,N_6092,N_4615);
and U11311 (N_11311,N_7741,N_5900);
and U11312 (N_11312,N_4038,N_7331);
and U11313 (N_11313,N_6812,N_4534);
xnor U11314 (N_11314,N_7160,N_6672);
or U11315 (N_11315,N_7412,N_6320);
nand U11316 (N_11316,N_5523,N_5718);
and U11317 (N_11317,N_4907,N_5223);
nor U11318 (N_11318,N_4087,N_7480);
xnor U11319 (N_11319,N_7176,N_7074);
xor U11320 (N_11320,N_6087,N_5038);
nor U11321 (N_11321,N_6806,N_6151);
nor U11322 (N_11322,N_7485,N_4398);
xor U11323 (N_11323,N_5726,N_6767);
nor U11324 (N_11324,N_5593,N_5890);
nor U11325 (N_11325,N_5356,N_6641);
or U11326 (N_11326,N_5923,N_7864);
nor U11327 (N_11327,N_6280,N_7077);
and U11328 (N_11328,N_4326,N_7201);
nand U11329 (N_11329,N_6319,N_5685);
and U11330 (N_11330,N_7328,N_6404);
nand U11331 (N_11331,N_5185,N_5545);
nor U11332 (N_11332,N_4020,N_6007);
xor U11333 (N_11333,N_5124,N_7732);
and U11334 (N_11334,N_4464,N_7827);
and U11335 (N_11335,N_5893,N_6761);
xor U11336 (N_11336,N_5740,N_7240);
or U11337 (N_11337,N_7531,N_7285);
nand U11338 (N_11338,N_5726,N_5512);
or U11339 (N_11339,N_4979,N_5632);
xor U11340 (N_11340,N_6655,N_6551);
and U11341 (N_11341,N_4386,N_5987);
xor U11342 (N_11342,N_5989,N_7083);
nor U11343 (N_11343,N_5915,N_7701);
nand U11344 (N_11344,N_4856,N_6163);
nand U11345 (N_11345,N_4064,N_5092);
nand U11346 (N_11346,N_7732,N_6561);
nand U11347 (N_11347,N_7814,N_7327);
nor U11348 (N_11348,N_4120,N_6570);
xnor U11349 (N_11349,N_7079,N_4311);
nor U11350 (N_11350,N_4085,N_7720);
or U11351 (N_11351,N_4011,N_6916);
and U11352 (N_11352,N_7833,N_5694);
and U11353 (N_11353,N_4548,N_5823);
or U11354 (N_11354,N_4979,N_6385);
nor U11355 (N_11355,N_4413,N_7072);
nor U11356 (N_11356,N_6306,N_7395);
nand U11357 (N_11357,N_6942,N_6114);
or U11358 (N_11358,N_6399,N_4876);
xnor U11359 (N_11359,N_5096,N_5900);
xor U11360 (N_11360,N_7867,N_4491);
xnor U11361 (N_11361,N_7983,N_5874);
nor U11362 (N_11362,N_7145,N_5210);
nor U11363 (N_11363,N_6880,N_7429);
xor U11364 (N_11364,N_5656,N_6363);
and U11365 (N_11365,N_6632,N_4208);
and U11366 (N_11366,N_4569,N_7427);
nor U11367 (N_11367,N_4616,N_7402);
nor U11368 (N_11368,N_4021,N_6994);
nand U11369 (N_11369,N_4913,N_4506);
and U11370 (N_11370,N_5970,N_6133);
nor U11371 (N_11371,N_7664,N_4731);
xor U11372 (N_11372,N_6699,N_5088);
and U11373 (N_11373,N_4608,N_5515);
nor U11374 (N_11374,N_5834,N_6734);
and U11375 (N_11375,N_4802,N_5417);
nand U11376 (N_11376,N_6765,N_7436);
and U11377 (N_11377,N_7331,N_4741);
nor U11378 (N_11378,N_5336,N_5489);
and U11379 (N_11379,N_7724,N_4776);
or U11380 (N_11380,N_7637,N_6375);
nand U11381 (N_11381,N_4086,N_5567);
nand U11382 (N_11382,N_6683,N_7888);
and U11383 (N_11383,N_7332,N_5658);
xnor U11384 (N_11384,N_6905,N_5891);
and U11385 (N_11385,N_4417,N_6149);
or U11386 (N_11386,N_6266,N_6818);
or U11387 (N_11387,N_6653,N_5758);
xor U11388 (N_11388,N_5046,N_7831);
or U11389 (N_11389,N_5224,N_6447);
nand U11390 (N_11390,N_6360,N_5073);
xor U11391 (N_11391,N_7954,N_4572);
or U11392 (N_11392,N_4374,N_5246);
and U11393 (N_11393,N_6442,N_7705);
nor U11394 (N_11394,N_4199,N_6363);
nor U11395 (N_11395,N_6995,N_4516);
nand U11396 (N_11396,N_4612,N_7016);
and U11397 (N_11397,N_7595,N_6319);
nand U11398 (N_11398,N_4197,N_4102);
or U11399 (N_11399,N_6343,N_6372);
xor U11400 (N_11400,N_4820,N_4399);
and U11401 (N_11401,N_5284,N_4502);
nor U11402 (N_11402,N_6384,N_7360);
or U11403 (N_11403,N_6475,N_4949);
or U11404 (N_11404,N_6307,N_6199);
xor U11405 (N_11405,N_6583,N_6972);
nand U11406 (N_11406,N_6474,N_4052);
nand U11407 (N_11407,N_4701,N_5433);
and U11408 (N_11408,N_4474,N_7363);
nand U11409 (N_11409,N_5000,N_7355);
or U11410 (N_11410,N_5992,N_5206);
or U11411 (N_11411,N_7396,N_6954);
or U11412 (N_11412,N_4826,N_7524);
xor U11413 (N_11413,N_7895,N_4276);
or U11414 (N_11414,N_7124,N_5821);
xor U11415 (N_11415,N_6443,N_4586);
nand U11416 (N_11416,N_6299,N_7507);
xor U11417 (N_11417,N_4714,N_7861);
and U11418 (N_11418,N_4313,N_7643);
xnor U11419 (N_11419,N_6276,N_4790);
nor U11420 (N_11420,N_6705,N_5301);
and U11421 (N_11421,N_6103,N_5398);
nand U11422 (N_11422,N_7965,N_5910);
xnor U11423 (N_11423,N_7669,N_6194);
xor U11424 (N_11424,N_4783,N_5524);
xor U11425 (N_11425,N_6164,N_7500);
or U11426 (N_11426,N_4727,N_6823);
or U11427 (N_11427,N_7327,N_4988);
or U11428 (N_11428,N_7490,N_5319);
or U11429 (N_11429,N_6308,N_4438);
xnor U11430 (N_11430,N_6898,N_4518);
xnor U11431 (N_11431,N_7465,N_7884);
nand U11432 (N_11432,N_6314,N_5178);
xor U11433 (N_11433,N_4445,N_7031);
nor U11434 (N_11434,N_6403,N_6151);
nand U11435 (N_11435,N_5701,N_4608);
nand U11436 (N_11436,N_7812,N_7859);
nand U11437 (N_11437,N_5252,N_5352);
or U11438 (N_11438,N_7713,N_5222);
and U11439 (N_11439,N_7002,N_6556);
nor U11440 (N_11440,N_7983,N_5971);
xnor U11441 (N_11441,N_4575,N_7381);
nand U11442 (N_11442,N_6115,N_5148);
xnor U11443 (N_11443,N_6530,N_5950);
nor U11444 (N_11444,N_6307,N_7623);
and U11445 (N_11445,N_5082,N_6683);
and U11446 (N_11446,N_4955,N_6090);
nor U11447 (N_11447,N_6814,N_7422);
nand U11448 (N_11448,N_5433,N_6158);
xnor U11449 (N_11449,N_5106,N_6192);
xnor U11450 (N_11450,N_4078,N_4927);
nand U11451 (N_11451,N_7003,N_7023);
xor U11452 (N_11452,N_6585,N_7232);
xnor U11453 (N_11453,N_7850,N_5876);
nor U11454 (N_11454,N_5490,N_4757);
nand U11455 (N_11455,N_7106,N_7350);
or U11456 (N_11456,N_4592,N_6269);
and U11457 (N_11457,N_4158,N_5180);
or U11458 (N_11458,N_7088,N_6615);
nand U11459 (N_11459,N_7026,N_5479);
nand U11460 (N_11460,N_4200,N_4374);
nor U11461 (N_11461,N_4268,N_7682);
or U11462 (N_11462,N_7877,N_4793);
xnor U11463 (N_11463,N_5971,N_7727);
xor U11464 (N_11464,N_7587,N_4410);
xor U11465 (N_11465,N_4850,N_7130);
nand U11466 (N_11466,N_5517,N_6087);
nand U11467 (N_11467,N_5146,N_4071);
xnor U11468 (N_11468,N_5048,N_4353);
and U11469 (N_11469,N_5297,N_6582);
or U11470 (N_11470,N_7004,N_5560);
nand U11471 (N_11471,N_5606,N_4990);
nor U11472 (N_11472,N_5136,N_5333);
xnor U11473 (N_11473,N_7464,N_7344);
xor U11474 (N_11474,N_7486,N_6170);
nand U11475 (N_11475,N_5656,N_5973);
nor U11476 (N_11476,N_7576,N_4523);
or U11477 (N_11477,N_6801,N_6722);
nand U11478 (N_11478,N_7514,N_5478);
xnor U11479 (N_11479,N_5934,N_7403);
nor U11480 (N_11480,N_6444,N_6173);
or U11481 (N_11481,N_4544,N_4261);
or U11482 (N_11482,N_7178,N_4545);
nor U11483 (N_11483,N_6651,N_7967);
and U11484 (N_11484,N_5076,N_5496);
nand U11485 (N_11485,N_7463,N_6651);
nand U11486 (N_11486,N_5001,N_6778);
and U11487 (N_11487,N_5117,N_7340);
nand U11488 (N_11488,N_5607,N_7591);
nand U11489 (N_11489,N_6074,N_7308);
nor U11490 (N_11490,N_5820,N_7518);
and U11491 (N_11491,N_7551,N_6165);
nand U11492 (N_11492,N_7229,N_7089);
nand U11493 (N_11493,N_5398,N_6012);
or U11494 (N_11494,N_7361,N_7359);
or U11495 (N_11495,N_7896,N_7257);
nor U11496 (N_11496,N_4304,N_5681);
nand U11497 (N_11497,N_6304,N_7264);
and U11498 (N_11498,N_5362,N_7434);
nor U11499 (N_11499,N_7518,N_4500);
nand U11500 (N_11500,N_5292,N_6956);
and U11501 (N_11501,N_6597,N_4121);
and U11502 (N_11502,N_6928,N_6444);
nor U11503 (N_11503,N_5120,N_4497);
nor U11504 (N_11504,N_7007,N_5305);
nor U11505 (N_11505,N_6562,N_4283);
nand U11506 (N_11506,N_5773,N_5373);
xnor U11507 (N_11507,N_7717,N_6813);
and U11508 (N_11508,N_7292,N_5465);
nor U11509 (N_11509,N_7744,N_7436);
and U11510 (N_11510,N_4958,N_6160);
xnor U11511 (N_11511,N_4864,N_5587);
or U11512 (N_11512,N_7599,N_6396);
xnor U11513 (N_11513,N_6676,N_4053);
or U11514 (N_11514,N_6289,N_7262);
xor U11515 (N_11515,N_5899,N_7754);
xnor U11516 (N_11516,N_4036,N_5500);
nand U11517 (N_11517,N_4712,N_7424);
nand U11518 (N_11518,N_4285,N_7942);
and U11519 (N_11519,N_7973,N_6180);
xnor U11520 (N_11520,N_7192,N_7935);
or U11521 (N_11521,N_6970,N_6375);
nand U11522 (N_11522,N_4842,N_5445);
and U11523 (N_11523,N_5037,N_4760);
and U11524 (N_11524,N_6373,N_4377);
nand U11525 (N_11525,N_4004,N_4894);
xor U11526 (N_11526,N_5847,N_4644);
and U11527 (N_11527,N_6035,N_5929);
or U11528 (N_11528,N_5852,N_4662);
xor U11529 (N_11529,N_6487,N_6042);
or U11530 (N_11530,N_5234,N_4232);
xnor U11531 (N_11531,N_6902,N_5693);
nor U11532 (N_11532,N_6666,N_4081);
and U11533 (N_11533,N_4521,N_7884);
and U11534 (N_11534,N_4290,N_7876);
xnor U11535 (N_11535,N_5601,N_7373);
nor U11536 (N_11536,N_7688,N_5106);
xnor U11537 (N_11537,N_6368,N_4694);
xnor U11538 (N_11538,N_6013,N_4761);
and U11539 (N_11539,N_6946,N_7983);
nand U11540 (N_11540,N_7103,N_5360);
nor U11541 (N_11541,N_5760,N_7421);
or U11542 (N_11542,N_7469,N_6227);
xnor U11543 (N_11543,N_7590,N_5416);
nand U11544 (N_11544,N_5876,N_5678);
nor U11545 (N_11545,N_7701,N_6926);
nor U11546 (N_11546,N_5428,N_4569);
and U11547 (N_11547,N_6709,N_6253);
and U11548 (N_11548,N_7694,N_6835);
nand U11549 (N_11549,N_5221,N_4538);
nand U11550 (N_11550,N_5428,N_6126);
and U11551 (N_11551,N_6547,N_4011);
nand U11552 (N_11552,N_7021,N_5185);
nand U11553 (N_11553,N_6331,N_6621);
nor U11554 (N_11554,N_4736,N_7476);
xnor U11555 (N_11555,N_7749,N_5067);
nand U11556 (N_11556,N_7611,N_6226);
or U11557 (N_11557,N_4195,N_4865);
xnor U11558 (N_11558,N_7865,N_6235);
or U11559 (N_11559,N_5798,N_4921);
or U11560 (N_11560,N_6552,N_5413);
xnor U11561 (N_11561,N_7417,N_4691);
nor U11562 (N_11562,N_4542,N_5959);
xor U11563 (N_11563,N_6224,N_6676);
nand U11564 (N_11564,N_4452,N_7721);
and U11565 (N_11565,N_7153,N_7617);
xnor U11566 (N_11566,N_4428,N_6916);
nand U11567 (N_11567,N_4289,N_6577);
xnor U11568 (N_11568,N_5816,N_5141);
xnor U11569 (N_11569,N_6098,N_5984);
xnor U11570 (N_11570,N_7446,N_5624);
nor U11571 (N_11571,N_6230,N_5709);
or U11572 (N_11572,N_4971,N_4122);
nor U11573 (N_11573,N_4237,N_7031);
xor U11574 (N_11574,N_4487,N_5017);
or U11575 (N_11575,N_7599,N_6536);
nand U11576 (N_11576,N_5348,N_4258);
xor U11577 (N_11577,N_4966,N_7368);
and U11578 (N_11578,N_7463,N_4625);
and U11579 (N_11579,N_6047,N_6736);
xor U11580 (N_11580,N_4727,N_7154);
or U11581 (N_11581,N_5414,N_6892);
nor U11582 (N_11582,N_5207,N_6881);
nand U11583 (N_11583,N_7527,N_6703);
and U11584 (N_11584,N_4940,N_4510);
or U11585 (N_11585,N_5879,N_7172);
xnor U11586 (N_11586,N_6897,N_5796);
nor U11587 (N_11587,N_4833,N_5198);
xnor U11588 (N_11588,N_7626,N_7402);
or U11589 (N_11589,N_7256,N_4029);
or U11590 (N_11590,N_4588,N_5686);
nor U11591 (N_11591,N_6603,N_5953);
or U11592 (N_11592,N_5699,N_7831);
nor U11593 (N_11593,N_7490,N_5796);
nand U11594 (N_11594,N_7717,N_7237);
nand U11595 (N_11595,N_4391,N_4484);
xnor U11596 (N_11596,N_7663,N_5285);
or U11597 (N_11597,N_4487,N_6239);
nor U11598 (N_11598,N_5427,N_6973);
nor U11599 (N_11599,N_4095,N_4671);
and U11600 (N_11600,N_4636,N_4398);
nor U11601 (N_11601,N_7314,N_5097);
or U11602 (N_11602,N_6861,N_4468);
xor U11603 (N_11603,N_7144,N_6316);
and U11604 (N_11604,N_7255,N_5136);
nor U11605 (N_11605,N_6171,N_6831);
nor U11606 (N_11606,N_4657,N_7347);
nor U11607 (N_11607,N_6658,N_6233);
or U11608 (N_11608,N_7773,N_5161);
and U11609 (N_11609,N_7046,N_4231);
xnor U11610 (N_11610,N_4588,N_4222);
and U11611 (N_11611,N_5443,N_7521);
or U11612 (N_11612,N_5481,N_4780);
nor U11613 (N_11613,N_6408,N_4202);
and U11614 (N_11614,N_7841,N_4413);
nor U11615 (N_11615,N_7049,N_6446);
nand U11616 (N_11616,N_6235,N_6309);
xnor U11617 (N_11617,N_4562,N_7067);
xor U11618 (N_11618,N_6830,N_6012);
nand U11619 (N_11619,N_7521,N_7032);
xnor U11620 (N_11620,N_7440,N_6461);
xnor U11621 (N_11621,N_4094,N_6809);
nor U11622 (N_11622,N_6485,N_7497);
or U11623 (N_11623,N_7478,N_4556);
or U11624 (N_11624,N_6265,N_6405);
nor U11625 (N_11625,N_4409,N_5537);
nor U11626 (N_11626,N_6363,N_5571);
nand U11627 (N_11627,N_4488,N_7331);
or U11628 (N_11628,N_7068,N_5408);
xor U11629 (N_11629,N_6307,N_6158);
or U11630 (N_11630,N_7004,N_4732);
nand U11631 (N_11631,N_4315,N_6151);
or U11632 (N_11632,N_5418,N_6933);
nor U11633 (N_11633,N_4262,N_4752);
or U11634 (N_11634,N_5664,N_6635);
or U11635 (N_11635,N_5599,N_4641);
xor U11636 (N_11636,N_7214,N_7217);
nor U11637 (N_11637,N_4051,N_5272);
xor U11638 (N_11638,N_4818,N_6905);
or U11639 (N_11639,N_4554,N_5619);
nor U11640 (N_11640,N_6708,N_7849);
and U11641 (N_11641,N_4175,N_7263);
nand U11642 (N_11642,N_5744,N_6101);
nand U11643 (N_11643,N_6791,N_4192);
xor U11644 (N_11644,N_6071,N_7828);
or U11645 (N_11645,N_5472,N_6691);
and U11646 (N_11646,N_4257,N_5042);
xnor U11647 (N_11647,N_6550,N_5237);
nor U11648 (N_11648,N_5582,N_7350);
and U11649 (N_11649,N_5749,N_4326);
or U11650 (N_11650,N_7438,N_4056);
nand U11651 (N_11651,N_6703,N_7573);
or U11652 (N_11652,N_7552,N_4936);
or U11653 (N_11653,N_4013,N_7148);
or U11654 (N_11654,N_6020,N_7214);
and U11655 (N_11655,N_4818,N_5080);
xnor U11656 (N_11656,N_6461,N_4478);
nand U11657 (N_11657,N_6379,N_7048);
nand U11658 (N_11658,N_6876,N_6545);
xnor U11659 (N_11659,N_7709,N_4217);
nor U11660 (N_11660,N_5752,N_6182);
xnor U11661 (N_11661,N_5705,N_6713);
nor U11662 (N_11662,N_4392,N_6412);
nand U11663 (N_11663,N_7163,N_7281);
or U11664 (N_11664,N_5041,N_6658);
xnor U11665 (N_11665,N_7089,N_6059);
and U11666 (N_11666,N_5952,N_6122);
xor U11667 (N_11667,N_6072,N_5439);
nand U11668 (N_11668,N_6797,N_4116);
xnor U11669 (N_11669,N_4976,N_7894);
nand U11670 (N_11670,N_7292,N_7354);
nor U11671 (N_11671,N_5589,N_4705);
and U11672 (N_11672,N_4156,N_7539);
nand U11673 (N_11673,N_4621,N_6302);
nor U11674 (N_11674,N_4466,N_4414);
or U11675 (N_11675,N_6678,N_4531);
nor U11676 (N_11676,N_7688,N_7650);
nor U11677 (N_11677,N_6867,N_6738);
and U11678 (N_11678,N_6747,N_5912);
nor U11679 (N_11679,N_4734,N_6310);
nor U11680 (N_11680,N_7678,N_4722);
nand U11681 (N_11681,N_7640,N_6778);
or U11682 (N_11682,N_4211,N_4288);
nor U11683 (N_11683,N_7059,N_4749);
nand U11684 (N_11684,N_5342,N_7211);
or U11685 (N_11685,N_4373,N_5972);
xnor U11686 (N_11686,N_5275,N_6823);
and U11687 (N_11687,N_6683,N_6695);
nand U11688 (N_11688,N_5183,N_4793);
and U11689 (N_11689,N_4063,N_4358);
or U11690 (N_11690,N_4938,N_6634);
or U11691 (N_11691,N_6037,N_5429);
xor U11692 (N_11692,N_4848,N_6884);
and U11693 (N_11693,N_4670,N_6323);
xor U11694 (N_11694,N_4408,N_5963);
nor U11695 (N_11695,N_6046,N_7785);
xor U11696 (N_11696,N_7211,N_6743);
nand U11697 (N_11697,N_6081,N_4200);
nor U11698 (N_11698,N_5550,N_4902);
or U11699 (N_11699,N_7519,N_5994);
and U11700 (N_11700,N_6825,N_4019);
or U11701 (N_11701,N_5840,N_5793);
xnor U11702 (N_11702,N_6034,N_5527);
or U11703 (N_11703,N_5438,N_6258);
nor U11704 (N_11704,N_5213,N_5558);
or U11705 (N_11705,N_4105,N_5312);
and U11706 (N_11706,N_5677,N_4580);
and U11707 (N_11707,N_4762,N_6669);
nor U11708 (N_11708,N_5212,N_5367);
xnor U11709 (N_11709,N_7928,N_7319);
and U11710 (N_11710,N_7632,N_6864);
and U11711 (N_11711,N_4190,N_4617);
xnor U11712 (N_11712,N_4347,N_4763);
or U11713 (N_11713,N_5407,N_6157);
or U11714 (N_11714,N_5530,N_6633);
or U11715 (N_11715,N_5178,N_7472);
xnor U11716 (N_11716,N_6185,N_6790);
xor U11717 (N_11717,N_6635,N_5860);
nand U11718 (N_11718,N_7256,N_7808);
or U11719 (N_11719,N_6342,N_7443);
or U11720 (N_11720,N_6529,N_5606);
nand U11721 (N_11721,N_5617,N_4236);
and U11722 (N_11722,N_6984,N_6978);
xor U11723 (N_11723,N_5268,N_5884);
xnor U11724 (N_11724,N_5383,N_6515);
nand U11725 (N_11725,N_5412,N_5815);
and U11726 (N_11726,N_6754,N_7801);
and U11727 (N_11727,N_7176,N_5554);
xnor U11728 (N_11728,N_4548,N_7238);
nand U11729 (N_11729,N_7933,N_6895);
or U11730 (N_11730,N_7046,N_7358);
or U11731 (N_11731,N_4528,N_4967);
and U11732 (N_11732,N_4848,N_5378);
nand U11733 (N_11733,N_7949,N_7329);
or U11734 (N_11734,N_6696,N_4969);
and U11735 (N_11735,N_4959,N_7275);
and U11736 (N_11736,N_5844,N_5503);
xnor U11737 (N_11737,N_7853,N_5336);
and U11738 (N_11738,N_7812,N_6346);
nand U11739 (N_11739,N_4565,N_7471);
nor U11740 (N_11740,N_6243,N_5523);
xnor U11741 (N_11741,N_5353,N_6888);
and U11742 (N_11742,N_5099,N_5032);
and U11743 (N_11743,N_5764,N_6725);
and U11744 (N_11744,N_6838,N_5757);
nor U11745 (N_11745,N_6285,N_4883);
nand U11746 (N_11746,N_5526,N_5287);
or U11747 (N_11747,N_4246,N_4712);
xnor U11748 (N_11748,N_5685,N_7600);
and U11749 (N_11749,N_5694,N_6431);
nand U11750 (N_11750,N_4752,N_7794);
xor U11751 (N_11751,N_7739,N_4232);
or U11752 (N_11752,N_7906,N_7770);
xnor U11753 (N_11753,N_5851,N_5105);
and U11754 (N_11754,N_5814,N_7898);
nand U11755 (N_11755,N_4131,N_6354);
and U11756 (N_11756,N_5722,N_6894);
nor U11757 (N_11757,N_7359,N_4758);
xnor U11758 (N_11758,N_5798,N_7960);
and U11759 (N_11759,N_5398,N_5789);
or U11760 (N_11760,N_5816,N_4716);
or U11761 (N_11761,N_4451,N_7818);
nor U11762 (N_11762,N_6270,N_6020);
nand U11763 (N_11763,N_6528,N_6630);
nor U11764 (N_11764,N_4747,N_7136);
or U11765 (N_11765,N_4498,N_6800);
xor U11766 (N_11766,N_4990,N_7434);
nor U11767 (N_11767,N_4395,N_4946);
nand U11768 (N_11768,N_5650,N_5112);
and U11769 (N_11769,N_4303,N_7278);
or U11770 (N_11770,N_5461,N_7223);
xnor U11771 (N_11771,N_5932,N_6773);
and U11772 (N_11772,N_4006,N_5258);
and U11773 (N_11773,N_5665,N_7858);
nand U11774 (N_11774,N_5397,N_5718);
xor U11775 (N_11775,N_4307,N_6357);
and U11776 (N_11776,N_7775,N_4941);
nand U11777 (N_11777,N_5915,N_7523);
and U11778 (N_11778,N_5895,N_4944);
xor U11779 (N_11779,N_5814,N_7258);
and U11780 (N_11780,N_4129,N_6159);
nor U11781 (N_11781,N_4690,N_7183);
nand U11782 (N_11782,N_5437,N_4348);
and U11783 (N_11783,N_6708,N_5328);
and U11784 (N_11784,N_7346,N_5934);
or U11785 (N_11785,N_5548,N_7158);
and U11786 (N_11786,N_4929,N_7113);
nor U11787 (N_11787,N_4365,N_5003);
nand U11788 (N_11788,N_5923,N_4369);
nor U11789 (N_11789,N_4883,N_4813);
and U11790 (N_11790,N_5321,N_6470);
nand U11791 (N_11791,N_7734,N_5417);
xor U11792 (N_11792,N_5782,N_7597);
and U11793 (N_11793,N_6914,N_7687);
nor U11794 (N_11794,N_6743,N_6036);
nand U11795 (N_11795,N_6959,N_5906);
or U11796 (N_11796,N_4042,N_4808);
nand U11797 (N_11797,N_5494,N_4517);
nand U11798 (N_11798,N_5458,N_4848);
or U11799 (N_11799,N_4984,N_7099);
and U11800 (N_11800,N_6312,N_6805);
and U11801 (N_11801,N_7492,N_4999);
nand U11802 (N_11802,N_4717,N_7089);
nor U11803 (N_11803,N_7406,N_6470);
nand U11804 (N_11804,N_5595,N_6954);
nand U11805 (N_11805,N_6470,N_6105);
nor U11806 (N_11806,N_6938,N_5854);
xnor U11807 (N_11807,N_6182,N_6603);
nand U11808 (N_11808,N_6430,N_7370);
and U11809 (N_11809,N_4303,N_7256);
and U11810 (N_11810,N_5448,N_6239);
and U11811 (N_11811,N_7645,N_5366);
nand U11812 (N_11812,N_6984,N_6699);
nand U11813 (N_11813,N_7353,N_6290);
and U11814 (N_11814,N_4215,N_5285);
nand U11815 (N_11815,N_7468,N_5738);
xor U11816 (N_11816,N_4618,N_5945);
or U11817 (N_11817,N_6297,N_6754);
nor U11818 (N_11818,N_4200,N_4877);
and U11819 (N_11819,N_5656,N_4302);
nand U11820 (N_11820,N_5405,N_4966);
nand U11821 (N_11821,N_7635,N_6362);
nand U11822 (N_11822,N_5631,N_7354);
nand U11823 (N_11823,N_7095,N_5055);
and U11824 (N_11824,N_7248,N_5850);
and U11825 (N_11825,N_7554,N_4095);
or U11826 (N_11826,N_6097,N_6101);
nand U11827 (N_11827,N_6947,N_7826);
and U11828 (N_11828,N_6157,N_5733);
nand U11829 (N_11829,N_7673,N_4330);
nor U11830 (N_11830,N_6843,N_7793);
and U11831 (N_11831,N_4398,N_4848);
and U11832 (N_11832,N_4369,N_4191);
xnor U11833 (N_11833,N_4742,N_4885);
nand U11834 (N_11834,N_7319,N_6781);
and U11835 (N_11835,N_7048,N_7773);
or U11836 (N_11836,N_5927,N_4292);
nor U11837 (N_11837,N_4639,N_7433);
and U11838 (N_11838,N_5061,N_6969);
and U11839 (N_11839,N_5741,N_5001);
xnor U11840 (N_11840,N_7506,N_5005);
or U11841 (N_11841,N_6883,N_6988);
or U11842 (N_11842,N_6276,N_5960);
nor U11843 (N_11843,N_6870,N_7917);
and U11844 (N_11844,N_4573,N_7815);
nand U11845 (N_11845,N_6376,N_6031);
nor U11846 (N_11846,N_5949,N_5632);
xor U11847 (N_11847,N_7420,N_6854);
or U11848 (N_11848,N_4217,N_6874);
nand U11849 (N_11849,N_4995,N_4569);
nor U11850 (N_11850,N_5299,N_5915);
or U11851 (N_11851,N_7205,N_6082);
or U11852 (N_11852,N_4012,N_6460);
nand U11853 (N_11853,N_6511,N_7284);
nand U11854 (N_11854,N_4980,N_4218);
and U11855 (N_11855,N_4834,N_5150);
nor U11856 (N_11856,N_7488,N_4563);
nor U11857 (N_11857,N_5143,N_5348);
or U11858 (N_11858,N_5359,N_5127);
xor U11859 (N_11859,N_6239,N_6093);
xnor U11860 (N_11860,N_5989,N_6060);
and U11861 (N_11861,N_6503,N_7536);
nand U11862 (N_11862,N_6917,N_7462);
nor U11863 (N_11863,N_5479,N_5146);
nand U11864 (N_11864,N_5517,N_6820);
nor U11865 (N_11865,N_6745,N_5324);
nand U11866 (N_11866,N_5085,N_4556);
xnor U11867 (N_11867,N_7109,N_6910);
and U11868 (N_11868,N_4452,N_7782);
nor U11869 (N_11869,N_7690,N_6004);
xnor U11870 (N_11870,N_5661,N_4194);
xnor U11871 (N_11871,N_7723,N_4485);
xor U11872 (N_11872,N_6100,N_5610);
or U11873 (N_11873,N_5937,N_6962);
xor U11874 (N_11874,N_7367,N_4651);
or U11875 (N_11875,N_6447,N_5970);
nand U11876 (N_11876,N_4360,N_7039);
or U11877 (N_11877,N_5484,N_5856);
and U11878 (N_11878,N_5303,N_6598);
xnor U11879 (N_11879,N_4268,N_6599);
xnor U11880 (N_11880,N_4058,N_7377);
or U11881 (N_11881,N_7471,N_4292);
xnor U11882 (N_11882,N_6929,N_7858);
and U11883 (N_11883,N_4876,N_4964);
or U11884 (N_11884,N_6219,N_4772);
nor U11885 (N_11885,N_7669,N_5058);
xor U11886 (N_11886,N_6057,N_6459);
nor U11887 (N_11887,N_4954,N_6637);
xnor U11888 (N_11888,N_7890,N_5158);
or U11889 (N_11889,N_7550,N_6081);
nor U11890 (N_11890,N_7048,N_6818);
nand U11891 (N_11891,N_5323,N_5163);
xnor U11892 (N_11892,N_5616,N_6737);
xnor U11893 (N_11893,N_4511,N_5369);
xor U11894 (N_11894,N_5265,N_6264);
nand U11895 (N_11895,N_4731,N_6927);
xor U11896 (N_11896,N_5162,N_7221);
xnor U11897 (N_11897,N_4894,N_6437);
and U11898 (N_11898,N_7758,N_6722);
xor U11899 (N_11899,N_4538,N_4349);
and U11900 (N_11900,N_5428,N_4299);
xor U11901 (N_11901,N_7034,N_4637);
xor U11902 (N_11902,N_6875,N_4153);
or U11903 (N_11903,N_5879,N_5000);
and U11904 (N_11904,N_5969,N_7790);
or U11905 (N_11905,N_6823,N_5552);
nor U11906 (N_11906,N_6565,N_7201);
or U11907 (N_11907,N_4177,N_5717);
nor U11908 (N_11908,N_7068,N_5624);
and U11909 (N_11909,N_7887,N_4257);
or U11910 (N_11910,N_7935,N_6934);
nor U11911 (N_11911,N_4873,N_6940);
xnor U11912 (N_11912,N_5015,N_7774);
and U11913 (N_11913,N_7323,N_7831);
nor U11914 (N_11914,N_5683,N_4975);
nand U11915 (N_11915,N_4665,N_5122);
nor U11916 (N_11916,N_5203,N_6842);
or U11917 (N_11917,N_4141,N_7902);
or U11918 (N_11918,N_4785,N_7534);
and U11919 (N_11919,N_4784,N_7292);
and U11920 (N_11920,N_6822,N_5058);
nand U11921 (N_11921,N_6383,N_5721);
or U11922 (N_11922,N_7740,N_6706);
xor U11923 (N_11923,N_5820,N_7369);
xnor U11924 (N_11924,N_6394,N_7413);
and U11925 (N_11925,N_6173,N_4134);
nor U11926 (N_11926,N_4340,N_5213);
and U11927 (N_11927,N_7308,N_5393);
nor U11928 (N_11928,N_7437,N_7434);
nor U11929 (N_11929,N_5242,N_6447);
xnor U11930 (N_11930,N_5717,N_6184);
nand U11931 (N_11931,N_4972,N_4256);
and U11932 (N_11932,N_4641,N_7778);
nor U11933 (N_11933,N_6182,N_7729);
xor U11934 (N_11934,N_4743,N_5489);
and U11935 (N_11935,N_4261,N_4357);
nor U11936 (N_11936,N_4751,N_7780);
xor U11937 (N_11937,N_4397,N_5544);
nor U11938 (N_11938,N_7023,N_5173);
nor U11939 (N_11939,N_4486,N_4506);
nand U11940 (N_11940,N_4469,N_5731);
nand U11941 (N_11941,N_7240,N_6104);
and U11942 (N_11942,N_7081,N_6467);
and U11943 (N_11943,N_5416,N_7783);
or U11944 (N_11944,N_7773,N_6062);
nand U11945 (N_11945,N_4903,N_4558);
and U11946 (N_11946,N_4162,N_7985);
and U11947 (N_11947,N_7792,N_4375);
nand U11948 (N_11948,N_7532,N_4822);
nand U11949 (N_11949,N_5593,N_6138);
or U11950 (N_11950,N_7772,N_6174);
nand U11951 (N_11951,N_4709,N_6319);
xor U11952 (N_11952,N_4925,N_6950);
and U11953 (N_11953,N_5676,N_5140);
nand U11954 (N_11954,N_6268,N_5427);
nand U11955 (N_11955,N_4327,N_6950);
or U11956 (N_11956,N_5949,N_6209);
xnor U11957 (N_11957,N_6235,N_6182);
and U11958 (N_11958,N_6693,N_7348);
or U11959 (N_11959,N_6906,N_7419);
or U11960 (N_11960,N_4487,N_7355);
xor U11961 (N_11961,N_6070,N_6383);
nand U11962 (N_11962,N_6805,N_6983);
nand U11963 (N_11963,N_4208,N_7437);
or U11964 (N_11964,N_6223,N_7718);
nor U11965 (N_11965,N_6807,N_5672);
or U11966 (N_11966,N_6041,N_4868);
or U11967 (N_11967,N_5322,N_5691);
and U11968 (N_11968,N_6295,N_6265);
xnor U11969 (N_11969,N_4005,N_7747);
xor U11970 (N_11970,N_4318,N_4553);
or U11971 (N_11971,N_4452,N_6452);
xnor U11972 (N_11972,N_4938,N_4750);
and U11973 (N_11973,N_6366,N_7347);
nor U11974 (N_11974,N_4726,N_5335);
and U11975 (N_11975,N_7793,N_7329);
nor U11976 (N_11976,N_7296,N_7319);
xnor U11977 (N_11977,N_6148,N_6096);
or U11978 (N_11978,N_6243,N_4628);
nand U11979 (N_11979,N_7999,N_7789);
or U11980 (N_11980,N_5600,N_7668);
and U11981 (N_11981,N_5762,N_4355);
nand U11982 (N_11982,N_5708,N_4333);
and U11983 (N_11983,N_6920,N_7667);
nor U11984 (N_11984,N_5696,N_6046);
xor U11985 (N_11985,N_7411,N_6009);
nor U11986 (N_11986,N_7591,N_5298);
nand U11987 (N_11987,N_5466,N_5333);
and U11988 (N_11988,N_7922,N_4740);
nor U11989 (N_11989,N_5850,N_5301);
xnor U11990 (N_11990,N_5498,N_7517);
nand U11991 (N_11991,N_4440,N_6456);
nor U11992 (N_11992,N_7681,N_6240);
xor U11993 (N_11993,N_7308,N_5204);
or U11994 (N_11994,N_6175,N_5299);
xnor U11995 (N_11995,N_6750,N_5645);
nor U11996 (N_11996,N_4974,N_4386);
or U11997 (N_11997,N_4503,N_7666);
or U11998 (N_11998,N_4035,N_7012);
nand U11999 (N_11999,N_7994,N_4081);
and U12000 (N_12000,N_9700,N_9288);
nor U12001 (N_12001,N_8576,N_10817);
nor U12002 (N_12002,N_8266,N_10371);
nor U12003 (N_12003,N_10483,N_8044);
nor U12004 (N_12004,N_9795,N_10310);
nand U12005 (N_12005,N_10760,N_8472);
nor U12006 (N_12006,N_10010,N_9245);
and U12007 (N_12007,N_8910,N_11957);
and U12008 (N_12008,N_8883,N_11497);
xnor U12009 (N_12009,N_10663,N_8520);
nand U12010 (N_12010,N_8285,N_8725);
xnor U12011 (N_12011,N_10505,N_10665);
xor U12012 (N_12012,N_8428,N_9389);
and U12013 (N_12013,N_8212,N_11103);
or U12014 (N_12014,N_9128,N_9423);
or U12015 (N_12015,N_8375,N_11825);
nand U12016 (N_12016,N_8496,N_8791);
and U12017 (N_12017,N_10195,N_8486);
nand U12018 (N_12018,N_10547,N_8696);
nand U12019 (N_12019,N_11819,N_10237);
and U12020 (N_12020,N_8831,N_9401);
nor U12021 (N_12021,N_10275,N_9167);
nand U12022 (N_12022,N_9521,N_10886);
nand U12023 (N_12023,N_9404,N_9102);
or U12024 (N_12024,N_10692,N_8835);
nand U12025 (N_12025,N_9494,N_10649);
and U12026 (N_12026,N_8545,N_8582);
and U12027 (N_12027,N_10640,N_8348);
nor U12028 (N_12028,N_8968,N_11105);
nor U12029 (N_12029,N_10900,N_8802);
nor U12030 (N_12030,N_11267,N_9991);
and U12031 (N_12031,N_11769,N_9859);
xnor U12032 (N_12032,N_9232,N_9169);
or U12033 (N_12033,N_8635,N_9522);
and U12034 (N_12034,N_11529,N_11830);
nand U12035 (N_12035,N_8389,N_9842);
and U12036 (N_12036,N_8532,N_8403);
nor U12037 (N_12037,N_10652,N_10311);
and U12038 (N_12038,N_8626,N_10482);
or U12039 (N_12039,N_9188,N_11712);
or U12040 (N_12040,N_10420,N_8634);
nand U12041 (N_12041,N_10438,N_11918);
and U12042 (N_12042,N_10851,N_10001);
nand U12043 (N_12043,N_9007,N_8652);
nor U12044 (N_12044,N_9878,N_10039);
or U12045 (N_12045,N_10688,N_11632);
nor U12046 (N_12046,N_9327,N_9472);
nor U12047 (N_12047,N_9109,N_9877);
nor U12048 (N_12048,N_8767,N_11652);
nand U12049 (N_12049,N_8839,N_8130);
nor U12050 (N_12050,N_8718,N_10631);
xnor U12051 (N_12051,N_8221,N_10047);
nand U12052 (N_12052,N_9125,N_8814);
nand U12053 (N_12053,N_10515,N_9962);
and U12054 (N_12054,N_11341,N_8892);
or U12055 (N_12055,N_10569,N_10784);
nor U12056 (N_12056,N_9014,N_11141);
nor U12057 (N_12057,N_8761,N_8733);
and U12058 (N_12058,N_8081,N_9609);
and U12059 (N_12059,N_8820,N_10374);
nand U12060 (N_12060,N_9292,N_10673);
xor U12061 (N_12061,N_10446,N_11000);
xnor U12062 (N_12062,N_9183,N_8329);
xor U12063 (N_12063,N_11506,N_10067);
or U12064 (N_12064,N_10377,N_10434);
xor U12065 (N_12065,N_10577,N_9776);
or U12066 (N_12066,N_8529,N_11390);
and U12067 (N_12067,N_9120,N_11575);
xor U12068 (N_12068,N_9174,N_11183);
nor U12069 (N_12069,N_9711,N_8257);
and U12070 (N_12070,N_10301,N_10818);
or U12071 (N_12071,N_11581,N_8919);
nand U12072 (N_12072,N_10883,N_9780);
nand U12073 (N_12073,N_9943,N_11455);
nand U12074 (N_12074,N_11223,N_8514);
or U12075 (N_12075,N_9093,N_11565);
or U12076 (N_12076,N_11944,N_10550);
and U12077 (N_12077,N_11049,N_11661);
nand U12078 (N_12078,N_11333,N_11534);
xnor U12079 (N_12079,N_9614,N_8448);
and U12080 (N_12080,N_11254,N_8141);
nand U12081 (N_12081,N_10060,N_9331);
nand U12082 (N_12082,N_8235,N_11771);
nor U12083 (N_12083,N_8322,N_8482);
or U12084 (N_12084,N_11943,N_11493);
xor U12085 (N_12085,N_11403,N_11259);
or U12086 (N_12086,N_9166,N_8539);
nand U12087 (N_12087,N_10607,N_8662);
and U12088 (N_12088,N_8692,N_11429);
xnor U12089 (N_12089,N_11278,N_11708);
nand U12090 (N_12090,N_8383,N_10308);
or U12091 (N_12091,N_11366,N_9193);
and U12092 (N_12092,N_9388,N_11723);
nor U12093 (N_12093,N_9145,N_11272);
nand U12094 (N_12094,N_9524,N_8845);
or U12095 (N_12095,N_11331,N_8060);
nor U12096 (N_12096,N_10299,N_8304);
or U12097 (N_12097,N_10270,N_8577);
nor U12098 (N_12098,N_9486,N_10812);
nand U12099 (N_12099,N_8785,N_11211);
nand U12100 (N_12100,N_9956,N_8591);
nand U12101 (N_12101,N_9872,N_11959);
nor U12102 (N_12102,N_8872,N_9335);
xnor U12103 (N_12103,N_8207,N_11874);
xor U12104 (N_12104,N_8985,N_8754);
nor U12105 (N_12105,N_9871,N_10266);
xnor U12106 (N_12106,N_8861,N_10739);
or U12107 (N_12107,N_10442,N_10257);
xnor U12108 (N_12108,N_9532,N_10525);
xnor U12109 (N_12109,N_8989,N_8700);
nand U12110 (N_12110,N_10924,N_10722);
nor U12111 (N_12111,N_8339,N_11379);
or U12112 (N_12112,N_9192,N_10633);
or U12113 (N_12113,N_9801,N_8611);
or U12114 (N_12114,N_11099,N_9605);
nand U12115 (N_12115,N_8302,N_11915);
or U12116 (N_12116,N_11227,N_11271);
or U12117 (N_12117,N_11371,N_9418);
or U12118 (N_12118,N_10976,N_10923);
and U12119 (N_12119,N_11710,N_11789);
and U12120 (N_12120,N_9505,N_11182);
xnor U12121 (N_12121,N_11679,N_8330);
or U12122 (N_12122,N_8984,N_9757);
and U12123 (N_12123,N_10381,N_11515);
xnor U12124 (N_12124,N_10020,N_8817);
nor U12125 (N_12125,N_11902,N_10655);
nor U12126 (N_12126,N_9530,N_10794);
nand U12127 (N_12127,N_8214,N_10155);
and U12128 (N_12128,N_9023,N_11650);
nand U12129 (N_12129,N_9152,N_11625);
nor U12130 (N_12130,N_10850,N_11124);
and U12131 (N_12131,N_9045,N_9274);
xor U12132 (N_12132,N_8753,N_9097);
xnor U12133 (N_12133,N_9812,N_10788);
xor U12134 (N_12134,N_8943,N_10090);
nor U12135 (N_12135,N_11420,N_8441);
nor U12136 (N_12136,N_9127,N_11243);
or U12137 (N_12137,N_11256,N_8321);
xor U12138 (N_12138,N_9493,N_8727);
and U12139 (N_12139,N_8227,N_8778);
and U12140 (N_12140,N_10548,N_9835);
nand U12141 (N_12141,N_11312,N_11042);
nand U12142 (N_12142,N_11633,N_9581);
nor U12143 (N_12143,N_8846,N_10925);
xnor U12144 (N_12144,N_11955,N_10524);
xnor U12145 (N_12145,N_9385,N_8209);
or U12146 (N_12146,N_9981,N_9623);
nor U12147 (N_12147,N_11725,N_10552);
and U12148 (N_12148,N_8877,N_10599);
or U12149 (N_12149,N_11010,N_10023);
xnor U12150 (N_12150,N_9630,N_8909);
or U12151 (N_12151,N_9194,N_9442);
xor U12152 (N_12152,N_10810,N_10680);
or U12153 (N_12153,N_8609,N_9864);
xor U12154 (N_12154,N_11500,N_8409);
xnor U12155 (N_12155,N_9387,N_11077);
nor U12156 (N_12156,N_10209,N_10297);
xor U12157 (N_12157,N_10877,N_11884);
or U12158 (N_12158,N_9363,N_10190);
and U12159 (N_12159,N_11548,N_8955);
xor U12160 (N_12160,N_11415,N_10595);
and U12161 (N_12161,N_9477,N_11871);
and U12162 (N_12162,N_11030,N_8790);
and U12163 (N_12163,N_9375,N_10054);
or U12164 (N_12164,N_10513,N_11011);
and U12165 (N_12165,N_8782,N_9811);
nand U12166 (N_12166,N_11310,N_8540);
or U12167 (N_12167,N_9879,N_10189);
nor U12168 (N_12168,N_9452,N_8586);
or U12169 (N_12169,N_9887,N_11114);
and U12170 (N_12170,N_8812,N_11121);
nor U12171 (N_12171,N_8323,N_11719);
xnor U12172 (N_12172,N_11168,N_8616);
or U12173 (N_12173,N_8109,N_10283);
or U12174 (N_12174,N_9715,N_11027);
xnor U12175 (N_12175,N_8675,N_10287);
or U12176 (N_12176,N_10026,N_11108);
or U12177 (N_12177,N_9690,N_10668);
nand U12178 (N_12178,N_11738,N_11167);
nor U12179 (N_12179,N_11586,N_11849);
nand U12180 (N_12180,N_9642,N_11537);
xor U12181 (N_12181,N_11145,N_11763);
nand U12182 (N_12182,N_10987,N_8037);
and U12183 (N_12183,N_10119,N_10272);
and U12184 (N_12184,N_11393,N_10651);
xnor U12185 (N_12185,N_8019,N_10841);
nor U12186 (N_12186,N_9203,N_9844);
nor U12187 (N_12187,N_11676,N_10022);
nand U12188 (N_12188,N_10413,N_9596);
xnor U12189 (N_12189,N_8705,N_9036);
and U12190 (N_12190,N_9511,N_8188);
and U12191 (N_12191,N_8464,N_11987);
xor U12192 (N_12192,N_9244,N_8865);
and U12193 (N_12193,N_11997,N_8874);
xor U12194 (N_12194,N_9116,N_9738);
or U12195 (N_12195,N_10499,N_10493);
nor U12196 (N_12196,N_10849,N_9090);
or U12197 (N_12197,N_10225,N_10559);
nor U12198 (N_12198,N_9393,N_11187);
or U12199 (N_12199,N_9408,N_10826);
and U12200 (N_12200,N_9399,N_11231);
xnor U12201 (N_12201,N_9555,N_8295);
nor U12202 (N_12202,N_8396,N_9115);
nand U12203 (N_12203,N_8074,N_8787);
and U12204 (N_12204,N_9638,N_8742);
nand U12205 (N_12205,N_8971,N_9495);
and U12206 (N_12206,N_8670,N_10880);
or U12207 (N_12207,N_11928,N_9114);
and U12208 (N_12208,N_11247,N_11040);
xor U12209 (N_12209,N_11948,N_9800);
and U12210 (N_12210,N_10008,N_11150);
xor U12211 (N_12211,N_8836,N_8604);
nor U12212 (N_12212,N_8837,N_10978);
or U12213 (N_12213,N_11592,N_9091);
and U12214 (N_12214,N_8864,N_10421);
nor U12215 (N_12215,N_9986,N_9656);
nor U12216 (N_12216,N_11360,N_10708);
xor U12217 (N_12217,N_11523,N_8116);
nor U12218 (N_12218,N_8058,N_10105);
and U12219 (N_12219,N_8051,N_8381);
xnor U12220 (N_12220,N_9652,N_11236);
and U12221 (N_12221,N_8771,N_10574);
nand U12222 (N_12222,N_10439,N_8365);
nand U12223 (N_12223,N_11270,N_8318);
nor U12224 (N_12224,N_8868,N_8160);
xnor U12225 (N_12225,N_10191,N_9894);
xnor U12226 (N_12226,N_10820,N_9980);
and U12227 (N_12227,N_9347,N_11604);
nand U12228 (N_12228,N_9883,N_11607);
nor U12229 (N_12229,N_8319,N_8028);
nor U12230 (N_12230,N_11845,N_9157);
nor U12231 (N_12231,N_10704,N_10306);
and U12232 (N_12232,N_9016,N_10048);
or U12233 (N_12233,N_10149,N_9682);
and U12234 (N_12234,N_11900,N_11307);
and U12235 (N_12235,N_11747,N_11917);
or U12236 (N_12236,N_11380,N_11002);
nor U12237 (N_12237,N_8101,N_11942);
nor U12238 (N_12238,N_9685,N_10435);
and U12239 (N_12239,N_8476,N_8309);
and U12240 (N_12240,N_9767,N_10447);
xnor U12241 (N_12241,N_10329,N_9163);
and U12242 (N_12242,N_10954,N_11337);
nor U12243 (N_12243,N_9551,N_10725);
nor U12244 (N_12244,N_8336,N_11752);
nand U12245 (N_12245,N_11234,N_11787);
and U12246 (N_12246,N_11125,N_10015);
or U12247 (N_12247,N_11136,N_10755);
nor U12248 (N_12248,N_8077,N_10669);
nor U12249 (N_12249,N_9606,N_11047);
nand U12250 (N_12250,N_9822,N_9969);
or U12251 (N_12251,N_10757,N_11894);
and U12252 (N_12252,N_10689,N_10252);
and U12253 (N_12253,N_9138,N_8653);
or U12254 (N_12254,N_9507,N_8848);
nand U12255 (N_12255,N_9600,N_10170);
nand U12256 (N_12256,N_8530,N_10638);
and U12257 (N_12257,N_8094,N_9316);
nand U12258 (N_12258,N_8584,N_11781);
nand U12259 (N_12259,N_9084,N_8583);
or U12260 (N_12260,N_11574,N_8988);
nand U12261 (N_12261,N_11190,N_8151);
nor U12262 (N_12262,N_10145,N_8786);
xor U12263 (N_12263,N_11153,N_10956);
nor U12264 (N_12264,N_9144,N_10215);
nor U12265 (N_12265,N_11945,N_9710);
or U12266 (N_12266,N_11767,N_8601);
nor U12267 (N_12267,N_9692,N_9197);
or U12268 (N_12268,N_11983,N_8260);
or U12269 (N_12269,N_9574,N_11981);
xor U12270 (N_12270,N_10417,N_8451);
nand U12271 (N_12271,N_10617,N_11303);
xor U12272 (N_12272,N_8363,N_11110);
nor U12273 (N_12273,N_8703,N_11930);
or U12274 (N_12274,N_11899,N_10815);
xor U12275 (N_12275,N_11806,N_10770);
xnor U12276 (N_12276,N_10713,N_8038);
nand U12277 (N_12277,N_9851,N_10071);
xor U12278 (N_12278,N_8813,N_11297);
nand U12279 (N_12279,N_9343,N_11300);
or U12280 (N_12280,N_9242,N_8970);
and U12281 (N_12281,N_10062,N_11465);
nor U12282 (N_12282,N_9467,N_9972);
xor U12283 (N_12283,N_9290,N_10608);
and U12284 (N_12284,N_9010,N_9271);
nor U12285 (N_12285,N_11573,N_11550);
and U12286 (N_12286,N_11582,N_11148);
xnor U12287 (N_12287,N_9924,N_11101);
xnor U12288 (N_12288,N_10452,N_8900);
and U12289 (N_12289,N_8983,N_9752);
xnor U12290 (N_12290,N_10829,N_10683);
nand U12291 (N_12291,N_10335,N_11605);
or U12292 (N_12292,N_9322,N_9382);
nand U12293 (N_12293,N_10902,N_11811);
nor U12294 (N_12294,N_10356,N_10120);
xnor U12295 (N_12295,N_11667,N_8738);
and U12296 (N_12296,N_9180,N_9698);
and U12297 (N_12297,N_11115,N_11513);
and U12298 (N_12298,N_10258,N_9243);
xnor U12299 (N_12299,N_8929,N_10543);
nand U12300 (N_12300,N_8132,N_9985);
nor U12301 (N_12301,N_10359,N_8867);
nand U12302 (N_12302,N_11196,N_9896);
nand U12303 (N_12303,N_10575,N_9797);
nor U12304 (N_12304,N_10063,N_10591);
nor U12305 (N_12305,N_10662,N_11893);
xor U12306 (N_12306,N_10657,N_8669);
and U12307 (N_12307,N_8268,N_9922);
or U12308 (N_12308,N_8393,N_9266);
xnor U12309 (N_12309,N_10797,N_11035);
xnor U12310 (N_12310,N_11986,N_8042);
or U12311 (N_12311,N_10744,N_10305);
xor U12312 (N_12312,N_9178,N_11502);
or U12313 (N_12313,N_11098,N_11896);
or U12314 (N_12314,N_9518,N_11599);
or U12315 (N_12315,N_8827,N_10217);
and U12316 (N_12316,N_10437,N_9182);
nor U12317 (N_12317,N_9639,N_8550);
and U12318 (N_12318,N_9989,N_9227);
and U12319 (N_12319,N_9337,N_10667);
xnor U12320 (N_12320,N_8041,N_10148);
nor U12321 (N_12321,N_8849,N_10791);
and U12322 (N_12322,N_10995,N_11804);
nand U12323 (N_12323,N_10949,N_9580);
nor U12324 (N_12324,N_9893,N_11503);
or U12325 (N_12325,N_9727,N_8800);
nor U12326 (N_12326,N_9351,N_11450);
xnor U12327 (N_12327,N_9504,N_9967);
or U12328 (N_12328,N_9542,N_8775);
xnor U12329 (N_12329,N_9264,N_8770);
xnor U12330 (N_12330,N_9817,N_9709);
and U12331 (N_12331,N_8713,N_8548);
nand U12332 (N_12332,N_10309,N_8199);
and U12333 (N_12333,N_9496,N_11364);
or U12334 (N_12334,N_10659,N_11239);
nor U12335 (N_12335,N_8695,N_9827);
nor U12336 (N_12336,N_10728,N_10496);
xor U12337 (N_12337,N_8245,N_8422);
xor U12338 (N_12338,N_9983,N_11613);
nor U12339 (N_12339,N_11144,N_8039);
or U12340 (N_12340,N_8862,N_11282);
xnor U12341 (N_12341,N_9329,N_8399);
or U12342 (N_12342,N_11316,N_8064);
nor U12343 (N_12343,N_10769,N_10616);
nand U12344 (N_12344,N_8471,N_8175);
nor U12345 (N_12345,N_10018,N_8829);
and U12346 (N_12346,N_8120,N_10862);
nor U12347 (N_12347,N_10584,N_10809);
and U12348 (N_12348,N_8842,N_9131);
nor U12349 (N_12349,N_11585,N_10402);
and U12350 (N_12350,N_10152,N_11936);
and U12351 (N_12351,N_10958,N_10520);
and U12352 (N_12352,N_11113,N_10471);
or U12353 (N_12353,N_11299,N_8522);
xor U12354 (N_12354,N_10490,N_11616);
nand U12355 (N_12355,N_8190,N_8907);
nor U12356 (N_12356,N_11219,N_11684);
and U12357 (N_12357,N_8618,N_11774);
xor U12358 (N_12358,N_11560,N_9056);
and U12359 (N_12359,N_11451,N_10619);
and U12360 (N_12360,N_8772,N_11858);
nor U12361 (N_12361,N_9763,N_8575);
or U12362 (N_12362,N_8587,N_9719);
or U12363 (N_12363,N_10064,N_8967);
and U12364 (N_12364,N_9675,N_11335);
nor U12365 (N_12365,N_11795,N_11623);
xnor U12366 (N_12366,N_10528,N_9620);
xor U12367 (N_12367,N_8431,N_8525);
nor U12368 (N_12368,N_8557,N_9468);
or U12369 (N_12369,N_11250,N_11396);
xnor U12370 (N_12370,N_11097,N_9425);
xnor U12371 (N_12371,N_9913,N_9592);
nor U12372 (N_12372,N_8882,N_11606);
nand U12373 (N_12373,N_11911,N_11185);
xnor U12374 (N_12374,N_11344,N_11966);
and U12375 (N_12375,N_10866,N_10178);
nor U12376 (N_12376,N_11290,N_9590);
nor U12377 (N_12377,N_9701,N_11904);
nand U12378 (N_12378,N_11218,N_8216);
nand U12379 (N_12379,N_10003,N_11559);
nor U12380 (N_12380,N_9736,N_8524);
or U12381 (N_12381,N_10768,N_8073);
and U12382 (N_12382,N_11547,N_11758);
nand U12383 (N_12383,N_10171,N_11742);
xor U12384 (N_12384,N_8826,N_9455);
xor U12385 (N_12385,N_9649,N_8721);
nor U12386 (N_12386,N_9315,N_8367);
nand U12387 (N_12387,N_10393,N_10321);
nor U12388 (N_12388,N_10994,N_8688);
and U12389 (N_12389,N_9750,N_9843);
and U12390 (N_12390,N_9489,N_8902);
nor U12391 (N_12391,N_10831,N_8492);
nand U12392 (N_12392,N_8405,N_8411);
and U12393 (N_12393,N_8208,N_9039);
nor U12394 (N_12394,N_11339,N_11776);
or U12395 (N_12395,N_11759,N_9965);
or U12396 (N_12396,N_10703,N_8292);
and U12397 (N_12397,N_8913,N_10967);
or U12398 (N_12398,N_8808,N_11055);
and U12399 (N_12399,N_11359,N_10984);
nor U12400 (N_12400,N_8086,N_9295);
nor U12401 (N_12401,N_9103,N_9629);
xnor U12402 (N_12402,N_9593,N_11628);
nor U12403 (N_12403,N_10121,N_8146);
xnor U12404 (N_12404,N_10615,N_10501);
or U12405 (N_12405,N_8599,N_11865);
or U12406 (N_12406,N_8340,N_8203);
xnor U12407 (N_12407,N_10303,N_10715);
xor U12408 (N_12408,N_11909,N_10772);
or U12409 (N_12409,N_10630,N_11844);
or U12410 (N_12410,N_10506,N_10202);
xnor U12411 (N_12411,N_11490,N_9995);
xnor U12412 (N_12412,N_10823,N_8716);
and U12413 (N_12413,N_10277,N_9668);
nor U12414 (N_12414,N_8608,N_10210);
nand U12415 (N_12415,N_10144,N_11260);
nor U12416 (N_12416,N_11674,N_8153);
xor U12417 (N_12417,N_11387,N_11539);
or U12418 (N_12418,N_11240,N_8498);
and U12419 (N_12419,N_9135,N_9436);
and U12420 (N_12420,N_9368,N_8597);
nor U12421 (N_12421,N_8694,N_10534);
nand U12422 (N_12422,N_10754,N_9435);
nor U12423 (N_12423,N_9526,N_9557);
nor U12424 (N_12424,N_8112,N_10491);
or U12425 (N_12425,N_10753,N_9004);
nor U12426 (N_12426,N_8751,N_8147);
and U12427 (N_12427,N_9903,N_9779);
or U12428 (N_12428,N_11139,N_8689);
nor U12429 (N_12429,N_11466,N_8654);
and U12430 (N_12430,N_10666,N_9235);
or U12431 (N_12431,N_11696,N_9523);
and U12432 (N_12432,N_9919,N_10106);
nand U12433 (N_12433,N_10636,N_10137);
and U12434 (N_12434,N_8730,N_9651);
and U12435 (N_12435,N_8225,N_9068);
xnor U12436 (N_12436,N_9134,N_9181);
and U12437 (N_12437,N_10610,N_11639);
or U12438 (N_12438,N_11249,N_8757);
nand U12439 (N_12439,N_9158,N_10096);
xnor U12440 (N_12440,N_9850,N_10750);
and U12441 (N_12441,N_8059,N_11651);
and U12442 (N_12442,N_11479,N_11274);
or U12443 (N_12443,N_11437,N_11717);
xnor U12444 (N_12444,N_9572,N_11951);
or U12445 (N_12445,N_8499,N_10674);
nand U12446 (N_12446,N_8085,N_10132);
or U12447 (N_12447,N_9305,N_9703);
nand U12448 (N_12448,N_11546,N_10672);
nand U12449 (N_12449,N_9895,N_11079);
and U12450 (N_12450,N_10223,N_11873);
xor U12451 (N_12451,N_9029,N_11089);
nor U12452 (N_12452,N_8824,N_8614);
xor U12453 (N_12453,N_9882,N_10970);
nor U12454 (N_12454,N_10360,N_10428);
nor U12455 (N_12455,N_10727,N_11238);
nor U12456 (N_12456,N_8966,N_10802);
nand U12457 (N_12457,N_10265,N_11475);
nand U12458 (N_12458,N_9326,N_11157);
or U12459 (N_12459,N_8159,N_8118);
or U12460 (N_12460,N_9793,N_11901);
nand U12461 (N_12461,N_11258,N_8815);
or U12462 (N_12462,N_8453,N_11666);
nand U12463 (N_12463,N_9549,N_10864);
or U12464 (N_12464,N_8394,N_11542);
or U12465 (N_12465,N_11705,N_11024);
nor U12466 (N_12466,N_10975,N_8495);
nand U12467 (N_12467,N_9345,N_10498);
and U12468 (N_12468,N_10024,N_10142);
xnor U12469 (N_12469,N_10783,N_9937);
and U12470 (N_12470,N_11660,N_9386);
or U12471 (N_12471,N_10611,N_8054);
or U12472 (N_12472,N_9622,N_9447);
xnor U12473 (N_12473,N_9589,N_9854);
or U12474 (N_12474,N_11469,N_10786);
and U12475 (N_12475,N_10706,N_8760);
nand U12476 (N_12476,N_8871,N_11384);
and U12477 (N_12477,N_10721,N_9766);
xor U12478 (N_12478,N_9256,N_11323);
and U12479 (N_12479,N_9976,N_10614);
nor U12480 (N_12480,N_8755,N_11749);
nor U12481 (N_12481,N_9405,N_9708);
or U12482 (N_12482,N_10656,N_11458);
nor U12483 (N_12483,N_9771,N_10541);
nor U12484 (N_12484,N_9011,N_9112);
or U12485 (N_12485,N_8707,N_11088);
xnor U12486 (N_12486,N_10028,N_10898);
or U12487 (N_12487,N_9813,N_8953);
nand U12488 (N_12488,N_11229,N_11486);
nand U12489 (N_12489,N_8274,N_10336);
and U12490 (N_12490,N_11756,N_8621);
or U12491 (N_12491,N_11378,N_11349);
and U12492 (N_12492,N_10184,N_10879);
and U12493 (N_12493,N_10077,N_8013);
xor U12494 (N_12494,N_9191,N_8043);
and U12495 (N_12495,N_8376,N_10946);
xnor U12496 (N_12496,N_9025,N_8334);
nor U12497 (N_12497,N_8513,N_9579);
nand U12498 (N_12498,N_10337,N_9664);
xor U12499 (N_12499,N_8898,N_11427);
or U12500 (N_12500,N_8969,N_10031);
nand U12501 (N_12501,N_11732,N_11212);
xor U12502 (N_12502,N_11281,N_8142);
nand U12503 (N_12503,N_10796,N_11886);
and U12504 (N_12504,N_8408,N_9753);
nor U12505 (N_12505,N_9217,N_9037);
xor U12506 (N_12506,N_8881,N_8179);
nor U12507 (N_12507,N_9647,N_9187);
and U12508 (N_12508,N_10100,N_8680);
nand U12509 (N_12509,N_9432,N_9395);
nand U12510 (N_12510,N_9540,N_11887);
nand U12511 (N_12511,N_9691,N_9100);
nor U12512 (N_12512,N_10445,N_10658);
xor U12513 (N_12513,N_8819,N_10322);
and U12514 (N_12514,N_11748,N_9765);
nor U12515 (N_12515,N_10295,N_8588);
nor U12516 (N_12516,N_10648,N_10733);
nor U12517 (N_12517,N_11956,N_9098);
or U12518 (N_12518,N_11368,N_10811);
xor U12519 (N_12519,N_11398,N_11135);
or U12520 (N_12520,N_9938,N_10718);
nand U12521 (N_12521,N_9643,N_9124);
and U12522 (N_12522,N_8645,N_9978);
xor U12523 (N_12523,N_8982,N_10370);
nor U12524 (N_12524,N_10396,N_9287);
nor U12525 (N_12525,N_10224,N_8361);
nand U12526 (N_12526,N_9428,N_11736);
or U12527 (N_12527,N_9870,N_9206);
and U12528 (N_12528,N_11257,N_10424);
nor U12529 (N_12529,N_9291,N_10418);
nor U12530 (N_12530,N_11785,N_10828);
nand U12531 (N_12531,N_11870,N_8267);
xnor U12532 (N_12532,N_11843,N_9728);
nor U12533 (N_12533,N_9360,N_10511);
and U12534 (N_12534,N_11609,N_8170);
nor U12535 (N_12535,N_8222,N_11095);
or U12536 (N_12536,N_10702,N_9755);
nor U12537 (N_12537,N_10578,N_11979);
and U12538 (N_12538,N_11799,N_11879);
and U12539 (N_12539,N_8417,N_10165);
nor U12540 (N_12540,N_9789,N_10682);
nor U12541 (N_12541,N_10992,N_10935);
nand U12542 (N_12542,N_9673,N_10176);
nor U12543 (N_12543,N_10017,N_8515);
nand U12544 (N_12544,N_11481,N_11764);
and U12545 (N_12545,N_9898,N_10572);
xnor U12546 (N_12546,N_8068,N_10212);
nor U12547 (N_12547,N_9480,N_8353);
and U12548 (N_12548,N_10123,N_11090);
xor U12549 (N_12549,N_8999,N_11025);
and U12550 (N_12550,N_8099,N_9267);
xor U12551 (N_12551,N_10670,N_8895);
nor U12552 (N_12552,N_11704,N_8371);
nor U12553 (N_12553,N_9143,N_8728);
nand U12554 (N_12554,N_11734,N_11375);
nor U12555 (N_12555,N_8182,N_11803);
nor U12556 (N_12556,N_11952,N_8676);
and U12557 (N_12557,N_9806,N_8136);
nor U12558 (N_12558,N_8928,N_9299);
nand U12559 (N_12559,N_11964,N_9044);
nand U12560 (N_12560,N_11078,N_8198);
or U12561 (N_12561,N_11060,N_9069);
nand U12562 (N_12562,N_8078,N_8241);
nor U12563 (N_12563,N_10453,N_8521);
and U12564 (N_12564,N_11087,N_10181);
and U12565 (N_12565,N_10153,N_9022);
nand U12566 (N_12566,N_11263,N_11891);
or U12567 (N_12567,N_11041,N_10825);
and U12568 (N_12568,N_10382,N_8287);
nand U12569 (N_12569,N_9324,N_10307);
nand U12570 (N_12570,N_10045,N_9311);
xor U12571 (N_12571,N_8853,N_11037);
or U12572 (N_12572,N_11831,N_11176);
nand U12573 (N_12573,N_8176,N_8445);
or U12574 (N_12574,N_8358,N_11975);
and U12575 (N_12575,N_9818,N_10516);
or U12576 (N_12576,N_8014,N_8594);
and U12577 (N_12577,N_8180,N_11394);
or U12578 (N_12578,N_10579,N_9446);
xor U12579 (N_12579,N_9807,N_9949);
or U12580 (N_12580,N_10450,N_10164);
and U12581 (N_12581,N_8400,N_10236);
or U12582 (N_12582,N_10111,N_11762);
xnor U12583 (N_12583,N_10455,N_10038);
and U12584 (N_12584,N_8140,N_10151);
and U12585 (N_12585,N_9501,N_8981);
and U12586 (N_12586,N_8878,N_11107);
nor U12587 (N_12587,N_10347,N_10238);
nor U12588 (N_12588,N_10957,N_11463);
or U12589 (N_12589,N_11841,N_8418);
nand U12590 (N_12590,N_8119,N_8466);
nand U12591 (N_12591,N_9377,N_8797);
or U12592 (N_12592,N_9908,N_9357);
nor U12593 (N_12593,N_8796,N_10332);
nand U12594 (N_12594,N_9198,N_11351);
and U12595 (N_12595,N_11483,N_11805);
or U12596 (N_12596,N_8254,N_8541);
nand U12597 (N_12597,N_8911,N_9048);
xnor U12598 (N_12598,N_11675,N_9831);
nand U12599 (N_12599,N_11611,N_8303);
nor U12600 (N_12600,N_8294,N_10005);
and U12601 (N_12601,N_11118,N_10875);
xor U12602 (N_12602,N_8229,N_10457);
or U12603 (N_12603,N_8788,N_8715);
xnor U12604 (N_12604,N_9249,N_9199);
xnor U12605 (N_12605,N_11972,N_10808);
nor U12606 (N_12606,N_9858,N_10404);
nand U12607 (N_12607,N_9019,N_11834);
or U12608 (N_12608,N_11817,N_11445);
nor U12609 (N_12609,N_11557,N_10495);
xor U12610 (N_12610,N_8185,N_10199);
or U12611 (N_12611,N_10074,N_11591);
or U12612 (N_12612,N_11596,N_10942);
xnor U12613 (N_12613,N_8997,N_9028);
and U12614 (N_12614,N_8975,N_11646);
and U12615 (N_12615,N_8595,N_10006);
nand U12616 (N_12616,N_9121,N_11851);
and U12617 (N_12617,N_10560,N_9735);
nor U12618 (N_12618,N_11988,N_10927);
nand U12619 (N_12619,N_11963,N_11718);
and U12620 (N_12620,N_11690,N_11004);
and U12621 (N_12621,N_9636,N_10486);
and U12622 (N_12622,N_8543,N_11301);
nand U12623 (N_12623,N_10571,N_9684);
nand U12624 (N_12624,N_8759,N_11677);
and U12625 (N_12625,N_10913,N_10154);
or U12626 (N_12626,N_10242,N_8901);
xnor U12627 (N_12627,N_9839,N_9954);
nor U12628 (N_12628,N_11318,N_9544);
nor U12629 (N_12629,N_11629,N_8379);
and U12630 (N_12630,N_9632,N_8017);
nor U12631 (N_12631,N_9313,N_11693);
or U12632 (N_12632,N_10863,N_10320);
nor U12633 (N_12633,N_9533,N_11104);
xnor U12634 (N_12634,N_11102,N_10546);
and U12635 (N_12635,N_11407,N_8333);
nor U12636 (N_12636,N_9886,N_10109);
xor U12637 (N_12637,N_10092,N_8327);
nand U12638 (N_12638,N_8110,N_11839);
and U12639 (N_12639,N_11698,N_8320);
nand U12640 (N_12640,N_9778,N_10107);
nand U12641 (N_12641,N_8991,N_11295);
or U12642 (N_12642,N_10385,N_9204);
nor U12643 (N_12643,N_11057,N_10333);
and U12644 (N_12644,N_9510,N_9334);
nand U12645 (N_12645,N_9814,N_8490);
nor U12646 (N_12646,N_8100,N_9852);
xor U12647 (N_12647,N_10160,N_11315);
or U12648 (N_12648,N_8995,N_9541);
and U12649 (N_12649,N_9396,N_10904);
nand U12650 (N_12650,N_8356,N_9796);
nor U12651 (N_12651,N_11823,N_9546);
nor U12652 (N_12652,N_8939,N_9402);
nor U12653 (N_12653,N_11262,N_9054);
or U12654 (N_12654,N_8506,N_10291);
and U12655 (N_12655,N_9671,N_8450);
xnor U12656 (N_12656,N_8938,N_11642);
nor U12657 (N_12657,N_8930,N_9231);
or U12658 (N_12658,N_9304,N_9672);
xnor U12659 (N_12659,N_8592,N_8380);
nor U12660 (N_12660,N_11638,N_10588);
nor U12661 (N_12661,N_11305,N_9724);
or U12662 (N_12662,N_11702,N_8818);
nor U12663 (N_12663,N_11641,N_9021);
or U12664 (N_12664,N_10403,N_10139);
and U12665 (N_12665,N_9448,N_10352);
and U12666 (N_12666,N_8007,N_11075);
xnor U12667 (N_12667,N_8841,N_10138);
nand U12668 (N_12668,N_9332,N_11489);
and U12669 (N_12669,N_9156,N_9319);
xor U12670 (N_12670,N_11554,N_8237);
xor U12671 (N_12671,N_8478,N_9861);
nor U12672 (N_12672,N_8672,N_9996);
nand U12673 (N_12673,N_10384,N_11132);
xor U12674 (N_12674,N_11369,N_9679);
xnor U12675 (N_12675,N_10081,N_10793);
xnor U12676 (N_12676,N_11399,N_11319);
nand U12677 (N_12677,N_8879,N_9699);
or U12678 (N_12678,N_10175,N_10029);
and U12679 (N_12679,N_9901,N_9035);
xor U12680 (N_12680,N_10792,N_9891);
or U12681 (N_12681,N_8963,N_11109);
and U12682 (N_12682,N_11189,N_10169);
nand U12683 (N_12683,N_9211,N_11014);
or U12684 (N_12684,N_11194,N_8364);
nor U12685 (N_12685,N_10785,N_9604);
and U12686 (N_12686,N_8480,N_10926);
or U12687 (N_12687,N_10613,N_10816);
nor U12688 (N_12688,N_9087,N_9838);
nor U12689 (N_12689,N_10763,N_9362);
and U12690 (N_12690,N_9759,N_11854);
nand U12691 (N_12691,N_8684,N_8157);
and U12692 (N_12692,N_10086,N_8507);
and U12693 (N_12693,N_9479,N_8870);
and U12694 (N_12694,N_11210,N_10530);
xnor U12695 (N_12695,N_8646,N_10351);
or U12696 (N_12696,N_11567,N_10980);
nand U12697 (N_12697,N_9429,N_9465);
or U12698 (N_12698,N_10500,N_11391);
nand U12699 (N_12699,N_8840,N_10255);
and U12700 (N_12700,N_8566,N_9856);
nor U12701 (N_12701,N_8003,N_10852);
nor U12702 (N_12702,N_11241,N_11017);
and U12703 (N_12703,N_10507,N_11919);
or U12704 (N_12704,N_10230,N_10587);
nor U12705 (N_12705,N_8942,N_9569);
nor U12706 (N_12706,N_11754,N_9619);
nor U12707 (N_12707,N_9437,N_8244);
xnor U12708 (N_12708,N_10914,N_8660);
nand U12709 (N_12709,N_11082,N_11232);
nand U12710 (N_12710,N_11877,N_9392);
and U12711 (N_12711,N_8792,N_8036);
nor U12712 (N_12712,N_9888,N_9020);
xor U12713 (N_12713,N_10625,N_9833);
and U12714 (N_12714,N_10947,N_11432);
and U12715 (N_12715,N_8378,N_8293);
or U12716 (N_12716,N_9960,N_10687);
xnor U12717 (N_12717,N_11119,N_11971);
or U12718 (N_12718,N_10734,N_8801);
or U12719 (N_12719,N_9660,N_8317);
nor U12720 (N_12720,N_11938,N_9669);
nor U12721 (N_12721,N_11400,N_11456);
and U12722 (N_12722,N_8573,N_8699);
nor U12723 (N_12723,N_11340,N_11989);
nor U12724 (N_12724,N_10477,N_11766);
xnor U12725 (N_12725,N_11084,N_9070);
or U12726 (N_12726,N_8325,N_9947);
and U12727 (N_12727,N_8986,N_8134);
or U12728 (N_12728,N_9566,N_11304);
xor U12729 (N_12729,N_10830,N_11541);
and U12730 (N_12730,N_10194,N_9519);
xor U12731 (N_12731,N_8427,N_10376);
and U12732 (N_12732,N_9265,N_11510);
nor U12733 (N_12733,N_9041,N_9052);
and U12734 (N_12734,N_9613,N_11026);
xor U12735 (N_12735,N_10628,N_8606);
or U12736 (N_12736,N_9565,N_10557);
or U12737 (N_12737,N_8816,N_8162);
and U12738 (N_12738,N_8342,N_8259);
xnor U12739 (N_12739,N_10991,N_11138);
or U12740 (N_12740,N_9380,N_11531);
and U12741 (N_12741,N_9902,N_8194);
or U12742 (N_12742,N_9676,N_11681);
and U12743 (N_12743,N_11740,N_11832);
nand U12744 (N_12744,N_9618,N_10889);
nand U12745 (N_12745,N_11786,N_11978);
nor U12746 (N_12746,N_11156,N_8264);
and U12747 (N_12747,N_8677,N_11430);
and U12748 (N_12748,N_11973,N_8226);
xor U12749 (N_12749,N_8423,N_10907);
or U12750 (N_12750,N_10399,N_8126);
or U12751 (N_12751,N_9038,N_10621);
and U12752 (N_12752,N_10315,N_9665);
nand U12753 (N_12753,N_8931,N_9200);
and U12754 (N_12754,N_9970,N_10545);
nor U12755 (N_12755,N_9516,N_9932);
xor U12756 (N_12756,N_10469,N_9161);
xor U12757 (N_12757,N_8163,N_10762);
and U12758 (N_12758,N_9439,N_11961);
or U12759 (N_12759,N_9279,N_9681);
nand U12760 (N_12760,N_8392,N_8904);
xor U12761 (N_12761,N_10627,N_11580);
xnor U12762 (N_12762,N_9648,N_9616);
nand U12763 (N_12763,N_8637,N_10917);
nor U12764 (N_12764,N_8166,N_10113);
nor U12765 (N_12765,N_9748,N_10639);
nand U12766 (N_12766,N_11248,N_10247);
and U12767 (N_12767,N_11706,N_9150);
xor U12768 (N_12768,N_10286,N_8781);
and U12769 (N_12769,N_9006,N_10853);
or U12770 (N_12770,N_9775,N_10700);
nand U12771 (N_12771,N_11610,N_10228);
nor U12772 (N_12772,N_9064,N_9223);
nand U12773 (N_12773,N_11790,N_10243);
xor U12774 (N_12774,N_10033,N_9430);
nor U12775 (N_12775,N_11169,N_10861);
xnor U12776 (N_12776,N_11205,N_11730);
nand U12777 (N_12777,N_9463,N_9086);
xor U12778 (N_12778,N_10943,N_9587);
xnor U12779 (N_12779,N_8996,N_9270);
xor U12780 (N_12780,N_10590,N_10362);
nand U12781 (N_12781,N_8069,N_8855);
and U12782 (N_12782,N_8647,N_8242);
nor U12783 (N_12783,N_11598,N_9189);
and U12784 (N_12784,N_10323,N_8769);
nand U12785 (N_12785,N_9973,N_11204);
or U12786 (N_12786,N_10521,N_9979);
xnor U12787 (N_12787,N_9234,N_9101);
nand U12788 (N_12788,N_8914,N_8178);
xor U12789 (N_12789,N_8620,N_9296);
or U12790 (N_12790,N_10245,N_11329);
nor U12791 (N_12791,N_8958,N_10531);
xor U12792 (N_12792,N_8823,N_8745);
nor U12793 (N_12793,N_9670,N_11492);
and U12794 (N_12794,N_8040,N_8799);
or U12795 (N_12795,N_8925,N_9015);
or U12796 (N_12796,N_10554,N_11411);
nor U12797 (N_12797,N_11967,N_9998);
or U12798 (N_12798,N_10431,N_11644);
or U12799 (N_12799,N_11233,N_8731);
and U12800 (N_12800,N_9365,N_11538);
nor U12801 (N_12801,N_10671,N_9900);
or U12802 (N_12802,N_8947,N_8402);
and U12803 (N_12803,N_8962,N_11452);
nand U12804 (N_12804,N_9214,N_8076);
and U12805 (N_12805,N_10114,N_8031);
xnor U12806 (N_12806,N_8297,N_8806);
nor U12807 (N_12807,N_10200,N_9769);
xor U12808 (N_12808,N_10989,N_10971);
nand U12809 (N_12809,N_11074,N_11768);
and U12810 (N_12810,N_9081,N_9939);
nor U12811 (N_12811,N_10776,N_8131);
and U12812 (N_12812,N_8300,N_8449);
and U12813 (N_12813,N_11755,N_8174);
nand U12814 (N_12814,N_10765,N_8127);
and U12815 (N_12815,N_11783,N_8406);
xor U12816 (N_12816,N_11470,N_10677);
xnor U12817 (N_12817,N_9828,N_10839);
or U12818 (N_12818,N_10800,N_10016);
nor U12819 (N_12819,N_8612,N_8204);
and U12820 (N_12820,N_11418,N_8171);
xnor U12821 (N_12821,N_8534,N_8215);
xor U12822 (N_12822,N_8169,N_10562);
and U12823 (N_12823,N_9403,N_9586);
nor U12824 (N_12824,N_11881,N_9904);
nand U12825 (N_12825,N_11720,N_8474);
nor U12826 (N_12826,N_9419,N_10182);
xnor U12827 (N_12827,N_10585,N_11005);
xor U12828 (N_12828,N_9050,N_10888);
or U12829 (N_12829,N_8385,N_9043);
xor U12830 (N_12830,N_8628,N_10643);
xnor U12831 (N_12831,N_8272,N_9534);
nor U12832 (N_12832,N_10146,N_8535);
and U12833 (N_12833,N_9737,N_11111);
nor U12834 (N_12834,N_10468,N_9030);
xnor U12835 (N_12835,N_8505,N_10833);
nand U12836 (N_12836,N_10881,N_11289);
xnor U12837 (N_12837,N_8331,N_10542);
and U12838 (N_12838,N_10514,N_10405);
and U12839 (N_12839,N_8066,N_11922);
nor U12840 (N_12840,N_11434,N_11965);
nor U12841 (N_12841,N_8168,N_11094);
xnor U12842 (N_12842,N_11921,N_8641);
or U12843 (N_12843,N_10475,N_11226);
and U12844 (N_12844,N_9367,N_11414);
xnor U12845 (N_12845,N_10098,N_8291);
nor U12846 (N_12846,N_11657,N_9009);
and U12847 (N_12847,N_9341,N_9469);
nand U12848 (N_12848,N_9889,N_8489);
or U12849 (N_12849,N_9603,N_10964);
and U12850 (N_12850,N_9230,N_11563);
nor U12851 (N_12851,N_10805,N_11746);
xnor U12852 (N_12852,N_9094,N_10398);
nor U12853 (N_12853,N_11269,N_11220);
or U12854 (N_12854,N_10279,N_10379);
nand U12855 (N_12855,N_10932,N_10462);
nor U12856 (N_12856,N_9957,N_10522);
xor U12857 (N_12857,N_8992,N_11009);
and U12858 (N_12858,N_9342,N_11330);
and U12859 (N_12859,N_8282,N_11086);
and U12860 (N_12860,N_9712,N_10085);
nor U12861 (N_12861,N_9293,N_8678);
and U12862 (N_12862,N_9697,N_10593);
nor U12863 (N_12863,N_10179,N_8223);
or U12864 (N_12864,N_10941,N_10460);
nand U12865 (N_12865,N_10642,N_9751);
and U12866 (N_12866,N_8789,N_9352);
xnor U12867 (N_12867,N_8565,N_9865);
nor U12868 (N_12868,N_9963,N_8298);
and U12869 (N_12869,N_10934,N_8714);
xor U12870 (N_12870,N_10216,N_8553);
and U12871 (N_12871,N_10289,N_8860);
nor U12872 (N_12872,N_11691,N_11927);
and U12873 (N_12873,N_11480,N_9720);
or U12874 (N_12874,N_10316,N_9866);
nand U12875 (N_12875,N_8465,N_10884);
nor U12876 (N_12876,N_8828,N_11031);
or U12877 (N_12877,N_9742,N_10489);
and U12878 (N_12878,N_8629,N_10174);
or U12879 (N_12879,N_11869,N_8564);
nand U12880 (N_12880,N_10869,N_11777);
xnor U12881 (N_12881,N_11334,N_8915);
nand U12882 (N_12882,N_8552,N_10448);
nor U12883 (N_12883,N_11727,N_11404);
nor U12884 (N_12884,N_10535,N_10618);
or U12885 (N_12885,N_11439,N_8916);
and U12886 (N_12886,N_10596,N_10361);
nor U12887 (N_12887,N_8708,N_10695);
nor U12888 (N_12888,N_8687,N_10425);
nand U12889 (N_12889,N_11525,N_10842);
nand U12890 (N_12890,N_10441,N_11286);
nor U12891 (N_12891,N_11350,N_9340);
and U12892 (N_12892,N_11630,N_10084);
xnor U12893 (N_12893,N_10766,N_11589);
nand U12894 (N_12894,N_10748,N_8726);
nor U12895 (N_12895,N_10632,N_9575);
nand U12896 (N_12896,N_8686,N_11590);
nor U12897 (N_12897,N_8516,N_9547);
nor U12898 (N_12898,N_9431,N_11279);
or U12899 (N_12899,N_10180,N_11615);
nor U12900 (N_12900,N_11903,N_8243);
xor U12901 (N_12901,N_8350,N_9845);
xnor U12902 (N_12902,N_9645,N_11744);
and U12903 (N_12903,N_8349,N_11687);
or U12904 (N_12904,N_11348,N_10478);
and U12905 (N_12905,N_9984,N_8519);
xnor U12906 (N_12906,N_9602,N_10916);
nand U12907 (N_12907,N_8404,N_8783);
nor U12908 (N_12908,N_10600,N_9303);
and U12909 (N_12909,N_8856,N_8590);
nor U12910 (N_12910,N_11409,N_11362);
or U12911 (N_12911,N_10999,N_9545);
nor U12912 (N_12912,N_9426,N_11096);
nand U12913 (N_12913,N_8424,N_9168);
or U12914 (N_12914,N_9280,N_9246);
nand U12915 (N_12915,N_9819,N_11253);
and U12916 (N_12916,N_8702,N_11837);
nor U12917 (N_12917,N_11029,N_11916);
nand U12918 (N_12918,N_8585,N_11228);
xnor U12919 (N_12919,N_8055,N_10340);
or U12920 (N_12920,N_9250,N_11284);
or U12921 (N_12921,N_11061,N_10366);
xor U12922 (N_12922,N_8657,N_10101);
nand U12923 (N_12923,N_10188,N_9594);
nand U12924 (N_12924,N_11052,N_10130);
nor U12925 (N_12925,N_9172,N_11937);
or U12926 (N_12926,N_8337,N_8310);
nor U12927 (N_12927,N_11587,N_8373);
nor U12928 (N_12928,N_8281,N_10040);
and U12929 (N_12929,N_10032,N_10664);
nor U12930 (N_12930,N_8301,N_9873);
nand U12931 (N_12931,N_8355,N_9353);
and U12932 (N_12932,N_11686,N_9107);
xnor U12933 (N_12933,N_8388,N_10124);
or U12934 (N_12934,N_9348,N_10167);
xor U12935 (N_12935,N_11015,N_8523);
nand U12936 (N_12936,N_9359,N_8477);
nor U12937 (N_12937,N_9968,N_11527);
nand U12938 (N_12938,N_8903,N_9987);
nand U12939 (N_12939,N_11812,N_11931);
and U12940 (N_12940,N_10394,N_11509);
nand U12941 (N_12941,N_10313,N_9237);
xnor U12942 (N_12942,N_10426,N_8978);
nand U12943 (N_12943,N_9553,N_11645);
and U12944 (N_12944,N_11522,N_10235);
nor U12945 (N_12945,N_9731,N_9941);
nand U12946 (N_12946,N_10523,N_8213);
nor U12947 (N_12947,N_10341,N_10948);
nor U12948 (N_12948,N_9027,N_11435);
nand U12949 (N_12949,N_8186,N_8261);
nand U12950 (N_12950,N_11022,N_9809);
nand U12951 (N_12951,N_10961,N_10566);
or U12952 (N_12952,N_10601,N_8603);
or U12953 (N_12953,N_8006,N_10273);
or U12954 (N_12954,N_8998,N_11365);
xor U12955 (N_12955,N_9820,N_10367);
nor U12956 (N_12956,N_9723,N_10711);
and U12957 (N_12957,N_11791,N_8458);
or U12958 (N_12958,N_10835,N_10896);
or U12959 (N_12959,N_10647,N_10726);
or U12960 (N_12960,N_11244,N_11142);
or U12961 (N_12961,N_9747,N_9663);
nor U12962 (N_12962,N_10944,N_10248);
and U12963 (N_12963,N_8275,N_8843);
or U12964 (N_12964,N_9907,N_9034);
xor U12965 (N_12965,N_10752,N_11314);
nor U12966 (N_12966,N_10774,N_11940);
xor U12967 (N_12967,N_8335,N_11083);
and U12968 (N_12968,N_11039,N_9096);
xnor U12969 (N_12969,N_10686,N_8650);
or U12970 (N_12970,N_11354,N_11080);
or U12971 (N_12971,N_11703,N_10091);
and U12972 (N_12972,N_9456,N_9307);
nor U12973 (N_12973,N_11558,N_11472);
or U12974 (N_12974,N_11495,N_9407);
nor U12975 (N_12975,N_9252,N_10264);
xor U12976 (N_12976,N_11291,N_10122);
nand U12977 (N_12977,N_8625,N_11143);
nor U12978 (N_12978,N_9358,N_9608);
xor U12979 (N_12979,N_11857,N_10246);
and U12980 (N_12980,N_9219,N_9869);
nor U12981 (N_12981,N_9626,N_10716);
xor U12982 (N_12982,N_11302,N_11324);
or U12983 (N_12983,N_10848,N_10056);
and U12984 (N_12984,N_9445,N_11753);
nor U12985 (N_12985,N_9159,N_9926);
nor U12986 (N_12986,N_11864,N_8426);
nor U12987 (N_12987,N_11714,N_11161);
xnor U12988 (N_12988,N_8344,N_9931);
and U12989 (N_12989,N_8944,N_10267);
nor U12990 (N_12990,N_10931,N_11117);
xnor U12991 (N_12991,N_9119,N_8063);
or U12992 (N_12992,N_8844,N_11346);
nand U12993 (N_12993,N_8290,N_11892);
nor U12994 (N_12994,N_11050,N_10973);
xnor U12995 (N_12995,N_8279,N_9786);
xor U12996 (N_12996,N_10058,N_10872);
and U12997 (N_12997,N_10919,N_10789);
and U12998 (N_12998,N_11172,N_11386);
nand U12999 (N_12999,N_10782,N_9912);
xnor U13000 (N_13000,N_11353,N_11171);
nand U13001 (N_13001,N_11820,N_10922);
and U13002 (N_13002,N_10485,N_10890);
xor U13003 (N_13003,N_9226,N_8205);
or U13004 (N_13004,N_11685,N_10082);
xor U13005 (N_13005,N_9890,N_8108);
nand U13006 (N_13006,N_10249,N_8830);
xnor U13007 (N_13007,N_11536,N_10391);
xnor U13008 (N_13008,N_10294,N_10538);
nand U13009 (N_13009,N_11508,N_8663);
xnor U13010 (N_13010,N_8822,N_8167);
or U13011 (N_13011,N_9040,N_11653);
nor U13012 (N_13012,N_10894,N_8369);
nand U13013 (N_13013,N_9104,N_11793);
nand U13014 (N_13014,N_10865,N_11835);
nand U13015 (N_13015,N_8030,N_10099);
and U13016 (N_13016,N_8993,N_11370);
nand U13017 (N_13017,N_8352,N_8952);
and U13018 (N_13018,N_9584,N_10945);
and U13019 (N_13019,N_9884,N_9803);
nand U13020 (N_13020,N_8581,N_11162);
or U13021 (N_13021,N_9933,N_8664);
nor U13022 (N_13022,N_11828,N_9153);
xnor U13023 (N_13023,N_8253,N_9961);
nand U13024 (N_13024,N_11484,N_10795);
or U13025 (N_13025,N_9646,N_10186);
xor U13026 (N_13026,N_9583,N_9722);
and U13027 (N_13027,N_11556,N_11517);
and U13028 (N_13028,N_8276,N_11612);
xnor U13029 (N_13029,N_9461,N_11342);
nand U13030 (N_13030,N_10979,N_9982);
or U13031 (N_13031,N_9971,N_10626);
and U13032 (N_13032,N_11397,N_8661);
or U13033 (N_13033,N_11895,N_10564);
nand U13034 (N_13034,N_8117,N_10602);
xnor U13035 (N_13035,N_9782,N_9881);
nor U13036 (N_13036,N_8129,N_8395);
or U13037 (N_13037,N_9003,N_8386);
nor U13038 (N_13038,N_10211,N_11198);
nand U13039 (N_13039,N_10043,N_9925);
and U13040 (N_13040,N_10847,N_11276);
and U13041 (N_13041,N_8920,N_8908);
and U13042 (N_13042,N_8712,N_11252);
nand U13043 (N_13043,N_8197,N_8270);
or U13044 (N_13044,N_11180,N_10814);
xor U13045 (N_13045,N_8559,N_11519);
or U13046 (N_13046,N_8430,N_8346);
or U13047 (N_13047,N_9424,N_9730);
and U13048 (N_13048,N_11514,N_10088);
or U13049 (N_13049,N_11137,N_10968);
nor U13050 (N_13050,N_8161,N_9218);
or U13051 (N_13051,N_11631,N_10549);
and U13052 (N_13052,N_8533,N_9123);
and U13053 (N_13053,N_11028,N_10963);
or U13054 (N_13054,N_11780,N_9275);
nand U13055 (N_13055,N_11471,N_10936);
nor U13056 (N_13056,N_9741,N_10871);
and U13057 (N_13057,N_10583,N_9470);
nor U13058 (N_13058,N_8184,N_8137);
nand U13059 (N_13059,N_8527,N_9175);
nor U13060 (N_13060,N_8082,N_10540);
nand U13061 (N_13061,N_10363,N_11946);
xnor U13062 (N_13062,N_11863,N_10203);
nand U13063 (N_13063,N_8265,N_9239);
or U13064 (N_13064,N_9849,N_9857);
xor U13065 (N_13065,N_10343,N_9777);
and U13066 (N_13066,N_9474,N_8021);
and U13067 (N_13067,N_11328,N_9958);
nand U13068 (N_13068,N_9661,N_8936);
or U13069 (N_13069,N_9862,N_10720);
nor U13070 (N_13070,N_9659,N_8758);
nand U13071 (N_13071,N_11699,N_11555);
nor U13072 (N_13072,N_8062,N_11417);
nand U13073 (N_13073,N_11802,N_11925);
nand U13074 (N_13074,N_8236,N_8894);
or U13075 (N_13075,N_11032,N_10002);
xor U13076 (N_13076,N_11163,N_8542);
nand U13077 (N_13077,N_11374,N_9815);
or U13078 (N_13078,N_9761,N_8632);
or U13079 (N_13079,N_11772,N_8284);
or U13080 (N_13080,N_10368,N_9298);
nor U13081 (N_13081,N_9935,N_10836);
and U13082 (N_13082,N_10536,N_8596);
or U13083 (N_13083,N_9847,N_8387);
xnor U13084 (N_13084,N_9787,N_8196);
or U13085 (N_13085,N_11827,N_11980);
nand U13086 (N_13086,N_8976,N_11838);
or U13087 (N_13087,N_11552,N_9610);
nand U13088 (N_13088,N_11292,N_11692);
and U13089 (N_13089,N_9837,N_11130);
xnor U13090 (N_13090,N_10073,N_8651);
or U13091 (N_13091,N_8918,N_10960);
and U13092 (N_13092,N_8324,N_9992);
xor U13093 (N_13093,N_10827,N_10253);
xnor U13094 (N_13094,N_10027,N_9768);
or U13095 (N_13095,N_11697,N_8278);
nand U13096 (N_13096,N_10690,N_9413);
nand U13097 (N_13097,N_9571,N_9483);
or U13098 (N_13098,N_9476,N_11859);
nor U13099 (N_13099,N_8766,N_11990);
and U13100 (N_13100,N_9110,N_8602);
xnor U13101 (N_13101,N_8067,N_10977);
and U13102 (N_13102,N_8809,N_8691);
xor U13103 (N_13103,N_11571,N_10832);
or U13104 (N_13104,N_10679,N_11127);
or U13105 (N_13105,N_11949,N_9988);
xor U13106 (N_13106,N_11408,N_10288);
nor U13107 (N_13107,N_10474,N_10806);
nand U13108 (N_13108,N_10895,N_10241);
xor U13109 (N_13109,N_8479,N_10969);
nor U13110 (N_13110,N_9770,N_11416);
or U13111 (N_13111,N_8050,N_10076);
nor U13112 (N_13112,N_11441,N_11707);
or U13113 (N_13113,N_11440,N_11505);
xnor U13114 (N_13114,N_8232,N_8048);
and U13115 (N_13115,N_10773,N_11543);
xnor U13116 (N_13116,N_9032,N_8457);
nor U13117 (N_13117,N_10078,N_8217);
or U13118 (N_13118,N_8027,N_11073);
nor U13119 (N_13119,N_11012,N_9233);
or U13120 (N_13120,N_11745,N_10208);
nand U13121 (N_13121,N_9918,N_10623);
nand U13122 (N_13122,N_9099,N_8219);
or U13123 (N_13123,N_9240,N_8834);
xor U13124 (N_13124,N_8610,N_8191);
and U13125 (N_13125,N_10380,N_11149);
nor U13126 (N_13126,N_9209,N_10419);
or U13127 (N_13127,N_11897,N_8810);
and U13128 (N_13128,N_11860,N_8884);
xnor U13129 (N_13129,N_10386,N_8090);
or U13130 (N_13130,N_9306,N_8328);
nand U13131 (N_13131,N_10854,N_8391);
nor U13132 (N_13132,N_8231,N_10057);
nor U13133 (N_13133,N_8876,N_10637);
nand U13134 (N_13134,N_10492,N_10915);
nand U13135 (N_13135,N_11929,N_9829);
xnor U13136 (N_13136,N_11672,N_11761);
nor U13137 (N_13137,N_9576,N_11512);
and U13138 (N_13138,N_9830,N_8667);
xnor U13139 (N_13139,N_11801,N_8412);
or U13140 (N_13140,N_11268,N_11602);
xnor U13141 (N_13141,N_10939,N_11833);
xnor U13142 (N_13142,N_8459,N_8026);
xor U13143 (N_13143,N_10196,N_10068);
nand U13144 (N_13144,N_11683,N_9310);
xnor U13145 (N_13145,N_11165,N_11357);
xnor U13146 (N_13146,N_11577,N_9876);
or U13147 (N_13147,N_9077,N_10244);
nor U13148 (N_13148,N_8390,N_11499);
nand U13149 (N_13149,N_8917,N_9667);
nand U13150 (N_13150,N_8922,N_9974);
and U13151 (N_13151,N_10214,N_8624);
nand U13152 (N_13152,N_9840,N_10346);
or U13153 (N_13153,N_10344,N_8311);
xnor U13154 (N_13154,N_10476,N_10738);
and U13155 (N_13155,N_11716,N_8128);
xnor U13156 (N_13156,N_11361,N_8434);
or U13157 (N_13157,N_8469,N_10580);
and U13158 (N_13158,N_10193,N_8092);
or U13159 (N_13159,N_9354,N_10644);
nand U13160 (N_13160,N_9141,N_9500);
nand U13161 (N_13161,N_10037,N_9049);
nand U13162 (N_13162,N_10375,N_8893);
xnor U13163 (N_13163,N_8659,N_10759);
xnor U13164 (N_13164,N_9412,N_11280);
xor U13165 (N_13165,N_10510,N_9598);
or U13166 (N_13166,N_9492,N_11023);
nor U13167 (N_13167,N_8343,N_11784);
or U13168 (N_13168,N_11584,N_10390);
xnor U13169 (N_13169,N_10897,N_10529);
or U13170 (N_13170,N_8382,N_10532);
nand U13171 (N_13171,N_9248,N_8719);
nor U13172 (N_13172,N_9460,N_11197);
nand U13173 (N_13173,N_11847,N_10276);
xnor U13174 (N_13174,N_10296,N_10254);
nor U13175 (N_13175,N_10061,N_10251);
or U13176 (N_13176,N_9946,N_11794);
and U13177 (N_13177,N_10484,N_10719);
nor U13178 (N_13178,N_11283,N_11528);
and U13179 (N_13179,N_10444,N_8072);
or U13180 (N_13180,N_10192,N_9105);
or U13181 (N_13181,N_11654,N_11737);
xor U13182 (N_13182,N_10260,N_10775);
or U13183 (N_13183,N_9176,N_9595);
or U13184 (N_13184,N_9564,N_11982);
or U13185 (N_13185,N_8454,N_10533);
or U13186 (N_13186,N_10781,N_8737);
nand U13187 (N_13187,N_9772,N_10928);
and U13188 (N_13188,N_11852,N_9260);
nand U13189 (N_13189,N_8681,N_10955);
and U13190 (N_13190,N_9001,N_9687);
and U13191 (N_13191,N_9808,N_8537);
and U13192 (N_13192,N_11235,N_8935);
and U13193 (N_13193,N_8446,N_8674);
nor U13194 (N_13194,N_9805,N_11775);
or U13195 (N_13195,N_8948,N_11072);
xnor U13196 (N_13196,N_10606,N_9289);
or U13197 (N_13197,N_11540,N_10870);
and U13198 (N_13198,N_10449,N_9585);
xor U13199 (N_13199,N_8921,N_10059);
nor U13200 (N_13200,N_8102,N_10729);
xor U13201 (N_13201,N_10758,N_10229);
xor U13202 (N_13202,N_9002,N_10609);
nand U13203 (N_13203,N_10166,N_11861);
xor U13204 (N_13204,N_11343,N_11689);
and U13205 (N_13205,N_9662,N_11482);
nor U13206 (N_13206,N_9863,N_9031);
xnor U13207 (N_13207,N_9253,N_9959);
nand U13208 (N_13208,N_8517,N_8673);
nor U13209 (N_13209,N_9411,N_10983);
xnor U13210 (N_13210,N_11824,N_9080);
and U13211 (N_13211,N_11154,N_10933);
or U13212 (N_13212,N_10036,N_11170);
and U13213 (N_13213,N_11207,N_9350);
xnor U13214 (N_13214,N_9860,N_10089);
and U13215 (N_13215,N_9294,N_9707);
nand U13216 (N_13216,N_8238,N_8113);
xnor U13217 (N_13217,N_8794,N_11298);
xor U13218 (N_13218,N_9760,N_8493);
or U13219 (N_13219,N_10044,N_10678);
or U13220 (N_13220,N_10876,N_11619);
and U13221 (N_13221,N_11665,N_11671);
nor U13222 (N_13222,N_9846,N_10813);
xor U13223 (N_13223,N_11213,N_8589);
nor U13224 (N_13224,N_10908,N_9207);
or U13225 (N_13225,N_8526,N_8671);
or U13226 (N_13226,N_10117,N_8071);
nand U13227 (N_13227,N_9376,N_8957);
xor U13228 (N_13228,N_11020,N_10378);
nor U13229 (N_13229,N_9302,N_11395);
or U13230 (N_13230,N_11561,N_11066);
nand U13231 (N_13231,N_9443,N_9517);
and U13232 (N_13232,N_9537,N_8251);
nor U13233 (N_13233,N_9126,N_10075);
xor U13234 (N_13234,N_9880,N_10746);
nand U13235 (N_13235,N_10087,N_10997);
nor U13236 (N_13236,N_8924,N_9222);
nor U13237 (N_13237,N_8481,N_9255);
nor U13238 (N_13238,N_11070,N_9936);
nand U13239 (N_13239,N_10654,N_9826);
or U13240 (N_13240,N_8444,N_8210);
or U13241 (N_13241,N_9251,N_11321);
or U13242 (N_13242,N_11152,N_8308);
and U13243 (N_13243,N_9548,N_10707);
or U13244 (N_13244,N_11193,N_9398);
nand U13245 (N_13245,N_9210,N_8397);
nand U13246 (N_13246,N_8022,N_8563);
nand U13247 (N_13247,N_10331,N_8262);
nor U13248 (N_13248,N_10221,N_10589);
xnor U13249 (N_13249,N_8648,N_10051);
nand U13250 (N_13250,N_10162,N_9804);
xor U13251 (N_13251,N_8838,N_10730);
xnor U13252 (N_13252,N_8734,N_11146);
or U13253 (N_13253,N_9017,N_11974);
nand U13254 (N_13254,N_11733,N_9824);
nand U13255 (N_13255,N_9349,N_8579);
nand U13256 (N_13256,N_9749,N_8091);
nor U13257 (N_13257,N_9921,N_8605);
nor U13258 (N_13258,N_8139,N_8189);
or U13259 (N_13259,N_8679,N_8570);
and U13260 (N_13260,N_8173,N_9562);
or U13261 (N_13261,N_9410,N_10412);
nor U13262 (N_13262,N_10620,N_9732);
and U13263 (N_13263,N_8933,N_10046);
nor U13264 (N_13264,N_8636,N_11242);
and U13265 (N_13265,N_10868,N_9550);
nand U13266 (N_13266,N_10779,N_8443);
or U13267 (N_13267,N_9012,N_10011);
xor U13268 (N_13268,N_10581,N_9414);
xor U13269 (N_13269,N_8723,N_8407);
and U13270 (N_13270,N_8617,N_10458);
and U13271 (N_13271,N_11478,N_11051);
nand U13272 (N_13272,N_10298,N_11842);
nand U13273 (N_13273,N_8722,N_9693);
and U13274 (N_13274,N_8468,N_11779);
or U13275 (N_13275,N_10177,N_11255);
and U13276 (N_13276,N_11782,N_11862);
nand U13277 (N_13277,N_10834,N_8246);
xnor U13278 (N_13278,N_9201,N_10339);
nor U13279 (N_13279,N_9739,N_10406);
nand U13280 (N_13280,N_10317,N_11112);
nand U13281 (N_13281,N_10415,N_9318);
nand U13282 (N_13282,N_11068,N_10972);
and U13283 (N_13283,N_9994,N_11428);
or U13284 (N_13284,N_11459,N_9790);
nor U13285 (N_13285,N_10034,N_10411);
nand U13286 (N_13286,N_9142,N_9825);
xnor U13287 (N_13287,N_10821,N_8047);
and U13288 (N_13288,N_10573,N_9057);
nand U13289 (N_13289,N_9073,N_11797);
nand U13290 (N_13290,N_8666,N_10126);
nor U13291 (N_13291,N_10116,N_11449);
and U13292 (N_13292,N_9567,N_9440);
nand U13293 (N_13293,N_10135,N_11553);
xnor U13294 (N_13294,N_10093,N_11621);
or U13295 (N_13295,N_9464,N_9784);
or U13296 (N_13296,N_10083,N_10042);
and U13297 (N_13297,N_8075,N_9942);
nor U13298 (N_13298,N_11421,N_10219);
or U13299 (N_13299,N_11494,N_11410);
xnor U13300 (N_13300,N_10597,N_11713);
or U13301 (N_13301,N_8470,N_8960);
nand U13302 (N_13302,N_8774,N_8432);
nand U13303 (N_13303,N_10355,N_8765);
xnor U13304 (N_13304,N_9905,N_8089);
and U13305 (N_13305,N_10891,N_8258);
and U13306 (N_13306,N_9356,N_9438);
and U13307 (N_13307,N_9897,N_10697);
and U13308 (N_13308,N_9745,N_8600);
xnor U13309 (N_13309,N_10840,N_8016);
and U13310 (N_13310,N_10519,N_9406);
and U13311 (N_13311,N_11336,N_9625);
nor U13312 (N_13312,N_8283,N_10407);
nor U13313 (N_13313,N_9802,N_11816);
and U13314 (N_13314,N_11424,N_9560);
and U13315 (N_13315,N_8024,N_9259);
nor U13316 (N_13316,N_10699,N_9951);
nand U13317 (N_13317,N_8220,N_8623);
nand U13318 (N_13318,N_11147,N_11266);
or U13319 (N_13319,N_10459,N_11800);
xor U13320 (N_13320,N_9173,N_10604);
or U13321 (N_13321,N_10749,N_9059);
and U13322 (N_13322,N_8312,N_9832);
and U13323 (N_13323,N_8923,N_9688);
xor U13324 (N_13324,N_11583,N_9531);
and U13325 (N_13325,N_8683,N_9083);
and U13326 (N_13326,N_8697,N_9067);
and U13327 (N_13327,N_11566,N_8442);
or U13328 (N_13328,N_8825,N_9258);
nand U13329 (N_13329,N_11846,N_10481);
nand U13330 (N_13330,N_8547,N_11422);
xnor U13331 (N_13331,N_11906,N_10456);
or U13332 (N_13332,N_10263,N_10996);
nor U13333 (N_13333,N_9149,N_10430);
nor U13334 (N_13334,N_8020,N_8857);
nand U13335 (N_13335,N_8668,N_11214);
nand U13336 (N_13336,N_11217,N_8850);
or U13337 (N_13337,N_10563,N_11969);
and U13338 (N_13338,N_9132,N_10860);
and U13339 (N_13339,N_9955,N_8551);
or U13340 (N_13340,N_10696,N_8247);
nand U13341 (N_13341,N_8811,N_9454);
nand U13342 (N_13342,N_8927,N_11063);
nand U13343 (N_13343,N_9617,N_9689);
and U13344 (N_13344,N_11709,N_8720);
and U13345 (N_13345,N_10986,N_10131);
xor U13346 (N_13346,N_8438,N_11443);
nor U13347 (N_13347,N_11603,N_11177);
nand U13348 (N_13348,N_10741,N_8106);
nor U13349 (N_13349,N_8240,N_8743);
nand U13350 (N_13350,N_11327,N_9379);
nor U13351 (N_13351,N_10079,N_10198);
or U13352 (N_13352,N_10624,N_9810);
nand U13353 (N_13353,N_9013,N_8165);
nor U13354 (N_13354,N_9421,N_9320);
nor U13355 (N_13355,N_10141,N_8080);
nand U13356 (N_13356,N_10414,N_9060);
nor U13357 (N_13357,N_10712,N_8181);
nor U13358 (N_13358,N_10143,N_8633);
and U13359 (N_13359,N_10856,N_9277);
nand U13360 (N_13360,N_8536,N_9384);
nand U13361 (N_13361,N_11092,N_8979);
and U13362 (N_13362,N_11019,N_11504);
nor U13363 (N_13363,N_11662,N_9346);
and U13364 (N_13364,N_10348,N_10846);
nand U13365 (N_13365,N_11890,N_11814);
or U13366 (N_13366,N_9058,N_8277);
nor U13367 (N_13367,N_10125,N_11680);
or U13368 (N_13368,N_8768,N_11184);
or U13369 (N_13369,N_10901,N_11230);
or U13370 (N_13370,N_8649,N_9923);
nor U13371 (N_13371,N_11829,N_11743);
or U13372 (N_13372,N_9338,N_10567);
or U13373 (N_13373,N_10205,N_10756);
xnor U13374 (N_13374,N_8439,N_11382);
and U13375 (N_13375,N_11815,N_11939);
nand U13376 (N_13376,N_8630,N_9582);
nand U13377 (N_13377,N_9195,N_9612);
xnor U13378 (N_13378,N_10000,N_8793);
and U13379 (N_13379,N_11995,N_9282);
or U13380 (N_13380,N_10675,N_11664);
nand U13381 (N_13381,N_8580,N_9018);
and U13382 (N_13382,N_10400,N_8858);
nor U13383 (N_13383,N_8143,N_8455);
nor U13384 (N_13384,N_8239,N_9066);
and U13385 (N_13385,N_11296,N_9321);
or U13386 (N_13386,N_8974,N_10857);
or U13387 (N_13387,N_11856,N_9914);
nand U13388 (N_13388,N_9911,N_11091);
nor U13389 (N_13389,N_9241,N_8665);
nor U13390 (N_13390,N_11352,N_11701);
nand U13391 (N_13391,N_11670,N_10112);
nand U13392 (N_13392,N_10742,N_11568);
nor U13393 (N_13393,N_8368,N_8224);
nor U13394 (N_13394,N_8416,N_10025);
xor U13395 (N_13395,N_9151,N_8429);
nand U13396 (N_13396,N_9713,N_11876);
xnor U13397 (N_13397,N_9934,N_9055);
or U13398 (N_13398,N_8735,N_9535);
nor U13399 (N_13399,N_11924,N_11188);
nor U13400 (N_13400,N_9920,N_11576);
nand U13401 (N_13401,N_8149,N_11406);
xor U13402 (N_13402,N_10128,N_11444);
and U13403 (N_13403,N_11237,N_11498);
xor U13404 (N_13404,N_11071,N_9948);
and U13405 (N_13405,N_11021,N_11208);
or U13406 (N_13406,N_8338,N_9906);
nand U13407 (N_13407,N_11912,N_9444);
and U13408 (N_13408,N_11760,N_9485);
and U13409 (N_13409,N_9484,N_10049);
and U13410 (N_13410,N_9644,N_11739);
nor U13411 (N_13411,N_9798,N_10537);
xor U13412 (N_13412,N_10740,N_10231);
xnor U13413 (N_13413,N_8859,N_8711);
xnor U13414 (N_13414,N_8949,N_8736);
and U13415 (N_13415,N_9514,N_10218);
nand U13416 (N_13416,N_9075,N_11122);
nor U13417 (N_13417,N_8750,N_9635);
or U13418 (N_13418,N_9033,N_8798);
nor U13419 (N_13419,N_11968,N_11356);
or U13420 (N_13420,N_11044,N_11724);
nand U13421 (N_13421,N_11947,N_8890);
nand U13422 (N_13422,N_11058,N_9089);
and U13423 (N_13423,N_10014,N_9047);
nand U13424 (N_13424,N_11317,N_8052);
nor U13425 (N_13425,N_8685,N_10349);
xnor U13426 (N_13426,N_9079,N_11181);
xnor U13427 (N_13427,N_9591,N_8345);
xnor U13428 (N_13428,N_8502,N_8640);
and U13429 (N_13429,N_9361,N_8639);
nand U13430 (N_13430,N_8578,N_8046);
or U13431 (N_13431,N_8107,N_8421);
xor U13432 (N_13432,N_8485,N_8362);
xnor U13433 (N_13433,N_10053,N_8508);
nand U13434 (N_13434,N_11174,N_9781);
nand U13435 (N_13435,N_10930,N_10508);
xnor U13436 (N_13436,N_10172,N_9397);
and U13437 (N_13437,N_9076,N_11325);
or U13438 (N_13438,N_11160,N_9706);
xnor U13439 (N_13439,N_10899,N_9216);
xor U13440 (N_13440,N_11116,N_10551);
xor U13441 (N_13441,N_11056,N_10156);
or U13442 (N_13442,N_9225,N_11715);
and U13443 (N_13443,N_8852,N_11601);
xnor U13444 (N_13444,N_8951,N_11544);
nor U13445 (N_13445,N_9374,N_11251);
and U13446 (N_13446,N_10837,N_10436);
xor U13447 (N_13447,N_8821,N_8704);
nor U13448 (N_13448,N_8315,N_11062);
xor U13449 (N_13449,N_10951,N_10129);
nand U13450 (N_13450,N_10807,N_9490);
xnor U13451 (N_13451,N_9179,N_8370);
nor U13452 (N_13452,N_10767,N_8035);
xnor U13453 (N_13453,N_11649,N_11306);
nor U13454 (N_13454,N_9637,N_9666);
and U13455 (N_13455,N_8413,N_9422);
xor U13456 (N_13456,N_9558,N_10440);
xnor U13457 (N_13457,N_9400,N_8111);
nand U13458 (N_13458,N_10250,N_9915);
nor U13459 (N_13459,N_8954,N_10292);
nand U13460 (N_13460,N_11721,N_9944);
or U13461 (N_13461,N_11726,N_11530);
xnor U13462 (N_13462,N_9821,N_11106);
or U13463 (N_13463,N_10497,N_9773);
nand U13464 (N_13464,N_8642,N_11412);
xnor U13465 (N_13465,N_8847,N_8105);
and U13466 (N_13466,N_8461,N_10822);
nor U13467 (N_13467,N_9208,N_8201);
nor U13468 (N_13468,N_8288,N_11436);
nor U13469 (N_13469,N_10938,N_10527);
nand U13470 (N_13470,N_11518,N_11960);
nand U13471 (N_13471,N_10685,N_10472);
and U13472 (N_13472,N_10594,N_10163);
xor U13473 (N_13473,N_10354,N_9085);
nand U13474 (N_13474,N_10576,N_10432);
xnor U13475 (N_13475,N_11626,N_10878);
nand U13476 (N_13476,N_8164,N_11984);
nor U13477 (N_13477,N_11045,N_8961);
nor U13478 (N_13478,N_11462,N_8777);
xnor U13479 (N_13479,N_10502,N_9314);
or U13480 (N_13480,N_8004,N_10570);
nor U13481 (N_13481,N_11402,N_11013);
and U13482 (N_13482,N_9409,N_10136);
or U13483 (N_13483,N_8631,N_9453);
and U13484 (N_13484,N_8706,N_8773);
nor U13485 (N_13485,N_10988,N_9155);
nand U13486 (N_13486,N_10388,N_10035);
or U13487 (N_13487,N_9184,N_10723);
xor U13488 (N_13488,N_8228,N_8415);
nand U13489 (N_13489,N_11614,N_10234);
xnor U13490 (N_13490,N_9624,N_11855);
xor U13491 (N_13491,N_10709,N_9848);
and U13492 (N_13492,N_9502,N_10903);
xor U13493 (N_13493,N_10845,N_9205);
nor U13494 (N_13494,N_9498,N_11273);
xnor U13495 (N_13495,N_9212,N_11507);
or U13496 (N_13496,N_8561,N_8504);
or U13497 (N_13497,N_8087,N_9641);
xor U13498 (N_13498,N_10693,N_11872);
xnor U13499 (N_13499,N_11579,N_8133);
xor U13500 (N_13500,N_10998,N_8682);
nor U13501 (N_13501,N_10464,N_8965);
and U13502 (N_13502,N_8572,N_8083);
nand U13503 (N_13503,N_9196,N_11985);
nor U13504 (N_13504,N_11043,N_8483);
or U13505 (N_13505,N_10327,N_8546);
nand U13506 (N_13506,N_9977,N_8172);
or U13507 (N_13507,N_10539,N_10724);
nand U13508 (N_13508,N_11848,N_8780);
or U13509 (N_13509,N_10328,N_10383);
nand U13510 (N_13510,N_11620,N_10004);
nand U13511 (N_13511,N_8475,N_11694);
xnor U13512 (N_13512,N_10201,N_11850);
nor U13513 (N_13513,N_8500,N_9220);
and U13514 (N_13514,N_9940,N_11751);
nand U13515 (N_13515,N_10159,N_11898);
nand U13516 (N_13516,N_11081,N_9855);
nand U13517 (N_13517,N_8888,N_9078);
nor U13518 (N_13518,N_10302,N_11923);
nand U13519 (N_13519,N_8114,N_9552);
xor U13520 (N_13520,N_8000,N_11688);
and U13521 (N_13521,N_9390,N_9952);
nor U13522 (N_13522,N_8398,N_11003);
and U13523 (N_13523,N_8010,N_11085);
or U13524 (N_13524,N_8644,N_8926);
nand U13525 (N_13525,N_8447,N_9284);
nand U13526 (N_13526,N_10646,N_8195);
xnor U13527 (N_13527,N_9718,N_11203);
and U13528 (N_13528,N_10052,N_10882);
or U13529 (N_13529,N_10940,N_11634);
and U13530 (N_13530,N_10133,N_8124);
nand U13531 (N_13531,N_11129,N_11950);
nand U13532 (N_13532,N_10921,N_9247);
or U13533 (N_13533,N_10735,N_10240);
and U13534 (N_13534,N_10157,N_9577);
xor U13535 (N_13535,N_9355,N_8934);
or U13536 (N_13536,N_8045,N_10747);
nor U13537 (N_13537,N_9945,N_11467);
and U13538 (N_13538,N_11221,N_11562);
and U13539 (N_13539,N_10650,N_8593);
nand U13540 (N_13540,N_8732,N_11178);
or U13541 (N_13541,N_9106,N_8187);
nor U13542 (N_13542,N_8473,N_9133);
xor U13543 (N_13543,N_9561,N_10227);
nor U13544 (N_13544,N_8152,N_10168);
and U13545 (N_13545,N_11622,N_10990);
and U13546 (N_13546,N_8549,N_9372);
and U13547 (N_13547,N_9111,N_11750);
xnor U13548 (N_13548,N_8057,N_11405);
or U13549 (N_13549,N_8347,N_10465);
nor U13550 (N_13550,N_9538,N_11033);
nor U13551 (N_13551,N_8135,N_10324);
nand U13552 (N_13552,N_11018,N_9147);
or U13553 (N_13553,N_11770,N_8230);
nor U13554 (N_13554,N_8156,N_11222);
nand U13555 (N_13555,N_11532,N_11908);
and U13556 (N_13556,N_10397,N_9631);
nand U13557 (N_13557,N_11320,N_11133);
xnor U13558 (N_13558,N_11464,N_9074);
and U13559 (N_13559,N_11419,N_8509);
nand U13560 (N_13560,N_9000,N_8070);
and U13561 (N_13561,N_10466,N_11496);
and U13562 (N_13562,N_8307,N_10330);
nand U13563 (N_13563,N_9929,N_8615);
and U13564 (N_13564,N_8729,N_10843);
and U13565 (N_13565,N_11448,N_8710);
and U13566 (N_13566,N_10959,N_11064);
nor U13567 (N_13567,N_10645,N_8701);
or U13568 (N_13568,N_10150,N_8656);
xnor U13569 (N_13569,N_11392,N_9714);
nor U13570 (N_13570,N_10269,N_8462);
or U13571 (N_13571,N_8795,N_9515);
nor U13572 (N_13572,N_11322,N_11728);
and U13573 (N_13573,N_8452,N_11958);
or U13574 (N_13574,N_10312,N_8497);
xnor U13575 (N_13575,N_11358,N_11545);
and U13576 (N_13576,N_8724,N_8627);
or U13577 (N_13577,N_9450,N_8097);
xnor U13578 (N_13578,N_11643,N_11826);
nor U13579 (N_13579,N_8144,N_11293);
and U13580 (N_13580,N_8001,N_10982);
nor U13581 (N_13581,N_10780,N_11878);
xnor U13582 (N_13582,N_11569,N_10586);
nor U13583 (N_13583,N_9634,N_9527);
nand U13584 (N_13584,N_8776,N_11332);
xor U13585 (N_13585,N_11648,N_8211);
xnor U13586 (N_13586,N_10844,N_11067);
and U13587 (N_13587,N_11202,N_9841);
nor U13588 (N_13588,N_10183,N_8115);
or U13589 (N_13589,N_11311,N_11446);
nand U13590 (N_13590,N_8556,N_10278);
or U13591 (N_13591,N_9257,N_10503);
xor U13592 (N_13592,N_10268,N_10387);
and U13593 (N_13593,N_11453,N_9975);
xor U13594 (N_13594,N_8752,N_11533);
xor U13595 (N_13595,N_9756,N_11798);
nor U13596 (N_13596,N_11735,N_11245);
or U13597 (N_13597,N_8248,N_11996);
or U13598 (N_13598,N_9301,N_8467);
nand U13599 (N_13599,N_9628,N_8762);
nor U13600 (N_13600,N_11520,N_11131);
xor U13601 (N_13601,N_11953,N_8012);
nor U13602 (N_13602,N_11447,N_8202);
nor U13603 (N_13603,N_9344,N_11275);
nand U13604 (N_13604,N_10953,N_9082);
xnor U13605 (N_13605,N_8896,N_11588);
nand U13606 (N_13606,N_8015,N_11008);
or U13607 (N_13607,N_8717,N_11549);
and U13608 (N_13608,N_10981,N_11164);
nor U13609 (N_13609,N_8891,N_10555);
nand U13610 (N_13610,N_11511,N_10185);
nand U13611 (N_13611,N_10824,N_11501);
or U13612 (N_13612,N_10893,N_9378);
or U13613 (N_13613,N_8183,N_11914);
xnor U13614 (N_13614,N_10612,N_11431);
xnor U13615 (N_13615,N_9366,N_10365);
and U13616 (N_13616,N_10918,N_9177);
and U13617 (N_13617,N_9008,N_11999);
and U13618 (N_13618,N_8832,N_10259);
nor U13619 (N_13619,N_10661,N_9263);
xnor U13620 (N_13620,N_8987,N_10423);
xor U13621 (N_13621,N_9686,N_8289);
xor U13622 (N_13622,N_9488,N_10676);
and U13623 (N_13623,N_11389,N_11423);
xnor U13624 (N_13624,N_8973,N_9588);
nand U13625 (N_13625,N_10873,N_11381);
xnor U13626 (N_13626,N_10285,N_10080);
nand U13627 (N_13627,N_10732,N_11206);
nand U13628 (N_13628,N_9221,N_9095);
nand U13629 (N_13629,N_11264,N_9543);
nand U13630 (N_13630,N_8622,N_8748);
nand U13631 (N_13631,N_9061,N_11913);
xor U13632 (N_13632,N_10745,N_8886);
and U13633 (N_13633,N_10072,N_8897);
xnor U13634 (N_13634,N_10874,N_9799);
and U13635 (N_13635,N_8033,N_9433);
or U13636 (N_13636,N_11564,N_9137);
nand U13637 (N_13637,N_9171,N_10701);
or U13638 (N_13638,N_9449,N_11962);
xor U13639 (N_13639,N_10461,N_9273);
xor U13640 (N_13640,N_9695,N_9466);
nand U13641 (N_13641,N_11460,N_10912);
and U13642 (N_13642,N_10350,N_11401);
xor U13643 (N_13643,N_8029,N_11977);
and U13644 (N_13644,N_9369,N_9481);
or U13645 (N_13645,N_9451,N_8741);
xor U13646 (N_13646,N_8273,N_8280);
or U13647 (N_13647,N_11309,N_9563);
and U13648 (N_13648,N_10314,N_10634);
nand U13649 (N_13649,N_9276,N_8419);
or U13650 (N_13650,N_10353,N_8980);
or U13651 (N_13651,N_10372,N_11191);
or U13652 (N_13652,N_9568,N_10443);
nor U13653 (N_13653,N_8538,N_10134);
or U13654 (N_13654,N_9457,N_10318);
nand U13655 (N_13655,N_11647,N_11076);
and U13656 (N_13656,N_11192,N_9694);
nor U13657 (N_13657,N_10544,N_8863);
nor U13658 (N_13658,N_8123,N_8138);
nand U13659 (N_13659,N_11597,N_9202);
and U13660 (N_13660,N_9702,N_8384);
xnor U13661 (N_13661,N_10118,N_11608);
xnor U13662 (N_13662,N_11875,N_10801);
and U13663 (N_13663,N_9615,N_11053);
and U13664 (N_13664,N_10256,N_10271);
nand U13665 (N_13665,N_9236,N_10629);
nand U13666 (N_13666,N_10284,N_11994);
and U13667 (N_13667,N_11373,N_9508);
xor U13668 (N_13668,N_11285,N_10717);
xor U13669 (N_13669,N_8643,N_9993);
or U13670 (N_13670,N_9071,N_10473);
xor U13671 (N_13671,N_11809,N_9285);
nor U13672 (N_13672,N_11840,N_8690);
xor U13673 (N_13673,N_10066,N_9497);
xnor U13674 (N_13674,N_9513,N_10905);
xnor U13675 (N_13675,N_11347,N_8956);
xnor U13676 (N_13676,N_10410,N_10684);
and U13677 (N_13677,N_10582,N_11659);
xor U13678 (N_13678,N_11173,N_10226);
nor U13679 (N_13679,N_11792,N_10304);
or U13680 (N_13680,N_9491,N_11516);
xnor U13681 (N_13681,N_8425,N_8906);
xor U13682 (N_13682,N_11700,N_9053);
nand U13683 (N_13683,N_10030,N_10790);
xor U13684 (N_13684,N_8049,N_11526);
xnor U13685 (N_13685,N_9046,N_10653);
and U13686 (N_13686,N_11976,N_10761);
nand U13687 (N_13687,N_10369,N_8093);
nor U13688 (N_13688,N_11807,N_8607);
and U13689 (N_13689,N_11200,N_9162);
nor U13690 (N_13690,N_8206,N_8372);
nand U13691 (N_13691,N_9657,N_9875);
nand U13692 (N_13692,N_11383,N_10290);
or U13693 (N_13693,N_8866,N_9459);
xor U13694 (N_13694,N_11438,N_10392);
and U13695 (N_13695,N_8749,N_8263);
or U13696 (N_13696,N_10338,N_10737);
nor U13697 (N_13697,N_8494,N_9286);
nand U13698 (N_13698,N_9910,N_10952);
and U13699 (N_13699,N_8959,N_8598);
or U13700 (N_13700,N_10910,N_10962);
nand U13701 (N_13701,N_11993,N_9371);
xor U13702 (N_13702,N_11246,N_11175);
nand U13703 (N_13703,N_8518,N_11036);
nand U13704 (N_13704,N_8945,N_10799);
and U13705 (N_13705,N_11158,N_8833);
and U13706 (N_13706,N_11048,N_9717);
xnor U13707 (N_13707,N_10007,N_11907);
nand U13708 (N_13708,N_9573,N_11678);
nand U13709 (N_13709,N_9042,N_10635);
and U13710 (N_13710,N_9254,N_8354);
nor U13711 (N_13711,N_10161,N_9658);
xor U13712 (N_13712,N_11134,N_9520);
nor U13713 (N_13713,N_9062,N_11377);
nor U13714 (N_13714,N_9721,N_11473);
nand U13715 (N_13715,N_9458,N_10282);
nand U13716 (N_13716,N_9113,N_10803);
nor U13717 (N_13717,N_8034,N_9140);
and U13718 (N_13718,N_9509,N_11065);
or U13719 (N_13719,N_10293,N_8571);
nand U13720 (N_13720,N_11578,N_10334);
or U13721 (N_13721,N_11215,N_11868);
or U13722 (N_13722,N_11468,N_10409);
nor U13723 (N_13723,N_9024,N_11059);
or U13724 (N_13724,N_11477,N_8905);
nor U13725 (N_13725,N_8510,N_10553);
or U13726 (N_13726,N_10787,N_8150);
or U13727 (N_13727,N_9364,N_8560);
or U13728 (N_13728,N_10867,N_9578);
nand U13729 (N_13729,N_10887,N_8747);
nand U13730 (N_13730,N_10021,N_11120);
nor U13731 (N_13731,N_9229,N_11669);
xor U13732 (N_13732,N_11457,N_11682);
or U13733 (N_13733,N_8512,N_10097);
nand U13734 (N_13734,N_10274,N_11920);
or U13735 (N_13735,N_9964,N_10558);
xor U13736 (N_13736,N_11425,N_11016);
xnor U13737 (N_13737,N_8088,N_9677);
or U13738 (N_13738,N_9383,N_9740);
and U13739 (N_13739,N_9278,N_10965);
or U13740 (N_13740,N_9381,N_11627);
nand U13741 (N_13741,N_8053,N_8249);
xor U13742 (N_13742,N_10065,N_11277);
and U13743 (N_13743,N_11551,N_11796);
and U13744 (N_13744,N_9117,N_10467);
and U13745 (N_13745,N_11600,N_9224);
or U13746 (N_13746,N_10517,N_9300);
nand U13747 (N_13747,N_10906,N_11656);
xnor U13748 (N_13748,N_8440,N_9836);
nor U13749 (N_13749,N_8658,N_10232);
nand U13750 (N_13750,N_10974,N_10300);
nor U13751 (N_13751,N_9373,N_9281);
xnor U13752 (N_13752,N_8410,N_11757);
and U13753 (N_13753,N_9139,N_9559);
or U13754 (N_13754,N_9705,N_9654);
xnor U13755 (N_13755,N_8460,N_8805);
or U13756 (N_13756,N_11729,N_9441);
and U13757 (N_13757,N_8256,N_8084);
xnor U13758 (N_13758,N_11166,N_8401);
and U13759 (N_13759,N_9678,N_8889);
xor U13760 (N_13760,N_10838,N_10714);
xor U13761 (N_13761,N_11535,N_10069);
nor U13762 (N_13762,N_9063,N_11595);
or U13763 (N_13763,N_11201,N_10892);
and U13764 (N_13764,N_9186,N_11313);
and U13765 (N_13765,N_8218,N_9868);
nand U13766 (N_13766,N_11140,N_11179);
xor U13767 (N_13767,N_10358,N_9154);
nand U13768 (N_13768,N_8018,N_8491);
and U13769 (N_13769,N_8456,N_10110);
xnor U13770 (N_13770,N_8155,N_9997);
nor U13771 (N_13771,N_8937,N_9621);
or U13772 (N_13772,N_11888,N_8487);
and U13773 (N_13773,N_10598,N_9170);
nor U13774 (N_13774,N_9539,N_8250);
nor U13775 (N_13775,N_11372,N_10158);
nor U13776 (N_13776,N_10681,N_10605);
and U13777 (N_13777,N_11880,N_8804);
and U13778 (N_13778,N_9570,N_10147);
or U13779 (N_13779,N_8360,N_10885);
xor U13780 (N_13780,N_10731,N_8807);
nand U13781 (N_13781,N_9317,N_10504);
xor U13782 (N_13782,N_10401,N_8964);
xnor U13783 (N_13783,N_10966,N_11970);
xor U13784 (N_13784,N_9650,N_9556);
xnor U13785 (N_13785,N_10055,N_8065);
nand U13786 (N_13786,N_11889,N_9312);
and U13787 (N_13787,N_8061,N_10013);
nor U13788 (N_13788,N_8374,N_9716);
xor U13789 (N_13789,N_8011,N_11822);
nand U13790 (N_13790,N_10127,N_9129);
xnor U13791 (N_13791,N_9148,N_11261);
and U13792 (N_13792,N_9917,N_8158);
or U13793 (N_13793,N_10357,N_9238);
xnor U13794 (N_13794,N_11818,N_11426);
and U13795 (N_13795,N_11123,N_10743);
xor U13796 (N_13796,N_9130,N_11294);
nor U13797 (N_13797,N_10262,N_9754);
and U13798 (N_13798,N_11345,N_9330);
and U13799 (N_13799,N_8555,N_8436);
nor U13800 (N_13800,N_8567,N_8887);
xnor U13801 (N_13801,N_11461,N_11038);
xor U13802 (N_13802,N_11054,N_8528);
or U13803 (N_13803,N_8932,N_9950);
xor U13804 (N_13804,N_8950,N_11637);
and U13805 (N_13805,N_8655,N_9916);
xor U13806 (N_13806,N_11265,N_10565);
or U13807 (N_13807,N_10280,N_9506);
nand U13808 (N_13808,N_11069,N_11933);
or U13809 (N_13809,N_8803,N_10568);
nor U13810 (N_13810,N_9269,N_8193);
nor U13811 (N_13811,N_10070,N_11126);
and U13812 (N_13812,N_9416,N_8756);
or U13813 (N_13813,N_8709,N_11765);
or U13814 (N_13814,N_9333,N_9528);
xor U13815 (N_13815,N_9607,N_11866);
and U13816 (N_13816,N_9554,N_9785);
nand U13817 (N_13817,N_11992,N_11773);
nor U13818 (N_13818,N_8332,N_8638);
xor U13819 (N_13819,N_11882,N_8875);
or U13820 (N_13820,N_11640,N_9471);
xnor U13821 (N_13821,N_11731,N_9953);
nor U13822 (N_13822,N_8122,N_8488);
and U13823 (N_13823,N_9892,N_8233);
or U13824 (N_13824,N_9475,N_10526);
xor U13825 (N_13825,N_9640,N_8023);
or U13826 (N_13826,N_10777,N_8946);
nor U13827 (N_13827,N_8851,N_9297);
or U13828 (N_13828,N_9823,N_9928);
or U13829 (N_13829,N_9512,N_8885);
and U13830 (N_13830,N_8558,N_8200);
nor U13831 (N_13831,N_11570,N_11991);
nand U13832 (N_13832,N_11905,N_8104);
nor U13833 (N_13833,N_11376,N_8562);
or U13834 (N_13834,N_8341,N_10855);
nor U13835 (N_13835,N_8056,N_8693);
and U13836 (N_13836,N_9190,N_8299);
or U13837 (N_13837,N_8252,N_10009);
nand U13838 (N_13838,N_10771,N_9478);
nand U13839 (N_13839,N_11941,N_9146);
nor U13840 (N_13840,N_9415,N_10512);
and U13841 (N_13841,N_11308,N_11910);
or U13842 (N_13842,N_11722,N_10325);
or U13843 (N_13843,N_10207,N_11521);
or U13844 (N_13844,N_9966,N_9005);
nand U13845 (N_13845,N_10751,N_11487);
and U13846 (N_13846,N_8357,N_9764);
or U13847 (N_13847,N_11385,N_9420);
xnor U13848 (N_13848,N_8784,N_8005);
nor U13849 (N_13849,N_10950,N_11885);
and U13850 (N_13850,N_11668,N_10094);
nor U13851 (N_13851,N_9746,N_11476);
xor U13852 (N_13852,N_10985,N_9118);
nand U13853 (N_13853,N_9899,N_11695);
nor U13854 (N_13854,N_10041,N_11673);
or U13855 (N_13855,N_8744,N_9165);
xnor U13856 (N_13856,N_11853,N_9261);
or U13857 (N_13857,N_9788,N_11618);
nor U13858 (N_13858,N_10102,N_8698);
nand U13859 (N_13859,N_9633,N_10463);
or U13860 (N_13860,N_9026,N_9136);
nor U13861 (N_13861,N_9601,N_11711);
nand U13862 (N_13862,N_10698,N_10115);
or U13863 (N_13863,N_10364,N_11093);
and U13864 (N_13864,N_9743,N_8351);
or U13865 (N_13865,N_10694,N_11046);
xor U13866 (N_13866,N_9744,N_10050);
nand U13867 (N_13867,N_9611,N_9339);
nor U13868 (N_13868,N_9427,N_10804);
nor U13869 (N_13869,N_11225,N_9336);
nand U13870 (N_13870,N_11954,N_9309);
nand U13871 (N_13871,N_9792,N_10233);
nand U13872 (N_13872,N_11934,N_10213);
nand U13873 (N_13873,N_8873,N_9108);
and U13874 (N_13874,N_10736,N_11636);
and U13875 (N_13875,N_11454,N_9783);
or U13876 (N_13876,N_9704,N_8269);
or U13877 (N_13877,N_10859,N_9683);
and U13878 (N_13878,N_10220,N_9482);
nand U13879 (N_13879,N_9473,N_11209);
and U13880 (N_13880,N_10012,N_8501);
nor U13881 (N_13881,N_8435,N_10108);
nor U13882 (N_13882,N_10342,N_8121);
nand U13883 (N_13883,N_11808,N_8574);
and U13884 (N_13884,N_8613,N_8032);
nand U13885 (N_13885,N_9228,N_8296);
and U13886 (N_13886,N_11007,N_8880);
nor U13887 (N_13887,N_8977,N_10239);
nor U13888 (N_13888,N_9088,N_11926);
or U13889 (N_13889,N_10389,N_9323);
or U13890 (N_13890,N_11216,N_10691);
and U13891 (N_13891,N_9065,N_9867);
or U13892 (N_13892,N_8554,N_8377);
and U13893 (N_13893,N_10345,N_8286);
xor U13894 (N_13894,N_8326,N_8746);
or U13895 (N_13895,N_10422,N_8779);
and U13896 (N_13896,N_8192,N_10429);
nor U13897 (N_13897,N_9834,N_8177);
nand U13898 (N_13898,N_11617,N_10319);
xor U13899 (N_13899,N_10103,N_9215);
nand U13900 (N_13900,N_9213,N_8463);
nand U13901 (N_13901,N_11338,N_9503);
or U13902 (N_13902,N_8940,N_11287);
and U13903 (N_13903,N_10592,N_10819);
and U13904 (N_13904,N_9597,N_8503);
nand U13905 (N_13905,N_8437,N_9391);
and U13906 (N_13906,N_9774,N_11491);
and U13907 (N_13907,N_9394,N_10929);
or U13908 (N_13908,N_8972,N_10858);
xnor U13909 (N_13909,N_10509,N_9874);
nand U13910 (N_13910,N_9325,N_9758);
xor U13911 (N_13911,N_8103,N_10641);
nand U13912 (N_13912,N_9370,N_9268);
nor U13913 (N_13913,N_8994,N_10470);
nor U13914 (N_13914,N_8313,N_9092);
and U13915 (N_13915,N_10556,N_11593);
and U13916 (N_13916,N_8854,N_11474);
nand U13917 (N_13917,N_10778,N_8096);
nand U13918 (N_13918,N_10518,N_9487);
and U13919 (N_13919,N_11658,N_9262);
nor U13920 (N_13920,N_11367,N_11034);
xnor U13921 (N_13921,N_11442,N_11741);
xor U13922 (N_13922,N_10488,N_10395);
or U13923 (N_13923,N_8763,N_11128);
xor U13924 (N_13924,N_9726,N_8025);
xnor U13925 (N_13925,N_10019,N_8740);
and U13926 (N_13926,N_10281,N_8002);
nor U13927 (N_13927,N_8008,N_8079);
and U13928 (N_13928,N_9283,N_9885);
xnor U13929 (N_13929,N_11821,N_11195);
nor U13930 (N_13930,N_8316,N_8366);
and U13931 (N_13931,N_11810,N_9930);
or U13932 (N_13932,N_10480,N_10433);
nand U13933 (N_13933,N_8125,N_10326);
and U13934 (N_13934,N_9909,N_10454);
xnor U13935 (N_13935,N_8154,N_10937);
nand U13936 (N_13936,N_9729,N_11001);
nor U13937 (N_13937,N_11100,N_11836);
xor U13938 (N_13938,N_10261,N_9990);
xnor U13939 (N_13939,N_10451,N_9725);
nor U13940 (N_13940,N_9525,N_8912);
or U13941 (N_13941,N_11155,N_10561);
nor U13942 (N_13942,N_11433,N_11655);
nor U13943 (N_13943,N_8314,N_11224);
nor U13944 (N_13944,N_8544,N_11488);
xnor U13945 (N_13945,N_11635,N_9791);
xor U13946 (N_13946,N_10705,N_10140);
xor U13947 (N_13947,N_8869,N_8306);
nand U13948 (N_13948,N_9122,N_10416);
or U13949 (N_13949,N_9816,N_10920);
and U13950 (N_13950,N_11572,N_8433);
xnor U13951 (N_13951,N_8619,N_11388);
nand U13952 (N_13952,N_10494,N_11159);
xnor U13953 (N_13953,N_10710,N_10206);
or U13954 (N_13954,N_9680,N_9674);
nand U13955 (N_13955,N_10909,N_11935);
xor U13956 (N_13956,N_8414,N_9462);
or U13957 (N_13957,N_8098,N_8305);
or U13958 (N_13958,N_8569,N_11151);
nor U13959 (N_13959,N_11326,N_10622);
xnor U13960 (N_13960,N_9696,N_11883);
or U13961 (N_13961,N_8009,N_8531);
xor U13962 (N_13962,N_11199,N_10487);
or U13963 (N_13963,N_11624,N_10095);
nor U13964 (N_13964,N_11485,N_11006);
nor U13965 (N_13965,N_10660,N_8899);
or U13966 (N_13966,N_11932,N_8420);
xnor U13967 (N_13967,N_11413,N_9272);
nand U13968 (N_13968,N_10187,N_9417);
xnor U13969 (N_13969,N_9762,N_11663);
nand U13970 (N_13970,N_8511,N_8990);
nor U13971 (N_13971,N_9499,N_8271);
xnor U13972 (N_13972,N_10798,N_11813);
nor U13973 (N_13973,N_11867,N_9794);
xnor U13974 (N_13974,N_8739,N_10204);
and U13975 (N_13975,N_9185,N_11186);
xor U13976 (N_13976,N_8941,N_9599);
or U13977 (N_13977,N_10408,N_9160);
and U13978 (N_13978,N_11998,N_9051);
nand U13979 (N_13979,N_11355,N_8095);
nor U13980 (N_13980,N_9653,N_10173);
xnor U13981 (N_13981,N_10104,N_11363);
nand U13982 (N_13982,N_11524,N_9999);
nand U13983 (N_13983,N_9927,N_11788);
and U13984 (N_13984,N_10222,N_9536);
nand U13985 (N_13985,N_9164,N_10911);
xnor U13986 (N_13986,N_8145,N_8234);
and U13987 (N_13987,N_8764,N_11778);
xnor U13988 (N_13988,N_9529,N_8484);
or U13989 (N_13989,N_9734,N_9328);
xor U13990 (N_13990,N_10479,N_9434);
xnor U13991 (N_13991,N_9733,N_10603);
nand U13992 (N_13992,N_11288,N_10197);
and U13993 (N_13993,N_8359,N_8255);
and U13994 (N_13994,N_10764,N_9072);
nor U13995 (N_13995,N_10373,N_8568);
nand U13996 (N_13996,N_10427,N_11594);
and U13997 (N_13997,N_8148,N_9853);
nand U13998 (N_13998,N_9308,N_9627);
xor U13999 (N_13999,N_9655,N_10993);
xor U14000 (N_14000,N_10698,N_11063);
or U14001 (N_14001,N_8167,N_9379);
nand U14002 (N_14002,N_10863,N_11553);
and U14003 (N_14003,N_9305,N_9121);
or U14004 (N_14004,N_11730,N_9222);
or U14005 (N_14005,N_9311,N_9506);
xor U14006 (N_14006,N_11206,N_9621);
nand U14007 (N_14007,N_11584,N_10491);
and U14008 (N_14008,N_11375,N_11693);
and U14009 (N_14009,N_11861,N_8531);
nand U14010 (N_14010,N_10338,N_9566);
nor U14011 (N_14011,N_9922,N_11041);
nand U14012 (N_14012,N_10980,N_9688);
or U14013 (N_14013,N_9422,N_11086);
nand U14014 (N_14014,N_10709,N_8808);
xor U14015 (N_14015,N_11848,N_10202);
xnor U14016 (N_14016,N_9257,N_11666);
xor U14017 (N_14017,N_11113,N_8096);
or U14018 (N_14018,N_9848,N_11654);
or U14019 (N_14019,N_10920,N_11408);
nor U14020 (N_14020,N_10980,N_11184);
and U14021 (N_14021,N_8099,N_10602);
nand U14022 (N_14022,N_8125,N_10146);
nor U14023 (N_14023,N_9402,N_11362);
nand U14024 (N_14024,N_8193,N_11173);
or U14025 (N_14025,N_9943,N_8948);
or U14026 (N_14026,N_10466,N_8425);
nor U14027 (N_14027,N_9783,N_10976);
or U14028 (N_14028,N_9809,N_9112);
nand U14029 (N_14029,N_10453,N_8702);
nand U14030 (N_14030,N_8771,N_10732);
or U14031 (N_14031,N_10775,N_8606);
xnor U14032 (N_14032,N_10810,N_10739);
xor U14033 (N_14033,N_9928,N_8099);
or U14034 (N_14034,N_9316,N_11489);
and U14035 (N_14035,N_11497,N_10575);
nor U14036 (N_14036,N_9582,N_8750);
nor U14037 (N_14037,N_9098,N_10041);
nor U14038 (N_14038,N_11465,N_11936);
nor U14039 (N_14039,N_11787,N_10293);
nor U14040 (N_14040,N_8441,N_8381);
or U14041 (N_14041,N_9037,N_11185);
xor U14042 (N_14042,N_8790,N_9516);
or U14043 (N_14043,N_11807,N_8082);
xor U14044 (N_14044,N_10620,N_9220);
and U14045 (N_14045,N_11569,N_8279);
and U14046 (N_14046,N_10341,N_8896);
nand U14047 (N_14047,N_11412,N_11877);
nand U14048 (N_14048,N_11406,N_10926);
or U14049 (N_14049,N_9390,N_9125);
or U14050 (N_14050,N_9116,N_8448);
nor U14051 (N_14051,N_9877,N_10122);
nor U14052 (N_14052,N_8416,N_10541);
xnor U14053 (N_14053,N_11828,N_10530);
nand U14054 (N_14054,N_10018,N_8311);
nand U14055 (N_14055,N_8719,N_8145);
nor U14056 (N_14056,N_10642,N_10019);
and U14057 (N_14057,N_10862,N_9047);
xor U14058 (N_14058,N_8835,N_11784);
nand U14059 (N_14059,N_8476,N_10477);
nor U14060 (N_14060,N_8768,N_10308);
and U14061 (N_14061,N_8758,N_9603);
xnor U14062 (N_14062,N_10810,N_10181);
nand U14063 (N_14063,N_11907,N_10298);
and U14064 (N_14064,N_9782,N_11952);
nand U14065 (N_14065,N_10157,N_11129);
xnor U14066 (N_14066,N_8117,N_10599);
nand U14067 (N_14067,N_8331,N_11579);
and U14068 (N_14068,N_8240,N_11184);
xnor U14069 (N_14069,N_9224,N_8084);
nand U14070 (N_14070,N_8433,N_9284);
and U14071 (N_14071,N_10086,N_8477);
xor U14072 (N_14072,N_9164,N_8874);
or U14073 (N_14073,N_10148,N_11275);
nor U14074 (N_14074,N_8947,N_8599);
nor U14075 (N_14075,N_11041,N_9727);
or U14076 (N_14076,N_11935,N_11418);
nor U14077 (N_14077,N_11367,N_11416);
nand U14078 (N_14078,N_9737,N_11584);
xor U14079 (N_14079,N_8517,N_9636);
and U14080 (N_14080,N_10977,N_11036);
or U14081 (N_14081,N_11176,N_8391);
nand U14082 (N_14082,N_11937,N_11242);
xnor U14083 (N_14083,N_8134,N_8235);
nand U14084 (N_14084,N_8228,N_11491);
and U14085 (N_14085,N_9147,N_10627);
and U14086 (N_14086,N_9881,N_10756);
nor U14087 (N_14087,N_9766,N_8332);
and U14088 (N_14088,N_10668,N_8145);
or U14089 (N_14089,N_9086,N_10238);
nand U14090 (N_14090,N_8672,N_8711);
nand U14091 (N_14091,N_11167,N_11065);
nand U14092 (N_14092,N_9825,N_8095);
nand U14093 (N_14093,N_11755,N_8887);
and U14094 (N_14094,N_8644,N_8937);
and U14095 (N_14095,N_10469,N_10959);
or U14096 (N_14096,N_9180,N_8015);
nand U14097 (N_14097,N_11644,N_11657);
nor U14098 (N_14098,N_8882,N_10471);
and U14099 (N_14099,N_11063,N_11670);
nand U14100 (N_14100,N_11895,N_11492);
or U14101 (N_14101,N_11615,N_10651);
nand U14102 (N_14102,N_9731,N_10243);
or U14103 (N_14103,N_11768,N_9731);
nor U14104 (N_14104,N_10803,N_8904);
xnor U14105 (N_14105,N_8962,N_8064);
nor U14106 (N_14106,N_11068,N_8289);
or U14107 (N_14107,N_8138,N_9767);
xnor U14108 (N_14108,N_11479,N_11251);
and U14109 (N_14109,N_8269,N_8801);
and U14110 (N_14110,N_10381,N_9093);
xor U14111 (N_14111,N_10109,N_9470);
nor U14112 (N_14112,N_9786,N_11063);
and U14113 (N_14113,N_8698,N_10383);
nor U14114 (N_14114,N_11976,N_9367);
nor U14115 (N_14115,N_8745,N_10403);
or U14116 (N_14116,N_9659,N_11365);
nor U14117 (N_14117,N_11373,N_10729);
nand U14118 (N_14118,N_11209,N_10745);
nand U14119 (N_14119,N_9716,N_10779);
xnor U14120 (N_14120,N_11221,N_11158);
and U14121 (N_14121,N_11147,N_10868);
or U14122 (N_14122,N_8422,N_10389);
nand U14123 (N_14123,N_10604,N_11106);
nand U14124 (N_14124,N_8141,N_9850);
and U14125 (N_14125,N_10255,N_11109);
and U14126 (N_14126,N_11326,N_10773);
nor U14127 (N_14127,N_10570,N_8706);
nand U14128 (N_14128,N_9619,N_9961);
or U14129 (N_14129,N_10777,N_10067);
nor U14130 (N_14130,N_8019,N_11025);
nor U14131 (N_14131,N_8075,N_9876);
nand U14132 (N_14132,N_9928,N_8911);
and U14133 (N_14133,N_11528,N_9384);
and U14134 (N_14134,N_10133,N_8425);
and U14135 (N_14135,N_11363,N_10484);
nand U14136 (N_14136,N_10906,N_8799);
xnor U14137 (N_14137,N_8829,N_9742);
and U14138 (N_14138,N_8600,N_10330);
or U14139 (N_14139,N_9369,N_9173);
and U14140 (N_14140,N_9875,N_9115);
xor U14141 (N_14141,N_10035,N_9423);
nor U14142 (N_14142,N_9825,N_8179);
xnor U14143 (N_14143,N_10873,N_9006);
nor U14144 (N_14144,N_8990,N_10233);
nand U14145 (N_14145,N_10424,N_11475);
xor U14146 (N_14146,N_11377,N_9825);
xnor U14147 (N_14147,N_10379,N_10300);
and U14148 (N_14148,N_8725,N_10883);
and U14149 (N_14149,N_9357,N_10406);
xor U14150 (N_14150,N_9094,N_10560);
or U14151 (N_14151,N_9720,N_10941);
xor U14152 (N_14152,N_9191,N_8432);
xnor U14153 (N_14153,N_11258,N_11875);
and U14154 (N_14154,N_10160,N_10730);
and U14155 (N_14155,N_11042,N_8510);
or U14156 (N_14156,N_9164,N_8679);
nor U14157 (N_14157,N_8378,N_8173);
and U14158 (N_14158,N_11753,N_10611);
or U14159 (N_14159,N_9396,N_8727);
and U14160 (N_14160,N_8610,N_9387);
xnor U14161 (N_14161,N_8297,N_9987);
or U14162 (N_14162,N_11084,N_9512);
or U14163 (N_14163,N_8211,N_8821);
nor U14164 (N_14164,N_8214,N_11641);
nand U14165 (N_14165,N_10977,N_10676);
or U14166 (N_14166,N_8326,N_11442);
xnor U14167 (N_14167,N_9524,N_8927);
or U14168 (N_14168,N_11883,N_10748);
nand U14169 (N_14169,N_11338,N_8643);
or U14170 (N_14170,N_9438,N_10373);
nor U14171 (N_14171,N_10554,N_9930);
nor U14172 (N_14172,N_11721,N_11383);
nor U14173 (N_14173,N_11404,N_10086);
nand U14174 (N_14174,N_11920,N_8985);
nor U14175 (N_14175,N_8321,N_8018);
nand U14176 (N_14176,N_11201,N_9246);
or U14177 (N_14177,N_10113,N_8466);
xnor U14178 (N_14178,N_11115,N_11006);
and U14179 (N_14179,N_9400,N_9915);
nor U14180 (N_14180,N_10960,N_10940);
and U14181 (N_14181,N_11418,N_9744);
nand U14182 (N_14182,N_10651,N_10965);
nor U14183 (N_14183,N_10226,N_9166);
nand U14184 (N_14184,N_11456,N_11120);
or U14185 (N_14185,N_9805,N_8406);
xnor U14186 (N_14186,N_10880,N_8481);
xnor U14187 (N_14187,N_8811,N_8662);
and U14188 (N_14188,N_11534,N_9924);
nand U14189 (N_14189,N_11133,N_11184);
nand U14190 (N_14190,N_9227,N_11370);
xnor U14191 (N_14191,N_9197,N_10823);
and U14192 (N_14192,N_9913,N_11197);
nor U14193 (N_14193,N_10095,N_8368);
xnor U14194 (N_14194,N_11584,N_9190);
and U14195 (N_14195,N_8130,N_8525);
xor U14196 (N_14196,N_11713,N_10555);
xnor U14197 (N_14197,N_11029,N_11578);
and U14198 (N_14198,N_10613,N_10931);
xor U14199 (N_14199,N_10646,N_8542);
nand U14200 (N_14200,N_9568,N_11661);
and U14201 (N_14201,N_11789,N_10082);
nand U14202 (N_14202,N_11093,N_11095);
or U14203 (N_14203,N_10097,N_11683);
nor U14204 (N_14204,N_11094,N_10676);
xnor U14205 (N_14205,N_11084,N_8655);
and U14206 (N_14206,N_11136,N_11309);
nor U14207 (N_14207,N_11449,N_11070);
nor U14208 (N_14208,N_9603,N_10527);
xor U14209 (N_14209,N_8365,N_8209);
xor U14210 (N_14210,N_9394,N_11686);
or U14211 (N_14211,N_8844,N_11991);
and U14212 (N_14212,N_8669,N_9351);
nand U14213 (N_14213,N_11013,N_9914);
or U14214 (N_14214,N_11616,N_11025);
nor U14215 (N_14215,N_11027,N_10514);
and U14216 (N_14216,N_9178,N_9314);
xor U14217 (N_14217,N_8590,N_11351);
or U14218 (N_14218,N_9956,N_10996);
xnor U14219 (N_14219,N_8513,N_10252);
xor U14220 (N_14220,N_9332,N_8010);
nor U14221 (N_14221,N_10495,N_9000);
xor U14222 (N_14222,N_10486,N_8205);
nand U14223 (N_14223,N_8136,N_11833);
nor U14224 (N_14224,N_9732,N_11853);
or U14225 (N_14225,N_9971,N_11843);
nand U14226 (N_14226,N_9411,N_10327);
or U14227 (N_14227,N_11977,N_11898);
and U14228 (N_14228,N_10950,N_10913);
xnor U14229 (N_14229,N_9885,N_11550);
xnor U14230 (N_14230,N_8264,N_8195);
and U14231 (N_14231,N_9240,N_11684);
xor U14232 (N_14232,N_11685,N_8516);
xor U14233 (N_14233,N_8543,N_11991);
or U14234 (N_14234,N_10403,N_11406);
nand U14235 (N_14235,N_8144,N_8250);
xor U14236 (N_14236,N_9742,N_8095);
xnor U14237 (N_14237,N_8386,N_8228);
nand U14238 (N_14238,N_9803,N_9435);
nand U14239 (N_14239,N_9618,N_8460);
nor U14240 (N_14240,N_9496,N_11092);
and U14241 (N_14241,N_11561,N_9209);
nand U14242 (N_14242,N_9503,N_10209);
xor U14243 (N_14243,N_10279,N_10069);
xnor U14244 (N_14244,N_8823,N_8216);
xor U14245 (N_14245,N_8226,N_8526);
and U14246 (N_14246,N_10509,N_9143);
nand U14247 (N_14247,N_10041,N_11308);
or U14248 (N_14248,N_8516,N_11469);
and U14249 (N_14249,N_11450,N_9591);
nor U14250 (N_14250,N_9262,N_10444);
xor U14251 (N_14251,N_11469,N_10087);
or U14252 (N_14252,N_10711,N_11065);
and U14253 (N_14253,N_11042,N_10965);
nand U14254 (N_14254,N_10698,N_10604);
or U14255 (N_14255,N_10692,N_9874);
or U14256 (N_14256,N_9572,N_10526);
and U14257 (N_14257,N_9330,N_10981);
xor U14258 (N_14258,N_9951,N_9684);
or U14259 (N_14259,N_9345,N_10416);
nor U14260 (N_14260,N_10270,N_11371);
nand U14261 (N_14261,N_9885,N_10080);
and U14262 (N_14262,N_11923,N_10385);
or U14263 (N_14263,N_10402,N_11214);
and U14264 (N_14264,N_9867,N_8806);
nand U14265 (N_14265,N_9762,N_11976);
or U14266 (N_14266,N_9636,N_9414);
xor U14267 (N_14267,N_10482,N_11213);
xor U14268 (N_14268,N_10336,N_9766);
xnor U14269 (N_14269,N_8867,N_10995);
and U14270 (N_14270,N_11292,N_11197);
and U14271 (N_14271,N_8520,N_11590);
nand U14272 (N_14272,N_11696,N_10929);
xor U14273 (N_14273,N_11178,N_11944);
or U14274 (N_14274,N_10285,N_9018);
nand U14275 (N_14275,N_8573,N_11580);
or U14276 (N_14276,N_8377,N_9706);
xnor U14277 (N_14277,N_11930,N_8224);
or U14278 (N_14278,N_11234,N_11523);
nand U14279 (N_14279,N_8532,N_11061);
and U14280 (N_14280,N_11436,N_8119);
and U14281 (N_14281,N_8305,N_8864);
nor U14282 (N_14282,N_8691,N_9360);
xor U14283 (N_14283,N_9310,N_10431);
or U14284 (N_14284,N_8938,N_10473);
and U14285 (N_14285,N_9768,N_11509);
nand U14286 (N_14286,N_10788,N_10354);
nand U14287 (N_14287,N_8518,N_11299);
and U14288 (N_14288,N_11112,N_11959);
nand U14289 (N_14289,N_8850,N_9715);
xnor U14290 (N_14290,N_9784,N_10127);
or U14291 (N_14291,N_11933,N_10097);
or U14292 (N_14292,N_9290,N_11046);
nor U14293 (N_14293,N_11090,N_8904);
and U14294 (N_14294,N_8453,N_11936);
nand U14295 (N_14295,N_9061,N_11941);
xnor U14296 (N_14296,N_11120,N_11003);
or U14297 (N_14297,N_10851,N_8627);
and U14298 (N_14298,N_9853,N_11596);
nand U14299 (N_14299,N_11738,N_9280);
nor U14300 (N_14300,N_8705,N_10955);
xor U14301 (N_14301,N_10333,N_8535);
nor U14302 (N_14302,N_10182,N_11713);
nand U14303 (N_14303,N_8167,N_8180);
or U14304 (N_14304,N_11676,N_9773);
xnor U14305 (N_14305,N_8976,N_10216);
nor U14306 (N_14306,N_9034,N_9609);
xnor U14307 (N_14307,N_8280,N_9431);
and U14308 (N_14308,N_11325,N_9098);
or U14309 (N_14309,N_10987,N_9532);
nand U14310 (N_14310,N_8242,N_9343);
nor U14311 (N_14311,N_10577,N_11864);
or U14312 (N_14312,N_9785,N_11193);
xnor U14313 (N_14313,N_9962,N_9087);
or U14314 (N_14314,N_8461,N_9956);
or U14315 (N_14315,N_8643,N_8604);
and U14316 (N_14316,N_8982,N_11178);
xnor U14317 (N_14317,N_9617,N_8935);
nor U14318 (N_14318,N_8930,N_10927);
and U14319 (N_14319,N_10368,N_11470);
or U14320 (N_14320,N_11123,N_11948);
or U14321 (N_14321,N_9315,N_8082);
nand U14322 (N_14322,N_9921,N_9560);
or U14323 (N_14323,N_10759,N_11800);
and U14324 (N_14324,N_11960,N_9956);
nor U14325 (N_14325,N_8692,N_10205);
and U14326 (N_14326,N_10644,N_11229);
and U14327 (N_14327,N_8071,N_9871);
or U14328 (N_14328,N_11010,N_9008);
xnor U14329 (N_14329,N_9247,N_10190);
or U14330 (N_14330,N_9539,N_10462);
xor U14331 (N_14331,N_11792,N_8014);
nor U14332 (N_14332,N_8593,N_9574);
and U14333 (N_14333,N_9773,N_11311);
or U14334 (N_14334,N_11041,N_11475);
nor U14335 (N_14335,N_10686,N_11718);
nor U14336 (N_14336,N_9798,N_8197);
nor U14337 (N_14337,N_8239,N_11310);
nand U14338 (N_14338,N_9952,N_9841);
nand U14339 (N_14339,N_9018,N_9226);
xor U14340 (N_14340,N_11442,N_10567);
nor U14341 (N_14341,N_8085,N_11625);
and U14342 (N_14342,N_8158,N_8243);
or U14343 (N_14343,N_11087,N_11259);
xor U14344 (N_14344,N_9020,N_11514);
or U14345 (N_14345,N_10307,N_8435);
nand U14346 (N_14346,N_8314,N_11775);
xor U14347 (N_14347,N_9292,N_9660);
and U14348 (N_14348,N_10943,N_9422);
and U14349 (N_14349,N_10434,N_9507);
and U14350 (N_14350,N_11182,N_10040);
and U14351 (N_14351,N_8802,N_9395);
nor U14352 (N_14352,N_8884,N_9304);
xor U14353 (N_14353,N_8917,N_9427);
nand U14354 (N_14354,N_9407,N_10383);
nor U14355 (N_14355,N_9736,N_11730);
and U14356 (N_14356,N_10382,N_11215);
or U14357 (N_14357,N_9901,N_8380);
and U14358 (N_14358,N_10174,N_9431);
and U14359 (N_14359,N_8551,N_10112);
xnor U14360 (N_14360,N_8680,N_8200);
or U14361 (N_14361,N_8814,N_8107);
nor U14362 (N_14362,N_9908,N_9933);
and U14363 (N_14363,N_10420,N_8838);
and U14364 (N_14364,N_9587,N_10956);
nand U14365 (N_14365,N_11049,N_8719);
xor U14366 (N_14366,N_10058,N_8276);
nor U14367 (N_14367,N_11136,N_8183);
nor U14368 (N_14368,N_11186,N_11263);
or U14369 (N_14369,N_10185,N_8286);
nand U14370 (N_14370,N_10560,N_11565);
and U14371 (N_14371,N_8721,N_8167);
or U14372 (N_14372,N_10533,N_9076);
xnor U14373 (N_14373,N_11636,N_8557);
or U14374 (N_14374,N_10475,N_11090);
xnor U14375 (N_14375,N_9814,N_8692);
and U14376 (N_14376,N_8899,N_10563);
nor U14377 (N_14377,N_8198,N_9968);
xor U14378 (N_14378,N_8593,N_8777);
nand U14379 (N_14379,N_10656,N_8145);
xnor U14380 (N_14380,N_11904,N_11284);
nand U14381 (N_14381,N_9569,N_10094);
and U14382 (N_14382,N_10426,N_8167);
or U14383 (N_14383,N_10159,N_10476);
xor U14384 (N_14384,N_11015,N_9161);
and U14385 (N_14385,N_10795,N_8256);
nand U14386 (N_14386,N_8390,N_10308);
or U14387 (N_14387,N_11049,N_10118);
nor U14388 (N_14388,N_10835,N_8767);
and U14389 (N_14389,N_9160,N_11385);
and U14390 (N_14390,N_11272,N_8271);
or U14391 (N_14391,N_8758,N_10819);
and U14392 (N_14392,N_11152,N_10709);
nor U14393 (N_14393,N_11618,N_10185);
nand U14394 (N_14394,N_8941,N_8066);
nor U14395 (N_14395,N_11719,N_9693);
nor U14396 (N_14396,N_9101,N_8011);
nand U14397 (N_14397,N_9331,N_9490);
nand U14398 (N_14398,N_11149,N_9719);
nor U14399 (N_14399,N_10414,N_9592);
and U14400 (N_14400,N_10051,N_8909);
xor U14401 (N_14401,N_9023,N_8883);
or U14402 (N_14402,N_11184,N_10235);
xnor U14403 (N_14403,N_11792,N_8977);
and U14404 (N_14404,N_9965,N_9108);
xor U14405 (N_14405,N_10297,N_9191);
and U14406 (N_14406,N_9594,N_10854);
nor U14407 (N_14407,N_11791,N_8347);
nand U14408 (N_14408,N_9077,N_11701);
nand U14409 (N_14409,N_10971,N_9304);
nand U14410 (N_14410,N_8711,N_8316);
nand U14411 (N_14411,N_8126,N_8353);
nor U14412 (N_14412,N_8619,N_10582);
xnor U14413 (N_14413,N_9355,N_11716);
or U14414 (N_14414,N_8046,N_11867);
nor U14415 (N_14415,N_8121,N_11615);
and U14416 (N_14416,N_10065,N_8107);
and U14417 (N_14417,N_11873,N_8877);
nor U14418 (N_14418,N_9210,N_8219);
or U14419 (N_14419,N_9993,N_10046);
or U14420 (N_14420,N_10749,N_10396);
or U14421 (N_14421,N_8900,N_10585);
and U14422 (N_14422,N_10459,N_10998);
and U14423 (N_14423,N_9397,N_11350);
nor U14424 (N_14424,N_9062,N_9605);
or U14425 (N_14425,N_10310,N_8319);
nor U14426 (N_14426,N_9276,N_11504);
nor U14427 (N_14427,N_11717,N_11948);
and U14428 (N_14428,N_8894,N_9006);
nor U14429 (N_14429,N_10213,N_9847);
nand U14430 (N_14430,N_9340,N_9281);
and U14431 (N_14431,N_10012,N_9238);
xnor U14432 (N_14432,N_9470,N_8410);
or U14433 (N_14433,N_10959,N_10196);
or U14434 (N_14434,N_11652,N_9687);
or U14435 (N_14435,N_9669,N_8944);
and U14436 (N_14436,N_8661,N_10184);
xor U14437 (N_14437,N_9540,N_8881);
and U14438 (N_14438,N_10940,N_11667);
nand U14439 (N_14439,N_9821,N_9565);
or U14440 (N_14440,N_11835,N_8600);
xnor U14441 (N_14441,N_10171,N_8518);
nand U14442 (N_14442,N_8498,N_11623);
nand U14443 (N_14443,N_9401,N_8443);
or U14444 (N_14444,N_8505,N_11655);
nor U14445 (N_14445,N_10102,N_10868);
xnor U14446 (N_14446,N_11295,N_10593);
or U14447 (N_14447,N_9448,N_9823);
and U14448 (N_14448,N_10404,N_11662);
and U14449 (N_14449,N_10440,N_10259);
and U14450 (N_14450,N_10220,N_11793);
nor U14451 (N_14451,N_9313,N_8176);
and U14452 (N_14452,N_10698,N_8453);
and U14453 (N_14453,N_8525,N_9495);
nand U14454 (N_14454,N_10224,N_8376);
nand U14455 (N_14455,N_9333,N_11200);
or U14456 (N_14456,N_8182,N_8723);
and U14457 (N_14457,N_10424,N_10890);
or U14458 (N_14458,N_9678,N_9179);
nand U14459 (N_14459,N_10790,N_11447);
xnor U14460 (N_14460,N_8148,N_8371);
nor U14461 (N_14461,N_9272,N_10456);
or U14462 (N_14462,N_10781,N_11193);
nand U14463 (N_14463,N_10778,N_8811);
nand U14464 (N_14464,N_11180,N_10186);
and U14465 (N_14465,N_8367,N_10263);
nor U14466 (N_14466,N_8063,N_10812);
nor U14467 (N_14467,N_10817,N_11092);
or U14468 (N_14468,N_11993,N_10099);
nand U14469 (N_14469,N_10830,N_9979);
xor U14470 (N_14470,N_9104,N_10576);
or U14471 (N_14471,N_10285,N_10332);
xor U14472 (N_14472,N_8479,N_10245);
nand U14473 (N_14473,N_8245,N_10289);
and U14474 (N_14474,N_8120,N_8575);
or U14475 (N_14475,N_11058,N_11548);
nand U14476 (N_14476,N_10040,N_8224);
or U14477 (N_14477,N_11902,N_9495);
and U14478 (N_14478,N_8092,N_9319);
xor U14479 (N_14479,N_9429,N_9536);
nand U14480 (N_14480,N_11994,N_9312);
and U14481 (N_14481,N_9371,N_8034);
and U14482 (N_14482,N_9571,N_11696);
xnor U14483 (N_14483,N_9047,N_10580);
nor U14484 (N_14484,N_9095,N_9282);
or U14485 (N_14485,N_8369,N_10168);
xor U14486 (N_14486,N_9609,N_9510);
xor U14487 (N_14487,N_11394,N_11871);
nand U14488 (N_14488,N_11323,N_9388);
xnor U14489 (N_14489,N_10122,N_10261);
nand U14490 (N_14490,N_8923,N_10447);
and U14491 (N_14491,N_10262,N_11100);
xnor U14492 (N_14492,N_8306,N_10019);
xor U14493 (N_14493,N_11713,N_9712);
nor U14494 (N_14494,N_10468,N_11973);
or U14495 (N_14495,N_8634,N_10946);
or U14496 (N_14496,N_11016,N_9432);
nor U14497 (N_14497,N_8147,N_9745);
or U14498 (N_14498,N_9028,N_9909);
xor U14499 (N_14499,N_8181,N_8614);
xnor U14500 (N_14500,N_8374,N_11224);
nor U14501 (N_14501,N_11414,N_8145);
or U14502 (N_14502,N_11940,N_11601);
xnor U14503 (N_14503,N_10751,N_11703);
xor U14504 (N_14504,N_10175,N_10998);
or U14505 (N_14505,N_8991,N_10826);
xor U14506 (N_14506,N_8262,N_9585);
nor U14507 (N_14507,N_8517,N_10625);
and U14508 (N_14508,N_11984,N_10728);
nand U14509 (N_14509,N_11848,N_11634);
nand U14510 (N_14510,N_10086,N_8351);
nor U14511 (N_14511,N_9029,N_11095);
or U14512 (N_14512,N_11547,N_10493);
and U14513 (N_14513,N_10820,N_9456);
xor U14514 (N_14514,N_10675,N_10358);
xnor U14515 (N_14515,N_9365,N_9848);
xnor U14516 (N_14516,N_8540,N_10360);
xnor U14517 (N_14517,N_9209,N_11627);
nand U14518 (N_14518,N_10330,N_11886);
nor U14519 (N_14519,N_9484,N_9490);
or U14520 (N_14520,N_10805,N_8580);
or U14521 (N_14521,N_11676,N_9961);
nand U14522 (N_14522,N_11659,N_10211);
or U14523 (N_14523,N_8189,N_10435);
nor U14524 (N_14524,N_8085,N_11227);
nand U14525 (N_14525,N_10071,N_9577);
nand U14526 (N_14526,N_9810,N_8570);
or U14527 (N_14527,N_11302,N_9732);
xnor U14528 (N_14528,N_9438,N_11917);
or U14529 (N_14529,N_11943,N_11751);
or U14530 (N_14530,N_8338,N_10695);
nor U14531 (N_14531,N_11215,N_10472);
nand U14532 (N_14532,N_8088,N_8751);
or U14533 (N_14533,N_8083,N_10140);
nand U14534 (N_14534,N_8496,N_8344);
or U14535 (N_14535,N_8675,N_8076);
nand U14536 (N_14536,N_10070,N_8101);
nand U14537 (N_14537,N_10355,N_10059);
nand U14538 (N_14538,N_8185,N_11637);
nor U14539 (N_14539,N_11743,N_10198);
xnor U14540 (N_14540,N_8327,N_10171);
and U14541 (N_14541,N_10635,N_8041);
or U14542 (N_14542,N_11974,N_9195);
nand U14543 (N_14543,N_11138,N_11620);
nand U14544 (N_14544,N_8530,N_8366);
xnor U14545 (N_14545,N_8410,N_10679);
or U14546 (N_14546,N_11007,N_11710);
nand U14547 (N_14547,N_9146,N_11483);
or U14548 (N_14548,N_11871,N_11724);
nand U14549 (N_14549,N_11143,N_9455);
or U14550 (N_14550,N_11048,N_9630);
or U14551 (N_14551,N_8469,N_8461);
or U14552 (N_14552,N_11325,N_10477);
xor U14553 (N_14553,N_9423,N_9816);
nand U14554 (N_14554,N_10871,N_10669);
nor U14555 (N_14555,N_8001,N_11159);
xor U14556 (N_14556,N_8415,N_10784);
xnor U14557 (N_14557,N_11454,N_8657);
and U14558 (N_14558,N_11309,N_10985);
nor U14559 (N_14559,N_8937,N_8232);
nand U14560 (N_14560,N_8941,N_10621);
nand U14561 (N_14561,N_8750,N_9740);
xor U14562 (N_14562,N_8716,N_11780);
nand U14563 (N_14563,N_11345,N_8008);
or U14564 (N_14564,N_8894,N_9364);
or U14565 (N_14565,N_11773,N_8089);
nand U14566 (N_14566,N_11332,N_10237);
and U14567 (N_14567,N_10240,N_8559);
and U14568 (N_14568,N_10620,N_10245);
xor U14569 (N_14569,N_11792,N_8707);
nand U14570 (N_14570,N_9123,N_11975);
nand U14571 (N_14571,N_10229,N_10829);
nor U14572 (N_14572,N_8582,N_8881);
and U14573 (N_14573,N_10910,N_8892);
nand U14574 (N_14574,N_8469,N_8556);
or U14575 (N_14575,N_8508,N_9620);
nor U14576 (N_14576,N_8643,N_11775);
and U14577 (N_14577,N_9921,N_10677);
or U14578 (N_14578,N_11666,N_11918);
or U14579 (N_14579,N_11341,N_9358);
or U14580 (N_14580,N_8507,N_11364);
and U14581 (N_14581,N_10889,N_10776);
nor U14582 (N_14582,N_9783,N_9685);
or U14583 (N_14583,N_11000,N_11279);
nor U14584 (N_14584,N_10143,N_9929);
nor U14585 (N_14585,N_9441,N_11283);
xnor U14586 (N_14586,N_10088,N_9075);
xor U14587 (N_14587,N_11999,N_10654);
or U14588 (N_14588,N_8348,N_11582);
nand U14589 (N_14589,N_10203,N_8138);
nor U14590 (N_14590,N_11013,N_10981);
nand U14591 (N_14591,N_11372,N_11060);
or U14592 (N_14592,N_8311,N_10991);
nand U14593 (N_14593,N_10093,N_8182);
nand U14594 (N_14594,N_11044,N_11081);
nor U14595 (N_14595,N_10625,N_9133);
and U14596 (N_14596,N_10398,N_9520);
xor U14597 (N_14597,N_10738,N_11073);
nand U14598 (N_14598,N_9223,N_8896);
nand U14599 (N_14599,N_8980,N_11854);
nand U14600 (N_14600,N_9662,N_8662);
xnor U14601 (N_14601,N_10614,N_10436);
nand U14602 (N_14602,N_10570,N_10465);
nand U14603 (N_14603,N_10637,N_11972);
nand U14604 (N_14604,N_9706,N_11483);
or U14605 (N_14605,N_9755,N_9199);
or U14606 (N_14606,N_11046,N_9778);
and U14607 (N_14607,N_9236,N_8719);
nor U14608 (N_14608,N_10711,N_9829);
nor U14609 (N_14609,N_10653,N_11156);
xor U14610 (N_14610,N_9084,N_9334);
or U14611 (N_14611,N_8611,N_11857);
and U14612 (N_14612,N_9646,N_10100);
nand U14613 (N_14613,N_10588,N_9821);
or U14614 (N_14614,N_9907,N_8387);
nor U14615 (N_14615,N_9836,N_11740);
nand U14616 (N_14616,N_11989,N_8716);
nand U14617 (N_14617,N_9704,N_9407);
or U14618 (N_14618,N_8434,N_11394);
and U14619 (N_14619,N_11832,N_10372);
nand U14620 (N_14620,N_8286,N_8385);
nand U14621 (N_14621,N_10931,N_10305);
and U14622 (N_14622,N_11065,N_10771);
nand U14623 (N_14623,N_8344,N_9400);
and U14624 (N_14624,N_9373,N_10362);
and U14625 (N_14625,N_9534,N_9169);
xnor U14626 (N_14626,N_11920,N_9248);
nand U14627 (N_14627,N_8377,N_10689);
nor U14628 (N_14628,N_8077,N_11325);
or U14629 (N_14629,N_8341,N_10560);
and U14630 (N_14630,N_8861,N_10740);
or U14631 (N_14631,N_11152,N_10545);
xnor U14632 (N_14632,N_8009,N_11741);
nand U14633 (N_14633,N_10233,N_10983);
and U14634 (N_14634,N_10650,N_8485);
or U14635 (N_14635,N_10204,N_9946);
xnor U14636 (N_14636,N_10407,N_9531);
nor U14637 (N_14637,N_9504,N_10365);
or U14638 (N_14638,N_10423,N_9662);
nand U14639 (N_14639,N_11803,N_11074);
and U14640 (N_14640,N_9421,N_9902);
and U14641 (N_14641,N_11797,N_11595);
xnor U14642 (N_14642,N_10217,N_11061);
nor U14643 (N_14643,N_11765,N_11663);
nor U14644 (N_14644,N_9493,N_10640);
nand U14645 (N_14645,N_11634,N_11615);
and U14646 (N_14646,N_10998,N_9693);
and U14647 (N_14647,N_8327,N_11826);
nand U14648 (N_14648,N_8878,N_11781);
nand U14649 (N_14649,N_8473,N_10734);
xor U14650 (N_14650,N_11639,N_9147);
nand U14651 (N_14651,N_10097,N_9435);
nor U14652 (N_14652,N_8253,N_11117);
nand U14653 (N_14653,N_11569,N_9983);
nor U14654 (N_14654,N_9858,N_8731);
xnor U14655 (N_14655,N_9580,N_9101);
and U14656 (N_14656,N_10974,N_9293);
and U14657 (N_14657,N_9110,N_10416);
nand U14658 (N_14658,N_9217,N_9897);
nor U14659 (N_14659,N_10805,N_9216);
nor U14660 (N_14660,N_11358,N_11753);
xnor U14661 (N_14661,N_11342,N_10360);
nand U14662 (N_14662,N_11807,N_11375);
nand U14663 (N_14663,N_9915,N_8002);
nand U14664 (N_14664,N_10109,N_9118);
nor U14665 (N_14665,N_8024,N_8672);
nand U14666 (N_14666,N_8943,N_8535);
nand U14667 (N_14667,N_10139,N_8989);
or U14668 (N_14668,N_8941,N_8722);
and U14669 (N_14669,N_8604,N_9931);
nor U14670 (N_14670,N_11337,N_9187);
xor U14671 (N_14671,N_9328,N_11520);
nor U14672 (N_14672,N_8625,N_9972);
xnor U14673 (N_14673,N_8182,N_10427);
nor U14674 (N_14674,N_8918,N_9478);
xor U14675 (N_14675,N_10614,N_9115);
or U14676 (N_14676,N_9996,N_11669);
xor U14677 (N_14677,N_10174,N_8179);
nor U14678 (N_14678,N_8520,N_10820);
and U14679 (N_14679,N_11753,N_11958);
nor U14680 (N_14680,N_11340,N_8632);
xnor U14681 (N_14681,N_8310,N_10563);
or U14682 (N_14682,N_11642,N_9425);
nor U14683 (N_14683,N_11984,N_8670);
and U14684 (N_14684,N_10571,N_10825);
nand U14685 (N_14685,N_8611,N_9805);
and U14686 (N_14686,N_10963,N_8678);
or U14687 (N_14687,N_11616,N_8390);
nor U14688 (N_14688,N_9679,N_10249);
xnor U14689 (N_14689,N_8720,N_11784);
xor U14690 (N_14690,N_11000,N_11568);
or U14691 (N_14691,N_10958,N_11388);
xor U14692 (N_14692,N_9054,N_10772);
and U14693 (N_14693,N_11348,N_10874);
xor U14694 (N_14694,N_8074,N_11827);
nand U14695 (N_14695,N_11219,N_8244);
nor U14696 (N_14696,N_11328,N_11653);
nand U14697 (N_14697,N_9977,N_11949);
or U14698 (N_14698,N_10261,N_10364);
nor U14699 (N_14699,N_11218,N_9370);
xor U14700 (N_14700,N_11009,N_11187);
xor U14701 (N_14701,N_9003,N_8741);
or U14702 (N_14702,N_11578,N_8400);
xnor U14703 (N_14703,N_10053,N_10920);
xnor U14704 (N_14704,N_10443,N_10438);
nor U14705 (N_14705,N_11041,N_8942);
xor U14706 (N_14706,N_11869,N_11364);
or U14707 (N_14707,N_10430,N_10737);
xor U14708 (N_14708,N_10470,N_9085);
nor U14709 (N_14709,N_10483,N_8304);
xor U14710 (N_14710,N_9860,N_9597);
or U14711 (N_14711,N_10531,N_8751);
and U14712 (N_14712,N_8309,N_10802);
xnor U14713 (N_14713,N_9090,N_9175);
or U14714 (N_14714,N_10461,N_10800);
or U14715 (N_14715,N_11614,N_11788);
or U14716 (N_14716,N_11674,N_9546);
nand U14717 (N_14717,N_9630,N_10220);
xnor U14718 (N_14718,N_10098,N_10169);
and U14719 (N_14719,N_8468,N_9885);
xor U14720 (N_14720,N_10267,N_9482);
nand U14721 (N_14721,N_10078,N_8728);
or U14722 (N_14722,N_10048,N_9463);
nor U14723 (N_14723,N_9971,N_11769);
nor U14724 (N_14724,N_9556,N_9967);
or U14725 (N_14725,N_10380,N_10231);
xnor U14726 (N_14726,N_10368,N_8791);
xor U14727 (N_14727,N_10301,N_8776);
nand U14728 (N_14728,N_10321,N_8861);
xnor U14729 (N_14729,N_8920,N_10313);
or U14730 (N_14730,N_9667,N_11486);
nand U14731 (N_14731,N_9186,N_8424);
and U14732 (N_14732,N_8173,N_10634);
nor U14733 (N_14733,N_9128,N_10241);
nand U14734 (N_14734,N_10725,N_10797);
xnor U14735 (N_14735,N_11434,N_11773);
or U14736 (N_14736,N_9811,N_11050);
and U14737 (N_14737,N_8391,N_9878);
nand U14738 (N_14738,N_9915,N_8530);
and U14739 (N_14739,N_8410,N_9517);
nor U14740 (N_14740,N_11453,N_8085);
xnor U14741 (N_14741,N_10749,N_10439);
or U14742 (N_14742,N_11970,N_8463);
nand U14743 (N_14743,N_8380,N_9502);
nand U14744 (N_14744,N_8512,N_9322);
or U14745 (N_14745,N_11880,N_8033);
xor U14746 (N_14746,N_8788,N_11480);
xor U14747 (N_14747,N_11835,N_9301);
nand U14748 (N_14748,N_11330,N_8383);
xor U14749 (N_14749,N_8725,N_8778);
nand U14750 (N_14750,N_9213,N_9408);
xor U14751 (N_14751,N_9890,N_9566);
or U14752 (N_14752,N_8741,N_11736);
or U14753 (N_14753,N_11602,N_11832);
and U14754 (N_14754,N_9191,N_10382);
nand U14755 (N_14755,N_11746,N_9527);
or U14756 (N_14756,N_9452,N_10853);
and U14757 (N_14757,N_11531,N_8899);
xnor U14758 (N_14758,N_10185,N_8016);
and U14759 (N_14759,N_10096,N_8772);
xor U14760 (N_14760,N_10896,N_11451);
nor U14761 (N_14761,N_11062,N_8254);
xnor U14762 (N_14762,N_10410,N_11047);
and U14763 (N_14763,N_9277,N_10848);
nor U14764 (N_14764,N_11598,N_9104);
or U14765 (N_14765,N_9930,N_10824);
or U14766 (N_14766,N_8861,N_8463);
or U14767 (N_14767,N_8410,N_11663);
and U14768 (N_14768,N_9295,N_10212);
or U14769 (N_14769,N_9685,N_11889);
or U14770 (N_14770,N_9932,N_11106);
nand U14771 (N_14771,N_10856,N_8039);
nand U14772 (N_14772,N_10021,N_11917);
xor U14773 (N_14773,N_11521,N_8873);
nand U14774 (N_14774,N_11956,N_8867);
and U14775 (N_14775,N_10762,N_10698);
nor U14776 (N_14776,N_8078,N_8321);
nor U14777 (N_14777,N_9880,N_8145);
and U14778 (N_14778,N_11908,N_10175);
nand U14779 (N_14779,N_11833,N_11771);
nand U14780 (N_14780,N_8722,N_10976);
xor U14781 (N_14781,N_10855,N_10184);
nor U14782 (N_14782,N_8939,N_10522);
nand U14783 (N_14783,N_8849,N_9853);
and U14784 (N_14784,N_9432,N_10153);
nand U14785 (N_14785,N_11277,N_11528);
or U14786 (N_14786,N_11567,N_9839);
nor U14787 (N_14787,N_11217,N_10148);
xnor U14788 (N_14788,N_11225,N_9550);
and U14789 (N_14789,N_10710,N_11955);
nor U14790 (N_14790,N_8797,N_8001);
xor U14791 (N_14791,N_10792,N_11677);
and U14792 (N_14792,N_10753,N_9195);
xor U14793 (N_14793,N_10540,N_11306);
and U14794 (N_14794,N_10138,N_11314);
xnor U14795 (N_14795,N_9105,N_9502);
xnor U14796 (N_14796,N_11254,N_8267);
nor U14797 (N_14797,N_8221,N_11389);
nor U14798 (N_14798,N_10454,N_11858);
and U14799 (N_14799,N_9319,N_10784);
and U14800 (N_14800,N_10902,N_10766);
or U14801 (N_14801,N_11991,N_8678);
xnor U14802 (N_14802,N_11206,N_9780);
nand U14803 (N_14803,N_9005,N_10917);
nor U14804 (N_14804,N_10321,N_10327);
xnor U14805 (N_14805,N_9741,N_11790);
or U14806 (N_14806,N_8721,N_9085);
and U14807 (N_14807,N_10681,N_10767);
xor U14808 (N_14808,N_11418,N_8084);
nor U14809 (N_14809,N_10324,N_8387);
nor U14810 (N_14810,N_9376,N_8051);
xor U14811 (N_14811,N_11804,N_11165);
or U14812 (N_14812,N_10526,N_8834);
nand U14813 (N_14813,N_8073,N_8349);
nor U14814 (N_14814,N_8023,N_10043);
nor U14815 (N_14815,N_11255,N_11615);
nor U14816 (N_14816,N_8817,N_11701);
nand U14817 (N_14817,N_9663,N_11305);
or U14818 (N_14818,N_11069,N_10327);
nand U14819 (N_14819,N_9151,N_11319);
xnor U14820 (N_14820,N_8931,N_9167);
or U14821 (N_14821,N_8944,N_9951);
nor U14822 (N_14822,N_9635,N_10176);
nor U14823 (N_14823,N_9588,N_11112);
xnor U14824 (N_14824,N_9164,N_9182);
or U14825 (N_14825,N_10181,N_10168);
or U14826 (N_14826,N_9034,N_11568);
or U14827 (N_14827,N_10444,N_10254);
nand U14828 (N_14828,N_10297,N_9292);
xnor U14829 (N_14829,N_8450,N_11322);
xor U14830 (N_14830,N_11056,N_9690);
and U14831 (N_14831,N_9723,N_8585);
nand U14832 (N_14832,N_10428,N_8850);
nor U14833 (N_14833,N_9630,N_9078);
and U14834 (N_14834,N_8592,N_9779);
xor U14835 (N_14835,N_9324,N_10762);
xor U14836 (N_14836,N_8255,N_9481);
and U14837 (N_14837,N_8398,N_11754);
nand U14838 (N_14838,N_11992,N_9023);
nor U14839 (N_14839,N_9181,N_10779);
nand U14840 (N_14840,N_9024,N_8624);
nor U14841 (N_14841,N_8279,N_8889);
nor U14842 (N_14842,N_10674,N_8174);
and U14843 (N_14843,N_8177,N_10824);
nor U14844 (N_14844,N_8739,N_11434);
and U14845 (N_14845,N_8841,N_9797);
or U14846 (N_14846,N_8967,N_10456);
xor U14847 (N_14847,N_8556,N_8918);
nor U14848 (N_14848,N_10808,N_11733);
and U14849 (N_14849,N_9821,N_10415);
nor U14850 (N_14850,N_10311,N_11861);
and U14851 (N_14851,N_10804,N_10679);
xnor U14852 (N_14852,N_10863,N_11621);
xnor U14853 (N_14853,N_11747,N_11118);
and U14854 (N_14854,N_11985,N_9611);
xnor U14855 (N_14855,N_10963,N_8033);
nand U14856 (N_14856,N_10131,N_11987);
nand U14857 (N_14857,N_9666,N_8938);
xnor U14858 (N_14858,N_8300,N_9628);
xor U14859 (N_14859,N_10623,N_11030);
xor U14860 (N_14860,N_9890,N_11479);
and U14861 (N_14861,N_9336,N_8456);
nor U14862 (N_14862,N_10384,N_9156);
nor U14863 (N_14863,N_11180,N_9128);
and U14864 (N_14864,N_11484,N_11114);
nor U14865 (N_14865,N_10214,N_11892);
nand U14866 (N_14866,N_9333,N_10081);
nor U14867 (N_14867,N_11080,N_10520);
xnor U14868 (N_14868,N_11881,N_11489);
or U14869 (N_14869,N_10365,N_11952);
xnor U14870 (N_14870,N_10871,N_8951);
nand U14871 (N_14871,N_11628,N_9297);
nor U14872 (N_14872,N_8717,N_9307);
nor U14873 (N_14873,N_11134,N_11497);
or U14874 (N_14874,N_10493,N_11227);
nand U14875 (N_14875,N_8832,N_10276);
and U14876 (N_14876,N_10586,N_9000);
nor U14877 (N_14877,N_11452,N_8318);
xnor U14878 (N_14878,N_9588,N_9080);
and U14879 (N_14879,N_9671,N_9097);
and U14880 (N_14880,N_9011,N_11245);
and U14881 (N_14881,N_9349,N_9493);
nand U14882 (N_14882,N_9872,N_11009);
nand U14883 (N_14883,N_9517,N_11195);
nor U14884 (N_14884,N_9310,N_10537);
xor U14885 (N_14885,N_10922,N_11279);
nor U14886 (N_14886,N_8319,N_10934);
xor U14887 (N_14887,N_10015,N_10038);
xor U14888 (N_14888,N_8941,N_9858);
or U14889 (N_14889,N_8887,N_8936);
or U14890 (N_14890,N_10136,N_9960);
xnor U14891 (N_14891,N_11726,N_11950);
xor U14892 (N_14892,N_11752,N_9880);
and U14893 (N_14893,N_10629,N_10218);
and U14894 (N_14894,N_8031,N_8068);
nand U14895 (N_14895,N_11615,N_8455);
nor U14896 (N_14896,N_9382,N_11640);
nand U14897 (N_14897,N_8300,N_11825);
or U14898 (N_14898,N_11715,N_10493);
nor U14899 (N_14899,N_10184,N_9125);
xor U14900 (N_14900,N_8550,N_9624);
and U14901 (N_14901,N_8903,N_9232);
nand U14902 (N_14902,N_11130,N_8960);
xor U14903 (N_14903,N_10400,N_9149);
xnor U14904 (N_14904,N_9247,N_9889);
nand U14905 (N_14905,N_11471,N_11557);
nand U14906 (N_14906,N_11566,N_11890);
xnor U14907 (N_14907,N_8716,N_10836);
and U14908 (N_14908,N_11455,N_8350);
nand U14909 (N_14909,N_11580,N_8263);
or U14910 (N_14910,N_9487,N_8650);
or U14911 (N_14911,N_11498,N_9625);
nand U14912 (N_14912,N_8577,N_9598);
xor U14913 (N_14913,N_10438,N_10100);
nand U14914 (N_14914,N_11048,N_11490);
nand U14915 (N_14915,N_11200,N_9129);
xnor U14916 (N_14916,N_8432,N_9023);
and U14917 (N_14917,N_11537,N_9101);
nor U14918 (N_14918,N_9766,N_11490);
nand U14919 (N_14919,N_10252,N_10125);
and U14920 (N_14920,N_8210,N_11986);
and U14921 (N_14921,N_11378,N_8207);
nor U14922 (N_14922,N_10165,N_10019);
xor U14923 (N_14923,N_10576,N_9680);
xor U14924 (N_14924,N_9353,N_8996);
or U14925 (N_14925,N_8948,N_10805);
xnor U14926 (N_14926,N_8266,N_10690);
or U14927 (N_14927,N_8140,N_9371);
nand U14928 (N_14928,N_9463,N_10428);
or U14929 (N_14929,N_9149,N_11922);
nor U14930 (N_14930,N_10105,N_9727);
xor U14931 (N_14931,N_8868,N_9257);
nor U14932 (N_14932,N_8713,N_8458);
or U14933 (N_14933,N_11788,N_9535);
xor U14934 (N_14934,N_9699,N_9338);
xor U14935 (N_14935,N_10006,N_10627);
xnor U14936 (N_14936,N_10710,N_10395);
xnor U14937 (N_14937,N_9774,N_8310);
or U14938 (N_14938,N_8824,N_8104);
and U14939 (N_14939,N_9541,N_8992);
or U14940 (N_14940,N_9894,N_10309);
and U14941 (N_14941,N_8538,N_11044);
nand U14942 (N_14942,N_11367,N_9095);
and U14943 (N_14943,N_10967,N_11044);
xor U14944 (N_14944,N_11774,N_11399);
nor U14945 (N_14945,N_11139,N_9905);
or U14946 (N_14946,N_11005,N_11976);
nor U14947 (N_14947,N_8218,N_9101);
nor U14948 (N_14948,N_9517,N_8532);
nor U14949 (N_14949,N_9605,N_8429);
xor U14950 (N_14950,N_9848,N_9517);
nand U14951 (N_14951,N_11230,N_9443);
or U14952 (N_14952,N_10019,N_10907);
xnor U14953 (N_14953,N_9473,N_10875);
xnor U14954 (N_14954,N_10271,N_10891);
and U14955 (N_14955,N_9527,N_9368);
xor U14956 (N_14956,N_8642,N_9036);
and U14957 (N_14957,N_8242,N_10030);
or U14958 (N_14958,N_11792,N_8030);
or U14959 (N_14959,N_10977,N_8403);
or U14960 (N_14960,N_11913,N_11715);
nand U14961 (N_14961,N_8103,N_11233);
xor U14962 (N_14962,N_9771,N_8698);
xnor U14963 (N_14963,N_9758,N_11262);
nand U14964 (N_14964,N_11640,N_10239);
nand U14965 (N_14965,N_9463,N_9678);
or U14966 (N_14966,N_11263,N_9463);
nor U14967 (N_14967,N_8454,N_8822);
nor U14968 (N_14968,N_8324,N_8325);
and U14969 (N_14969,N_11148,N_11428);
and U14970 (N_14970,N_8854,N_9212);
or U14971 (N_14971,N_11316,N_8346);
xor U14972 (N_14972,N_8288,N_11946);
nand U14973 (N_14973,N_9764,N_9419);
nor U14974 (N_14974,N_10767,N_10920);
and U14975 (N_14975,N_10739,N_10735);
nor U14976 (N_14976,N_8468,N_9761);
nand U14977 (N_14977,N_9889,N_11855);
nand U14978 (N_14978,N_11616,N_10057);
nor U14979 (N_14979,N_8857,N_9556);
xor U14980 (N_14980,N_11163,N_9120);
nor U14981 (N_14981,N_11737,N_10524);
nand U14982 (N_14982,N_8160,N_8679);
and U14983 (N_14983,N_10059,N_11608);
xor U14984 (N_14984,N_9328,N_8336);
and U14985 (N_14985,N_11529,N_8216);
xnor U14986 (N_14986,N_9344,N_9224);
and U14987 (N_14987,N_10954,N_10668);
and U14988 (N_14988,N_8294,N_11415);
nor U14989 (N_14989,N_11502,N_8351);
xnor U14990 (N_14990,N_11996,N_10451);
nand U14991 (N_14991,N_9258,N_8867);
nor U14992 (N_14992,N_10548,N_10285);
nand U14993 (N_14993,N_10029,N_10901);
nor U14994 (N_14994,N_9685,N_8605);
nand U14995 (N_14995,N_11986,N_8623);
nor U14996 (N_14996,N_10669,N_10097);
xor U14997 (N_14997,N_9330,N_11478);
nand U14998 (N_14998,N_9528,N_9948);
xor U14999 (N_14999,N_11006,N_8806);
and U15000 (N_15000,N_10957,N_10460);
nor U15001 (N_15001,N_8264,N_9339);
xnor U15002 (N_15002,N_11722,N_8255);
xor U15003 (N_15003,N_8378,N_10865);
or U15004 (N_15004,N_9360,N_8041);
nand U15005 (N_15005,N_8556,N_9324);
or U15006 (N_15006,N_10618,N_8707);
and U15007 (N_15007,N_10850,N_9796);
nor U15008 (N_15008,N_8214,N_9156);
xnor U15009 (N_15009,N_11048,N_8768);
or U15010 (N_15010,N_10563,N_9321);
xnor U15011 (N_15011,N_8861,N_11415);
or U15012 (N_15012,N_9144,N_9311);
nor U15013 (N_15013,N_8711,N_11717);
and U15014 (N_15014,N_9104,N_10675);
or U15015 (N_15015,N_11102,N_9747);
nor U15016 (N_15016,N_11642,N_10821);
or U15017 (N_15017,N_11355,N_10868);
xnor U15018 (N_15018,N_8593,N_11917);
nor U15019 (N_15019,N_9703,N_9906);
nor U15020 (N_15020,N_10265,N_9052);
nand U15021 (N_15021,N_9407,N_8991);
nor U15022 (N_15022,N_8209,N_8046);
xor U15023 (N_15023,N_11698,N_8651);
and U15024 (N_15024,N_10524,N_9294);
nand U15025 (N_15025,N_9294,N_9744);
or U15026 (N_15026,N_11950,N_11793);
xnor U15027 (N_15027,N_9924,N_9256);
and U15028 (N_15028,N_9444,N_8947);
nor U15029 (N_15029,N_9833,N_9010);
nand U15030 (N_15030,N_9810,N_11451);
nor U15031 (N_15031,N_9372,N_9822);
nand U15032 (N_15032,N_9935,N_11861);
nand U15033 (N_15033,N_11188,N_11155);
or U15034 (N_15034,N_8317,N_8089);
and U15035 (N_15035,N_11863,N_8248);
xor U15036 (N_15036,N_11299,N_11612);
and U15037 (N_15037,N_11036,N_8530);
or U15038 (N_15038,N_9088,N_9734);
and U15039 (N_15039,N_11429,N_9858);
nand U15040 (N_15040,N_10735,N_11947);
nand U15041 (N_15041,N_9564,N_8373);
nand U15042 (N_15042,N_10429,N_8535);
nor U15043 (N_15043,N_8361,N_8091);
nor U15044 (N_15044,N_8444,N_10325);
xor U15045 (N_15045,N_10718,N_10072);
or U15046 (N_15046,N_10048,N_11575);
and U15047 (N_15047,N_9670,N_8417);
nor U15048 (N_15048,N_11309,N_11524);
nand U15049 (N_15049,N_9309,N_11642);
nor U15050 (N_15050,N_9729,N_10064);
nor U15051 (N_15051,N_8591,N_11193);
or U15052 (N_15052,N_8259,N_11242);
xnor U15053 (N_15053,N_10270,N_9711);
and U15054 (N_15054,N_10775,N_10822);
xor U15055 (N_15055,N_11951,N_9717);
nor U15056 (N_15056,N_9931,N_11293);
xnor U15057 (N_15057,N_8920,N_9605);
nand U15058 (N_15058,N_10746,N_9593);
nor U15059 (N_15059,N_11655,N_10171);
nor U15060 (N_15060,N_11243,N_9418);
and U15061 (N_15061,N_9527,N_8213);
or U15062 (N_15062,N_10622,N_9739);
nor U15063 (N_15063,N_8413,N_9652);
xnor U15064 (N_15064,N_8343,N_8780);
and U15065 (N_15065,N_11176,N_9635);
nand U15066 (N_15066,N_8357,N_8319);
xnor U15067 (N_15067,N_9229,N_8931);
or U15068 (N_15068,N_9465,N_11032);
xnor U15069 (N_15069,N_9842,N_8391);
nor U15070 (N_15070,N_9589,N_8631);
and U15071 (N_15071,N_9669,N_9065);
or U15072 (N_15072,N_10610,N_8284);
xor U15073 (N_15073,N_8655,N_9392);
nor U15074 (N_15074,N_11730,N_10517);
nand U15075 (N_15075,N_9804,N_9011);
nor U15076 (N_15076,N_11628,N_11414);
or U15077 (N_15077,N_10453,N_11390);
nand U15078 (N_15078,N_9928,N_9658);
xor U15079 (N_15079,N_11800,N_8811);
and U15080 (N_15080,N_11284,N_9044);
xnor U15081 (N_15081,N_8923,N_9860);
and U15082 (N_15082,N_10529,N_10784);
nand U15083 (N_15083,N_11658,N_8546);
or U15084 (N_15084,N_8156,N_11013);
nor U15085 (N_15085,N_10227,N_10107);
nand U15086 (N_15086,N_9145,N_10439);
nor U15087 (N_15087,N_9225,N_10680);
xor U15088 (N_15088,N_8148,N_9874);
nor U15089 (N_15089,N_8086,N_8848);
nor U15090 (N_15090,N_8581,N_8792);
nand U15091 (N_15091,N_9363,N_8959);
or U15092 (N_15092,N_9949,N_9248);
xor U15093 (N_15093,N_11002,N_9662);
or U15094 (N_15094,N_9295,N_8031);
nor U15095 (N_15095,N_10905,N_11798);
xor U15096 (N_15096,N_8983,N_8554);
xor U15097 (N_15097,N_9365,N_10146);
nor U15098 (N_15098,N_8909,N_8446);
xnor U15099 (N_15099,N_10907,N_10791);
nand U15100 (N_15100,N_9561,N_11534);
and U15101 (N_15101,N_8405,N_11704);
nor U15102 (N_15102,N_9568,N_10223);
nor U15103 (N_15103,N_8433,N_11560);
and U15104 (N_15104,N_8533,N_9521);
nor U15105 (N_15105,N_8219,N_10041);
and U15106 (N_15106,N_9924,N_9679);
or U15107 (N_15107,N_8110,N_11983);
nor U15108 (N_15108,N_11439,N_9499);
and U15109 (N_15109,N_10695,N_10966);
or U15110 (N_15110,N_8372,N_9285);
and U15111 (N_15111,N_8800,N_8651);
or U15112 (N_15112,N_8900,N_10263);
or U15113 (N_15113,N_10883,N_10813);
xor U15114 (N_15114,N_11369,N_11530);
nor U15115 (N_15115,N_11612,N_11763);
and U15116 (N_15116,N_10654,N_9594);
nand U15117 (N_15117,N_8074,N_8422);
or U15118 (N_15118,N_9522,N_9933);
and U15119 (N_15119,N_8611,N_8168);
and U15120 (N_15120,N_8144,N_11171);
nor U15121 (N_15121,N_11172,N_9230);
nor U15122 (N_15122,N_9064,N_8719);
or U15123 (N_15123,N_8376,N_10751);
xor U15124 (N_15124,N_8258,N_9840);
and U15125 (N_15125,N_8822,N_10895);
nor U15126 (N_15126,N_10338,N_10499);
xnor U15127 (N_15127,N_11441,N_10506);
nand U15128 (N_15128,N_10063,N_8730);
and U15129 (N_15129,N_11816,N_8174);
nand U15130 (N_15130,N_10740,N_10354);
xor U15131 (N_15131,N_9630,N_9697);
nor U15132 (N_15132,N_9013,N_10854);
nand U15133 (N_15133,N_10827,N_8196);
nand U15134 (N_15134,N_9913,N_9057);
and U15135 (N_15135,N_11672,N_11813);
or U15136 (N_15136,N_9908,N_9215);
and U15137 (N_15137,N_9392,N_11064);
nor U15138 (N_15138,N_11851,N_11746);
and U15139 (N_15139,N_8018,N_8717);
and U15140 (N_15140,N_8885,N_10119);
nor U15141 (N_15141,N_10902,N_8632);
nor U15142 (N_15142,N_9424,N_8791);
nor U15143 (N_15143,N_10670,N_9231);
xnor U15144 (N_15144,N_10931,N_9399);
and U15145 (N_15145,N_9027,N_11840);
and U15146 (N_15146,N_10707,N_9370);
nor U15147 (N_15147,N_10780,N_9407);
or U15148 (N_15148,N_9517,N_8794);
xor U15149 (N_15149,N_11601,N_10052);
xor U15150 (N_15150,N_10056,N_8261);
xnor U15151 (N_15151,N_9714,N_10530);
nor U15152 (N_15152,N_11550,N_11812);
or U15153 (N_15153,N_10253,N_10099);
or U15154 (N_15154,N_8519,N_9087);
nand U15155 (N_15155,N_8543,N_9000);
nor U15156 (N_15156,N_8844,N_8687);
xor U15157 (N_15157,N_9448,N_8897);
nand U15158 (N_15158,N_11469,N_8180);
nor U15159 (N_15159,N_9304,N_9806);
or U15160 (N_15160,N_10886,N_8346);
or U15161 (N_15161,N_8066,N_11766);
nor U15162 (N_15162,N_11827,N_8036);
xnor U15163 (N_15163,N_9336,N_11069);
or U15164 (N_15164,N_10673,N_8167);
and U15165 (N_15165,N_8741,N_11101);
nand U15166 (N_15166,N_8887,N_8399);
and U15167 (N_15167,N_11028,N_9439);
nand U15168 (N_15168,N_11405,N_11247);
or U15169 (N_15169,N_10721,N_11653);
or U15170 (N_15170,N_9064,N_8452);
or U15171 (N_15171,N_9664,N_8572);
nand U15172 (N_15172,N_11549,N_8504);
xor U15173 (N_15173,N_11713,N_8395);
and U15174 (N_15174,N_11641,N_10103);
or U15175 (N_15175,N_8863,N_8816);
and U15176 (N_15176,N_10438,N_11264);
nand U15177 (N_15177,N_11221,N_11544);
and U15178 (N_15178,N_11716,N_11509);
nand U15179 (N_15179,N_10486,N_10562);
and U15180 (N_15180,N_10578,N_8296);
or U15181 (N_15181,N_11536,N_9662);
xnor U15182 (N_15182,N_10720,N_9202);
nand U15183 (N_15183,N_8711,N_10789);
and U15184 (N_15184,N_11014,N_11767);
and U15185 (N_15185,N_11278,N_11120);
and U15186 (N_15186,N_10059,N_9274);
or U15187 (N_15187,N_9682,N_8735);
nor U15188 (N_15188,N_10390,N_9499);
and U15189 (N_15189,N_9637,N_11839);
or U15190 (N_15190,N_8648,N_11128);
xnor U15191 (N_15191,N_9125,N_11098);
or U15192 (N_15192,N_10402,N_8888);
and U15193 (N_15193,N_8624,N_8867);
or U15194 (N_15194,N_9277,N_11267);
xnor U15195 (N_15195,N_8161,N_8136);
or U15196 (N_15196,N_10955,N_8935);
xnor U15197 (N_15197,N_8286,N_9928);
xnor U15198 (N_15198,N_8051,N_11162);
nand U15199 (N_15199,N_9566,N_10932);
or U15200 (N_15200,N_11483,N_11489);
nor U15201 (N_15201,N_11185,N_8509);
nor U15202 (N_15202,N_9088,N_9066);
and U15203 (N_15203,N_11068,N_8725);
or U15204 (N_15204,N_8474,N_10430);
or U15205 (N_15205,N_8478,N_8505);
nand U15206 (N_15206,N_8717,N_11869);
nand U15207 (N_15207,N_9697,N_10520);
or U15208 (N_15208,N_8964,N_10412);
xor U15209 (N_15209,N_9574,N_11301);
and U15210 (N_15210,N_10990,N_11178);
nor U15211 (N_15211,N_11639,N_10120);
or U15212 (N_15212,N_10148,N_10646);
nor U15213 (N_15213,N_11621,N_9634);
xnor U15214 (N_15214,N_9006,N_10888);
nor U15215 (N_15215,N_11120,N_9580);
or U15216 (N_15216,N_10741,N_10940);
nand U15217 (N_15217,N_9049,N_8901);
nand U15218 (N_15218,N_8894,N_9126);
or U15219 (N_15219,N_11200,N_9140);
xor U15220 (N_15220,N_9545,N_11090);
nand U15221 (N_15221,N_8313,N_10609);
xor U15222 (N_15222,N_11979,N_10546);
nand U15223 (N_15223,N_11948,N_8632);
xor U15224 (N_15224,N_11978,N_8668);
nand U15225 (N_15225,N_9402,N_11242);
nand U15226 (N_15226,N_8768,N_8561);
and U15227 (N_15227,N_9103,N_9796);
nand U15228 (N_15228,N_10345,N_10996);
xor U15229 (N_15229,N_8967,N_8063);
nor U15230 (N_15230,N_8391,N_8907);
xnor U15231 (N_15231,N_11475,N_10066);
nand U15232 (N_15232,N_8686,N_10616);
nand U15233 (N_15233,N_10591,N_9638);
nand U15234 (N_15234,N_8068,N_10034);
or U15235 (N_15235,N_8106,N_10739);
xnor U15236 (N_15236,N_11549,N_8351);
nor U15237 (N_15237,N_8128,N_10334);
and U15238 (N_15238,N_11942,N_11797);
or U15239 (N_15239,N_9146,N_11645);
and U15240 (N_15240,N_9237,N_11783);
nor U15241 (N_15241,N_11172,N_8637);
or U15242 (N_15242,N_11688,N_8249);
nand U15243 (N_15243,N_10055,N_9715);
and U15244 (N_15244,N_11213,N_9893);
and U15245 (N_15245,N_11250,N_11043);
nor U15246 (N_15246,N_8657,N_9155);
or U15247 (N_15247,N_11575,N_11372);
or U15248 (N_15248,N_11451,N_10859);
nand U15249 (N_15249,N_10223,N_11001);
nand U15250 (N_15250,N_9043,N_11860);
and U15251 (N_15251,N_8478,N_9053);
nor U15252 (N_15252,N_9134,N_11091);
or U15253 (N_15253,N_10773,N_8426);
or U15254 (N_15254,N_8777,N_11308);
nand U15255 (N_15255,N_10617,N_9400);
and U15256 (N_15256,N_10065,N_9400);
and U15257 (N_15257,N_8111,N_11157);
nand U15258 (N_15258,N_8309,N_11867);
and U15259 (N_15259,N_10364,N_11931);
xor U15260 (N_15260,N_10068,N_8849);
or U15261 (N_15261,N_11327,N_8249);
or U15262 (N_15262,N_9401,N_9578);
nor U15263 (N_15263,N_10473,N_9693);
nor U15264 (N_15264,N_10746,N_8086);
xor U15265 (N_15265,N_11809,N_9640);
nor U15266 (N_15266,N_11334,N_11234);
and U15267 (N_15267,N_9535,N_8564);
and U15268 (N_15268,N_11874,N_8511);
nand U15269 (N_15269,N_9752,N_9924);
and U15270 (N_15270,N_8469,N_10004);
and U15271 (N_15271,N_10788,N_10523);
nor U15272 (N_15272,N_10611,N_9639);
xnor U15273 (N_15273,N_8309,N_9472);
and U15274 (N_15274,N_8795,N_10335);
xor U15275 (N_15275,N_11390,N_10669);
and U15276 (N_15276,N_9657,N_10306);
and U15277 (N_15277,N_10493,N_10004);
or U15278 (N_15278,N_10244,N_8552);
and U15279 (N_15279,N_9710,N_10697);
xnor U15280 (N_15280,N_10671,N_11965);
or U15281 (N_15281,N_8855,N_11993);
or U15282 (N_15282,N_10319,N_11066);
xor U15283 (N_15283,N_9729,N_8703);
and U15284 (N_15284,N_11159,N_8526);
nor U15285 (N_15285,N_10259,N_9603);
and U15286 (N_15286,N_9955,N_10738);
nand U15287 (N_15287,N_8607,N_10411);
xor U15288 (N_15288,N_11985,N_10448);
or U15289 (N_15289,N_11130,N_8658);
and U15290 (N_15290,N_9926,N_11622);
nand U15291 (N_15291,N_8310,N_10281);
or U15292 (N_15292,N_9266,N_8907);
and U15293 (N_15293,N_11412,N_9297);
nand U15294 (N_15294,N_11390,N_11092);
and U15295 (N_15295,N_11839,N_11298);
nand U15296 (N_15296,N_8066,N_8042);
or U15297 (N_15297,N_9293,N_9038);
nor U15298 (N_15298,N_9028,N_11926);
and U15299 (N_15299,N_10800,N_10496);
or U15300 (N_15300,N_9066,N_8919);
nand U15301 (N_15301,N_11238,N_11478);
and U15302 (N_15302,N_9251,N_10380);
or U15303 (N_15303,N_9276,N_11766);
and U15304 (N_15304,N_8249,N_9923);
xor U15305 (N_15305,N_10565,N_11636);
nand U15306 (N_15306,N_10567,N_10547);
nand U15307 (N_15307,N_8729,N_11782);
nor U15308 (N_15308,N_11168,N_10761);
or U15309 (N_15309,N_8005,N_9340);
nand U15310 (N_15310,N_11826,N_8499);
nand U15311 (N_15311,N_9363,N_11338);
and U15312 (N_15312,N_8330,N_10476);
nand U15313 (N_15313,N_9004,N_10694);
and U15314 (N_15314,N_8817,N_8030);
or U15315 (N_15315,N_9001,N_10532);
nand U15316 (N_15316,N_11813,N_9595);
and U15317 (N_15317,N_11302,N_8822);
and U15318 (N_15318,N_8840,N_9955);
and U15319 (N_15319,N_11377,N_10440);
and U15320 (N_15320,N_9159,N_10903);
and U15321 (N_15321,N_8467,N_11286);
or U15322 (N_15322,N_11459,N_9928);
xnor U15323 (N_15323,N_9661,N_10484);
or U15324 (N_15324,N_9331,N_9784);
or U15325 (N_15325,N_10600,N_8306);
nor U15326 (N_15326,N_10310,N_11707);
xnor U15327 (N_15327,N_9885,N_9694);
nor U15328 (N_15328,N_9183,N_9527);
xnor U15329 (N_15329,N_10905,N_9128);
and U15330 (N_15330,N_8207,N_8202);
and U15331 (N_15331,N_8422,N_8848);
xnor U15332 (N_15332,N_8786,N_11925);
and U15333 (N_15333,N_10545,N_10365);
nand U15334 (N_15334,N_10722,N_10790);
and U15335 (N_15335,N_9462,N_8666);
and U15336 (N_15336,N_8939,N_8679);
or U15337 (N_15337,N_11206,N_9420);
nor U15338 (N_15338,N_10308,N_8585);
nor U15339 (N_15339,N_8165,N_8052);
or U15340 (N_15340,N_11790,N_8868);
or U15341 (N_15341,N_8824,N_8319);
or U15342 (N_15342,N_8103,N_10200);
nand U15343 (N_15343,N_9241,N_10822);
xor U15344 (N_15344,N_9610,N_8480);
nor U15345 (N_15345,N_9319,N_10264);
or U15346 (N_15346,N_8292,N_11823);
nor U15347 (N_15347,N_11317,N_11895);
nand U15348 (N_15348,N_8818,N_9903);
nor U15349 (N_15349,N_11888,N_9151);
nand U15350 (N_15350,N_9256,N_9969);
and U15351 (N_15351,N_10509,N_11808);
nand U15352 (N_15352,N_9617,N_9696);
or U15353 (N_15353,N_11422,N_11864);
xor U15354 (N_15354,N_9037,N_11980);
xnor U15355 (N_15355,N_11112,N_9139);
nor U15356 (N_15356,N_11493,N_8769);
nand U15357 (N_15357,N_10989,N_10149);
or U15358 (N_15358,N_11183,N_8150);
nor U15359 (N_15359,N_8001,N_9861);
and U15360 (N_15360,N_8930,N_10318);
and U15361 (N_15361,N_10348,N_10443);
nor U15362 (N_15362,N_9880,N_10321);
and U15363 (N_15363,N_9265,N_11945);
and U15364 (N_15364,N_8768,N_9765);
and U15365 (N_15365,N_11235,N_9714);
or U15366 (N_15366,N_10362,N_11956);
or U15367 (N_15367,N_11531,N_9736);
nor U15368 (N_15368,N_10811,N_10154);
xor U15369 (N_15369,N_9171,N_10076);
or U15370 (N_15370,N_10079,N_9549);
xnor U15371 (N_15371,N_9141,N_11967);
nand U15372 (N_15372,N_10907,N_10704);
and U15373 (N_15373,N_8075,N_10610);
nand U15374 (N_15374,N_8034,N_10595);
nor U15375 (N_15375,N_10085,N_9686);
xor U15376 (N_15376,N_9850,N_9973);
xnor U15377 (N_15377,N_11944,N_11187);
nand U15378 (N_15378,N_10740,N_8777);
and U15379 (N_15379,N_10931,N_8496);
nor U15380 (N_15380,N_9590,N_11610);
and U15381 (N_15381,N_11096,N_8726);
and U15382 (N_15382,N_11300,N_11794);
or U15383 (N_15383,N_9245,N_10529);
or U15384 (N_15384,N_11671,N_8665);
nor U15385 (N_15385,N_8204,N_10251);
or U15386 (N_15386,N_10395,N_11775);
and U15387 (N_15387,N_10296,N_11992);
nand U15388 (N_15388,N_11261,N_9047);
nor U15389 (N_15389,N_11794,N_9774);
nor U15390 (N_15390,N_10829,N_10757);
or U15391 (N_15391,N_11447,N_10767);
nor U15392 (N_15392,N_8898,N_11453);
or U15393 (N_15393,N_8108,N_10388);
and U15394 (N_15394,N_11178,N_9079);
nor U15395 (N_15395,N_10427,N_9586);
or U15396 (N_15396,N_11890,N_8996);
nand U15397 (N_15397,N_9652,N_9271);
and U15398 (N_15398,N_9253,N_10236);
nand U15399 (N_15399,N_10812,N_10425);
nand U15400 (N_15400,N_8623,N_10217);
xnor U15401 (N_15401,N_10438,N_9104);
and U15402 (N_15402,N_9915,N_11191);
nand U15403 (N_15403,N_11660,N_10945);
or U15404 (N_15404,N_9277,N_11424);
or U15405 (N_15405,N_10693,N_8917);
and U15406 (N_15406,N_11781,N_9254);
nand U15407 (N_15407,N_11611,N_9605);
or U15408 (N_15408,N_10880,N_10712);
nor U15409 (N_15409,N_11937,N_9162);
nand U15410 (N_15410,N_9456,N_8627);
xor U15411 (N_15411,N_9376,N_10277);
or U15412 (N_15412,N_10800,N_8485);
or U15413 (N_15413,N_8583,N_10970);
and U15414 (N_15414,N_11668,N_9784);
nand U15415 (N_15415,N_9203,N_8863);
nand U15416 (N_15416,N_11195,N_9639);
or U15417 (N_15417,N_8980,N_10946);
xor U15418 (N_15418,N_9669,N_9631);
and U15419 (N_15419,N_9602,N_10144);
nor U15420 (N_15420,N_10303,N_10610);
nor U15421 (N_15421,N_11365,N_8556);
or U15422 (N_15422,N_8370,N_8193);
xnor U15423 (N_15423,N_9739,N_9984);
and U15424 (N_15424,N_8151,N_9160);
nand U15425 (N_15425,N_10740,N_8387);
or U15426 (N_15426,N_11150,N_9122);
and U15427 (N_15427,N_11904,N_8641);
nor U15428 (N_15428,N_10554,N_9498);
and U15429 (N_15429,N_11676,N_11734);
and U15430 (N_15430,N_10285,N_10279);
xnor U15431 (N_15431,N_9633,N_11197);
or U15432 (N_15432,N_10683,N_8743);
nand U15433 (N_15433,N_9231,N_9854);
or U15434 (N_15434,N_8571,N_8850);
or U15435 (N_15435,N_11210,N_11568);
nand U15436 (N_15436,N_9857,N_11087);
nor U15437 (N_15437,N_11703,N_10017);
and U15438 (N_15438,N_9087,N_8326);
and U15439 (N_15439,N_10530,N_8727);
nor U15440 (N_15440,N_10015,N_11265);
and U15441 (N_15441,N_10586,N_8125);
xnor U15442 (N_15442,N_8270,N_10623);
nand U15443 (N_15443,N_11389,N_10215);
xor U15444 (N_15444,N_10445,N_11383);
or U15445 (N_15445,N_8216,N_10645);
nand U15446 (N_15446,N_10780,N_8988);
xnor U15447 (N_15447,N_11513,N_10481);
nor U15448 (N_15448,N_9482,N_8634);
nor U15449 (N_15449,N_11189,N_11843);
nor U15450 (N_15450,N_10686,N_11680);
or U15451 (N_15451,N_8405,N_11734);
nand U15452 (N_15452,N_10242,N_11459);
and U15453 (N_15453,N_11672,N_10021);
or U15454 (N_15454,N_10145,N_8931);
and U15455 (N_15455,N_8924,N_9324);
and U15456 (N_15456,N_8058,N_10785);
or U15457 (N_15457,N_9887,N_10116);
nor U15458 (N_15458,N_8077,N_9999);
nand U15459 (N_15459,N_11867,N_9202);
nor U15460 (N_15460,N_11553,N_8795);
and U15461 (N_15461,N_8802,N_10859);
and U15462 (N_15462,N_11000,N_8393);
xnor U15463 (N_15463,N_10591,N_9720);
nand U15464 (N_15464,N_10258,N_10319);
or U15465 (N_15465,N_9124,N_10172);
nor U15466 (N_15466,N_9256,N_10380);
and U15467 (N_15467,N_8074,N_11610);
xor U15468 (N_15468,N_10651,N_10108);
and U15469 (N_15469,N_8543,N_10008);
nor U15470 (N_15470,N_8972,N_10855);
xor U15471 (N_15471,N_9520,N_9487);
nor U15472 (N_15472,N_9142,N_11639);
nand U15473 (N_15473,N_11104,N_8482);
or U15474 (N_15474,N_8221,N_11105);
xor U15475 (N_15475,N_8376,N_9207);
nand U15476 (N_15476,N_9403,N_11462);
nand U15477 (N_15477,N_8621,N_10099);
nor U15478 (N_15478,N_10064,N_10593);
xnor U15479 (N_15479,N_10316,N_8501);
or U15480 (N_15480,N_10770,N_9291);
and U15481 (N_15481,N_10620,N_9634);
or U15482 (N_15482,N_11406,N_11811);
nor U15483 (N_15483,N_8374,N_9579);
nor U15484 (N_15484,N_11422,N_10829);
or U15485 (N_15485,N_8603,N_10435);
xor U15486 (N_15486,N_9204,N_8974);
or U15487 (N_15487,N_8522,N_11877);
nand U15488 (N_15488,N_9324,N_11697);
or U15489 (N_15489,N_8556,N_11720);
and U15490 (N_15490,N_8960,N_10147);
xor U15491 (N_15491,N_11795,N_9166);
nand U15492 (N_15492,N_8500,N_10054);
nand U15493 (N_15493,N_10715,N_9930);
and U15494 (N_15494,N_9029,N_11280);
or U15495 (N_15495,N_8150,N_8009);
nand U15496 (N_15496,N_11485,N_10783);
nand U15497 (N_15497,N_8376,N_10924);
xnor U15498 (N_15498,N_11590,N_11722);
nand U15499 (N_15499,N_11797,N_11470);
nor U15500 (N_15500,N_10970,N_8885);
nand U15501 (N_15501,N_8167,N_9065);
nand U15502 (N_15502,N_9463,N_10182);
nor U15503 (N_15503,N_10002,N_9219);
nor U15504 (N_15504,N_9009,N_10991);
or U15505 (N_15505,N_11424,N_8095);
nor U15506 (N_15506,N_10265,N_10461);
xor U15507 (N_15507,N_8433,N_8068);
and U15508 (N_15508,N_8703,N_9069);
xnor U15509 (N_15509,N_9542,N_8764);
xor U15510 (N_15510,N_9345,N_11599);
nand U15511 (N_15511,N_8351,N_10821);
nor U15512 (N_15512,N_11896,N_9519);
xnor U15513 (N_15513,N_9705,N_9833);
and U15514 (N_15514,N_11557,N_10542);
and U15515 (N_15515,N_9622,N_10064);
xor U15516 (N_15516,N_8773,N_9765);
and U15517 (N_15517,N_11586,N_8785);
nand U15518 (N_15518,N_11986,N_8786);
and U15519 (N_15519,N_8474,N_8189);
nand U15520 (N_15520,N_8545,N_9664);
and U15521 (N_15521,N_10495,N_9486);
and U15522 (N_15522,N_9141,N_8047);
nor U15523 (N_15523,N_11180,N_8085);
nor U15524 (N_15524,N_10938,N_10271);
xnor U15525 (N_15525,N_8666,N_8251);
xnor U15526 (N_15526,N_10845,N_9632);
xnor U15527 (N_15527,N_10394,N_9707);
nor U15528 (N_15528,N_8465,N_10881);
or U15529 (N_15529,N_10264,N_8195);
or U15530 (N_15530,N_11739,N_9811);
xor U15531 (N_15531,N_8164,N_8463);
xor U15532 (N_15532,N_11006,N_9180);
xnor U15533 (N_15533,N_11502,N_8726);
nor U15534 (N_15534,N_11072,N_11739);
and U15535 (N_15535,N_10649,N_11417);
or U15536 (N_15536,N_11545,N_9857);
xor U15537 (N_15537,N_11200,N_11309);
nor U15538 (N_15538,N_9482,N_11057);
or U15539 (N_15539,N_9010,N_8306);
xnor U15540 (N_15540,N_8300,N_8186);
nand U15541 (N_15541,N_10787,N_9786);
nor U15542 (N_15542,N_10102,N_11433);
and U15543 (N_15543,N_10874,N_11746);
nor U15544 (N_15544,N_9690,N_8627);
and U15545 (N_15545,N_10542,N_11715);
nand U15546 (N_15546,N_9821,N_9384);
nand U15547 (N_15547,N_10869,N_8965);
nand U15548 (N_15548,N_11381,N_11548);
nor U15549 (N_15549,N_8006,N_11355);
nor U15550 (N_15550,N_8907,N_8947);
nand U15551 (N_15551,N_9813,N_9149);
nor U15552 (N_15552,N_8326,N_9847);
and U15553 (N_15553,N_9497,N_10016);
or U15554 (N_15554,N_10104,N_9188);
nor U15555 (N_15555,N_11494,N_11758);
or U15556 (N_15556,N_10200,N_11638);
nand U15557 (N_15557,N_8024,N_10476);
and U15558 (N_15558,N_11711,N_10337);
nor U15559 (N_15559,N_11672,N_11241);
or U15560 (N_15560,N_9186,N_9251);
and U15561 (N_15561,N_11469,N_11833);
nand U15562 (N_15562,N_11300,N_8948);
nor U15563 (N_15563,N_10661,N_9740);
xnor U15564 (N_15564,N_8799,N_8805);
nand U15565 (N_15565,N_10294,N_11145);
nand U15566 (N_15566,N_10339,N_10309);
and U15567 (N_15567,N_8355,N_8680);
and U15568 (N_15568,N_10453,N_9863);
nand U15569 (N_15569,N_11904,N_8902);
or U15570 (N_15570,N_8876,N_11026);
and U15571 (N_15571,N_9678,N_9533);
or U15572 (N_15572,N_11760,N_11468);
nand U15573 (N_15573,N_9595,N_11083);
nand U15574 (N_15574,N_9796,N_11263);
xnor U15575 (N_15575,N_8677,N_11285);
nor U15576 (N_15576,N_9693,N_11256);
nand U15577 (N_15577,N_10682,N_11031);
xnor U15578 (N_15578,N_9888,N_10788);
xor U15579 (N_15579,N_8362,N_11320);
and U15580 (N_15580,N_9954,N_10692);
or U15581 (N_15581,N_10884,N_10549);
and U15582 (N_15582,N_11938,N_9766);
and U15583 (N_15583,N_8438,N_8023);
nand U15584 (N_15584,N_8177,N_8486);
or U15585 (N_15585,N_9211,N_9230);
xor U15586 (N_15586,N_8996,N_11589);
xnor U15587 (N_15587,N_11451,N_11915);
nor U15588 (N_15588,N_8420,N_9280);
xnor U15589 (N_15589,N_11691,N_10436);
or U15590 (N_15590,N_8516,N_10066);
nand U15591 (N_15591,N_11882,N_8062);
or U15592 (N_15592,N_8597,N_9488);
or U15593 (N_15593,N_8679,N_8511);
xor U15594 (N_15594,N_8284,N_11990);
or U15595 (N_15595,N_10982,N_10786);
xnor U15596 (N_15596,N_10725,N_11039);
nor U15597 (N_15597,N_9766,N_8647);
nor U15598 (N_15598,N_10087,N_9951);
nand U15599 (N_15599,N_8524,N_11746);
xnor U15600 (N_15600,N_10658,N_11330);
xor U15601 (N_15601,N_8734,N_8838);
and U15602 (N_15602,N_11346,N_9973);
nand U15603 (N_15603,N_9406,N_9911);
or U15604 (N_15604,N_11258,N_10730);
and U15605 (N_15605,N_10719,N_10912);
xor U15606 (N_15606,N_9471,N_8585);
xor U15607 (N_15607,N_10385,N_11614);
or U15608 (N_15608,N_8701,N_9754);
nor U15609 (N_15609,N_9723,N_11068);
and U15610 (N_15610,N_11270,N_11857);
xor U15611 (N_15611,N_8489,N_9361);
nor U15612 (N_15612,N_10961,N_9495);
and U15613 (N_15613,N_9161,N_9779);
or U15614 (N_15614,N_10221,N_10056);
nand U15615 (N_15615,N_8929,N_11382);
and U15616 (N_15616,N_8584,N_9649);
xor U15617 (N_15617,N_8472,N_10960);
nor U15618 (N_15618,N_10059,N_8444);
xor U15619 (N_15619,N_9024,N_10859);
nand U15620 (N_15620,N_9595,N_10118);
nand U15621 (N_15621,N_9900,N_10316);
or U15622 (N_15622,N_11052,N_8436);
xnor U15623 (N_15623,N_10094,N_9855);
or U15624 (N_15624,N_8343,N_11394);
or U15625 (N_15625,N_9517,N_9008);
nor U15626 (N_15626,N_8823,N_9267);
nand U15627 (N_15627,N_8867,N_10889);
or U15628 (N_15628,N_11843,N_11827);
or U15629 (N_15629,N_10287,N_9279);
nand U15630 (N_15630,N_11235,N_10281);
and U15631 (N_15631,N_11732,N_10105);
and U15632 (N_15632,N_10370,N_11774);
or U15633 (N_15633,N_8737,N_9259);
nand U15634 (N_15634,N_8141,N_10448);
nand U15635 (N_15635,N_9341,N_9130);
nor U15636 (N_15636,N_11569,N_8082);
or U15637 (N_15637,N_8647,N_9825);
nor U15638 (N_15638,N_8967,N_9689);
nor U15639 (N_15639,N_9567,N_11834);
and U15640 (N_15640,N_11160,N_10298);
nand U15641 (N_15641,N_10823,N_9815);
nor U15642 (N_15642,N_9817,N_9387);
xnor U15643 (N_15643,N_8584,N_10708);
nor U15644 (N_15644,N_9088,N_9928);
and U15645 (N_15645,N_11986,N_9710);
nand U15646 (N_15646,N_11720,N_9440);
xnor U15647 (N_15647,N_9185,N_11865);
and U15648 (N_15648,N_10665,N_9136);
or U15649 (N_15649,N_8331,N_8859);
nor U15650 (N_15650,N_8328,N_8939);
or U15651 (N_15651,N_9643,N_11035);
or U15652 (N_15652,N_9512,N_9594);
xor U15653 (N_15653,N_8846,N_11476);
nand U15654 (N_15654,N_8444,N_10511);
nand U15655 (N_15655,N_10521,N_11273);
and U15656 (N_15656,N_10005,N_8180);
nand U15657 (N_15657,N_10714,N_10377);
and U15658 (N_15658,N_8229,N_8932);
or U15659 (N_15659,N_9599,N_11368);
and U15660 (N_15660,N_9821,N_9890);
nor U15661 (N_15661,N_11248,N_8346);
nand U15662 (N_15662,N_8031,N_11182);
and U15663 (N_15663,N_11728,N_11282);
nor U15664 (N_15664,N_8114,N_11426);
or U15665 (N_15665,N_9928,N_8221);
or U15666 (N_15666,N_11922,N_9859);
and U15667 (N_15667,N_9468,N_11945);
and U15668 (N_15668,N_11257,N_8360);
and U15669 (N_15669,N_10933,N_11761);
nand U15670 (N_15670,N_9804,N_8052);
xor U15671 (N_15671,N_11622,N_10646);
or U15672 (N_15672,N_8078,N_8238);
xnor U15673 (N_15673,N_10693,N_10611);
or U15674 (N_15674,N_9464,N_9425);
nand U15675 (N_15675,N_11497,N_10688);
and U15676 (N_15676,N_8224,N_8499);
nand U15677 (N_15677,N_10478,N_11984);
nor U15678 (N_15678,N_10389,N_11541);
and U15679 (N_15679,N_11878,N_10257);
or U15680 (N_15680,N_9750,N_10326);
and U15681 (N_15681,N_9613,N_9368);
or U15682 (N_15682,N_9122,N_9743);
nor U15683 (N_15683,N_11783,N_9612);
or U15684 (N_15684,N_8747,N_9324);
nor U15685 (N_15685,N_9385,N_10785);
xor U15686 (N_15686,N_10719,N_11032);
and U15687 (N_15687,N_11840,N_10259);
or U15688 (N_15688,N_9191,N_10543);
nor U15689 (N_15689,N_11938,N_10232);
nor U15690 (N_15690,N_10909,N_10732);
and U15691 (N_15691,N_9124,N_10259);
nor U15692 (N_15692,N_10913,N_8232);
and U15693 (N_15693,N_11046,N_11619);
or U15694 (N_15694,N_8223,N_8049);
nor U15695 (N_15695,N_11082,N_8928);
nand U15696 (N_15696,N_10378,N_10928);
or U15697 (N_15697,N_11956,N_10435);
nor U15698 (N_15698,N_9747,N_11600);
nor U15699 (N_15699,N_9818,N_9895);
nor U15700 (N_15700,N_9082,N_10556);
or U15701 (N_15701,N_9945,N_11381);
nor U15702 (N_15702,N_9892,N_9858);
or U15703 (N_15703,N_8759,N_9970);
nor U15704 (N_15704,N_11076,N_11013);
nor U15705 (N_15705,N_11021,N_11817);
xor U15706 (N_15706,N_11690,N_10081);
nor U15707 (N_15707,N_9667,N_9254);
and U15708 (N_15708,N_8798,N_9934);
or U15709 (N_15709,N_9463,N_11943);
xor U15710 (N_15710,N_10232,N_11020);
xor U15711 (N_15711,N_11510,N_10535);
and U15712 (N_15712,N_11174,N_9738);
or U15713 (N_15713,N_8789,N_10261);
or U15714 (N_15714,N_10308,N_8615);
nand U15715 (N_15715,N_10654,N_11660);
and U15716 (N_15716,N_11702,N_9988);
nand U15717 (N_15717,N_11369,N_11713);
or U15718 (N_15718,N_8487,N_8096);
and U15719 (N_15719,N_10565,N_11212);
and U15720 (N_15720,N_11887,N_10715);
or U15721 (N_15721,N_10628,N_11754);
nand U15722 (N_15722,N_11159,N_11652);
nor U15723 (N_15723,N_9036,N_8852);
xor U15724 (N_15724,N_8511,N_9684);
nand U15725 (N_15725,N_8731,N_10908);
or U15726 (N_15726,N_8408,N_9903);
xor U15727 (N_15727,N_8176,N_10419);
or U15728 (N_15728,N_10765,N_9784);
and U15729 (N_15729,N_11245,N_11306);
or U15730 (N_15730,N_10869,N_8411);
xor U15731 (N_15731,N_11837,N_11054);
and U15732 (N_15732,N_10555,N_9340);
nand U15733 (N_15733,N_10852,N_8894);
or U15734 (N_15734,N_10010,N_8785);
nand U15735 (N_15735,N_9868,N_8356);
xor U15736 (N_15736,N_9689,N_11474);
xnor U15737 (N_15737,N_8366,N_11731);
or U15738 (N_15738,N_10455,N_10786);
and U15739 (N_15739,N_9367,N_9411);
or U15740 (N_15740,N_10288,N_8098);
nand U15741 (N_15741,N_9209,N_9037);
and U15742 (N_15742,N_9291,N_10930);
xnor U15743 (N_15743,N_9155,N_9356);
nor U15744 (N_15744,N_8444,N_10560);
and U15745 (N_15745,N_8358,N_9521);
xnor U15746 (N_15746,N_8542,N_8621);
xor U15747 (N_15747,N_8085,N_9082);
nand U15748 (N_15748,N_11950,N_8817);
or U15749 (N_15749,N_8105,N_11797);
nand U15750 (N_15750,N_8941,N_11094);
xor U15751 (N_15751,N_8033,N_8369);
xor U15752 (N_15752,N_8225,N_9502);
nand U15753 (N_15753,N_9784,N_10495);
nand U15754 (N_15754,N_8976,N_8404);
xor U15755 (N_15755,N_10288,N_10733);
or U15756 (N_15756,N_10739,N_10656);
nand U15757 (N_15757,N_8922,N_10827);
nand U15758 (N_15758,N_11078,N_11466);
xor U15759 (N_15759,N_9106,N_9092);
nor U15760 (N_15760,N_10836,N_9631);
or U15761 (N_15761,N_10655,N_10631);
nand U15762 (N_15762,N_9615,N_11044);
and U15763 (N_15763,N_8302,N_9740);
and U15764 (N_15764,N_11893,N_8770);
and U15765 (N_15765,N_9020,N_9109);
nor U15766 (N_15766,N_9317,N_10184);
and U15767 (N_15767,N_10704,N_9829);
and U15768 (N_15768,N_11174,N_10353);
nand U15769 (N_15769,N_11628,N_8456);
nand U15770 (N_15770,N_11013,N_11182);
xor U15771 (N_15771,N_10643,N_8197);
and U15772 (N_15772,N_9715,N_11654);
or U15773 (N_15773,N_11081,N_9274);
or U15774 (N_15774,N_9647,N_11862);
xnor U15775 (N_15775,N_11304,N_10264);
nor U15776 (N_15776,N_9990,N_10564);
and U15777 (N_15777,N_8304,N_10941);
nor U15778 (N_15778,N_9232,N_8168);
or U15779 (N_15779,N_10061,N_10696);
and U15780 (N_15780,N_10636,N_11062);
and U15781 (N_15781,N_8770,N_11848);
or U15782 (N_15782,N_11870,N_8835);
or U15783 (N_15783,N_11127,N_11256);
nand U15784 (N_15784,N_10491,N_8658);
or U15785 (N_15785,N_11484,N_8097);
xnor U15786 (N_15786,N_8154,N_8307);
nor U15787 (N_15787,N_10764,N_11828);
nor U15788 (N_15788,N_10121,N_9096);
and U15789 (N_15789,N_11484,N_11598);
and U15790 (N_15790,N_11536,N_8017);
nor U15791 (N_15791,N_9093,N_9664);
xor U15792 (N_15792,N_9958,N_11519);
nor U15793 (N_15793,N_11543,N_9254);
and U15794 (N_15794,N_11440,N_11980);
nand U15795 (N_15795,N_8237,N_9522);
xor U15796 (N_15796,N_9894,N_9276);
or U15797 (N_15797,N_11429,N_9477);
or U15798 (N_15798,N_10899,N_8576);
or U15799 (N_15799,N_11739,N_8266);
nand U15800 (N_15800,N_9232,N_11629);
and U15801 (N_15801,N_11922,N_9082);
and U15802 (N_15802,N_10619,N_9876);
or U15803 (N_15803,N_10563,N_9230);
nor U15804 (N_15804,N_10722,N_8528);
and U15805 (N_15805,N_11265,N_8614);
xor U15806 (N_15806,N_11636,N_11122);
or U15807 (N_15807,N_10458,N_9652);
xor U15808 (N_15808,N_9478,N_8212);
or U15809 (N_15809,N_9224,N_9867);
or U15810 (N_15810,N_10509,N_8129);
nor U15811 (N_15811,N_11626,N_10308);
xor U15812 (N_15812,N_9539,N_8594);
and U15813 (N_15813,N_8291,N_11430);
or U15814 (N_15814,N_10445,N_10986);
nor U15815 (N_15815,N_9949,N_11010);
nor U15816 (N_15816,N_9240,N_8131);
nor U15817 (N_15817,N_9628,N_8636);
or U15818 (N_15818,N_10102,N_8949);
nand U15819 (N_15819,N_11970,N_8411);
xor U15820 (N_15820,N_10616,N_10565);
xnor U15821 (N_15821,N_8662,N_8262);
and U15822 (N_15822,N_8335,N_10792);
xnor U15823 (N_15823,N_8226,N_8271);
xor U15824 (N_15824,N_8096,N_10505);
nor U15825 (N_15825,N_11766,N_10701);
nand U15826 (N_15826,N_8851,N_8823);
nand U15827 (N_15827,N_9242,N_10669);
and U15828 (N_15828,N_10753,N_8886);
nor U15829 (N_15829,N_9746,N_10761);
nor U15830 (N_15830,N_8647,N_11989);
nand U15831 (N_15831,N_9819,N_8958);
nand U15832 (N_15832,N_8481,N_11037);
nand U15833 (N_15833,N_9335,N_10978);
or U15834 (N_15834,N_10932,N_8615);
and U15835 (N_15835,N_8360,N_10524);
xor U15836 (N_15836,N_8862,N_9543);
nand U15837 (N_15837,N_9888,N_9276);
xor U15838 (N_15838,N_9132,N_11895);
xnor U15839 (N_15839,N_8450,N_11467);
nor U15840 (N_15840,N_10802,N_11754);
and U15841 (N_15841,N_11861,N_11137);
nand U15842 (N_15842,N_9691,N_11240);
nor U15843 (N_15843,N_8451,N_11024);
or U15844 (N_15844,N_10517,N_10619);
and U15845 (N_15845,N_9845,N_11478);
nand U15846 (N_15846,N_9630,N_10799);
xnor U15847 (N_15847,N_10962,N_11627);
or U15848 (N_15848,N_10881,N_10052);
nor U15849 (N_15849,N_10787,N_11461);
or U15850 (N_15850,N_11179,N_11428);
xor U15851 (N_15851,N_8005,N_11787);
or U15852 (N_15852,N_9248,N_10581);
nand U15853 (N_15853,N_8794,N_9778);
xnor U15854 (N_15854,N_9619,N_10298);
xor U15855 (N_15855,N_9430,N_10595);
nand U15856 (N_15856,N_8109,N_11684);
xor U15857 (N_15857,N_10934,N_9352);
xor U15858 (N_15858,N_9491,N_10894);
xor U15859 (N_15859,N_9057,N_8463);
nand U15860 (N_15860,N_11427,N_11730);
nand U15861 (N_15861,N_10478,N_10633);
xnor U15862 (N_15862,N_9940,N_8282);
nand U15863 (N_15863,N_8694,N_10765);
nand U15864 (N_15864,N_9900,N_11660);
nand U15865 (N_15865,N_9171,N_10794);
nand U15866 (N_15866,N_10433,N_9055);
nand U15867 (N_15867,N_11461,N_9159);
and U15868 (N_15868,N_11262,N_9133);
xnor U15869 (N_15869,N_8565,N_11164);
nand U15870 (N_15870,N_9562,N_8759);
xnor U15871 (N_15871,N_8284,N_9037);
nand U15872 (N_15872,N_11000,N_11622);
xnor U15873 (N_15873,N_8491,N_10165);
and U15874 (N_15874,N_8825,N_8438);
xnor U15875 (N_15875,N_11304,N_8257);
xor U15876 (N_15876,N_9512,N_9432);
nor U15877 (N_15877,N_11970,N_10071);
nor U15878 (N_15878,N_9146,N_9253);
nor U15879 (N_15879,N_9902,N_10949);
nand U15880 (N_15880,N_10341,N_8486);
or U15881 (N_15881,N_8584,N_9342);
xor U15882 (N_15882,N_11419,N_8368);
and U15883 (N_15883,N_8939,N_9814);
or U15884 (N_15884,N_10496,N_8929);
xnor U15885 (N_15885,N_9044,N_11114);
or U15886 (N_15886,N_9982,N_9359);
xor U15887 (N_15887,N_10095,N_9750);
and U15888 (N_15888,N_9131,N_9536);
xnor U15889 (N_15889,N_10836,N_8421);
nor U15890 (N_15890,N_9770,N_8252);
xor U15891 (N_15891,N_10309,N_8416);
nand U15892 (N_15892,N_11399,N_11238);
or U15893 (N_15893,N_11281,N_8102);
xor U15894 (N_15894,N_10329,N_8635);
nor U15895 (N_15895,N_11942,N_9899);
and U15896 (N_15896,N_9072,N_11901);
xnor U15897 (N_15897,N_10542,N_8450);
nor U15898 (N_15898,N_10330,N_10747);
nor U15899 (N_15899,N_9263,N_11401);
nor U15900 (N_15900,N_8394,N_9108);
nand U15901 (N_15901,N_9814,N_11879);
nand U15902 (N_15902,N_8673,N_11589);
nand U15903 (N_15903,N_8700,N_9596);
or U15904 (N_15904,N_9505,N_11598);
nor U15905 (N_15905,N_9909,N_11263);
and U15906 (N_15906,N_11886,N_9205);
nand U15907 (N_15907,N_11176,N_8040);
xnor U15908 (N_15908,N_11820,N_9829);
and U15909 (N_15909,N_8670,N_10828);
nor U15910 (N_15910,N_10457,N_9186);
xnor U15911 (N_15911,N_9978,N_9359);
nor U15912 (N_15912,N_9801,N_8588);
or U15913 (N_15913,N_8022,N_9226);
or U15914 (N_15914,N_11006,N_9095);
and U15915 (N_15915,N_9814,N_10614);
and U15916 (N_15916,N_8670,N_11718);
nor U15917 (N_15917,N_11584,N_11671);
or U15918 (N_15918,N_10866,N_10959);
or U15919 (N_15919,N_10146,N_11524);
nor U15920 (N_15920,N_11652,N_10668);
xor U15921 (N_15921,N_10370,N_8085);
xor U15922 (N_15922,N_10839,N_10482);
nand U15923 (N_15923,N_8085,N_11285);
nor U15924 (N_15924,N_9008,N_9117);
or U15925 (N_15925,N_8785,N_8092);
or U15926 (N_15926,N_11427,N_11590);
or U15927 (N_15927,N_8279,N_8742);
nor U15928 (N_15928,N_10929,N_9501);
xnor U15929 (N_15929,N_9383,N_10608);
and U15930 (N_15930,N_11372,N_10615);
and U15931 (N_15931,N_8041,N_11959);
nand U15932 (N_15932,N_9108,N_8881);
and U15933 (N_15933,N_11535,N_11132);
or U15934 (N_15934,N_8248,N_9858);
nor U15935 (N_15935,N_11739,N_9011);
xor U15936 (N_15936,N_8496,N_9115);
xnor U15937 (N_15937,N_8524,N_11441);
xnor U15938 (N_15938,N_10894,N_11292);
xnor U15939 (N_15939,N_10977,N_10390);
nand U15940 (N_15940,N_8801,N_11550);
nand U15941 (N_15941,N_8192,N_8979);
xnor U15942 (N_15942,N_9116,N_9253);
nand U15943 (N_15943,N_8356,N_8368);
xnor U15944 (N_15944,N_9951,N_8785);
nand U15945 (N_15945,N_10160,N_9246);
nor U15946 (N_15946,N_8055,N_9440);
xor U15947 (N_15947,N_8599,N_8285);
or U15948 (N_15948,N_8556,N_11348);
and U15949 (N_15949,N_11031,N_10397);
nor U15950 (N_15950,N_8892,N_9054);
and U15951 (N_15951,N_8276,N_8491);
nor U15952 (N_15952,N_9908,N_9544);
or U15953 (N_15953,N_9291,N_8605);
xnor U15954 (N_15954,N_8178,N_10032);
and U15955 (N_15955,N_9627,N_10849);
nand U15956 (N_15956,N_9997,N_11204);
nand U15957 (N_15957,N_11633,N_11374);
nor U15958 (N_15958,N_9057,N_10841);
nand U15959 (N_15959,N_11672,N_11253);
and U15960 (N_15960,N_8092,N_8600);
and U15961 (N_15961,N_8033,N_9003);
nand U15962 (N_15962,N_9956,N_8635);
nand U15963 (N_15963,N_9811,N_9131);
nor U15964 (N_15964,N_10547,N_11808);
xor U15965 (N_15965,N_10347,N_11601);
and U15966 (N_15966,N_8336,N_9741);
nor U15967 (N_15967,N_8275,N_11004);
xor U15968 (N_15968,N_11512,N_8421);
xnor U15969 (N_15969,N_11390,N_9361);
nand U15970 (N_15970,N_8203,N_8481);
nand U15971 (N_15971,N_10635,N_10860);
and U15972 (N_15972,N_9853,N_11702);
or U15973 (N_15973,N_11488,N_9323);
nor U15974 (N_15974,N_10778,N_10521);
nor U15975 (N_15975,N_9523,N_10508);
nor U15976 (N_15976,N_8401,N_11301);
and U15977 (N_15977,N_11703,N_8862);
or U15978 (N_15978,N_10021,N_11535);
nor U15979 (N_15979,N_10076,N_8626);
and U15980 (N_15980,N_8800,N_10824);
nor U15981 (N_15981,N_9674,N_8526);
xnor U15982 (N_15982,N_8748,N_11170);
and U15983 (N_15983,N_9859,N_11532);
or U15984 (N_15984,N_10854,N_10935);
and U15985 (N_15985,N_8589,N_10167);
or U15986 (N_15986,N_8377,N_11267);
nand U15987 (N_15987,N_9642,N_10970);
xor U15988 (N_15988,N_10855,N_9926);
xor U15989 (N_15989,N_9115,N_8026);
and U15990 (N_15990,N_11716,N_10796);
or U15991 (N_15991,N_9518,N_9187);
nand U15992 (N_15992,N_9028,N_8658);
xor U15993 (N_15993,N_9592,N_10347);
or U15994 (N_15994,N_10458,N_10692);
xnor U15995 (N_15995,N_8940,N_11316);
and U15996 (N_15996,N_11296,N_11494);
nor U15997 (N_15997,N_10049,N_8367);
nor U15998 (N_15998,N_9804,N_11192);
nand U15999 (N_15999,N_9688,N_10922);
xnor U16000 (N_16000,N_12066,N_14331);
nor U16001 (N_16001,N_15986,N_12860);
nor U16002 (N_16002,N_14369,N_15070);
nand U16003 (N_16003,N_12109,N_13807);
and U16004 (N_16004,N_12030,N_12168);
xor U16005 (N_16005,N_13906,N_15798);
nor U16006 (N_16006,N_13384,N_13857);
xor U16007 (N_16007,N_14405,N_12247);
xor U16008 (N_16008,N_12347,N_12282);
and U16009 (N_16009,N_14920,N_15424);
xor U16010 (N_16010,N_15859,N_12164);
nor U16011 (N_16011,N_14915,N_12616);
or U16012 (N_16012,N_14825,N_15998);
and U16013 (N_16013,N_15925,N_14417);
and U16014 (N_16014,N_13977,N_13856);
nand U16015 (N_16015,N_13218,N_14322);
xor U16016 (N_16016,N_13047,N_14004);
nor U16017 (N_16017,N_14802,N_14321);
nor U16018 (N_16018,N_15526,N_14737);
nor U16019 (N_16019,N_12734,N_15778);
and U16020 (N_16020,N_15226,N_14413);
xor U16021 (N_16021,N_13204,N_15606);
nand U16022 (N_16022,N_13706,N_15076);
and U16023 (N_16023,N_13037,N_15217);
or U16024 (N_16024,N_12565,N_15899);
or U16025 (N_16025,N_15811,N_12926);
and U16026 (N_16026,N_12851,N_13871);
nor U16027 (N_16027,N_15551,N_15101);
or U16028 (N_16028,N_14037,N_15609);
nor U16029 (N_16029,N_15637,N_13736);
and U16030 (N_16030,N_14766,N_13006);
and U16031 (N_16031,N_14008,N_13644);
xnor U16032 (N_16032,N_13525,N_15722);
or U16033 (N_16033,N_14309,N_12686);
xnor U16034 (N_16034,N_15398,N_12158);
xor U16035 (N_16035,N_12106,N_12888);
nand U16036 (N_16036,N_14010,N_13827);
nand U16037 (N_16037,N_15168,N_13855);
nand U16038 (N_16038,N_12610,N_15997);
or U16039 (N_16039,N_15454,N_15981);
and U16040 (N_16040,N_12972,N_12014);
nand U16041 (N_16041,N_15565,N_14348);
or U16042 (N_16042,N_12508,N_15384);
nand U16043 (N_16043,N_15336,N_13143);
or U16044 (N_16044,N_15535,N_15490);
or U16045 (N_16045,N_14900,N_12986);
and U16046 (N_16046,N_13165,N_12693);
xor U16047 (N_16047,N_13010,N_14217);
nand U16048 (N_16048,N_13067,N_14127);
xnor U16049 (N_16049,N_12436,N_13998);
xnor U16050 (N_16050,N_15635,N_12017);
nand U16051 (N_16051,N_12403,N_12024);
or U16052 (N_16052,N_15307,N_12391);
nand U16053 (N_16053,N_15060,N_13149);
and U16054 (N_16054,N_13030,N_12800);
and U16055 (N_16055,N_15321,N_12053);
nor U16056 (N_16056,N_13792,N_12067);
nand U16057 (N_16057,N_12887,N_14157);
xor U16058 (N_16058,N_14657,N_14717);
nor U16059 (N_16059,N_15913,N_12601);
nand U16060 (N_16060,N_14082,N_13338);
nand U16061 (N_16061,N_15770,N_12228);
nand U16062 (N_16062,N_15466,N_15977);
and U16063 (N_16063,N_12358,N_13873);
nand U16064 (N_16064,N_12397,N_15359);
nand U16065 (N_16065,N_13043,N_13563);
xor U16066 (N_16066,N_15086,N_15935);
nor U16067 (N_16067,N_12945,N_13130);
nand U16068 (N_16068,N_14169,N_14958);
xnor U16069 (N_16069,N_12160,N_12351);
or U16070 (N_16070,N_13958,N_12617);
or U16071 (N_16071,N_13119,N_12513);
nand U16072 (N_16072,N_14660,N_13232);
and U16073 (N_16073,N_12793,N_14675);
or U16074 (N_16074,N_12473,N_13961);
nor U16075 (N_16075,N_12520,N_13612);
or U16076 (N_16076,N_15430,N_13800);
nor U16077 (N_16077,N_12544,N_13409);
xnor U16078 (N_16078,N_12789,N_13317);
and U16079 (N_16079,N_12037,N_12438);
and U16080 (N_16080,N_13478,N_13724);
nor U16081 (N_16081,N_12779,N_13840);
xor U16082 (N_16082,N_13224,N_13781);
and U16083 (N_16083,N_13948,N_14954);
xnor U16084 (N_16084,N_12833,N_13131);
nor U16085 (N_16085,N_14424,N_12556);
xnor U16086 (N_16086,N_13164,N_15559);
or U16087 (N_16087,N_12129,N_14077);
or U16088 (N_16088,N_15143,N_15381);
xor U16089 (N_16089,N_13760,N_12339);
xor U16090 (N_16090,N_13234,N_12704);
nand U16091 (N_16091,N_14682,N_13445);
or U16092 (N_16092,N_13475,N_15516);
nand U16093 (N_16093,N_13682,N_12019);
or U16094 (N_16094,N_15041,N_13400);
nor U16095 (N_16095,N_15073,N_12469);
and U16096 (N_16096,N_15427,N_15180);
xnor U16097 (N_16097,N_14941,N_15806);
and U16098 (N_16098,N_13930,N_13254);
and U16099 (N_16099,N_13088,N_14994);
and U16100 (N_16100,N_12794,N_15155);
nor U16101 (N_16101,N_15318,N_15577);
and U16102 (N_16102,N_12707,N_15158);
nor U16103 (N_16103,N_13056,N_12294);
nor U16104 (N_16104,N_12760,N_14389);
and U16105 (N_16105,N_12232,N_15580);
nand U16106 (N_16106,N_15269,N_15819);
nor U16107 (N_16107,N_12356,N_12212);
nor U16108 (N_16108,N_15405,N_14517);
or U16109 (N_16109,N_15149,N_14306);
nor U16110 (N_16110,N_14045,N_12973);
nor U16111 (N_16111,N_12879,N_14176);
and U16112 (N_16112,N_15259,N_14299);
and U16113 (N_16113,N_12426,N_12906);
and U16114 (N_16114,N_14252,N_15864);
nand U16115 (N_16115,N_14735,N_14133);
and U16116 (N_16116,N_13122,N_12865);
and U16117 (N_16117,N_15994,N_12861);
xor U16118 (N_16118,N_12036,N_14788);
xor U16119 (N_16119,N_13878,N_15782);
nor U16120 (N_16120,N_15726,N_12183);
or U16121 (N_16121,N_13801,N_13548);
xor U16122 (N_16122,N_12303,N_14151);
nand U16123 (N_16123,N_12984,N_13513);
and U16124 (N_16124,N_14233,N_15173);
nor U16125 (N_16125,N_13009,N_13341);
xor U16126 (N_16126,N_15162,N_12603);
nand U16127 (N_16127,N_13701,N_12392);
nand U16128 (N_16128,N_15825,N_12802);
and U16129 (N_16129,N_14962,N_14659);
nor U16130 (N_16130,N_14633,N_13619);
or U16131 (N_16131,N_13744,N_12839);
xor U16132 (N_16132,N_13918,N_12065);
nor U16133 (N_16133,N_13888,N_14241);
nand U16134 (N_16134,N_13872,N_12235);
nor U16135 (N_16135,N_13019,N_14960);
and U16136 (N_16136,N_12411,N_15129);
and U16137 (N_16137,N_14130,N_14070);
nor U16138 (N_16138,N_13710,N_14815);
nand U16139 (N_16139,N_15447,N_15995);
and U16140 (N_16140,N_13649,N_15821);
nand U16141 (N_16141,N_13516,N_13770);
nor U16142 (N_16142,N_12107,N_14810);
and U16143 (N_16143,N_15274,N_14845);
and U16144 (N_16144,N_14315,N_14724);
nor U16145 (N_16145,N_13875,N_15252);
xor U16146 (N_16146,N_15013,N_15902);
xor U16147 (N_16147,N_14428,N_13725);
xor U16148 (N_16148,N_12846,N_14198);
nand U16149 (N_16149,N_12821,N_13117);
nand U16150 (N_16150,N_12165,N_14163);
and U16151 (N_16151,N_12652,N_12157);
xor U16152 (N_16152,N_13665,N_13246);
or U16153 (N_16153,N_14086,N_14154);
xor U16154 (N_16154,N_13837,N_15246);
nand U16155 (N_16155,N_15063,N_15970);
nor U16156 (N_16156,N_13315,N_13798);
xor U16157 (N_16157,N_15633,N_14449);
xnor U16158 (N_16158,N_13713,N_15377);
nand U16159 (N_16159,N_12390,N_15685);
or U16160 (N_16160,N_13116,N_12174);
and U16161 (N_16161,N_14692,N_15542);
nor U16162 (N_16162,N_14100,N_12614);
nor U16163 (N_16163,N_15955,N_14518);
xor U16164 (N_16164,N_14083,N_12340);
nand U16165 (N_16165,N_14279,N_12316);
and U16166 (N_16166,N_12700,N_14113);
or U16167 (N_16167,N_13309,N_13370);
xor U16168 (N_16168,N_13076,N_13499);
xnor U16169 (N_16169,N_15059,N_13180);
or U16170 (N_16170,N_13344,N_13676);
nor U16171 (N_16171,N_14333,N_13062);
and U16172 (N_16172,N_15718,N_13205);
and U16173 (N_16173,N_14214,N_15746);
nand U16174 (N_16174,N_12337,N_12239);
nor U16175 (N_16175,N_14658,N_14245);
nand U16176 (N_16176,N_15593,N_12499);
nor U16177 (N_16177,N_15844,N_13284);
nand U16178 (N_16178,N_13380,N_14789);
and U16179 (N_16179,N_15378,N_14770);
or U16180 (N_16180,N_15368,N_13568);
and U16181 (N_16181,N_13610,N_12699);
nand U16182 (N_16182,N_12357,N_14543);
xor U16183 (N_16183,N_15800,N_15115);
nor U16184 (N_16184,N_14505,N_15411);
xor U16185 (N_16185,N_14227,N_14533);
nand U16186 (N_16186,N_13882,N_14809);
nor U16187 (N_16187,N_14503,N_12737);
nor U16188 (N_16188,N_14952,N_12990);
nor U16189 (N_16189,N_12214,N_14351);
nor U16190 (N_16190,N_14025,N_13763);
or U16191 (N_16191,N_12702,N_13401);
and U16192 (N_16192,N_15191,N_12830);
or U16193 (N_16193,N_13783,N_13280);
nor U16194 (N_16194,N_12754,N_14251);
nor U16195 (N_16195,N_14913,N_13040);
nand U16196 (N_16196,N_14561,N_15497);
xnor U16197 (N_16197,N_13864,N_15001);
xnor U16198 (N_16198,N_12903,N_12582);
and U16199 (N_16199,N_14160,N_14730);
or U16200 (N_16200,N_14071,N_15097);
nand U16201 (N_16201,N_15938,N_13477);
nor U16202 (N_16202,N_14653,N_13161);
xor U16203 (N_16203,N_12971,N_14884);
or U16204 (N_16204,N_13427,N_12177);
nor U16205 (N_16205,N_14338,N_13843);
xnor U16206 (N_16206,N_14515,N_15761);
xor U16207 (N_16207,N_15521,N_13994);
nor U16208 (N_16208,N_14409,N_13025);
and U16209 (N_16209,N_15412,N_13520);
xnor U16210 (N_16210,N_13667,N_14755);
and U16211 (N_16211,N_15894,N_13543);
xor U16212 (N_16212,N_13313,N_13751);
nor U16213 (N_16213,N_12344,N_15507);
nor U16214 (N_16214,N_12795,N_12723);
or U16215 (N_16215,N_13891,N_15583);
and U16216 (N_16216,N_12824,N_15476);
or U16217 (N_16217,N_15029,N_13290);
xnor U16218 (N_16218,N_14972,N_15895);
nand U16219 (N_16219,N_15716,N_13029);
or U16220 (N_16220,N_15792,N_13426);
nor U16221 (N_16221,N_15199,N_15174);
nand U16222 (N_16222,N_15966,N_12034);
nand U16223 (N_16223,N_14065,N_14850);
xor U16224 (N_16224,N_14525,N_15514);
xor U16225 (N_16225,N_14075,N_14950);
or U16226 (N_16226,N_12204,N_13109);
nor U16227 (N_16227,N_14656,N_15181);
nand U16228 (N_16228,N_13432,N_13822);
nor U16229 (N_16229,N_13894,N_14641);
nor U16230 (N_16230,N_12048,N_14150);
xor U16231 (N_16231,N_13080,N_12078);
or U16232 (N_16232,N_12904,N_13892);
xnor U16233 (N_16233,N_14666,N_13386);
nand U16234 (N_16234,N_12983,N_12180);
or U16235 (N_16235,N_14786,N_12277);
or U16236 (N_16236,N_12470,N_13461);
nor U16237 (N_16237,N_13422,N_14228);
nor U16238 (N_16238,N_14537,N_15508);
and U16239 (N_16239,N_12678,N_13887);
nand U16240 (N_16240,N_14566,N_15779);
and U16241 (N_16241,N_12364,N_13579);
xor U16242 (N_16242,N_15627,N_15592);
and U16243 (N_16243,N_13262,N_14420);
or U16244 (N_16244,N_15908,N_15728);
xnor U16245 (N_16245,N_13046,N_12332);
nand U16246 (N_16246,N_12877,N_15028);
and U16247 (N_16247,N_14317,N_13836);
nand U16248 (N_16248,N_14775,N_15492);
nand U16249 (N_16249,N_12598,N_15758);
and U16250 (N_16250,N_14883,N_14598);
nor U16251 (N_16251,N_14545,N_12694);
nor U16252 (N_16252,N_15022,N_15103);
nor U16253 (N_16253,N_15896,N_12421);
nand U16254 (N_16254,N_15564,N_12121);
nor U16255 (N_16255,N_12629,N_12864);
or U16256 (N_16256,N_12871,N_13115);
nand U16257 (N_16257,N_14337,N_14250);
or U16258 (N_16258,N_14795,N_13472);
nand U16259 (N_16259,N_13811,N_14425);
nand U16260 (N_16260,N_15735,N_15413);
xnor U16261 (N_16261,N_14934,N_12122);
and U16262 (N_16262,N_15144,N_13362);
xor U16263 (N_16263,N_12855,N_12590);
xnor U16264 (N_16264,N_14190,N_12060);
xor U16265 (N_16265,N_14710,N_13852);
nor U16266 (N_16266,N_12703,N_15153);
nor U16267 (N_16267,N_12536,N_12105);
or U16268 (N_16268,N_15085,N_14205);
xor U16269 (N_16269,N_14437,N_13349);
and U16270 (N_16270,N_15419,N_15275);
nand U16271 (N_16271,N_14536,N_15932);
nand U16272 (N_16272,N_14534,N_12008);
nand U16273 (N_16273,N_14196,N_12335);
and U16274 (N_16274,N_13403,N_12216);
or U16275 (N_16275,N_12203,N_15812);
and U16276 (N_16276,N_14864,N_14164);
nand U16277 (N_16277,N_12382,N_12462);
or U16278 (N_16278,N_13421,N_13850);
and U16279 (N_16279,N_12938,N_13297);
and U16280 (N_16280,N_12127,N_12234);
nand U16281 (N_16281,N_15946,N_12994);
xnor U16282 (N_16282,N_14370,N_13990);
and U16283 (N_16283,N_12831,N_14118);
nor U16284 (N_16284,N_13417,N_13718);
xor U16285 (N_16285,N_12052,N_13708);
nand U16286 (N_16286,N_12044,N_13042);
xor U16287 (N_16287,N_13127,N_15442);
nand U16288 (N_16288,N_12817,N_13176);
or U16289 (N_16289,N_12405,N_15750);
nand U16290 (N_16290,N_15841,N_13668);
nand U16291 (N_16291,N_13263,N_14297);
xnor U16292 (N_16292,N_12095,N_13787);
or U16293 (N_16293,N_15433,N_13883);
and U16294 (N_16294,N_14155,N_15455);
nand U16295 (N_16295,N_15629,N_12498);
nand U16296 (N_16296,N_14387,N_15373);
or U16297 (N_16297,N_14436,N_12862);
or U16298 (N_16298,N_12563,N_12491);
and U16299 (N_16299,N_15300,N_12759);
nand U16300 (N_16300,N_12051,N_14401);
or U16301 (N_16301,N_15224,N_12135);
and U16302 (N_16302,N_12479,N_14927);
xor U16303 (N_16303,N_14649,N_15051);
nor U16304 (N_16304,N_13346,N_15035);
nor U16305 (N_16305,N_12352,N_13705);
nor U16306 (N_16306,N_12452,N_13425);
and U16307 (N_16307,N_13778,N_12837);
xor U16308 (N_16308,N_14516,N_13919);
nor U16309 (N_16309,N_14341,N_13993);
or U16310 (N_16310,N_14930,N_15372);
nor U16311 (N_16311,N_13173,N_15872);
xnor U16312 (N_16312,N_14925,N_14942);
and U16313 (N_16313,N_15450,N_15467);
or U16314 (N_16314,N_13527,N_14197);
or U16315 (N_16315,N_15288,N_15401);
nor U16316 (N_16316,N_13617,N_14628);
xnor U16317 (N_16317,N_12149,N_15148);
nand U16318 (N_16318,N_14290,N_12534);
nor U16319 (N_16319,N_13199,N_14679);
nor U16320 (N_16320,N_12557,N_15416);
or U16321 (N_16321,N_14115,N_15944);
or U16322 (N_16322,N_14288,N_13483);
xor U16323 (N_16323,N_14350,N_15404);
and U16324 (N_16324,N_14731,N_13106);
nor U16325 (N_16325,N_15658,N_14318);
xor U16326 (N_16326,N_14922,N_13820);
nand U16327 (N_16327,N_13632,N_12928);
and U16328 (N_16328,N_14207,N_12959);
xor U16329 (N_16329,N_12957,N_15712);
or U16330 (N_16330,N_13625,N_15566);
nor U16331 (N_16331,N_15376,N_14423);
or U16332 (N_16332,N_12688,N_12538);
or U16333 (N_16333,N_12844,N_14109);
and U16334 (N_16334,N_12002,N_12675);
xnor U16335 (N_16335,N_14044,N_14550);
nor U16336 (N_16336,N_15860,N_13305);
nand U16337 (N_16337,N_13847,N_13711);
xor U16338 (N_16338,N_12627,N_15027);
and U16339 (N_16339,N_14806,N_14800);
or U16340 (N_16340,N_13321,N_15396);
and U16341 (N_16341,N_12960,N_15688);
xnor U16342 (N_16342,N_13323,N_13589);
and U16343 (N_16343,N_12432,N_14271);
or U16344 (N_16344,N_15822,N_13438);
or U16345 (N_16345,N_12345,N_14732);
xnor U16346 (N_16346,N_14796,N_15287);
or U16347 (N_16347,N_14528,N_14531);
nand U16348 (N_16348,N_12854,N_14498);
xor U16349 (N_16349,N_12799,N_14946);
xnor U16350 (N_16350,N_13907,N_14439);
and U16351 (N_16351,N_15117,N_15748);
nand U16352 (N_16352,N_15574,N_15383);
xnor U16353 (N_16353,N_13938,N_12920);
xnor U16354 (N_16354,N_15885,N_15988);
nand U16355 (N_16355,N_15581,N_15655);
nand U16356 (N_16356,N_12043,N_14846);
nor U16357 (N_16357,N_14791,N_14638);
and U16358 (N_16358,N_13904,N_15717);
and U16359 (N_16359,N_13788,N_12246);
nor U16360 (N_16360,N_12417,N_13739);
or U16361 (N_16361,N_13740,N_15588);
nand U16362 (N_16362,N_12620,N_14608);
or U16363 (N_16363,N_14548,N_14509);
or U16364 (N_16364,N_13183,N_12684);
nand U16365 (N_16365,N_13576,N_13108);
nand U16366 (N_16366,N_13437,N_13156);
nor U16367 (N_16367,N_14339,N_15694);
or U16368 (N_16368,N_14132,N_12481);
nand U16369 (N_16369,N_14159,N_14346);
or U16370 (N_16370,N_13345,N_15867);
nor U16371 (N_16371,N_12057,N_14602);
nor U16372 (N_16372,N_12101,N_12161);
nor U16373 (N_16373,N_13562,N_12213);
and U16374 (N_16374,N_13749,N_12826);
nor U16375 (N_16375,N_13113,N_14092);
and U16376 (N_16376,N_14480,N_15838);
or U16377 (N_16377,N_14836,N_12097);
and U16378 (N_16378,N_14126,N_13310);
or U16379 (N_16379,N_12896,N_13210);
and U16380 (N_16380,N_14215,N_14576);
nor U16381 (N_16381,N_14764,N_15011);
or U16382 (N_16382,N_12064,N_15068);
nand U16383 (N_16383,N_15094,N_12338);
xor U16384 (N_16384,N_13782,N_12979);
nor U16385 (N_16385,N_15686,N_12633);
or U16386 (N_16386,N_13174,N_13936);
xnor U16387 (N_16387,N_14816,N_13842);
xor U16388 (N_16388,N_14275,N_14995);
nand U16389 (N_16389,N_15711,N_15484);
nor U16390 (N_16390,N_13796,N_13353);
xnor U16391 (N_16391,N_12768,N_13126);
xnor U16392 (N_16392,N_15904,N_14054);
nand U16393 (N_16393,N_13142,N_14374);
or U16394 (N_16394,N_12948,N_12395);
xnor U16395 (N_16395,N_13986,N_12114);
nor U16396 (N_16396,N_15532,N_14671);
nor U16397 (N_16397,N_15941,N_14378);
xor U16398 (N_16398,N_13399,N_12041);
nor U16399 (N_16399,N_12517,N_13652);
or U16400 (N_16400,N_12910,N_13066);
and U16401 (N_16401,N_12708,N_12753);
nand U16402 (N_16402,N_13479,N_14277);
or U16403 (N_16403,N_14352,N_13187);
or U16404 (N_16404,N_15693,N_14293);
xor U16405 (N_16405,N_13954,N_14371);
and U16406 (N_16406,N_12267,N_14097);
nand U16407 (N_16407,N_14161,N_14728);
or U16408 (N_16408,N_15671,N_15370);
nor U16409 (N_16409,N_14382,N_14918);
and U16410 (N_16410,N_15910,N_15256);
nor U16411 (N_16411,N_13012,N_15053);
or U16412 (N_16412,N_15724,N_14752);
and U16413 (N_16413,N_13190,N_12825);
xnor U16414 (N_16414,N_14460,N_15539);
xnor U16415 (N_16415,N_14327,N_15408);
nor U16416 (N_16416,N_12515,N_15803);
nor U16417 (N_16417,N_12714,N_15952);
xor U16418 (N_16418,N_12297,N_12327);
nor U16419 (N_16419,N_14396,N_12223);
and U16420 (N_16420,N_15323,N_13249);
nor U16421 (N_16421,N_14998,N_13523);
xnor U16422 (N_16422,N_12574,N_14146);
xnor U16423 (N_16423,N_12859,N_13584);
and U16424 (N_16424,N_14639,N_12219);
or U16425 (N_16425,N_15348,N_14385);
nor U16426 (N_16426,N_12163,N_13570);
nor U16427 (N_16427,N_14074,N_13044);
or U16428 (N_16428,N_14103,N_13935);
or U16429 (N_16429,N_12309,N_15641);
and U16430 (N_16430,N_12413,N_15087);
xnor U16431 (N_16431,N_12288,N_15834);
and U16432 (N_16432,N_15017,N_13077);
or U16433 (N_16433,N_15345,N_13188);
xor U16434 (N_16434,N_12231,N_12250);
nor U16435 (N_16435,N_14880,N_12883);
or U16436 (N_16436,N_15884,N_14397);
xor U16437 (N_16437,N_14373,N_15030);
or U16438 (N_16438,N_15346,N_13406);
nor U16439 (N_16439,N_13420,N_12806);
xnor U16440 (N_16440,N_15617,N_15190);
or U16441 (N_16441,N_12343,N_12878);
and U16442 (N_16442,N_12090,N_13726);
nor U16443 (N_16443,N_13152,N_15487);
xnor U16444 (N_16444,N_12644,N_13829);
or U16445 (N_16445,N_15605,N_15084);
xor U16446 (N_16446,N_14458,N_13003);
nor U16447 (N_16447,N_13022,N_12415);
nand U16448 (N_16448,N_13326,N_15483);
or U16449 (N_16449,N_15393,N_13671);
xnor U16450 (N_16450,N_14364,N_14664);
xor U16451 (N_16451,N_12068,N_14254);
nor U16452 (N_16452,N_13503,N_15285);
nor U16453 (N_16453,N_13566,N_13357);
nor U16454 (N_16454,N_15648,N_15969);
xor U16455 (N_16455,N_14344,N_13910);
or U16456 (N_16456,N_12656,N_14342);
and U16457 (N_16457,N_14591,N_12669);
and U16458 (N_16458,N_14136,N_13695);
nand U16459 (N_16459,N_12419,N_15296);
nor U16460 (N_16460,N_14665,N_12460);
or U16461 (N_16461,N_12384,N_12492);
xnor U16462 (N_16462,N_13685,N_14780);
or U16463 (N_16463,N_13236,N_13070);
xnor U16464 (N_16464,N_15261,N_13079);
nor U16465 (N_16465,N_14587,N_14099);
xor U16466 (N_16466,N_14655,N_15554);
nand U16467 (N_16467,N_14211,N_15156);
and U16468 (N_16468,N_15620,N_14137);
nor U16469 (N_16469,N_15328,N_15293);
and U16470 (N_16470,N_15951,N_12319);
nor U16471 (N_16471,N_13244,N_13239);
or U16472 (N_16472,N_13825,N_13269);
nand U16473 (N_16473,N_14944,N_15082);
xor U16474 (N_16474,N_12162,N_12027);
and U16475 (N_16475,N_13163,N_13243);
xor U16476 (N_16476,N_14812,N_13608);
or U16477 (N_16477,N_12398,N_14708);
nor U16478 (N_16478,N_13858,N_12747);
xor U16479 (N_16479,N_12437,N_12665);
nor U16480 (N_16480,N_14347,N_13352);
or U16481 (N_16481,N_13583,N_14723);
and U16482 (N_16482,N_15108,N_14859);
and U16483 (N_16483,N_13699,N_12061);
or U16484 (N_16484,N_13927,N_13064);
or U16485 (N_16485,N_12716,N_12431);
or U16486 (N_16486,N_13517,N_14018);
xor U16487 (N_16487,N_12981,N_12238);
or U16488 (N_16488,N_15081,N_15015);
and U16489 (N_16489,N_15876,N_14016);
xor U16490 (N_16490,N_15584,N_15773);
nand U16491 (N_16491,N_15267,N_14226);
or U16492 (N_16492,N_13946,N_14175);
xnor U16493 (N_16493,N_15525,N_15680);
nand U16494 (N_16494,N_12892,N_14570);
and U16495 (N_16495,N_12275,N_15311);
or U16496 (N_16496,N_14209,N_12512);
nand U16497 (N_16497,N_15996,N_15471);
or U16498 (N_16498,N_13550,N_14138);
xor U16499 (N_16499,N_14158,N_13953);
and U16500 (N_16500,N_12776,N_12805);
nor U16501 (N_16501,N_15116,N_15481);
nand U16502 (N_16502,N_13752,N_12112);
nand U16503 (N_16503,N_14208,N_14560);
xor U16504 (N_16504,N_13206,N_12369);
and U16505 (N_16505,N_14466,N_13446);
xnor U16506 (N_16506,N_14117,N_15298);
nor U16507 (N_16507,N_15244,N_13075);
or U16508 (N_16508,N_15582,N_14484);
nor U16509 (N_16509,N_14242,N_14779);
and U16510 (N_16510,N_14911,N_13600);
nor U16511 (N_16511,N_12638,N_15830);
nor U16512 (N_16512,N_13081,N_14544);
nand U16513 (N_16513,N_13496,N_13507);
nor U16514 (N_16514,N_13675,N_14538);
and U16515 (N_16515,N_12485,N_13248);
and U16516 (N_16516,N_13331,N_15184);
nor U16517 (N_16517,N_12350,N_12880);
xor U16518 (N_16518,N_15172,N_12023);
and U16519 (N_16519,N_15861,N_15796);
nor U16520 (N_16520,N_14381,N_12439);
and U16521 (N_16521,N_13912,N_14868);
and U16522 (N_16522,N_13967,N_15982);
nand U16523 (N_16523,N_15506,N_14052);
nor U16524 (N_16524,N_14617,N_15745);
or U16525 (N_16525,N_14741,N_14360);
nor U16526 (N_16526,N_13678,N_13350);
and U16527 (N_16527,N_13340,N_14002);
xor U16528 (N_16528,N_12608,N_13880);
xnor U16529 (N_16529,N_14578,N_14557);
and U16530 (N_16530,N_12552,N_14267);
xor U16531 (N_16531,N_13831,N_15573);
nor U16532 (N_16532,N_14192,N_14345);
or U16533 (N_16533,N_15211,N_14087);
nand U16534 (N_16534,N_14062,N_12522);
or U16535 (N_16535,N_12039,N_15410);
and U16536 (N_16536,N_13158,N_14896);
and U16537 (N_16537,N_13048,N_13114);
nor U16538 (N_16538,N_13237,N_14687);
xor U16539 (N_16539,N_12689,N_12989);
or U16540 (N_16540,N_12474,N_14854);
or U16541 (N_16541,N_14798,N_12809);
nand U16542 (N_16542,N_13182,N_13952);
nand U16543 (N_16543,N_12933,N_15183);
xnor U16544 (N_16544,N_13041,N_13714);
and U16545 (N_16545,N_14905,N_13133);
xor U16546 (N_16546,N_12650,N_14527);
or U16547 (N_16547,N_13092,N_13287);
xnor U16548 (N_16548,N_15239,N_14580);
nor U16549 (N_16549,N_15472,N_13963);
nand U16550 (N_16550,N_14066,N_15768);
nor U16551 (N_16551,N_13201,N_13459);
nor U16552 (N_16552,N_13832,N_15600);
nand U16553 (N_16553,N_15194,N_13700);
or U16554 (N_16554,N_12328,N_14221);
xor U16555 (N_16555,N_14829,N_12530);
nand U16556 (N_16556,N_12077,N_15003);
or U16557 (N_16557,N_13674,N_12968);
xor U16558 (N_16558,N_13603,N_13036);
nand U16559 (N_16559,N_15851,N_12494);
nand U16560 (N_16560,N_12919,N_12209);
nor U16561 (N_16561,N_14268,N_14224);
nor U16562 (N_16562,N_15349,N_13428);
nand U16563 (N_16563,N_12434,N_14316);
nor U16564 (N_16564,N_14935,N_12978);
nand U16565 (N_16565,N_15047,N_14199);
or U16566 (N_16566,N_15327,N_15391);
nor U16567 (N_16567,N_12224,N_15984);
xor U16568 (N_16568,N_15795,N_15868);
xor U16569 (N_16569,N_12843,N_12393);
nand U16570 (N_16570,N_12424,N_13096);
xor U16571 (N_16571,N_14431,N_14419);
and U16572 (N_16572,N_13696,N_13488);
xor U16573 (N_16573,N_12602,N_15824);
or U16574 (N_16574,N_12088,N_14650);
nand U16575 (N_16575,N_12728,N_12982);
and U16576 (N_16576,N_14050,N_13677);
nand U16577 (N_16577,N_15354,N_14957);
nor U16578 (N_16578,N_14760,N_12283);
xor U16579 (N_16579,N_15380,N_13686);
and U16580 (N_16580,N_13213,N_14114);
and U16581 (N_16581,N_12526,N_12930);
nor U16582 (N_16582,N_14468,N_14477);
nand U16583 (N_16583,N_14607,N_12256);
or U16584 (N_16584,N_12546,N_14408);
xnor U16585 (N_16585,N_15220,N_14494);
nand U16586 (N_16586,N_14343,N_13304);
xnor U16587 (N_16587,N_12706,N_13813);
and U16588 (N_16588,N_13526,N_15808);
nor U16589 (N_16589,N_14430,N_14844);
xnor U16590 (N_16590,N_12087,N_13853);
nand U16591 (N_16591,N_12894,N_14429);
nand U16592 (N_16592,N_14624,N_14003);
xnor U16593 (N_16593,N_12588,N_12171);
or U16594 (N_16594,N_12814,N_12543);
or U16595 (N_16595,N_12942,N_12649);
or U16596 (N_16596,N_15495,N_12189);
nor U16597 (N_16597,N_15294,N_13288);
xnor U16598 (N_16598,N_12265,N_13229);
and U16599 (N_16599,N_15690,N_15324);
and U16600 (N_16600,N_13616,N_13884);
nor U16601 (N_16601,N_14028,N_13535);
and U16602 (N_16602,N_14698,N_14212);
xor U16603 (N_16603,N_15901,N_15703);
or U16604 (N_16604,N_15734,N_12455);
or U16605 (N_16605,N_14610,N_12550);
xnor U16606 (N_16606,N_13226,N_13580);
nand U16607 (N_16607,N_15077,N_15891);
xor U16608 (N_16608,N_14451,N_12254);
nand U16609 (N_16609,N_13463,N_13172);
nand U16610 (N_16610,N_13251,N_15446);
xnor U16611 (N_16611,N_15095,N_12570);
or U16612 (N_16612,N_12985,N_13945);
xor U16613 (N_16613,N_12807,N_15738);
xor U16614 (N_16614,N_14124,N_13055);
or U16615 (N_16615,N_14597,N_14740);
and U16616 (N_16616,N_13318,N_15105);
nor U16617 (N_16617,N_14276,N_14223);
nor U16618 (N_16618,N_12225,N_15740);
and U16619 (N_16619,N_15132,N_15216);
xnor U16620 (N_16620,N_14349,N_15119);
and U16621 (N_16621,N_12924,N_13135);
nand U16622 (N_16622,N_12482,N_13679);
or U16623 (N_16623,N_12872,N_13402);
or U16624 (N_16624,N_12028,N_13195);
xnor U16625 (N_16625,N_13324,N_13322);
nor U16626 (N_16626,N_13377,N_14507);
nand U16627 (N_16627,N_13376,N_13124);
nand U16628 (N_16628,N_12341,N_14238);
nand U16629 (N_16629,N_15415,N_13735);
xor U16630 (N_16630,N_15587,N_14482);
xnor U16631 (N_16631,N_12987,N_12577);
or U16632 (N_16632,N_13059,N_15873);
nor U16633 (N_16633,N_12853,N_14121);
nor U16634 (N_16634,N_15515,N_14490);
xnor U16635 (N_16635,N_12869,N_12922);
nor U16636 (N_16636,N_12748,N_15263);
or U16637 (N_16637,N_13957,N_12278);
nand U16638 (N_16638,N_15665,N_14488);
and U16639 (N_16639,N_12736,N_13120);
and U16640 (N_16640,N_14693,N_12022);
and U16641 (N_16641,N_14783,N_14266);
and U16642 (N_16642,N_13024,N_12657);
or U16643 (N_16643,N_12296,N_12671);
or U16644 (N_16644,N_15668,N_14799);
nand U16645 (N_16645,N_13759,N_12909);
nor U16646 (N_16646,N_12190,N_12558);
and U16647 (N_16647,N_15485,N_13732);
and U16648 (N_16648,N_14089,N_13865);
nand U16649 (N_16649,N_15929,N_15004);
nand U16650 (N_16650,N_14464,N_13768);
nand U16651 (N_16651,N_12927,N_15038);
nor U16652 (N_16652,N_14601,N_14586);
xnor U16653 (N_16653,N_15254,N_15664);
xor U16654 (N_16654,N_15755,N_12311);
nor U16655 (N_16655,N_13090,N_12642);
xnor U16656 (N_16656,N_13007,N_15794);
and U16657 (N_16657,N_15061,N_13298);
or U16658 (N_16658,N_15854,N_12360);
xor U16659 (N_16659,N_14936,N_13118);
nand U16660 (N_16660,N_12863,N_15603);
xnor U16661 (N_16661,N_13111,N_15281);
xnor U16662 (N_16662,N_14851,N_12780);
nand U16663 (N_16663,N_15503,N_12893);
or U16664 (N_16664,N_13016,N_14990);
and U16665 (N_16665,N_15777,N_15963);
nand U16666 (N_16666,N_12944,N_15741);
and U16667 (N_16667,N_12816,N_14001);
nand U16668 (N_16668,N_15019,N_14811);
nand U16669 (N_16669,N_13052,N_13460);
xor U16670 (N_16670,N_14383,N_13032);
nor U16671 (N_16671,N_12132,N_13797);
nor U16672 (N_16672,N_15159,N_14231);
or U16673 (N_16673,N_12585,N_15639);
or U16674 (N_16674,N_14032,N_15089);
nand U16675 (N_16675,N_15698,N_13308);
or U16676 (N_16676,N_12032,N_12484);
nor U16677 (N_16677,N_14873,N_15943);
nor U16678 (N_16678,N_15678,N_14305);
and U16679 (N_16679,N_12443,N_14502);
or U16680 (N_16680,N_14453,N_14933);
nand U16681 (N_16681,N_15974,N_14067);
nand U16682 (N_16682,N_13968,N_14784);
nand U16683 (N_16683,N_15200,N_15541);
or U16684 (N_16684,N_14970,N_12266);
or U16685 (N_16685,N_15856,N_15531);
nand U16686 (N_16686,N_15660,N_13771);
xor U16687 (N_16687,N_14901,N_12739);
xnor U16688 (N_16688,N_14095,N_13659);
xor U16689 (N_16689,N_15486,N_12082);
xnor U16690 (N_16690,N_15783,N_13767);
or U16691 (N_16691,N_14107,N_12539);
nand U16692 (N_16692,N_12130,N_13301);
and U16693 (N_16693,N_14571,N_13559);
or U16694 (N_16694,N_13314,N_14746);
nor U16695 (N_16695,N_13762,N_15807);
nor U16696 (N_16696,N_14726,N_12306);
xor U16697 (N_16697,N_12026,N_12456);
or U16698 (N_16698,N_15793,N_13159);
nor U16699 (N_16699,N_13327,N_12466);
nor U16700 (N_16700,N_12867,N_14835);
and U16701 (N_16701,N_12478,N_12412);
xor U16702 (N_16702,N_12540,N_14651);
nor U16703 (N_16703,N_13508,N_15142);
xnor U16704 (N_16704,N_15202,N_14187);
and U16705 (N_16705,N_15947,N_14286);
xor U16706 (N_16706,N_14493,N_13049);
nor U16707 (N_16707,N_12778,N_15444);
and U16708 (N_16708,N_15598,N_12774);
nor U16709 (N_16709,N_12321,N_12169);
or U16710 (N_16710,N_14618,N_15529);
and U16711 (N_16711,N_14719,N_12752);
nor U16712 (N_16712,N_14572,N_13793);
or U16713 (N_16713,N_15742,N_12004);
or U16714 (N_16714,N_15537,N_14300);
xor U16715 (N_16715,N_13690,N_15670);
or U16716 (N_16716,N_15043,N_12006);
or U16717 (N_16717,N_14733,N_13011);
nand U16718 (N_16718,N_15139,N_15356);
xor U16719 (N_16719,N_13844,N_13898);
xnor U16720 (N_16720,N_15379,N_15233);
nand U16721 (N_16721,N_13890,N_14000);
or U16722 (N_16722,N_13502,N_13920);
nand U16723 (N_16723,N_14862,N_14718);
xnor U16724 (N_16724,N_13125,N_15306);
and U16725 (N_16725,N_14104,N_13521);
or U16726 (N_16726,N_14860,N_12848);
nand U16727 (N_16727,N_14013,N_13424);
nor U16728 (N_16728,N_15953,N_15374);
nor U16729 (N_16729,N_14128,N_15152);
or U16730 (N_16730,N_12820,N_15230);
xor U16731 (N_16731,N_14485,N_13207);
or U16732 (N_16732,N_13947,N_14532);
or U16733 (N_16733,N_15126,N_12712);
nand U16734 (N_16734,N_14782,N_13974);
nor U16735 (N_16735,N_14703,N_15937);
nand U16736 (N_16736,N_13596,N_15849);
nand U16737 (N_16737,N_12690,N_12808);
nor U16738 (N_16738,N_15169,N_14856);
or U16739 (N_16739,N_13748,N_15604);
nor U16740 (N_16740,N_15196,N_12819);
and U16741 (N_16741,N_13531,N_15021);
xor U16742 (N_16742,N_12144,N_14274);
and U16743 (N_16743,N_15700,N_13529);
and U16744 (N_16744,N_14459,N_13001);
nor U16745 (N_16745,N_12676,N_15502);
and U16746 (N_16746,N_12682,N_13150);
nand U16747 (N_16747,N_15787,N_12139);
and U16748 (N_16748,N_13670,N_13162);
nor U16749 (N_16749,N_13330,N_12458);
and U16750 (N_16750,N_15754,N_14840);
nor U16751 (N_16751,N_12658,N_14600);
and U16752 (N_16752,N_12010,N_13501);
xor U16753 (N_16753,N_15916,N_15343);
xor U16754 (N_16754,N_13467,N_15057);
nand U16755 (N_16755,N_13093,N_15002);
or U16756 (N_16756,N_15820,N_14049);
xnor U16757 (N_16757,N_14079,N_12647);
nor U16758 (N_16758,N_15314,N_14289);
and U16759 (N_16759,N_12348,N_13316);
nor U16760 (N_16760,N_12746,N_15441);
nand U16761 (N_16761,N_12882,N_12454);
xnor U16762 (N_16762,N_15826,N_14388);
and U16763 (N_16763,N_12471,N_12612);
xor U16764 (N_16764,N_15026,N_12104);
nand U16765 (N_16765,N_14295,N_14596);
xnor U16766 (N_16766,N_15651,N_12075);
and U16767 (N_16767,N_13312,N_15209);
or U16768 (N_16768,N_12804,N_15114);
xor U16769 (N_16769,N_15561,N_12423);
nand U16770 (N_16770,N_15187,N_12717);
nor U16771 (N_16771,N_13099,N_12749);
and U16772 (N_16772,N_14590,N_15034);
or U16773 (N_16773,N_13524,N_15301);
nand U16774 (N_16774,N_14674,N_13339);
and U16775 (N_16775,N_15972,N_12373);
xor U16776 (N_16776,N_15674,N_12009);
or U16777 (N_16777,N_15753,N_15928);
nor U16778 (N_16778,N_12085,N_13546);
xor U16779 (N_16779,N_15575,N_14876);
or U16780 (N_16780,N_15386,N_12493);
nand U16781 (N_16781,N_14014,N_15113);
and U16782 (N_16782,N_14186,N_14912);
nand U16783 (N_16783,N_14749,N_13630);
xor U16784 (N_16784,N_14887,N_14402);
nor U16785 (N_16785,N_12935,N_12187);
and U16786 (N_16786,N_14902,N_12934);
or U16787 (N_16787,N_14511,N_12634);
and U16788 (N_16788,N_14988,N_14686);
nand U16789 (N_16789,N_14747,N_14029);
xor U16790 (N_16790,N_12038,N_13756);
xor U16791 (N_16791,N_15647,N_15546);
and U16792 (N_16792,N_15638,N_13789);
nand U16793 (N_16793,N_12858,N_14777);
xnor U16794 (N_16794,N_13221,N_13964);
or U16795 (N_16795,N_14035,N_13281);
or U16796 (N_16796,N_13628,N_13664);
nand U16797 (N_16797,N_13247,N_15253);
or U16798 (N_16798,N_14611,N_12131);
and U16799 (N_16799,N_14986,N_13528);
or U16800 (N_16800,N_12497,N_13145);
nor U16801 (N_16801,N_14261,N_12307);
nor U16802 (N_16802,N_13476,N_13045);
xor U16803 (N_16803,N_14984,N_15903);
or U16804 (N_16804,N_14031,N_12366);
xor U16805 (N_16805,N_13069,N_12274);
nor U16806 (N_16806,N_12194,N_13571);
nand U16807 (N_16807,N_13896,N_12308);
and U16808 (N_16808,N_14465,N_15110);
nor U16809 (N_16809,N_12428,N_13971);
xnor U16810 (N_16810,N_13200,N_12091);
or U16811 (N_16811,N_13495,N_12151);
nand U16812 (N_16812,N_14996,N_12476);
xnor U16813 (N_16813,N_15482,N_13777);
and U16814 (N_16814,N_12042,N_15479);
and U16815 (N_16815,N_14736,N_12284);
and U16816 (N_16816,N_15397,N_12564);
nand U16817 (N_16817,N_13368,N_14603);
or U16818 (N_16818,N_14781,N_15900);
and U16819 (N_16819,N_15643,N_13439);
and U16820 (N_16820,N_14020,N_12133);
nor U16821 (N_16821,N_15610,N_14091);
and U16822 (N_16822,N_15775,N_14053);
and U16823 (N_16823,N_12607,N_14379);
nor U16824 (N_16824,N_13038,N_13379);
xnor U16825 (N_16825,N_15962,N_13388);
or U16826 (N_16826,N_12630,N_15048);
xor U16827 (N_16827,N_12029,N_14916);
and U16828 (N_16828,N_14881,N_14562);
xnor U16829 (N_16829,N_14145,N_14615);
and U16830 (N_16830,N_14555,N_13275);
nand U16831 (N_16831,N_15990,N_13110);
xor U16832 (N_16832,N_13806,N_14278);
and U16833 (N_16833,N_15614,N_15536);
and U16834 (N_16834,N_13063,N_14929);
or U16835 (N_16835,N_12613,N_15350);
and U16836 (N_16836,N_13219,N_15337);
or U16837 (N_16837,N_14218,N_12071);
nand U16838 (N_16838,N_14125,N_14235);
xor U16839 (N_16839,N_15931,N_13015);
and U16840 (N_16840,N_13720,N_13879);
xor U16841 (N_16841,N_14582,N_14372);
nor U16842 (N_16842,N_12389,N_12589);
xor U16843 (N_16843,N_13307,N_13217);
xor U16844 (N_16844,N_13058,N_13289);
xnor U16845 (N_16845,N_15358,N_15832);
nand U16846 (N_16846,N_14090,N_12711);
and U16847 (N_16847,N_13876,N_15530);
or U16848 (N_16848,N_13712,N_12276);
or U16849 (N_16849,N_14512,N_15823);
nor U16850 (N_16850,N_14377,N_15074);
nor U16851 (N_16851,N_14541,N_12622);
nor U16852 (N_16852,N_13824,N_15692);
or U16853 (N_16853,N_12870,N_15785);
and U16854 (N_16854,N_15499,N_12592);
and U16855 (N_16855,N_15579,N_15453);
nand U16856 (N_16856,N_12249,N_15666);
xor U16857 (N_16857,N_13466,N_15392);
or U16858 (N_16858,N_12416,N_12697);
nor U16859 (N_16859,N_13347,N_14059);
nor U16860 (N_16860,N_12788,N_15802);
nor U16861 (N_16861,N_15434,N_15240);
xnor U16862 (N_16862,N_13845,N_14320);
and U16863 (N_16863,N_12631,N_15672);
xnor U16864 (N_16864,N_13928,N_14263);
or U16865 (N_16865,N_15862,N_12913);
xnor U16866 (N_16866,N_12280,N_13471);
and U16867 (N_16867,N_14948,N_12380);
and U16868 (N_16868,N_14855,N_12418);
and U16869 (N_16869,N_13306,N_12359);
or U16870 (N_16870,N_15695,N_13572);
or U16871 (N_16871,N_14179,N_13480);
nor U16872 (N_16872,N_15338,N_13996);
and U16873 (N_16873,N_14017,N_12372);
or U16874 (N_16874,N_15707,N_15960);
or U16875 (N_16875,N_15524,N_13605);
nor U16876 (N_16876,N_15385,N_12202);
or U16877 (N_16877,N_13877,N_13389);
or U16878 (N_16878,N_13923,N_13104);
or U16879 (N_16879,N_14354,N_13899);
nand U16880 (N_16880,N_13351,N_14200);
xnor U16881 (N_16881,N_13728,N_14967);
or U16882 (N_16882,N_13071,N_13859);
nor U16883 (N_16883,N_15757,N_13833);
or U16884 (N_16884,N_12721,N_12301);
or U16885 (N_16885,N_12624,N_14027);
xnor U16886 (N_16886,N_15790,N_14885);
or U16887 (N_16887,N_12797,N_14206);
and U16888 (N_16888,N_15636,N_13364);
nor U16889 (N_16889,N_13555,N_15364);
and U16890 (N_16890,N_12365,N_14715);
and U16891 (N_16891,N_13569,N_13916);
xor U16892 (N_16892,N_13293,N_14400);
nand U16893 (N_16893,N_13002,N_13026);
or U16894 (N_16894,N_14501,N_15677);
nand U16895 (N_16895,N_15786,N_12094);
and U16896 (N_16896,N_13905,N_15302);
or U16897 (N_16897,N_15682,N_12488);
nor U16898 (N_16898,N_13083,N_13614);
or U16899 (N_16899,N_12295,N_13692);
nor U16900 (N_16900,N_13311,N_13268);
nand U16901 (N_16901,N_12475,N_13592);
or U16902 (N_16902,N_13929,N_12453);
xnor U16903 (N_16903,N_13490,N_15979);
xnor U16904 (N_16904,N_12324,N_13348);
xor U16905 (N_16905,N_15662,N_14893);
or U16906 (N_16906,N_13319,N_12400);
xor U16907 (N_16907,N_15000,N_13758);
or U16908 (N_16908,N_14926,N_14219);
xnor U16909 (N_16909,N_12782,N_13689);
and U16910 (N_16910,N_15265,N_14432);
xnor U16911 (N_16911,N_15518,N_13277);
xnor U16912 (N_16912,N_15615,N_12541);
nor U16913 (N_16913,N_13557,N_15069);
or U16914 (N_16914,N_15406,N_12535);
nor U16915 (N_16915,N_14976,N_14298);
or U16916 (N_16916,N_12762,N_15669);
nand U16917 (N_16917,N_14270,N_14961);
or U16918 (N_16918,N_12936,N_12641);
nand U16919 (N_16919,N_12062,N_13854);
or U16920 (N_16920,N_13641,N_14909);
and U16921 (N_16921,N_12584,N_15743);
nor U16922 (N_16922,N_13487,N_12353);
or U16923 (N_16923,N_15767,N_12977);
nand U16924 (N_16924,N_15954,N_13624);
nand U16925 (N_16925,N_15942,N_14433);
nand U16926 (N_16926,N_14974,N_15791);
and U16927 (N_16927,N_12567,N_13452);
nand U16928 (N_16928,N_13440,N_15890);
nand U16929 (N_16929,N_14191,N_14504);
xor U16930 (N_16930,N_15247,N_14999);
nand U16931 (N_16931,N_15663,N_15303);
and U16932 (N_16932,N_12595,N_14026);
and U16933 (N_16933,N_12783,N_13900);
or U16934 (N_16934,N_13542,N_15251);
nand U16935 (N_16935,N_14015,N_13112);
nand U16936 (N_16936,N_14963,N_14642);
nor U16937 (N_16937,N_13622,N_14551);
nand U16938 (N_16938,N_14471,N_13917);
xor U16939 (N_16939,N_12537,N_15046);
nand U16940 (N_16940,N_15918,N_14821);
xor U16941 (N_16941,N_15320,N_13585);
or U16942 (N_16942,N_13510,N_14684);
and U16943 (N_16943,N_12198,N_12001);
xnor U16944 (N_16944,N_12420,N_12035);
and U16945 (N_16945,N_13851,N_15527);
nor U16946 (N_16946,N_15175,N_14808);
nand U16947 (N_16947,N_12025,N_13536);
nor U16948 (N_16948,N_14997,N_14768);
nand U16949 (N_16949,N_14609,N_14807);
or U16950 (N_16950,N_15595,N_15654);
and U16951 (N_16951,N_15178,N_12937);
and U16952 (N_16952,N_12379,N_15075);
and U16953 (N_16953,N_14529,N_12170);
and U16954 (N_16954,N_12270,N_15552);
nor U16955 (N_16955,N_14332,N_15964);
nor U16956 (N_16956,N_12505,N_15353);
nand U16957 (N_16957,N_14030,N_14714);
nor U16958 (N_16958,N_14691,N_12683);
nand U16959 (N_16959,N_14861,N_14253);
and U16960 (N_16960,N_15684,N_14985);
and U16961 (N_16961,N_13469,N_14897);
xor U16962 (N_16962,N_12667,N_14403);
nor U16963 (N_16963,N_14847,N_15206);
nand U16964 (N_16964,N_12679,N_15585);
xor U16965 (N_16965,N_12487,N_15730);
nand U16966 (N_16966,N_14051,N_12070);
xor U16967 (N_16967,N_14949,N_14404);
or U16968 (N_16968,N_12113,N_15456);
or U16969 (N_16969,N_12445,N_13814);
and U16970 (N_16970,N_13635,N_14753);
xor U16971 (N_16971,N_12521,N_14398);
or U16972 (N_16972,N_14131,N_14474);
or U16973 (N_16973,N_15429,N_13636);
nand U16974 (N_16974,N_15725,N_12378);
xnor U16975 (N_16975,N_14772,N_15400);
or U16976 (N_16976,N_12179,N_14945);
and U16977 (N_16977,N_12336,N_14526);
xnor U16978 (N_16978,N_15237,N_12349);
nand U16979 (N_16979,N_12674,N_15435);
nand U16980 (N_16980,N_14889,N_14589);
or U16981 (N_16981,N_15548,N_14787);
or U16982 (N_16982,N_12229,N_12063);
and U16983 (N_16983,N_15681,N_13443);
or U16984 (N_16984,N_12072,N_14785);
and U16985 (N_16985,N_14778,N_13681);
nand U16986 (N_16986,N_12655,N_12695);
nor U16987 (N_16987,N_12199,N_14193);
nor U16988 (N_16988,N_12929,N_12596);
and U16989 (N_16989,N_15882,N_15489);
xnor U16990 (N_16990,N_15171,N_14406);
xor U16991 (N_16991,N_13484,N_15547);
or U16992 (N_16992,N_12111,N_14757);
or U16993 (N_16993,N_12905,N_14358);
nand U16994 (N_16994,N_12786,N_13586);
nand U16995 (N_16995,N_13766,N_13737);
or U16996 (N_16996,N_15649,N_13296);
and U16997 (N_16997,N_14444,N_15907);
or U16998 (N_16998,N_15198,N_14294);
and U16999 (N_16999,N_12516,N_14695);
xor U17000 (N_17000,N_14462,N_13072);
xnor U17001 (N_17001,N_13554,N_12868);
and U17002 (N_17002,N_12672,N_12940);
and U17003 (N_17003,N_14712,N_15733);
xor U17004 (N_17004,N_14265,N_12138);
or U17005 (N_17005,N_12586,N_13716);
nor U17006 (N_17006,N_13779,N_15312);
or U17007 (N_17007,N_13795,N_13654);
nand U17008 (N_17008,N_14699,N_13601);
nand U17009 (N_17009,N_14794,N_14564);
nor U17010 (N_17010,N_13153,N_12079);
nand U17011 (N_17011,N_15815,N_15090);
nand U17012 (N_17012,N_13802,N_12668);
or U17013 (N_17013,N_12320,N_12733);
xor U17014 (N_17014,N_14106,N_12841);
and U17015 (N_17015,N_14247,N_12765);
xor U17016 (N_17016,N_13374,N_13776);
nor U17017 (N_17017,N_13123,N_13129);
or U17018 (N_17018,N_13441,N_13168);
xor U17019 (N_17019,N_12873,N_15919);
nand U17020 (N_17020,N_14475,N_13522);
and U17021 (N_17021,N_15008,N_15273);
nor U17022 (N_17022,N_12255,N_13950);
or U17023 (N_17023,N_15563,N_13282);
nand U17024 (N_17024,N_12643,N_13942);
and U17025 (N_17025,N_14301,N_13506);
nand U17026 (N_17026,N_13738,N_13178);
and U17027 (N_17027,N_13984,N_12175);
or U17028 (N_17028,N_12766,N_13573);
or U17029 (N_17029,N_14055,N_15056);
nand U17030 (N_17030,N_14407,N_15999);
nand U17031 (N_17031,N_12333,N_13978);
nor U17032 (N_17032,N_15213,N_12215);
and U17033 (N_17033,N_15967,N_15276);
xnor U17034 (N_17034,N_15831,N_15612);
or U17035 (N_17035,N_14773,N_13757);
and U17036 (N_17036,N_15550,N_15394);
and U17037 (N_17037,N_13274,N_13509);
or U17038 (N_17038,N_12823,N_13196);
and U17039 (N_17039,N_14355,N_12110);
nand U17040 (N_17040,N_12430,N_12691);
nor U17041 (N_17041,N_15399,N_14148);
and U17042 (N_17042,N_15329,N_13860);
nand U17043 (N_17043,N_15150,N_12680);
nor U17044 (N_17044,N_12315,N_12547);
or U17045 (N_17045,N_14380,N_12148);
and U17046 (N_17046,N_14647,N_14047);
nand U17047 (N_17047,N_13193,N_13564);
nor U17048 (N_17048,N_13455,N_15290);
and U17049 (N_17049,N_15555,N_15623);
xnor U17050 (N_17050,N_12529,N_13609);
or U17051 (N_17051,N_14758,N_15853);
or U17052 (N_17052,N_13444,N_13869);
xnor U17053 (N_17053,N_15204,N_12941);
nand U17054 (N_17054,N_15474,N_13336);
or U17055 (N_17055,N_14487,N_12116);
nor U17056 (N_17056,N_12890,N_13491);
or U17057 (N_17057,N_15009,N_14230);
and U17058 (N_17058,N_13587,N_14319);
nand U17059 (N_17059,N_13299,N_13742);
nand U17060 (N_17060,N_12472,N_13214);
nand U17061 (N_17061,N_12735,N_14024);
xor U17062 (N_17062,N_13588,N_14328);
xor U17063 (N_17063,N_12325,N_13393);
nor U17064 (N_17064,N_13468,N_12137);
nand U17065 (N_17065,N_13966,N_15452);
xnor U17066 (N_17066,N_14801,N_12367);
and U17067 (N_17067,N_15185,N_15134);
xnor U17068 (N_17068,N_15375,N_15863);
nand U17069 (N_17069,N_15299,N_13997);
or U17070 (N_17070,N_13581,N_13447);
and U17071 (N_17071,N_15704,N_12237);
nand U17072 (N_17072,N_14272,N_12623);
nand U17073 (N_17073,N_14705,N_14980);
or U17074 (N_17074,N_14139,N_15799);
xnor U17075 (N_17075,N_15421,N_12599);
and U17076 (N_17076,N_15067,N_14837);
xor U17077 (N_17077,N_13582,N_13132);
xnor U17078 (N_17078,N_13607,N_12102);
and U17079 (N_17079,N_15477,N_14057);
nor U17080 (N_17080,N_14392,N_13233);
xor U17081 (N_17081,N_13492,N_15597);
xnor U17082 (N_17082,N_12069,N_15628);
nand U17083 (N_17083,N_13435,N_12618);
nor U17084 (N_17084,N_15965,N_14142);
and U17085 (N_17085,N_15140,N_14575);
and U17086 (N_17086,N_14790,N_13841);
nor U17087 (N_17087,N_15468,N_15939);
xnor U17088 (N_17088,N_12468,N_12632);
or U17089 (N_17089,N_15297,N_13673);
or U17090 (N_17090,N_14848,N_12965);
nand U17091 (N_17091,N_14565,N_15661);
and U17092 (N_17092,N_13360,N_15335);
and U17093 (N_17093,N_13074,N_15215);
or U17094 (N_17094,N_15622,N_12233);
or U17095 (N_17095,N_14895,N_14102);
or U17096 (N_17096,N_15189,N_12889);
nor U17097 (N_17097,N_12211,N_13897);
nor U17098 (N_17098,N_12988,N_12500);
and U17099 (N_17099,N_14184,N_15837);
nor U17100 (N_17100,N_13745,N_15207);
nor U17101 (N_17101,N_14522,N_15163);
and U17102 (N_17102,N_14048,N_13211);
nand U17103 (N_17103,N_15958,N_12523);
or U17104 (N_17104,N_15367,N_15018);
nand U17105 (N_17105,N_13100,N_13060);
and U17106 (N_17106,N_14910,N_12015);
xnor U17107 (N_17107,N_13138,N_13932);
or U17108 (N_17108,N_15167,N_13240);
or U17109 (N_17109,N_13027,N_15272);
nor U17110 (N_17110,N_12261,N_12461);
or U17111 (N_17111,N_15286,N_13623);
or U17112 (N_17112,N_15195,N_15403);
xnor U17113 (N_17113,N_13629,N_12518);
nor U17114 (N_17114,N_14956,N_12943);
xnor U17115 (N_17115,N_13098,N_15238);
xnor U17116 (N_17116,N_14907,N_12829);
or U17117 (N_17117,N_12591,N_12835);
nor U17118 (N_17118,N_15208,N_13672);
nor U17119 (N_17119,N_12049,N_15214);
nand U17120 (N_17120,N_13773,N_14225);
nor U17121 (N_17121,N_12376,N_14975);
and U17122 (N_17122,N_15333,N_15607);
xor U17123 (N_17123,N_13086,N_15589);
and U17124 (N_17124,N_15843,N_15729);
and U17125 (N_17125,N_15880,N_14882);
and U17126 (N_17126,N_12840,N_12124);
and U17127 (N_17127,N_14663,N_13754);
and U17128 (N_17128,N_14112,N_15912);
nor U17129 (N_17129,N_15264,N_13683);
and U17130 (N_17130,N_12790,N_14216);
or U17131 (N_17131,N_14450,N_13599);
or U17132 (N_17132,N_12096,N_15062);
xnor U17133 (N_17133,N_15657,N_13943);
nand U17134 (N_17134,N_15014,N_13355);
nand U17135 (N_17135,N_15042,N_13028);
or U17136 (N_17136,N_14256,N_14852);
or U17137 (N_17137,N_15945,N_14672);
nor U17138 (N_17138,N_14415,N_12555);
nor U17139 (N_17139,N_13926,N_14734);
nand U17140 (N_17140,N_13208,N_15519);
nor U17141 (N_17141,N_12951,N_13839);
or U17142 (N_17142,N_12388,N_13537);
and U17143 (N_17143,N_12252,N_14236);
or U17144 (N_17144,N_13838,N_15534);
nand U17145 (N_17145,N_15016,N_14992);
nand U17146 (N_17146,N_12300,N_13354);
or U17147 (N_17147,N_12134,N_12031);
nor U17148 (N_17148,N_15927,N_15500);
or U17149 (N_17149,N_13337,N_12849);
nor U17150 (N_17150,N_15496,N_15460);
or U17151 (N_17151,N_12317,N_14937);
xnor U17152 (N_17152,N_14676,N_15749);
nor U17153 (N_17153,N_15228,N_12742);
xor U17154 (N_17154,N_13626,N_15810);
and U17155 (N_17155,N_14819,N_15141);
xnor U17156 (N_17156,N_13097,N_15619);
nand U17157 (N_17157,N_13018,N_15147);
xor U17158 (N_17158,N_13809,N_14585);
xnor U17159 (N_17159,N_13637,N_15850);
or U17160 (N_17160,N_14899,N_12975);
nand U17161 (N_17161,N_12917,N_12218);
nor U17162 (N_17162,N_14359,N_13398);
nor U17163 (N_17163,N_15512,N_15262);
xnor U17164 (N_17164,N_15305,N_12572);
nor U17165 (N_17165,N_13500,N_13128);
nand U17166 (N_17166,N_12726,N_15744);
xnor U17167 (N_17167,N_13741,N_14875);
or U17168 (N_17168,N_13486,N_12173);
nand U17169 (N_17169,N_13255,N_14039);
and U17170 (N_17170,N_15715,N_13552);
or U17171 (N_17171,N_14616,N_14888);
or U17172 (N_17172,N_13260,N_12553);
nand U17173 (N_17173,N_14237,N_15109);
nand U17174 (N_17174,N_12673,N_15369);
xor U17175 (N_17175,N_14688,N_15591);
nand U17176 (N_17176,N_14491,N_15780);
and U17177 (N_17177,N_15111,N_14756);
or U17178 (N_17178,N_15462,N_12245);
nor U17179 (N_17179,N_12086,N_15473);
xor U17180 (N_17180,N_14496,N_13979);
and U17181 (N_17181,N_15341,N_13988);
nand U17182 (N_17182,N_13965,N_15540);
nand U17183 (N_17183,N_14792,N_12661);
and U17184 (N_17184,N_15160,N_12210);
xnor U17185 (N_17185,N_14652,N_13411);
and U17186 (N_17186,N_14078,N_13658);
and U17187 (N_17187,N_15203,N_13215);
nor U17188 (N_17188,N_15621,N_15222);
or U17189 (N_17189,N_14765,N_15634);
and U17190 (N_17190,N_14412,N_13363);
xnor U17191 (N_17191,N_14685,N_13885);
and U17192 (N_17192,N_12081,N_13212);
xnor U17193 (N_17193,N_14061,N_12178);
nand U17194 (N_17194,N_12013,N_12312);
or U17195 (N_17195,N_12875,N_14966);
nor U17196 (N_17196,N_15776,N_12646);
and U17197 (N_17197,N_14149,N_15839);
or U17198 (N_17198,N_13387,N_15227);
or U17199 (N_17199,N_15351,N_13359);
nand U17200 (N_17200,N_15510,N_13371);
and U17201 (N_17201,N_13731,N_12963);
or U17202 (N_17202,N_13765,N_13369);
nor U17203 (N_17203,N_14367,N_12322);
and U17204 (N_17204,N_15006,N_13874);
and U17205 (N_17205,N_15304,N_13191);
and U17206 (N_17206,N_15065,N_15764);
nand U17207 (N_17207,N_12128,N_15135);
or U17208 (N_17208,N_14890,N_12236);
nand U17209 (N_17209,N_14626,N_12318);
xor U17210 (N_17210,N_12581,N_15756);
or U17211 (N_17211,N_15282,N_12639);
nor U17212 (N_17212,N_14234,N_13230);
nor U17213 (N_17213,N_15829,N_12763);
or U17214 (N_17214,N_14506,N_14524);
or U17215 (N_17215,N_13567,N_13512);
xor U17216 (N_17216,N_15079,N_12709);
nor U17217 (N_17217,N_13680,N_12561);
nor U17218 (N_17218,N_13515,N_12153);
nor U17219 (N_17219,N_13821,N_15594);
and U17220 (N_17220,N_13270,N_14751);
or U17221 (N_17221,N_15713,N_14620);
nor U17222 (N_17222,N_13094,N_15992);
xor U17223 (N_17223,N_15691,N_12386);
nand U17224 (N_17224,N_14716,N_14479);
nor U17225 (N_17225,N_14643,N_15432);
nand U17226 (N_17226,N_14291,N_13051);
or U17227 (N_17227,N_14619,N_14689);
nand U17228 (N_17228,N_13786,N_15395);
nand U17229 (N_17229,N_15897,N_15488);
nor U17230 (N_17230,N_12504,N_12510);
or U17231 (N_17231,N_14421,N_12744);
xor U17232 (N_17232,N_13687,N_13812);
nor U17233 (N_17233,N_13846,N_15449);
and U17234 (N_17234,N_12902,N_14877);
xor U17235 (N_17235,N_12402,N_15340);
xor U17236 (N_17236,N_15464,N_13551);
nand U17237 (N_17237,N_12201,N_15737);
xor U17238 (N_17238,N_13578,N_12958);
and U17239 (N_17239,N_12666,N_13334);
or U17240 (N_17240,N_12046,N_15509);
xor U17241 (N_17241,N_12970,N_13078);
and U17242 (N_17242,N_14632,N_12775);
xor U17243 (N_17243,N_12304,N_15361);
nor U17244 (N_17244,N_15789,N_12334);
nor U17245 (N_17245,N_12383,N_14308);
xor U17246 (N_17246,N_13082,N_12740);
and U17247 (N_17247,N_12346,N_13982);
nand U17248 (N_17248,N_15223,N_13575);
or U17249 (N_17249,N_14390,N_12757);
or U17250 (N_17250,N_12387,N_13390);
and U17251 (N_17251,N_14973,N_13252);
nand U17252 (N_17252,N_15578,N_13457);
or U17253 (N_17253,N_14644,N_13273);
and U17254 (N_17254,N_15719,N_12205);
or U17255 (N_17255,N_12777,N_14769);
or U17256 (N_17256,N_15797,N_14667);
nor U17257 (N_17257,N_15675,N_13454);
nor U17258 (N_17258,N_13704,N_14183);
nor U17259 (N_17259,N_14162,N_12285);
nand U17260 (N_17260,N_15991,N_12609);
nor U17261 (N_17261,N_13121,N_14069);
and U17262 (N_17262,N_13709,N_13901);
nor U17263 (N_17263,N_12677,N_14823);
nand U17264 (N_17264,N_15052,N_14174);
nand U17265 (N_17265,N_15985,N_15705);
nand U17266 (N_17266,N_14375,N_14068);
and U17267 (N_17267,N_15987,N_13107);
and U17268 (N_17268,N_13225,N_12847);
nand U17269 (N_17269,N_12362,N_13474);
and U17270 (N_17270,N_14427,N_15039);
nor U17271 (N_17271,N_13803,N_13358);
nand U17272 (N_17272,N_12696,N_14483);
xor U17273 (N_17273,N_12242,N_13005);
or U17274 (N_17274,N_15545,N_15520);
nor U17275 (N_17275,N_12191,N_15235);
nand U17276 (N_17276,N_15814,N_15128);
nand U17277 (N_17277,N_14426,N_12483);
nand U17278 (N_17278,N_15165,N_13057);
nand U17279 (N_17279,N_15122,N_13995);
and U17280 (N_17280,N_12093,N_14080);
nand U17281 (N_17281,N_14129,N_12743);
nand U17282 (N_17282,N_14523,N_12845);
nor U17283 (N_17283,N_15801,N_12597);
xnor U17284 (N_17284,N_12956,N_12490);
or U17285 (N_17285,N_15322,N_14336);
nand U17286 (N_17286,N_12636,N_14573);
and U17287 (N_17287,N_15940,N_12076);
xnor U17288 (N_17288,N_14613,N_13707);
or U17289 (N_17289,N_14776,N_12832);
xor U17290 (N_17290,N_14931,N_15866);
or U17291 (N_17291,N_13017,N_15950);
nand U17292 (N_17292,N_15382,N_12154);
nand U17293 (N_17293,N_13342,N_14923);
nor U17294 (N_17294,N_14977,N_14376);
xnor U17295 (N_17295,N_14042,N_13646);
xor U17296 (N_17296,N_15523,N_12289);
or U17297 (N_17297,N_12594,N_13688);
xor U17298 (N_17298,N_15093,N_12099);
nand U17299 (N_17299,N_13648,N_15766);
and U17300 (N_17300,N_15092,N_13259);
xnor U17301 (N_17301,N_15922,N_14156);
nand U17302 (N_17302,N_14478,N_13023);
and U17303 (N_17303,N_14438,N_12891);
xor U17304 (N_17304,N_13976,N_13639);
nand U17305 (N_17305,N_12897,N_15760);
nor U17306 (N_17306,N_14979,N_14476);
and U17307 (N_17307,N_15326,N_14094);
and U17308 (N_17308,N_14621,N_13328);
or U17309 (N_17309,N_15888,N_14177);
nor U17310 (N_17310,N_15154,N_14188);
nand U17311 (N_17311,N_14793,N_15193);
nor U17312 (N_17312,N_14356,N_12573);
nand U17313 (N_17313,N_12000,N_14292);
and U17314 (N_17314,N_14454,N_14928);
xnor U17315 (N_17315,N_15418,N_15242);
and U17316 (N_17316,N_14009,N_15557);
nand U17317 (N_17317,N_13747,N_15978);
xnor U17318 (N_17318,N_12269,N_14750);
nor U17319 (N_17319,N_12767,N_15961);
nor U17320 (N_17320,N_15221,N_13647);
nor U17321 (N_17321,N_14853,N_12626);
xnor U17322 (N_17322,N_15313,N_15846);
or U17323 (N_17323,N_13848,N_12331);
xnor U17324 (N_17324,N_14513,N_12464);
xor U17325 (N_17325,N_12811,N_13638);
and U17326 (N_17326,N_14727,N_12524);
and U17327 (N_17327,N_15145,N_12615);
nor U17328 (N_17328,N_12857,N_15845);
or U17329 (N_17329,N_12302,N_13914);
and U17330 (N_17330,N_14908,N_13410);
nand U17331 (N_17331,N_14368,N_14285);
or U17332 (N_17332,N_14834,N_14434);
and U17333 (N_17333,N_14324,N_13407);
and U17334 (N_17334,N_12192,N_13395);
or U17335 (N_17335,N_15357,N_15650);
or U17336 (N_17336,N_15886,N_15816);
xnor U17337 (N_17337,N_14640,N_15818);
xor U17338 (N_17338,N_12954,N_13294);
and U17339 (N_17339,N_14556,N_12103);
or U17340 (N_17340,N_14729,N_15917);
or U17341 (N_17341,N_12230,N_14817);
and U17342 (N_17342,N_12147,N_14366);
or U17343 (N_17343,N_13556,N_14063);
nand U17344 (N_17344,N_14500,N_13033);
or U17345 (N_17345,N_13902,N_15602);
and U17346 (N_17346,N_14058,N_12007);
and U17347 (N_17347,N_12018,N_13769);
nand U17348 (N_17348,N_12701,N_15599);
nand U17349 (N_17349,N_12184,N_13889);
nor U17350 (N_17350,N_14968,N_12444);
and U17351 (N_17351,N_14282,N_13717);
xor U17352 (N_17352,N_15892,N_15762);
or U17353 (N_17353,N_14857,N_14046);
and U17354 (N_17354,N_13519,N_15146);
or U17355 (N_17355,N_14022,N_14614);
nor U17356 (N_17356,N_15804,N_15673);
or U17357 (N_17357,N_14334,N_12506);
nor U17358 (N_17358,N_14754,N_14869);
nand U17359 (N_17359,N_12542,N_14243);
or U17360 (N_17360,N_15099,N_13504);
or U17361 (N_17361,N_14340,N_13450);
and U17362 (N_17362,N_12881,N_13332);
xor U17363 (N_17363,N_13245,N_14143);
nand U17364 (N_17364,N_12528,N_14635);
and U17365 (N_17365,N_15388,N_12549);
nor U17366 (N_17366,N_12408,N_13511);
nor U17367 (N_17367,N_14625,N_15709);
nor U17368 (N_17368,N_14255,N_14034);
and U17369 (N_17369,N_14457,N_13743);
nor U17370 (N_17370,N_13283,N_15905);
or U17371 (N_17371,N_13934,N_13238);
xor U17372 (N_17372,N_14194,N_12167);
nor U17373 (N_17373,N_14567,N_15983);
or U17374 (N_17374,N_15611,N_14919);
nor U17375 (N_17375,N_15250,N_13722);
nor U17376 (N_17376,N_13913,N_13590);
nor U17377 (N_17377,N_12287,N_14721);
or U17378 (N_17378,N_12401,N_13361);
nor U17379 (N_17379,N_13750,N_12758);
nor U17380 (N_17380,N_12580,N_12719);
and U17381 (N_17381,N_12142,N_14210);
nor U17382 (N_17382,N_14076,N_12874);
nand U17383 (N_17383,N_12822,N_15513);
or U17384 (N_17384,N_14213,N_12185);
nand U17385 (N_17385,N_13727,N_13549);
xnor U17386 (N_17386,N_14495,N_13456);
nor U17387 (N_17387,N_13167,N_14947);
nor U17388 (N_17388,N_15874,N_12852);
nand U17389 (N_17389,N_15511,N_14410);
or U17390 (N_17390,N_12217,N_13169);
or U17391 (N_17391,N_13834,N_14720);
xor U17392 (N_17392,N_12660,N_14144);
nand U17393 (N_17393,N_15549,N_15875);
nand U17394 (N_17394,N_13642,N_13202);
xor U17395 (N_17395,N_12394,N_14167);
nand U17396 (N_17396,N_14553,N_12196);
xnor U17397 (N_17397,N_14084,N_13973);
nor U17398 (N_17398,N_12292,N_12812);
or U17399 (N_17399,N_15443,N_12264);
nand U17400 (N_17400,N_12206,N_13192);
nand U17401 (N_17401,N_15570,N_13356);
or U17402 (N_17402,N_13909,N_13085);
nor U17403 (N_17403,N_14743,N_12115);
nand U17404 (N_17404,N_13241,N_12451);
nor U17405 (N_17405,N_15448,N_13220);
nor U17406 (N_17406,N_15098,N_12999);
xnor U17407 (N_17407,N_12222,N_15833);
nand U17408 (N_17408,N_15218,N_12692);
nand U17409 (N_17409,N_15334,N_14033);
xnor U17410 (N_17410,N_14514,N_15852);
nand U17411 (N_17411,N_12003,N_12056);
or U17412 (N_17412,N_14599,N_12911);
or U17413 (N_17413,N_13539,N_13560);
nor U17414 (N_17414,N_14745,N_14870);
xor U17415 (N_17415,N_13819,N_12243);
and U17416 (N_17416,N_12885,N_15553);
nand U17417 (N_17417,N_13956,N_12286);
nand U17418 (N_17418,N_12803,N_13780);
xnor U17419 (N_17419,N_15360,N_15417);
nand U17420 (N_17420,N_12329,N_15100);
xor U17421 (N_17421,N_12145,N_12792);
nor U17422 (N_17422,N_13102,N_12080);
or U17423 (N_17423,N_13203,N_14648);
nor U17424 (N_17424,N_13774,N_13325);
nor U17425 (N_17425,N_13481,N_12370);
xor U17426 (N_17426,N_14357,N_14939);
nand U17427 (N_17427,N_15558,N_12117);
nor U17428 (N_17428,N_12193,N_14713);
and U17429 (N_17429,N_13866,N_15121);
or U17430 (N_17430,N_14871,N_14311);
nand U17431 (N_17431,N_15344,N_15387);
and U17432 (N_17432,N_13621,N_15025);
and U17433 (N_17433,N_12750,N_14280);
or U17434 (N_17434,N_12773,N_14762);
or U17435 (N_17435,N_13235,N_13105);
nor U17436 (N_17436,N_14443,N_13433);
xnor U17437 (N_17437,N_12548,N_14304);
or U17438 (N_17438,N_13394,N_13442);
xor U17439 (N_17439,N_13547,N_13367);
and U17440 (N_17440,N_14260,N_12651);
xor U17441 (N_17441,N_14418,N_13949);
nor U17442 (N_17442,N_13141,N_13136);
nand U17443 (N_17443,N_14924,N_12900);
xor U17444 (N_17444,N_13861,N_12996);
or U17445 (N_17445,N_12092,N_15817);
nor U17446 (N_17446,N_13134,N_14222);
nand U17447 (N_17447,N_14668,N_12005);
nor U17448 (N_17448,N_14361,N_15243);
nor U17449 (N_17449,N_15260,N_15980);
nor U17450 (N_17450,N_15151,N_12449);
nand U17451 (N_17451,N_14012,N_14414);
xor U17452 (N_17452,N_13415,N_14558);
or U17453 (N_17453,N_13295,N_15390);
and U17454 (N_17454,N_15137,N_13228);
or U17455 (N_17455,N_13955,N_12375);
and U17456 (N_17456,N_15624,N_13050);
nand U17457 (N_17457,N_13258,N_13412);
nand U17458 (N_17458,N_12974,N_12791);
nor U17459 (N_17459,N_13715,N_15567);
or U17460 (N_17460,N_15271,N_13186);
nor U17461 (N_17461,N_12271,N_14581);
nor U17462 (N_17462,N_15277,N_12625);
xor U17463 (N_17463,N_14469,N_15697);
xor U17464 (N_17464,N_14830,N_13514);
nor U17465 (N_17465,N_12681,N_12725);
xnor U17466 (N_17466,N_15428,N_14771);
or U17467 (N_17467,N_13396,N_14043);
or U17468 (N_17468,N_13004,N_12226);
and U17469 (N_17469,N_15268,N_15440);
nand U17470 (N_17470,N_12787,N_14818);
nand U17471 (N_17471,N_12648,N_12098);
or U17472 (N_17472,N_13137,N_13498);
nor U17473 (N_17473,N_14486,N_15310);
nor U17474 (N_17474,N_14951,N_14122);
xor U17475 (N_17475,N_14711,N_14326);
and U17476 (N_17476,N_12054,N_12040);
nand U17477 (N_17477,N_12047,N_15083);
and U17478 (N_17478,N_12489,N_14365);
xor U17479 (N_17479,N_12914,N_12425);
and U17480 (N_17480,N_15855,N_14804);
xnor U17481 (N_17481,N_15702,N_15355);
or U17482 (N_17482,N_13975,N_13666);
nand U17483 (N_17483,N_14463,N_12221);
xnor U17484 (N_17484,N_12976,N_14258);
nand U17485 (N_17485,N_13931,N_15102);
and U17486 (N_17486,N_12912,N_15805);
or U17487 (N_17487,N_15278,N_14441);
nor U17488 (N_17488,N_15136,N_12698);
nand U17489 (N_17489,N_13453,N_14629);
nor U17490 (N_17490,N_14814,N_13992);
nand U17491 (N_17491,N_13154,N_12898);
or U17492 (N_17492,N_15231,N_14312);
or U17493 (N_17493,N_15280,N_15317);
or U17494 (N_17494,N_13227,N_14422);
and U17495 (N_17495,N_14240,N_13830);
or U17496 (N_17496,N_13084,N_13181);
or U17497 (N_17497,N_15010,N_15869);
nand U17498 (N_17498,N_15881,N_13595);
nand U17499 (N_17499,N_14828,N_13631);
nor U17500 (N_17500,N_13697,N_13087);
and U17501 (N_17501,N_13404,N_15212);
or U17502 (N_17502,N_12932,N_13532);
nor U17503 (N_17503,N_15044,N_13216);
and U17504 (N_17504,N_14546,N_15170);
nand U17505 (N_17505,N_12785,N_12012);
xnor U17506 (N_17506,N_12918,N_15878);
and U17507 (N_17507,N_13271,N_12730);
nand U17508 (N_17508,N_14147,N_12525);
nand U17509 (N_17509,N_12207,N_14574);
or U17510 (N_17510,N_13693,N_15608);
and U17511 (N_17511,N_14722,N_14310);
and U17512 (N_17512,N_14694,N_14577);
nor U17513 (N_17513,N_13179,N_14767);
xnor U17514 (N_17514,N_13615,N_13761);
or U17515 (N_17515,N_14314,N_14774);
or U17516 (N_17516,N_12713,N_15696);
xnor U17517 (N_17517,N_12143,N_14072);
or U17518 (N_17518,N_12554,N_15091);
or U17519 (N_17519,N_13895,N_14168);
and U17520 (N_17520,N_15934,N_15835);
nand U17521 (N_17521,N_13534,N_14455);
nand U17522 (N_17522,N_12654,N_14803);
and U17523 (N_17523,N_15522,N_14748);
and U17524 (N_17524,N_15130,N_12579);
xor U17525 (N_17525,N_15176,N_13266);
or U17526 (N_17526,N_14872,N_12818);
xnor U17527 (N_17527,N_15036,N_12409);
nor U17528 (N_17528,N_12459,N_12741);
or U17529 (N_17529,N_14991,N_15828);
or U17530 (N_17530,N_13962,N_12263);
or U17531 (N_17531,N_14583,N_15568);
nor U17532 (N_17532,N_14262,N_12253);
and U17533 (N_17533,N_14302,N_12220);
or U17534 (N_17534,N_15763,N_14152);
xor U17535 (N_17535,N_15459,N_12856);
or U17536 (N_17536,N_12290,N_12374);
or U17537 (N_17537,N_13553,N_15078);
and U17538 (N_17538,N_14101,N_14552);
nand U17539 (N_17539,N_12724,N_14867);
nor U17540 (N_17540,N_13014,N_12998);
nor U17541 (N_17541,N_14110,N_15045);
nand U17542 (N_17542,N_12126,N_15701);
nor U17543 (N_17543,N_14739,N_15133);
nor U17544 (N_17544,N_14971,N_13746);
nor U17545 (N_17545,N_12119,N_15714);
or U17546 (N_17546,N_14284,N_15957);
or U17547 (N_17547,N_13651,N_15315);
or U17548 (N_17548,N_12118,N_13999);
nor U17549 (N_17549,N_14244,N_13940);
and U17550 (N_17550,N_12964,N_14116);
or U17551 (N_17551,N_15475,N_13222);
or U17552 (N_17552,N_14669,N_12901);
nor U17553 (N_17553,N_12195,N_14189);
and U17554 (N_17554,N_13286,N_15667);
xor U17555 (N_17555,N_13209,N_14021);
or U17556 (N_17556,N_12640,N_14489);
nor U17557 (N_17557,N_12921,N_15071);
nor U17558 (N_17558,N_14232,N_13416);
and U17559 (N_17559,N_13408,N_12244);
nand U17560 (N_17560,N_15993,N_14898);
nor U17561 (N_17561,N_14363,N_12310);
nor U17562 (N_17562,N_14447,N_13723);
and U17563 (N_17563,N_12176,N_13020);
and U17564 (N_17564,N_12815,N_13000);
nor U17565 (N_17565,N_13969,N_15528);
nor U17566 (N_17566,N_15182,N_13591);
and U17567 (N_17567,N_14257,N_12435);
xnor U17568 (N_17568,N_14202,N_14906);
nand U17569 (N_17569,N_14539,N_13139);
or U17570 (N_17570,N_12448,N_15723);
nor U17571 (N_17571,N_14700,N_15236);
nand U17572 (N_17572,N_12441,N_12761);
and U17573 (N_17573,N_15308,N_13753);
nor U17574 (N_17574,N_12463,N_13721);
nor U17575 (N_17575,N_14645,N_13465);
nor U17576 (N_17576,N_14038,N_15255);
and U17577 (N_17577,N_13698,N_15848);
nor U17578 (N_17578,N_15054,N_14886);
xor U17579 (N_17579,N_15138,N_12083);
xor U17580 (N_17580,N_12146,N_13470);
nand U17581 (N_17581,N_15023,N_12227);
xor U17582 (N_17582,N_14416,N_15504);
and U17583 (N_17583,N_12182,N_13921);
xor U17584 (N_17584,N_12446,N_14993);
nand U17585 (N_17585,N_13985,N_15596);
and U17586 (N_17586,N_14041,N_13320);
and U17587 (N_17587,N_13397,N_12715);
xnor U17588 (N_17588,N_14981,N_14903);
nor U17589 (N_17589,N_12705,N_14683);
nor U17590 (N_17590,N_13790,N_12955);
nor U17591 (N_17591,N_13497,N_12659);
and U17592 (N_17592,N_12123,N_13493);
nand U17593 (N_17593,N_13385,N_14662);
and U17594 (N_17594,N_12279,N_15024);
and U17595 (N_17595,N_14195,N_14510);
and U17596 (N_17596,N_15781,N_13634);
and U17597 (N_17597,N_14273,N_14858);
nor U17598 (N_17598,N_15316,N_13784);
and U17599 (N_17599,N_15616,N_15560);
xor U17600 (N_17600,N_14134,N_14863);
and U17601 (N_17601,N_14822,N_12876);
xor U17602 (N_17602,N_12377,N_13558);
or U17603 (N_17603,N_15731,N_13925);
xor U17604 (N_17604,N_13146,N_12731);
and U17605 (N_17605,N_12465,N_15007);
nand U17606 (N_17606,N_14220,N_13140);
xnor U17607 (N_17607,N_14283,N_13494);
or U17608 (N_17608,N_13886,N_12952);
nor U17609 (N_17609,N_12200,N_13292);
xnor U17610 (N_17610,N_12020,N_13151);
nand U17611 (N_17611,N_12141,N_15232);
nor U17612 (N_17612,N_14701,N_13375);
and U17613 (N_17613,N_12687,N_15569);
or U17614 (N_17614,N_13540,N_14088);
or U17615 (N_17615,N_15330,N_13627);
or U17616 (N_17616,N_15088,N_14831);
xor U17617 (N_17617,N_13981,N_15571);
nand U17618 (N_17618,N_13155,N_15445);
xor U17619 (N_17619,N_13937,N_15118);
nand U17620 (N_17620,N_14904,N_15414);
nor U17621 (N_17621,N_15721,N_13147);
nand U17622 (N_17622,N_14759,N_15229);
and U17623 (N_17623,N_14461,N_13922);
nor U17624 (N_17624,N_14108,N_13816);
nor U17625 (N_17625,N_14399,N_15425);
and U17626 (N_17626,N_13267,N_14023);
nand U17627 (N_17627,N_12410,N_13868);
nor U17628 (N_17628,N_13184,N_14182);
or U17629 (N_17629,N_15342,N_13485);
nor U17630 (N_17630,N_13611,N_15883);
nand U17631 (N_17631,N_13870,N_13285);
or U17632 (N_17632,N_15423,N_12354);
and U17633 (N_17633,N_13863,N_14678);
and U17634 (N_17634,N_14470,N_12884);
nand U17635 (N_17635,N_14520,N_13473);
xor U17636 (N_17636,N_15909,N_14456);
nand U17637 (N_17637,N_14742,N_12583);
and U17638 (N_17638,N_15923,N_15270);
or U17639 (N_17639,N_15124,N_15752);
xnor U17640 (N_17640,N_13482,N_14568);
or U17641 (N_17641,N_12992,N_12969);
nor U17642 (N_17642,N_14955,N_13924);
or U17643 (N_17643,N_15652,N_15538);
and U17644 (N_17644,N_14841,N_14060);
and U17645 (N_17645,N_14843,N_15736);
nand U17646 (N_17646,N_15123,N_15104);
nor U17647 (N_17647,N_13261,N_14677);
nor U17648 (N_17648,N_15933,N_13065);
xor U17649 (N_17649,N_12509,N_14335);
and U17650 (N_17650,N_13061,N_15973);
or U17651 (N_17651,N_15865,N_15948);
nand U17652 (N_17652,N_14965,N_13413);
nand U17653 (N_17653,N_12755,N_14827);
or U17654 (N_17654,N_15708,N_12533);
or U17655 (N_17655,N_15465,N_12248);
or U17656 (N_17656,N_15005,N_12727);
nor U17657 (N_17657,N_12653,N_14914);
nor U17658 (N_17658,N_15339,N_13755);
nor U17659 (N_17659,N_12850,N_12838);
nor U17660 (N_17660,N_14654,N_12496);
xor U17661 (N_17661,N_12414,N_12058);
xnor U17662 (N_17662,N_12732,N_14987);
and U17663 (N_17663,N_14559,N_12427);
or U17664 (N_17664,N_14824,N_15989);
or U17665 (N_17665,N_13799,N_14442);
nor U17666 (N_17666,N_15292,N_13987);
or U17667 (N_17667,N_13650,N_15420);
nor U17668 (N_17668,N_12507,N_13810);
nand U17669 (N_17669,N_15480,N_14673);
nor U17670 (N_17670,N_13458,N_14634);
nor U17671 (N_17671,N_13633,N_14384);
nand U17672 (N_17672,N_15458,N_14120);
nor U17673 (N_17673,N_15188,N_15072);
and U17674 (N_17674,N_12155,N_13035);
and U17675 (N_17675,N_14932,N_13170);
and U17676 (N_17676,N_14056,N_14246);
and U17677 (N_17677,N_15625,N_12635);
xnor U17678 (N_17678,N_14011,N_14019);
nand U17679 (N_17679,N_12527,N_12895);
xor U17680 (N_17680,N_13941,N_13602);
or U17681 (N_17681,N_14891,N_14866);
and U17682 (N_17682,N_14323,N_15431);
nand U17683 (N_17683,N_15037,N_13970);
and U17684 (N_17684,N_15956,N_12442);
xor U17685 (N_17685,N_15679,N_12293);
xor U17686 (N_17686,N_15501,N_13983);
nand U17687 (N_17687,N_12729,N_13734);
xnor U17688 (N_17688,N_13594,N_14592);
or U17689 (N_17689,N_15911,N_15562);
or U17690 (N_17690,N_15080,N_13021);
nand U17691 (N_17691,N_14081,N_13574);
and U17692 (N_17692,N_13593,N_14329);
and U17693 (N_17693,N_15319,N_12980);
xnor U17694 (N_17694,N_14964,N_12241);
and U17695 (N_17695,N_12503,N_15544);
nor U17696 (N_17696,N_15642,N_15470);
and U17697 (N_17697,N_13381,N_15493);
and U17698 (N_17698,N_15031,N_12260);
nor U17699 (N_17699,N_15857,N_15436);
nor U17700 (N_17700,N_14085,N_13073);
xor U17701 (N_17701,N_13505,N_13794);
or U17702 (N_17702,N_14563,N_14549);
nand U17703 (N_17703,N_12371,N_14171);
and U17704 (N_17704,N_15689,N_12422);
nand U17705 (N_17705,N_12021,N_12156);
nor U17706 (N_17706,N_13089,N_12240);
and U17707 (N_17707,N_13972,N_15127);
nor U17708 (N_17708,N_15457,N_13656);
nor U17709 (N_17709,N_12514,N_14878);
nand U17710 (N_17710,N_13733,N_12531);
and U17711 (N_17711,N_13175,N_13694);
and U17712 (N_17712,N_15219,N_14605);
or U17713 (N_17713,N_13291,N_14172);
and U17714 (N_17714,N_15659,N_15871);
or U17715 (N_17715,N_15644,N_12188);
nand U17716 (N_17716,N_12997,N_14702);
or U17717 (N_17717,N_12257,N_14744);
nor U17718 (N_17718,N_15366,N_13008);
nor U17719 (N_17719,N_14435,N_12916);
nand U17720 (N_17720,N_12810,N_15106);
or U17721 (N_17721,N_14473,N_12059);
nor U17722 (N_17722,N_14391,N_14073);
xnor U17723 (N_17723,N_14865,N_13091);
xnor U17724 (N_17724,N_15058,N_13643);
nand U17725 (N_17725,N_14036,N_15258);
xor U17726 (N_17726,N_13157,N_13545);
and U17727 (N_17727,N_13817,N_14140);
and U17728 (N_17728,N_14725,N_14249);
and U17729 (N_17729,N_15788,N_13278);
xnor U17730 (N_17730,N_15491,N_12770);
and U17731 (N_17731,N_13729,N_14849);
and U17732 (N_17732,N_15975,N_15630);
and U17733 (N_17733,N_15439,N_12560);
nor U17734 (N_17734,N_14832,N_15613);
nor U17735 (N_17735,N_12172,N_12150);
and U17736 (N_17736,N_14838,N_13256);
xor U17737 (N_17737,N_15422,N_12915);
and U17738 (N_17738,N_13302,N_12361);
nand U17739 (N_17739,N_12961,N_13242);
or U17740 (N_17740,N_14584,N_15257);
and U17741 (N_17741,N_13565,N_13908);
nor U17742 (N_17742,N_13148,N_15739);
nand U17743 (N_17743,N_14530,N_14007);
or U17744 (N_17744,N_13791,N_13253);
nand U17745 (N_17745,N_14874,N_14006);
nor U17746 (N_17746,N_13185,N_15295);
or U17747 (N_17747,N_15192,N_13101);
or U17748 (N_17748,N_12606,N_12313);
nand U17749 (N_17749,N_14969,N_13405);
xnor U17750 (N_17750,N_14646,N_14229);
and U17751 (N_17751,N_12258,N_15469);
and U17752 (N_17752,N_13231,N_14978);
nand U17753 (N_17753,N_12947,N_12407);
xnor U17754 (N_17754,N_15626,N_14982);
and U17755 (N_17755,N_12396,N_13436);
and U17756 (N_17756,N_14820,N_14670);
nor U17757 (N_17757,N_15478,N_13429);
nor U17758 (N_17758,N_12575,N_13418);
nor U17759 (N_17759,N_13177,N_14595);
or U17760 (N_17760,N_14508,N_13194);
nand U17761 (N_17761,N_13272,N_15050);
xor U17762 (N_17762,N_13991,N_13434);
and U17763 (N_17763,N_15177,N_12628);
or U17764 (N_17764,N_14394,N_13691);
xor U17765 (N_17765,N_15131,N_15727);
nand U17766 (N_17766,N_12251,N_15161);
or U17767 (N_17767,N_14296,N_15283);
nor U17768 (N_17768,N_12745,N_12718);
nand U17769 (N_17769,N_15096,N_12828);
or U17770 (N_17770,N_12450,N_15631);
nand U17771 (N_17771,N_14307,N_14630);
nor U17772 (N_17772,N_13382,N_14989);
xor U17773 (N_17773,N_14953,N_12262);
or U17774 (N_17774,N_15710,N_13329);
or U17775 (N_17775,N_12949,N_13604);
or U17776 (N_17776,N_14894,N_12764);
and U17777 (N_17777,N_12152,N_12769);
xnor U17778 (N_17778,N_14170,N_15889);
and U17779 (N_17779,N_15813,N_15205);
xnor U17780 (N_17780,N_15769,N_15971);
xor U17781 (N_17781,N_12605,N_13606);
nand U17782 (N_17782,N_12084,N_14141);
or U17783 (N_17783,N_12268,N_12950);
xnor U17784 (N_17784,N_14940,N_12566);
xnor U17785 (N_17785,N_13265,N_15157);
or U17786 (N_17786,N_14239,N_15930);
xor U17787 (N_17787,N_15906,N_15249);
nand U17788 (N_17788,N_13980,N_14763);
or U17789 (N_17789,N_15451,N_13366);
nand U17790 (N_17790,N_12055,N_15576);
nor U17791 (N_17791,N_15402,N_15676);
nand U17792 (N_17792,N_14706,N_13618);
and U17793 (N_17793,N_12953,N_12662);
nor U17794 (N_17794,N_12568,N_15774);
xnor U17795 (N_17795,N_15505,N_14938);
nor U17796 (N_17796,N_15543,N_12519);
nand U17797 (N_17797,N_13103,N_15836);
xor U17798 (N_17798,N_13419,N_14264);
or U17799 (N_17799,N_13951,N_13662);
or U17800 (N_17800,N_14178,N_13597);
or U17801 (N_17801,N_12486,N_13335);
xor U17802 (N_17802,N_15656,N_13881);
and U17803 (N_17803,N_13703,N_13835);
nor U17804 (N_17804,N_12298,N_15618);
nand U17805 (N_17805,N_12108,N_12368);
nor U17806 (N_17806,N_13449,N_12074);
nand U17807 (N_17807,N_15291,N_15632);
nor U17808 (N_17808,N_15033,N_13257);
nor U17809 (N_17809,N_14631,N_13279);
nand U17810 (N_17810,N_12836,N_15107);
and U17811 (N_17811,N_14064,N_12866);
nor U17812 (N_17812,N_14111,N_13198);
xor U17813 (N_17813,N_12545,N_15289);
xor U17814 (N_17814,N_13464,N_14540);
nand U17815 (N_17815,N_13598,N_15936);
or U17816 (N_17816,N_13719,N_15125);
nor U17817 (N_17817,N_15407,N_15347);
or U17818 (N_17818,N_15032,N_13530);
nor U17819 (N_17819,N_15179,N_13653);
and U17820 (N_17820,N_15245,N_14105);
nand U17821 (N_17821,N_12381,N_15809);
xnor U17822 (N_17822,N_14497,N_13538);
nand U17823 (N_17823,N_14697,N_14166);
xnor U17824 (N_17824,N_12159,N_14353);
and U17825 (N_17825,N_14547,N_15325);
nand U17826 (N_17826,N_14201,N_12645);
and U17827 (N_17827,N_15926,N_13764);
nand U17828 (N_17828,N_13544,N_14704);
nand U17829 (N_17829,N_13815,N_15921);
nand U17830 (N_17830,N_12967,N_12355);
or U17831 (N_17831,N_12073,N_13160);
and U17832 (N_17832,N_13518,N_12197);
nand U17833 (N_17833,N_12467,N_15784);
nor U17834 (N_17834,N_13684,N_15893);
xor U17835 (N_17835,N_12842,N_13068);
nor U17836 (N_17836,N_12710,N_15064);
nand U17837 (N_17837,N_15210,N_13197);
xnor U17838 (N_17838,N_14259,N_14521);
and U17839 (N_17839,N_14096,N_13013);
xor U17840 (N_17840,N_12399,N_14472);
or U17841 (N_17841,N_12751,N_15186);
nor U17842 (N_17842,N_12939,N_13730);
nand U17843 (N_17843,N_15898,N_12925);
or U17844 (N_17844,N_14879,N_12281);
and U17845 (N_17845,N_14203,N_15645);
and U17846 (N_17846,N_15687,N_15949);
and U17847 (N_17847,N_12511,N_15201);
nor U17848 (N_17848,N_12050,N_12140);
or U17849 (N_17849,N_15879,N_13300);
nand U17850 (N_17850,N_15197,N_15870);
and U17851 (N_17851,N_15959,N_15225);
nor U17852 (N_17852,N_15924,N_14594);
xor U17853 (N_17853,N_15517,N_12796);
and U17854 (N_17854,N_14452,N_12722);
nor U17855 (N_17855,N_13303,N_14579);
and U17856 (N_17856,N_12995,N_12323);
and U17857 (N_17857,N_12562,N_14690);
xnor U17858 (N_17858,N_14606,N_14535);
or U17859 (N_17859,N_14467,N_12326);
and U17860 (N_17860,N_14681,N_12480);
xor U17861 (N_17861,N_15055,N_13264);
xor U17862 (N_17862,N_13171,N_15847);
nand U17863 (N_17863,N_15968,N_15683);
and U17864 (N_17864,N_12120,N_13533);
xnor U17865 (N_17865,N_15840,N_12440);
and U17866 (N_17866,N_12756,N_15120);
and U17867 (N_17867,N_13818,N_13657);
nand U17868 (N_17868,N_13414,N_14313);
xor U17869 (N_17869,N_15732,N_12136);
nor U17870 (N_17870,N_14709,N_15706);
or U17871 (N_17871,N_12433,N_13392);
xnor U17872 (N_17872,N_13561,N_12272);
nand U17873 (N_17873,N_12551,N_14448);
nand U17874 (N_17874,N_12619,N_14287);
xor U17875 (N_17875,N_15365,N_14921);
nor U17876 (N_17876,N_12991,N_15409);
and U17877 (N_17877,N_12363,N_13378);
nor U17878 (N_17878,N_15331,N_14623);
nand U17879 (N_17879,N_15309,N_15590);
and U17880 (N_17880,N_14330,N_13373);
nand U17881 (N_17881,N_14519,N_13431);
xnor U17882 (N_17882,N_12772,N_15877);
or U17883 (N_17883,N_13805,N_12559);
nor U17884 (N_17884,N_13655,N_14098);
or U17885 (N_17885,N_13826,N_13144);
nor U17886 (N_17886,N_12798,N_12801);
xor U17887 (N_17887,N_12604,N_15241);
nand U17888 (N_17888,N_12611,N_12305);
and U17889 (N_17889,N_13333,N_12600);
xnor U17890 (N_17890,N_13944,N_12784);
xor U17891 (N_17891,N_12720,N_15040);
or U17892 (N_17892,N_13430,N_13862);
nor U17893 (N_17893,N_14943,N_14248);
and U17894 (N_17894,N_12593,N_13448);
nand U17895 (N_17895,N_15066,N_15751);
and U17896 (N_17896,N_14492,N_13031);
nor U17897 (N_17897,N_13893,N_13661);
or U17898 (N_17898,N_13669,N_15842);
or U17899 (N_17899,N_15572,N_12406);
nand U17900 (N_17900,N_14386,N_12125);
or U17901 (N_17901,N_13772,N_15248);
nor U17902 (N_17902,N_14707,N_13489);
and U17903 (N_17903,N_12495,N_14839);
and U17904 (N_17904,N_12429,N_12886);
and U17905 (N_17905,N_14123,N_13911);
or U17906 (N_17906,N_13383,N_13095);
nor U17907 (N_17907,N_14761,N_14696);
or U17908 (N_17908,N_13054,N_13828);
or U17909 (N_17909,N_12016,N_13804);
or U17910 (N_17910,N_12738,N_15858);
nand U17911 (N_17911,N_12962,N_15914);
and U17912 (N_17912,N_14680,N_15012);
nor U17913 (N_17913,N_12501,N_12899);
nor U17914 (N_17914,N_13577,N_15653);
or U17915 (N_17915,N_14593,N_12578);
nor U17916 (N_17916,N_15371,N_15640);
and U17917 (N_17917,N_15266,N_15765);
xnor U17918 (N_17918,N_13343,N_15771);
xnor U17919 (N_17919,N_12670,N_14181);
xnor U17920 (N_17920,N_14119,N_14135);
and U17921 (N_17921,N_13250,N_15112);
and U17922 (N_17922,N_15279,N_13960);
nand U17923 (N_17923,N_13660,N_14569);
nand U17924 (N_17924,N_15747,N_13365);
nor U17925 (N_17925,N_14362,N_14622);
or U17926 (N_17926,N_14917,N_13423);
and U17927 (N_17927,N_14446,N_14269);
or U17928 (N_17928,N_14842,N_14040);
xnor U17929 (N_17929,N_14165,N_15772);
and U17930 (N_17930,N_12813,N_13189);
or U17931 (N_17931,N_12571,N_15915);
nand U17932 (N_17932,N_12045,N_15699);
or U17933 (N_17933,N_13276,N_15498);
xnor U17934 (N_17934,N_12273,N_13915);
nor U17935 (N_17935,N_13849,N_14411);
nand U17936 (N_17936,N_14303,N_14833);
nand U17937 (N_17937,N_12966,N_14005);
nand U17938 (N_17938,N_14281,N_12033);
nor U17939 (N_17939,N_13959,N_15759);
nand U17940 (N_17940,N_12186,N_12685);
nor U17941 (N_17941,N_12314,N_13775);
and U17942 (N_17942,N_15352,N_14813);
and U17943 (N_17943,N_14959,N_14185);
or U17944 (N_17944,N_15887,N_12931);
nand U17945 (N_17945,N_15234,N_14612);
nor U17946 (N_17946,N_12181,N_15166);
and U17947 (N_17947,N_12946,N_12907);
nand U17948 (N_17948,N_14797,N_13451);
or U17949 (N_17949,N_14588,N_12827);
or U17950 (N_17950,N_15533,N_14636);
or U17951 (N_17951,N_15920,N_15556);
and U17952 (N_17952,N_13039,N_13933);
or U17953 (N_17953,N_12330,N_15389);
xnor U17954 (N_17954,N_14153,N_12208);
nor U17955 (N_17955,N_12457,N_13663);
nand U17956 (N_17956,N_12342,N_13785);
nor U17957 (N_17957,N_14395,N_12637);
nor U17958 (N_17958,N_15426,N_14738);
xnor U17959 (N_17959,N_13541,N_15049);
nand U17960 (N_17960,N_14180,N_13391);
xnor U17961 (N_17961,N_13989,N_12100);
nand U17962 (N_17962,N_12781,N_14604);
nor U17963 (N_17963,N_13808,N_14499);
and U17964 (N_17964,N_15720,N_12477);
xnor U17965 (N_17965,N_13867,N_15164);
xor U17966 (N_17966,N_13939,N_15494);
nor U17967 (N_17967,N_13462,N_12569);
nor U17968 (N_17968,N_15461,N_14661);
nor U17969 (N_17969,N_15362,N_13903);
xnor U17970 (N_17970,N_14393,N_12621);
nor U17971 (N_17971,N_12587,N_15601);
nand U17972 (N_17972,N_14637,N_12834);
and U17973 (N_17973,N_15438,N_15827);
and U17974 (N_17974,N_13640,N_15586);
xnor U17975 (N_17975,N_12447,N_12089);
nor U17976 (N_17976,N_12291,N_12576);
nor U17977 (N_17977,N_15363,N_15646);
and U17978 (N_17978,N_13223,N_13645);
and U17979 (N_17979,N_14826,N_13372);
nor U17980 (N_17980,N_14445,N_14627);
or U17981 (N_17981,N_15437,N_12299);
and U17982 (N_17982,N_14983,N_12771);
xnor U17983 (N_17983,N_12166,N_12923);
nand U17984 (N_17984,N_13823,N_12502);
and U17985 (N_17985,N_15332,N_14093);
nor U17986 (N_17986,N_12532,N_13053);
and U17987 (N_17987,N_13702,N_12385);
or U17988 (N_17988,N_12011,N_14805);
xnor U17989 (N_17989,N_12664,N_13034);
nand U17990 (N_17990,N_12663,N_12908);
nor U17991 (N_17991,N_13613,N_14173);
or U17992 (N_17992,N_14204,N_14440);
nor U17993 (N_17993,N_12404,N_12993);
and U17994 (N_17994,N_14554,N_14892);
or U17995 (N_17995,N_13620,N_13166);
and U17996 (N_17996,N_12259,N_15284);
or U17997 (N_17997,N_14325,N_14481);
and U17998 (N_17998,N_15463,N_14542);
xnor U17999 (N_17999,N_15020,N_15976);
xor U18000 (N_18000,N_15504,N_15587);
xnor U18001 (N_18001,N_13201,N_15778);
xnor U18002 (N_18002,N_12016,N_14890);
or U18003 (N_18003,N_13577,N_15250);
nand U18004 (N_18004,N_14512,N_12068);
nand U18005 (N_18005,N_14163,N_13686);
or U18006 (N_18006,N_15546,N_14898);
and U18007 (N_18007,N_15139,N_12454);
and U18008 (N_18008,N_13506,N_15184);
nand U18009 (N_18009,N_15462,N_15158);
nand U18010 (N_18010,N_12161,N_13069);
nor U18011 (N_18011,N_15678,N_14499);
nor U18012 (N_18012,N_14883,N_14955);
nand U18013 (N_18013,N_13267,N_15152);
or U18014 (N_18014,N_14641,N_15638);
and U18015 (N_18015,N_14458,N_15110);
nor U18016 (N_18016,N_12401,N_13316);
and U18017 (N_18017,N_15414,N_15539);
xnor U18018 (N_18018,N_14811,N_12919);
or U18019 (N_18019,N_12003,N_12519);
xor U18020 (N_18020,N_12984,N_12650);
and U18021 (N_18021,N_13273,N_14705);
and U18022 (N_18022,N_13051,N_15134);
and U18023 (N_18023,N_14322,N_13994);
nand U18024 (N_18024,N_14017,N_12236);
and U18025 (N_18025,N_15306,N_14320);
or U18026 (N_18026,N_14473,N_13307);
nand U18027 (N_18027,N_13712,N_12055);
nor U18028 (N_18028,N_12900,N_12916);
nand U18029 (N_18029,N_14958,N_14898);
and U18030 (N_18030,N_14566,N_14702);
or U18031 (N_18031,N_13368,N_12714);
or U18032 (N_18032,N_13580,N_14735);
nor U18033 (N_18033,N_12348,N_13068);
and U18034 (N_18034,N_12440,N_13356);
xnor U18035 (N_18035,N_14132,N_15459);
xor U18036 (N_18036,N_14419,N_12988);
nand U18037 (N_18037,N_14277,N_15552);
xor U18038 (N_18038,N_12119,N_12093);
nor U18039 (N_18039,N_13100,N_13649);
nor U18040 (N_18040,N_12120,N_13974);
or U18041 (N_18041,N_14206,N_13562);
nand U18042 (N_18042,N_14339,N_12365);
and U18043 (N_18043,N_15348,N_14460);
or U18044 (N_18044,N_13077,N_13176);
xor U18045 (N_18045,N_14704,N_12524);
nand U18046 (N_18046,N_15400,N_13350);
nand U18047 (N_18047,N_15781,N_13779);
xnor U18048 (N_18048,N_12424,N_15036);
and U18049 (N_18049,N_12358,N_14289);
nor U18050 (N_18050,N_14114,N_15434);
nand U18051 (N_18051,N_15389,N_14773);
nand U18052 (N_18052,N_12008,N_14065);
nand U18053 (N_18053,N_14359,N_15062);
or U18054 (N_18054,N_13286,N_14032);
and U18055 (N_18055,N_12286,N_15849);
nor U18056 (N_18056,N_12663,N_15445);
and U18057 (N_18057,N_14756,N_14387);
or U18058 (N_18058,N_14901,N_14229);
or U18059 (N_18059,N_13840,N_12686);
xnor U18060 (N_18060,N_13029,N_15036);
nor U18061 (N_18061,N_15578,N_12832);
or U18062 (N_18062,N_13230,N_12112);
and U18063 (N_18063,N_12763,N_15558);
xnor U18064 (N_18064,N_14076,N_14905);
nor U18065 (N_18065,N_12887,N_14841);
or U18066 (N_18066,N_13526,N_14265);
nand U18067 (N_18067,N_13174,N_14148);
or U18068 (N_18068,N_12267,N_12791);
and U18069 (N_18069,N_13533,N_12164);
or U18070 (N_18070,N_13820,N_13704);
nor U18071 (N_18071,N_13059,N_15544);
nand U18072 (N_18072,N_15110,N_13403);
and U18073 (N_18073,N_12929,N_15225);
nand U18074 (N_18074,N_13553,N_15910);
or U18075 (N_18075,N_13128,N_12965);
or U18076 (N_18076,N_14720,N_12535);
and U18077 (N_18077,N_12571,N_12233);
and U18078 (N_18078,N_12573,N_12925);
and U18079 (N_18079,N_13973,N_14064);
nor U18080 (N_18080,N_13410,N_15252);
or U18081 (N_18081,N_14211,N_15524);
xnor U18082 (N_18082,N_14180,N_12134);
nand U18083 (N_18083,N_15108,N_13339);
nand U18084 (N_18084,N_15667,N_14142);
or U18085 (N_18085,N_14802,N_14435);
nor U18086 (N_18086,N_12628,N_12255);
xor U18087 (N_18087,N_14266,N_14243);
nand U18088 (N_18088,N_12536,N_15664);
or U18089 (N_18089,N_13145,N_12188);
xor U18090 (N_18090,N_15959,N_14832);
xnor U18091 (N_18091,N_14168,N_12582);
or U18092 (N_18092,N_13123,N_13642);
nand U18093 (N_18093,N_13598,N_15055);
nand U18094 (N_18094,N_14226,N_12609);
and U18095 (N_18095,N_12603,N_13404);
nor U18096 (N_18096,N_14766,N_15664);
nand U18097 (N_18097,N_12083,N_13679);
nor U18098 (N_18098,N_14571,N_12996);
nor U18099 (N_18099,N_12353,N_12150);
xor U18100 (N_18100,N_14856,N_14405);
nor U18101 (N_18101,N_15902,N_15616);
or U18102 (N_18102,N_13013,N_13430);
nand U18103 (N_18103,N_14957,N_15032);
xor U18104 (N_18104,N_13387,N_12489);
nand U18105 (N_18105,N_14775,N_13313);
nand U18106 (N_18106,N_13549,N_15249);
or U18107 (N_18107,N_14845,N_14739);
nand U18108 (N_18108,N_13474,N_12224);
and U18109 (N_18109,N_14148,N_15108);
or U18110 (N_18110,N_14826,N_14974);
and U18111 (N_18111,N_12369,N_14488);
nand U18112 (N_18112,N_15589,N_15494);
and U18113 (N_18113,N_12320,N_14805);
xnor U18114 (N_18114,N_15237,N_13062);
xor U18115 (N_18115,N_15776,N_15511);
or U18116 (N_18116,N_15915,N_15139);
xor U18117 (N_18117,N_13195,N_13452);
nor U18118 (N_18118,N_13383,N_12835);
xor U18119 (N_18119,N_12158,N_13472);
nand U18120 (N_18120,N_13009,N_15199);
xnor U18121 (N_18121,N_12610,N_14054);
xnor U18122 (N_18122,N_13825,N_15830);
xor U18123 (N_18123,N_13599,N_15513);
and U18124 (N_18124,N_14373,N_13829);
or U18125 (N_18125,N_13341,N_13350);
nand U18126 (N_18126,N_13426,N_15291);
nor U18127 (N_18127,N_15824,N_12985);
xor U18128 (N_18128,N_14146,N_13307);
or U18129 (N_18129,N_15793,N_13346);
xnor U18130 (N_18130,N_14788,N_12278);
nand U18131 (N_18131,N_14207,N_12429);
nor U18132 (N_18132,N_15945,N_15705);
nand U18133 (N_18133,N_14394,N_13304);
xor U18134 (N_18134,N_15209,N_12876);
and U18135 (N_18135,N_12566,N_13135);
xor U18136 (N_18136,N_15033,N_12696);
or U18137 (N_18137,N_15743,N_14500);
and U18138 (N_18138,N_14633,N_12920);
and U18139 (N_18139,N_12076,N_13224);
or U18140 (N_18140,N_15495,N_15440);
nand U18141 (N_18141,N_14879,N_12098);
nand U18142 (N_18142,N_13929,N_15900);
nand U18143 (N_18143,N_12162,N_14147);
xnor U18144 (N_18144,N_13771,N_15770);
xor U18145 (N_18145,N_15582,N_15370);
or U18146 (N_18146,N_15855,N_13917);
or U18147 (N_18147,N_14071,N_15425);
nand U18148 (N_18148,N_14365,N_15401);
nor U18149 (N_18149,N_12834,N_13475);
and U18150 (N_18150,N_12192,N_13142);
nor U18151 (N_18151,N_15985,N_13055);
nand U18152 (N_18152,N_12434,N_13225);
and U18153 (N_18153,N_13259,N_13782);
and U18154 (N_18154,N_13258,N_14205);
xnor U18155 (N_18155,N_15717,N_15225);
and U18156 (N_18156,N_13922,N_15837);
and U18157 (N_18157,N_12895,N_14287);
nand U18158 (N_18158,N_15271,N_14490);
nor U18159 (N_18159,N_13916,N_15311);
and U18160 (N_18160,N_12221,N_14206);
nor U18161 (N_18161,N_14727,N_15424);
or U18162 (N_18162,N_12030,N_14358);
nand U18163 (N_18163,N_12185,N_15502);
or U18164 (N_18164,N_15733,N_14795);
and U18165 (N_18165,N_12333,N_14128);
or U18166 (N_18166,N_12535,N_15260);
xor U18167 (N_18167,N_13047,N_12678);
and U18168 (N_18168,N_12118,N_15551);
xnor U18169 (N_18169,N_14237,N_14291);
and U18170 (N_18170,N_14378,N_15374);
xnor U18171 (N_18171,N_12291,N_13679);
nand U18172 (N_18172,N_13356,N_13030);
nor U18173 (N_18173,N_15415,N_12302);
xor U18174 (N_18174,N_14005,N_14998);
and U18175 (N_18175,N_14670,N_13934);
or U18176 (N_18176,N_13959,N_13777);
and U18177 (N_18177,N_15134,N_15997);
and U18178 (N_18178,N_12584,N_14228);
nand U18179 (N_18179,N_13749,N_13773);
nand U18180 (N_18180,N_14155,N_13280);
nor U18181 (N_18181,N_14898,N_15075);
and U18182 (N_18182,N_14739,N_15346);
nand U18183 (N_18183,N_12696,N_12027);
and U18184 (N_18184,N_12165,N_15557);
or U18185 (N_18185,N_13483,N_14777);
and U18186 (N_18186,N_14033,N_13217);
or U18187 (N_18187,N_15937,N_12021);
nand U18188 (N_18188,N_14700,N_13006);
xor U18189 (N_18189,N_13917,N_13334);
nand U18190 (N_18190,N_13179,N_15498);
nor U18191 (N_18191,N_14764,N_13868);
nand U18192 (N_18192,N_13508,N_15817);
nor U18193 (N_18193,N_13691,N_12604);
nor U18194 (N_18194,N_12930,N_15845);
nand U18195 (N_18195,N_14444,N_12477);
xnor U18196 (N_18196,N_14949,N_14181);
nor U18197 (N_18197,N_13508,N_13227);
xnor U18198 (N_18198,N_15506,N_15026);
and U18199 (N_18199,N_13604,N_12390);
or U18200 (N_18200,N_14113,N_12923);
or U18201 (N_18201,N_14489,N_12342);
nand U18202 (N_18202,N_15077,N_15892);
nor U18203 (N_18203,N_13397,N_12598);
nor U18204 (N_18204,N_15571,N_12625);
xnor U18205 (N_18205,N_15444,N_15129);
nor U18206 (N_18206,N_13540,N_12868);
nand U18207 (N_18207,N_14221,N_12160);
xor U18208 (N_18208,N_14115,N_12142);
nor U18209 (N_18209,N_15252,N_15001);
or U18210 (N_18210,N_13279,N_14827);
nand U18211 (N_18211,N_14021,N_14512);
nor U18212 (N_18212,N_14991,N_15570);
and U18213 (N_18213,N_15044,N_15685);
or U18214 (N_18214,N_12171,N_13262);
nor U18215 (N_18215,N_15709,N_13994);
or U18216 (N_18216,N_15664,N_13424);
nand U18217 (N_18217,N_14728,N_12341);
nand U18218 (N_18218,N_13750,N_13156);
xnor U18219 (N_18219,N_14275,N_12917);
nand U18220 (N_18220,N_15792,N_15140);
and U18221 (N_18221,N_15317,N_14626);
or U18222 (N_18222,N_14898,N_14605);
nand U18223 (N_18223,N_13542,N_14630);
nor U18224 (N_18224,N_15438,N_15148);
xor U18225 (N_18225,N_15682,N_13357);
or U18226 (N_18226,N_15153,N_15501);
nor U18227 (N_18227,N_15282,N_15350);
nand U18228 (N_18228,N_12105,N_12952);
or U18229 (N_18229,N_15094,N_13972);
and U18230 (N_18230,N_14895,N_13454);
or U18231 (N_18231,N_12726,N_15385);
nand U18232 (N_18232,N_14110,N_13897);
xor U18233 (N_18233,N_14799,N_14215);
nor U18234 (N_18234,N_15743,N_15078);
nand U18235 (N_18235,N_13496,N_12916);
and U18236 (N_18236,N_12432,N_12939);
xor U18237 (N_18237,N_15120,N_15898);
and U18238 (N_18238,N_12075,N_13987);
and U18239 (N_18239,N_14023,N_15428);
xor U18240 (N_18240,N_13035,N_15674);
nand U18241 (N_18241,N_15233,N_15668);
nor U18242 (N_18242,N_15692,N_15344);
nand U18243 (N_18243,N_12066,N_15526);
or U18244 (N_18244,N_13841,N_15559);
and U18245 (N_18245,N_12703,N_13990);
nand U18246 (N_18246,N_14496,N_15114);
and U18247 (N_18247,N_15438,N_12900);
and U18248 (N_18248,N_15634,N_15136);
or U18249 (N_18249,N_14621,N_14731);
nor U18250 (N_18250,N_14307,N_12796);
or U18251 (N_18251,N_12301,N_14319);
xor U18252 (N_18252,N_14790,N_12901);
nand U18253 (N_18253,N_12380,N_12992);
and U18254 (N_18254,N_14362,N_12640);
nand U18255 (N_18255,N_14765,N_12889);
and U18256 (N_18256,N_14210,N_12998);
xor U18257 (N_18257,N_13803,N_15125);
and U18258 (N_18258,N_13228,N_15948);
and U18259 (N_18259,N_13177,N_14207);
xnor U18260 (N_18260,N_12869,N_14189);
nor U18261 (N_18261,N_15466,N_12904);
nor U18262 (N_18262,N_13296,N_15107);
or U18263 (N_18263,N_15519,N_12533);
or U18264 (N_18264,N_13633,N_15372);
nor U18265 (N_18265,N_15388,N_15266);
or U18266 (N_18266,N_13182,N_13611);
nand U18267 (N_18267,N_14577,N_12218);
nor U18268 (N_18268,N_14468,N_13147);
nor U18269 (N_18269,N_15947,N_15374);
nor U18270 (N_18270,N_15722,N_12518);
nand U18271 (N_18271,N_12327,N_14009);
and U18272 (N_18272,N_13691,N_13716);
nand U18273 (N_18273,N_15920,N_14647);
xnor U18274 (N_18274,N_13969,N_12799);
or U18275 (N_18275,N_15807,N_13238);
nand U18276 (N_18276,N_13667,N_12058);
or U18277 (N_18277,N_12961,N_12666);
or U18278 (N_18278,N_15481,N_13783);
xnor U18279 (N_18279,N_15421,N_13910);
xnor U18280 (N_18280,N_14901,N_13602);
xor U18281 (N_18281,N_12251,N_13891);
or U18282 (N_18282,N_13809,N_13879);
nor U18283 (N_18283,N_15808,N_15957);
or U18284 (N_18284,N_14437,N_13609);
nand U18285 (N_18285,N_15149,N_12183);
and U18286 (N_18286,N_12494,N_14447);
nand U18287 (N_18287,N_13206,N_13078);
and U18288 (N_18288,N_14942,N_12959);
xor U18289 (N_18289,N_12891,N_13682);
or U18290 (N_18290,N_14394,N_15241);
nand U18291 (N_18291,N_12282,N_15611);
nand U18292 (N_18292,N_12490,N_13768);
xnor U18293 (N_18293,N_15578,N_13260);
and U18294 (N_18294,N_14218,N_14610);
xor U18295 (N_18295,N_12018,N_12947);
xor U18296 (N_18296,N_14867,N_13672);
xnor U18297 (N_18297,N_14173,N_12242);
nor U18298 (N_18298,N_15509,N_12939);
nand U18299 (N_18299,N_13786,N_14916);
xnor U18300 (N_18300,N_14930,N_13299);
nor U18301 (N_18301,N_12041,N_14090);
and U18302 (N_18302,N_13784,N_12204);
nand U18303 (N_18303,N_12506,N_12650);
nor U18304 (N_18304,N_15101,N_14545);
nor U18305 (N_18305,N_14638,N_12588);
nor U18306 (N_18306,N_13109,N_15630);
nand U18307 (N_18307,N_14817,N_14527);
nor U18308 (N_18308,N_15626,N_14515);
nor U18309 (N_18309,N_13026,N_14288);
xor U18310 (N_18310,N_12723,N_13388);
xor U18311 (N_18311,N_14375,N_14484);
and U18312 (N_18312,N_12438,N_12687);
or U18313 (N_18313,N_14926,N_13469);
or U18314 (N_18314,N_14062,N_13637);
nand U18315 (N_18315,N_13237,N_15797);
xor U18316 (N_18316,N_15520,N_15684);
nand U18317 (N_18317,N_15378,N_14565);
nor U18318 (N_18318,N_12718,N_12283);
and U18319 (N_18319,N_12949,N_12950);
xnor U18320 (N_18320,N_13471,N_13430);
xnor U18321 (N_18321,N_15367,N_12498);
or U18322 (N_18322,N_12022,N_12660);
nor U18323 (N_18323,N_12804,N_12139);
nor U18324 (N_18324,N_15329,N_14642);
xnor U18325 (N_18325,N_12096,N_13471);
xnor U18326 (N_18326,N_12717,N_13288);
nor U18327 (N_18327,N_15474,N_12114);
and U18328 (N_18328,N_14471,N_14461);
nand U18329 (N_18329,N_12433,N_13431);
nand U18330 (N_18330,N_14694,N_15315);
or U18331 (N_18331,N_13621,N_15792);
and U18332 (N_18332,N_13338,N_15040);
and U18333 (N_18333,N_12428,N_14863);
nor U18334 (N_18334,N_13057,N_14371);
nand U18335 (N_18335,N_15424,N_12973);
and U18336 (N_18336,N_14598,N_14892);
xor U18337 (N_18337,N_12594,N_14296);
nor U18338 (N_18338,N_14925,N_12460);
or U18339 (N_18339,N_15192,N_13967);
nand U18340 (N_18340,N_12183,N_13994);
or U18341 (N_18341,N_15202,N_12633);
xor U18342 (N_18342,N_12253,N_12432);
nand U18343 (N_18343,N_12831,N_14013);
and U18344 (N_18344,N_13719,N_15982);
or U18345 (N_18345,N_15405,N_15007);
nand U18346 (N_18346,N_14763,N_13452);
and U18347 (N_18347,N_12860,N_15541);
nor U18348 (N_18348,N_13071,N_13165);
nand U18349 (N_18349,N_12986,N_14257);
or U18350 (N_18350,N_14651,N_13477);
and U18351 (N_18351,N_15955,N_14372);
nand U18352 (N_18352,N_14423,N_15319);
xor U18353 (N_18353,N_13729,N_14653);
xnor U18354 (N_18354,N_15025,N_13663);
or U18355 (N_18355,N_14971,N_13857);
and U18356 (N_18356,N_15123,N_13867);
nor U18357 (N_18357,N_15770,N_15583);
or U18358 (N_18358,N_14366,N_13006);
nand U18359 (N_18359,N_12442,N_12608);
or U18360 (N_18360,N_15656,N_12269);
or U18361 (N_18361,N_12395,N_13619);
nor U18362 (N_18362,N_13734,N_14738);
nor U18363 (N_18363,N_12693,N_13946);
nand U18364 (N_18364,N_14125,N_12415);
nand U18365 (N_18365,N_12176,N_15501);
and U18366 (N_18366,N_13175,N_15580);
or U18367 (N_18367,N_13024,N_15493);
or U18368 (N_18368,N_12514,N_14807);
or U18369 (N_18369,N_14746,N_12266);
nor U18370 (N_18370,N_14955,N_14593);
or U18371 (N_18371,N_12561,N_14591);
nor U18372 (N_18372,N_14750,N_15215);
or U18373 (N_18373,N_13063,N_13132);
xor U18374 (N_18374,N_13361,N_13178);
or U18375 (N_18375,N_13604,N_12384);
nor U18376 (N_18376,N_15448,N_15483);
and U18377 (N_18377,N_12528,N_12961);
or U18378 (N_18378,N_15455,N_15879);
and U18379 (N_18379,N_15932,N_12067);
xor U18380 (N_18380,N_14855,N_12270);
xor U18381 (N_18381,N_15109,N_14052);
nand U18382 (N_18382,N_15189,N_14168);
or U18383 (N_18383,N_12606,N_14150);
nor U18384 (N_18384,N_15205,N_14795);
nand U18385 (N_18385,N_15951,N_13724);
or U18386 (N_18386,N_15221,N_12081);
nand U18387 (N_18387,N_13525,N_12861);
nand U18388 (N_18388,N_12730,N_13491);
nor U18389 (N_18389,N_14235,N_15922);
nor U18390 (N_18390,N_12572,N_12236);
xor U18391 (N_18391,N_14490,N_14240);
or U18392 (N_18392,N_13576,N_15155);
and U18393 (N_18393,N_12276,N_13472);
or U18394 (N_18394,N_13594,N_12477);
and U18395 (N_18395,N_12731,N_14132);
and U18396 (N_18396,N_14211,N_12798);
and U18397 (N_18397,N_13524,N_12871);
or U18398 (N_18398,N_14943,N_12340);
or U18399 (N_18399,N_14287,N_13169);
nand U18400 (N_18400,N_13033,N_15419);
and U18401 (N_18401,N_12229,N_13671);
nor U18402 (N_18402,N_14027,N_15143);
nor U18403 (N_18403,N_12582,N_12956);
nor U18404 (N_18404,N_15732,N_14820);
nand U18405 (N_18405,N_14290,N_12403);
or U18406 (N_18406,N_12723,N_12242);
and U18407 (N_18407,N_15564,N_13573);
and U18408 (N_18408,N_15698,N_15436);
or U18409 (N_18409,N_13040,N_12717);
and U18410 (N_18410,N_15026,N_13226);
and U18411 (N_18411,N_13101,N_12324);
and U18412 (N_18412,N_15116,N_13436);
nand U18413 (N_18413,N_15818,N_14534);
nand U18414 (N_18414,N_15210,N_14624);
nor U18415 (N_18415,N_12075,N_12510);
nor U18416 (N_18416,N_12457,N_13887);
nand U18417 (N_18417,N_14469,N_12361);
or U18418 (N_18418,N_13549,N_13992);
nand U18419 (N_18419,N_15571,N_12158);
xor U18420 (N_18420,N_14039,N_12644);
and U18421 (N_18421,N_12058,N_12463);
nand U18422 (N_18422,N_14292,N_13421);
xnor U18423 (N_18423,N_12857,N_15261);
xor U18424 (N_18424,N_13291,N_12602);
nor U18425 (N_18425,N_14683,N_13809);
nand U18426 (N_18426,N_14945,N_12103);
or U18427 (N_18427,N_12081,N_14745);
nand U18428 (N_18428,N_12740,N_15102);
and U18429 (N_18429,N_14332,N_12620);
xor U18430 (N_18430,N_15115,N_14121);
and U18431 (N_18431,N_15858,N_13601);
nor U18432 (N_18432,N_13332,N_15237);
and U18433 (N_18433,N_15144,N_12603);
or U18434 (N_18434,N_14442,N_12862);
nor U18435 (N_18435,N_15484,N_15402);
nor U18436 (N_18436,N_15793,N_14414);
or U18437 (N_18437,N_13646,N_13162);
and U18438 (N_18438,N_13148,N_12629);
nand U18439 (N_18439,N_15565,N_14289);
or U18440 (N_18440,N_12721,N_13772);
nor U18441 (N_18441,N_12186,N_15566);
xnor U18442 (N_18442,N_12486,N_12533);
nand U18443 (N_18443,N_12813,N_14771);
xor U18444 (N_18444,N_12527,N_12285);
nor U18445 (N_18445,N_14743,N_14979);
xnor U18446 (N_18446,N_15274,N_15844);
or U18447 (N_18447,N_12647,N_14946);
and U18448 (N_18448,N_13976,N_12859);
and U18449 (N_18449,N_13807,N_15014);
or U18450 (N_18450,N_12499,N_14200);
nand U18451 (N_18451,N_13889,N_12886);
or U18452 (N_18452,N_13756,N_13394);
or U18453 (N_18453,N_12618,N_12356);
and U18454 (N_18454,N_13981,N_13517);
nor U18455 (N_18455,N_14961,N_12506);
nand U18456 (N_18456,N_13708,N_12626);
and U18457 (N_18457,N_14364,N_13923);
or U18458 (N_18458,N_15696,N_13645);
nor U18459 (N_18459,N_12416,N_12824);
xnor U18460 (N_18460,N_12780,N_14175);
or U18461 (N_18461,N_14130,N_14263);
nor U18462 (N_18462,N_15349,N_12347);
nand U18463 (N_18463,N_13125,N_14585);
or U18464 (N_18464,N_13011,N_12207);
and U18465 (N_18465,N_15173,N_14414);
or U18466 (N_18466,N_12651,N_13000);
xor U18467 (N_18467,N_13010,N_15016);
xnor U18468 (N_18468,N_14304,N_14840);
nand U18469 (N_18469,N_12200,N_13873);
and U18470 (N_18470,N_15862,N_15979);
xnor U18471 (N_18471,N_13721,N_14965);
or U18472 (N_18472,N_12041,N_13385);
and U18473 (N_18473,N_15132,N_15965);
and U18474 (N_18474,N_12867,N_14872);
and U18475 (N_18475,N_12127,N_12540);
nor U18476 (N_18476,N_15840,N_14144);
nand U18477 (N_18477,N_15271,N_13700);
xnor U18478 (N_18478,N_13468,N_12839);
nor U18479 (N_18479,N_12119,N_15830);
xor U18480 (N_18480,N_14777,N_13476);
or U18481 (N_18481,N_14888,N_15865);
xnor U18482 (N_18482,N_13416,N_14170);
nor U18483 (N_18483,N_15249,N_12800);
nor U18484 (N_18484,N_13434,N_14031);
or U18485 (N_18485,N_15583,N_13061);
or U18486 (N_18486,N_15663,N_13422);
nand U18487 (N_18487,N_13253,N_13789);
and U18488 (N_18488,N_13970,N_14848);
nand U18489 (N_18489,N_14766,N_15198);
nand U18490 (N_18490,N_15109,N_12637);
and U18491 (N_18491,N_15260,N_15042);
nor U18492 (N_18492,N_13554,N_15940);
and U18493 (N_18493,N_13935,N_12520);
or U18494 (N_18494,N_14097,N_14157);
and U18495 (N_18495,N_13111,N_12678);
xor U18496 (N_18496,N_15279,N_13235);
and U18497 (N_18497,N_12830,N_14263);
xnor U18498 (N_18498,N_13423,N_12210);
and U18499 (N_18499,N_15445,N_12322);
xnor U18500 (N_18500,N_15265,N_13451);
xor U18501 (N_18501,N_14171,N_12018);
or U18502 (N_18502,N_14404,N_14469);
or U18503 (N_18503,N_12497,N_13366);
nor U18504 (N_18504,N_12077,N_15937);
and U18505 (N_18505,N_13819,N_12073);
xor U18506 (N_18506,N_13279,N_12185);
nor U18507 (N_18507,N_15249,N_12845);
and U18508 (N_18508,N_12637,N_14476);
nand U18509 (N_18509,N_12238,N_14188);
nor U18510 (N_18510,N_15604,N_12010);
or U18511 (N_18511,N_14175,N_15259);
nand U18512 (N_18512,N_15805,N_14272);
or U18513 (N_18513,N_14667,N_14299);
nor U18514 (N_18514,N_15507,N_14930);
nor U18515 (N_18515,N_12668,N_13711);
nand U18516 (N_18516,N_15660,N_12061);
xor U18517 (N_18517,N_12889,N_14463);
xor U18518 (N_18518,N_14108,N_13856);
nor U18519 (N_18519,N_13436,N_15402);
or U18520 (N_18520,N_13370,N_15245);
xnor U18521 (N_18521,N_12495,N_14747);
and U18522 (N_18522,N_12886,N_12329);
nand U18523 (N_18523,N_12088,N_12831);
nand U18524 (N_18524,N_14434,N_14692);
nand U18525 (N_18525,N_12265,N_12529);
xor U18526 (N_18526,N_14512,N_12153);
or U18527 (N_18527,N_14867,N_15900);
nor U18528 (N_18528,N_13420,N_12647);
and U18529 (N_18529,N_14358,N_12004);
nand U18530 (N_18530,N_13255,N_13986);
nor U18531 (N_18531,N_12024,N_14596);
or U18532 (N_18532,N_14210,N_15280);
xnor U18533 (N_18533,N_13984,N_15501);
nand U18534 (N_18534,N_15409,N_13236);
or U18535 (N_18535,N_15762,N_15289);
nand U18536 (N_18536,N_15389,N_14718);
or U18537 (N_18537,N_12702,N_12727);
nand U18538 (N_18538,N_14839,N_12003);
and U18539 (N_18539,N_12047,N_13079);
nand U18540 (N_18540,N_15391,N_15996);
nor U18541 (N_18541,N_12516,N_14853);
or U18542 (N_18542,N_15316,N_15521);
xnor U18543 (N_18543,N_12214,N_15989);
nand U18544 (N_18544,N_14568,N_13849);
or U18545 (N_18545,N_15545,N_14519);
xnor U18546 (N_18546,N_13839,N_14080);
nand U18547 (N_18547,N_14270,N_14645);
or U18548 (N_18548,N_13295,N_14334);
or U18549 (N_18549,N_13504,N_13200);
nor U18550 (N_18550,N_14402,N_13957);
nand U18551 (N_18551,N_15498,N_15038);
xor U18552 (N_18552,N_12859,N_14380);
nand U18553 (N_18553,N_13137,N_12549);
nand U18554 (N_18554,N_13083,N_15952);
nand U18555 (N_18555,N_12322,N_14679);
and U18556 (N_18556,N_15117,N_13052);
or U18557 (N_18557,N_14752,N_13180);
xor U18558 (N_18558,N_12783,N_12447);
nor U18559 (N_18559,N_15814,N_12501);
nor U18560 (N_18560,N_15683,N_12903);
xnor U18561 (N_18561,N_13151,N_13951);
or U18562 (N_18562,N_14351,N_14992);
xnor U18563 (N_18563,N_14412,N_12877);
nand U18564 (N_18564,N_12589,N_12686);
xor U18565 (N_18565,N_13660,N_15896);
xnor U18566 (N_18566,N_14263,N_13793);
or U18567 (N_18567,N_12078,N_12437);
and U18568 (N_18568,N_15904,N_12902);
xor U18569 (N_18569,N_14704,N_12142);
nor U18570 (N_18570,N_15061,N_14948);
or U18571 (N_18571,N_15678,N_14221);
nand U18572 (N_18572,N_15135,N_15399);
and U18573 (N_18573,N_12674,N_14184);
and U18574 (N_18574,N_14413,N_12790);
nor U18575 (N_18575,N_15470,N_14440);
nor U18576 (N_18576,N_12202,N_14091);
xor U18577 (N_18577,N_15868,N_14124);
xor U18578 (N_18578,N_12026,N_12759);
and U18579 (N_18579,N_12139,N_13018);
nor U18580 (N_18580,N_12420,N_13854);
and U18581 (N_18581,N_13462,N_14570);
nor U18582 (N_18582,N_15454,N_12131);
xnor U18583 (N_18583,N_13212,N_13626);
or U18584 (N_18584,N_14636,N_15810);
and U18585 (N_18585,N_15801,N_14754);
and U18586 (N_18586,N_15775,N_14544);
and U18587 (N_18587,N_12748,N_14983);
or U18588 (N_18588,N_13840,N_13024);
and U18589 (N_18589,N_14476,N_13458);
or U18590 (N_18590,N_12744,N_13186);
or U18591 (N_18591,N_15058,N_13836);
xnor U18592 (N_18592,N_14007,N_15138);
nand U18593 (N_18593,N_15475,N_14881);
or U18594 (N_18594,N_13601,N_14044);
nor U18595 (N_18595,N_14419,N_12360);
nor U18596 (N_18596,N_12113,N_15379);
and U18597 (N_18597,N_13497,N_12505);
nor U18598 (N_18598,N_15733,N_12420);
xor U18599 (N_18599,N_14789,N_15386);
nand U18600 (N_18600,N_14479,N_14241);
or U18601 (N_18601,N_12249,N_14076);
xor U18602 (N_18602,N_13844,N_15103);
xnor U18603 (N_18603,N_15849,N_14614);
nand U18604 (N_18604,N_13338,N_12894);
nand U18605 (N_18605,N_15154,N_13778);
nor U18606 (N_18606,N_15478,N_15154);
nor U18607 (N_18607,N_15221,N_13498);
nand U18608 (N_18608,N_15763,N_15398);
or U18609 (N_18609,N_15923,N_12174);
nor U18610 (N_18610,N_12733,N_15194);
or U18611 (N_18611,N_14997,N_14523);
and U18612 (N_18612,N_12046,N_12056);
nor U18613 (N_18613,N_14685,N_14740);
xor U18614 (N_18614,N_13713,N_13565);
nand U18615 (N_18615,N_14692,N_12366);
and U18616 (N_18616,N_13836,N_14083);
xnor U18617 (N_18617,N_12368,N_12636);
xor U18618 (N_18618,N_12626,N_12999);
xor U18619 (N_18619,N_15292,N_13411);
and U18620 (N_18620,N_12492,N_14726);
nor U18621 (N_18621,N_14045,N_15462);
and U18622 (N_18622,N_15812,N_15705);
and U18623 (N_18623,N_15304,N_15931);
nor U18624 (N_18624,N_15922,N_13290);
and U18625 (N_18625,N_12114,N_12822);
xnor U18626 (N_18626,N_13152,N_13917);
and U18627 (N_18627,N_15072,N_14046);
nor U18628 (N_18628,N_13659,N_13746);
nor U18629 (N_18629,N_15162,N_12628);
and U18630 (N_18630,N_15981,N_15874);
nor U18631 (N_18631,N_12625,N_14145);
and U18632 (N_18632,N_12369,N_14461);
nor U18633 (N_18633,N_15098,N_12904);
xor U18634 (N_18634,N_15749,N_15754);
nand U18635 (N_18635,N_12382,N_15045);
nor U18636 (N_18636,N_13481,N_13343);
nor U18637 (N_18637,N_14147,N_13511);
or U18638 (N_18638,N_15932,N_14121);
and U18639 (N_18639,N_12790,N_14500);
or U18640 (N_18640,N_15115,N_14991);
nand U18641 (N_18641,N_12736,N_15989);
xnor U18642 (N_18642,N_15085,N_14685);
xor U18643 (N_18643,N_12272,N_13680);
nand U18644 (N_18644,N_12827,N_15293);
xnor U18645 (N_18645,N_15262,N_12415);
and U18646 (N_18646,N_14890,N_13779);
nand U18647 (N_18647,N_12161,N_14538);
nand U18648 (N_18648,N_12051,N_13949);
xnor U18649 (N_18649,N_14628,N_14011);
or U18650 (N_18650,N_12381,N_15288);
and U18651 (N_18651,N_13948,N_12045);
and U18652 (N_18652,N_12291,N_15457);
xnor U18653 (N_18653,N_13395,N_15025);
nand U18654 (N_18654,N_13605,N_15437);
or U18655 (N_18655,N_14609,N_14263);
xnor U18656 (N_18656,N_15713,N_12769);
nor U18657 (N_18657,N_12607,N_14040);
xor U18658 (N_18658,N_15967,N_14369);
nand U18659 (N_18659,N_13797,N_12820);
nor U18660 (N_18660,N_13084,N_13868);
or U18661 (N_18661,N_13136,N_15999);
xnor U18662 (N_18662,N_13769,N_13348);
xor U18663 (N_18663,N_13405,N_13936);
nor U18664 (N_18664,N_13851,N_13135);
or U18665 (N_18665,N_14569,N_13006);
nand U18666 (N_18666,N_15961,N_14112);
and U18667 (N_18667,N_15524,N_15771);
nand U18668 (N_18668,N_15357,N_12991);
or U18669 (N_18669,N_12054,N_13352);
or U18670 (N_18670,N_14360,N_12053);
xnor U18671 (N_18671,N_14883,N_12973);
xor U18672 (N_18672,N_15813,N_15969);
xnor U18673 (N_18673,N_13815,N_13249);
or U18674 (N_18674,N_14233,N_15399);
nand U18675 (N_18675,N_13333,N_14998);
nand U18676 (N_18676,N_13038,N_12118);
and U18677 (N_18677,N_13265,N_14403);
nand U18678 (N_18678,N_12658,N_14143);
nand U18679 (N_18679,N_13362,N_13420);
or U18680 (N_18680,N_15993,N_12309);
nand U18681 (N_18681,N_15707,N_15802);
or U18682 (N_18682,N_12112,N_14743);
and U18683 (N_18683,N_13558,N_13883);
xnor U18684 (N_18684,N_15397,N_15351);
or U18685 (N_18685,N_15815,N_15018);
nor U18686 (N_18686,N_15621,N_12305);
nand U18687 (N_18687,N_13943,N_12054);
nor U18688 (N_18688,N_14190,N_15236);
xnor U18689 (N_18689,N_14027,N_14803);
nand U18690 (N_18690,N_15905,N_14396);
nor U18691 (N_18691,N_15950,N_13656);
or U18692 (N_18692,N_12550,N_13963);
nand U18693 (N_18693,N_14292,N_13634);
nand U18694 (N_18694,N_13212,N_15420);
and U18695 (N_18695,N_12813,N_12971);
nand U18696 (N_18696,N_13169,N_13132);
nand U18697 (N_18697,N_13752,N_14316);
and U18698 (N_18698,N_15894,N_14975);
nor U18699 (N_18699,N_14107,N_12862);
or U18700 (N_18700,N_13816,N_12301);
nand U18701 (N_18701,N_14476,N_12925);
nand U18702 (N_18702,N_14878,N_13242);
nor U18703 (N_18703,N_12311,N_12821);
and U18704 (N_18704,N_13327,N_14257);
nor U18705 (N_18705,N_12655,N_14822);
nand U18706 (N_18706,N_13206,N_12985);
and U18707 (N_18707,N_12347,N_14001);
and U18708 (N_18708,N_14722,N_13766);
and U18709 (N_18709,N_14913,N_15098);
and U18710 (N_18710,N_15024,N_15504);
nor U18711 (N_18711,N_15532,N_12506);
or U18712 (N_18712,N_14756,N_15019);
and U18713 (N_18713,N_15315,N_13159);
nor U18714 (N_18714,N_15292,N_15845);
nor U18715 (N_18715,N_13188,N_13259);
nor U18716 (N_18716,N_15694,N_14925);
and U18717 (N_18717,N_12136,N_12869);
xnor U18718 (N_18718,N_14525,N_15093);
nand U18719 (N_18719,N_12796,N_12659);
and U18720 (N_18720,N_13439,N_12030);
nand U18721 (N_18721,N_13695,N_13119);
and U18722 (N_18722,N_12267,N_12354);
nor U18723 (N_18723,N_14759,N_13984);
or U18724 (N_18724,N_13259,N_15793);
nor U18725 (N_18725,N_13218,N_13143);
xnor U18726 (N_18726,N_15908,N_13372);
nand U18727 (N_18727,N_15397,N_15512);
and U18728 (N_18728,N_13939,N_13482);
and U18729 (N_18729,N_13966,N_12731);
or U18730 (N_18730,N_12825,N_15124);
xor U18731 (N_18731,N_12978,N_12126);
nor U18732 (N_18732,N_15871,N_12366);
nand U18733 (N_18733,N_14813,N_12470);
or U18734 (N_18734,N_13607,N_15795);
nor U18735 (N_18735,N_14258,N_12792);
and U18736 (N_18736,N_12191,N_13789);
nor U18737 (N_18737,N_12627,N_13114);
and U18738 (N_18738,N_15760,N_14430);
or U18739 (N_18739,N_13762,N_15882);
and U18740 (N_18740,N_12581,N_12685);
xnor U18741 (N_18741,N_14383,N_15431);
nand U18742 (N_18742,N_12499,N_12093);
or U18743 (N_18743,N_15770,N_14597);
or U18744 (N_18744,N_15539,N_15760);
nor U18745 (N_18745,N_12607,N_14107);
and U18746 (N_18746,N_13742,N_15600);
and U18747 (N_18747,N_15969,N_12345);
nand U18748 (N_18748,N_13037,N_14121);
or U18749 (N_18749,N_13920,N_14929);
xnor U18750 (N_18750,N_14912,N_13029);
or U18751 (N_18751,N_14551,N_12515);
nand U18752 (N_18752,N_14240,N_14374);
nor U18753 (N_18753,N_13518,N_13249);
and U18754 (N_18754,N_15510,N_13817);
nor U18755 (N_18755,N_12927,N_12557);
nor U18756 (N_18756,N_12334,N_15854);
and U18757 (N_18757,N_12085,N_12102);
nand U18758 (N_18758,N_13327,N_14200);
and U18759 (N_18759,N_13981,N_13875);
or U18760 (N_18760,N_13939,N_15995);
and U18761 (N_18761,N_15463,N_12716);
xnor U18762 (N_18762,N_12712,N_13253);
nor U18763 (N_18763,N_12636,N_12154);
or U18764 (N_18764,N_14605,N_14034);
and U18765 (N_18765,N_13778,N_15702);
nand U18766 (N_18766,N_13428,N_13415);
nor U18767 (N_18767,N_12557,N_15273);
or U18768 (N_18768,N_14964,N_15211);
nand U18769 (N_18769,N_13401,N_13357);
xnor U18770 (N_18770,N_14646,N_12782);
nor U18771 (N_18771,N_13638,N_14677);
or U18772 (N_18772,N_12335,N_12474);
xnor U18773 (N_18773,N_15227,N_15600);
and U18774 (N_18774,N_15545,N_13288);
xor U18775 (N_18775,N_14322,N_13096);
xnor U18776 (N_18776,N_13055,N_13561);
or U18777 (N_18777,N_12891,N_12549);
xnor U18778 (N_18778,N_15729,N_12124);
xor U18779 (N_18779,N_13571,N_13988);
or U18780 (N_18780,N_13655,N_13698);
nand U18781 (N_18781,N_14172,N_14190);
or U18782 (N_18782,N_13360,N_14656);
or U18783 (N_18783,N_14274,N_14768);
xnor U18784 (N_18784,N_15617,N_14543);
nor U18785 (N_18785,N_12688,N_13435);
nor U18786 (N_18786,N_12899,N_13771);
and U18787 (N_18787,N_15919,N_13101);
xnor U18788 (N_18788,N_12173,N_15051);
nand U18789 (N_18789,N_15512,N_14073);
nand U18790 (N_18790,N_13778,N_12098);
xnor U18791 (N_18791,N_14616,N_13691);
xnor U18792 (N_18792,N_12479,N_13627);
and U18793 (N_18793,N_12106,N_13368);
nand U18794 (N_18794,N_13262,N_15104);
or U18795 (N_18795,N_14916,N_14454);
nor U18796 (N_18796,N_14130,N_15518);
nand U18797 (N_18797,N_15781,N_13465);
or U18798 (N_18798,N_14605,N_12059);
nand U18799 (N_18799,N_12906,N_12129);
nor U18800 (N_18800,N_13016,N_15738);
xor U18801 (N_18801,N_13084,N_15895);
nand U18802 (N_18802,N_13585,N_13114);
nand U18803 (N_18803,N_15022,N_12995);
nand U18804 (N_18804,N_15281,N_14575);
nor U18805 (N_18805,N_12912,N_14317);
and U18806 (N_18806,N_12710,N_14872);
and U18807 (N_18807,N_15207,N_14891);
or U18808 (N_18808,N_13098,N_14468);
nor U18809 (N_18809,N_12026,N_12539);
nor U18810 (N_18810,N_12432,N_14223);
nand U18811 (N_18811,N_14833,N_12665);
nor U18812 (N_18812,N_13920,N_14707);
xor U18813 (N_18813,N_12038,N_15260);
nand U18814 (N_18814,N_15508,N_14925);
and U18815 (N_18815,N_15579,N_15424);
nor U18816 (N_18816,N_13526,N_12484);
and U18817 (N_18817,N_13366,N_13631);
xnor U18818 (N_18818,N_12587,N_13833);
xor U18819 (N_18819,N_15180,N_14423);
nand U18820 (N_18820,N_13633,N_14971);
xor U18821 (N_18821,N_13082,N_15884);
and U18822 (N_18822,N_14405,N_15467);
or U18823 (N_18823,N_12969,N_15927);
or U18824 (N_18824,N_14265,N_12074);
nor U18825 (N_18825,N_12520,N_13959);
or U18826 (N_18826,N_15385,N_13727);
or U18827 (N_18827,N_12090,N_15322);
nor U18828 (N_18828,N_14428,N_13151);
nor U18829 (N_18829,N_12515,N_15539);
nand U18830 (N_18830,N_14892,N_12046);
xnor U18831 (N_18831,N_14888,N_12417);
or U18832 (N_18832,N_15967,N_12966);
nand U18833 (N_18833,N_13547,N_15384);
nor U18834 (N_18834,N_15945,N_13856);
nand U18835 (N_18835,N_15915,N_14117);
nand U18836 (N_18836,N_12250,N_13317);
or U18837 (N_18837,N_14839,N_13233);
xor U18838 (N_18838,N_12802,N_14720);
nor U18839 (N_18839,N_12266,N_14906);
xor U18840 (N_18840,N_13028,N_13130);
and U18841 (N_18841,N_13591,N_13485);
nor U18842 (N_18842,N_13962,N_15045);
or U18843 (N_18843,N_15333,N_13556);
nor U18844 (N_18844,N_15799,N_15945);
nor U18845 (N_18845,N_15078,N_15471);
or U18846 (N_18846,N_12896,N_15741);
nor U18847 (N_18847,N_13474,N_12014);
and U18848 (N_18848,N_14957,N_13528);
and U18849 (N_18849,N_15457,N_15266);
xor U18850 (N_18850,N_13447,N_15213);
or U18851 (N_18851,N_12592,N_15201);
nand U18852 (N_18852,N_12210,N_12947);
nand U18853 (N_18853,N_12811,N_12664);
xnor U18854 (N_18854,N_14876,N_13426);
and U18855 (N_18855,N_13860,N_14599);
xor U18856 (N_18856,N_14917,N_12301);
or U18857 (N_18857,N_15322,N_15800);
or U18858 (N_18858,N_12826,N_15320);
and U18859 (N_18859,N_15554,N_13630);
nor U18860 (N_18860,N_15462,N_13682);
or U18861 (N_18861,N_15857,N_14731);
and U18862 (N_18862,N_13285,N_13836);
nor U18863 (N_18863,N_12626,N_13629);
or U18864 (N_18864,N_14051,N_13690);
and U18865 (N_18865,N_12476,N_14042);
nand U18866 (N_18866,N_13069,N_14845);
nand U18867 (N_18867,N_14706,N_12817);
and U18868 (N_18868,N_15089,N_13481);
or U18869 (N_18869,N_12572,N_13431);
or U18870 (N_18870,N_13549,N_14528);
xor U18871 (N_18871,N_14376,N_12765);
xnor U18872 (N_18872,N_15465,N_14650);
nor U18873 (N_18873,N_14832,N_13515);
xnor U18874 (N_18874,N_15900,N_15084);
xnor U18875 (N_18875,N_15165,N_15488);
nand U18876 (N_18876,N_15598,N_12925);
nor U18877 (N_18877,N_13209,N_14034);
or U18878 (N_18878,N_14168,N_15801);
nor U18879 (N_18879,N_12689,N_12998);
and U18880 (N_18880,N_13061,N_15740);
and U18881 (N_18881,N_13047,N_12935);
xnor U18882 (N_18882,N_15776,N_13351);
xor U18883 (N_18883,N_13359,N_13760);
xor U18884 (N_18884,N_13939,N_12340);
or U18885 (N_18885,N_12810,N_15785);
or U18886 (N_18886,N_15391,N_12245);
nor U18887 (N_18887,N_13239,N_12732);
nand U18888 (N_18888,N_13355,N_13730);
or U18889 (N_18889,N_12341,N_14929);
nor U18890 (N_18890,N_13739,N_15708);
xor U18891 (N_18891,N_15977,N_12964);
xnor U18892 (N_18892,N_13550,N_15115);
nand U18893 (N_18893,N_15567,N_12573);
nor U18894 (N_18894,N_14358,N_14412);
nand U18895 (N_18895,N_14614,N_12189);
and U18896 (N_18896,N_15529,N_13321);
nor U18897 (N_18897,N_15357,N_13057);
nand U18898 (N_18898,N_15197,N_13650);
nand U18899 (N_18899,N_15058,N_13759);
and U18900 (N_18900,N_14969,N_14139);
nand U18901 (N_18901,N_15649,N_12929);
nand U18902 (N_18902,N_15099,N_12107);
nor U18903 (N_18903,N_12289,N_14045);
nor U18904 (N_18904,N_15599,N_13518);
nand U18905 (N_18905,N_12282,N_13004);
and U18906 (N_18906,N_12164,N_15761);
nand U18907 (N_18907,N_15921,N_12872);
and U18908 (N_18908,N_12599,N_12027);
xnor U18909 (N_18909,N_13140,N_13709);
xor U18910 (N_18910,N_15119,N_13575);
xor U18911 (N_18911,N_14801,N_12225);
nor U18912 (N_18912,N_15396,N_12022);
and U18913 (N_18913,N_13867,N_12273);
nand U18914 (N_18914,N_12924,N_14492);
or U18915 (N_18915,N_12957,N_15610);
xnor U18916 (N_18916,N_14270,N_12908);
nor U18917 (N_18917,N_13146,N_12718);
nand U18918 (N_18918,N_14292,N_14593);
nand U18919 (N_18919,N_13401,N_13776);
nand U18920 (N_18920,N_15091,N_13233);
nand U18921 (N_18921,N_13478,N_14931);
or U18922 (N_18922,N_12991,N_14937);
xor U18923 (N_18923,N_15275,N_12619);
and U18924 (N_18924,N_13634,N_14495);
nand U18925 (N_18925,N_13575,N_14801);
and U18926 (N_18926,N_13488,N_12938);
nand U18927 (N_18927,N_13055,N_13050);
nand U18928 (N_18928,N_12194,N_14829);
and U18929 (N_18929,N_13392,N_13936);
xnor U18930 (N_18930,N_13992,N_12005);
nand U18931 (N_18931,N_12715,N_15048);
or U18932 (N_18932,N_14787,N_15344);
nand U18933 (N_18933,N_15901,N_15848);
nor U18934 (N_18934,N_14821,N_14890);
or U18935 (N_18935,N_14389,N_12143);
nor U18936 (N_18936,N_15672,N_13546);
and U18937 (N_18937,N_15368,N_14473);
and U18938 (N_18938,N_14796,N_14657);
or U18939 (N_18939,N_14731,N_15641);
and U18940 (N_18940,N_15522,N_15065);
and U18941 (N_18941,N_13662,N_14431);
nand U18942 (N_18942,N_13663,N_15934);
and U18943 (N_18943,N_13370,N_12021);
nor U18944 (N_18944,N_14746,N_15868);
or U18945 (N_18945,N_14922,N_13981);
nand U18946 (N_18946,N_14321,N_12092);
nand U18947 (N_18947,N_13156,N_15694);
and U18948 (N_18948,N_13881,N_15834);
and U18949 (N_18949,N_12783,N_15402);
and U18950 (N_18950,N_12480,N_13510);
xor U18951 (N_18951,N_14695,N_14819);
xor U18952 (N_18952,N_13937,N_14539);
or U18953 (N_18953,N_15856,N_12633);
and U18954 (N_18954,N_14553,N_12898);
and U18955 (N_18955,N_12905,N_14944);
xnor U18956 (N_18956,N_13506,N_12739);
and U18957 (N_18957,N_12936,N_15217);
and U18958 (N_18958,N_14970,N_15376);
nand U18959 (N_18959,N_14041,N_15857);
xor U18960 (N_18960,N_15892,N_13541);
nand U18961 (N_18961,N_15268,N_13792);
nand U18962 (N_18962,N_13658,N_13243);
and U18963 (N_18963,N_15785,N_12704);
nor U18964 (N_18964,N_12364,N_15598);
and U18965 (N_18965,N_13039,N_13402);
nand U18966 (N_18966,N_15429,N_15802);
nor U18967 (N_18967,N_15931,N_14410);
nand U18968 (N_18968,N_14705,N_12815);
or U18969 (N_18969,N_13122,N_12664);
and U18970 (N_18970,N_14568,N_14378);
and U18971 (N_18971,N_12868,N_12022);
and U18972 (N_18972,N_12721,N_12277);
nor U18973 (N_18973,N_14587,N_14517);
nor U18974 (N_18974,N_13230,N_15797);
nand U18975 (N_18975,N_12563,N_14135);
nand U18976 (N_18976,N_14584,N_14292);
xor U18977 (N_18977,N_12331,N_12335);
nor U18978 (N_18978,N_14334,N_13264);
nor U18979 (N_18979,N_12838,N_13608);
or U18980 (N_18980,N_15390,N_13094);
xor U18981 (N_18981,N_14121,N_14972);
xnor U18982 (N_18982,N_15077,N_15695);
xor U18983 (N_18983,N_12570,N_13420);
or U18984 (N_18984,N_14201,N_13751);
and U18985 (N_18985,N_13953,N_15440);
xnor U18986 (N_18986,N_13272,N_13754);
and U18987 (N_18987,N_15326,N_12359);
or U18988 (N_18988,N_15098,N_12645);
or U18989 (N_18989,N_15631,N_14455);
nor U18990 (N_18990,N_15881,N_14072);
xor U18991 (N_18991,N_15821,N_13786);
and U18992 (N_18992,N_14642,N_14668);
or U18993 (N_18993,N_12882,N_14139);
and U18994 (N_18994,N_13158,N_12248);
xnor U18995 (N_18995,N_14993,N_13207);
xnor U18996 (N_18996,N_13291,N_13603);
nor U18997 (N_18997,N_14222,N_14596);
nor U18998 (N_18998,N_15007,N_15195);
xnor U18999 (N_18999,N_13427,N_13061);
and U19000 (N_19000,N_13865,N_12944);
xnor U19001 (N_19001,N_12226,N_15673);
xor U19002 (N_19002,N_12819,N_12487);
and U19003 (N_19003,N_13411,N_13296);
or U19004 (N_19004,N_14310,N_14643);
nand U19005 (N_19005,N_13370,N_13942);
and U19006 (N_19006,N_13840,N_14495);
and U19007 (N_19007,N_12240,N_14171);
or U19008 (N_19008,N_12986,N_14647);
and U19009 (N_19009,N_14467,N_12769);
or U19010 (N_19010,N_13289,N_14365);
xor U19011 (N_19011,N_12617,N_15539);
nand U19012 (N_19012,N_13902,N_14717);
nand U19013 (N_19013,N_12977,N_13362);
nand U19014 (N_19014,N_12842,N_12260);
or U19015 (N_19015,N_13777,N_14753);
xnor U19016 (N_19016,N_12117,N_12635);
nand U19017 (N_19017,N_14203,N_14965);
xnor U19018 (N_19018,N_14006,N_14077);
nand U19019 (N_19019,N_12636,N_12098);
nor U19020 (N_19020,N_15031,N_12866);
nor U19021 (N_19021,N_12156,N_15213);
and U19022 (N_19022,N_12187,N_15977);
or U19023 (N_19023,N_12848,N_13727);
xor U19024 (N_19024,N_14426,N_13067);
xor U19025 (N_19025,N_14468,N_15799);
or U19026 (N_19026,N_15056,N_13659);
nand U19027 (N_19027,N_14936,N_13401);
and U19028 (N_19028,N_12267,N_15414);
or U19029 (N_19029,N_13758,N_14837);
or U19030 (N_19030,N_14981,N_15379);
nor U19031 (N_19031,N_12647,N_12845);
nand U19032 (N_19032,N_14057,N_13956);
and U19033 (N_19033,N_14009,N_12471);
or U19034 (N_19034,N_15417,N_14653);
xor U19035 (N_19035,N_14172,N_13005);
and U19036 (N_19036,N_15395,N_12808);
and U19037 (N_19037,N_15277,N_14511);
xor U19038 (N_19038,N_13598,N_15003);
or U19039 (N_19039,N_12457,N_12548);
nand U19040 (N_19040,N_14888,N_15593);
nand U19041 (N_19041,N_15021,N_13236);
nand U19042 (N_19042,N_13479,N_14366);
nand U19043 (N_19043,N_15043,N_15126);
nand U19044 (N_19044,N_14055,N_12498);
or U19045 (N_19045,N_13316,N_14637);
or U19046 (N_19046,N_14666,N_15185);
or U19047 (N_19047,N_12829,N_15595);
and U19048 (N_19048,N_14046,N_12547);
xor U19049 (N_19049,N_14920,N_12639);
nand U19050 (N_19050,N_15284,N_15757);
nor U19051 (N_19051,N_13591,N_14291);
or U19052 (N_19052,N_14387,N_12024);
nor U19053 (N_19053,N_12204,N_15968);
and U19054 (N_19054,N_15310,N_14706);
or U19055 (N_19055,N_13317,N_13217);
and U19056 (N_19056,N_14323,N_13579);
nand U19057 (N_19057,N_14456,N_14610);
or U19058 (N_19058,N_13370,N_14754);
nor U19059 (N_19059,N_13652,N_12778);
or U19060 (N_19060,N_13586,N_13900);
nor U19061 (N_19061,N_13906,N_12600);
nand U19062 (N_19062,N_12084,N_15625);
nor U19063 (N_19063,N_14950,N_15420);
nand U19064 (N_19064,N_12117,N_13164);
or U19065 (N_19065,N_12166,N_12828);
xnor U19066 (N_19066,N_14173,N_13327);
nor U19067 (N_19067,N_14472,N_14120);
nor U19068 (N_19068,N_13010,N_13879);
and U19069 (N_19069,N_14585,N_15140);
xor U19070 (N_19070,N_14656,N_12144);
nand U19071 (N_19071,N_13840,N_12350);
and U19072 (N_19072,N_13070,N_15745);
nand U19073 (N_19073,N_14079,N_13249);
and U19074 (N_19074,N_12252,N_12764);
and U19075 (N_19075,N_14066,N_14914);
nand U19076 (N_19076,N_12751,N_12670);
or U19077 (N_19077,N_13180,N_12019);
nor U19078 (N_19078,N_13260,N_15168);
nor U19079 (N_19079,N_13854,N_12533);
and U19080 (N_19080,N_13940,N_13565);
or U19081 (N_19081,N_13282,N_13919);
nor U19082 (N_19082,N_14803,N_12134);
and U19083 (N_19083,N_15982,N_15768);
nor U19084 (N_19084,N_12065,N_13993);
nand U19085 (N_19085,N_15044,N_15109);
nor U19086 (N_19086,N_12102,N_12467);
xnor U19087 (N_19087,N_15629,N_13249);
or U19088 (N_19088,N_12912,N_13506);
or U19089 (N_19089,N_14832,N_13453);
and U19090 (N_19090,N_13166,N_12745);
nand U19091 (N_19091,N_14574,N_14076);
or U19092 (N_19092,N_15228,N_13787);
nor U19093 (N_19093,N_14142,N_14111);
nand U19094 (N_19094,N_12730,N_12324);
nand U19095 (N_19095,N_15951,N_15971);
xnor U19096 (N_19096,N_14545,N_13872);
nor U19097 (N_19097,N_13161,N_15407);
nand U19098 (N_19098,N_15948,N_12067);
nand U19099 (N_19099,N_15115,N_14998);
or U19100 (N_19100,N_15572,N_15792);
nand U19101 (N_19101,N_12572,N_15044);
xor U19102 (N_19102,N_12002,N_15731);
nor U19103 (N_19103,N_15933,N_15857);
and U19104 (N_19104,N_15186,N_12274);
nand U19105 (N_19105,N_12667,N_14462);
nor U19106 (N_19106,N_15426,N_12949);
xnor U19107 (N_19107,N_15035,N_15646);
nand U19108 (N_19108,N_13941,N_15641);
or U19109 (N_19109,N_12790,N_12924);
nand U19110 (N_19110,N_15405,N_12616);
or U19111 (N_19111,N_13357,N_15232);
nand U19112 (N_19112,N_14424,N_13770);
or U19113 (N_19113,N_13511,N_15575);
nor U19114 (N_19114,N_14487,N_13691);
xnor U19115 (N_19115,N_13878,N_12882);
nor U19116 (N_19116,N_15686,N_15037);
nand U19117 (N_19117,N_14316,N_13370);
and U19118 (N_19118,N_14981,N_14478);
xor U19119 (N_19119,N_15137,N_13152);
and U19120 (N_19120,N_13713,N_15393);
or U19121 (N_19121,N_14219,N_15679);
xor U19122 (N_19122,N_13576,N_15795);
xnor U19123 (N_19123,N_15610,N_13077);
nand U19124 (N_19124,N_12424,N_13961);
and U19125 (N_19125,N_15519,N_15250);
xnor U19126 (N_19126,N_13816,N_13909);
nor U19127 (N_19127,N_15207,N_14252);
xnor U19128 (N_19128,N_15508,N_13587);
and U19129 (N_19129,N_14626,N_14302);
nand U19130 (N_19130,N_12690,N_14722);
xnor U19131 (N_19131,N_14727,N_12745);
or U19132 (N_19132,N_13666,N_15365);
xor U19133 (N_19133,N_14203,N_14543);
nand U19134 (N_19134,N_12535,N_13387);
nor U19135 (N_19135,N_14640,N_12246);
xnor U19136 (N_19136,N_12495,N_14518);
xor U19137 (N_19137,N_15256,N_13197);
or U19138 (N_19138,N_14901,N_14136);
nor U19139 (N_19139,N_15668,N_12460);
xor U19140 (N_19140,N_15624,N_12552);
and U19141 (N_19141,N_14492,N_13646);
xnor U19142 (N_19142,N_15871,N_15206);
or U19143 (N_19143,N_13424,N_13233);
and U19144 (N_19144,N_12230,N_13556);
and U19145 (N_19145,N_14790,N_12283);
or U19146 (N_19146,N_13370,N_12956);
and U19147 (N_19147,N_13710,N_12053);
or U19148 (N_19148,N_15723,N_15371);
or U19149 (N_19149,N_14695,N_13194);
xor U19150 (N_19150,N_12979,N_15212);
xnor U19151 (N_19151,N_13639,N_12278);
and U19152 (N_19152,N_15555,N_12085);
and U19153 (N_19153,N_14614,N_13108);
nand U19154 (N_19154,N_14179,N_14506);
xnor U19155 (N_19155,N_15305,N_15805);
nor U19156 (N_19156,N_15192,N_15239);
or U19157 (N_19157,N_13839,N_14986);
nor U19158 (N_19158,N_14265,N_13454);
xnor U19159 (N_19159,N_13036,N_15102);
or U19160 (N_19160,N_13825,N_14659);
xnor U19161 (N_19161,N_12121,N_14751);
nor U19162 (N_19162,N_15615,N_15329);
xor U19163 (N_19163,N_12601,N_13167);
and U19164 (N_19164,N_12339,N_14936);
nand U19165 (N_19165,N_14902,N_13185);
or U19166 (N_19166,N_12781,N_13557);
xnor U19167 (N_19167,N_15823,N_12478);
or U19168 (N_19168,N_15276,N_14814);
nand U19169 (N_19169,N_13055,N_12116);
xor U19170 (N_19170,N_14400,N_14402);
xnor U19171 (N_19171,N_14941,N_12205);
nand U19172 (N_19172,N_15547,N_13508);
xor U19173 (N_19173,N_13529,N_14926);
and U19174 (N_19174,N_15312,N_12525);
or U19175 (N_19175,N_14890,N_13340);
nand U19176 (N_19176,N_14468,N_13606);
and U19177 (N_19177,N_15235,N_12504);
and U19178 (N_19178,N_13605,N_15459);
nor U19179 (N_19179,N_15331,N_15049);
nand U19180 (N_19180,N_14731,N_13943);
xnor U19181 (N_19181,N_13373,N_15765);
nand U19182 (N_19182,N_14592,N_12163);
nand U19183 (N_19183,N_13644,N_12945);
nand U19184 (N_19184,N_15848,N_14564);
nand U19185 (N_19185,N_15165,N_12729);
nand U19186 (N_19186,N_15719,N_15346);
nand U19187 (N_19187,N_15030,N_13794);
xor U19188 (N_19188,N_12992,N_15431);
or U19189 (N_19189,N_14314,N_13754);
or U19190 (N_19190,N_12257,N_12912);
and U19191 (N_19191,N_12547,N_13887);
and U19192 (N_19192,N_14169,N_13264);
nand U19193 (N_19193,N_14471,N_12366);
nand U19194 (N_19194,N_13486,N_13972);
xnor U19195 (N_19195,N_12962,N_15840);
nand U19196 (N_19196,N_13549,N_13628);
xor U19197 (N_19197,N_13372,N_13181);
and U19198 (N_19198,N_13965,N_13021);
or U19199 (N_19199,N_15686,N_13361);
xor U19200 (N_19200,N_14403,N_13623);
and U19201 (N_19201,N_13748,N_12707);
nand U19202 (N_19202,N_12549,N_12405);
nand U19203 (N_19203,N_13613,N_12782);
nor U19204 (N_19204,N_12636,N_12628);
xor U19205 (N_19205,N_14332,N_15453);
xnor U19206 (N_19206,N_13173,N_13192);
nand U19207 (N_19207,N_15834,N_15703);
nand U19208 (N_19208,N_14774,N_14681);
nor U19209 (N_19209,N_14111,N_12312);
nor U19210 (N_19210,N_12324,N_15686);
nor U19211 (N_19211,N_15931,N_13376);
or U19212 (N_19212,N_13575,N_14152);
and U19213 (N_19213,N_15492,N_14337);
and U19214 (N_19214,N_15280,N_14940);
nor U19215 (N_19215,N_13678,N_13431);
nor U19216 (N_19216,N_15617,N_12497);
xor U19217 (N_19217,N_13791,N_13101);
nor U19218 (N_19218,N_14147,N_15691);
nor U19219 (N_19219,N_12949,N_12181);
or U19220 (N_19220,N_13981,N_15303);
or U19221 (N_19221,N_14644,N_15472);
xor U19222 (N_19222,N_13406,N_12495);
and U19223 (N_19223,N_13541,N_14507);
nand U19224 (N_19224,N_13770,N_13816);
xnor U19225 (N_19225,N_13704,N_12809);
nand U19226 (N_19226,N_14819,N_13466);
or U19227 (N_19227,N_14246,N_15468);
and U19228 (N_19228,N_12306,N_14815);
and U19229 (N_19229,N_15933,N_14194);
nor U19230 (N_19230,N_15953,N_15302);
and U19231 (N_19231,N_15511,N_14683);
and U19232 (N_19232,N_12569,N_12940);
and U19233 (N_19233,N_13657,N_13724);
xnor U19234 (N_19234,N_12141,N_15668);
xnor U19235 (N_19235,N_15089,N_14640);
nor U19236 (N_19236,N_13983,N_14320);
nand U19237 (N_19237,N_12886,N_14128);
xnor U19238 (N_19238,N_14128,N_12252);
and U19239 (N_19239,N_13520,N_14339);
xor U19240 (N_19240,N_15425,N_13503);
or U19241 (N_19241,N_12580,N_12073);
or U19242 (N_19242,N_13404,N_12323);
nor U19243 (N_19243,N_13534,N_15243);
xor U19244 (N_19244,N_12485,N_14183);
xor U19245 (N_19245,N_13201,N_14751);
or U19246 (N_19246,N_12256,N_12679);
nand U19247 (N_19247,N_13081,N_12582);
nand U19248 (N_19248,N_14058,N_15996);
and U19249 (N_19249,N_14754,N_13861);
or U19250 (N_19250,N_13903,N_12980);
or U19251 (N_19251,N_15690,N_14375);
nand U19252 (N_19252,N_13442,N_14637);
nand U19253 (N_19253,N_15691,N_15560);
nand U19254 (N_19254,N_15554,N_13281);
and U19255 (N_19255,N_15347,N_15210);
xor U19256 (N_19256,N_15352,N_15787);
nor U19257 (N_19257,N_13495,N_13633);
and U19258 (N_19258,N_12087,N_13303);
xnor U19259 (N_19259,N_15965,N_12249);
or U19260 (N_19260,N_14448,N_13109);
nand U19261 (N_19261,N_15599,N_15520);
nor U19262 (N_19262,N_13343,N_12102);
nor U19263 (N_19263,N_13484,N_15017);
xnor U19264 (N_19264,N_15042,N_13574);
or U19265 (N_19265,N_12897,N_13584);
nand U19266 (N_19266,N_15352,N_12740);
or U19267 (N_19267,N_14533,N_14154);
and U19268 (N_19268,N_13651,N_12233);
xor U19269 (N_19269,N_13006,N_12053);
nand U19270 (N_19270,N_15591,N_13787);
or U19271 (N_19271,N_13705,N_12154);
or U19272 (N_19272,N_13420,N_14769);
xor U19273 (N_19273,N_15410,N_13815);
and U19274 (N_19274,N_12799,N_13834);
or U19275 (N_19275,N_14072,N_14531);
and U19276 (N_19276,N_13213,N_14423);
and U19277 (N_19277,N_13005,N_14720);
nand U19278 (N_19278,N_12145,N_13834);
xor U19279 (N_19279,N_14529,N_13438);
xor U19280 (N_19280,N_14714,N_12077);
nor U19281 (N_19281,N_14164,N_14599);
and U19282 (N_19282,N_13568,N_13243);
nand U19283 (N_19283,N_14490,N_15330);
and U19284 (N_19284,N_13294,N_15477);
or U19285 (N_19285,N_13226,N_14928);
xor U19286 (N_19286,N_12167,N_13528);
and U19287 (N_19287,N_15011,N_14156);
and U19288 (N_19288,N_15923,N_12636);
nand U19289 (N_19289,N_14268,N_14091);
or U19290 (N_19290,N_15444,N_15569);
nor U19291 (N_19291,N_12598,N_13577);
or U19292 (N_19292,N_14035,N_13426);
or U19293 (N_19293,N_15580,N_15522);
nand U19294 (N_19294,N_12829,N_13621);
nand U19295 (N_19295,N_12693,N_15086);
xor U19296 (N_19296,N_14316,N_15907);
nor U19297 (N_19297,N_13460,N_13380);
or U19298 (N_19298,N_15100,N_15378);
nand U19299 (N_19299,N_14091,N_14005);
nor U19300 (N_19300,N_14446,N_15939);
nor U19301 (N_19301,N_14949,N_15694);
and U19302 (N_19302,N_12368,N_13177);
nand U19303 (N_19303,N_15548,N_14357);
nand U19304 (N_19304,N_15000,N_12261);
xor U19305 (N_19305,N_13670,N_13725);
xnor U19306 (N_19306,N_13972,N_15882);
and U19307 (N_19307,N_15999,N_14894);
xnor U19308 (N_19308,N_12064,N_13991);
nor U19309 (N_19309,N_15776,N_12404);
and U19310 (N_19310,N_15859,N_14150);
xnor U19311 (N_19311,N_15860,N_13550);
nor U19312 (N_19312,N_13870,N_15920);
or U19313 (N_19313,N_13660,N_14202);
nand U19314 (N_19314,N_15706,N_13921);
or U19315 (N_19315,N_13606,N_15529);
xor U19316 (N_19316,N_15639,N_12001);
nand U19317 (N_19317,N_12620,N_12017);
or U19318 (N_19318,N_13537,N_14335);
nand U19319 (N_19319,N_12894,N_14639);
nand U19320 (N_19320,N_15021,N_14762);
xor U19321 (N_19321,N_15802,N_13040);
and U19322 (N_19322,N_15112,N_14729);
xnor U19323 (N_19323,N_15652,N_13231);
nand U19324 (N_19324,N_12990,N_12810);
and U19325 (N_19325,N_13741,N_12672);
nor U19326 (N_19326,N_12396,N_15646);
nor U19327 (N_19327,N_15352,N_14717);
xor U19328 (N_19328,N_14447,N_14514);
xor U19329 (N_19329,N_14731,N_14103);
nand U19330 (N_19330,N_15752,N_12224);
nor U19331 (N_19331,N_15104,N_15776);
nand U19332 (N_19332,N_15966,N_12277);
nor U19333 (N_19333,N_12467,N_13462);
and U19334 (N_19334,N_14990,N_12781);
nor U19335 (N_19335,N_12279,N_12733);
xnor U19336 (N_19336,N_13143,N_14328);
nor U19337 (N_19337,N_13303,N_12090);
and U19338 (N_19338,N_14888,N_13638);
and U19339 (N_19339,N_14107,N_12079);
or U19340 (N_19340,N_12717,N_14136);
xnor U19341 (N_19341,N_15324,N_12194);
nor U19342 (N_19342,N_15390,N_14278);
nor U19343 (N_19343,N_15266,N_13918);
or U19344 (N_19344,N_12369,N_15147);
nor U19345 (N_19345,N_14153,N_14240);
nor U19346 (N_19346,N_12389,N_14100);
nor U19347 (N_19347,N_15316,N_14565);
nand U19348 (N_19348,N_15605,N_15297);
and U19349 (N_19349,N_13379,N_15428);
xor U19350 (N_19350,N_14475,N_14655);
nor U19351 (N_19351,N_15026,N_13534);
nor U19352 (N_19352,N_12352,N_13950);
or U19353 (N_19353,N_15568,N_12014);
nand U19354 (N_19354,N_14551,N_12520);
xnor U19355 (N_19355,N_12906,N_15690);
and U19356 (N_19356,N_13689,N_12548);
nor U19357 (N_19357,N_14923,N_14910);
or U19358 (N_19358,N_13776,N_14678);
xor U19359 (N_19359,N_13285,N_15034);
xor U19360 (N_19360,N_15902,N_15325);
nor U19361 (N_19361,N_15422,N_14804);
xnor U19362 (N_19362,N_12215,N_14854);
nor U19363 (N_19363,N_15508,N_15229);
nand U19364 (N_19364,N_13466,N_15547);
xnor U19365 (N_19365,N_12037,N_12529);
and U19366 (N_19366,N_13634,N_15488);
or U19367 (N_19367,N_15212,N_12996);
or U19368 (N_19368,N_14248,N_13402);
xor U19369 (N_19369,N_13550,N_12675);
xor U19370 (N_19370,N_15392,N_12603);
or U19371 (N_19371,N_15154,N_13929);
or U19372 (N_19372,N_14557,N_14429);
and U19373 (N_19373,N_15147,N_12701);
or U19374 (N_19374,N_15488,N_15620);
or U19375 (N_19375,N_12012,N_14351);
or U19376 (N_19376,N_13871,N_12270);
or U19377 (N_19377,N_13469,N_15420);
nand U19378 (N_19378,N_15535,N_14141);
xor U19379 (N_19379,N_12370,N_13138);
or U19380 (N_19380,N_15630,N_12150);
and U19381 (N_19381,N_12931,N_15472);
xnor U19382 (N_19382,N_12410,N_13930);
nor U19383 (N_19383,N_13524,N_14469);
or U19384 (N_19384,N_14419,N_13347);
nand U19385 (N_19385,N_14817,N_12480);
and U19386 (N_19386,N_12379,N_15084);
or U19387 (N_19387,N_13491,N_14921);
nand U19388 (N_19388,N_13396,N_15923);
xnor U19389 (N_19389,N_13500,N_13231);
or U19390 (N_19390,N_14537,N_12592);
and U19391 (N_19391,N_15723,N_14583);
and U19392 (N_19392,N_15859,N_13926);
and U19393 (N_19393,N_15509,N_15785);
or U19394 (N_19394,N_12411,N_12496);
or U19395 (N_19395,N_13043,N_14144);
xor U19396 (N_19396,N_13006,N_12339);
and U19397 (N_19397,N_13158,N_14616);
xor U19398 (N_19398,N_13965,N_12916);
or U19399 (N_19399,N_14165,N_12261);
nor U19400 (N_19400,N_12523,N_13484);
nand U19401 (N_19401,N_12927,N_13013);
nor U19402 (N_19402,N_12988,N_13584);
xnor U19403 (N_19403,N_13970,N_12036);
xor U19404 (N_19404,N_13716,N_12105);
xor U19405 (N_19405,N_13564,N_14755);
or U19406 (N_19406,N_12142,N_12339);
xnor U19407 (N_19407,N_12860,N_12552);
nand U19408 (N_19408,N_14659,N_13152);
and U19409 (N_19409,N_14477,N_12440);
or U19410 (N_19410,N_14036,N_13600);
or U19411 (N_19411,N_13906,N_13595);
nand U19412 (N_19412,N_14316,N_12575);
nand U19413 (N_19413,N_12493,N_13819);
nor U19414 (N_19414,N_13461,N_14770);
and U19415 (N_19415,N_13909,N_12828);
nor U19416 (N_19416,N_15867,N_13138);
xor U19417 (N_19417,N_12508,N_12520);
xnor U19418 (N_19418,N_12075,N_14441);
nand U19419 (N_19419,N_15352,N_13381);
or U19420 (N_19420,N_13518,N_12859);
and U19421 (N_19421,N_12643,N_12911);
nor U19422 (N_19422,N_15688,N_14168);
and U19423 (N_19423,N_14228,N_14255);
xor U19424 (N_19424,N_13443,N_14094);
nand U19425 (N_19425,N_14971,N_14890);
nor U19426 (N_19426,N_13307,N_13340);
or U19427 (N_19427,N_13982,N_14394);
nand U19428 (N_19428,N_14501,N_14727);
nor U19429 (N_19429,N_13849,N_12366);
xnor U19430 (N_19430,N_14013,N_13762);
and U19431 (N_19431,N_15978,N_12938);
or U19432 (N_19432,N_13295,N_15178);
and U19433 (N_19433,N_13154,N_12531);
or U19434 (N_19434,N_15334,N_12842);
xor U19435 (N_19435,N_12574,N_12084);
nand U19436 (N_19436,N_13156,N_12906);
xor U19437 (N_19437,N_12862,N_14739);
nor U19438 (N_19438,N_13276,N_15934);
xnor U19439 (N_19439,N_15460,N_14000);
xnor U19440 (N_19440,N_14952,N_15845);
nand U19441 (N_19441,N_14940,N_15059);
xnor U19442 (N_19442,N_12349,N_13058);
nor U19443 (N_19443,N_12195,N_14355);
xnor U19444 (N_19444,N_14239,N_15733);
and U19445 (N_19445,N_15934,N_14014);
nand U19446 (N_19446,N_14259,N_12741);
nor U19447 (N_19447,N_15004,N_15197);
xnor U19448 (N_19448,N_14861,N_15500);
and U19449 (N_19449,N_15122,N_14649);
and U19450 (N_19450,N_14308,N_15442);
or U19451 (N_19451,N_15010,N_14589);
and U19452 (N_19452,N_12742,N_15667);
nand U19453 (N_19453,N_12204,N_15196);
nand U19454 (N_19454,N_15231,N_14978);
xor U19455 (N_19455,N_15661,N_14830);
nor U19456 (N_19456,N_14619,N_12085);
or U19457 (N_19457,N_14647,N_13497);
xnor U19458 (N_19458,N_15307,N_13898);
or U19459 (N_19459,N_12589,N_13790);
nor U19460 (N_19460,N_14151,N_14115);
or U19461 (N_19461,N_15231,N_14634);
nor U19462 (N_19462,N_15937,N_13966);
or U19463 (N_19463,N_14252,N_12962);
or U19464 (N_19464,N_13100,N_14698);
or U19465 (N_19465,N_15756,N_13224);
xnor U19466 (N_19466,N_12298,N_14124);
xnor U19467 (N_19467,N_15461,N_12556);
nor U19468 (N_19468,N_13413,N_15116);
or U19469 (N_19469,N_12771,N_13873);
nor U19470 (N_19470,N_14675,N_14600);
or U19471 (N_19471,N_15221,N_12995);
or U19472 (N_19472,N_13483,N_13739);
nand U19473 (N_19473,N_13078,N_14303);
nor U19474 (N_19474,N_12492,N_13681);
xor U19475 (N_19475,N_14144,N_15796);
nor U19476 (N_19476,N_12656,N_12103);
nor U19477 (N_19477,N_14318,N_14305);
or U19478 (N_19478,N_12952,N_15079);
nor U19479 (N_19479,N_12263,N_13417);
nor U19480 (N_19480,N_13113,N_13212);
nor U19481 (N_19481,N_13011,N_12475);
xnor U19482 (N_19482,N_14275,N_12973);
or U19483 (N_19483,N_14012,N_12759);
xor U19484 (N_19484,N_15222,N_15053);
xor U19485 (N_19485,N_14833,N_13555);
or U19486 (N_19486,N_13564,N_14260);
and U19487 (N_19487,N_13269,N_14182);
or U19488 (N_19488,N_12824,N_15220);
nor U19489 (N_19489,N_12285,N_13816);
and U19490 (N_19490,N_13401,N_14505);
or U19491 (N_19491,N_14569,N_12170);
nor U19492 (N_19492,N_14531,N_15684);
and U19493 (N_19493,N_13012,N_15406);
xnor U19494 (N_19494,N_14565,N_14098);
or U19495 (N_19495,N_14819,N_15190);
or U19496 (N_19496,N_13257,N_13955);
nor U19497 (N_19497,N_12591,N_15302);
or U19498 (N_19498,N_15290,N_12338);
nand U19499 (N_19499,N_14716,N_13291);
xor U19500 (N_19500,N_15535,N_14810);
or U19501 (N_19501,N_14581,N_14073);
xor U19502 (N_19502,N_12688,N_12624);
nand U19503 (N_19503,N_12433,N_15844);
nor U19504 (N_19504,N_13144,N_14627);
xnor U19505 (N_19505,N_13275,N_13650);
and U19506 (N_19506,N_14176,N_14647);
nor U19507 (N_19507,N_12518,N_14207);
or U19508 (N_19508,N_14506,N_13639);
and U19509 (N_19509,N_14773,N_13207);
nor U19510 (N_19510,N_13719,N_13533);
nor U19511 (N_19511,N_12089,N_14405);
and U19512 (N_19512,N_13194,N_15483);
nand U19513 (N_19513,N_12985,N_15247);
and U19514 (N_19514,N_14184,N_12508);
xnor U19515 (N_19515,N_12605,N_12489);
nor U19516 (N_19516,N_14972,N_14966);
xor U19517 (N_19517,N_15019,N_15974);
and U19518 (N_19518,N_13079,N_14262);
xnor U19519 (N_19519,N_14606,N_15184);
xor U19520 (N_19520,N_13012,N_13435);
nand U19521 (N_19521,N_13567,N_12297);
nor U19522 (N_19522,N_12828,N_12450);
nor U19523 (N_19523,N_14804,N_12535);
or U19524 (N_19524,N_15098,N_14837);
nand U19525 (N_19525,N_12190,N_15669);
nor U19526 (N_19526,N_13923,N_13513);
and U19527 (N_19527,N_13460,N_15555);
nor U19528 (N_19528,N_13042,N_15959);
and U19529 (N_19529,N_15677,N_15944);
xnor U19530 (N_19530,N_15673,N_15347);
nand U19531 (N_19531,N_14171,N_15212);
and U19532 (N_19532,N_15222,N_14296);
xnor U19533 (N_19533,N_15333,N_14850);
or U19534 (N_19534,N_13411,N_15426);
and U19535 (N_19535,N_14040,N_15199);
nand U19536 (N_19536,N_15134,N_14744);
and U19537 (N_19537,N_13797,N_14843);
and U19538 (N_19538,N_12966,N_13277);
and U19539 (N_19539,N_12126,N_13198);
nor U19540 (N_19540,N_14924,N_12063);
nand U19541 (N_19541,N_13281,N_15454);
and U19542 (N_19542,N_14622,N_12819);
or U19543 (N_19543,N_15187,N_12029);
nor U19544 (N_19544,N_12209,N_14166);
and U19545 (N_19545,N_14738,N_12432);
and U19546 (N_19546,N_13919,N_12310);
or U19547 (N_19547,N_12518,N_12849);
and U19548 (N_19548,N_13972,N_12927);
or U19549 (N_19549,N_12851,N_14097);
and U19550 (N_19550,N_15597,N_12648);
nand U19551 (N_19551,N_15731,N_13050);
nor U19552 (N_19552,N_13974,N_13643);
xor U19553 (N_19553,N_14621,N_14150);
and U19554 (N_19554,N_15898,N_14126);
nor U19555 (N_19555,N_13519,N_15233);
and U19556 (N_19556,N_13703,N_15193);
nor U19557 (N_19557,N_14510,N_13599);
and U19558 (N_19558,N_15874,N_12272);
or U19559 (N_19559,N_15915,N_14172);
xnor U19560 (N_19560,N_14207,N_13007);
and U19561 (N_19561,N_14167,N_12948);
nor U19562 (N_19562,N_14120,N_12208);
or U19563 (N_19563,N_12338,N_14938);
or U19564 (N_19564,N_15632,N_13011);
or U19565 (N_19565,N_15138,N_15487);
nand U19566 (N_19566,N_13004,N_13681);
nor U19567 (N_19567,N_12033,N_15123);
nand U19568 (N_19568,N_14835,N_15057);
nand U19569 (N_19569,N_12327,N_13774);
and U19570 (N_19570,N_15219,N_12305);
and U19571 (N_19571,N_13191,N_15363);
nor U19572 (N_19572,N_12040,N_14434);
and U19573 (N_19573,N_12395,N_12834);
or U19574 (N_19574,N_12843,N_13974);
nor U19575 (N_19575,N_14908,N_14478);
nor U19576 (N_19576,N_12100,N_12856);
xor U19577 (N_19577,N_13813,N_15691);
and U19578 (N_19578,N_13583,N_14569);
nand U19579 (N_19579,N_13991,N_14640);
or U19580 (N_19580,N_15767,N_14614);
or U19581 (N_19581,N_14508,N_14056);
nand U19582 (N_19582,N_13611,N_15219);
or U19583 (N_19583,N_15113,N_13484);
or U19584 (N_19584,N_14335,N_14903);
nor U19585 (N_19585,N_13843,N_14554);
or U19586 (N_19586,N_12784,N_13261);
or U19587 (N_19587,N_13125,N_13957);
and U19588 (N_19588,N_15264,N_15941);
and U19589 (N_19589,N_12112,N_14792);
and U19590 (N_19590,N_15515,N_12940);
xor U19591 (N_19591,N_13009,N_15925);
and U19592 (N_19592,N_14707,N_12963);
nor U19593 (N_19593,N_15142,N_14639);
or U19594 (N_19594,N_14714,N_15900);
nand U19595 (N_19595,N_12931,N_14341);
nand U19596 (N_19596,N_14271,N_15749);
and U19597 (N_19597,N_13543,N_13029);
nor U19598 (N_19598,N_13641,N_13007);
nand U19599 (N_19599,N_15381,N_12612);
and U19600 (N_19600,N_15509,N_13984);
xor U19601 (N_19601,N_14739,N_13357);
or U19602 (N_19602,N_13622,N_15201);
nand U19603 (N_19603,N_15692,N_15223);
nand U19604 (N_19604,N_15822,N_13795);
and U19605 (N_19605,N_14283,N_15829);
xnor U19606 (N_19606,N_15945,N_12700);
or U19607 (N_19607,N_14656,N_13933);
xnor U19608 (N_19608,N_15809,N_13456);
nand U19609 (N_19609,N_14823,N_14625);
nor U19610 (N_19610,N_14361,N_12969);
nor U19611 (N_19611,N_12986,N_12486);
xnor U19612 (N_19612,N_12488,N_12890);
nor U19613 (N_19613,N_15645,N_15749);
xnor U19614 (N_19614,N_14944,N_15186);
nand U19615 (N_19615,N_13425,N_14984);
and U19616 (N_19616,N_14351,N_13311);
nor U19617 (N_19617,N_12024,N_14284);
xnor U19618 (N_19618,N_14376,N_15460);
nand U19619 (N_19619,N_13111,N_14900);
nand U19620 (N_19620,N_14630,N_12368);
nand U19621 (N_19621,N_15856,N_15593);
xor U19622 (N_19622,N_14076,N_12894);
or U19623 (N_19623,N_15821,N_12621);
and U19624 (N_19624,N_13452,N_12832);
nand U19625 (N_19625,N_13895,N_14026);
nor U19626 (N_19626,N_13289,N_14494);
nor U19627 (N_19627,N_12288,N_12372);
and U19628 (N_19628,N_12748,N_15308);
nor U19629 (N_19629,N_15375,N_15143);
or U19630 (N_19630,N_14651,N_12388);
nor U19631 (N_19631,N_15021,N_14050);
and U19632 (N_19632,N_13081,N_15236);
nand U19633 (N_19633,N_14388,N_13554);
or U19634 (N_19634,N_15819,N_12431);
xnor U19635 (N_19635,N_13838,N_15960);
nand U19636 (N_19636,N_15886,N_13470);
and U19637 (N_19637,N_14645,N_14224);
nand U19638 (N_19638,N_14525,N_14512);
xor U19639 (N_19639,N_14430,N_14750);
or U19640 (N_19640,N_13933,N_12363);
and U19641 (N_19641,N_14462,N_14456);
and U19642 (N_19642,N_15485,N_12474);
and U19643 (N_19643,N_13691,N_15847);
nor U19644 (N_19644,N_15251,N_15394);
nand U19645 (N_19645,N_12278,N_12730);
nor U19646 (N_19646,N_15572,N_15026);
or U19647 (N_19647,N_15526,N_12590);
xor U19648 (N_19648,N_13604,N_15542);
or U19649 (N_19649,N_14866,N_14587);
and U19650 (N_19650,N_15284,N_15733);
or U19651 (N_19651,N_12051,N_13926);
nand U19652 (N_19652,N_14986,N_15321);
nor U19653 (N_19653,N_13119,N_15343);
nand U19654 (N_19654,N_15347,N_14004);
nor U19655 (N_19655,N_13778,N_14993);
and U19656 (N_19656,N_14205,N_13352);
or U19657 (N_19657,N_14365,N_14790);
nor U19658 (N_19658,N_13025,N_12127);
nor U19659 (N_19659,N_13720,N_13944);
and U19660 (N_19660,N_15993,N_13028);
nor U19661 (N_19661,N_12146,N_12872);
or U19662 (N_19662,N_14552,N_12076);
xor U19663 (N_19663,N_14896,N_12601);
nand U19664 (N_19664,N_12502,N_15128);
and U19665 (N_19665,N_14843,N_14331);
xnor U19666 (N_19666,N_12848,N_15364);
xnor U19667 (N_19667,N_13430,N_14628);
xnor U19668 (N_19668,N_15439,N_14611);
xnor U19669 (N_19669,N_12207,N_15187);
or U19670 (N_19670,N_12667,N_13880);
xnor U19671 (N_19671,N_15431,N_13028);
nand U19672 (N_19672,N_14291,N_14517);
xnor U19673 (N_19673,N_15317,N_15631);
and U19674 (N_19674,N_15919,N_14721);
nand U19675 (N_19675,N_15510,N_12147);
nand U19676 (N_19676,N_14116,N_12594);
or U19677 (N_19677,N_14979,N_12569);
and U19678 (N_19678,N_12095,N_12777);
nand U19679 (N_19679,N_12051,N_12315);
and U19680 (N_19680,N_13852,N_12328);
nor U19681 (N_19681,N_12955,N_12051);
nand U19682 (N_19682,N_13875,N_14707);
nor U19683 (N_19683,N_12046,N_14037);
nand U19684 (N_19684,N_12826,N_12171);
or U19685 (N_19685,N_15607,N_12372);
xor U19686 (N_19686,N_15274,N_14536);
xnor U19687 (N_19687,N_15061,N_13596);
nand U19688 (N_19688,N_15016,N_13576);
or U19689 (N_19689,N_13139,N_15174);
or U19690 (N_19690,N_15244,N_14644);
and U19691 (N_19691,N_15685,N_14013);
nor U19692 (N_19692,N_15929,N_12172);
nor U19693 (N_19693,N_15168,N_13166);
or U19694 (N_19694,N_13433,N_12598);
nand U19695 (N_19695,N_15941,N_13040);
and U19696 (N_19696,N_15296,N_15513);
xnor U19697 (N_19697,N_14700,N_14825);
xnor U19698 (N_19698,N_14655,N_15925);
and U19699 (N_19699,N_12878,N_13498);
xor U19700 (N_19700,N_15147,N_14268);
or U19701 (N_19701,N_13784,N_14872);
nand U19702 (N_19702,N_14509,N_15083);
nand U19703 (N_19703,N_13382,N_15915);
xor U19704 (N_19704,N_12529,N_14735);
or U19705 (N_19705,N_13844,N_15627);
and U19706 (N_19706,N_12007,N_15003);
xnor U19707 (N_19707,N_12540,N_14174);
or U19708 (N_19708,N_13040,N_15657);
and U19709 (N_19709,N_12937,N_15313);
and U19710 (N_19710,N_14877,N_13879);
nor U19711 (N_19711,N_13078,N_14885);
and U19712 (N_19712,N_12463,N_15468);
and U19713 (N_19713,N_15271,N_14095);
or U19714 (N_19714,N_15038,N_15866);
nand U19715 (N_19715,N_15173,N_14212);
xor U19716 (N_19716,N_15355,N_14885);
nor U19717 (N_19717,N_12305,N_15542);
xnor U19718 (N_19718,N_15665,N_14976);
nor U19719 (N_19719,N_14619,N_15849);
xnor U19720 (N_19720,N_14993,N_15984);
nand U19721 (N_19721,N_14821,N_13893);
and U19722 (N_19722,N_14469,N_15961);
nor U19723 (N_19723,N_14818,N_14070);
nor U19724 (N_19724,N_13052,N_15501);
nor U19725 (N_19725,N_15053,N_14149);
xnor U19726 (N_19726,N_14121,N_13889);
xnor U19727 (N_19727,N_14674,N_13226);
or U19728 (N_19728,N_15346,N_15294);
and U19729 (N_19729,N_13489,N_15146);
and U19730 (N_19730,N_15466,N_15709);
xnor U19731 (N_19731,N_12255,N_13548);
or U19732 (N_19732,N_13924,N_12030);
nor U19733 (N_19733,N_15624,N_14995);
or U19734 (N_19734,N_15513,N_13900);
or U19735 (N_19735,N_14076,N_14068);
and U19736 (N_19736,N_12358,N_14658);
nor U19737 (N_19737,N_13261,N_15014);
xnor U19738 (N_19738,N_12456,N_15929);
or U19739 (N_19739,N_13156,N_13375);
nor U19740 (N_19740,N_14543,N_12913);
xor U19741 (N_19741,N_14125,N_15796);
nor U19742 (N_19742,N_15525,N_12937);
or U19743 (N_19743,N_14835,N_12076);
xor U19744 (N_19744,N_15772,N_15835);
nor U19745 (N_19745,N_12702,N_14300);
xor U19746 (N_19746,N_12487,N_12439);
nand U19747 (N_19747,N_13719,N_13553);
nand U19748 (N_19748,N_12991,N_13692);
nand U19749 (N_19749,N_12359,N_14095);
and U19750 (N_19750,N_13680,N_14358);
or U19751 (N_19751,N_15656,N_13496);
or U19752 (N_19752,N_14155,N_14525);
nand U19753 (N_19753,N_13782,N_14291);
nor U19754 (N_19754,N_13125,N_13930);
or U19755 (N_19755,N_14027,N_15325);
nand U19756 (N_19756,N_15949,N_15207);
and U19757 (N_19757,N_15242,N_14484);
xnor U19758 (N_19758,N_12528,N_13153);
or U19759 (N_19759,N_14586,N_12697);
nand U19760 (N_19760,N_15814,N_15979);
or U19761 (N_19761,N_15384,N_13292);
or U19762 (N_19762,N_13360,N_12562);
nand U19763 (N_19763,N_15260,N_12973);
nor U19764 (N_19764,N_12893,N_13214);
nand U19765 (N_19765,N_15589,N_15247);
nand U19766 (N_19766,N_15996,N_12937);
or U19767 (N_19767,N_14524,N_15950);
or U19768 (N_19768,N_12219,N_12567);
nand U19769 (N_19769,N_14259,N_12081);
or U19770 (N_19770,N_13692,N_12990);
xor U19771 (N_19771,N_13245,N_12773);
and U19772 (N_19772,N_12835,N_13542);
and U19773 (N_19773,N_15415,N_15084);
or U19774 (N_19774,N_14876,N_14776);
nor U19775 (N_19775,N_14995,N_15220);
or U19776 (N_19776,N_13288,N_15600);
nand U19777 (N_19777,N_12794,N_13213);
or U19778 (N_19778,N_13518,N_13852);
or U19779 (N_19779,N_13850,N_12655);
xnor U19780 (N_19780,N_13077,N_13830);
nor U19781 (N_19781,N_15400,N_12836);
nand U19782 (N_19782,N_12980,N_13976);
or U19783 (N_19783,N_13792,N_14702);
and U19784 (N_19784,N_14740,N_14403);
or U19785 (N_19785,N_15610,N_13810);
nand U19786 (N_19786,N_14701,N_14054);
nand U19787 (N_19787,N_12485,N_12075);
nand U19788 (N_19788,N_14330,N_13849);
and U19789 (N_19789,N_12521,N_15681);
and U19790 (N_19790,N_12855,N_14812);
nand U19791 (N_19791,N_13881,N_12517);
nor U19792 (N_19792,N_15915,N_12625);
xnor U19793 (N_19793,N_15259,N_15551);
nand U19794 (N_19794,N_15697,N_14526);
nor U19795 (N_19795,N_14850,N_14100);
or U19796 (N_19796,N_14777,N_15180);
and U19797 (N_19797,N_13501,N_13699);
and U19798 (N_19798,N_12336,N_14624);
and U19799 (N_19799,N_14353,N_15975);
or U19800 (N_19800,N_15193,N_15962);
xor U19801 (N_19801,N_12127,N_12598);
nand U19802 (N_19802,N_13367,N_13307);
and U19803 (N_19803,N_13555,N_14033);
and U19804 (N_19804,N_13319,N_14284);
nand U19805 (N_19805,N_14008,N_13420);
and U19806 (N_19806,N_13420,N_14313);
nor U19807 (N_19807,N_13622,N_15218);
and U19808 (N_19808,N_12998,N_14876);
xnor U19809 (N_19809,N_14649,N_15271);
and U19810 (N_19810,N_15133,N_12183);
and U19811 (N_19811,N_15662,N_15194);
and U19812 (N_19812,N_14055,N_13556);
and U19813 (N_19813,N_14835,N_15113);
nor U19814 (N_19814,N_13445,N_12257);
xor U19815 (N_19815,N_13650,N_15935);
or U19816 (N_19816,N_15989,N_14145);
xnor U19817 (N_19817,N_13270,N_13149);
xor U19818 (N_19818,N_12929,N_13630);
and U19819 (N_19819,N_12418,N_14219);
or U19820 (N_19820,N_12882,N_14194);
and U19821 (N_19821,N_12672,N_13200);
or U19822 (N_19822,N_15495,N_12804);
and U19823 (N_19823,N_13688,N_15650);
nand U19824 (N_19824,N_14780,N_12742);
or U19825 (N_19825,N_15542,N_12953);
nand U19826 (N_19826,N_15405,N_15158);
or U19827 (N_19827,N_13893,N_14064);
nor U19828 (N_19828,N_15447,N_12489);
xor U19829 (N_19829,N_15538,N_13680);
or U19830 (N_19830,N_14110,N_12810);
or U19831 (N_19831,N_13685,N_14319);
and U19832 (N_19832,N_13079,N_12629);
and U19833 (N_19833,N_14711,N_15141);
nand U19834 (N_19834,N_15682,N_13964);
nand U19835 (N_19835,N_13182,N_12173);
nand U19836 (N_19836,N_15820,N_13140);
xnor U19837 (N_19837,N_13974,N_14836);
and U19838 (N_19838,N_12432,N_15106);
and U19839 (N_19839,N_13818,N_14781);
nor U19840 (N_19840,N_14096,N_12435);
or U19841 (N_19841,N_15919,N_13638);
nand U19842 (N_19842,N_14760,N_13905);
nand U19843 (N_19843,N_15292,N_15694);
nand U19844 (N_19844,N_12587,N_12688);
and U19845 (N_19845,N_12888,N_12546);
xnor U19846 (N_19846,N_13614,N_13261);
nor U19847 (N_19847,N_12532,N_12089);
or U19848 (N_19848,N_12667,N_15228);
and U19849 (N_19849,N_13288,N_12695);
nand U19850 (N_19850,N_12963,N_13521);
or U19851 (N_19851,N_12355,N_15751);
and U19852 (N_19852,N_14504,N_14969);
nor U19853 (N_19853,N_13447,N_14048);
nand U19854 (N_19854,N_15637,N_13445);
and U19855 (N_19855,N_15825,N_15779);
nor U19856 (N_19856,N_14367,N_13584);
nor U19857 (N_19857,N_12252,N_13162);
nor U19858 (N_19858,N_12975,N_12503);
nand U19859 (N_19859,N_13657,N_12581);
nor U19860 (N_19860,N_12653,N_12195);
or U19861 (N_19861,N_14328,N_12845);
and U19862 (N_19862,N_12152,N_13505);
xnor U19863 (N_19863,N_15856,N_13190);
and U19864 (N_19864,N_13500,N_13012);
and U19865 (N_19865,N_12383,N_13676);
xnor U19866 (N_19866,N_12049,N_14943);
or U19867 (N_19867,N_13496,N_12260);
or U19868 (N_19868,N_12454,N_13670);
nand U19869 (N_19869,N_14500,N_13497);
and U19870 (N_19870,N_15792,N_12888);
and U19871 (N_19871,N_13131,N_15310);
nand U19872 (N_19872,N_14301,N_12825);
or U19873 (N_19873,N_14549,N_14570);
xnor U19874 (N_19874,N_13757,N_13335);
or U19875 (N_19875,N_14130,N_14281);
or U19876 (N_19876,N_15023,N_13210);
or U19877 (N_19877,N_12264,N_12731);
and U19878 (N_19878,N_15863,N_12038);
or U19879 (N_19879,N_14000,N_15854);
and U19880 (N_19880,N_13970,N_12826);
nand U19881 (N_19881,N_13422,N_14890);
xor U19882 (N_19882,N_14968,N_14442);
nand U19883 (N_19883,N_15614,N_14707);
and U19884 (N_19884,N_12431,N_14417);
nand U19885 (N_19885,N_14135,N_14092);
nor U19886 (N_19886,N_12901,N_14231);
nor U19887 (N_19887,N_12411,N_15258);
and U19888 (N_19888,N_12884,N_15494);
or U19889 (N_19889,N_14056,N_12455);
nand U19890 (N_19890,N_12348,N_13562);
nor U19891 (N_19891,N_12012,N_13038);
nand U19892 (N_19892,N_13843,N_13624);
nor U19893 (N_19893,N_15429,N_12524);
nand U19894 (N_19894,N_13697,N_13901);
or U19895 (N_19895,N_13435,N_12436);
nand U19896 (N_19896,N_14960,N_15186);
xor U19897 (N_19897,N_14724,N_12743);
or U19898 (N_19898,N_14750,N_13359);
and U19899 (N_19899,N_15313,N_14056);
xor U19900 (N_19900,N_14850,N_14465);
nand U19901 (N_19901,N_12473,N_15153);
nand U19902 (N_19902,N_15353,N_14877);
nand U19903 (N_19903,N_12701,N_12211);
nor U19904 (N_19904,N_13936,N_12030);
nand U19905 (N_19905,N_15836,N_14538);
or U19906 (N_19906,N_14386,N_13164);
xor U19907 (N_19907,N_13328,N_12523);
nor U19908 (N_19908,N_13710,N_12102);
xor U19909 (N_19909,N_12177,N_13175);
or U19910 (N_19910,N_13966,N_13040);
nor U19911 (N_19911,N_13952,N_15422);
or U19912 (N_19912,N_12944,N_14630);
or U19913 (N_19913,N_14281,N_15765);
nand U19914 (N_19914,N_15343,N_15997);
xor U19915 (N_19915,N_12236,N_12207);
and U19916 (N_19916,N_13434,N_12834);
xnor U19917 (N_19917,N_12072,N_12587);
xnor U19918 (N_19918,N_14206,N_13616);
xnor U19919 (N_19919,N_12889,N_15685);
or U19920 (N_19920,N_15386,N_15504);
xnor U19921 (N_19921,N_13019,N_12547);
nor U19922 (N_19922,N_15572,N_13340);
nor U19923 (N_19923,N_12996,N_14953);
nor U19924 (N_19924,N_15616,N_12472);
nand U19925 (N_19925,N_14147,N_13682);
or U19926 (N_19926,N_14220,N_13325);
nor U19927 (N_19927,N_15171,N_12593);
xor U19928 (N_19928,N_15829,N_14896);
xor U19929 (N_19929,N_13091,N_14395);
nor U19930 (N_19930,N_15744,N_14743);
nor U19931 (N_19931,N_12352,N_12437);
xor U19932 (N_19932,N_14448,N_13283);
nand U19933 (N_19933,N_14104,N_13928);
and U19934 (N_19934,N_13815,N_12607);
xnor U19935 (N_19935,N_13587,N_12667);
nand U19936 (N_19936,N_12671,N_12376);
nand U19937 (N_19937,N_12963,N_15789);
or U19938 (N_19938,N_15558,N_12790);
nand U19939 (N_19939,N_15818,N_14310);
xnor U19940 (N_19940,N_13970,N_12167);
xor U19941 (N_19941,N_12852,N_14331);
nor U19942 (N_19942,N_15359,N_12042);
nor U19943 (N_19943,N_14639,N_13599);
xnor U19944 (N_19944,N_12631,N_12478);
nand U19945 (N_19945,N_14746,N_12791);
xnor U19946 (N_19946,N_14286,N_14441);
xnor U19947 (N_19947,N_12986,N_15371);
or U19948 (N_19948,N_13300,N_15862);
nand U19949 (N_19949,N_12203,N_12740);
and U19950 (N_19950,N_14988,N_15498);
nand U19951 (N_19951,N_13691,N_14947);
or U19952 (N_19952,N_12626,N_13262);
nand U19953 (N_19953,N_15803,N_14196);
xor U19954 (N_19954,N_15552,N_12277);
nor U19955 (N_19955,N_14539,N_14693);
or U19956 (N_19956,N_13275,N_14426);
nor U19957 (N_19957,N_14282,N_14126);
nand U19958 (N_19958,N_15215,N_15030);
nor U19959 (N_19959,N_14090,N_15058);
or U19960 (N_19960,N_13710,N_15563);
nand U19961 (N_19961,N_12499,N_12686);
nor U19962 (N_19962,N_14579,N_15819);
or U19963 (N_19963,N_12131,N_14072);
and U19964 (N_19964,N_15114,N_15937);
nor U19965 (N_19965,N_12424,N_13809);
or U19966 (N_19966,N_13860,N_12301);
nand U19967 (N_19967,N_14973,N_15423);
nor U19968 (N_19968,N_13122,N_15028);
or U19969 (N_19969,N_15881,N_13064);
xnor U19970 (N_19970,N_12758,N_15668);
nand U19971 (N_19971,N_15706,N_15762);
xnor U19972 (N_19972,N_12574,N_15389);
nand U19973 (N_19973,N_15349,N_14673);
or U19974 (N_19974,N_13085,N_13463);
nand U19975 (N_19975,N_12265,N_14267);
nor U19976 (N_19976,N_15725,N_15348);
and U19977 (N_19977,N_14072,N_15703);
or U19978 (N_19978,N_15574,N_12087);
and U19979 (N_19979,N_15514,N_13415);
nor U19980 (N_19980,N_13187,N_14216);
xnor U19981 (N_19981,N_12147,N_15290);
nor U19982 (N_19982,N_12037,N_12373);
nand U19983 (N_19983,N_15815,N_14469);
nor U19984 (N_19984,N_13794,N_12569);
and U19985 (N_19985,N_13632,N_14763);
xor U19986 (N_19986,N_12944,N_14009);
xnor U19987 (N_19987,N_14315,N_15375);
nor U19988 (N_19988,N_14425,N_15279);
xnor U19989 (N_19989,N_15068,N_15908);
or U19990 (N_19990,N_13934,N_12390);
xor U19991 (N_19991,N_15846,N_14559);
xnor U19992 (N_19992,N_15620,N_15480);
nor U19993 (N_19993,N_15034,N_15452);
nand U19994 (N_19994,N_14302,N_12372);
nand U19995 (N_19995,N_12761,N_13171);
nor U19996 (N_19996,N_14928,N_14408);
xor U19997 (N_19997,N_14286,N_15366);
nand U19998 (N_19998,N_15695,N_12115);
or U19999 (N_19999,N_15883,N_13020);
xnor UO_0 (O_0,N_18873,N_17602);
nand UO_1 (O_1,N_18072,N_16669);
nor UO_2 (O_2,N_16338,N_18636);
nand UO_3 (O_3,N_18026,N_19184);
nor UO_4 (O_4,N_16800,N_17910);
xor UO_5 (O_5,N_17543,N_18939);
or UO_6 (O_6,N_18104,N_18685);
or UO_7 (O_7,N_17030,N_19829);
nand UO_8 (O_8,N_18421,N_19549);
or UO_9 (O_9,N_17811,N_16605);
nor UO_10 (O_10,N_16103,N_16494);
nand UO_11 (O_11,N_17717,N_16365);
nand UO_12 (O_12,N_19617,N_19582);
xor UO_13 (O_13,N_18438,N_19873);
xnor UO_14 (O_14,N_18342,N_16948);
nor UO_15 (O_15,N_19440,N_16563);
nand UO_16 (O_16,N_17260,N_19914);
xor UO_17 (O_17,N_17677,N_17705);
xor UO_18 (O_18,N_16364,N_17386);
nor UO_19 (O_19,N_18220,N_17970);
nand UO_20 (O_20,N_18721,N_16144);
or UO_21 (O_21,N_16612,N_17274);
or UO_22 (O_22,N_16092,N_19010);
xor UO_23 (O_23,N_19232,N_17762);
nor UO_24 (O_24,N_17001,N_16936);
and UO_25 (O_25,N_19331,N_17091);
nor UO_26 (O_26,N_18248,N_18491);
xnor UO_27 (O_27,N_18573,N_17204);
nor UO_28 (O_28,N_19485,N_18098);
or UO_29 (O_29,N_18890,N_19187);
or UO_30 (O_30,N_17381,N_17066);
xnor UO_31 (O_31,N_16055,N_16792);
nand UO_32 (O_32,N_16396,N_16973);
nor UO_33 (O_33,N_18510,N_16705);
or UO_34 (O_34,N_17930,N_17799);
or UO_35 (O_35,N_16916,N_16772);
nand UO_36 (O_36,N_17002,N_18879);
nor UO_37 (O_37,N_19385,N_19124);
xnor UO_38 (O_38,N_17610,N_17908);
or UO_39 (O_39,N_19116,N_19195);
nor UO_40 (O_40,N_16725,N_17258);
xor UO_41 (O_41,N_16521,N_18909);
and UO_42 (O_42,N_16013,N_18087);
or UO_43 (O_43,N_17807,N_18019);
and UO_44 (O_44,N_17335,N_17311);
or UO_45 (O_45,N_17620,N_18336);
nor UO_46 (O_46,N_19981,N_17332);
or UO_47 (O_47,N_19655,N_17409);
or UO_48 (O_48,N_17178,N_18004);
or UO_49 (O_49,N_16397,N_17388);
nand UO_50 (O_50,N_19310,N_17545);
or UO_51 (O_51,N_17623,N_16188);
or UO_52 (O_52,N_16529,N_17429);
xnor UO_53 (O_53,N_18828,N_16415);
nor UO_54 (O_54,N_16880,N_19021);
xor UO_55 (O_55,N_18807,N_19588);
nor UO_56 (O_56,N_16052,N_19567);
xor UO_57 (O_57,N_16440,N_19715);
nand UO_58 (O_58,N_17188,N_17995);
or UO_59 (O_59,N_16629,N_19785);
xor UO_60 (O_60,N_16147,N_19740);
xor UO_61 (O_61,N_17529,N_18758);
or UO_62 (O_62,N_17627,N_19418);
nor UO_63 (O_63,N_16582,N_17794);
or UO_64 (O_64,N_16622,N_19692);
nand UO_65 (O_65,N_16630,N_18922);
xnor UO_66 (O_66,N_17916,N_19060);
xor UO_67 (O_67,N_16924,N_16565);
nor UO_68 (O_68,N_18221,N_16340);
or UO_69 (O_69,N_19201,N_17975);
xor UO_70 (O_70,N_19601,N_17730);
or UO_71 (O_71,N_18040,N_19275);
or UO_72 (O_72,N_18205,N_17185);
nor UO_73 (O_73,N_16229,N_16568);
xor UO_74 (O_74,N_16575,N_17537);
xnor UO_75 (O_75,N_19085,N_17437);
and UO_76 (O_76,N_18419,N_19545);
nand UO_77 (O_77,N_19600,N_18151);
nand UO_78 (O_78,N_18899,N_17798);
nor UO_79 (O_79,N_17329,N_18688);
or UO_80 (O_80,N_17160,N_17723);
or UO_81 (O_81,N_16865,N_16222);
nor UO_82 (O_82,N_17552,N_16555);
xor UO_83 (O_83,N_17861,N_19780);
nand UO_84 (O_84,N_19927,N_17046);
nor UO_85 (O_85,N_18167,N_16448);
and UO_86 (O_86,N_18918,N_17391);
nand UO_87 (O_87,N_16495,N_16053);
nor UO_88 (O_88,N_19076,N_19098);
nor UO_89 (O_89,N_19609,N_16118);
and UO_90 (O_90,N_18191,N_16993);
nand UO_91 (O_91,N_18207,N_17561);
nor UO_92 (O_92,N_19965,N_18204);
nor UO_93 (O_93,N_16351,N_16295);
or UO_94 (O_94,N_19604,N_18484);
and UO_95 (O_95,N_19226,N_19828);
and UO_96 (O_96,N_17064,N_16580);
and UO_97 (O_97,N_17467,N_18679);
nor UO_98 (O_98,N_17588,N_19401);
nor UO_99 (O_99,N_16171,N_18812);
and UO_100 (O_100,N_19213,N_17351);
and UO_101 (O_101,N_18306,N_18970);
and UO_102 (O_102,N_16766,N_16095);
and UO_103 (O_103,N_18780,N_18941);
or UO_104 (O_104,N_16793,N_17431);
and UO_105 (O_105,N_19050,N_17031);
nand UO_106 (O_106,N_18340,N_17748);
and UO_107 (O_107,N_19728,N_19653);
and UO_108 (O_108,N_19228,N_16806);
or UO_109 (O_109,N_17683,N_18494);
xor UO_110 (O_110,N_18990,N_19411);
nand UO_111 (O_111,N_19542,N_17816);
and UO_112 (O_112,N_18471,N_17339);
nand UO_113 (O_113,N_18328,N_19413);
nand UO_114 (O_114,N_16434,N_16400);
or UO_115 (O_115,N_18163,N_17344);
and UO_116 (O_116,N_19796,N_18963);
or UO_117 (O_117,N_18566,N_17096);
nor UO_118 (O_118,N_16598,N_17439);
or UO_119 (O_119,N_16911,N_16818);
and UO_120 (O_120,N_18582,N_17461);
xnor UO_121 (O_121,N_16848,N_16492);
and UO_122 (O_122,N_19465,N_16234);
nor UO_123 (O_123,N_16411,N_19649);
or UO_124 (O_124,N_16853,N_19886);
or UO_125 (O_125,N_17896,N_19838);
and UO_126 (O_126,N_16301,N_16697);
and UO_127 (O_127,N_18614,N_17215);
and UO_128 (O_128,N_18876,N_19816);
and UO_129 (O_129,N_17474,N_18991);
nand UO_130 (O_130,N_19335,N_16657);
or UO_131 (O_131,N_18803,N_16695);
nand UO_132 (O_132,N_17140,N_19526);
xnor UO_133 (O_133,N_17590,N_19951);
and UO_134 (O_134,N_17352,N_17769);
nor UO_135 (O_135,N_16442,N_19803);
nand UO_136 (O_136,N_18794,N_17507);
nand UO_137 (O_137,N_19598,N_17736);
xor UO_138 (O_138,N_17019,N_17987);
nand UO_139 (O_139,N_16341,N_19665);
or UO_140 (O_140,N_19267,N_16775);
nor UO_141 (O_141,N_19845,N_17435);
nor UO_142 (O_142,N_18028,N_16759);
and UO_143 (O_143,N_17129,N_19202);
nand UO_144 (O_144,N_18635,N_19778);
and UO_145 (O_145,N_16783,N_16162);
xnor UO_146 (O_146,N_19141,N_19521);
xor UO_147 (O_147,N_16734,N_19972);
xnor UO_148 (O_148,N_16843,N_16032);
or UO_149 (O_149,N_18293,N_19954);
and UO_150 (O_150,N_19580,N_17781);
nand UO_151 (O_151,N_19307,N_19462);
nor UO_152 (O_152,N_16597,N_17396);
nor UO_153 (O_153,N_18746,N_19039);
xnor UO_154 (O_154,N_18795,N_17950);
and UO_155 (O_155,N_18784,N_19475);
nand UO_156 (O_156,N_17082,N_18574);
nand UO_157 (O_157,N_16919,N_19057);
xnor UO_158 (O_158,N_19662,N_19742);
xor UO_159 (O_159,N_18928,N_18280);
and UO_160 (O_160,N_19253,N_19702);
and UO_161 (O_161,N_19594,N_16861);
nand UO_162 (O_162,N_17826,N_17061);
nor UO_163 (O_163,N_18558,N_18198);
xnor UO_164 (O_164,N_18196,N_18069);
xor UO_165 (O_165,N_19164,N_16438);
xnor UO_166 (O_166,N_17808,N_19833);
nor UO_167 (O_167,N_16077,N_17733);
nor UO_168 (O_168,N_16286,N_18039);
or UO_169 (O_169,N_17323,N_18545);
or UO_170 (O_170,N_16586,N_17279);
nand UO_171 (O_171,N_19309,N_16285);
nor UO_172 (O_172,N_17532,N_16296);
and UO_173 (O_173,N_18121,N_18531);
nand UO_174 (O_174,N_16639,N_17731);
and UO_175 (O_175,N_19717,N_17138);
nor UO_176 (O_176,N_17810,N_19325);
or UO_177 (O_177,N_18470,N_16422);
or UO_178 (O_178,N_19033,N_17951);
nand UO_179 (O_179,N_19864,N_19221);
nor UO_180 (O_180,N_17199,N_16302);
and UO_181 (O_181,N_17593,N_19119);
and UO_182 (O_182,N_16500,N_19952);
or UO_183 (O_183,N_19442,N_17221);
nand UO_184 (O_184,N_17471,N_17098);
and UO_185 (O_185,N_16029,N_18715);
and UO_186 (O_186,N_18355,N_19009);
xnor UO_187 (O_187,N_17051,N_16122);
nor UO_188 (O_188,N_17747,N_18144);
nor UO_189 (O_189,N_19509,N_19049);
nand UO_190 (O_190,N_19869,N_17516);
or UO_191 (O_191,N_19245,N_16215);
nor UO_192 (O_192,N_18923,N_19476);
xor UO_193 (O_193,N_17006,N_19751);
and UO_194 (O_194,N_16617,N_19459);
or UO_195 (O_195,N_16857,N_18997);
nor UO_196 (O_196,N_18010,N_17058);
or UO_197 (O_197,N_17139,N_18792);
nand UO_198 (O_198,N_17008,N_16659);
xnor UO_199 (O_199,N_17553,N_18388);
xnor UO_200 (O_200,N_18366,N_16418);
nand UO_201 (O_201,N_18849,N_19054);
nand UO_202 (O_202,N_16814,N_18783);
or UO_203 (O_203,N_18360,N_19846);
xor UO_204 (O_204,N_16967,N_17976);
nor UO_205 (O_205,N_17034,N_17792);
or UO_206 (O_206,N_16955,N_18641);
nand UO_207 (O_207,N_19678,N_16940);
nand UO_208 (O_208,N_19095,N_18344);
xor UO_209 (O_209,N_16807,N_17660);
or UO_210 (O_210,N_16128,N_17982);
nand UO_211 (O_211,N_18983,N_19059);
xor UO_212 (O_212,N_16483,N_19387);
nand UO_213 (O_213,N_17394,N_19613);
or UO_214 (O_214,N_19020,N_17174);
or UO_215 (O_215,N_17420,N_17918);
xor UO_216 (O_216,N_16124,N_16196);
nor UO_217 (O_217,N_19908,N_19987);
and UO_218 (O_218,N_16997,N_17067);
xnor UO_219 (O_219,N_19859,N_18933);
xnor UO_220 (O_220,N_17922,N_16975);
nor UO_221 (O_221,N_19641,N_18393);
or UO_222 (O_222,N_16879,N_19605);
xnor UO_223 (O_223,N_19384,N_18569);
nor UO_224 (O_224,N_16712,N_19279);
nor UO_225 (O_225,N_16675,N_17669);
nor UO_226 (O_226,N_16871,N_16211);
nand UO_227 (O_227,N_19166,N_18521);
and UO_228 (O_228,N_18414,N_16877);
and UO_229 (O_229,N_16497,N_16511);
xnor UO_230 (O_230,N_17121,N_19262);
and UO_231 (O_231,N_19224,N_18498);
or UO_232 (O_232,N_16944,N_17497);
nand UO_233 (O_233,N_16540,N_19007);
nand UO_234 (O_234,N_19808,N_17978);
nor UO_235 (O_235,N_17889,N_17354);
nand UO_236 (O_236,N_19817,N_18013);
nand UO_237 (O_237,N_17741,N_18593);
xnor UO_238 (O_238,N_16904,N_17618);
xnor UO_239 (O_239,N_19676,N_18822);
nand UO_240 (O_240,N_16374,N_16874);
or UO_241 (O_241,N_17390,N_17210);
xor UO_242 (O_242,N_18063,N_18088);
nor UO_243 (O_243,N_17812,N_16887);
and UO_244 (O_244,N_18297,N_19337);
xor UO_245 (O_245,N_18245,N_16932);
nand UO_246 (O_246,N_18985,N_17648);
or UO_247 (O_247,N_18691,N_19243);
or UO_248 (O_248,N_16031,N_16724);
nand UO_249 (O_249,N_18612,N_18678);
and UO_250 (O_250,N_16957,N_18870);
xnor UO_251 (O_251,N_19242,N_17696);
and UO_252 (O_252,N_18423,N_18193);
or UO_253 (O_253,N_16961,N_17301);
nand UO_254 (O_254,N_17007,N_17206);
xnor UO_255 (O_255,N_16729,N_16140);
or UO_256 (O_256,N_18056,N_18606);
and UO_257 (O_257,N_17992,N_16832);
and UO_258 (O_258,N_17321,N_17688);
xnor UO_259 (O_259,N_19455,N_17695);
nor UO_260 (O_260,N_18134,N_16007);
nand UO_261 (O_261,N_17805,N_17433);
and UO_262 (O_262,N_17374,N_18238);
or UO_263 (O_263,N_17789,N_19703);
and UO_264 (O_264,N_19278,N_19274);
xor UO_265 (O_265,N_16737,N_19830);
nor UO_266 (O_266,N_16674,N_18886);
or UO_267 (O_267,N_16363,N_16572);
or UO_268 (O_268,N_17740,N_19088);
xnor UO_269 (O_269,N_19506,N_18829);
xnor UO_270 (O_270,N_19924,N_18848);
or UO_271 (O_271,N_17631,N_17614);
nor UO_272 (O_272,N_18754,N_19394);
and UO_273 (O_273,N_18620,N_16837);
nor UO_274 (O_274,N_18047,N_18753);
and UO_275 (O_275,N_16966,N_17304);
xnor UO_276 (O_276,N_17299,N_17528);
nand UO_277 (O_277,N_18321,N_19848);
nor UO_278 (O_278,N_18960,N_18251);
nand UO_279 (O_279,N_17824,N_19937);
and UO_280 (O_280,N_16036,N_19448);
nand UO_281 (O_281,N_16349,N_18206);
and UO_282 (O_282,N_16123,N_17542);
and UO_283 (O_283,N_16048,N_17270);
or UO_284 (O_284,N_18506,N_16256);
nor UO_285 (O_285,N_16370,N_18209);
nor UO_286 (O_286,N_16947,N_16163);
nand UO_287 (O_287,N_16509,N_18239);
or UO_288 (O_288,N_16548,N_16361);
nor UO_289 (O_289,N_17447,N_19263);
nand UO_290 (O_290,N_16709,N_17926);
and UO_291 (O_291,N_16010,N_18046);
and UO_292 (O_292,N_17925,N_19167);
nor UO_293 (O_293,N_19212,N_16628);
or UO_294 (O_294,N_19332,N_18045);
or UO_295 (O_295,N_16112,N_17266);
nor UO_296 (O_296,N_19031,N_18347);
and UO_297 (O_297,N_17856,N_17653);
nand UO_298 (O_298,N_17906,N_19960);
xor UO_299 (O_299,N_16332,N_16569);
and UO_300 (O_300,N_19921,N_17591);
nor UO_301 (O_301,N_19823,N_17452);
xor UO_302 (O_302,N_18623,N_16551);
or UO_303 (O_303,N_18589,N_16658);
xor UO_304 (O_304,N_19342,N_17133);
xnor UO_305 (O_305,N_19392,N_16868);
and UO_306 (O_306,N_18392,N_18730);
nand UO_307 (O_307,N_19423,N_16412);
nor UO_308 (O_308,N_17693,N_19273);
nor UO_309 (O_309,N_16337,N_19416);
nand UO_310 (O_310,N_16428,N_18843);
nand UO_311 (O_311,N_19320,N_17687);
nand UO_312 (O_312,N_17005,N_17626);
xnor UO_313 (O_313,N_18583,N_18952);
nor UO_314 (O_314,N_17904,N_16938);
xor UO_315 (O_315,N_17276,N_17905);
nor UO_316 (O_316,N_18290,N_16976);
nand UO_317 (O_317,N_18698,N_19318);
or UO_318 (O_318,N_17087,N_16891);
nor UO_319 (O_319,N_17974,N_17491);
xnor UO_320 (O_320,N_19438,N_18141);
or UO_321 (O_321,N_16039,N_17080);
xnor UO_322 (O_322,N_19074,N_18402);
xor UO_323 (O_323,N_18676,N_16684);
nor UO_324 (O_324,N_19984,N_18846);
and UO_325 (O_325,N_19659,N_18858);
or UO_326 (O_326,N_17745,N_16860);
nor UO_327 (O_327,N_18362,N_18428);
or UO_328 (O_328,N_16149,N_16813);
nand UO_329 (O_329,N_17913,N_16009);
or UO_330 (O_330,N_18109,N_17343);
and UO_331 (O_331,N_18756,N_18687);
xnor UO_332 (O_332,N_17057,N_18027);
xor UO_333 (O_333,N_19541,N_19001);
nand UO_334 (O_334,N_16290,N_19053);
or UO_335 (O_335,N_18229,N_19186);
nor UO_336 (O_336,N_16786,N_18572);
nor UO_337 (O_337,N_17103,N_16210);
and UO_338 (O_338,N_19566,N_19943);
and UO_339 (O_339,N_17457,N_19695);
nand UO_340 (O_340,N_16405,N_16816);
or UO_341 (O_341,N_17242,N_18301);
and UO_342 (O_342,N_16246,N_18811);
or UO_343 (O_343,N_16012,N_17010);
or UO_344 (O_344,N_18618,N_16959);
nor UO_345 (O_345,N_17192,N_19866);
and UO_346 (O_346,N_17795,N_17700);
or UO_347 (O_347,N_18009,N_19317);
nand UO_348 (O_348,N_17999,N_18259);
and UO_349 (O_349,N_16858,N_17126);
xnor UO_350 (O_350,N_16579,N_18775);
xor UO_351 (O_351,N_18814,N_17981);
nand UO_352 (O_352,N_17797,N_16672);
or UO_353 (O_353,N_16269,N_18008);
nand UO_354 (O_354,N_18078,N_18339);
nand UO_355 (O_355,N_17224,N_18197);
nor UO_356 (O_356,N_19065,N_17081);
xor UO_357 (O_357,N_17099,N_16476);
or UO_358 (O_358,N_17013,N_17621);
nand UO_359 (O_359,N_17630,N_16040);
and UO_360 (O_360,N_17572,N_18847);
or UO_361 (O_361,N_19732,N_17968);
and UO_362 (O_362,N_19764,N_18439);
xor UO_363 (O_363,N_16272,N_19302);
and UO_364 (O_364,N_18090,N_19269);
nor UO_365 (O_365,N_16063,N_19922);
nand UO_366 (O_366,N_18714,N_16541);
nand UO_367 (O_367,N_18469,N_18995);
nand UO_368 (O_368,N_19532,N_18560);
nor UO_369 (O_369,N_19435,N_19109);
nor UO_370 (O_370,N_16232,N_19086);
or UO_371 (O_371,N_19963,N_16248);
nand UO_372 (O_372,N_19658,N_18967);
or UO_373 (O_373,N_19040,N_17229);
nor UO_374 (O_374,N_19348,N_18595);
or UO_375 (O_375,N_16304,N_16158);
or UO_376 (O_376,N_19589,N_16207);
nand UO_377 (O_377,N_17763,N_17036);
nor UO_378 (O_378,N_19378,N_18869);
nand UO_379 (O_379,N_16965,N_17619);
nand UO_380 (O_380,N_17316,N_16869);
and UO_381 (O_381,N_19622,N_18789);
xnor UO_382 (O_382,N_19953,N_19755);
nor UO_383 (O_383,N_19078,N_18271);
nand UO_384 (O_384,N_17165,N_17211);
xnor UO_385 (O_385,N_17181,N_18645);
nand UO_386 (O_386,N_18683,N_18946);
nor UO_387 (O_387,N_17832,N_16165);
or UO_388 (O_388,N_18887,N_17681);
xnor UO_389 (O_389,N_17047,N_17800);
or UO_390 (O_390,N_16291,N_16485);
or UO_391 (O_391,N_18845,N_16173);
xor UO_392 (O_392,N_18661,N_16864);
or UO_393 (O_393,N_18124,N_16836);
nor UO_394 (O_394,N_16876,N_17515);
or UO_395 (O_395,N_18894,N_16604);
and UO_396 (O_396,N_18526,N_16022);
nor UO_397 (O_397,N_18628,N_17370);
nor UO_398 (O_398,N_17408,N_16177);
xor UO_399 (O_399,N_16567,N_16120);
nand UO_400 (O_400,N_19868,N_17407);
or UO_401 (O_401,N_19806,N_17074);
nor UO_402 (O_402,N_16473,N_17658);
or UO_403 (O_403,N_17387,N_17715);
and UO_404 (O_404,N_19569,N_18020);
nand UO_405 (O_405,N_19558,N_17149);
nor UO_406 (O_406,N_19290,N_16688);
nand UO_407 (O_407,N_16606,N_19568);
or UO_408 (O_408,N_17871,N_18559);
nor UO_409 (O_409,N_16525,N_17060);
xnor UO_410 (O_410,N_16518,N_18189);
nand UO_411 (O_411,N_16257,N_18318);
xnor UO_412 (O_412,N_19469,N_19134);
xnor UO_413 (O_413,N_17110,N_16827);
nor UO_414 (O_414,N_16757,N_19013);
nand UO_415 (O_415,N_19673,N_18652);
nor UO_416 (O_416,N_16047,N_16206);
or UO_417 (O_417,N_18910,N_19259);
and UO_418 (O_418,N_17540,N_18654);
nand UO_419 (O_419,N_16951,N_19068);
and UO_420 (O_420,N_16648,N_18773);
xnor UO_421 (O_421,N_16192,N_18330);
xnor UO_422 (O_422,N_17783,N_16321);
and UO_423 (O_423,N_16401,N_19019);
or UO_424 (O_424,N_19241,N_18587);
nor UO_425 (O_425,N_17845,N_18668);
nor UO_426 (O_426,N_18865,N_18584);
and UO_427 (O_427,N_17765,N_17434);
and UO_428 (O_428,N_19888,N_19280);
nand UO_429 (O_429,N_19883,N_16949);
and UO_430 (O_430,N_17840,N_19794);
nor UO_431 (O_431,N_18455,N_18424);
nor UO_432 (O_432,N_19524,N_18037);
nand UO_433 (O_433,N_16941,N_17701);
nand UO_434 (O_434,N_19691,N_18103);
nor UO_435 (O_435,N_16897,N_16933);
nand UO_436 (O_436,N_16150,N_18123);
nand UO_437 (O_437,N_17377,N_17484);
and UO_438 (O_438,N_18228,N_19386);
or UO_439 (O_439,N_19327,N_19998);
or UO_440 (O_440,N_17719,N_17654);
nand UO_441 (O_441,N_19672,N_17600);
or UO_442 (O_442,N_19235,N_17865);
xor UO_443 (O_443,N_17038,N_17668);
and UO_444 (O_444,N_18079,N_18361);
or UO_445 (O_445,N_17548,N_19491);
xnor UO_446 (O_446,N_19895,N_18354);
nand UO_447 (O_447,N_17170,N_19284);
nor UO_448 (O_448,N_16530,N_17326);
and UO_449 (O_449,N_16570,N_18317);
xnor UO_450 (O_450,N_18826,N_19457);
xor UO_451 (O_451,N_19204,N_18519);
nor UO_452 (O_452,N_18703,N_19536);
and UO_453 (O_453,N_18158,N_19766);
xnor UO_454 (O_454,N_17971,N_19073);
nor UO_455 (O_455,N_19412,N_16840);
xor UO_456 (O_456,N_19777,N_17694);
xnor UO_457 (O_457,N_19756,N_17450);
nor UO_458 (O_458,N_18182,N_18252);
or UO_459 (O_459,N_16381,N_19490);
and UO_460 (O_460,N_17283,N_19807);
or UO_461 (O_461,N_16693,N_19648);
nor UO_462 (O_462,N_18854,N_18500);
nor UO_463 (O_463,N_18278,N_17116);
nor UO_464 (O_464,N_16716,N_19852);
or UO_465 (O_465,N_16805,N_19961);
or UO_466 (O_466,N_19391,N_17936);
nand UO_467 (O_467,N_18649,N_16991);
nor UO_468 (O_468,N_18647,N_18254);
nor UO_469 (O_469,N_19495,N_16421);
xnor UO_470 (O_470,N_16611,N_17559);
xnor UO_471 (O_471,N_18324,N_17164);
or UO_472 (O_472,N_19429,N_19281);
nand UO_473 (O_473,N_18266,N_18375);
and UO_474 (O_474,N_18700,N_18871);
and UO_475 (O_475,N_19393,N_17369);
nor UO_476 (O_476,N_17606,N_17834);
or UO_477 (O_477,N_18808,N_17758);
xnor UO_478 (O_478,N_19017,N_19805);
and UO_479 (O_479,N_17493,N_18949);
nor UO_480 (O_480,N_16602,N_17337);
and UO_481 (O_481,N_16527,N_18187);
nand UO_482 (O_482,N_16553,N_17020);
xnor UO_483 (O_483,N_19379,N_16803);
and UO_484 (O_484,N_19355,N_19107);
nor UO_485 (O_485,N_19901,N_16952);
or UO_486 (O_486,N_16252,N_16204);
nand UO_487 (O_487,N_17703,N_17359);
xnor UO_488 (O_488,N_16668,N_19688);
and UO_489 (O_489,N_19158,N_18068);
and UO_490 (O_490,N_16559,N_18260);
and UO_491 (O_491,N_17044,N_19191);
and UO_492 (O_492,N_17893,N_19419);
and UO_493 (O_493,N_16119,N_17287);
and UO_494 (O_494,N_16892,N_17252);
or UO_495 (O_495,N_18660,N_18077);
and UO_496 (O_496,N_18003,N_16956);
nor UO_497 (O_497,N_19697,N_18288);
nor UO_498 (O_498,N_18666,N_19163);
or UO_499 (O_499,N_17857,N_17514);
nand UO_500 (O_500,N_18214,N_16596);
or UO_501 (O_501,N_16532,N_19559);
and UO_502 (O_502,N_17280,N_18931);
nor UO_503 (O_503,N_17836,N_17644);
nand UO_504 (O_504,N_19523,N_18480);
xnor UO_505 (O_505,N_18371,N_19140);
and UO_506 (O_506,N_18255,N_16578);
xnor UO_507 (O_507,N_18993,N_18749);
and UO_508 (O_508,N_16071,N_18049);
and UO_509 (O_509,N_17285,N_18166);
and UO_510 (O_510,N_18016,N_16576);
nor UO_511 (O_511,N_19397,N_17888);
xnor UO_512 (O_512,N_17458,N_19510);
and UO_513 (O_513,N_17937,N_16319);
and UO_514 (O_514,N_17053,N_16213);
or UO_515 (O_515,N_17817,N_16846);
nor UO_516 (O_516,N_18707,N_16652);
xor UO_517 (O_517,N_16809,N_18951);
or UO_518 (O_518,N_19103,N_17293);
xnor UO_519 (O_519,N_18674,N_19871);
nand UO_520 (O_520,N_19497,N_18523);
xor UO_521 (O_521,N_18074,N_16076);
nand UO_522 (O_522,N_18955,N_17646);
and UO_523 (O_523,N_17468,N_16732);
nand UO_524 (O_524,N_19718,N_16318);
nand UO_525 (O_525,N_19209,N_18102);
nand UO_526 (O_526,N_16186,N_19400);
and UO_527 (O_527,N_16808,N_16661);
xor UO_528 (O_528,N_17163,N_18242);
nand UO_529 (O_529,N_19389,N_19360);
nand UO_530 (O_530,N_16486,N_18508);
nor UO_531 (O_531,N_16627,N_18053);
nand UO_532 (O_532,N_16034,N_16902);
or UO_533 (O_533,N_18834,N_17508);
or UO_534 (O_534,N_16056,N_18289);
and UO_535 (O_535,N_16739,N_19652);
xnor UO_536 (O_536,N_16758,N_18801);
nand UO_537 (O_537,N_19159,N_19251);
or UO_538 (O_538,N_19172,N_18724);
nand UO_539 (O_539,N_16852,N_16574);
nor UO_540 (O_540,N_16680,N_18790);
xor UO_541 (O_541,N_19029,N_17902);
and UO_542 (O_542,N_18999,N_17297);
or UO_543 (O_543,N_16824,N_18409);
nor UO_544 (O_544,N_19923,N_19002);
xnor UO_545 (O_545,N_16741,N_18201);
nor UO_546 (O_546,N_18374,N_17362);
nor UO_547 (O_547,N_18132,N_17613);
and UO_548 (O_548,N_17510,N_16273);
xor UO_549 (O_549,N_18607,N_16182);
or UO_550 (O_550,N_17428,N_19727);
and UO_551 (O_551,N_19881,N_18296);
xor UO_552 (O_552,N_16426,N_18334);
nand UO_553 (O_553,N_17547,N_17504);
nor UO_554 (O_554,N_17023,N_18917);
and UO_555 (O_555,N_16898,N_17453);
and UO_556 (O_556,N_19441,N_18203);
xnor UO_557 (O_557,N_19080,N_18598);
nor UO_558 (O_558,N_17322,N_17875);
xnor UO_559 (O_559,N_16603,N_19346);
xor UO_560 (O_560,N_17942,N_19032);
and UO_561 (O_561,N_18195,N_18373);
and UO_562 (O_562,N_19878,N_18675);
or UO_563 (O_563,N_18954,N_16375);
nor UO_564 (O_564,N_19978,N_19237);
or UO_565 (O_565,N_19716,N_17526);
or UO_566 (O_566,N_17330,N_17151);
and UO_567 (O_567,N_18934,N_16749);
nor UO_568 (O_568,N_16624,N_18329);
and UO_569 (O_569,N_18957,N_16691);
xor UO_570 (O_570,N_17897,N_18530);
xnor UO_571 (O_571,N_19528,N_16625);
xnor UO_572 (O_572,N_19576,N_17112);
and UO_573 (O_573,N_19783,N_16581);
xor UO_574 (O_574,N_18611,N_16347);
and UO_575 (O_575,N_17194,N_19350);
and UO_576 (O_576,N_16125,N_17900);
xor UO_577 (O_577,N_18128,N_18541);
nand UO_578 (O_578,N_18307,N_17774);
nand UO_579 (O_579,N_17785,N_16398);
nor UO_580 (O_580,N_17964,N_16504);
and UO_581 (O_581,N_18457,N_17488);
nor UO_582 (O_582,N_18819,N_19449);
or UO_583 (O_583,N_17403,N_19862);
or UO_584 (O_584,N_17259,N_17402);
xnor UO_585 (O_585,N_18425,N_19198);
or UO_586 (O_586,N_16673,N_19188);
xnor UO_587 (O_587,N_16255,N_17635);
nand UO_588 (O_588,N_19724,N_17176);
or UO_589 (O_589,N_18552,N_19644);
and UO_590 (O_590,N_18921,N_16353);
or UO_591 (O_591,N_17177,N_19127);
and UO_592 (O_592,N_16804,N_16621);
or UO_593 (O_593,N_18322,N_16084);
xnor UO_594 (O_594,N_18720,N_18627);
nor UO_595 (O_595,N_17024,N_19847);
xor UO_596 (O_596,N_16240,N_18159);
xnor UO_597 (O_597,N_18616,N_16841);
xnor UO_598 (O_598,N_17440,N_18608);
or UO_599 (O_599,N_16945,N_19211);
or UO_600 (O_600,N_16449,N_18442);
or UO_601 (O_601,N_16798,N_17130);
and UO_602 (O_602,N_17048,N_18356);
nor UO_603 (O_603,N_19131,N_18578);
xnor UO_604 (O_604,N_19737,N_18629);
and UO_605 (O_605,N_17539,N_16091);
or UO_606 (O_606,N_19940,N_17699);
nand UO_607 (O_607,N_19339,N_16566);
or UO_608 (O_608,N_17432,N_18436);
and UO_609 (O_609,N_18224,N_16154);
and UO_610 (O_610,N_17436,N_16849);
and UO_611 (O_611,N_18925,N_19774);
nor UO_612 (O_612,N_16782,N_18429);
nand UO_613 (O_613,N_16514,N_17869);
nor UO_614 (O_614,N_17784,N_18460);
and UO_615 (O_615,N_19679,N_16030);
xor UO_616 (O_616,N_17645,N_16645);
nand UO_617 (O_617,N_17833,N_19169);
and UO_618 (O_618,N_16850,N_19421);
nor UO_619 (O_619,N_16523,N_18095);
nor UO_620 (O_620,N_19602,N_18903);
xor UO_621 (O_621,N_16435,N_16503);
nand UO_622 (O_622,N_18748,N_16002);
and UO_623 (O_623,N_16552,N_18913);
and UO_624 (O_624,N_16802,N_18656);
nor UO_625 (O_625,N_18091,N_16972);
and UO_626 (O_626,N_17813,N_19514);
and UO_627 (O_627,N_16126,N_19261);
nor UO_628 (O_628,N_18139,N_18417);
nand UO_629 (O_629,N_19955,N_16696);
and UO_630 (O_630,N_16038,N_17568);
or UO_631 (O_631,N_18152,N_19283);
nand UO_632 (O_632,N_19061,N_19512);
nand UO_633 (O_633,N_17237,N_16512);
or UO_634 (O_634,N_17698,N_16133);
nor UO_635 (O_635,N_18855,N_19534);
xnor UO_636 (O_636,N_17441,N_17073);
nor UO_637 (O_637,N_16233,N_18810);
nor UO_638 (O_638,N_17234,N_18462);
or UO_639 (O_639,N_17257,N_17375);
xnor UO_640 (O_640,N_16294,N_18813);
xor UO_641 (O_641,N_19821,N_19011);
xnor UO_642 (O_642,N_18272,N_17595);
or UO_643 (O_643,N_16930,N_17534);
xnor UO_644 (O_644,N_18453,N_18000);
xnor UO_645 (O_645,N_19082,N_16795);
and UO_646 (O_646,N_16698,N_18542);
nand UO_647 (O_647,N_17090,N_16781);
and UO_648 (O_648,N_19236,N_16193);
nor UO_649 (O_649,N_16239,N_17659);
or UO_650 (O_650,N_17822,N_19882);
or UO_651 (O_651,N_18835,N_17424);
and UO_652 (O_652,N_18131,N_16482);
nand UO_653 (O_653,N_17230,N_18926);
xnor UO_654 (O_654,N_16313,N_18670);
and UO_655 (O_655,N_16946,N_18975);
and UO_656 (O_656,N_17609,N_17986);
or UO_657 (O_657,N_18496,N_18609);
or UO_658 (O_658,N_16108,N_19561);
nor UO_659 (O_659,N_18509,N_16427);
xnor UO_660 (O_660,N_17773,N_16379);
nand UO_661 (O_661,N_16466,N_18982);
nand UO_662 (O_662,N_17216,N_17037);
nor UO_663 (O_663,N_17943,N_19041);
nor UO_664 (O_664,N_19178,N_16170);
xnor UO_665 (O_665,N_16003,N_17255);
and UO_666 (O_666,N_18263,N_17949);
and UO_667 (O_667,N_16130,N_19450);
xor UO_668 (O_668,N_19511,N_19255);
and UO_669 (O_669,N_17924,N_16542);
and UO_670 (O_670,N_16028,N_19220);
or UO_671 (O_671,N_16019,N_17570);
xnor UO_672 (O_672,N_19776,N_16886);
nand UO_673 (O_673,N_17616,N_19364);
nor UO_674 (O_674,N_18919,N_18908);
nand UO_675 (O_675,N_17768,N_16533);
xnor UO_676 (O_676,N_18927,N_18015);
nor UO_677 (O_677,N_16223,N_17704);
nand UO_678 (O_678,N_16817,N_19734);
nor UO_679 (O_679,N_19956,N_19231);
and UO_680 (O_680,N_17127,N_17877);
nor UO_681 (O_681,N_17541,N_18316);
nor UO_682 (O_682,N_18093,N_19948);
nand UO_683 (O_683,N_19887,N_18269);
nor UO_684 (O_684,N_17158,N_19968);
xnor UO_685 (O_685,N_17578,N_19404);
nand UO_686 (O_686,N_16113,N_16583);
nand UO_687 (O_687,N_19047,N_17756);
nor UO_688 (O_688,N_16134,N_18797);
nor UO_689 (O_689,N_19949,N_19052);
nand UO_690 (O_690,N_16198,N_16329);
nor UO_691 (O_691,N_19603,N_17778);
nand UO_692 (O_692,N_18840,N_18274);
nor UO_693 (O_693,N_19753,N_19877);
xor UO_694 (O_694,N_17678,N_17573);
nor UO_695 (O_695,N_19176,N_18237);
nor UO_696 (O_696,N_16609,N_18367);
or UO_697 (O_697,N_18989,N_17716);
and UO_698 (O_698,N_16237,N_17850);
xor UO_699 (O_699,N_17239,N_18327);
or UO_700 (O_700,N_16742,N_19750);
and UO_701 (O_701,N_19791,N_17638);
nand UO_702 (O_702,N_18839,N_16591);
and UO_703 (O_703,N_18505,N_17718);
nand UO_704 (O_704,N_18648,N_16189);
and UO_705 (O_705,N_16984,N_16263);
and UO_706 (O_706,N_19430,N_16711);
or UO_707 (O_707,N_18430,N_16231);
nor UO_708 (O_708,N_18256,N_18458);
and UO_709 (O_709,N_19494,N_18432);
and UO_710 (O_710,N_16027,N_16926);
nand UO_711 (O_711,N_16241,N_17207);
xnor UO_712 (O_712,N_17275,N_19062);
nand UO_713 (O_713,N_17022,N_19112);
nand UO_714 (O_714,N_17469,N_18738);
or UO_715 (O_715,N_19976,N_18437);
and UO_716 (O_716,N_19352,N_18446);
and UO_717 (O_717,N_19930,N_19046);
nor UO_718 (O_718,N_18064,N_19874);
xor UO_719 (O_719,N_18633,N_18665);
nor UO_720 (O_720,N_17070,N_19544);
or UO_721 (O_721,N_16143,N_18492);
and UO_722 (O_722,N_16856,N_16595);
or UO_723 (O_723,N_19548,N_19525);
xnor UO_724 (O_724,N_19230,N_19056);
xnor UO_725 (O_725,N_16547,N_17446);
or UO_726 (O_726,N_16011,N_16977);
nand UO_727 (O_727,N_19624,N_18408);
or UO_728 (O_728,N_16592,N_17666);
nor UO_729 (O_729,N_17045,N_16999);
and UO_730 (O_730,N_16169,N_16155);
nand UO_731 (O_731,N_18716,N_16895);
xnor UO_732 (O_732,N_19744,N_17764);
nor UO_733 (O_733,N_17029,N_17102);
or UO_734 (O_734,N_17796,N_17486);
xnor UO_735 (O_735,N_17015,N_19626);
xor UO_736 (O_736,N_18023,N_19729);
and UO_737 (O_737,N_18482,N_18905);
or UO_738 (O_738,N_17639,N_17517);
nand UO_739 (O_739,N_19944,N_17998);
and UO_740 (O_740,N_17931,N_19218);
xor UO_741 (O_741,N_18314,N_18287);
nor UO_742 (O_742,N_19282,N_16703);
and UO_743 (O_743,N_19075,N_19483);
or UO_744 (O_744,N_17934,N_19995);
or UO_745 (O_745,N_19865,N_16183);
xor UO_746 (O_746,N_18977,N_19489);
nor UO_747 (O_747,N_19143,N_18841);
or UO_748 (O_748,N_16888,N_19957);
and UO_749 (O_749,N_18465,N_18085);
and UO_750 (O_750,N_17509,N_17050);
or UO_751 (O_751,N_16043,N_18284);
xor UO_752 (O_752,N_16253,N_17744);
nand UO_753 (O_753,N_17209,N_16714);
or UO_754 (O_754,N_16138,N_16060);
nand UO_755 (O_755,N_16588,N_18844);
nor UO_756 (O_756,N_17788,N_19781);
and UO_757 (O_757,N_16594,N_19014);
nand UO_758 (O_758,N_16528,N_18524);
nand UO_759 (O_759,N_18893,N_16083);
xnor UO_760 (O_760,N_17247,N_16367);
nand UO_761 (O_761,N_18889,N_16436);
nor UO_762 (O_762,N_19910,N_16167);
and UO_763 (O_763,N_17345,N_18549);
nand UO_764 (O_764,N_16878,N_18570);
nor UO_765 (O_765,N_16179,N_16501);
xor UO_766 (O_766,N_19834,N_18022);
and UO_767 (O_767,N_18638,N_18148);
or UO_768 (O_768,N_19633,N_19097);
nor UO_769 (O_769,N_16600,N_19366);
nand UO_770 (O_770,N_18769,N_18451);
and UO_771 (O_771,N_19912,N_19444);
nor UO_772 (O_772,N_17191,N_19493);
nor UO_773 (O_773,N_17708,N_19936);
or UO_774 (O_774,N_16502,N_19329);
nand UO_775 (O_775,N_19363,N_19991);
and UO_776 (O_776,N_18359,N_19773);
nand UO_777 (O_777,N_19686,N_19634);
nand UO_778 (O_778,N_18137,N_16881);
nand UO_779 (O_779,N_17605,N_18682);
nor UO_780 (O_780,N_18684,N_18705);
or UO_781 (O_781,N_18395,N_19900);
and UO_782 (O_782,N_17772,N_17767);
nand UO_783 (O_783,N_19170,N_19890);
nand UO_784 (O_784,N_19436,N_17641);
nand UO_785 (O_785,N_17475,N_16107);
xor UO_786 (O_786,N_18050,N_18177);
or UO_787 (O_787,N_18082,N_17366);
and UO_788 (O_788,N_18901,N_18175);
and UO_789 (O_789,N_19303,N_16172);
nor UO_790 (O_790,N_19156,N_19373);
or UO_791 (O_791,N_17128,N_17072);
and UO_792 (O_792,N_18188,N_18739);
nor UO_793 (O_793,N_17947,N_17025);
or UO_794 (O_794,N_18378,N_19486);
nand UO_795 (O_795,N_16970,N_18605);
xor UO_796 (O_796,N_16046,N_19621);
nor UO_797 (O_797,N_18621,N_18619);
or UO_798 (O_798,N_19831,N_17268);
nand UO_799 (O_799,N_19706,N_18325);
and UO_800 (O_800,N_19616,N_16653);
or UO_801 (O_801,N_17208,N_17166);
or UO_802 (O_802,N_17611,N_19880);
or UO_803 (O_803,N_18782,N_16326);
xnor UO_804 (O_804,N_19028,N_18940);
nand UO_805 (O_805,N_18533,N_19216);
and UO_806 (O_806,N_18702,N_17093);
nor UO_807 (O_807,N_18279,N_17115);
nor UO_808 (O_808,N_17713,N_18213);
nor UO_809 (O_809,N_17780,N_18514);
or UO_810 (O_810,N_19492,N_19974);
and UO_811 (O_811,N_17983,N_19959);
nor UO_812 (O_812,N_19434,N_18986);
nor UO_813 (O_813,N_18503,N_19067);
and UO_814 (O_814,N_17675,N_19674);
and UO_815 (O_815,N_19809,N_19051);
or UO_816 (O_816,N_18757,N_16985);
and UO_817 (O_817,N_19822,N_18744);
nand UO_818 (O_818,N_18295,N_16489);
xor UO_819 (O_819,N_19382,N_19063);
or UO_820 (O_820,N_18692,N_16796);
and UO_821 (O_821,N_19175,N_18838);
nor UO_822 (O_822,N_18190,N_16045);
xor UO_823 (O_823,N_18979,N_18149);
nor UO_824 (O_824,N_16283,N_19272);
nor UO_825 (O_825,N_16344,N_17265);
and UO_826 (O_826,N_16117,N_19515);
nor UO_827 (O_827,N_18275,N_17136);
or UO_828 (O_828,N_17786,N_19977);
or UO_829 (O_829,N_16531,N_19712);
nand UO_830 (O_830,N_17125,N_19907);
nor UO_831 (O_831,N_18448,N_18345);
and UO_832 (O_832,N_18302,N_18231);
and UO_833 (O_833,N_16339,N_16175);
xor UO_834 (O_834,N_19735,N_16707);
nand UO_835 (O_835,N_18634,N_16354);
xnor UO_836 (O_836,N_16799,N_18126);
or UO_837 (O_837,N_16776,N_19553);
and UO_838 (O_838,N_19077,N_16613);
nor UO_839 (O_839,N_19367,N_16590);
and UO_840 (O_840,N_16267,N_16220);
nor UO_841 (O_841,N_18529,N_17120);
and UO_842 (O_842,N_17302,N_16907);
nand UO_843 (O_843,N_17725,N_19518);
and UO_844 (O_844,N_17250,N_17101);
xnor UO_845 (O_845,N_18713,N_17624);
and UO_846 (O_846,N_16025,N_19513);
nand UO_847 (O_847,N_19699,N_17145);
nor UO_848 (O_848,N_19316,N_18456);
nor UO_849 (O_849,N_16777,N_18394);
nand UO_850 (O_850,N_16676,N_18267);
and UO_851 (O_851,N_19472,N_19305);
and UO_852 (O_852,N_18298,N_16914);
and UO_853 (O_853,N_17324,N_16480);
nand UO_854 (O_854,N_17766,N_19970);
nor UO_855 (O_855,N_18740,N_19012);
or UO_856 (O_856,N_19101,N_18625);
or UO_857 (O_857,N_16690,N_16560);
nor UO_858 (O_858,N_16450,N_18034);
nor UO_859 (O_859,N_17243,N_18029);
nor UO_860 (O_860,N_16068,N_16278);
nor UO_861 (O_861,N_17576,N_18885);
and UO_862 (O_862,N_17742,N_18681);
nor UO_863 (O_863,N_19114,N_18192);
nor UO_864 (O_864,N_17225,N_19048);
xor UO_865 (O_865,N_17317,N_18096);
nand UO_866 (O_866,N_19872,N_17991);
xnor UO_867 (O_867,N_18896,N_16292);
or UO_868 (O_868,N_19696,N_17596);
xor UO_869 (O_869,N_17162,N_19142);
xor UO_870 (O_870,N_19861,N_16180);
xnor UO_871 (O_871,N_17445,N_18485);
or UO_872 (O_872,N_18697,N_18644);
and UO_873 (O_873,N_17069,N_17182);
and UO_874 (O_874,N_19157,N_19826);
xor UO_875 (O_875,N_19396,N_18059);
and UO_876 (O_876,N_16148,N_16327);
or UO_877 (O_877,N_16336,N_18771);
xnor UO_878 (O_878,N_17751,N_18171);
nor UO_879 (O_879,N_17847,N_18836);
and UO_880 (O_880,N_17738,N_18164);
nor UO_881 (O_881,N_19249,N_16141);
nand UO_882 (O_882,N_17583,N_18817);
and UO_883 (O_883,N_19710,N_18712);
xor UO_884 (O_884,N_17088,N_19286);
xnor UO_885 (O_885,N_19784,N_18591);
nand UO_886 (O_886,N_16953,N_18875);
or UO_887 (O_887,N_17231,N_18323);
and UO_888 (O_888,N_17560,N_16406);
nor UO_889 (O_889,N_18639,N_17410);
nand UO_890 (O_890,N_17672,N_18837);
nand UO_891 (O_891,N_19203,N_16457);
xor UO_892 (O_892,N_19669,N_17078);
nand UO_893 (O_893,N_18557,N_17531);
nand UO_894 (O_894,N_19507,N_18938);
and UO_895 (O_895,N_17804,N_18127);
or UO_896 (O_896,N_17470,N_17131);
nor UO_897 (O_897,N_16730,N_17750);
xnor UO_898 (O_898,N_18319,N_17056);
or UO_899 (O_899,N_18169,N_16293);
xor UO_900 (O_900,N_17820,N_19122);
nand UO_901 (O_901,N_17680,N_18830);
xnor UO_902 (O_902,N_17404,N_19005);
nor UO_903 (O_903,N_18737,N_18372);
nor UO_904 (O_904,N_16244,N_19301);
nor UO_905 (O_905,N_18689,N_19663);
xor UO_906 (O_906,N_19470,N_17109);
xnor UO_907 (O_907,N_19707,N_17292);
and UO_908 (O_908,N_16979,N_19452);
xor UO_909 (O_909,N_18236,N_19760);
xnor UO_910 (O_910,N_18051,N_17267);
xor UO_911 (O_911,N_17018,N_16033);
nor UO_912 (O_912,N_19264,N_16978);
nor UO_913 (O_913,N_19925,N_17953);
and UO_914 (O_914,N_19177,N_16593);
xnor UO_915 (O_915,N_16829,N_19840);
and UO_916 (O_916,N_17313,N_18831);
nor UO_917 (O_917,N_17122,N_18403);
and UO_918 (O_918,N_19250,N_17957);
or UO_919 (O_919,N_16059,N_17592);
nand UO_920 (O_920,N_16626,N_19814);
nor UO_921 (O_921,N_19579,N_19906);
and UO_922 (O_922,N_17180,N_17522);
or UO_923 (O_923,N_19208,N_16385);
nor UO_924 (O_924,N_19501,N_16847);
and UO_925 (O_925,N_19000,N_19743);
or UO_926 (O_926,N_18718,N_16416);
and UO_927 (O_927,N_16872,N_17456);
xnor UO_928 (O_928,N_17202,N_19628);
nand UO_929 (O_929,N_19820,N_17707);
nand UO_930 (O_930,N_18398,N_16670);
xnor UO_931 (O_931,N_18821,N_16284);
nor UO_932 (O_932,N_16663,N_16383);
and UO_933 (O_933,N_18929,N_16275);
or UO_934 (O_934,N_16903,N_19454);
nand UO_935 (O_935,N_17124,N_19636);
and UO_936 (O_936,N_16736,N_17887);
and UO_937 (O_937,N_17779,N_17017);
and UO_938 (O_938,N_18701,N_16303);
nor UO_939 (O_939,N_18805,N_19667);
xnor UO_940 (O_940,N_19867,N_17821);
or UO_941 (O_941,N_16101,N_16110);
nor UO_942 (O_942,N_18562,N_17240);
or UO_943 (O_943,N_19551,N_19420);
nor UO_944 (O_944,N_19361,N_19538);
or UO_945 (O_945,N_16994,N_16647);
or UO_946 (O_946,N_17155,N_16251);
nand UO_947 (O_947,N_19642,N_16135);
or UO_948 (O_948,N_18443,N_17640);
and UO_949 (O_949,N_19200,N_16014);
nor UO_950 (O_950,N_18454,N_16589);
and UO_951 (O_951,N_19324,N_16828);
xor UO_952 (O_952,N_16281,N_18891);
nand UO_953 (O_953,N_17482,N_18140);
and UO_954 (O_954,N_16465,N_18435);
and UO_955 (O_955,N_16616,N_18170);
nand UO_956 (O_956,N_19081,N_16990);
nand UO_957 (O_957,N_19680,N_18217);
xnor UO_958 (O_958,N_19117,N_18368);
nand UO_959 (O_959,N_16312,N_17289);
and UO_960 (O_960,N_19913,N_19786);
nand UO_961 (O_961,N_16931,N_18262);
nor UO_962 (O_962,N_19619,N_17028);
nand UO_963 (O_963,N_16104,N_17524);
xnor UO_964 (O_964,N_16297,N_16218);
and UO_965 (O_965,N_16368,N_18604);
and UO_966 (O_966,N_18226,N_16980);
and UO_967 (O_967,N_17186,N_17585);
and UO_968 (O_968,N_17135,N_16601);
or UO_969 (O_969,N_16200,N_16640);
nand UO_970 (O_970,N_18969,N_16342);
or UO_971 (O_971,N_16748,N_18972);
nand UO_972 (O_972,N_16635,N_17643);
xor UO_973 (O_973,N_17538,N_19503);
nor UO_974 (O_974,N_16610,N_17876);
nand UO_975 (O_975,N_18488,N_19225);
xnor UO_976 (O_976,N_17898,N_16429);
and UO_977 (O_977,N_16662,N_16274);
or UO_978 (O_978,N_17423,N_18081);
or UO_979 (O_979,N_19330,N_16470);
or UO_980 (O_980,N_16667,N_19488);
or UO_981 (O_981,N_18704,N_17063);
nand UO_982 (O_982,N_18764,N_18335);
or UO_983 (O_983,N_19271,N_17903);
xnor UO_984 (O_984,N_16556,N_16390);
nor UO_985 (O_985,N_16105,N_17527);
nand UO_986 (O_986,N_16199,N_19254);
nor UO_987 (O_987,N_16859,N_16664);
and UO_988 (O_988,N_17684,N_18075);
nand UO_989 (O_989,N_16510,N_17642);
nand UO_990 (O_990,N_16694,N_18401);
xnor UO_991 (O_991,N_17218,N_17040);
or UO_992 (O_992,N_17097,N_16484);
nor UO_993 (O_993,N_16201,N_19406);
and UO_994 (O_994,N_19410,N_18332);
and UO_995 (O_995,N_18950,N_17331);
xor UO_996 (O_996,N_16998,N_19093);
nand UO_997 (O_997,N_17291,N_16115);
nor UO_998 (O_998,N_19289,N_16195);
nor UO_999 (O_999,N_19745,N_18472);
or UO_1000 (O_1000,N_18881,N_17205);
nand UO_1001 (O_1001,N_17598,N_18113);
and UO_1002 (O_1002,N_17485,N_17365);
xor UO_1003 (O_1003,N_17965,N_19287);
or UO_1004 (O_1004,N_18427,N_19248);
and UO_1005 (O_1005,N_19427,N_18657);
xnor UO_1006 (O_1006,N_18215,N_19100);
xor UO_1007 (O_1007,N_18249,N_18115);
xor UO_1008 (O_1008,N_19388,N_17392);
nor UO_1009 (O_1009,N_18544,N_17233);
nand UO_1010 (O_1010,N_17993,N_18357);
or UO_1011 (O_1011,N_16160,N_19635);
nor UO_1012 (O_1012,N_17157,N_19070);
and UO_1013 (O_1013,N_18551,N_17625);
xnor UO_1014 (O_1014,N_19675,N_16764);
or UO_1015 (O_1015,N_16087,N_19409);
or UO_1016 (O_1016,N_18690,N_18122);
nand UO_1017 (O_1017,N_18842,N_16683);
and UO_1018 (O_1018,N_18663,N_19726);
or UO_1019 (O_1019,N_19022,N_18014);
nand UO_1020 (O_1020,N_18343,N_18779);
and UO_1021 (O_1021,N_17477,N_19468);
or UO_1022 (O_1022,N_16515,N_17187);
nand UO_1023 (O_1023,N_18497,N_17895);
or UO_1024 (O_1024,N_18160,N_18776);
or UO_1025 (O_1025,N_17052,N_19091);
nor UO_1026 (O_1026,N_18862,N_16665);
xor UO_1027 (O_1027,N_18253,N_16811);
nand UO_1028 (O_1028,N_19719,N_17341);
and UO_1029 (O_1029,N_17557,N_19573);
and UO_1030 (O_1030,N_18389,N_18067);
nor UO_1031 (O_1031,N_18311,N_19761);
and UO_1032 (O_1032,N_16194,N_16227);
and UO_1033 (O_1033,N_16479,N_19130);
or UO_1034 (O_1034,N_16355,N_18413);
nand UO_1035 (O_1035,N_18346,N_16561);
nand UO_1036 (O_1036,N_19148,N_18232);
or UO_1037 (O_1037,N_17159,N_17823);
nor UO_1038 (O_1038,N_19904,N_16774);
nand UO_1039 (O_1039,N_16867,N_16266);
and UO_1040 (O_1040,N_17880,N_18397);
or UO_1041 (O_1041,N_19747,N_17442);
nor UO_1042 (O_1042,N_19917,N_17612);
xnor UO_1043 (O_1043,N_17153,N_17938);
xor UO_1044 (O_1044,N_17183,N_19947);
and UO_1045 (O_1045,N_16638,N_16004);
xor UO_1046 (O_1046,N_16410,N_18358);
xor UO_1047 (O_1047,N_16432,N_17959);
or UO_1048 (O_1048,N_17184,N_17284);
or UO_1049 (O_1049,N_18878,N_16085);
xnor UO_1050 (O_1050,N_18399,N_16522);
xnor UO_1051 (O_1051,N_18948,N_16102);
or UO_1052 (O_1052,N_19671,N_19759);
or UO_1053 (O_1053,N_17161,N_18277);
nand UO_1054 (O_1054,N_19522,N_19405);
and UO_1055 (O_1055,N_18406,N_18962);
nand UO_1056 (O_1056,N_16969,N_18532);
nand UO_1057 (O_1057,N_16623,N_19818);
nand UO_1058 (O_1058,N_16403,N_19478);
and UO_1059 (O_1059,N_16769,N_19351);
and UO_1060 (O_1060,N_17932,N_18765);
and UO_1061 (O_1061,N_16909,N_19298);
and UO_1062 (O_1062,N_16376,N_17227);
xnor UO_1063 (O_1063,N_18791,N_19722);
and UO_1064 (O_1064,N_16715,N_18507);
xor UO_1065 (O_1065,N_19376,N_19362);
and UO_1066 (O_1066,N_17803,N_19104);
or UO_1067 (O_1067,N_16554,N_18150);
nor UO_1068 (O_1068,N_17384,N_17914);
and UO_1069 (O_1069,N_19990,N_18300);
xnor UO_1070 (O_1070,N_19853,N_19238);
nand UO_1071 (O_1071,N_19643,N_19466);
nand UO_1072 (O_1072,N_18035,N_17523);
and UO_1073 (O_1073,N_16474,N_18286);
or UO_1074 (O_1074,N_16395,N_17244);
and UO_1075 (O_1075,N_19560,N_19851);
xnor UO_1076 (O_1076,N_17706,N_19615);
nand UO_1077 (O_1077,N_18669,N_19035);
nor UO_1078 (O_1078,N_16137,N_16789);
or UO_1079 (O_1079,N_16812,N_17253);
or UO_1080 (O_1080,N_16743,N_18564);
xor UO_1081 (O_1081,N_17347,N_19746);
nand UO_1082 (O_1082,N_18066,N_19666);
nor UO_1083 (O_1083,N_18352,N_18766);
nor UO_1084 (O_1084,N_16751,N_16546);
or UO_1085 (O_1085,N_19240,N_19985);
nor UO_1086 (O_1086,N_18971,N_19788);
nor UO_1087 (O_1087,N_16908,N_17582);
or UO_1088 (O_1088,N_16356,N_16153);
xnor UO_1089 (O_1089,N_17518,N_18247);
or UO_1090 (O_1090,N_18270,N_18381);
or UO_1091 (O_1091,N_18048,N_18741);
nand UO_1092 (O_1092,N_19983,N_16360);
nand UO_1093 (O_1093,N_16538,N_19196);
nor UO_1094 (O_1094,N_17647,N_19358);
xnor UO_1095 (O_1095,N_17739,N_16562);
nand UO_1096 (O_1096,N_19945,N_18501);
xor UO_1097 (O_1097,N_16139,N_18006);
or UO_1098 (O_1098,N_18129,N_17886);
nand UO_1099 (O_1099,N_18219,N_16704);
and UO_1100 (O_1100,N_18535,N_16900);
and UO_1101 (O_1101,N_19721,N_16488);
xor UO_1102 (O_1102,N_17628,N_19789);
and UO_1103 (O_1103,N_18653,N_18119);
xor UO_1104 (O_1104,N_16890,N_17878);
or UO_1105 (O_1105,N_16399,N_18291);
xnor UO_1106 (O_1106,N_19584,N_16520);
nand UO_1107 (O_1107,N_16633,N_16762);
and UO_1108 (O_1108,N_19610,N_17132);
nor UO_1109 (O_1109,N_18884,N_18489);
nand UO_1110 (O_1110,N_17263,N_18735);
xor UO_1111 (O_1111,N_16333,N_18958);
nor UO_1112 (O_1112,N_17220,N_18832);
nor UO_1113 (O_1113,N_17219,N_17575);
nand UO_1114 (O_1114,N_16114,N_18240);
xnor UO_1115 (O_1115,N_16723,N_16954);
and UO_1116 (O_1116,N_16722,N_19979);
or UO_1117 (O_1117,N_17262,N_16078);
nand UO_1118 (O_1118,N_17306,N_19018);
or UO_1119 (O_1119,N_17894,N_17460);
xnor UO_1120 (O_1120,N_16306,N_19425);
xnor UO_1121 (O_1121,N_16317,N_18180);
nand UO_1122 (O_1122,N_18110,N_17062);
or UO_1123 (O_1123,N_19260,N_18114);
nand UO_1124 (O_1124,N_17819,N_18590);
nor UO_1125 (O_1125,N_17782,N_18602);
or UO_1126 (O_1126,N_18490,N_19660);
xor UO_1127 (O_1127,N_18310,N_19295);
xor UO_1128 (O_1128,N_16490,N_16960);
or UO_1129 (O_1129,N_17360,N_17368);
or UO_1130 (O_1130,N_17586,N_18751);
nand UO_1131 (O_1131,N_19690,N_16516);
nand UO_1132 (O_1132,N_16768,N_16208);
nor UO_1133 (O_1133,N_19587,N_19832);
nor UO_1134 (O_1134,N_16735,N_19399);
or UO_1135 (O_1135,N_16689,N_17814);
and UO_1136 (O_1136,N_17920,N_18915);
or UO_1137 (O_1137,N_17272,N_17449);
xor UO_1138 (O_1138,N_18382,N_17505);
and UO_1139 (O_1139,N_16851,N_16780);
or UO_1140 (O_1140,N_19811,N_17496);
xnor UO_1141 (O_1141,N_16472,N_16446);
or UO_1142 (O_1142,N_17892,N_16842);
nand UO_1143 (O_1143,N_17011,N_18032);
nor UO_1144 (O_1144,N_19736,N_17197);
or UO_1145 (O_1145,N_16464,N_19096);
nor UO_1146 (O_1146,N_17476,N_18729);
or UO_1147 (O_1147,N_19664,N_16430);
or UO_1148 (O_1148,N_16058,N_18727);
nand UO_1149 (O_1149,N_18473,N_17147);
or UO_1150 (O_1150,N_17406,N_19802);
and UO_1151 (O_1151,N_19102,N_19445);
and UO_1152 (O_1152,N_18043,N_18222);
and UO_1153 (O_1153,N_16156,N_19477);
and UO_1154 (O_1154,N_17712,N_17483);
nand UO_1155 (O_1155,N_16389,N_18613);
or UO_1156 (O_1156,N_17413,N_19899);
nand UO_1157 (O_1157,N_18083,N_16190);
xor UO_1158 (O_1158,N_19118,N_17085);
and UO_1159 (O_1159,N_18133,N_19768);
nor UO_1160 (O_1160,N_17479,N_16838);
xor UO_1161 (O_1161,N_16923,N_17172);
and UO_1162 (O_1162,N_16226,N_19115);
or UO_1163 (O_1163,N_18184,N_17422);
xnor UO_1164 (O_1164,N_17113,N_17720);
nor UO_1165 (O_1165,N_19258,N_18943);
nor UO_1166 (O_1166,N_18426,N_16513);
nor UO_1167 (O_1167,N_19244,N_19748);
and UO_1168 (O_1168,N_18643,N_16614);
xnor UO_1169 (O_1169,N_18550,N_19571);
nand UO_1170 (O_1170,N_16072,N_17035);
and UO_1171 (O_1171,N_19897,N_18555);
and UO_1172 (O_1172,N_19689,N_17414);
nor UO_1173 (O_1173,N_19918,N_17809);
xnor UO_1174 (O_1174,N_16987,N_19502);
nor UO_1175 (O_1175,N_17118,N_17670);
nand UO_1176 (O_1176,N_16618,N_17864);
or UO_1177 (O_1177,N_17851,N_16094);
or UO_1178 (O_1178,N_17649,N_19407);
and UO_1179 (O_1179,N_16823,N_18495);
nor UO_1180 (O_1180,N_19138,N_18477);
or UO_1181 (O_1181,N_19487,N_18575);
nor UO_1182 (O_1182,N_16896,N_16348);
xor UO_1183 (O_1183,N_17086,N_16797);
or UO_1184 (O_1184,N_19992,N_17312);
and UO_1185 (O_1185,N_19875,N_16679);
xor UO_1186 (O_1186,N_18980,N_18007);
nor UO_1187 (O_1187,N_16447,N_17513);
nand UO_1188 (O_1188,N_17849,N_18363);
nand UO_1189 (O_1189,N_17065,N_19849);
nor UO_1190 (O_1190,N_18733,N_16109);
nor UO_1191 (O_1191,N_17334,N_19596);
xor UO_1192 (O_1192,N_16377,N_17997);
xor UO_1193 (O_1193,N_16651,N_17462);
and UO_1194 (O_1194,N_19150,N_19467);
nand UO_1195 (O_1195,N_19543,N_19614);
nor UO_1196 (O_1196,N_18033,N_19517);
xor UO_1197 (O_1197,N_18804,N_18135);
and UO_1198 (O_1198,N_17691,N_18181);
or UO_1199 (O_1199,N_17771,N_18312);
nand UO_1200 (O_1200,N_17917,N_19443);
and UO_1201 (O_1201,N_19839,N_19372);
xor UO_1202 (O_1202,N_16731,N_17430);
and UO_1203 (O_1203,N_16044,N_16282);
nand UO_1204 (O_1204,N_16016,N_19293);
or UO_1205 (O_1205,N_17885,N_17776);
or UO_1206 (O_1206,N_16086,N_18418);
nand UO_1207 (O_1207,N_19437,N_17866);
and UO_1208 (O_1208,N_17963,N_17385);
nor UO_1209 (O_1209,N_18900,N_17714);
xor UO_1210 (O_1210,N_17464,N_19915);
or UO_1211 (O_1211,N_16096,N_18199);
nor UO_1212 (O_1212,N_17100,N_16462);
nand UO_1213 (O_1213,N_16437,N_18018);
nand UO_1214 (O_1214,N_18597,N_19036);
xor UO_1215 (O_1215,N_19090,N_17511);
or UO_1216 (O_1216,N_16499,N_19016);
and UO_1217 (O_1217,N_19996,N_19334);
or UO_1218 (O_1218,N_18646,N_19606);
nand UO_1219 (O_1219,N_17148,N_19535);
xnor UO_1220 (O_1220,N_19799,N_16487);
or UO_1221 (O_1221,N_18536,N_19206);
nand UO_1222 (O_1222,N_16320,N_18370);
or UO_1223 (O_1223,N_17907,N_18143);
or UO_1224 (O_1224,N_18974,N_17146);
nand UO_1225 (O_1225,N_18157,N_18273);
nand UO_1226 (O_1226,N_19276,N_19723);
and UO_1227 (O_1227,N_19210,N_19625);
nor UO_1228 (O_1228,N_17427,N_16378);
nand UO_1229 (O_1229,N_18305,N_18799);
nor UO_1230 (O_1230,N_17489,N_18155);
nand UO_1231 (O_1231,N_18664,N_19989);
xor UO_1232 (O_1232,N_19591,N_19291);
or UO_1233 (O_1233,N_19181,N_17068);
nand UO_1234 (O_1234,N_17697,N_17855);
nor UO_1235 (O_1235,N_17743,N_16202);
nand UO_1236 (O_1236,N_18416,N_18539);
nor UO_1237 (O_1237,N_19498,N_19227);
nor UO_1238 (O_1238,N_17296,N_17835);
nand UO_1239 (O_1239,N_17490,N_19006);
nor UO_1240 (O_1240,N_19876,N_19234);
and UO_1241 (O_1241,N_19775,N_18534);
or UO_1242 (O_1242,N_17955,N_18173);
and UO_1243 (O_1243,N_17095,N_18383);
nand UO_1244 (O_1244,N_16371,N_17336);
xnor UO_1245 (O_1245,N_16280,N_17994);
and UO_1246 (O_1246,N_19647,N_16964);
nand UO_1247 (O_1247,N_18863,N_19779);
nand UO_1248 (O_1248,N_16392,N_19733);
xnor UO_1249 (O_1249,N_17245,N_17839);
or UO_1250 (O_1250,N_19460,N_19854);
and UO_1251 (O_1251,N_17361,N_19354);
nor UO_1252 (O_1252,N_16454,N_18024);
xnor UO_1253 (O_1253,N_18850,N_16131);
nand UO_1254 (O_1254,N_18787,N_19607);
xor UO_1255 (O_1255,N_16962,N_17179);
nor UO_1256 (O_1256,N_17043,N_19426);
xor UO_1257 (O_1257,N_16913,N_18308);
nor UO_1258 (O_1258,N_16884,N_17581);
nor UO_1259 (O_1259,N_19997,N_17286);
or UO_1260 (O_1260,N_17382,N_18282);
and UO_1261 (O_1261,N_16459,N_18673);
xor UO_1262 (O_1262,N_17232,N_17929);
and UO_1263 (O_1263,N_17603,N_17921);
xnor UO_1264 (O_1264,N_17499,N_16845);
nor UO_1265 (O_1265,N_17246,N_16644);
and UO_1266 (O_1266,N_18385,N_19246);
xor UO_1267 (O_1267,N_16719,N_19824);
nor UO_1268 (O_1268,N_19812,N_16311);
and UO_1269 (O_1269,N_19687,N_16414);
xnor UO_1270 (O_1270,N_19964,N_16564);
xor UO_1271 (O_1271,N_17966,N_18655);
nand UO_1272 (O_1272,N_17249,N_17661);
or UO_1273 (O_1273,N_17519,N_19958);
nor UO_1274 (O_1274,N_19980,N_18380);
nand UO_1275 (O_1275,N_18142,N_16756);
or UO_1276 (O_1276,N_16268,N_16330);
nand UO_1277 (O_1277,N_18031,N_17944);
nand UO_1278 (O_1278,N_19620,N_18786);
xnor UO_1279 (O_1279,N_18662,N_18030);
or UO_1280 (O_1280,N_16265,N_19171);
and UO_1281 (O_1281,N_19105,N_19153);
or UO_1282 (O_1282,N_17405,N_17502);
or UO_1283 (O_1283,N_16000,N_17459);
xor UO_1284 (O_1284,N_18719,N_19108);
or UO_1285 (O_1285,N_19552,N_17860);
and UO_1286 (O_1286,N_17295,N_18387);
and UO_1287 (O_1287,N_16407,N_16585);
and UO_1288 (O_1288,N_17348,N_16537);
and UO_1289 (O_1289,N_19357,N_18601);
or UO_1290 (O_1290,N_18732,N_16247);
and UO_1291 (O_1291,N_16615,N_17355);
or UO_1292 (O_1292,N_17426,N_19640);
nand UO_1293 (O_1293,N_19288,N_16721);
nand UO_1294 (O_1294,N_16619,N_18561);
nor UO_1295 (O_1295,N_17114,N_18728);
xor UO_1296 (O_1296,N_16767,N_18225);
xnor UO_1297 (O_1297,N_18897,N_18659);
or UO_1298 (O_1298,N_16350,N_16706);
nand UO_1299 (O_1299,N_17308,N_19681);
nor UO_1300 (O_1300,N_19292,N_19147);
or UO_1301 (O_1301,N_18283,N_18246);
or UO_1302 (O_1302,N_16820,N_16982);
or UO_1303 (O_1303,N_19094,N_19668);
and UO_1304 (O_1304,N_19714,N_18833);
or UO_1305 (O_1305,N_19030,N_16166);
nand UO_1306 (O_1306,N_19257,N_18723);
or UO_1307 (O_1307,N_19950,N_18599);
xnor UO_1308 (O_1308,N_19003,N_16760);
or UO_1309 (O_1309,N_16974,N_16423);
nand UO_1310 (O_1310,N_17746,N_18877);
xnor UO_1311 (O_1311,N_18709,N_17251);
and UO_1312 (O_1312,N_18478,N_18021);
xor UO_1313 (O_1313,N_18218,N_17655);
nand UO_1314 (O_1314,N_16587,N_19092);
and UO_1315 (O_1315,N_18261,N_18080);
nor UO_1316 (O_1316,N_16322,N_16021);
nor UO_1317 (O_1317,N_18631,N_19089);
xnor UO_1318 (O_1318,N_17761,N_18880);
and UO_1319 (O_1319,N_17142,N_17506);
nor UO_1320 (O_1320,N_17254,N_16708);
and UO_1321 (O_1321,N_17867,N_19656);
xor UO_1322 (O_1322,N_18686,N_19547);
and UO_1323 (O_1323,N_19162,N_16496);
nor UO_1324 (O_1324,N_19123,N_17935);
nor UO_1325 (O_1325,N_17189,N_18902);
or UO_1326 (O_1326,N_19711,N_19795);
and UO_1327 (O_1327,N_16755,N_18556);
nand UO_1328 (O_1328,N_19338,N_18571);
and UO_1329 (O_1329,N_17622,N_16373);
xor UO_1330 (O_1330,N_19583,N_19461);
xor UO_1331 (O_1331,N_16111,N_17664);
or UO_1332 (O_1332,N_18859,N_16097);
xor UO_1333 (O_1333,N_16219,N_17150);
nand UO_1334 (O_1334,N_16720,N_19343);
or UO_1335 (O_1335,N_19390,N_17500);
xor UO_1336 (O_1336,N_17156,N_18176);
or UO_1337 (O_1337,N_18851,N_17941);
xor UO_1338 (O_1338,N_16191,N_17558);
xnor UO_1339 (O_1339,N_18116,N_18680);
or UO_1340 (O_1340,N_18400,N_16536);
nand UO_1341 (O_1341,N_19801,N_19758);
or UO_1342 (O_1342,N_17173,N_18517);
nand UO_1343 (O_1343,N_16791,N_16445);
or UO_1344 (O_1344,N_18434,N_17421);
and UO_1345 (O_1345,N_19612,N_18244);
or UO_1346 (O_1346,N_18547,N_18852);
nor UO_1347 (O_1347,N_17089,N_19941);
and UO_1348 (O_1348,N_17915,N_16433);
and UO_1349 (O_1349,N_17735,N_17379);
and UO_1350 (O_1350,N_16245,N_19479);
and UO_1351 (O_1351,N_16885,N_16015);
or UO_1352 (O_1352,N_16986,N_16478);
xnor UO_1353 (O_1353,N_17217,N_16844);
or UO_1354 (O_1354,N_18956,N_17222);
nand UO_1355 (O_1355,N_17829,N_18106);
nor UO_1356 (O_1356,N_16471,N_16677);
or UO_1357 (O_1357,N_19938,N_16833);
or UO_1358 (O_1358,N_17167,N_17307);
and UO_1359 (O_1359,N_17152,N_19837);
or UO_1360 (O_1360,N_16481,N_16910);
nand UO_1361 (O_1361,N_19973,N_17927);
xnor UO_1362 (O_1362,N_19787,N_17682);
nand UO_1363 (O_1363,N_19256,N_17979);
or UO_1364 (O_1364,N_18044,N_16249);
and UO_1365 (O_1365,N_19935,N_18745);
or UO_1366 (O_1366,N_18338,N_18752);
nand UO_1367 (O_1367,N_17567,N_16452);
nor UO_1368 (O_1368,N_17049,N_17651);
or UO_1369 (O_1369,N_17990,N_17473);
xnor UO_1370 (O_1370,N_17389,N_16309);
and UO_1371 (O_1371,N_19557,N_19205);
and UO_1372 (O_1372,N_18493,N_17077);
nor UO_1373 (O_1373,N_17196,N_18258);
nor UO_1374 (O_1374,N_17465,N_17945);
nor UO_1375 (O_1375,N_16221,N_18976);
nor UO_1376 (O_1376,N_17632,N_17777);
and UO_1377 (O_1377,N_17123,N_19929);
and UO_1378 (O_1378,N_19819,N_17503);
nand UO_1379 (O_1379,N_18208,N_16830);
nand UO_1380 (O_1380,N_19464,N_17501);
xor UO_1381 (O_1381,N_17940,N_17928);
and UO_1382 (O_1382,N_18349,N_19306);
nand UO_1383 (O_1383,N_18717,N_17397);
nor UO_1384 (O_1384,N_16391,N_19574);
nand UO_1385 (O_1385,N_18420,N_17555);
nor UO_1386 (O_1386,N_19328,N_16067);
and UO_1387 (O_1387,N_17198,N_18449);
or UO_1388 (O_1388,N_19207,N_18386);
xnor UO_1389 (O_1389,N_16666,N_19402);
nand UO_1390 (O_1390,N_18626,N_18825);
nand UO_1391 (O_1391,N_17734,N_17300);
and UO_1392 (O_1392,N_19738,N_16081);
nor UO_1393 (O_1393,N_18100,N_19199);
xor UO_1394 (O_1394,N_19684,N_16372);
and UO_1395 (O_1395,N_19349,N_17569);
xnor UO_1396 (O_1396,N_16098,N_18042);
xnor UO_1397 (O_1397,N_17972,N_19593);
xnor UO_1398 (O_1398,N_18892,N_18292);
nand UO_1399 (O_1399,N_17417,N_19135);
and UO_1400 (O_1400,N_19844,N_16261);
xor UO_1401 (O_1401,N_18099,N_17689);
xnor UO_1402 (O_1402,N_16099,N_19064);
xnor UO_1403 (O_1403,N_18445,N_16023);
or UO_1404 (O_1404,N_17549,N_17831);
and UO_1405 (O_1405,N_16958,N_18827);
or UO_1406 (O_1406,N_19752,N_17604);
xnor UO_1407 (O_1407,N_18964,N_16006);
xor UO_1408 (O_1408,N_17562,N_19315);
nor UO_1409 (O_1409,N_17358,N_18802);
xnor UO_1410 (O_1410,N_16270,N_16784);
and UO_1411 (O_1411,N_19700,N_16819);
nor UO_1412 (O_1412,N_18818,N_16989);
nor UO_1413 (O_1413,N_17380,N_18094);
xnor UO_1414 (O_1414,N_16307,N_16176);
and UO_1415 (O_1415,N_17988,N_16413);
nand UO_1416 (O_1416,N_16692,N_19069);
and UO_1417 (O_1417,N_17753,N_17587);
or UO_1418 (O_1418,N_17883,N_18672);
xnor UO_1419 (O_1419,N_18281,N_19377);
or UO_1420 (O_1420,N_19044,N_17563);
xnor UO_1421 (O_1421,N_18978,N_19537);
or UO_1422 (O_1422,N_16788,N_16100);
xor UO_1423 (O_1423,N_16905,N_18117);
or UO_1424 (O_1424,N_19982,N_17346);
xor UO_1425 (O_1425,N_18162,N_16785);
or UO_1426 (O_1426,N_16577,N_19739);
or UO_1427 (O_1427,N_18806,N_17787);
nand UO_1428 (O_1428,N_18017,N_16573);
xor UO_1429 (O_1429,N_19045,N_17055);
and UO_1430 (O_1430,N_18384,N_16380);
nand UO_1431 (O_1431,N_16106,N_17933);
nor UO_1432 (O_1432,N_17607,N_17977);
and UO_1433 (O_1433,N_18097,N_18651);
nor UO_1434 (O_1434,N_19297,N_16262);
or UO_1435 (O_1435,N_16608,N_16825);
xor UO_1436 (O_1436,N_18565,N_19403);
xor UO_1437 (O_1437,N_16761,N_16650);
or UO_1438 (O_1438,N_18968,N_17195);
or UO_1439 (O_1439,N_17340,N_17891);
and UO_1440 (O_1440,N_16771,N_18174);
xnor UO_1441 (O_1441,N_19709,N_18512);
nand UO_1442 (O_1442,N_16259,N_17168);
or UO_1443 (O_1443,N_19870,N_18650);
nor UO_1444 (O_1444,N_16899,N_16185);
xnor UO_1445 (O_1445,N_18179,N_19359);
and UO_1446 (O_1446,N_19590,N_18936);
or UO_1447 (O_1447,N_16671,N_19988);
or UO_1448 (O_1448,N_17104,N_18441);
or UO_1449 (O_1449,N_19180,N_19066);
nor UO_1450 (O_1450,N_17608,N_16402);
and UO_1451 (O_1451,N_16352,N_17752);
and UO_1452 (O_1452,N_18762,N_18959);
xor UO_1453 (O_1453,N_18461,N_19160);
or UO_1454 (O_1454,N_19125,N_17662);
nor UO_1455 (O_1455,N_16300,N_19592);
xnor UO_1456 (O_1456,N_19670,N_17844);
nand UO_1457 (O_1457,N_18136,N_19375);
nand UO_1458 (O_1458,N_16093,N_18326);
and UO_1459 (O_1459,N_17882,N_19500);
nand UO_1460 (O_1460,N_19137,N_16534);
nor UO_1461 (O_1461,N_18185,N_17117);
nor UO_1462 (O_1462,N_19189,N_19219);
and UO_1463 (O_1463,N_17948,N_16127);
xor UO_1464 (O_1464,N_19369,N_18904);
xnor UO_1465 (O_1465,N_19128,N_16152);
nor UO_1466 (O_1466,N_18798,N_16228);
nor UO_1467 (O_1467,N_18763,N_16539);
or UO_1468 (O_1468,N_17325,N_19456);
xnor UO_1469 (O_1469,N_17577,N_18823);
nor UO_1470 (O_1470,N_18906,N_19265);
nand UO_1471 (O_1471,N_16089,N_19347);
or UO_1472 (O_1472,N_17710,N_16943);
or UO_1473 (O_1473,N_17665,N_18916);
nand UO_1474 (O_1474,N_18466,N_19155);
nand UO_1475 (O_1475,N_17273,N_19975);
nand UO_1476 (O_1476,N_16507,N_18364);
or UO_1477 (O_1477,N_19311,N_16287);
nor UO_1478 (O_1478,N_18054,N_18857);
and UO_1479 (O_1479,N_16386,N_17393);
and UO_1480 (O_1480,N_18543,N_16549);
and UO_1481 (O_1481,N_18788,N_18212);
xor UO_1482 (O_1482,N_19126,N_17599);
nor UO_1483 (O_1483,N_17472,N_16920);
or UO_1484 (O_1484,N_18984,N_18463);
and UO_1485 (O_1485,N_16325,N_16699);
nand UO_1486 (O_1486,N_18667,N_19113);
nand UO_1487 (O_1487,N_16863,N_18475);
and UO_1488 (O_1488,N_16642,N_18061);
and UO_1489 (O_1489,N_17256,N_18468);
and UO_1490 (O_1490,N_16197,N_19424);
and UO_1491 (O_1491,N_17212,N_17137);
and UO_1492 (O_1492,N_19136,N_17961);
or UO_1493 (O_1493,N_19173,N_18487);
nand UO_1494 (O_1494,N_19790,N_16369);
nand UO_1495 (O_1495,N_18722,N_17967);
and UO_1496 (O_1496,N_17853,N_16906);
or UO_1497 (O_1497,N_17448,N_18658);
nor UO_1498 (O_1498,N_18981,N_19037);
and UO_1499 (O_1499,N_18696,N_16726);
nand UO_1500 (O_1500,N_19730,N_17973);
xnor UO_1501 (O_1501,N_18474,N_18867);
and UO_1502 (O_1502,N_16835,N_19725);
and UO_1503 (O_1503,N_16187,N_17328);
and UO_1504 (O_1504,N_16159,N_16790);
or UO_1505 (O_1505,N_16305,N_19885);
xor UO_1506 (O_1506,N_18861,N_19815);
nor UO_1507 (O_1507,N_16524,N_16468);
nand UO_1508 (O_1508,N_16184,N_16508);
or UO_1509 (O_1509,N_16451,N_18165);
or UO_1510 (O_1510,N_19408,N_19798);
xnor UO_1511 (O_1511,N_17367,N_19835);
xor UO_1512 (O_1512,N_19858,N_17801);
nand UO_1513 (O_1513,N_18444,N_18987);
or UO_1514 (O_1514,N_18778,N_17830);
or UO_1515 (O_1515,N_19767,N_17438);
or UO_1516 (O_1516,N_16718,N_19967);
nand UO_1517 (O_1517,N_19539,N_19529);
and UO_1518 (O_1518,N_19161,N_19884);
nand UO_1519 (O_1519,N_16066,N_16366);
or UO_1520 (O_1520,N_19353,N_17667);
and UO_1521 (O_1521,N_18734,N_16632);
xor UO_1522 (O_1522,N_19934,N_18750);
or UO_1523 (O_1523,N_19705,N_17909);
or UO_1524 (O_1524,N_17228,N_16054);
nor UO_1525 (O_1525,N_17416,N_18911);
and UO_1526 (O_1526,N_16264,N_16461);
or UO_1527 (O_1527,N_17079,N_19446);
nand UO_1528 (O_1528,N_18953,N_17012);
nand UO_1529 (O_1529,N_17213,N_17879);
nand UO_1530 (O_1530,N_16925,N_18377);
or UO_1531 (O_1531,N_17732,N_17838);
nand UO_1532 (O_1532,N_17989,N_19004);
nor UO_1533 (O_1533,N_16236,N_17884);
nor UO_1534 (O_1534,N_16883,N_17303);
nand UO_1535 (O_1535,N_18479,N_19563);
nor UO_1536 (O_1536,N_18592,N_18770);
nor UO_1537 (O_1537,N_19825,N_18961);
nand UO_1538 (O_1538,N_19296,N_17349);
or UO_1539 (O_1539,N_18168,N_16425);
and UO_1540 (O_1540,N_18452,N_17843);
nor UO_1541 (O_1541,N_18693,N_16388);
or UO_1542 (O_1542,N_18052,N_18945);
nand UO_1543 (O_1543,N_17363,N_19530);
xor UO_1544 (O_1544,N_17565,N_18125);
xor UO_1545 (O_1545,N_16174,N_19683);
nand UO_1546 (O_1546,N_18567,N_19693);
xnor UO_1547 (O_1547,N_19827,N_19023);
or UO_1548 (O_1548,N_16543,N_18736);
or UO_1549 (O_1549,N_18777,N_17241);
or UO_1550 (O_1550,N_18640,N_19654);
xnor UO_1551 (O_1551,N_17685,N_17353);
nor UO_1552 (O_1552,N_16057,N_16328);
nand UO_1553 (O_1553,N_18005,N_19939);
xnor UO_1554 (O_1554,N_18520,N_17679);
and UO_1555 (O_1555,N_16493,N_18412);
or UO_1556 (O_1556,N_19916,N_17318);
xnor UO_1557 (O_1557,N_18747,N_18145);
and UO_1558 (O_1558,N_18824,N_19556);
nand UO_1559 (O_1559,N_16620,N_19519);
xnor UO_1560 (O_1560,N_17193,N_16599);
xnor UO_1561 (O_1561,N_18767,N_17418);
and UO_1562 (O_1562,N_16687,N_19810);
nand UO_1563 (O_1563,N_16419,N_19368);
nor UO_1564 (O_1564,N_19966,N_16161);
nand UO_1565 (O_1565,N_16873,N_17032);
nor UO_1566 (O_1566,N_19926,N_18111);
nor UO_1567 (O_1567,N_19099,N_18341);
nand UO_1568 (O_1568,N_16116,N_16357);
and UO_1569 (O_1569,N_16937,N_18996);
nand UO_1570 (O_1570,N_19504,N_18603);
nand UO_1571 (O_1571,N_16209,N_17842);
and UO_1572 (O_1572,N_19942,N_19026);
or UO_1573 (O_1573,N_17277,N_19239);
and UO_1574 (O_1574,N_18772,N_19447);
and UO_1575 (O_1575,N_18130,N_19151);
nor UO_1576 (O_1576,N_18216,N_16080);
nand UO_1577 (O_1577,N_16928,N_18499);
nand UO_1578 (O_1578,N_19546,N_19804);
and UO_1579 (O_1579,N_18230,N_18333);
or UO_1580 (O_1580,N_16637,N_18411);
or UO_1581 (O_1581,N_18742,N_17071);
or UO_1582 (O_1582,N_16681,N_16750);
or UO_1583 (O_1583,N_19645,N_18235);
xor UO_1584 (O_1584,N_16358,N_18433);
xnor UO_1585 (O_1585,N_19555,N_16345);
xor UO_1586 (O_1586,N_18476,N_16700);
and UO_1587 (O_1587,N_17310,N_18816);
and UO_1588 (O_1588,N_18108,N_17214);
nor UO_1589 (O_1589,N_16212,N_16020);
nor UO_1590 (O_1590,N_18153,N_17564);
xnor UO_1591 (O_1591,N_19565,N_19024);
nand UO_1592 (O_1592,N_19395,N_19340);
xor UO_1593 (O_1593,N_19371,N_18586);
or UO_1594 (O_1594,N_19145,N_16343);
nand UO_1595 (O_1595,N_16717,N_16550);
nand UO_1596 (O_1596,N_17141,N_19677);
xnor UO_1597 (O_1597,N_18467,N_18725);
or UO_1598 (O_1598,N_16996,N_17003);
and UO_1599 (O_1599,N_16394,N_19304);
nand UO_1600 (O_1600,N_19496,N_18285);
and UO_1601 (O_1601,N_19891,N_18294);
xor UO_1602 (O_1602,N_17868,N_17356);
or UO_1603 (O_1603,N_16168,N_16214);
nor UO_1604 (O_1604,N_18671,N_19651);
nor UO_1605 (O_1605,N_17802,N_16654);
and UO_1606 (O_1606,N_19540,N_18073);
nand UO_1607 (O_1607,N_17401,N_18422);
and UO_1608 (O_1608,N_19380,N_19083);
xnor UO_1609 (O_1609,N_16324,N_16710);
and UO_1610 (O_1610,N_19439,N_17862);
nor UO_1611 (O_1611,N_19152,N_18243);
xnor UO_1612 (O_1612,N_18303,N_19698);
nand UO_1613 (O_1613,N_18515,N_19836);
nand UO_1614 (O_1614,N_16701,N_18146);
nor UO_1615 (O_1615,N_16308,N_18576);
and UO_1616 (O_1616,N_19508,N_16145);
nand UO_1617 (O_1617,N_17288,N_19894);
nor UO_1618 (O_1618,N_19174,N_17319);
and UO_1619 (O_1619,N_16747,N_18642);
nand UO_1620 (O_1620,N_19920,N_18186);
or UO_1621 (O_1621,N_17790,N_18233);
xnor UO_1622 (O_1622,N_17760,N_17729);
and UO_1623 (O_1623,N_16912,N_18070);
nand UO_1624 (O_1624,N_19685,N_19474);
nor UO_1625 (O_1625,N_18883,N_17415);
nor UO_1626 (O_1626,N_16181,N_16362);
xnor UO_1627 (O_1627,N_16074,N_19971);
and UO_1628 (O_1628,N_16408,N_17984);
or UO_1629 (O_1629,N_18785,N_16151);
xor UO_1630 (O_1630,N_19182,N_17727);
xor UO_1631 (O_1631,N_19898,N_16713);
or UO_1632 (O_1632,N_18546,N_17248);
or UO_1633 (O_1633,N_19428,N_18194);
nand UO_1634 (O_1634,N_19133,N_17264);
xnor UO_1635 (O_1635,N_19027,N_18554);
xnor UO_1636 (O_1636,N_16927,N_17033);
nor UO_1637 (O_1637,N_17226,N_17818);
nand UO_1638 (O_1638,N_19299,N_19499);
and UO_1639 (O_1639,N_18440,N_17837);
nor UO_1640 (O_1640,N_19623,N_19144);
nor UO_1641 (O_1641,N_19192,N_18241);
nand UO_1642 (O_1642,N_16477,N_17076);
and UO_1643 (O_1643,N_19345,N_19841);
and UO_1644 (O_1644,N_17134,N_16702);
or UO_1645 (O_1645,N_19562,N_16458);
or UO_1646 (O_1646,N_16519,N_18537);
xor UO_1647 (O_1647,N_19084,N_17890);
nor UO_1648 (O_1648,N_16299,N_16069);
xor UO_1649 (O_1649,N_17525,N_19326);
nand UO_1650 (O_1650,N_18853,N_19855);
nor UO_1651 (O_1651,N_19058,N_16136);
xor UO_1652 (O_1652,N_17333,N_17455);
nand UO_1653 (O_1653,N_17000,N_19165);
xor UO_1654 (O_1654,N_17848,N_17236);
nor UO_1655 (O_1655,N_18055,N_17874);
nand UO_1656 (O_1656,N_19294,N_18868);
and UO_1657 (O_1657,N_16815,N_16754);
and UO_1658 (O_1658,N_16641,N_19682);
xor UO_1659 (O_1659,N_17342,N_17863);
nor UO_1660 (O_1660,N_19962,N_17383);
nand UO_1661 (O_1661,N_16008,N_18874);
nand UO_1662 (O_1662,N_16235,N_18486);
xnor UO_1663 (O_1663,N_18057,N_19661);
and UO_1664 (O_1664,N_17084,N_17495);
nor UO_1665 (O_1665,N_18264,N_17298);
nand UO_1666 (O_1666,N_18617,N_19146);
or UO_1667 (O_1667,N_19183,N_18309);
or UO_1668 (O_1668,N_19585,N_17203);
xor UO_1669 (O_1669,N_17901,N_18888);
or UO_1670 (O_1670,N_17912,N_17395);
or UO_1671 (O_1671,N_19919,N_18060);
or UO_1672 (O_1672,N_19905,N_16404);
xor UO_1673 (O_1673,N_18390,N_17657);
nand UO_1674 (O_1674,N_18250,N_16656);
and UO_1675 (O_1675,N_18563,N_19193);
nand UO_1676 (O_1676,N_17466,N_17594);
and UO_1677 (O_1677,N_16866,N_17663);
or UO_1678 (O_1678,N_19471,N_17806);
nor UO_1679 (O_1679,N_16424,N_19704);
xor UO_1680 (O_1680,N_19374,N_17027);
xnor UO_1681 (O_1681,N_19793,N_18118);
nor UO_1682 (O_1682,N_19902,N_18548);
nand UO_1683 (O_1683,N_16935,N_16526);
xor UO_1684 (O_1684,N_18907,N_18615);
nand UO_1685 (O_1685,N_16745,N_18760);
xnor UO_1686 (O_1686,N_18404,N_18610);
nand UO_1687 (O_1687,N_16517,N_16205);
nor UO_1688 (O_1688,N_16607,N_18415);
and UO_1689 (O_1689,N_16968,N_19247);
nor UO_1690 (O_1690,N_16506,N_17411);
xor UO_1691 (O_1691,N_19533,N_18796);
and UO_1692 (O_1692,N_18768,N_19481);
or UO_1693 (O_1693,N_17223,N_17881);
nor UO_1694 (O_1694,N_18058,N_17579);
nand UO_1695 (O_1695,N_17487,N_17533);
nor UO_1696 (O_1696,N_19333,N_18726);
nor UO_1697 (O_1697,N_19650,N_19194);
nor UO_1698 (O_1698,N_16431,N_18743);
nand UO_1699 (O_1699,N_19741,N_19889);
nor UO_1700 (O_1700,N_16915,N_16634);
or UO_1701 (O_1701,N_18304,N_18947);
xor UO_1702 (O_1702,N_18866,N_18200);
nor UO_1703 (O_1703,N_19595,N_17544);
nand UO_1704 (O_1704,N_19071,N_16921);
nor UO_1705 (O_1705,N_18350,N_17550);
nor UO_1706 (O_1706,N_16744,N_18459);
nand UO_1707 (O_1707,N_17702,N_16981);
nor UO_1708 (O_1708,N_19550,N_18513);
nand UO_1709 (O_1709,N_19079,N_16064);
or UO_1710 (O_1710,N_18407,N_18706);
xnor UO_1711 (O_1711,N_19233,N_19038);
or UO_1712 (O_1712,N_19433,N_17969);
or UO_1713 (O_1713,N_18708,N_19185);
nand UO_1714 (O_1714,N_19570,N_19417);
or UO_1715 (O_1715,N_16384,N_18761);
xnor UO_1716 (O_1716,N_16050,N_18538);
and UO_1717 (O_1717,N_19797,N_16334);
or UO_1718 (O_1718,N_17676,N_16254);
xor UO_1719 (O_1719,N_16443,N_16917);
nand UO_1720 (O_1720,N_18774,N_17371);
nand UO_1721 (O_1721,N_18622,N_17290);
xnor UO_1722 (O_1722,N_17828,N_17650);
and UO_1723 (O_1723,N_17690,N_16276);
xor UO_1724 (O_1724,N_19229,N_19843);
and UO_1725 (O_1725,N_18234,N_18348);
or UO_1726 (O_1726,N_16558,N_18579);
xnor UO_1727 (O_1727,N_18935,N_19800);
nand UO_1728 (O_1728,N_18431,N_17512);
xnor UO_1729 (O_1729,N_17615,N_16387);
nand UO_1730 (O_1730,N_19322,N_19757);
or UO_1731 (O_1731,N_16950,N_18596);
or UO_1732 (O_1732,N_17494,N_19214);
and UO_1733 (O_1733,N_17419,N_18630);
nor UO_1734 (O_1734,N_16535,N_18930);
and UO_1735 (O_1735,N_16643,N_16746);
nand UO_1736 (O_1736,N_17314,N_19572);
xor UO_1737 (O_1737,N_19132,N_18107);
nand UO_1738 (O_1738,N_19577,N_19611);
nor UO_1739 (O_1739,N_19933,N_17144);
nand UO_1740 (O_1740,N_16121,N_16439);
nor UO_1741 (O_1741,N_18464,N_18105);
nand UO_1742 (O_1742,N_19581,N_18577);
or UO_1743 (O_1743,N_18011,N_19414);
nand UO_1744 (O_1744,N_17092,N_16893);
nand UO_1745 (O_1745,N_17722,N_18992);
and UO_1746 (O_1746,N_17364,N_18677);
nor UO_1747 (O_1747,N_16971,N_18800);
xnor UO_1748 (O_1748,N_19484,N_17858);
nor UO_1749 (O_1749,N_19856,N_17980);
nand UO_1750 (O_1750,N_17556,N_19111);
or UO_1751 (O_1751,N_16070,N_17551);
and UO_1752 (O_1752,N_16005,N_19994);
nor UO_1753 (O_1753,N_17200,N_17692);
xor UO_1754 (O_1754,N_18522,N_19879);
xor UO_1755 (O_1755,N_18365,N_16740);
nand UO_1756 (O_1756,N_18315,N_19415);
or UO_1757 (O_1757,N_19932,N_18481);
nand UO_1758 (O_1758,N_19765,N_18872);
or UO_1759 (O_1759,N_17956,N_17238);
or UO_1760 (O_1760,N_18156,N_19222);
and UO_1761 (O_1761,N_18937,N_17041);
and UO_1762 (O_1762,N_18138,N_16065);
or UO_1763 (O_1763,N_17021,N_18594);
nand UO_1764 (O_1764,N_18257,N_16765);
and UO_1765 (O_1765,N_17400,N_19639);
and UO_1766 (O_1766,N_16646,N_19986);
or UO_1767 (O_1767,N_16164,N_16752);
nand UO_1768 (O_1768,N_16017,N_17014);
or UO_1769 (O_1769,N_19482,N_17674);
or UO_1770 (O_1770,N_17119,N_18710);
nor UO_1771 (O_1771,N_19034,N_16678);
or UO_1772 (O_1772,N_17536,N_16733);
nor UO_1773 (O_1773,N_16298,N_18101);
xnor UO_1774 (O_1774,N_17278,N_18516);
and UO_1775 (O_1775,N_19432,N_17309);
and UO_1776 (O_1776,N_16794,N_18178);
nand UO_1777 (O_1777,N_19564,N_18585);
and UO_1778 (O_1778,N_17852,N_17535);
or UO_1779 (O_1779,N_19344,N_16049);
nor UO_1780 (O_1780,N_16035,N_16157);
xnor UO_1781 (O_1781,N_17282,N_19575);
nor UO_1782 (O_1782,N_19422,N_17652);
nor UO_1783 (O_1783,N_19129,N_18966);
xnor UO_1784 (O_1784,N_18183,N_18071);
nand UO_1785 (O_1785,N_18001,N_19813);
xnor UO_1786 (O_1786,N_18504,N_19638);
nand UO_1787 (O_1787,N_18038,N_17169);
xnor UO_1788 (O_1788,N_17305,N_19215);
and UO_1789 (O_1789,N_18405,N_16062);
nand UO_1790 (O_1790,N_17870,N_16831);
or UO_1791 (O_1791,N_18895,N_16655);
xor UO_1792 (O_1792,N_16834,N_16826);
and UO_1793 (O_1793,N_19631,N_16216);
or UO_1794 (O_1794,N_19190,N_18268);
nand UO_1795 (O_1795,N_18632,N_16088);
or UO_1796 (O_1796,N_19599,N_16289);
xnor UO_1797 (O_1797,N_18820,N_18988);
xnor UO_1798 (O_1798,N_17711,N_16243);
nand UO_1799 (O_1799,N_18860,N_16469);
nand UO_1800 (O_1800,N_17899,N_18062);
or UO_1801 (O_1801,N_17960,N_18410);
and UO_1802 (O_1802,N_16346,N_18912);
xor UO_1803 (O_1803,N_17521,N_16584);
nand UO_1804 (O_1804,N_17580,N_17759);
nor UO_1805 (O_1805,N_16146,N_19708);
or UO_1806 (O_1806,N_18084,N_17728);
and UO_1807 (O_1807,N_18914,N_17954);
or UO_1808 (O_1808,N_19321,N_17261);
nor UO_1809 (O_1809,N_18265,N_17143);
and UO_1810 (O_1810,N_18376,N_19197);
nand UO_1811 (O_1811,N_19763,N_16636);
or UO_1812 (O_1812,N_17633,N_16225);
nor UO_1813 (O_1813,N_19505,N_16763);
and UO_1814 (O_1814,N_17054,N_19608);
nor UO_1815 (O_1815,N_16685,N_19473);
and UO_1816 (O_1816,N_19928,N_16870);
nand UO_1817 (O_1817,N_17175,N_19308);
nand UO_1818 (O_1818,N_18815,N_16260);
xnor UO_1819 (O_1819,N_16051,N_17338);
or UO_1820 (O_1820,N_17154,N_16918);
xnor UO_1821 (O_1821,N_16463,N_18932);
or UO_1822 (O_1822,N_18447,N_19336);
nand UO_1823 (O_1823,N_17498,N_18320);
or UO_1824 (O_1824,N_17589,N_19312);
xor UO_1825 (O_1825,N_18699,N_19453);
nand UO_1826 (O_1826,N_17571,N_19313);
nand UO_1827 (O_1827,N_19527,N_16821);
nor UO_1828 (O_1828,N_17320,N_16238);
xnor UO_1829 (O_1829,N_19657,N_18161);
xnor UO_1830 (O_1830,N_18227,N_16271);
xnor UO_1831 (O_1831,N_16875,N_18759);
xor UO_1832 (O_1832,N_16409,N_17566);
and UO_1833 (O_1833,N_17721,N_18568);
and UO_1834 (O_1834,N_19383,N_19627);
or UO_1835 (O_1835,N_16037,N_19139);
nor UO_1836 (O_1836,N_17754,N_17791);
and UO_1837 (O_1837,N_17671,N_19072);
and UO_1838 (O_1838,N_19015,N_16453);
xor UO_1839 (O_1839,N_19792,N_17398);
xnor UO_1840 (O_1840,N_19381,N_19713);
and UO_1841 (O_1841,N_16217,N_19520);
and UO_1842 (O_1842,N_16773,N_18092);
and UO_1843 (O_1843,N_19008,N_19597);
xnor UO_1844 (O_1844,N_19701,N_16079);
nand UO_1845 (O_1845,N_16753,N_16779);
xor UO_1846 (O_1846,N_16082,N_16258);
xor UO_1847 (O_1847,N_17873,N_16075);
or UO_1848 (O_1848,N_16393,N_17271);
nor UO_1849 (O_1849,N_18065,N_16631);
xor UO_1850 (O_1850,N_16382,N_18353);
or UO_1851 (O_1851,N_16279,N_19754);
or UO_1852 (O_1852,N_19458,N_17350);
nand UO_1853 (O_1853,N_19121,N_18518);
and UO_1854 (O_1854,N_19993,N_17939);
or UO_1855 (O_1855,N_18313,N_16889);
nor UO_1856 (O_1856,N_18731,N_18944);
and UO_1857 (O_1857,N_18154,N_17546);
and UO_1858 (O_1858,N_17601,N_18965);
nand UO_1859 (O_1859,N_16018,N_17946);
and UO_1860 (O_1860,N_16335,N_17059);
and UO_1861 (O_1861,N_18223,N_19270);
and UO_1862 (O_1862,N_17315,N_16315);
xor UO_1863 (O_1863,N_17235,N_16787);
and UO_1864 (O_1864,N_19946,N_19629);
nand UO_1865 (O_1865,N_17854,N_17039);
nand UO_1866 (O_1866,N_17399,N_18396);
nor UO_1867 (O_1867,N_18369,N_16855);
xor UO_1868 (O_1868,N_17520,N_16649);
nor UO_1869 (O_1869,N_19025,N_16995);
or UO_1870 (O_1870,N_16314,N_17996);
nor UO_1871 (O_1871,N_16323,N_16862);
and UO_1872 (O_1872,N_19646,N_17737);
or UO_1873 (O_1873,N_19770,N_19268);
or UO_1874 (O_1874,N_17958,N_17083);
nor UO_1875 (O_1875,N_16882,N_19637);
and UO_1876 (O_1876,N_19149,N_17016);
and UO_1877 (O_1877,N_16224,N_16230);
and UO_1878 (O_1878,N_16810,N_19749);
nor UO_1879 (O_1879,N_19771,N_17327);
and UO_1880 (O_1880,N_18624,N_19999);
nand UO_1881 (O_1881,N_16203,N_17480);
and UO_1882 (O_1882,N_18637,N_16250);
and UO_1883 (O_1883,N_16682,N_17952);
nor UO_1884 (O_1884,N_17075,N_17106);
nand UO_1885 (O_1885,N_18025,N_19903);
nand UO_1886 (O_1886,N_18202,N_17846);
and UO_1887 (O_1887,N_18120,N_18502);
and UO_1888 (O_1888,N_18211,N_19266);
nand UO_1889 (O_1889,N_18540,N_19285);
nand UO_1890 (O_1890,N_16942,N_19110);
and UO_1891 (O_1891,N_19586,N_17859);
or UO_1892 (O_1892,N_19120,N_19720);
xor UO_1893 (O_1893,N_17372,N_17574);
xor UO_1894 (O_1894,N_18781,N_18920);
xnor UO_1895 (O_1895,N_17911,N_16498);
nand UO_1896 (O_1896,N_19179,N_19893);
xor UO_1897 (O_1897,N_19896,N_17357);
nand UO_1898 (O_1898,N_17554,N_18086);
xor UO_1899 (O_1899,N_19892,N_17755);
xor UO_1900 (O_1900,N_17919,N_16417);
nor UO_1901 (O_1901,N_18210,N_16894);
xor UO_1902 (O_1902,N_17629,N_16686);
xor UO_1903 (O_1903,N_18525,N_17444);
nor UO_1904 (O_1904,N_17042,N_17378);
and UO_1905 (O_1905,N_19772,N_18511);
xor UO_1906 (O_1906,N_16288,N_16929);
xor UO_1907 (O_1907,N_18793,N_17171);
nand UO_1908 (O_1908,N_16061,N_18856);
xor UO_1909 (O_1909,N_17673,N_19314);
or UO_1910 (O_1910,N_17617,N_16983);
nand UO_1911 (O_1911,N_17281,N_18942);
nand UO_1912 (O_1912,N_16505,N_19578);
and UO_1913 (O_1913,N_18089,N_16316);
or UO_1914 (O_1914,N_17770,N_18002);
or UO_1915 (O_1915,N_17825,N_18924);
nor UO_1916 (O_1916,N_18711,N_18809);
and UO_1917 (O_1917,N_16242,N_19463);
nand UO_1918 (O_1918,N_19168,N_18994);
and UO_1919 (O_1919,N_16728,N_17841);
and UO_1920 (O_1920,N_16090,N_19931);
nand UO_1921 (O_1921,N_16727,N_18528);
or UO_1922 (O_1922,N_19782,N_16963);
nand UO_1923 (O_1923,N_18036,N_19531);
or UO_1924 (O_1924,N_17478,N_18331);
and UO_1925 (O_1925,N_18450,N_16901);
xor UO_1926 (O_1926,N_17190,N_19323);
nor UO_1927 (O_1927,N_16024,N_16660);
nor UO_1928 (O_1928,N_16042,N_16475);
xnor UO_1929 (O_1929,N_19769,N_17709);
nor UO_1930 (O_1930,N_16441,N_16839);
xor UO_1931 (O_1931,N_19398,N_17463);
and UO_1932 (O_1932,N_16854,N_16738);
and UO_1933 (O_1933,N_19909,N_17726);
or UO_1934 (O_1934,N_16142,N_19842);
nor UO_1935 (O_1935,N_19554,N_16801);
or UO_1936 (O_1936,N_19370,N_16359);
nand UO_1937 (O_1937,N_19223,N_16545);
nor UO_1938 (O_1938,N_17775,N_19762);
nand UO_1939 (O_1939,N_16460,N_17923);
xnor UO_1940 (O_1940,N_17009,N_19694);
and UO_1941 (O_1941,N_18012,N_17108);
and UO_1942 (O_1942,N_16277,N_18076);
nor UO_1943 (O_1943,N_16001,N_17815);
nand UO_1944 (O_1944,N_19087,N_16129);
or UO_1945 (O_1945,N_17827,N_18391);
and UO_1946 (O_1946,N_19480,N_16934);
and UO_1947 (O_1947,N_17443,N_19154);
or UO_1948 (O_1948,N_18553,N_16939);
and UO_1949 (O_1949,N_19055,N_16822);
nor UO_1950 (O_1950,N_19969,N_18041);
nor UO_1951 (O_1951,N_19850,N_17026);
and UO_1952 (O_1952,N_18276,N_16922);
xnor UO_1953 (O_1953,N_17107,N_19300);
xnor UO_1954 (O_1954,N_18694,N_18973);
and UO_1955 (O_1955,N_18337,N_19252);
nand UO_1956 (O_1956,N_19106,N_17376);
nor UO_1957 (O_1957,N_19319,N_16455);
and UO_1958 (O_1958,N_17269,N_18882);
and UO_1959 (O_1959,N_17636,N_17656);
xor UO_1960 (O_1960,N_16132,N_16544);
nor UO_1961 (O_1961,N_16770,N_18580);
or UO_1962 (O_1962,N_19632,N_19731);
xor UO_1963 (O_1963,N_17530,N_16178);
or UO_1964 (O_1964,N_18600,N_17492);
nor UO_1965 (O_1965,N_19630,N_18299);
nand UO_1966 (O_1966,N_16310,N_19857);
nand UO_1967 (O_1967,N_16026,N_17584);
nand UO_1968 (O_1968,N_19341,N_17454);
xnor UO_1969 (O_1969,N_16073,N_18147);
or UO_1970 (O_1970,N_18864,N_17686);
nor UO_1971 (O_1971,N_19365,N_16467);
or UO_1972 (O_1972,N_19217,N_18581);
xnor UO_1973 (O_1973,N_17412,N_16420);
and UO_1974 (O_1974,N_19277,N_19516);
xnor UO_1975 (O_1975,N_19042,N_16444);
or UO_1976 (O_1976,N_17425,N_16778);
and UO_1977 (O_1977,N_17597,N_18755);
nor UO_1978 (O_1978,N_16456,N_18527);
xnor UO_1979 (O_1979,N_17294,N_16557);
or UO_1980 (O_1980,N_16331,N_17985);
xor UO_1981 (O_1981,N_17634,N_18379);
nor UO_1982 (O_1982,N_16571,N_16041);
nand UO_1983 (O_1983,N_18588,N_17793);
nand UO_1984 (O_1984,N_16491,N_17004);
xnor UO_1985 (O_1985,N_19860,N_18695);
and UO_1986 (O_1986,N_17481,N_17111);
nor UO_1987 (O_1987,N_16988,N_17201);
nand UO_1988 (O_1988,N_18172,N_18898);
and UO_1989 (O_1989,N_17637,N_19356);
or UO_1990 (O_1990,N_17757,N_19618);
nor UO_1991 (O_1991,N_17094,N_17451);
xnor UO_1992 (O_1992,N_18998,N_18112);
nand UO_1993 (O_1993,N_17105,N_18483);
nor UO_1994 (O_1994,N_16992,N_19431);
xor UO_1995 (O_1995,N_19043,N_19911);
and UO_1996 (O_1996,N_19863,N_17872);
and UO_1997 (O_1997,N_19451,N_17373);
nand UO_1998 (O_1998,N_17724,N_18351);
nand UO_1999 (O_1999,N_17962,N_17749);
nand UO_2000 (O_2000,N_18831,N_17414);
and UO_2001 (O_2001,N_16183,N_19125);
nor UO_2002 (O_2002,N_18695,N_18401);
nor UO_2003 (O_2003,N_19570,N_18297);
or UO_2004 (O_2004,N_16463,N_19998);
xor UO_2005 (O_2005,N_17255,N_18967);
or UO_2006 (O_2006,N_17469,N_19542);
or UO_2007 (O_2007,N_19783,N_19138);
or UO_2008 (O_2008,N_16033,N_18527);
nand UO_2009 (O_2009,N_17552,N_16947);
and UO_2010 (O_2010,N_16108,N_17465);
nand UO_2011 (O_2011,N_19937,N_19217);
nor UO_2012 (O_2012,N_19059,N_18577);
xnor UO_2013 (O_2013,N_16200,N_18366);
xor UO_2014 (O_2014,N_19180,N_17570);
or UO_2015 (O_2015,N_18575,N_16962);
nor UO_2016 (O_2016,N_17197,N_17089);
nor UO_2017 (O_2017,N_17060,N_18508);
or UO_2018 (O_2018,N_16786,N_18626);
or UO_2019 (O_2019,N_17257,N_18364);
nand UO_2020 (O_2020,N_18944,N_17284);
and UO_2021 (O_2021,N_16977,N_16839);
xor UO_2022 (O_2022,N_19080,N_17289);
nor UO_2023 (O_2023,N_17594,N_17458);
xor UO_2024 (O_2024,N_17605,N_17448);
xnor UO_2025 (O_2025,N_18483,N_18557);
xnor UO_2026 (O_2026,N_16258,N_19058);
nand UO_2027 (O_2027,N_16683,N_17193);
nor UO_2028 (O_2028,N_19072,N_19219);
nand UO_2029 (O_2029,N_17216,N_19216);
nand UO_2030 (O_2030,N_16015,N_16022);
or UO_2031 (O_2031,N_17865,N_19202);
nor UO_2032 (O_2032,N_17563,N_16113);
nand UO_2033 (O_2033,N_17825,N_16227);
nor UO_2034 (O_2034,N_18401,N_18479);
nor UO_2035 (O_2035,N_16015,N_18098);
nor UO_2036 (O_2036,N_16773,N_16547);
nor UO_2037 (O_2037,N_16190,N_16118);
or UO_2038 (O_2038,N_19538,N_17046);
nand UO_2039 (O_2039,N_16755,N_19293);
nand UO_2040 (O_2040,N_19451,N_16273);
xnor UO_2041 (O_2041,N_16661,N_17015);
nor UO_2042 (O_2042,N_16021,N_19884);
and UO_2043 (O_2043,N_17622,N_19263);
xor UO_2044 (O_2044,N_19372,N_17000);
xnor UO_2045 (O_2045,N_16338,N_17578);
and UO_2046 (O_2046,N_17866,N_19518);
nor UO_2047 (O_2047,N_19479,N_18218);
xnor UO_2048 (O_2048,N_17941,N_16008);
nand UO_2049 (O_2049,N_17197,N_18197);
xnor UO_2050 (O_2050,N_16784,N_16884);
and UO_2051 (O_2051,N_17487,N_17979);
or UO_2052 (O_2052,N_16982,N_16623);
nand UO_2053 (O_2053,N_17826,N_19584);
xnor UO_2054 (O_2054,N_16870,N_19811);
nor UO_2055 (O_2055,N_17793,N_19291);
nor UO_2056 (O_2056,N_16333,N_18230);
nor UO_2057 (O_2057,N_17438,N_19550);
or UO_2058 (O_2058,N_17552,N_17050);
nor UO_2059 (O_2059,N_16298,N_17536);
and UO_2060 (O_2060,N_18699,N_17593);
nor UO_2061 (O_2061,N_19780,N_19990);
nor UO_2062 (O_2062,N_18086,N_17079);
nand UO_2063 (O_2063,N_16040,N_17774);
or UO_2064 (O_2064,N_18987,N_18190);
nor UO_2065 (O_2065,N_16411,N_17589);
or UO_2066 (O_2066,N_19954,N_17623);
xnor UO_2067 (O_2067,N_18665,N_19328);
or UO_2068 (O_2068,N_19994,N_19153);
xor UO_2069 (O_2069,N_19033,N_16626);
and UO_2070 (O_2070,N_19531,N_16695);
xor UO_2071 (O_2071,N_16383,N_16563);
and UO_2072 (O_2072,N_17118,N_17169);
and UO_2073 (O_2073,N_16496,N_19760);
or UO_2074 (O_2074,N_16230,N_16235);
or UO_2075 (O_2075,N_16007,N_17711);
nand UO_2076 (O_2076,N_18606,N_18555);
and UO_2077 (O_2077,N_19579,N_16601);
nor UO_2078 (O_2078,N_16295,N_17553);
and UO_2079 (O_2079,N_19556,N_16554);
and UO_2080 (O_2080,N_17384,N_18407);
or UO_2081 (O_2081,N_19470,N_16493);
xnor UO_2082 (O_2082,N_17482,N_16462);
and UO_2083 (O_2083,N_16912,N_19876);
and UO_2084 (O_2084,N_18084,N_18664);
and UO_2085 (O_2085,N_19716,N_16883);
nor UO_2086 (O_2086,N_19532,N_19486);
nor UO_2087 (O_2087,N_16904,N_18461);
and UO_2088 (O_2088,N_16816,N_17455);
nor UO_2089 (O_2089,N_16893,N_18100);
nand UO_2090 (O_2090,N_18092,N_18900);
nor UO_2091 (O_2091,N_16652,N_16593);
and UO_2092 (O_2092,N_18789,N_17772);
nand UO_2093 (O_2093,N_17135,N_18006);
nand UO_2094 (O_2094,N_16203,N_16794);
nand UO_2095 (O_2095,N_17646,N_18931);
xor UO_2096 (O_2096,N_19360,N_18829);
or UO_2097 (O_2097,N_16251,N_17797);
xor UO_2098 (O_2098,N_18546,N_19900);
or UO_2099 (O_2099,N_17153,N_18744);
or UO_2100 (O_2100,N_16007,N_17074);
nor UO_2101 (O_2101,N_19368,N_17016);
or UO_2102 (O_2102,N_16606,N_16846);
nor UO_2103 (O_2103,N_16655,N_17744);
nand UO_2104 (O_2104,N_16796,N_19646);
or UO_2105 (O_2105,N_16687,N_17167);
and UO_2106 (O_2106,N_17818,N_17038);
or UO_2107 (O_2107,N_17840,N_19761);
and UO_2108 (O_2108,N_18774,N_17986);
and UO_2109 (O_2109,N_17498,N_19051);
nor UO_2110 (O_2110,N_16049,N_18289);
nor UO_2111 (O_2111,N_16142,N_17680);
or UO_2112 (O_2112,N_18535,N_16647);
nand UO_2113 (O_2113,N_19319,N_18865);
nand UO_2114 (O_2114,N_16134,N_16088);
or UO_2115 (O_2115,N_16323,N_16007);
nor UO_2116 (O_2116,N_16499,N_19685);
nand UO_2117 (O_2117,N_16553,N_18287);
xor UO_2118 (O_2118,N_17885,N_16787);
or UO_2119 (O_2119,N_19471,N_19928);
or UO_2120 (O_2120,N_19750,N_19827);
nor UO_2121 (O_2121,N_17894,N_17029);
nor UO_2122 (O_2122,N_18871,N_17641);
xnor UO_2123 (O_2123,N_18772,N_16994);
nand UO_2124 (O_2124,N_18644,N_16699);
nand UO_2125 (O_2125,N_19677,N_16061);
or UO_2126 (O_2126,N_18674,N_18473);
or UO_2127 (O_2127,N_18228,N_16512);
and UO_2128 (O_2128,N_19378,N_19963);
nor UO_2129 (O_2129,N_19300,N_16574);
or UO_2130 (O_2130,N_19357,N_17537);
xor UO_2131 (O_2131,N_17179,N_19069);
and UO_2132 (O_2132,N_18044,N_18914);
and UO_2133 (O_2133,N_18402,N_17926);
nor UO_2134 (O_2134,N_16683,N_18208);
or UO_2135 (O_2135,N_18059,N_19983);
or UO_2136 (O_2136,N_16675,N_17412);
nand UO_2137 (O_2137,N_18161,N_19601);
nor UO_2138 (O_2138,N_18322,N_18671);
xor UO_2139 (O_2139,N_17754,N_18422);
nor UO_2140 (O_2140,N_17180,N_16319);
xor UO_2141 (O_2141,N_17239,N_16598);
xor UO_2142 (O_2142,N_19099,N_17607);
xnor UO_2143 (O_2143,N_19718,N_17508);
nor UO_2144 (O_2144,N_17213,N_19824);
nand UO_2145 (O_2145,N_16655,N_16485);
xnor UO_2146 (O_2146,N_19083,N_19594);
or UO_2147 (O_2147,N_17419,N_16315);
or UO_2148 (O_2148,N_16816,N_18092);
or UO_2149 (O_2149,N_18108,N_18706);
xnor UO_2150 (O_2150,N_19594,N_18720);
and UO_2151 (O_2151,N_19066,N_19724);
nand UO_2152 (O_2152,N_16198,N_18002);
and UO_2153 (O_2153,N_19752,N_16522);
xor UO_2154 (O_2154,N_16833,N_16190);
nor UO_2155 (O_2155,N_17347,N_17613);
and UO_2156 (O_2156,N_17520,N_19216);
xor UO_2157 (O_2157,N_16310,N_18313);
nand UO_2158 (O_2158,N_17899,N_19259);
and UO_2159 (O_2159,N_19782,N_16719);
xor UO_2160 (O_2160,N_18604,N_19191);
and UO_2161 (O_2161,N_16191,N_16081);
nor UO_2162 (O_2162,N_17099,N_17727);
nor UO_2163 (O_2163,N_17008,N_18679);
nor UO_2164 (O_2164,N_18474,N_19700);
and UO_2165 (O_2165,N_18707,N_17973);
xnor UO_2166 (O_2166,N_17337,N_19374);
xnor UO_2167 (O_2167,N_18485,N_18541);
nor UO_2168 (O_2168,N_16456,N_18450);
nand UO_2169 (O_2169,N_16260,N_19646);
nor UO_2170 (O_2170,N_19224,N_16347);
nor UO_2171 (O_2171,N_16995,N_16987);
xnor UO_2172 (O_2172,N_19830,N_19477);
xnor UO_2173 (O_2173,N_19293,N_18720);
nor UO_2174 (O_2174,N_17403,N_16485);
nand UO_2175 (O_2175,N_19600,N_19234);
xor UO_2176 (O_2176,N_17618,N_16730);
xor UO_2177 (O_2177,N_18255,N_17071);
nand UO_2178 (O_2178,N_17581,N_17330);
nand UO_2179 (O_2179,N_17817,N_17302);
nand UO_2180 (O_2180,N_19369,N_18877);
nor UO_2181 (O_2181,N_18433,N_17044);
nand UO_2182 (O_2182,N_19923,N_16368);
nor UO_2183 (O_2183,N_17776,N_19709);
nand UO_2184 (O_2184,N_16244,N_19935);
nor UO_2185 (O_2185,N_16531,N_17454);
xor UO_2186 (O_2186,N_19510,N_18513);
nand UO_2187 (O_2187,N_16238,N_18412);
xnor UO_2188 (O_2188,N_16972,N_18442);
xor UO_2189 (O_2189,N_18388,N_17554);
nand UO_2190 (O_2190,N_17455,N_17858);
nand UO_2191 (O_2191,N_19984,N_17288);
or UO_2192 (O_2192,N_18981,N_16434);
nand UO_2193 (O_2193,N_18645,N_19807);
xnor UO_2194 (O_2194,N_17962,N_17292);
or UO_2195 (O_2195,N_18275,N_18424);
nand UO_2196 (O_2196,N_18572,N_19370);
xnor UO_2197 (O_2197,N_19402,N_19350);
nor UO_2198 (O_2198,N_17767,N_19724);
and UO_2199 (O_2199,N_19203,N_18757);
or UO_2200 (O_2200,N_17228,N_17571);
nand UO_2201 (O_2201,N_16951,N_16510);
nand UO_2202 (O_2202,N_17682,N_19907);
nand UO_2203 (O_2203,N_18419,N_19974);
or UO_2204 (O_2204,N_18071,N_19505);
nand UO_2205 (O_2205,N_19206,N_19340);
xnor UO_2206 (O_2206,N_19519,N_16636);
nand UO_2207 (O_2207,N_16646,N_16198);
and UO_2208 (O_2208,N_16464,N_19274);
and UO_2209 (O_2209,N_18944,N_16580);
or UO_2210 (O_2210,N_18602,N_17682);
nor UO_2211 (O_2211,N_16215,N_17466);
nand UO_2212 (O_2212,N_16380,N_18770);
or UO_2213 (O_2213,N_16654,N_16748);
and UO_2214 (O_2214,N_16429,N_17963);
nand UO_2215 (O_2215,N_18434,N_19738);
nor UO_2216 (O_2216,N_16858,N_18227);
nor UO_2217 (O_2217,N_17804,N_16017);
or UO_2218 (O_2218,N_19531,N_17982);
nand UO_2219 (O_2219,N_17985,N_18144);
nor UO_2220 (O_2220,N_16012,N_17338);
nor UO_2221 (O_2221,N_16228,N_18471);
and UO_2222 (O_2222,N_19306,N_19652);
or UO_2223 (O_2223,N_16206,N_19120);
xor UO_2224 (O_2224,N_17275,N_19617);
xor UO_2225 (O_2225,N_17185,N_18624);
or UO_2226 (O_2226,N_16878,N_19718);
xnor UO_2227 (O_2227,N_19365,N_16868);
nor UO_2228 (O_2228,N_18018,N_19149);
nand UO_2229 (O_2229,N_19955,N_19996);
nor UO_2230 (O_2230,N_17537,N_17010);
nand UO_2231 (O_2231,N_18906,N_18765);
xnor UO_2232 (O_2232,N_17948,N_16545);
or UO_2233 (O_2233,N_18321,N_19171);
nand UO_2234 (O_2234,N_19292,N_16234);
nor UO_2235 (O_2235,N_17165,N_19982);
and UO_2236 (O_2236,N_17060,N_16669);
or UO_2237 (O_2237,N_17241,N_18668);
or UO_2238 (O_2238,N_16630,N_16463);
nand UO_2239 (O_2239,N_19726,N_19493);
xnor UO_2240 (O_2240,N_16114,N_18312);
xnor UO_2241 (O_2241,N_19182,N_16992);
xnor UO_2242 (O_2242,N_17937,N_18119);
and UO_2243 (O_2243,N_19566,N_19870);
nand UO_2244 (O_2244,N_17325,N_16518);
xor UO_2245 (O_2245,N_19081,N_18251);
nand UO_2246 (O_2246,N_19594,N_17569);
xnor UO_2247 (O_2247,N_19415,N_17372);
nand UO_2248 (O_2248,N_19952,N_16029);
xnor UO_2249 (O_2249,N_19329,N_16744);
or UO_2250 (O_2250,N_16297,N_17015);
nor UO_2251 (O_2251,N_18570,N_16168);
or UO_2252 (O_2252,N_18107,N_16169);
and UO_2253 (O_2253,N_16905,N_19336);
or UO_2254 (O_2254,N_18559,N_19362);
and UO_2255 (O_2255,N_18309,N_18276);
nand UO_2256 (O_2256,N_17093,N_18613);
xor UO_2257 (O_2257,N_19720,N_16569);
and UO_2258 (O_2258,N_18666,N_18005);
and UO_2259 (O_2259,N_16679,N_16287);
nand UO_2260 (O_2260,N_19001,N_17646);
or UO_2261 (O_2261,N_16533,N_18861);
nand UO_2262 (O_2262,N_18112,N_16726);
xor UO_2263 (O_2263,N_17326,N_18468);
and UO_2264 (O_2264,N_17827,N_16863);
nor UO_2265 (O_2265,N_18554,N_18734);
xnor UO_2266 (O_2266,N_18450,N_19645);
nand UO_2267 (O_2267,N_18122,N_17650);
xor UO_2268 (O_2268,N_16503,N_16780);
nand UO_2269 (O_2269,N_19831,N_18145);
xnor UO_2270 (O_2270,N_17563,N_19043);
xor UO_2271 (O_2271,N_16339,N_18419);
or UO_2272 (O_2272,N_18217,N_18656);
or UO_2273 (O_2273,N_18719,N_16234);
xor UO_2274 (O_2274,N_19446,N_19471);
nor UO_2275 (O_2275,N_17839,N_18346);
and UO_2276 (O_2276,N_16151,N_18307);
xnor UO_2277 (O_2277,N_16066,N_19873);
nor UO_2278 (O_2278,N_18118,N_18639);
or UO_2279 (O_2279,N_19894,N_18636);
nand UO_2280 (O_2280,N_16643,N_19223);
or UO_2281 (O_2281,N_17880,N_16834);
nor UO_2282 (O_2282,N_19770,N_19535);
xnor UO_2283 (O_2283,N_18203,N_17173);
or UO_2284 (O_2284,N_18418,N_17596);
or UO_2285 (O_2285,N_18272,N_17768);
nor UO_2286 (O_2286,N_19928,N_19011);
nor UO_2287 (O_2287,N_19136,N_19034);
nor UO_2288 (O_2288,N_17767,N_17922);
nand UO_2289 (O_2289,N_18037,N_19529);
or UO_2290 (O_2290,N_17188,N_16164);
xnor UO_2291 (O_2291,N_17628,N_16824);
nand UO_2292 (O_2292,N_17990,N_18747);
or UO_2293 (O_2293,N_16087,N_16066);
nor UO_2294 (O_2294,N_16139,N_17121);
nor UO_2295 (O_2295,N_16109,N_19290);
and UO_2296 (O_2296,N_16836,N_16089);
xor UO_2297 (O_2297,N_18437,N_19994);
or UO_2298 (O_2298,N_17664,N_16745);
nand UO_2299 (O_2299,N_18459,N_19703);
xor UO_2300 (O_2300,N_17111,N_17939);
nor UO_2301 (O_2301,N_19130,N_18779);
and UO_2302 (O_2302,N_19316,N_16592);
xor UO_2303 (O_2303,N_17677,N_17016);
nor UO_2304 (O_2304,N_19499,N_16555);
nor UO_2305 (O_2305,N_16895,N_19290);
or UO_2306 (O_2306,N_16499,N_17042);
nand UO_2307 (O_2307,N_17122,N_16447);
and UO_2308 (O_2308,N_19637,N_19841);
nor UO_2309 (O_2309,N_16440,N_19228);
xor UO_2310 (O_2310,N_18065,N_18599);
and UO_2311 (O_2311,N_19291,N_16549);
nor UO_2312 (O_2312,N_17714,N_19486);
or UO_2313 (O_2313,N_17251,N_19418);
nand UO_2314 (O_2314,N_19179,N_16667);
or UO_2315 (O_2315,N_19795,N_17790);
nor UO_2316 (O_2316,N_18451,N_17143);
xor UO_2317 (O_2317,N_19933,N_19380);
nand UO_2318 (O_2318,N_17604,N_18335);
nand UO_2319 (O_2319,N_19310,N_18026);
nor UO_2320 (O_2320,N_18478,N_18291);
xor UO_2321 (O_2321,N_17893,N_18255);
and UO_2322 (O_2322,N_16251,N_16400);
and UO_2323 (O_2323,N_19053,N_16199);
nand UO_2324 (O_2324,N_16790,N_18674);
and UO_2325 (O_2325,N_18525,N_19607);
xnor UO_2326 (O_2326,N_17344,N_18544);
or UO_2327 (O_2327,N_17036,N_16749);
nor UO_2328 (O_2328,N_16568,N_18492);
nand UO_2329 (O_2329,N_17322,N_17669);
xnor UO_2330 (O_2330,N_18827,N_16284);
nand UO_2331 (O_2331,N_17221,N_18384);
nor UO_2332 (O_2332,N_18842,N_17588);
xnor UO_2333 (O_2333,N_16544,N_17045);
and UO_2334 (O_2334,N_18198,N_16625);
and UO_2335 (O_2335,N_16933,N_19551);
xnor UO_2336 (O_2336,N_16092,N_18407);
nand UO_2337 (O_2337,N_18716,N_16322);
nand UO_2338 (O_2338,N_17337,N_19787);
xnor UO_2339 (O_2339,N_17498,N_18454);
nor UO_2340 (O_2340,N_18767,N_16764);
or UO_2341 (O_2341,N_19968,N_19989);
or UO_2342 (O_2342,N_19982,N_18505);
nand UO_2343 (O_2343,N_17451,N_18189);
and UO_2344 (O_2344,N_16806,N_16088);
xor UO_2345 (O_2345,N_16938,N_16025);
and UO_2346 (O_2346,N_17293,N_17012);
or UO_2347 (O_2347,N_19907,N_19791);
and UO_2348 (O_2348,N_18051,N_19372);
nor UO_2349 (O_2349,N_19585,N_16758);
xnor UO_2350 (O_2350,N_19458,N_16617);
or UO_2351 (O_2351,N_16103,N_16444);
nand UO_2352 (O_2352,N_18963,N_19587);
nor UO_2353 (O_2353,N_19653,N_16949);
or UO_2354 (O_2354,N_19481,N_18206);
and UO_2355 (O_2355,N_18596,N_16347);
and UO_2356 (O_2356,N_17027,N_18201);
nor UO_2357 (O_2357,N_18677,N_18376);
xor UO_2358 (O_2358,N_19641,N_18707);
nor UO_2359 (O_2359,N_17296,N_17052);
or UO_2360 (O_2360,N_17562,N_16107);
nor UO_2361 (O_2361,N_16061,N_16478);
nor UO_2362 (O_2362,N_16973,N_17932);
or UO_2363 (O_2363,N_18392,N_17748);
nor UO_2364 (O_2364,N_19565,N_19556);
or UO_2365 (O_2365,N_19128,N_19196);
or UO_2366 (O_2366,N_19946,N_19375);
or UO_2367 (O_2367,N_16138,N_16650);
and UO_2368 (O_2368,N_17639,N_18236);
or UO_2369 (O_2369,N_17619,N_18200);
and UO_2370 (O_2370,N_16428,N_18650);
xnor UO_2371 (O_2371,N_19372,N_17784);
nor UO_2372 (O_2372,N_19122,N_19998);
or UO_2373 (O_2373,N_19175,N_19197);
nand UO_2374 (O_2374,N_19195,N_19005);
nor UO_2375 (O_2375,N_19371,N_17218);
and UO_2376 (O_2376,N_18176,N_16897);
xnor UO_2377 (O_2377,N_16316,N_17331);
nor UO_2378 (O_2378,N_19059,N_17589);
xnor UO_2379 (O_2379,N_16689,N_18554);
or UO_2380 (O_2380,N_19424,N_18080);
or UO_2381 (O_2381,N_18485,N_17821);
nand UO_2382 (O_2382,N_19510,N_19981);
and UO_2383 (O_2383,N_18141,N_16113);
or UO_2384 (O_2384,N_17405,N_19115);
nor UO_2385 (O_2385,N_16505,N_16355);
and UO_2386 (O_2386,N_16341,N_18789);
nand UO_2387 (O_2387,N_19795,N_16448);
or UO_2388 (O_2388,N_19931,N_16738);
nand UO_2389 (O_2389,N_16391,N_18244);
and UO_2390 (O_2390,N_18730,N_19609);
nor UO_2391 (O_2391,N_19321,N_17292);
nor UO_2392 (O_2392,N_17630,N_16898);
or UO_2393 (O_2393,N_17276,N_19979);
xor UO_2394 (O_2394,N_17034,N_16914);
or UO_2395 (O_2395,N_19131,N_17214);
xor UO_2396 (O_2396,N_18311,N_17429);
and UO_2397 (O_2397,N_19785,N_16597);
nor UO_2398 (O_2398,N_18551,N_18905);
xor UO_2399 (O_2399,N_18913,N_17997);
nor UO_2400 (O_2400,N_17860,N_18903);
nand UO_2401 (O_2401,N_16420,N_16556);
nor UO_2402 (O_2402,N_17226,N_16853);
nand UO_2403 (O_2403,N_18406,N_18011);
or UO_2404 (O_2404,N_16402,N_16445);
or UO_2405 (O_2405,N_18951,N_19957);
and UO_2406 (O_2406,N_19319,N_19614);
or UO_2407 (O_2407,N_17537,N_18561);
nor UO_2408 (O_2408,N_17753,N_18432);
xor UO_2409 (O_2409,N_16487,N_17847);
and UO_2410 (O_2410,N_19541,N_16959);
or UO_2411 (O_2411,N_16148,N_18589);
or UO_2412 (O_2412,N_19795,N_17232);
nor UO_2413 (O_2413,N_19591,N_17345);
xnor UO_2414 (O_2414,N_19785,N_19084);
nand UO_2415 (O_2415,N_17665,N_18998);
nor UO_2416 (O_2416,N_18381,N_19977);
or UO_2417 (O_2417,N_17193,N_18551);
and UO_2418 (O_2418,N_19262,N_18735);
nand UO_2419 (O_2419,N_19543,N_18889);
xor UO_2420 (O_2420,N_19255,N_16522);
or UO_2421 (O_2421,N_17390,N_18769);
xor UO_2422 (O_2422,N_18901,N_16343);
nor UO_2423 (O_2423,N_19122,N_18625);
and UO_2424 (O_2424,N_19243,N_19235);
or UO_2425 (O_2425,N_16290,N_19335);
or UO_2426 (O_2426,N_16372,N_16670);
and UO_2427 (O_2427,N_16435,N_16881);
nand UO_2428 (O_2428,N_18802,N_19990);
nor UO_2429 (O_2429,N_18986,N_19318);
and UO_2430 (O_2430,N_18024,N_19715);
or UO_2431 (O_2431,N_18856,N_16486);
or UO_2432 (O_2432,N_18338,N_19550);
and UO_2433 (O_2433,N_19943,N_16938);
xor UO_2434 (O_2434,N_16116,N_19989);
nand UO_2435 (O_2435,N_19456,N_18229);
and UO_2436 (O_2436,N_18109,N_17937);
xnor UO_2437 (O_2437,N_16937,N_18198);
and UO_2438 (O_2438,N_17061,N_16652);
xnor UO_2439 (O_2439,N_19637,N_19653);
nand UO_2440 (O_2440,N_16791,N_19650);
nor UO_2441 (O_2441,N_17252,N_17563);
xnor UO_2442 (O_2442,N_16799,N_18950);
or UO_2443 (O_2443,N_17305,N_18969);
or UO_2444 (O_2444,N_19171,N_17632);
nand UO_2445 (O_2445,N_17533,N_17718);
or UO_2446 (O_2446,N_16204,N_18383);
nor UO_2447 (O_2447,N_17367,N_16861);
xnor UO_2448 (O_2448,N_17772,N_18350);
nor UO_2449 (O_2449,N_19359,N_18113);
nand UO_2450 (O_2450,N_16392,N_16442);
xor UO_2451 (O_2451,N_16886,N_16570);
xor UO_2452 (O_2452,N_19406,N_17135);
nor UO_2453 (O_2453,N_16100,N_19576);
xor UO_2454 (O_2454,N_19305,N_19258);
nor UO_2455 (O_2455,N_19070,N_17769);
xnor UO_2456 (O_2456,N_16938,N_19442);
xnor UO_2457 (O_2457,N_16135,N_19835);
nand UO_2458 (O_2458,N_19973,N_16522);
and UO_2459 (O_2459,N_17452,N_16632);
or UO_2460 (O_2460,N_19280,N_16793);
or UO_2461 (O_2461,N_18701,N_17673);
xnor UO_2462 (O_2462,N_16384,N_16209);
or UO_2463 (O_2463,N_18118,N_19644);
xnor UO_2464 (O_2464,N_18155,N_18929);
nand UO_2465 (O_2465,N_16017,N_16824);
xnor UO_2466 (O_2466,N_18536,N_17637);
nand UO_2467 (O_2467,N_17736,N_18669);
or UO_2468 (O_2468,N_17503,N_17787);
nand UO_2469 (O_2469,N_16620,N_18924);
xnor UO_2470 (O_2470,N_19833,N_18558);
and UO_2471 (O_2471,N_16744,N_19024);
nand UO_2472 (O_2472,N_16238,N_17971);
and UO_2473 (O_2473,N_17487,N_16502);
or UO_2474 (O_2474,N_17728,N_16825);
xnor UO_2475 (O_2475,N_19783,N_19040);
or UO_2476 (O_2476,N_16471,N_18122);
xnor UO_2477 (O_2477,N_16342,N_19713);
or UO_2478 (O_2478,N_18620,N_16450);
xor UO_2479 (O_2479,N_18219,N_19152);
nor UO_2480 (O_2480,N_17593,N_17321);
nor UO_2481 (O_2481,N_17030,N_16959);
and UO_2482 (O_2482,N_16957,N_18569);
or UO_2483 (O_2483,N_16416,N_17660);
nor UO_2484 (O_2484,N_18270,N_19227);
nor UO_2485 (O_2485,N_16166,N_18917);
xnor UO_2486 (O_2486,N_19312,N_16269);
nand UO_2487 (O_2487,N_19477,N_16724);
and UO_2488 (O_2488,N_19281,N_19198);
nor UO_2489 (O_2489,N_17374,N_16109);
nor UO_2490 (O_2490,N_18180,N_16497);
xnor UO_2491 (O_2491,N_19476,N_18246);
or UO_2492 (O_2492,N_18780,N_19904);
or UO_2493 (O_2493,N_17897,N_17189);
xnor UO_2494 (O_2494,N_17477,N_19650);
nor UO_2495 (O_2495,N_16381,N_19799);
or UO_2496 (O_2496,N_16867,N_17582);
xnor UO_2497 (O_2497,N_19861,N_18444);
nor UO_2498 (O_2498,N_19017,N_19209);
nor UO_2499 (O_2499,N_16010,N_19555);
endmodule